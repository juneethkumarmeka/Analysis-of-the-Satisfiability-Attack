module basic_2500_25000_3000_100_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
nand U0 (N_0,In_2478,In_869);
or U1 (N_1,In_2363,In_51);
nand U2 (N_2,In_1566,In_1558);
or U3 (N_3,In_2146,In_1503);
and U4 (N_4,In_850,In_749);
nor U5 (N_5,In_475,In_574);
xor U6 (N_6,In_1,In_2339);
xnor U7 (N_7,In_2380,In_2193);
xor U8 (N_8,In_1904,In_1509);
nand U9 (N_9,In_54,In_1237);
and U10 (N_10,In_569,In_1907);
xor U11 (N_11,In_201,In_317);
nand U12 (N_12,In_577,In_1268);
and U13 (N_13,In_2358,In_2004);
or U14 (N_14,In_163,In_623);
nand U15 (N_15,In_557,In_937);
nand U16 (N_16,In_810,In_2011);
nor U17 (N_17,In_2170,In_1931);
nand U18 (N_18,In_556,In_396);
xor U19 (N_19,In_1909,In_584);
or U20 (N_20,In_558,In_1598);
or U21 (N_21,In_1230,In_490);
and U22 (N_22,In_1589,In_2452);
nand U23 (N_23,In_1720,In_1660);
nor U24 (N_24,In_843,In_1078);
nand U25 (N_25,In_1400,In_478);
xnor U26 (N_26,In_1814,In_1073);
or U27 (N_27,In_2332,In_1471);
nor U28 (N_28,In_976,In_74);
nor U29 (N_29,In_1472,In_1447);
nand U30 (N_30,In_1187,In_2469);
nor U31 (N_31,In_2191,In_56);
or U32 (N_32,In_2364,In_637);
and U33 (N_33,In_1286,In_1012);
and U34 (N_34,In_708,In_667);
and U35 (N_35,In_2225,In_2054);
xor U36 (N_36,In_890,In_499);
nor U37 (N_37,In_412,In_1665);
and U38 (N_38,In_2185,In_1090);
or U39 (N_39,In_2323,In_1360);
nand U40 (N_40,In_150,In_2049);
and U41 (N_41,In_17,In_2474);
or U42 (N_42,In_2172,In_1853);
nand U43 (N_43,In_2485,In_709);
nand U44 (N_44,In_1719,In_564);
nand U45 (N_45,In_2127,In_1937);
nor U46 (N_46,In_189,In_1725);
and U47 (N_47,In_1065,In_818);
and U48 (N_48,In_315,In_756);
nand U49 (N_49,In_1809,In_1573);
or U50 (N_50,In_991,In_2247);
or U51 (N_51,In_1932,In_862);
or U52 (N_52,In_1748,In_1759);
or U53 (N_53,In_479,In_1109);
nand U54 (N_54,In_73,In_1161);
nor U55 (N_55,In_1269,In_665);
or U56 (N_56,In_1359,In_1403);
nand U57 (N_57,In_1704,In_318);
nand U58 (N_58,In_591,In_820);
or U59 (N_59,In_70,In_1765);
nor U60 (N_60,In_1977,In_449);
and U61 (N_61,In_1987,In_539);
xnor U62 (N_62,In_37,In_249);
nand U63 (N_63,In_887,In_1256);
nand U64 (N_64,In_901,In_2278);
xor U65 (N_65,In_1523,In_1584);
xor U66 (N_66,In_1140,In_1219);
xor U67 (N_67,In_870,In_715);
or U68 (N_68,In_1319,In_982);
and U69 (N_69,In_1167,In_83);
nand U70 (N_70,In_421,In_1839);
nor U71 (N_71,In_40,In_1114);
nor U72 (N_72,In_759,In_2436);
nand U73 (N_73,In_128,In_1204);
and U74 (N_74,In_302,In_2265);
or U75 (N_75,In_1735,In_1992);
nand U76 (N_76,In_1985,In_1887);
xnor U77 (N_77,In_1612,In_649);
or U78 (N_78,In_305,In_2166);
or U79 (N_79,In_2472,In_2309);
and U80 (N_80,In_751,In_536);
nand U81 (N_81,In_1976,In_491);
and U82 (N_82,In_214,In_130);
nand U83 (N_83,In_778,In_1934);
nand U84 (N_84,In_774,In_2388);
nand U85 (N_85,In_394,In_1636);
or U86 (N_86,In_2280,In_95);
nor U87 (N_87,In_388,In_1724);
or U88 (N_88,In_198,In_1994);
or U89 (N_89,In_959,In_1946);
nand U90 (N_90,In_180,In_2184);
xnor U91 (N_91,In_2200,In_97);
xnor U92 (N_92,In_1036,In_1231);
nand U93 (N_93,In_1241,In_1867);
nor U94 (N_94,In_2208,In_2121);
nor U95 (N_95,In_808,In_393);
nor U96 (N_96,In_1914,In_96);
or U97 (N_97,In_1832,In_2350);
and U98 (N_98,In_213,In_2490);
nor U99 (N_99,In_866,In_2284);
xor U100 (N_100,In_1440,In_469);
nor U101 (N_101,In_607,In_1702);
and U102 (N_102,In_1410,In_670);
nor U103 (N_103,In_178,In_2091);
xnor U104 (N_104,In_2017,In_793);
or U105 (N_105,In_1479,In_1613);
xor U106 (N_106,In_790,In_11);
xor U107 (N_107,In_691,In_831);
nand U108 (N_108,In_1182,In_171);
nor U109 (N_109,In_1330,In_1189);
nor U110 (N_110,In_1718,In_1142);
or U111 (N_111,In_2105,In_605);
and U112 (N_112,In_1708,In_68);
or U113 (N_113,In_1491,In_237);
xor U114 (N_114,In_983,In_158);
or U115 (N_115,In_1557,In_1654);
or U116 (N_116,In_2095,In_1437);
nor U117 (N_117,In_1647,In_521);
or U118 (N_118,In_1006,In_616);
nor U119 (N_119,In_1138,In_878);
nand U120 (N_120,In_2142,In_1101);
or U121 (N_121,In_1004,In_1877);
nor U122 (N_122,In_100,In_2032);
and U123 (N_123,In_63,In_1037);
xnor U124 (N_124,In_739,In_524);
nand U125 (N_125,In_1155,In_1973);
or U126 (N_126,In_1068,In_60);
nor U127 (N_127,In_1502,In_1644);
nor U128 (N_128,In_1171,In_608);
nor U129 (N_129,In_1295,In_1056);
and U130 (N_130,In_1574,In_1726);
nor U131 (N_131,In_265,In_132);
and U132 (N_132,In_207,In_1981);
nand U133 (N_133,In_657,In_441);
xor U134 (N_134,In_1944,In_1581);
and U135 (N_135,In_142,In_534);
nand U136 (N_136,In_2356,In_2186);
and U137 (N_137,In_471,In_2212);
and U138 (N_138,In_1760,In_2286);
nand U139 (N_139,In_826,In_66);
xor U140 (N_140,In_10,In_2051);
nand U141 (N_141,In_1422,In_1250);
nor U142 (N_142,In_529,In_1721);
nand U143 (N_143,In_1104,In_2366);
and U144 (N_144,In_1420,In_1924);
xor U145 (N_145,In_2390,In_543);
and U146 (N_146,In_281,In_155);
nor U147 (N_147,In_755,In_275);
and U148 (N_148,In_1482,In_1692);
xnor U149 (N_149,In_382,In_138);
xnor U150 (N_150,In_2048,In_635);
or U151 (N_151,In_477,In_1510);
nand U152 (N_152,In_1605,In_190);
nand U153 (N_153,In_1465,In_1080);
nand U154 (N_154,In_466,In_512);
nor U155 (N_155,In_955,In_1445);
or U156 (N_156,In_1433,In_410);
nand U157 (N_157,In_414,In_447);
xnor U158 (N_158,In_392,In_1274);
nand U159 (N_159,In_234,In_1102);
nand U160 (N_160,In_294,In_2113);
and U161 (N_161,In_2025,In_2440);
xnor U162 (N_162,In_2168,In_485);
or U163 (N_163,In_398,In_1648);
nor U164 (N_164,In_596,In_288);
and U165 (N_165,In_454,In_1733);
nor U166 (N_166,In_404,In_2458);
nand U167 (N_167,In_2376,In_1087);
nor U168 (N_168,In_1556,In_1333);
or U169 (N_169,In_1264,In_2112);
xnor U170 (N_170,In_2345,In_659);
or U171 (N_171,In_2318,In_2209);
and U172 (N_172,In_359,In_2169);
or U173 (N_173,In_600,In_99);
and U174 (N_174,In_1882,In_687);
nand U175 (N_175,In_886,In_1480);
or U176 (N_176,In_450,In_1788);
and U177 (N_177,In_2154,In_1808);
nand U178 (N_178,In_1508,In_2279);
or U179 (N_179,In_719,In_496);
nand U180 (N_180,In_1632,In_2241);
and U181 (N_181,In_2438,In_1857);
nor U182 (N_182,In_1134,In_2414);
nor U183 (N_183,In_1300,In_1528);
nand U184 (N_184,In_2373,In_1540);
nand U185 (N_185,In_1011,In_1031);
nor U186 (N_186,In_2374,In_2282);
xor U187 (N_187,In_409,In_323);
nor U188 (N_188,In_758,In_2214);
and U189 (N_189,In_1880,In_1982);
xnor U190 (N_190,In_763,In_2306);
or U191 (N_191,In_996,In_2258);
and U192 (N_192,In_2470,In_241);
or U193 (N_193,In_2274,In_645);
xor U194 (N_194,In_1616,In_2220);
xor U195 (N_195,In_453,In_2281);
xnor U196 (N_196,In_62,In_990);
or U197 (N_197,In_981,In_1916);
nor U198 (N_198,In_986,In_1940);
nor U199 (N_199,In_2013,In_1734);
xnor U200 (N_200,In_1792,In_1892);
nor U201 (N_201,In_1336,In_892);
or U202 (N_202,In_979,In_2068);
or U203 (N_203,In_1969,In_695);
nand U204 (N_204,In_278,In_916);
nor U205 (N_205,In_231,In_2222);
or U206 (N_206,In_1518,In_854);
nand U207 (N_207,In_1507,In_333);
or U208 (N_208,In_2368,In_2346);
nand U209 (N_209,In_1213,In_1545);
nand U210 (N_210,In_2404,In_978);
nor U211 (N_211,In_295,In_1257);
xor U212 (N_212,In_296,In_2125);
xor U213 (N_213,In_112,In_788);
and U214 (N_214,In_2389,In_434);
nand U215 (N_215,In_2211,In_1374);
and U216 (N_216,In_837,In_1623);
nand U217 (N_217,In_357,In_2114);
nor U218 (N_218,In_140,In_134);
xor U219 (N_219,In_773,In_517);
or U220 (N_220,In_1630,In_2322);
and U221 (N_221,In_2023,In_2147);
nand U222 (N_222,In_1381,In_1035);
nand U223 (N_223,In_1675,In_290);
or U224 (N_224,In_2256,In_2045);
xor U225 (N_225,In_1930,In_1520);
or U226 (N_226,In_841,In_1607);
nor U227 (N_227,In_965,In_1332);
xnor U228 (N_228,In_1239,In_125);
nand U229 (N_229,In_331,In_1772);
and U230 (N_230,In_436,In_1764);
or U231 (N_231,In_1337,In_1975);
nand U232 (N_232,In_971,In_1423);
xnor U233 (N_233,In_697,In_85);
or U234 (N_234,In_1628,In_1272);
nand U235 (N_235,In_1150,In_1267);
nor U236 (N_236,In_585,In_2161);
xor U237 (N_237,In_1711,In_643);
xor U238 (N_238,In_1145,In_1293);
nor U239 (N_239,In_2443,In_2480);
nor U240 (N_240,In_121,In_2029);
nand U241 (N_241,In_219,In_1048);
nor U242 (N_242,In_2402,In_67);
or U243 (N_243,In_1835,In_1417);
nand U244 (N_244,In_170,In_2198);
and U245 (N_245,In_304,In_2295);
and U246 (N_246,In_1024,In_2031);
xor U247 (N_247,In_771,In_1536);
nand U248 (N_248,In_1798,In_379);
and U249 (N_249,In_444,In_1296);
and U250 (N_250,In_1008,In_606);
or U251 (N_251,In_849,In_2109);
nand U252 (N_252,In_350,In_1081);
and U253 (N_253,In_1836,In_2027);
nor U254 (N_254,In_2075,In_2255);
and U255 (N_255,In_2,In_1871);
xor U256 (N_256,In_1326,In_277);
xnor U257 (N_257,In_2233,In_1678);
nor U258 (N_258,In_2468,In_2341);
and U259 (N_259,In_2344,N_184);
or U260 (N_260,In_1587,In_2412);
nand U261 (N_261,In_1959,In_511);
nor U262 (N_262,In_1478,In_1179);
or U263 (N_263,In_86,In_386);
and U264 (N_264,In_1232,In_1637);
and U265 (N_265,N_52,In_1328);
and U266 (N_266,N_108,In_356);
xnor U267 (N_267,In_1668,In_897);
nand U268 (N_268,In_930,In_527);
nor U269 (N_269,In_2300,In_384);
xnor U270 (N_270,N_35,In_615);
nand U271 (N_271,In_1752,In_1365);
xnor U272 (N_272,In_1045,In_2488);
or U273 (N_273,In_1898,In_1986);
xor U274 (N_274,In_151,In_133);
nand U275 (N_275,In_1289,In_238);
nor U276 (N_276,In_2174,In_452);
nor U277 (N_277,In_507,In_2144);
and U278 (N_278,In_2021,In_2329);
nor U279 (N_279,In_914,N_238);
and U280 (N_280,In_126,In_334);
or U281 (N_281,In_1622,In_1217);
and U282 (N_282,In_933,In_860);
or U283 (N_283,In_1758,In_680);
nor U284 (N_284,In_924,In_1355);
and U285 (N_285,In_13,In_631);
or U286 (N_286,In_1271,In_2403);
and U287 (N_287,In_2081,In_1072);
or U288 (N_288,N_242,In_1196);
nor U289 (N_289,In_119,In_614);
and U290 (N_290,In_1162,In_1818);
and U291 (N_291,N_188,In_1354);
nor U292 (N_292,In_1136,In_169);
nand U293 (N_293,In_2087,In_1164);
nand U294 (N_294,In_1228,In_272);
and U295 (N_295,In_1304,In_2423);
xor U296 (N_296,In_1902,In_194);
or U297 (N_297,In_953,N_115);
nand U298 (N_298,In_791,N_90);
and U299 (N_299,In_1497,In_242);
and U300 (N_300,In_2044,In_1694);
nand U301 (N_301,In_1099,In_2413);
nor U302 (N_302,In_424,In_1310);
xnor U303 (N_303,In_338,In_1691);
xor U304 (N_304,In_2242,In_1338);
or U305 (N_305,In_1461,In_256);
or U306 (N_306,In_830,In_989);
nor U307 (N_307,In_2289,In_1383);
xor U308 (N_308,In_2024,In_704);
nand U309 (N_309,In_28,In_291);
xnor U310 (N_310,In_2287,In_1125);
nor U311 (N_311,N_162,In_1156);
or U312 (N_312,In_2427,In_1340);
and U313 (N_313,In_2138,In_191);
and U314 (N_314,In_319,In_1989);
xor U315 (N_315,In_813,N_190);
and U316 (N_316,In_1178,In_613);
xor U317 (N_317,In_640,In_1192);
or U318 (N_318,N_237,In_1091);
xnor U319 (N_319,In_619,In_1797);
and U320 (N_320,N_221,In_825);
or U321 (N_321,In_941,In_1816);
or U322 (N_322,N_197,In_355);
or U323 (N_323,In_1493,In_2386);
nor U324 (N_324,In_2076,In_1190);
and U325 (N_325,In_16,In_1591);
nor U326 (N_326,In_34,N_215);
or U327 (N_327,In_2426,In_710);
xor U328 (N_328,N_5,In_1077);
nand U329 (N_329,N_39,In_202);
or U330 (N_330,In_1728,In_1784);
and U331 (N_331,In_852,In_1917);
xnor U332 (N_332,In_2057,In_815);
or U333 (N_333,In_271,In_1103);
or U334 (N_334,In_1253,In_2003);
nand U335 (N_335,In_1018,In_2418);
and U336 (N_336,In_1639,In_224);
or U337 (N_337,In_1195,In_124);
nor U338 (N_338,In_2206,In_1657);
nand U339 (N_339,In_1224,In_2001);
nand U340 (N_340,In_737,In_2179);
or U341 (N_341,In_590,In_1499);
nor U342 (N_342,In_2082,In_2262);
or U343 (N_343,In_27,In_1896);
and U344 (N_344,In_806,In_1999);
and U345 (N_345,In_1496,In_280);
or U346 (N_346,In_373,N_138);
or U347 (N_347,In_1525,In_728);
nand U348 (N_348,In_2123,In_904);
nor U349 (N_349,In_2463,In_1655);
xnor U350 (N_350,In_1830,In_362);
xor U351 (N_351,In_2006,In_1893);
and U352 (N_352,In_2464,In_2187);
and U353 (N_353,In_836,In_1088);
or U354 (N_354,In_839,In_1597);
nor U355 (N_355,In_1667,In_786);
and U356 (N_356,In_1700,N_148);
xnor U357 (N_357,In_420,In_2271);
nand U358 (N_358,In_1848,In_2159);
or U359 (N_359,In_977,In_153);
nor U360 (N_360,In_53,In_2498);
nand U361 (N_361,In_429,In_1512);
nand U362 (N_362,In_805,In_1876);
nor U363 (N_363,In_1463,In_2064);
nor U364 (N_364,N_118,In_555);
nor U365 (N_365,N_239,In_1534);
xor U366 (N_366,In_423,In_248);
xor U367 (N_367,In_2145,In_1351);
nand U368 (N_368,N_105,In_566);
nor U369 (N_369,In_2367,In_1858);
nor U370 (N_370,In_993,N_172);
or U371 (N_371,In_395,In_1677);
nor U372 (N_372,In_2340,In_2007);
or U373 (N_373,In_1550,In_1869);
nand U374 (N_374,In_2129,In_2157);
xor U375 (N_375,In_1137,In_724);
nand U376 (N_376,In_612,In_1375);
or U377 (N_377,In_369,In_1292);
nor U378 (N_378,In_2108,In_1922);
and U379 (N_379,In_1823,In_1096);
nand U380 (N_380,In_243,N_186);
or U381 (N_381,In_208,N_211);
nand U382 (N_382,In_293,N_24);
and U383 (N_383,In_2182,In_209);
nand U384 (N_384,In_1915,In_2425);
xnor U385 (N_385,In_1070,In_467);
and U386 (N_386,In_2450,In_2387);
nand U387 (N_387,In_1113,In_1427);
or U388 (N_388,In_1385,In_1026);
nand U389 (N_389,In_1131,In_1448);
nor U390 (N_390,N_116,In_2334);
nor U391 (N_391,In_538,In_1276);
nor U392 (N_392,In_2448,In_1756);
or U393 (N_393,In_954,In_223);
and U394 (N_394,In_948,In_2128);
or U395 (N_395,In_1817,N_227);
nor U396 (N_396,In_1277,In_668);
or U397 (N_397,N_65,In_1701);
nand U398 (N_398,In_1742,N_246);
nor U399 (N_399,In_1970,N_192);
xnor U400 (N_400,In_2477,In_1363);
nor U401 (N_401,In_1707,In_1266);
and U402 (N_402,In_729,In_1543);
or U403 (N_403,In_1686,In_1933);
and U404 (N_404,In_225,In_1886);
or U405 (N_405,In_1949,In_671);
and U406 (N_406,In_935,In_1601);
nor U407 (N_407,In_840,In_995);
nand U408 (N_408,In_722,In_2041);
nor U409 (N_409,In_1233,In_1527);
xnor U410 (N_410,In_1392,In_1910);
nor U411 (N_411,In_1430,In_1789);
xor U412 (N_412,N_111,In_1715);
nor U413 (N_413,In_1172,In_1066);
nand U414 (N_414,In_2089,In_1373);
or U415 (N_415,In_713,N_174);
and U416 (N_416,In_928,In_1653);
xnor U417 (N_417,In_921,In_65);
nand U418 (N_418,In_405,In_164);
nor U419 (N_419,In_972,N_95);
and U420 (N_420,In_655,In_365);
nand U421 (N_421,In_1820,In_675);
and U422 (N_422,In_1807,In_1058);
xnor U423 (N_423,In_274,In_797);
xnor U424 (N_424,In_1649,In_515);
or U425 (N_425,In_1315,In_459);
nand U426 (N_426,In_1846,In_1954);
nand U427 (N_427,In_23,In_21);
nor U428 (N_428,In_1442,In_1827);
and U429 (N_429,In_32,In_1082);
or U430 (N_430,In_1242,In_2415);
xnor U431 (N_431,N_69,In_663);
or U432 (N_432,In_641,N_230);
nand U433 (N_433,In_1569,In_523);
or U434 (N_434,In_1390,In_1919);
nand U435 (N_435,N_34,In_2400);
and U436 (N_436,N_3,N_241);
xor U437 (N_437,In_1317,In_216);
nor U438 (N_438,In_525,In_2092);
xor U439 (N_439,In_2139,N_201);
nand U440 (N_440,In_2457,In_1438);
nor U441 (N_441,In_910,In_102);
or U442 (N_442,In_1851,In_162);
or U443 (N_443,In_2397,In_266);
xnor U444 (N_444,In_1439,In_1565);
or U445 (N_445,In_1731,N_129);
and U446 (N_446,In_332,In_879);
nand U447 (N_447,In_1100,In_2176);
nor U448 (N_448,In_537,In_1019);
nand U449 (N_449,N_178,In_2487);
and U450 (N_450,In_1248,In_464);
nand U451 (N_451,In_787,In_642);
and U452 (N_452,In_123,In_1169);
nand U453 (N_453,In_1663,In_1918);
nand U454 (N_454,In_1819,In_1111);
or U455 (N_455,In_2351,N_71);
or U456 (N_456,In_1806,In_1779);
and U457 (N_457,In_1469,In_1378);
nand U458 (N_458,In_519,In_1316);
or U459 (N_459,N_8,In_970);
or U460 (N_460,In_1768,In_1651);
or U461 (N_461,In_915,In_514);
and U462 (N_462,In_385,N_79);
and U463 (N_463,N_123,In_1168);
or U464 (N_464,In_2201,In_1582);
nor U465 (N_465,N_66,In_1229);
and U466 (N_466,In_1530,N_214);
or U467 (N_467,In_835,In_1038);
nor U468 (N_468,In_431,In_44);
nand U469 (N_469,In_2078,In_1216);
and U470 (N_470,In_572,In_1221);
and U471 (N_471,In_211,In_681);
xnor U472 (N_472,In_316,In_2355);
nand U473 (N_473,In_1732,In_312);
xnor U474 (N_474,In_765,N_53);
or U475 (N_475,In_1034,In_1098);
xor U476 (N_476,In_792,N_74);
nor U477 (N_477,In_313,In_2202);
or U478 (N_478,In_1791,In_2009);
and U479 (N_479,In_2014,In_378);
and U480 (N_480,In_1255,N_125);
nand U481 (N_481,In_1766,In_87);
nor U482 (N_482,N_206,In_1388);
and U483 (N_483,In_2194,In_1382);
xnor U484 (N_484,In_1901,In_1243);
and U485 (N_485,In_1952,In_2455);
nand U486 (N_486,In_301,In_1926);
xor U487 (N_487,In_336,In_310);
and U488 (N_488,N_126,In_2093);
nor U489 (N_489,In_1214,In_812);
xor U490 (N_490,In_1174,In_578);
and U491 (N_491,In_958,In_1855);
or U492 (N_492,In_799,In_361);
or U493 (N_493,In_1425,N_85);
nand U494 (N_494,In_817,In_401);
or U495 (N_495,In_530,In_1906);
nand U496 (N_496,In_480,In_2126);
or U497 (N_497,In_602,In_2462);
xnor U498 (N_498,In_1312,In_859);
or U499 (N_499,In_846,In_458);
and U500 (N_500,In_1370,In_78);
xor U501 (N_501,In_2084,N_497);
or U502 (N_502,In_1435,In_1135);
and U503 (N_503,In_1025,In_349);
nand U504 (N_504,N_20,N_328);
or U505 (N_505,In_2038,In_2270);
nor U506 (N_506,In_533,In_1712);
or U507 (N_507,In_803,In_82);
xor U508 (N_508,In_780,In_1297);
and U509 (N_509,In_2328,In_116);
nor U510 (N_510,In_2035,N_119);
or U511 (N_511,N_75,In_565);
nand U512 (N_512,In_45,In_1866);
xnor U513 (N_513,N_360,In_366);
or U514 (N_514,In_2330,In_1258);
or U515 (N_515,In_1629,In_1457);
nand U516 (N_516,In_1996,In_1652);
nor U517 (N_517,In_1181,In_2034);
nand U518 (N_518,In_1662,In_516);
and U519 (N_519,In_617,In_2324);
xnor U520 (N_520,N_399,In_2132);
xor U521 (N_521,N_314,In_625);
nand U522 (N_522,In_822,In_1318);
nand U523 (N_523,In_907,In_1003);
and U524 (N_524,In_1210,N_351);
xnor U525 (N_525,In_283,N_391);
or U526 (N_526,N_309,In_206);
nand U527 (N_527,In_1881,In_1202);
nor U528 (N_528,In_1962,In_1927);
xnor U529 (N_529,In_1251,In_15);
or U530 (N_530,In_662,In_1621);
or U531 (N_531,In_1804,N_175);
or U532 (N_532,In_2476,In_1695);
or U533 (N_533,In_2232,In_1245);
and U534 (N_534,In_2088,N_251);
and U535 (N_535,In_2310,In_1331);
xnor U536 (N_536,In_2365,In_2055);
nand U537 (N_537,N_357,In_2028);
nand U538 (N_538,In_199,In_2395);
and U539 (N_539,In_1001,In_416);
nor U540 (N_540,N_14,In_1209);
nand U541 (N_541,In_513,In_204);
and U542 (N_542,In_1722,In_2473);
nand U543 (N_543,In_250,N_291);
and U544 (N_544,N_410,In_1419);
xor U545 (N_545,In_1366,In_1782);
or U546 (N_546,N_473,N_367);
and U547 (N_547,N_370,In_1929);
xor U548 (N_548,N_340,In_147);
nor U549 (N_549,In_347,In_1737);
nand U550 (N_550,In_2337,N_18);
nor U551 (N_551,In_2177,In_1234);
or U552 (N_552,N_216,N_67);
xor U553 (N_553,In_648,In_743);
xor U554 (N_554,In_1555,In_750);
xnor U555 (N_555,N_139,In_196);
xor U556 (N_556,In_828,In_2251);
and U557 (N_557,N_428,In_483);
xnor U558 (N_558,In_898,In_2417);
xor U559 (N_559,N_350,In_961);
nand U560 (N_560,In_1021,In_227);
and U561 (N_561,In_1394,In_1413);
xnor U562 (N_562,In_2012,In_2040);
and U563 (N_563,In_2276,In_744);
nor U564 (N_564,N_416,In_1222);
and U565 (N_565,N_471,In_2033);
and U566 (N_566,N_312,In_876);
xor U567 (N_567,N_305,In_1751);
or U568 (N_568,In_2444,In_55);
nor U569 (N_569,N_440,In_1452);
nand U570 (N_570,In_639,In_36);
nand U571 (N_571,In_1495,In_1801);
xnor U572 (N_572,In_1280,N_277);
xnor U573 (N_573,In_270,In_285);
and U574 (N_574,N_465,In_72);
and U575 (N_575,In_2430,In_2333);
or U576 (N_576,N_398,N_414);
and U577 (N_577,In_108,N_245);
or U578 (N_578,In_923,N_341);
nand U579 (N_579,In_1710,In_2460);
and U580 (N_580,In_1713,In_1047);
nor U581 (N_581,In_98,N_493);
xnor U582 (N_582,In_1714,In_2424);
xnor U583 (N_583,In_919,In_769);
nor U584 (N_584,N_265,In_320);
or U585 (N_585,In_1016,In_573);
or U586 (N_586,In_422,In_807);
and U587 (N_587,In_652,In_2396);
nor U588 (N_588,In_936,In_1041);
and U589 (N_589,In_1455,In_1158);
nand U590 (N_590,In_149,In_1864);
xnor U591 (N_591,In_1467,In_2090);
and U592 (N_592,In_166,In_1468);
or U593 (N_593,In_1307,In_845);
nor U594 (N_594,In_322,In_811);
or U595 (N_595,In_2319,In_946);
nor U596 (N_596,In_762,N_110);
and U597 (N_597,In_1415,In_2459);
or U598 (N_598,N_259,In_968);
nand U599 (N_599,N_262,In_120);
or U600 (N_600,In_258,In_856);
xnor U601 (N_601,In_2171,In_800);
xor U602 (N_602,In_183,In_802);
xnor U603 (N_603,In_2316,In_727);
nor U604 (N_604,In_1859,In_1030);
or U605 (N_605,In_205,In_2297);
or U606 (N_606,In_348,In_2204);
and U607 (N_607,In_252,In_908);
nand U608 (N_608,In_541,In_1826);
nand U609 (N_609,In_1407,In_1885);
or U610 (N_610,N_22,In_1746);
and U611 (N_611,In_809,N_356);
nand U612 (N_612,N_250,In_1854);
and U613 (N_613,In_1118,N_157);
xnor U614 (N_614,N_161,N_210);
nand U615 (N_615,In_1399,In_1097);
nand U616 (N_616,In_2349,In_1744);
nand U617 (N_617,In_1615,In_1335);
and U618 (N_618,N_136,In_920);
nand U619 (N_619,In_2118,N_273);
nand U620 (N_620,In_1339,In_35);
and U621 (N_621,N_483,In_2435);
or U622 (N_622,In_2362,N_33);
nand U623 (N_623,In_403,In_1603);
and U624 (N_624,In_1444,N_293);
xnor U625 (N_625,In_1046,In_2314);
nand U626 (N_626,In_1320,N_423);
nor U627 (N_627,In_604,In_716);
nor U628 (N_628,In_1769,In_1620);
and U629 (N_629,In_1112,N_13);
nand U630 (N_630,In_903,In_2197);
nor U631 (N_631,In_1506,In_609);
or U632 (N_632,In_1180,N_431);
nand U633 (N_633,In_2060,In_2348);
or U634 (N_634,In_844,In_2454);
and U635 (N_635,In_1429,In_335);
xnor U636 (N_636,In_428,In_442);
and U637 (N_637,N_92,In_913);
nor U638 (N_638,In_186,N_49);
nand U639 (N_639,In_2313,In_900);
nand U640 (N_640,In_2010,In_706);
nand U641 (N_641,N_427,In_71);
nand U642 (N_642,In_611,In_1165);
nand U643 (N_643,In_254,N_420);
and U644 (N_644,In_618,In_2305);
nor U645 (N_645,N_317,In_863);
or U646 (N_646,In_1050,In_711);
or U647 (N_647,In_284,N_217);
and U648 (N_648,N_443,In_650);
xnor U649 (N_649,N_320,In_1093);
nor U650 (N_650,In_1567,In_554);
nand U651 (N_651,In_474,In_1094);
nand U652 (N_652,In_381,In_2016);
nand U653 (N_653,In_3,N_469);
or U654 (N_654,In_2065,In_1634);
nor U655 (N_655,N_229,In_1578);
and U656 (N_656,N_283,In_1757);
nand U657 (N_657,In_1522,In_24);
xnor U658 (N_658,In_167,N_359);
and U659 (N_659,N_375,In_1055);
and U660 (N_660,In_1284,In_505);
or U661 (N_661,In_1958,N_487);
or U662 (N_662,In_251,In_1747);
and U663 (N_663,In_1369,In_372);
nand U664 (N_664,In_210,N_382);
xor U665 (N_665,In_1993,In_2335);
nor U666 (N_666,N_441,In_1750);
xor U667 (N_667,In_2331,In_417);
xnor U668 (N_668,In_1755,N_476);
nor U669 (N_669,In_33,In_1703);
or U670 (N_670,In_1197,In_1485);
and U671 (N_671,N_271,In_712);
or U672 (N_672,In_1013,In_1456);
xnor U673 (N_673,In_1128,N_103);
or U674 (N_674,N_321,N_372);
or U675 (N_675,N_422,N_218);
nand U676 (N_676,In_1560,In_1998);
nor U677 (N_677,N_47,In_2261);
or U678 (N_678,N_308,In_2231);
or U679 (N_679,In_1261,In_526);
or U680 (N_680,In_1729,N_352);
nor U681 (N_681,In_2369,In_465);
nand U682 (N_682,In_2115,In_1515);
nand U683 (N_683,In_1017,In_875);
or U684 (N_684,In_2210,In_1436);
nor U685 (N_685,In_2293,In_580);
nor U686 (N_686,In_1865,In_1843);
nor U687 (N_687,In_1529,In_664);
or U688 (N_688,N_87,In_1658);
nor U689 (N_689,In_2327,In_1398);
and U690 (N_690,In_2224,N_289);
xor U691 (N_691,In_1120,In_1965);
or U692 (N_692,N_297,In_535);
xnor U693 (N_693,In_2098,In_1585);
nor U694 (N_694,In_1551,In_2236);
nand U695 (N_695,In_1043,In_377);
and U696 (N_696,In_783,In_2456);
nand U697 (N_697,In_161,In_592);
and U698 (N_698,N_302,In_798);
xor U699 (N_699,In_597,In_1738);
or U700 (N_700,In_804,N_209);
and U701 (N_701,In_647,In_882);
nand U702 (N_702,N_330,N_269);
xor U703 (N_703,N_54,In_371);
or U704 (N_704,In_430,In_456);
or U705 (N_705,In_877,In_1441);
nor U706 (N_706,In_1201,In_1563);
xnor U707 (N_707,In_1611,In_1803);
xnor U708 (N_708,In_1022,In_2252);
xnor U709 (N_709,In_2370,N_156);
or U710 (N_710,In_2283,In_157);
and U711 (N_711,In_939,N_109);
nand U712 (N_712,N_279,N_248);
xnor U713 (N_713,In_563,In_766);
and U714 (N_714,N_28,N_484);
nand U715 (N_715,In_628,In_1541);
or U716 (N_716,N_147,N_355);
xnor U717 (N_717,In_966,In_181);
and U718 (N_718,In_1207,In_2240);
nand U719 (N_719,In_2077,In_343);
or U720 (N_720,In_666,In_2493);
or U721 (N_721,N_329,In_2219);
nand U722 (N_722,In_2361,In_684);
nor U723 (N_723,In_38,In_353);
and U724 (N_724,N_73,N_41);
and U725 (N_725,In_1028,In_31);
and U726 (N_726,In_1314,In_2353);
nor U727 (N_727,N_433,N_258);
nor U728 (N_728,In_2285,In_1428);
or U729 (N_729,In_1531,In_247);
nand U730 (N_730,In_1535,In_1626);
nand U731 (N_731,In_2047,In_693);
and U732 (N_732,In_1849,In_857);
nor U733 (N_733,In_2149,In_2239);
nor U734 (N_734,In_1343,N_72);
xnor U735 (N_735,N_371,N_385);
nor U736 (N_736,N_267,In_1938);
xor U737 (N_737,N_429,In_1576);
xnor U738 (N_738,In_1200,In_952);
nand U739 (N_739,In_25,N_80);
or U740 (N_740,In_1872,In_2158);
and U741 (N_741,In_2183,In_1874);
nand U742 (N_742,In_79,In_1313);
xnor U743 (N_743,N_120,N_358);
nand U744 (N_744,In_1347,In_1309);
and U745 (N_745,N_145,In_1199);
xnor U746 (N_746,In_145,N_389);
nand U747 (N_747,In_1119,In_20);
xnor U748 (N_748,N_386,N_62);
nand U749 (N_749,In_1380,In_2133);
xnor U750 (N_750,In_374,In_2453);
and U751 (N_751,N_78,N_45);
or U752 (N_752,In_1595,In_823);
or U753 (N_753,In_1602,N_364);
or U754 (N_754,N_491,N_623);
nand U755 (N_755,N_529,N_582);
and U756 (N_756,In_2384,N_96);
or U757 (N_757,N_586,In_1811);
nor U758 (N_758,In_437,In_2015);
nor U759 (N_759,In_2431,In_212);
nor U760 (N_760,In_630,In_2165);
and U761 (N_761,N_10,N_228);
nor U762 (N_762,In_1526,In_1943);
nand U763 (N_763,N_635,N_58);
xor U764 (N_764,In_2491,N_524);
xnor U765 (N_765,In_929,In_1840);
nand U766 (N_766,In_638,N_51);
or U767 (N_767,N_518,In_1740);
or U768 (N_768,N_101,In_508);
nand U769 (N_769,N_442,In_1489);
or U770 (N_770,N_527,In_984);
or U771 (N_771,N_739,In_2215);
and U772 (N_772,N_12,In_909);
and U773 (N_773,N_628,N_368);
or U774 (N_774,In_1641,N_622);
nand U775 (N_775,N_697,In_103);
xor U776 (N_776,In_177,In_1481);
and U777 (N_777,In_1484,In_1888);
and U778 (N_778,N_736,N_601);
nor U779 (N_779,In_30,N_30);
and U780 (N_780,In_101,In_1810);
and U781 (N_781,In_2441,N_453);
nand U782 (N_782,N_226,N_369);
xor U783 (N_783,In_726,In_732);
nor U784 (N_784,In_1060,N_354);
xor U785 (N_785,In_2140,N_573);
xnor U786 (N_786,N_597,N_616);
and U787 (N_787,In_1223,In_1847);
xor U788 (N_788,In_380,In_1588);
nand U789 (N_789,N_603,In_375);
xor U790 (N_790,In_1762,N_97);
nand U791 (N_791,In_314,N_337);
nor U792 (N_792,In_1492,In_2227);
nand U793 (N_793,N_725,In_2303);
or U794 (N_794,In_1014,In_2486);
or U795 (N_795,In_796,In_1575);
nor U796 (N_796,N_629,N_32);
nand U797 (N_797,In_76,In_7);
xnor U798 (N_798,In_1583,N_208);
nor U799 (N_799,In_917,In_2205);
or U800 (N_800,N_652,N_159);
or U801 (N_801,N_496,In_327);
or U802 (N_802,In_784,In_2238);
and U803 (N_803,N_749,N_553);
and U804 (N_804,In_337,N_198);
xor U805 (N_805,In_1083,N_160);
nor U806 (N_806,In_1990,In_2495);
or U807 (N_807,In_300,In_889);
nand U808 (N_808,In_1727,N_574);
and U809 (N_809,In_2073,In_733);
and U810 (N_810,In_2475,N_706);
and U811 (N_811,In_776,In_692);
nor U812 (N_812,In_1614,In_1948);
xor U813 (N_813,In_998,N_84);
nand U814 (N_814,In_775,In_1521);
nand U815 (N_815,In_1379,In_1913);
and U816 (N_816,In_752,In_1608);
nor U817 (N_817,In_1776,N_68);
or U818 (N_818,N_632,N_104);
nor U819 (N_819,In_506,In_218);
nor U820 (N_820,In_139,In_1116);
nor U821 (N_821,N_560,In_1693);
nand U822 (N_822,N_135,N_82);
nor U823 (N_823,N_55,In_2226);
nor U824 (N_824,In_240,In_1105);
and U825 (N_825,In_1329,N_280);
and U826 (N_826,N_155,N_114);
or U827 (N_827,In_1263,In_1771);
nand U828 (N_828,In_2381,N_298);
nand U829 (N_829,In_1084,In_861);
nor U830 (N_830,In_2137,In_1236);
xor U831 (N_831,N_438,N_718);
nand U832 (N_832,In_1829,In_1322);
nor U833 (N_833,N_282,N_704);
and U834 (N_834,N_322,In_351);
nor U835 (N_835,In_2002,N_687);
or U836 (N_836,In_1544,In_1879);
nand U837 (N_837,In_88,In_880);
xor U838 (N_838,N_479,In_951);
or U839 (N_839,N_505,N_510);
and U840 (N_840,N_439,In_2342);
xor U841 (N_841,N_133,In_899);
xnor U842 (N_842,In_1153,In_2189);
and U843 (N_843,In_906,N_381);
xnor U844 (N_844,In_997,In_1580);
or U845 (N_845,In_193,In_432);
or U846 (N_846,N_183,In_1203);
nand U847 (N_847,N_464,In_1273);
nand U848 (N_848,In_2026,In_172);
and U849 (N_849,In_896,In_2234);
nand U850 (N_850,In_2086,N_673);
xnor U851 (N_851,In_2235,N_475);
and U852 (N_852,In_451,N_694);
xor U853 (N_853,In_1281,In_545);
and U854 (N_854,N_686,In_768);
nor U855 (N_855,In_2074,N_36);
and U856 (N_856,In_131,In_731);
and U857 (N_857,In_1815,N_538);
and U858 (N_858,In_397,N_633);
nand U859 (N_859,N_252,N_285);
and U860 (N_860,In_884,N_685);
nor U861 (N_861,In_1953,N_301);
nor U862 (N_862,In_2447,N_182);
xor U863 (N_863,N_677,N_418);
and U864 (N_864,In_1795,In_1283);
or U865 (N_865,N_402,In_255);
nor U866 (N_866,In_286,In_1064);
and U867 (N_867,N_490,In_1838);
and U868 (N_868,N_383,In_470);
nor U869 (N_869,N_703,N_223);
and U870 (N_870,In_1571,In_1015);
nor U871 (N_871,N_268,In_891);
nor U872 (N_872,In_1773,In_203);
nor U873 (N_873,In_1126,In_1443);
nand U874 (N_874,In_1173,In_938);
or U875 (N_875,In_1144,In_2484);
and U876 (N_876,In_705,In_2378);
and U877 (N_877,In_2408,In_1303);
xnor U878 (N_878,In_1431,N_455);
xnor U879 (N_879,N_711,N_342);
or U880 (N_880,N_77,In_352);
nand U881 (N_881,N_661,N_194);
nor U882 (N_882,N_690,In_1361);
nor U883 (N_883,In_1548,In_660);
and U884 (N_884,In_1432,N_567);
or U885 (N_885,In_760,In_1053);
or U886 (N_886,N_195,In_1434);
or U887 (N_887,N_584,N_401);
nand U888 (N_888,In_969,In_80);
nor U889 (N_889,N_76,N_646);
or U890 (N_890,N_193,In_1323);
or U891 (N_891,In_932,N_191);
xor U892 (N_892,N_688,N_729);
and U893 (N_893,N_571,In_2178);
and U894 (N_894,In_1951,In_626);
nand U895 (N_895,In_2196,In_949);
or U896 (N_896,In_653,In_2203);
xnor U897 (N_897,In_562,In_730);
nand U898 (N_898,In_1672,In_686);
nor U899 (N_899,In_2410,N_618);
xor U900 (N_900,N_142,In_1044);
nand U901 (N_901,In_1824,N_274);
nand U902 (N_902,N_392,N_682);
nand U903 (N_903,In_1852,N_286);
xnor U904 (N_904,In_1107,In_2434);
nor U905 (N_905,N_645,In_1504);
nor U906 (N_906,In_2100,N_668);
and U907 (N_907,N_189,In_1821);
or U908 (N_908,N_555,In_548);
or U909 (N_909,In_588,In_814);
nand U910 (N_910,In_551,In_1743);
nand U911 (N_911,N_577,N_593);
nand U912 (N_912,In_987,In_184);
nor U913 (N_913,In_2244,N_659);
nor U914 (N_914,In_698,In_2291);
or U915 (N_915,In_141,N_508);
or U916 (N_916,In_1767,In_1076);
or U917 (N_917,N_591,In_2085);
or U918 (N_918,In_325,N_456);
or U919 (N_919,In_43,In_1408);
xor U920 (N_920,N_444,In_1635);
nand U921 (N_921,In_1505,In_1516);
or U922 (N_922,N_642,In_601);
xnor U923 (N_923,In_746,In_2246);
nor U924 (N_924,In_2264,N_315);
xor U925 (N_925,In_1009,In_2292);
nor U926 (N_926,In_2352,N_311);
nor U927 (N_927,N_554,N_702);
xor U928 (N_928,N_365,N_545);
nor U929 (N_929,In_2148,In_644);
and U930 (N_930,In_488,N_98);
and U931 (N_931,In_463,In_957);
nor U932 (N_932,In_57,In_419);
and U933 (N_933,In_115,N_461);
or U934 (N_934,In_944,In_2290);
nor U935 (N_935,N_40,N_256);
nor U936 (N_936,In_159,In_84);
nor U937 (N_937,In_260,N_533);
nand U938 (N_938,N_565,In_182);
nand U939 (N_939,In_1561,In_433);
nand U940 (N_940,In_1894,In_1396);
and U941 (N_941,In_1476,In_2135);
xor U942 (N_942,In_2416,In_1844);
and U943 (N_943,In_2419,In_1205);
and U944 (N_944,In_1324,In_1069);
and U945 (N_945,In_18,N_663);
nor U946 (N_946,In_690,In_58);
and U947 (N_947,In_2122,N_130);
or U948 (N_948,In_1148,In_156);
nor U949 (N_949,N_467,N_558);
nand U950 (N_950,In_1352,In_598);
or U951 (N_951,N_397,In_438);
or U952 (N_952,In_1878,In_117);
nand U953 (N_953,In_1450,In_1961);
xor U954 (N_954,In_540,N_167);
nor U955 (N_955,In_144,In_222);
xnor U956 (N_956,In_2111,N_339);
and U957 (N_957,In_2499,In_503);
xnor U958 (N_958,N_205,In_1356);
xor U959 (N_959,In_1397,In_975);
nand U960 (N_960,In_829,In_1498);
and U961 (N_961,N_288,In_457);
nor U962 (N_962,N_451,In_518);
or U963 (N_963,In_1592,In_1108);
nor U964 (N_964,In_902,N_260);
or U965 (N_965,In_559,N_627);
xor U966 (N_966,In_1486,In_931);
xnor U967 (N_967,N_589,N_570);
and U968 (N_968,In_1903,In_1524);
or U969 (N_969,N_700,N_701);
nand U970 (N_970,In_1669,In_1288);
or U971 (N_971,N_353,In_871);
and U972 (N_972,N_548,In_2101);
or U973 (N_973,In_2497,N_379);
nor U974 (N_974,N_562,N_621);
nand U975 (N_975,In_2061,In_1925);
xor U976 (N_976,N_362,In_2156);
nor U977 (N_977,N_25,In_1968);
or U978 (N_978,In_303,In_367);
xnor U979 (N_979,In_1950,In_443);
and U980 (N_980,In_1487,N_166);
xor U981 (N_981,In_197,In_2217);
and U982 (N_982,N_290,In_2326);
nand U983 (N_983,In_1238,In_1547);
nand U984 (N_984,N_395,In_1717);
nor U985 (N_985,N_313,In_339);
and U986 (N_986,N_117,In_2461);
xnor U987 (N_987,In_838,In_561);
or U988 (N_988,In_493,In_2243);
nand U989 (N_989,In_725,In_2107);
or U990 (N_990,In_1291,N_390);
and U991 (N_991,N_486,N_662);
nand U992 (N_992,In_2405,N_549);
or U993 (N_993,In_1183,In_2080);
xnor U994 (N_994,In_113,In_1368);
nor U995 (N_995,In_1796,In_781);
or U996 (N_996,In_29,N_411);
nand U997 (N_997,In_1813,In_1054);
nor U998 (N_998,In_2311,In_1834);
or U999 (N_999,In_1294,N_6);
and U1000 (N_1000,N_604,N_681);
or U1001 (N_1001,N_575,In_795);
or U1002 (N_1002,N_946,N_348);
and U1003 (N_1003,N_331,In_344);
nand U1004 (N_1004,N_669,In_1689);
nor U1005 (N_1005,In_49,N_149);
or U1006 (N_1006,N_716,N_827);
xor U1007 (N_1007,In_912,In_509);
and U1008 (N_1008,In_2050,N_744);
xnor U1009 (N_1009,In_905,In_894);
or U1010 (N_1010,In_1357,In_1074);
or U1011 (N_1011,N_818,In_455);
or U1012 (N_1012,In_363,In_2446);
or U1013 (N_1013,In_627,In_2466);
nor U1014 (N_1014,N_997,N_415);
and U1015 (N_1015,In_2094,N_839);
and U1016 (N_1016,N_692,In_2269);
nand U1017 (N_1017,N_501,In_1327);
nor U1018 (N_1018,In_2377,N_934);
nor U1019 (N_1019,In_2391,In_495);
nand U1020 (N_1020,N_134,In_868);
nand U1021 (N_1021,In_2019,N_199);
xnor U1022 (N_1022,N_599,N_278);
nand U1023 (N_1023,In_2063,In_2042);
or U1024 (N_1024,N_671,N_844);
nor U1025 (N_1025,In_2155,N_187);
and U1026 (N_1026,N_742,In_1110);
or U1027 (N_1027,In_2259,In_1802);
nor U1028 (N_1028,In_1184,N_874);
nand U1029 (N_1029,In_1553,In_779);
nand U1030 (N_1030,N_474,In_1920);
and U1031 (N_1031,In_701,In_200);
nand U1032 (N_1032,In_2037,N_805);
and U1033 (N_1033,In_1685,In_1889);
or U1034 (N_1034,In_1393,In_439);
and U1035 (N_1035,In_1177,In_1650);
or U1036 (N_1036,N_743,In_2036);
nor U1037 (N_1037,In_587,In_427);
xnor U1038 (N_1038,N_880,N_150);
and U1039 (N_1039,N_463,In_152);
xor U1040 (N_1040,In_2173,In_1991);
or U1041 (N_1041,In_12,In_426);
xor U1042 (N_1042,In_368,N_800);
nand U1043 (N_1043,In_594,N_641);
nand U1044 (N_1044,In_794,In_1389);
nor U1045 (N_1045,In_922,In_1391);
and U1046 (N_1046,In_239,N_580);
and U1047 (N_1047,N_634,In_2357);
nand U1048 (N_1048,N_781,In_261);
or U1049 (N_1049,In_1841,N_989);
nor U1050 (N_1050,N_132,In_1151);
nor U1051 (N_1051,N_541,In_1980);
or U1052 (N_1052,N_546,N_310);
or U1053 (N_1053,In_1549,In_2496);
nor U1054 (N_1054,In_2052,In_2260);
or U1055 (N_1055,In_1633,In_1186);
xor U1056 (N_1056,N_225,In_1863);
nand U1057 (N_1057,N_377,N_956);
nand U1058 (N_1058,N_612,N_517);
nor U1059 (N_1059,In_985,N_519);
or U1060 (N_1060,N_81,In_2302);
xnor U1061 (N_1061,N_326,In_1624);
and U1062 (N_1062,In_2449,In_2120);
and U1063 (N_1063,N_902,N_904);
nand U1064 (N_1064,In_2354,In_187);
nor U1065 (N_1065,In_735,In_633);
nand U1066 (N_1066,N_976,In_64);
and U1067 (N_1067,In_1761,In_321);
and U1068 (N_1068,In_1032,In_236);
nand U1069 (N_1069,N_709,In_960);
nand U1070 (N_1070,In_1754,N_724);
nor U1071 (N_1071,In_342,N_988);
nor U1072 (N_1072,N_950,In_945);
nor U1073 (N_1073,N_834,In_1115);
xnor U1074 (N_1074,In_1458,N_503);
and U1075 (N_1075,N_823,N_295);
nand U1076 (N_1076,N_349,N_941);
and U1077 (N_1077,N_180,N_387);
nor U1078 (N_1078,In_2254,N_234);
and U1079 (N_1079,In_136,In_1311);
and U1080 (N_1080,In_1371,In_226);
nor U1081 (N_1081,N_695,In_576);
nand U1082 (N_1082,N_605,In_2071);
xnor U1083 (N_1083,N_412,N_504);
xor U1084 (N_1084,N_869,In_2325);
and U1085 (N_1085,In_2338,In_1842);
xnor U1086 (N_1086,N_204,N_448);
and U1087 (N_1087,In_888,N_715);
or U1088 (N_1088,In_2421,N_992);
or U1089 (N_1089,In_154,In_2131);
xor U1090 (N_1090,In_2471,In_105);
nand U1091 (N_1091,In_1941,In_1459);
nor U1092 (N_1092,N_609,In_188);
nand U1093 (N_1093,In_221,In_1298);
and U1094 (N_1094,In_2312,N_815);
nor U1095 (N_1095,N_789,N_607);
xnor U1096 (N_1096,In_279,N_909);
nand U1097 (N_1097,In_926,N_859);
and U1098 (N_1098,In_676,In_460);
nor U1099 (N_1099,In_1163,In_1086);
nand U1100 (N_1100,N_521,In_2096);
xor U1101 (N_1101,N_747,In_757);
nand U1102 (N_1102,In_2304,N_696);
or U1103 (N_1103,N_264,In_1617);
and U1104 (N_1104,N_944,N_220);
xor U1105 (N_1105,In_2428,In_330);
or U1106 (N_1106,In_2152,N_380);
or U1107 (N_1107,In_1146,In_1850);
nor U1108 (N_1108,In_1942,In_2492);
xnor U1109 (N_1109,N_858,N_666);
nand U1110 (N_1110,N_705,In_531);
and U1111 (N_1111,N_772,N_878);
and U1112 (N_1112,N_836,N_2);
xor U1113 (N_1113,N_856,N_843);
and U1114 (N_1114,N_421,In_824);
nor U1115 (N_1115,N_176,N_816);
and U1116 (N_1116,N_863,N_790);
or U1117 (N_1117,N_99,N_845);
and U1118 (N_1118,In_122,N_862);
nor U1119 (N_1119,In_46,N_945);
or U1120 (N_1120,N_889,In_1279);
xnor U1121 (N_1121,N_986,In_2143);
and U1122 (N_1122,In_311,In_2383);
and U1123 (N_1123,In_387,In_678);
and U1124 (N_1124,In_308,In_2124);
or U1125 (N_1125,In_425,N_454);
nor U1126 (N_1126,In_764,In_328);
and U1127 (N_1127,In_114,In_19);
nor U1128 (N_1128,N_778,In_93);
nand U1129 (N_1129,In_2130,N_121);
nor U1130 (N_1130,N_756,In_407);
and U1131 (N_1131,In_2104,N_996);
nor U1132 (N_1132,In_1040,N_803);
xnor U1133 (N_1133,In_1546,In_688);
and U1134 (N_1134,In_1960,N_376);
nand U1135 (N_1135,N_179,N_817);
and U1136 (N_1136,N_38,In_1418);
and U1137 (N_1137,In_1971,N_670);
nor U1138 (N_1138,In_341,In_1411);
or U1139 (N_1139,In_2097,In_160);
nand U1140 (N_1140,N_207,N_63);
and U1141 (N_1141,In_677,In_1325);
nor U1142 (N_1142,N_667,N_48);
xnor U1143 (N_1143,In_137,N_737);
nand U1144 (N_1144,N_942,N_822);
and U1145 (N_1145,In_2046,In_287);
xnor U1146 (N_1146,In_1538,In_1483);
nor U1147 (N_1147,In_391,In_92);
nor U1148 (N_1148,N_296,N_768);
nand U1149 (N_1149,In_2409,N_678);
or U1150 (N_1150,N_472,N_324);
or U1151 (N_1151,In_2099,N_164);
nand U1152 (N_1152,N_957,N_0);
and U1153 (N_1153,In_110,In_745);
nand U1154 (N_1154,N_617,In_1935);
or U1155 (N_1155,In_581,In_575);
or U1156 (N_1156,In_106,N_511);
or U1157 (N_1157,N_939,N_613);
nor U1158 (N_1158,In_175,In_1453);
xnor U1159 (N_1159,In_1845,N_625);
or U1160 (N_1160,N_16,N_323);
nand U1161 (N_1161,N_973,In_192);
nor U1162 (N_1162,N_432,N_361);
nand U1163 (N_1163,N_606,N_979);
xor U1164 (N_1164,N_528,N_203);
nand U1165 (N_1165,N_600,N_564);
nand U1166 (N_1166,N_275,N_689);
nand U1167 (N_1167,In_1683,N_169);
nor U1168 (N_1168,In_1997,In_1570);
nand U1169 (N_1169,N_452,In_1265);
nor U1170 (N_1170,N_543,In_2119);
xnor U1171 (N_1171,N_11,In_1260);
and U1172 (N_1172,N_222,In_1194);
nand U1173 (N_1173,In_217,N_763);
nand U1174 (N_1174,In_674,In_52);
or U1175 (N_1175,In_1384,N_826);
or U1176 (N_1176,In_176,N_885);
or U1177 (N_1177,In_9,In_2022);
nand U1178 (N_1178,In_1979,In_685);
nand U1179 (N_1179,In_41,N_866);
xnor U1180 (N_1180,N_542,N_637);
nand U1181 (N_1181,N_766,N_470);
and U1182 (N_1182,In_494,In_2134);
nand U1183 (N_1183,In_872,In_91);
and U1184 (N_1184,In_462,In_2008);
nand U1185 (N_1185,In_785,In_1862);
nor U1186 (N_1186,In_1631,N_615);
xor U1187 (N_1187,N_384,In_672);
xor U1188 (N_1188,In_973,In_1220);
nand U1189 (N_1189,N_755,N_526);
nor U1190 (N_1190,In_26,N_21);
nand U1191 (N_1191,N_419,In_42);
nand U1192 (N_1192,N_809,N_44);
and U1193 (N_1193,In_721,N_966);
nand U1194 (N_1194,In_1753,In_770);
nor U1195 (N_1195,N_294,In_1462);
xor U1196 (N_1196,N_581,N_828);
and U1197 (N_1197,N_579,N_219);
or U1198 (N_1198,N_984,In_1642);
nand U1199 (N_1199,In_552,In_1908);
nor U1200 (N_1200,N_266,N_699);
nor U1201 (N_1201,N_761,In_1349);
or U1202 (N_1202,In_992,In_610);
nor U1203 (N_1203,In_827,N_891);
xnor U1204 (N_1204,In_2245,In_2360);
nor U1205 (N_1205,N_679,N_462);
nand U1206 (N_1206,N_213,N_721);
or U1207 (N_1207,In_104,In_329);
or U1208 (N_1208,N_720,In_734);
nand U1209 (N_1209,In_864,In_694);
and U1210 (N_1210,In_2379,In_498);
nor U1211 (N_1211,In_885,In_1488);
nor U1212 (N_1212,N_911,In_742);
or U1213 (N_1213,N_870,In_947);
xnor U1214 (N_1214,In_501,In_47);
nand U1215 (N_1215,In_2164,In_560);
xor U1216 (N_1216,N_753,N_231);
nand U1217 (N_1217,In_1891,In_2223);
nor U1218 (N_1218,In_2230,In_411);
and U1219 (N_1219,In_2162,In_1687);
nand U1220 (N_1220,In_1249,In_229);
and U1221 (N_1221,N_602,N_850);
and U1222 (N_1222,In_542,In_2070);
or U1223 (N_1223,In_309,In_1141);
or U1224 (N_1224,N_478,N_128);
nand U1225 (N_1225,N_15,In_1215);
nand U1226 (N_1226,N_127,In_1395);
xnor U1227 (N_1227,N_343,In_1680);
xor U1228 (N_1228,In_714,N_745);
xnor U1229 (N_1229,In_445,N_684);
xor U1230 (N_1230,In_1763,In_415);
and U1231 (N_1231,In_1978,N_466);
or U1232 (N_1232,N_748,N_948);
nand U1233 (N_1233,In_2192,In_1052);
nand U1234 (N_1234,In_267,N_760);
and U1235 (N_1235,In_6,In_988);
or U1236 (N_1236,In_689,N_631);
nand U1237 (N_1237,In_257,N_921);
or U1238 (N_1238,N_572,In_1124);
and U1239 (N_1239,N_947,N_417);
or U1240 (N_1240,In_2467,In_1405);
xnor U1241 (N_1241,In_165,In_2451);
or U1242 (N_1242,In_1367,N_513);
xnor U1243 (N_1243,In_262,In_1235);
xor U1244 (N_1244,In_1572,In_2195);
or U1245 (N_1245,N_243,In_81);
nand U1246 (N_1246,N_281,In_2268);
or U1247 (N_1247,In_2106,N_994);
or U1248 (N_1248,N_37,In_244);
nand U1249 (N_1249,In_1500,N_767);
nand U1250 (N_1250,N_1136,N_644);
xor U1251 (N_1251,N_303,N_675);
or U1252 (N_1252,N_757,N_1047);
nor U1253 (N_1253,In_2347,N_544);
or U1254 (N_1254,In_2298,N_665);
nor U1255 (N_1255,In_168,In_1928);
or U1256 (N_1256,N_1109,N_525);
xor U1257 (N_1257,In_1334,N_1224);
and U1258 (N_1258,In_2059,N_884);
and U1259 (N_1259,In_2401,N_1061);
xor U1260 (N_1260,In_1640,In_956);
nor U1261 (N_1261,In_461,In_1023);
xor U1262 (N_1262,N_1059,N_782);
xor U1263 (N_1263,N_917,N_658);
nand U1264 (N_1264,N_393,In_2216);
or U1265 (N_1265,N_758,N_244);
or U1266 (N_1266,N_708,N_514);
or U1267 (N_1267,N_913,In_1449);
xor U1268 (N_1268,In_253,In_1301);
xnor U1269 (N_1269,In_1905,N_853);
or U1270 (N_1270,N_797,In_1377);
xor U1271 (N_1271,In_1609,N_751);
and U1272 (N_1272,In_1071,In_848);
xnor U1273 (N_1273,N_1036,In_282);
and U1274 (N_1274,N_1177,N_842);
and U1275 (N_1275,In_497,N_1110);
xnor U1276 (N_1276,N_1009,In_418);
nand U1277 (N_1277,In_832,N_916);
nand U1278 (N_1278,In_1656,N_912);
xnor U1279 (N_1279,N_568,N_801);
and U1280 (N_1280,N_1053,In_1175);
nand U1281 (N_1281,N_1238,In_1837);
or U1282 (N_1282,In_1618,In_2167);
or U1283 (N_1283,In_107,N_94);
nor U1284 (N_1284,In_656,In_1812);
nor U1285 (N_1285,N_888,N_1153);
xor U1286 (N_1286,In_1706,N_907);
nand U1287 (N_1287,N_960,In_834);
xor U1288 (N_1288,N_656,In_489);
nor U1289 (N_1289,In_1659,In_1166);
nor U1290 (N_1290,N_9,In_881);
xor U1291 (N_1291,N_489,N_893);
xor U1292 (N_1292,N_1058,N_587);
and U1293 (N_1293,N_177,In_1610);
nor U1294 (N_1294,In_2058,N_1218);
xor U1295 (N_1295,N_733,In_1321);
and U1296 (N_1296,N_873,In_1278);
nand U1297 (N_1297,In_2207,N_143);
and U1298 (N_1298,In_967,In_1474);
nor U1299 (N_1299,N_1170,N_61);
nor U1300 (N_1300,N_1120,In_1939);
nor U1301 (N_1301,In_2218,N_1065);
xor U1302 (N_1302,In_1984,In_1661);
nor U1303 (N_1303,In_14,N_1052);
xor U1304 (N_1304,N_1183,In_2288);
nand U1305 (N_1305,In_510,In_1666);
or U1306 (N_1306,In_1122,N_1215);
and U1307 (N_1307,N_1051,N_363);
xnor U1308 (N_1308,In_1406,N_212);
nand U1309 (N_1309,N_900,N_1155);
nor U1310 (N_1310,N_931,N_963);
nor U1311 (N_1311,N_1222,In_2433);
and U1312 (N_1312,In_632,N_59);
nand U1313 (N_1313,N_1174,In_1299);
nand U1314 (N_1314,N_898,N_886);
nor U1315 (N_1315,N_1084,In_1800);
nor U1316 (N_1316,In_1923,In_1778);
or U1317 (N_1317,N_1242,N_970);
or U1318 (N_1318,N_872,N_468);
and U1319 (N_1319,N_892,In_980);
or U1320 (N_1320,In_1671,N_1208);
and U1321 (N_1321,N_1220,In_1473);
or U1322 (N_1322,N_1099,In_360);
xnor U1323 (N_1323,N_1054,In_1594);
nor U1324 (N_1324,N_928,N_978);
nand U1325 (N_1325,In_1247,In_472);
xor U1326 (N_1326,N_512,In_1127);
or U1327 (N_1327,In_1404,N_786);
or U1328 (N_1328,N_1032,In_487);
nand U1329 (N_1329,N_424,N_550);
xnor U1330 (N_1330,N_374,N_804);
nor U1331 (N_1331,N_969,N_1133);
nor U1332 (N_1332,N_883,In_1259);
nor U1333 (N_1333,N_999,In_1532);
nor U1334 (N_1334,N_50,In_1974);
nor U1335 (N_1335,In_1160,N_894);
nor U1336 (N_1336,N_594,In_2181);
and U1337 (N_1337,In_2317,In_1828);
xnor U1338 (N_1338,In_1514,N_732);
or U1339 (N_1339,N_1121,In_1227);
nand U1340 (N_1340,In_1152,N_1031);
and U1341 (N_1341,N_539,N_967);
nand U1342 (N_1342,N_1165,In_532);
or U1343 (N_1343,N_1198,N_1185);
nor U1344 (N_1344,In_1275,In_1884);
xnor U1345 (N_1345,N_409,In_546);
xnor U1346 (N_1346,N_1130,N_1161);
and U1347 (N_1347,In_1133,N_272);
nand U1348 (N_1348,N_408,In_230);
nor U1349 (N_1349,N_791,N_1168);
xnor U1350 (N_1350,In_358,In_1709);
nor U1351 (N_1351,In_1783,N_638);
nand U1352 (N_1352,N_1240,In_59);
xnor U1353 (N_1353,In_484,In_718);
nor U1354 (N_1354,In_1376,N_1191);
xor U1355 (N_1355,In_1682,In_2199);
or U1356 (N_1356,In_2067,In_1387);
xor U1357 (N_1357,N_672,In_1344);
nand U1358 (N_1358,In_408,N_814);
xnor U1359 (N_1359,N_154,In_406);
xnor U1360 (N_1360,In_1619,In_399);
or U1361 (N_1361,N_1069,In_1416);
nand U1362 (N_1362,In_1897,In_1029);
nand U1363 (N_1363,N_1034,N_1026);
nor U1364 (N_1364,N_100,N_1145);
and U1365 (N_1365,N_784,N_1140);
nor U1366 (N_1366,N_1017,N_1148);
nand U1367 (N_1367,In_761,In_1198);
nand U1368 (N_1368,N_520,In_2272);
and U1369 (N_1369,In_934,N_233);
and U1370 (N_1370,N_1201,In_593);
and U1371 (N_1371,N_46,N_710);
nand U1372 (N_1372,N_1232,In_2371);
xnor U1373 (N_1373,N_735,N_1236);
or U1374 (N_1374,N_626,N_70);
or U1375 (N_1375,In_1559,N_838);
nand U1376 (N_1376,In_2483,In_1945);
nor U1377 (N_1377,In_215,In_999);
nand U1378 (N_1378,N_1105,N_1092);
or U1379 (N_1379,In_1519,N_1107);
nor U1380 (N_1380,N_1007,N_1171);
xor U1381 (N_1381,In_1697,In_1218);
nand U1382 (N_1382,In_481,N_57);
nor U1383 (N_1383,In_747,N_1129);
or U1384 (N_1384,N_1164,N_788);
and U1385 (N_1385,N_1046,In_39);
xnor U1386 (N_1386,In_1287,N_1094);
or U1387 (N_1387,N_557,N_610);
nand U1388 (N_1388,In_1121,N_1076);
nand U1389 (N_1389,N_1075,N_1016);
and U1390 (N_1390,In_1646,In_1586);
xnor U1391 (N_1391,In_1059,In_1781);
xnor U1392 (N_1392,N_1,N_620);
and U1393 (N_1393,N_924,In_853);
and U1394 (N_1394,In_2422,In_389);
xor U1395 (N_1395,N_1122,N_776);
nor U1396 (N_1396,N_263,N_936);
nand U1397 (N_1397,In_940,In_942);
and U1398 (N_1398,N_596,N_1115);
nand U1399 (N_1399,In_683,N_1202);
or U1400 (N_1400,N_86,N_158);
nor U1401 (N_1401,N_935,In_1345);
or U1402 (N_1402,N_307,In_1007);
nand U1403 (N_1403,N_654,In_1825);
or U1404 (N_1404,N_406,In_1770);
or U1405 (N_1405,N_102,In_77);
xnor U1406 (N_1406,In_446,N_1087);
or U1407 (N_1407,N_1149,In_603);
or U1408 (N_1408,N_759,N_802);
xor U1409 (N_1409,In_1664,N_552);
and U1410 (N_1410,N_316,In_1302);
nor U1411 (N_1411,In_1793,N_1096);
or U1412 (N_1412,In_476,In_1833);
or U1413 (N_1413,In_354,N_561);
nand U1414 (N_1414,N_1213,N_1050);
or U1415 (N_1415,N_595,N_1089);
or U1416 (N_1416,In_127,In_658);
nor U1417 (N_1417,N_707,N_923);
or U1418 (N_1418,In_1000,N_405);
or U1419 (N_1419,In_622,In_717);
nand U1420 (N_1420,In_2429,In_174);
xnor U1421 (N_1421,N_1123,N_1249);
nor U1422 (N_1422,In_1554,N_833);
nor U1423 (N_1423,N_1248,In_1599);
or U1424 (N_1424,In_468,N_1081);
nand U1425 (N_1425,N_547,N_1028);
nand U1426 (N_1426,In_2228,N_1166);
or U1427 (N_1427,N_257,In_1537);
xor U1428 (N_1428,N_1231,N_962);
or U1429 (N_1429,In_1206,N_1211);
xor U1430 (N_1430,N_434,N_578);
xor U1431 (N_1431,In_2411,In_582);
nand U1432 (N_1432,In_346,N_146);
xnor U1433 (N_1433,In_143,In_963);
xnor U1434 (N_1434,N_1005,In_2188);
or U1435 (N_1435,N_1018,N_890);
and U1436 (N_1436,N_1124,In_2175);
and U1437 (N_1437,N_877,N_1015);
xor U1438 (N_1438,N_977,N_1066);
and U1439 (N_1439,In_1414,N_819);
nand U1440 (N_1440,N_1068,N_447);
nand U1441 (N_1441,In_1132,In_1342);
nor U1442 (N_1442,N_413,In_568);
xnor U1443 (N_1443,N_793,In_504);
and U1444 (N_1444,N_482,In_549);
xnor U1445 (N_1445,In_1856,In_402);
nor U1446 (N_1446,N_446,In_69);
xor U1447 (N_1447,In_2151,In_1673);
and U1448 (N_1448,In_1057,In_1154);
or U1449 (N_1449,N_855,N_1055);
and U1450 (N_1450,N_985,In_2407);
nand U1451 (N_1451,N_651,N_959);
xnor U1452 (N_1452,N_754,N_643);
nand U1453 (N_1453,N_691,In_1562);
xor U1454 (N_1454,In_2482,N_1228);
and U1455 (N_1455,N_284,In_185);
or U1456 (N_1456,N_163,N_388);
or U1457 (N_1457,N_1226,In_1900);
nand U1458 (N_1458,In_1157,N_1063);
nand U1459 (N_1459,In_1777,N_502);
nand U1460 (N_1460,N_500,In_1470);
and U1461 (N_1461,N_664,N_1188);
or U1462 (N_1462,N_837,N_940);
nand U1463 (N_1463,N_852,N_731);
nor U1464 (N_1464,In_502,In_179);
and U1465 (N_1465,N_499,N_373);
nand U1466 (N_1466,In_0,N_1118);
nor U1467 (N_1467,In_636,N_563);
xor U1468 (N_1468,N_1132,N_1138);
nor U1469 (N_1469,N_779,In_855);
nor U1470 (N_1470,In_1643,N_933);
xnor U1471 (N_1471,N_1135,N_304);
xnor U1472 (N_1472,In_1674,N_619);
or U1473 (N_1473,N_811,N_1013);
xnor U1474 (N_1474,In_232,N_29);
or U1475 (N_1475,In_2494,In_1955);
and U1476 (N_1476,In_1730,In_1645);
or U1477 (N_1477,N_1175,N_847);
or U1478 (N_1478,In_1117,N_1103);
nor U1479 (N_1479,N_824,In_1577);
nand U1480 (N_1480,N_832,N_653);
and U1481 (N_1481,In_1539,In_173);
xor U1482 (N_1482,N_831,In_2489);
or U1483 (N_1483,N_879,N_535);
nor U1484 (N_1484,N_559,N_1209);
nand U1485 (N_1485,In_1822,N_764);
and U1486 (N_1486,N_1243,N_1074);
nor U1487 (N_1487,N_723,N_1239);
nor U1488 (N_1488,In_440,In_2315);
nand U1489 (N_1489,N_346,In_2018);
or U1490 (N_1490,N_657,N_1203);
nand U1491 (N_1491,N_1150,N_247);
nand U1492 (N_1492,In_2294,N_1119);
and U1493 (N_1493,N_436,In_1831);
and U1494 (N_1494,In_1625,In_974);
xor U1495 (N_1495,N_722,N_1025);
xor U1496 (N_1496,N_955,In_1188);
xnor U1497 (N_1497,In_1039,In_1106);
nand U1498 (N_1498,In_1736,In_1947);
nand U1499 (N_1499,In_2237,In_1067);
xor U1500 (N_1500,N_1447,In_782);
or U1501 (N_1501,In_2420,In_522);
and U1502 (N_1502,N_611,In_259);
and U1503 (N_1503,N_165,N_1444);
nand U1504 (N_1504,In_1446,In_2301);
or U1505 (N_1505,N_1446,In_500);
or U1506 (N_1506,N_1196,N_1090);
xnor U1507 (N_1507,N_1237,N_835);
xor U1508 (N_1508,N_585,N_813);
or U1509 (N_1509,N_897,N_1478);
xor U1510 (N_1510,In_2229,N_583);
nor U1511 (N_1511,N_1156,In_553);
nor U1512 (N_1512,N_1382,N_769);
nand U1513 (N_1513,N_1178,N_1338);
and U1514 (N_1514,N_1040,N_1411);
or U1515 (N_1515,In_2153,N_1060);
nand U1516 (N_1516,N_1030,N_1284);
nand U1517 (N_1517,N_1400,N_459);
nor U1518 (N_1518,N_719,In_2249);
nor U1519 (N_1519,In_383,N_975);
and U1520 (N_1520,N_530,In_1143);
nor U1521 (N_1521,N_1113,In_646);
and U1522 (N_1522,N_325,In_1049);
xnor U1523 (N_1523,In_1787,N_1042);
and U1524 (N_1524,In_816,N_1290);
and U1525 (N_1525,In_1412,N_630);
nand U1526 (N_1526,N_980,In_2043);
xnor U1527 (N_1527,N_60,N_1386);
xnor U1528 (N_1528,N_1414,N_693);
nand U1529 (N_1529,In_1676,N_1483);
nand U1530 (N_1530,In_741,In_1285);
and U1531 (N_1531,N_1375,N_608);
nor U1532 (N_1532,In_550,N_810);
and U1533 (N_1533,In_1475,In_679);
nor U1534 (N_1534,N_1359,N_1184);
or U1535 (N_1535,N_648,N_1485);
nor U1536 (N_1536,N_137,In_1749);
xnor U1537 (N_1537,N_23,In_1246);
nand U1538 (N_1538,In_2266,N_590);
nor U1539 (N_1539,N_1383,In_1627);
and U1540 (N_1540,In_245,In_1606);
nand U1541 (N_1541,In_2465,In_1696);
nand U1542 (N_1542,N_124,N_875);
nand U1543 (N_1543,In_777,In_1254);
or U1544 (N_1544,In_1020,In_738);
and U1545 (N_1545,N_840,In_1670);
xor U1546 (N_1546,In_1170,N_1479);
nor U1547 (N_1547,N_1160,N_712);
and U1548 (N_1548,N_336,In_2066);
xnor U1549 (N_1549,In_1860,N_995);
and U1550 (N_1550,In_819,N_89);
or U1551 (N_1551,In_340,In_1350);
nand U1552 (N_1552,N_1426,In_1873);
and U1553 (N_1553,In_2248,In_2190);
nand U1554 (N_1554,N_556,N_1429);
nand U1555 (N_1555,N_1128,N_1043);
or U1556 (N_1556,In_146,In_1358);
xor U1557 (N_1557,N_43,In_390);
nor U1558 (N_1558,In_1638,N_200);
nor U1559 (N_1559,N_17,N_292);
xor U1560 (N_1560,N_1163,N_334);
nand U1561 (N_1561,In_2307,In_595);
nand U1562 (N_1562,In_1372,N_1278);
nor U1563 (N_1563,N_1337,In_1593);
or U1564 (N_1564,N_868,In_544);
or U1565 (N_1565,N_785,In_1062);
nor U1566 (N_1566,N_1271,N_1308);
nor U1567 (N_1567,In_1956,N_1112);
nor U1568 (N_1568,N_1001,N_1495);
and U1569 (N_1569,In_2056,In_1402);
and U1570 (N_1570,N_812,N_1085);
nand U1571 (N_1571,In_1967,In_1185);
and U1572 (N_1572,N_777,N_1323);
nand U1573 (N_1573,N_1420,N_407);
nand U1574 (N_1574,In_2250,N_1259);
nor U1575 (N_1575,N_492,In_2385);
xor U1576 (N_1576,N_1012,N_551);
or U1577 (N_1577,In_2481,N_507);
and U1578 (N_1578,In_851,In_2321);
and U1579 (N_1579,N_1438,In_2263);
nor U1580 (N_1580,N_841,N_1481);
nor U1581 (N_1581,In_634,In_2213);
xor U1582 (N_1582,N_864,N_1080);
xor U1583 (N_1583,N_106,N_153);
nor U1584 (N_1584,In_1921,N_1306);
xor U1585 (N_1585,N_181,N_952);
nand U1586 (N_1586,N_140,In_1911);
xor U1587 (N_1587,In_1027,N_1274);
xnor U1588 (N_1588,N_922,In_298);
nor U1589 (N_1589,N_1206,N_1403);
nor U1590 (N_1590,N_1314,In_1010);
nand U1591 (N_1591,N_1281,In_400);
xor U1592 (N_1592,N_1442,N_430);
or U1593 (N_1593,N_783,N_1397);
nand U1594 (N_1594,N_1082,In_1895);
or U1595 (N_1595,N_639,N_366);
nor U1596 (N_1596,N_750,In_2117);
xor U1597 (N_1597,In_1460,In_621);
or U1598 (N_1598,N_1435,N_1488);
or U1599 (N_1599,N_1179,In_129);
and U1600 (N_1600,N_253,N_1225);
and U1601 (N_1601,N_1456,In_1936);
nand U1602 (N_1602,In_1341,In_1774);
nand U1603 (N_1603,N_1341,In_1095);
and U1604 (N_1604,N_915,In_233);
nor U1605 (N_1605,In_586,N_982);
nand U1606 (N_1606,N_1360,N_1300);
nand U1607 (N_1607,In_118,N_1173);
nand U1608 (N_1608,In_1454,N_276);
nor U1609 (N_1609,N_1317,In_2160);
and U1610 (N_1610,In_492,N_1246);
or U1611 (N_1611,In_1699,N_1455);
or U1612 (N_1612,N_1471,In_1564);
xor U1613 (N_1613,In_1424,N_1292);
xnor U1614 (N_1614,N_319,In_661);
nand U1615 (N_1615,N_1086,In_94);
or U1616 (N_1616,N_1340,In_2336);
or U1617 (N_1617,In_1386,In_1348);
nand U1618 (N_1618,N_636,N_1408);
nand U1619 (N_1619,N_1095,In_246);
nor U1620 (N_1620,N_435,N_318);
nand U1621 (N_1621,In_370,N_974);
nand U1622 (N_1622,N_1044,In_345);
nand U1623 (N_1623,N_426,In_2375);
and U1624 (N_1624,N_1390,In_1149);
nand U1625 (N_1625,N_914,N_1297);
xor U1626 (N_1626,N_1335,In_1494);
or U1627 (N_1627,N_1358,N_920);
or U1628 (N_1628,N_1077,N_1487);
or U1629 (N_1629,N_740,N_1402);
or U1630 (N_1630,In_624,N_1428);
nand U1631 (N_1631,N_1440,N_1320);
and U1632 (N_1632,In_1861,In_1306);
or U1633 (N_1633,In_2308,N_1474);
and U1634 (N_1634,In_1409,N_1321);
nor U1635 (N_1635,N_4,N_640);
xnor U1636 (N_1636,N_1356,N_1493);
and U1637 (N_1637,N_794,N_532);
xnor U1638 (N_1638,In_801,N_458);
nor U1639 (N_1639,N_235,In_950);
or U1640 (N_1640,N_1264,In_2394);
or U1641 (N_1641,In_1308,N_345);
nand U1642 (N_1642,In_2180,N_887);
xor U1643 (N_1643,In_111,N_1385);
nor U1644 (N_1644,In_599,N_1365);
or U1645 (N_1645,N_943,In_48);
nor U1646 (N_1646,N_1433,In_833);
or U1647 (N_1647,In_1679,N_224);
nor U1648 (N_1648,In_1716,N_1366);
and U1649 (N_1649,In_1890,N_1205);
nand U1650 (N_1650,N_1258,In_1983);
nand U1651 (N_1651,In_754,In_50);
and U1652 (N_1652,In_1092,N_1024);
nor U1653 (N_1653,In_1252,In_482);
nand U1654 (N_1654,N_1457,N_1431);
nand U1655 (N_1655,N_796,N_1336);
or U1656 (N_1656,In_2079,N_717);
nand U1657 (N_1657,N_1022,N_1369);
nor U1658 (N_1658,N_1169,N_1079);
nor U1659 (N_1659,N_287,N_983);
nand U1660 (N_1660,N_901,N_1045);
or U1661 (N_1661,N_576,In_874);
nand U1662 (N_1662,N_1212,In_1533);
or U1663 (N_1663,N_1158,N_1295);
or U1664 (N_1664,N_1352,N_806);
or U1665 (N_1665,N_1014,N_1418);
xor U1666 (N_1666,N_1280,N_1137);
xor U1667 (N_1667,N_825,N_951);
nor U1668 (N_1668,N_1371,In_1513);
nor U1669 (N_1669,N_1421,N_1217);
xnor U1670 (N_1670,In_2267,N_792);
nand U1671 (N_1671,In_1790,In_1139);
nand U1672 (N_1672,N_1116,In_2432);
nand U1673 (N_1673,In_1421,N_1460);
nand U1674 (N_1674,In_2398,N_1270);
nand U1675 (N_1675,N_378,N_1393);
or U1676 (N_1676,N_647,N_1322);
nand U1677 (N_1677,In_1346,N_1011);
nor U1678 (N_1678,In_1875,N_1454);
and U1679 (N_1679,N_1354,In_1005);
or U1680 (N_1680,N_1473,In_2257);
and U1681 (N_1681,N_1003,N_1357);
or U1682 (N_1682,N_1453,In_22);
or U1683 (N_1683,In_1870,N_1468);
xnor U1684 (N_1684,In_2277,N_1362);
or U1685 (N_1685,In_1305,N_1497);
or U1686 (N_1686,In_964,N_403);
nand U1687 (N_1687,In_1775,N_1344);
nand U1688 (N_1688,N_1125,In_228);
or U1689 (N_1689,N_1412,In_2343);
and U1690 (N_1690,N_1364,N_1318);
nand U1691 (N_1691,In_1002,N_865);
and U1692 (N_1692,N_196,In_911);
xnor U1693 (N_1693,N_1033,N_899);
or U1694 (N_1694,N_1305,In_1033);
or U1695 (N_1695,N_987,N_741);
nand U1696 (N_1696,N_1376,N_131);
or U1697 (N_1697,In_994,N_1372);
or U1698 (N_1698,In_4,N_1367);
and U1699 (N_1699,N_1332,N_498);
and U1700 (N_1700,N_1253,N_1041);
and U1701 (N_1701,N_698,In_2020);
and U1702 (N_1702,N_170,N_1368);
nor U1703 (N_1703,N_1327,N_144);
nand U1704 (N_1704,N_1229,N_1396);
and U1705 (N_1705,In_1745,In_1262);
or U1706 (N_1706,N_1269,N_795);
or U1707 (N_1707,In_2296,N_1247);
nand U1708 (N_1708,N_1381,In_1688);
nand U1709 (N_1709,In_2116,In_2110);
nor U1710 (N_1710,N_1190,In_1741);
xor U1711 (N_1711,N_1039,N_919);
or U1712 (N_1712,In_1426,N_1325);
or U1713 (N_1713,N_787,N_993);
or U1714 (N_1714,N_771,In_867);
nand U1715 (N_1715,N_1293,In_1681);
nand U1716 (N_1716,N_1291,N_333);
xnor U1717 (N_1717,N_1415,N_1216);
nor U1718 (N_1718,N_968,In_5);
nand U1719 (N_1719,N_1282,In_748);
nor U1720 (N_1720,N_728,N_141);
nor U1721 (N_1721,N_1151,In_1042);
nand U1722 (N_1722,In_736,N_88);
and U1723 (N_1723,In_669,N_770);
nor U1724 (N_1724,N_1250,N_1091);
or U1725 (N_1725,In_700,N_1000);
xnor U1726 (N_1726,N_714,N_335);
and U1727 (N_1727,N_270,In_307);
nand U1728 (N_1728,N_1349,In_1063);
xor U1729 (N_1729,N_1154,N_425);
and U1730 (N_1730,N_1498,N_1230);
and U1731 (N_1731,N_1283,N_1370);
or U1732 (N_1732,N_1277,N_445);
and U1733 (N_1733,In_2000,In_1517);
xnor U1734 (N_1734,N_1285,In_2392);
nor U1735 (N_1735,In_148,N_522);
or U1736 (N_1736,N_683,In_1123);
or U1737 (N_1737,N_1021,N_1252);
nor U1738 (N_1738,N_1267,N_1223);
nand U1739 (N_1739,N_857,N_1159);
or U1740 (N_1740,In_289,In_1159);
and U1741 (N_1741,In_520,In_893);
or U1742 (N_1742,N_1439,In_1466);
nor U1743 (N_1743,N_26,N_1353);
nand U1744 (N_1744,In_1604,N_1469);
and U1745 (N_1745,N_31,N_1221);
and U1746 (N_1746,N_1445,N_236);
and U1747 (N_1747,N_1117,N_1329);
and U1748 (N_1748,N_1263,N_1200);
nand U1749 (N_1749,N_457,N_1157);
or U1750 (N_1750,N_1600,N_1450);
and U1751 (N_1751,N_1547,In_1596);
nand U1752 (N_1752,N_1740,N_460);
and U1753 (N_1753,N_1062,N_1152);
or U1754 (N_1754,N_1576,In_2275);
nor U1755 (N_1755,N_752,In_579);
nand U1756 (N_1756,N_1592,N_1127);
nand U1757 (N_1757,N_1738,N_1275);
or U1758 (N_1758,In_673,N_1593);
and U1759 (N_1759,N_1507,In_567);
nand U1760 (N_1760,N_1537,N_1687);
nor U1761 (N_1761,N_1570,N_1027);
and U1762 (N_1762,N_953,N_1131);
nor U1763 (N_1763,N_1665,N_746);
nor U1764 (N_1764,N_1539,N_910);
nor U1765 (N_1765,N_1699,N_1565);
nand U1766 (N_1766,N_1348,N_1560);
nand U1767 (N_1767,N_849,N_1134);
nor U1768 (N_1768,In_571,N_1611);
and U1769 (N_1769,N_1588,In_2320);
or U1770 (N_1770,N_42,In_2069);
and U1771 (N_1771,In_486,In_865);
nor U1772 (N_1772,In_1212,N_1744);
nand U1773 (N_1773,In_1600,N_64);
nor U1774 (N_1774,In_1362,N_27);
nand U1775 (N_1775,N_523,In_109);
xnor U1776 (N_1776,N_1342,In_2437);
nand U1777 (N_1777,N_1683,N_1484);
or U1778 (N_1778,N_1476,In_1353);
or U1779 (N_1779,N_1416,N_1298);
nand U1780 (N_1780,N_1696,In_1147);
nand U1781 (N_1781,In_1966,N_1727);
nor U1782 (N_1782,N_1670,N_1573);
nand U1783 (N_1783,N_1605,N_1346);
xor U1784 (N_1784,N_660,N_1745);
and U1785 (N_1785,N_1666,In_1290);
nand U1786 (N_1786,N_1635,N_509);
and U1787 (N_1787,N_1279,N_19);
xnor U1788 (N_1788,N_1698,N_1502);
or U1789 (N_1789,In_1079,N_1741);
xnor U1790 (N_1790,N_1413,N_1591);
nor U1791 (N_1791,In_821,N_1647);
and U1792 (N_1792,In_2273,In_772);
nand U1793 (N_1793,N_727,N_1747);
xor U1794 (N_1794,In_2299,N_1345);
nand U1795 (N_1795,N_1363,N_1723);
and U1796 (N_1796,In_276,N_676);
nor U1797 (N_1797,N_1374,N_1580);
nand U1798 (N_1798,N_537,N_1603);
xnor U1799 (N_1799,N_1489,In_324);
nor U1800 (N_1800,N_1722,N_1608);
or U1801 (N_1801,N_1430,N_1561);
and U1802 (N_1802,N_906,N_1615);
nor U1803 (N_1803,N_650,In_1883);
and U1804 (N_1804,In_1698,N_1577);
xor U1805 (N_1805,N_1659,N_93);
xor U1806 (N_1806,N_1564,N_932);
xnor U1807 (N_1807,N_1527,N_1690);
or U1808 (N_1808,N_1679,In_299);
xnor U1809 (N_1809,N_1002,N_255);
or U1810 (N_1810,N_1581,In_1511);
xnor U1811 (N_1811,N_1186,N_1310);
and U1812 (N_1812,In_1240,N_1715);
nor U1813 (N_1813,In_273,N_1181);
nor U1814 (N_1814,N_1008,N_1695);
xnor U1815 (N_1815,N_1713,N_1401);
or U1816 (N_1816,N_1452,N_1301);
nand U1817 (N_1817,N_540,In_1191);
or U1818 (N_1818,N_1563,N_1669);
and U1819 (N_1819,N_1541,N_930);
nor U1820 (N_1820,N_1227,N_516);
nor U1821 (N_1821,N_1552,N_829);
nor U1822 (N_1822,N_1097,In_707);
nor U1823 (N_1823,N_1162,N_1704);
xnor U1824 (N_1824,N_937,N_1590);
or U1825 (N_1825,N_1141,N_1522);
and U1826 (N_1826,In_2062,In_2406);
or U1827 (N_1827,N_991,N_1568);
and U1828 (N_1828,N_1422,In_8);
xor U1829 (N_1829,In_842,N_1709);
nand U1830 (N_1830,N_1494,N_1614);
xnor U1831 (N_1831,N_762,N_1671);
or U1832 (N_1832,N_1689,N_1071);
and U1833 (N_1833,N_1392,N_1101);
and U1834 (N_1834,N_614,N_1607);
and U1835 (N_1835,N_1667,N_1648);
nor U1836 (N_1836,In_1193,N_1579);
and U1837 (N_1837,N_1718,N_1712);
and U1838 (N_1838,N_1730,N_1705);
nor U1839 (N_1839,N_1651,N_1549);
xnor U1840 (N_1840,N_1302,In_847);
nand U1841 (N_1841,In_1723,N_1287);
nor U1842 (N_1842,N_1531,N_1645);
nand U1843 (N_1843,N_1637,N_1700);
xor U1844 (N_1844,N_1543,N_1313);
xor U1845 (N_1845,N_954,N_1143);
nand U1846 (N_1846,In_1364,N_926);
or U1847 (N_1847,N_1328,N_1571);
xor U1848 (N_1848,N_1417,N_83);
xnor U1849 (N_1849,N_1503,N_929);
xor U1850 (N_1850,N_927,In_682);
nand U1851 (N_1851,N_1538,N_1621);
nor U1852 (N_1852,N_1574,N_1004);
xor U1853 (N_1853,N_1703,N_91);
xnor U1854 (N_1854,N_998,N_1424);
xnor U1855 (N_1855,N_1628,N_1601);
xnor U1856 (N_1856,N_726,N_1048);
xor U1857 (N_1857,N_1406,N_773);
nand U1858 (N_1858,N_1387,In_1899);
nand U1859 (N_1859,N_896,In_1490);
xnor U1860 (N_1860,N_1404,N_1187);
nor U1861 (N_1861,N_1681,N_1664);
and U1862 (N_1862,N_1521,N_1180);
nor U1863 (N_1863,N_1299,N_1104);
nand U1864 (N_1864,N_1589,In_2445);
or U1865 (N_1865,N_1199,N_1437);
or U1866 (N_1866,N_1739,N_1254);
xnor U1867 (N_1867,N_1304,In_528);
nor U1868 (N_1868,In_589,In_2253);
or U1869 (N_1869,In_297,N_1195);
xor U1870 (N_1870,N_1146,N_1093);
or U1871 (N_1871,N_1204,In_2163);
and U1872 (N_1872,N_1307,In_702);
xor U1873 (N_1873,N_1613,In_1225);
xor U1874 (N_1874,N_480,N_1674);
or U1875 (N_1875,N_1622,N_1147);
nor U1876 (N_1876,In_1226,N_494);
or U1877 (N_1877,N_1644,In_1912);
or U1878 (N_1878,N_332,In_2030);
nor U1879 (N_1879,N_1643,In_1501);
nor U1880 (N_1880,N_1525,In_654);
nor U1881 (N_1881,N_1049,N_1554);
or U1882 (N_1882,N_1661,N_1691);
nand U1883 (N_1883,N_1654,N_1490);
and U1884 (N_1884,N_1569,In_703);
and U1885 (N_1885,N_1189,N_1624);
nor U1886 (N_1886,N_1673,N_1423);
xor U1887 (N_1887,In_570,In_1401);
or U1888 (N_1888,N_1334,N_1662);
nor U1889 (N_1889,N_347,N_1266);
and U1890 (N_1890,N_1126,N_338);
or U1891 (N_1891,N_1315,N_112);
nor U1892 (N_1892,N_477,N_1518);
xnor U1893 (N_1893,In_376,N_1678);
xor U1894 (N_1894,N_1466,N_168);
or U1895 (N_1895,N_1725,N_1652);
nor U1896 (N_1896,N_1556,N_506);
nor U1897 (N_1897,N_1532,N_569);
or U1898 (N_1898,N_1514,N_1655);
xor U1899 (N_1899,N_1558,N_1316);
nor U1900 (N_1900,N_1692,In_1690);
nand U1901 (N_1901,N_1509,N_1035);
or U1902 (N_1902,In_1579,N_1587);
nand U1903 (N_1903,N_1330,N_1214);
and U1904 (N_1904,N_1144,In_962);
or U1905 (N_1905,N_1114,N_1377);
and U1906 (N_1906,In_220,N_1708);
xor U1907 (N_1907,N_1639,N_938);
and U1908 (N_1908,N_449,N_1496);
xor U1909 (N_1909,N_1395,N_1710);
nand U1910 (N_1910,N_1536,N_1660);
and U1911 (N_1911,N_1410,N_1331);
nor U1912 (N_1912,N_1482,In_1085);
xor U1913 (N_1913,N_1504,N_624);
and U1914 (N_1914,N_1480,N_1653);
xnor U1915 (N_1915,In_263,In_883);
xor U1916 (N_1916,N_1542,N_1734);
and U1917 (N_1917,N_1407,N_1510);
or U1918 (N_1918,N_1519,N_1088);
xnor U1919 (N_1919,N_1501,In_268);
nor U1920 (N_1920,N_1398,N_107);
nand U1921 (N_1921,N_1584,N_1630);
and U1922 (N_1922,N_1530,N_1567);
xor U1923 (N_1923,N_1343,In_1542);
nor U1924 (N_1924,N_1257,N_1486);
xor U1925 (N_1925,In_326,N_1272);
or U1926 (N_1926,N_1078,N_1702);
nor U1927 (N_1927,In_2141,N_655);
nor U1928 (N_1928,N_1067,N_1550);
and U1929 (N_1929,N_1492,N_1534);
or U1930 (N_1930,In_547,N_1288);
nand U1931 (N_1931,N_674,In_2072);
and U1932 (N_1932,In_2372,In_292);
or U1933 (N_1933,N_1139,N_1706);
and U1934 (N_1934,N_774,N_1056);
nand U1935 (N_1935,N_1557,N_971);
xor U1936 (N_1936,N_775,In_364);
xor U1937 (N_1937,In_740,N_1646);
nor U1938 (N_1938,N_990,N_1618);
nand U1939 (N_1939,In_943,N_1355);
nand U1940 (N_1940,N_1737,N_730);
xor U1941 (N_1941,In_925,N_1599);
nand U1942 (N_1942,N_152,N_876);
or U1943 (N_1943,N_1451,N_734);
or U1944 (N_1944,N_680,N_1535);
or U1945 (N_1945,In_2479,N_1658);
or U1946 (N_1946,N_1720,In_2083);
and U1947 (N_1947,N_1566,N_871);
and U1948 (N_1948,In_2103,N_1436);
nand U1949 (N_1949,In_1590,In_1786);
or U1950 (N_1950,N_1555,N_1023);
nand U1951 (N_1951,In_2053,In_2382);
xnor U1952 (N_1952,N_1234,N_1642);
and U1953 (N_1953,N_1668,In_1799);
nor U1954 (N_1954,In_1705,N_1684);
and U1955 (N_1955,N_1207,N_1721);
and U1956 (N_1956,N_1586,N_854);
nor U1957 (N_1957,In_1988,N_1072);
nand U1958 (N_1958,N_1736,N_173);
nor U1959 (N_1959,N_1256,N_566);
and U1960 (N_1960,N_821,N_1749);
and U1961 (N_1961,N_1729,N_1006);
nand U1962 (N_1962,N_1499,N_958);
xnor U1963 (N_1963,In_620,N_1038);
nor U1964 (N_1964,In_1051,N_1609);
nor U1965 (N_1965,In_135,N_981);
nor U1966 (N_1966,N_1688,N_1513);
and U1967 (N_1967,N_1477,N_400);
xnor U1968 (N_1968,N_1623,N_820);
and U1969 (N_1969,N_598,N_1373);
and U1970 (N_1970,N_1582,In_2136);
nor U1971 (N_1971,N_861,N_1019);
or U1972 (N_1972,N_738,N_1508);
and U1973 (N_1973,In_2150,In_1552);
xor U1974 (N_1974,N_808,N_1606);
and U1975 (N_1975,N_1548,N_1467);
or U1976 (N_1976,N_592,N_799);
nand U1977 (N_1977,In_1129,N_488);
or U1978 (N_1978,In_1451,In_696);
and U1979 (N_1979,N_404,N_1462);
and U1980 (N_1980,N_1261,N_122);
and U1981 (N_1981,N_1449,N_807);
and U1982 (N_1982,N_1620,N_534);
or U1983 (N_1983,N_1512,N_1102);
xor U1984 (N_1984,N_1575,N_232);
xnor U1985 (N_1985,N_1172,N_588);
xnor U1986 (N_1986,N_1731,N_1638);
nor U1987 (N_1987,In_235,N_185);
or U1988 (N_1988,N_299,In_1868);
and U1989 (N_1989,N_972,N_1732);
or U1990 (N_1990,N_1309,N_1350);
nand U1991 (N_1991,N_1167,N_202);
xor U1992 (N_1992,In_858,N_1241);
and U1993 (N_1993,N_1333,N_903);
or U1994 (N_1994,N_1636,N_961);
and U1995 (N_1995,N_1443,N_1551);
and U1996 (N_1996,In_1739,N_1578);
nand U1997 (N_1997,N_1726,In_1780);
nor U1998 (N_1998,N_905,N_918);
or U1999 (N_1999,N_1632,In_269);
nor U2000 (N_2000,N_1545,In_306);
nor U2001 (N_2001,N_1617,In_1794);
nor U2002 (N_2002,N_495,N_1768);
or U2003 (N_2003,N_1929,N_1733);
and U2004 (N_2004,N_1798,N_1742);
nand U2005 (N_2005,N_1846,N_1759);
and U2006 (N_2006,N_1906,N_1901);
xnor U2007 (N_2007,N_1993,In_895);
or U2008 (N_2008,N_1711,N_1952);
and U2009 (N_2009,N_1470,N_1553);
or U2010 (N_2010,N_1904,N_1935);
or U2011 (N_2011,N_1070,N_1676);
and U2012 (N_2012,N_1235,N_249);
nand U2013 (N_2013,N_895,N_1656);
nor U2014 (N_2014,N_1845,N_1852);
xnor U2015 (N_2015,In_61,N_1735);
nand U2016 (N_2016,In_1785,N_1182);
or U2017 (N_2017,N_1289,N_1836);
nand U2018 (N_2018,N_1245,N_1625);
xor U2019 (N_2019,N_1766,N_1192);
or U2020 (N_2020,N_1793,N_1763);
xnor U2021 (N_2021,N_1980,N_1441);
nor U2022 (N_2022,N_1037,N_1544);
and U2023 (N_2023,N_1758,N_1529);
nand U2024 (N_2024,N_1819,N_1516);
nor U2025 (N_2025,N_1934,N_1627);
nand U2026 (N_2026,N_1379,In_720);
xor U2027 (N_2027,N_1251,N_1860);
nand U2028 (N_2028,N_1779,N_1851);
or U2029 (N_2029,N_1319,In_2039);
nand U2030 (N_2030,N_1461,N_1890);
xor U2031 (N_2031,N_1783,N_1506);
xor U2032 (N_2032,N_1850,In_767);
and U2033 (N_2033,N_713,In_264);
xor U2034 (N_2034,N_1693,N_1546);
or U2035 (N_2035,N_1864,N_536);
xnor U2036 (N_2036,N_1391,N_1210);
xor U2037 (N_2037,In_629,N_1965);
nor U2038 (N_2038,In_90,N_515);
xnor U2039 (N_2039,N_1663,N_1524);
or U2040 (N_2040,N_1882,N_1932);
nand U2041 (N_2041,N_1106,N_1871);
nand U2042 (N_2042,N_1878,N_1859);
or U2043 (N_2043,N_1863,N_1986);
and U2044 (N_2044,N_1883,N_1631);
xor U2045 (N_2045,N_1974,N_1719);
and U2046 (N_2046,In_1963,N_1312);
nand U2047 (N_2047,N_1848,N_1459);
or U2048 (N_2048,N_1855,N_1835);
nand U2049 (N_2049,N_1957,N_1815);
nor U2050 (N_2050,N_1953,N_300);
or U2051 (N_2051,N_1602,N_1812);
and U2052 (N_2052,In_1568,N_1910);
or U2053 (N_2053,N_531,N_1806);
and U2054 (N_2054,N_1427,N_1785);
and U2055 (N_2055,N_1870,N_1955);
xor U2056 (N_2056,N_1083,N_1672);
xnor U2057 (N_2057,N_1533,N_450);
or U2058 (N_2058,In_1089,N_1978);
and U2059 (N_2059,In_2102,N_151);
nand U2060 (N_2060,N_1982,In_1464);
and U2061 (N_2061,N_1912,In_651);
or U2062 (N_2062,N_1865,N_1276);
xor U2063 (N_2063,N_1784,N_1800);
nor U2064 (N_2064,N_1448,In_723);
or U2065 (N_2065,N_485,N_1751);
xnor U2066 (N_2066,In_1176,N_1597);
nor U2067 (N_2067,N_1964,N_1142);
and U2068 (N_2068,N_1832,N_1820);
or U2069 (N_2069,N_1787,In_1684);
xnor U2070 (N_2070,N_1892,N_1849);
nand U2071 (N_2071,N_1598,N_1996);
xnor U2072 (N_2072,In_89,N_1831);
nor U2073 (N_2073,N_1425,N_1791);
and U2074 (N_2074,N_1020,N_1924);
or U2075 (N_2075,N_56,N_1802);
nand U2076 (N_2076,N_1515,N_1724);
nand U2077 (N_2077,N_1987,N_1959);
xnor U2078 (N_2078,N_1389,N_1778);
nor U2079 (N_2079,N_1286,N_830);
and U2080 (N_2080,N_1891,N_1828);
xor U2081 (N_2081,N_1975,N_1844);
xnor U2082 (N_2082,N_1823,N_1193);
nor U2083 (N_2083,N_1682,N_1794);
and U2084 (N_2084,N_1889,N_1840);
xnor U2085 (N_2085,In_2442,In_2005);
nor U2086 (N_2086,N_1874,N_1967);
nor U2087 (N_2087,N_1777,N_1866);
and U2088 (N_2088,N_882,N_1838);
nand U2089 (N_2089,N_780,N_1754);
and U2090 (N_2090,N_1789,N_1686);
xnor U2091 (N_2091,N_1098,In_1957);
and U2092 (N_2092,N_1817,N_1985);
xor U2093 (N_2093,N_1931,N_1813);
xnor U2094 (N_2094,N_1528,In_927);
xnor U2095 (N_2095,N_1176,N_1991);
xnor U2096 (N_2096,N_1361,N_1790);
nand U2097 (N_2097,N_1233,N_1807);
or U2098 (N_2098,N_1916,N_394);
and U2099 (N_2099,N_1970,N_1463);
nor U2100 (N_2100,N_1979,N_1886);
or U2101 (N_2101,N_1983,N_437);
or U2102 (N_2102,N_1936,N_1797);
nand U2103 (N_2103,N_1219,N_1853);
nand U2104 (N_2104,N_949,N_1833);
and U2105 (N_2105,N_1940,N_1816);
and U2106 (N_2106,N_1895,N_1857);
xnor U2107 (N_2107,N_344,N_1994);
and U2108 (N_2108,N_1294,In_448);
nand U2109 (N_2109,In_1964,N_1010);
and U2110 (N_2110,N_1933,N_1707);
nor U2111 (N_2111,N_1100,N_7);
xnor U2112 (N_2112,N_1847,N_1971);
nor U2113 (N_2113,N_327,N_1756);
xnor U2114 (N_2114,N_1868,N_1938);
and U2115 (N_2115,N_1902,N_1939);
or U2116 (N_2116,N_1755,N_261);
nand U2117 (N_2117,N_1827,N_1872);
or U2118 (N_2118,N_1887,N_1907);
nand U2119 (N_2119,N_1780,N_1595);
nor U2120 (N_2120,N_1057,N_649);
xnor U2121 (N_2121,N_1594,N_867);
nand U2122 (N_2122,N_1896,N_1399);
xnor U2123 (N_2123,In_1477,In_873);
and U2124 (N_2124,N_1612,In_1130);
nand U2125 (N_2125,N_1394,N_1714);
nand U2126 (N_2126,N_1562,N_1753);
xor U2127 (N_2127,N_1884,N_1856);
nor U2128 (N_2128,N_1610,N_1818);
or U2129 (N_2129,N_1905,N_1900);
xor U2130 (N_2130,N_1804,N_1701);
and U2131 (N_2131,N_1771,N_1262);
or U2132 (N_2132,In_1995,N_1743);
nor U2133 (N_2133,N_1409,In_2393);
and U2134 (N_2134,N_1776,N_1619);
nor U2135 (N_2135,N_1908,N_860);
or U2136 (N_2136,N_1862,N_1717);
nor U2137 (N_2137,In_1211,N_1825);
and U2138 (N_2138,N_1511,N_1893);
xor U2139 (N_2139,N_846,N_1941);
and U2140 (N_2140,N_1491,In_789);
nand U2141 (N_2141,In_753,N_1943);
nand U2142 (N_2142,N_1772,N_1927);
or U2143 (N_2143,In_473,N_798);
nand U2144 (N_2144,N_1604,N_1926);
nand U2145 (N_2145,N_1918,N_1990);
nor U2146 (N_2146,In_435,N_1244);
nor U2147 (N_2147,N_1919,N_1821);
nor U2148 (N_2148,N_1822,In_1972);
xnor U2149 (N_2149,N_1748,N_1572);
nand U2150 (N_2150,N_1111,N_1757);
xor U2151 (N_2151,N_1716,N_1914);
or U2152 (N_2152,In_1208,N_925);
or U2153 (N_2153,N_1949,N_1951);
nand U2154 (N_2154,N_1500,N_1803);
and U2155 (N_2155,N_1903,N_1786);
nor U2156 (N_2156,N_1347,N_1770);
nand U2157 (N_2157,N_1894,N_1762);
xor U2158 (N_2158,N_1255,N_1915);
or U2159 (N_2159,N_1326,N_1775);
xor U2160 (N_2160,N_1782,N_1311);
nand U2161 (N_2161,In_699,N_1945);
and U2162 (N_2162,N_1956,In_1282);
xnor U2163 (N_2163,N_1958,N_1464);
and U2164 (N_2164,N_1829,N_240);
nand U2165 (N_2165,N_881,In_2221);
nand U2166 (N_2166,N_1999,N_1273);
xnor U2167 (N_2167,N_1378,N_1843);
nor U2168 (N_2168,N_1881,N_1963);
or U2169 (N_2169,N_1922,N_1928);
or U2170 (N_2170,N_1750,N_1826);
xor U2171 (N_2171,N_1858,N_1774);
nor U2172 (N_2172,N_1830,N_1942);
or U2173 (N_2173,N_1675,N_1616);
nor U2174 (N_2174,In_2359,N_1995);
xor U2175 (N_2175,N_1432,N_1434);
nor U2176 (N_2176,N_1897,N_1997);
and U2177 (N_2177,N_1977,N_1876);
nor U2178 (N_2178,N_1268,N_1765);
xor U2179 (N_2179,N_1801,N_1640);
xor U2180 (N_2180,N_1197,N_1339);
and U2181 (N_2181,N_1961,N_1966);
or U2182 (N_2182,N_1808,N_1805);
xnor U2183 (N_2183,N_1517,N_1944);
or U2184 (N_2184,N_1540,N_306);
or U2185 (N_2185,N_1954,N_113);
and U2186 (N_2186,N_1388,N_1913);
xor U2187 (N_2187,N_1968,N_1898);
xor U2188 (N_2188,N_1885,N_1324);
and U2189 (N_2189,N_1880,N_851);
xor U2190 (N_2190,N_1962,N_1969);
or U2191 (N_2191,N_1925,N_1472);
or U2192 (N_2192,N_1680,N_1405);
nand U2193 (N_2193,In_195,N_1626);
xnor U2194 (N_2194,In_1244,N_1923);
nor U2195 (N_2195,N_1988,N_171);
xor U2196 (N_2196,N_1781,N_1649);
or U2197 (N_2197,N_1984,N_1937);
nand U2198 (N_2198,N_1769,N_1930);
or U2199 (N_2199,N_1909,N_1920);
nor U2200 (N_2200,N_254,N_1760);
nor U2201 (N_2201,N_1950,N_765);
or U2202 (N_2202,N_1384,N_1073);
nand U2203 (N_2203,N_1869,N_1911);
nor U2204 (N_2204,N_1505,N_1788);
and U2205 (N_2205,N_965,N_1657);
and U2206 (N_2206,N_1877,N_1998);
nor U2207 (N_2207,N_1972,In_918);
xor U2208 (N_2208,N_1260,N_1921);
xnor U2209 (N_2209,N_1583,N_1559);
nor U2210 (N_2210,N_1792,N_1989);
and U2211 (N_2211,N_1746,N_481);
and U2212 (N_2212,N_1694,N_1351);
or U2213 (N_2213,In_1061,N_1811);
xnor U2214 (N_2214,N_1773,N_1265);
or U2215 (N_2215,N_1520,N_1960);
and U2216 (N_2216,N_1475,N_1796);
nor U2217 (N_2217,N_1834,N_1899);
or U2218 (N_2218,N_1981,N_1685);
nand U2219 (N_2219,N_1992,N_1947);
nor U2220 (N_2220,In_1075,N_1839);
and U2221 (N_2221,N_1795,N_1633);
and U2222 (N_2222,N_964,N_1824);
or U2223 (N_2223,N_1629,N_1641);
nand U2224 (N_2224,N_1875,In_75);
nand U2225 (N_2225,N_1380,In_1805);
or U2226 (N_2226,N_1809,N_1767);
or U2227 (N_2227,In_1270,N_1650);
nor U2228 (N_2228,N_908,N_1029);
xnor U2229 (N_2229,N_848,N_1064);
nor U2230 (N_2230,N_1108,N_1526);
or U2231 (N_2231,N_1728,N_1296);
nand U2232 (N_2232,N_1973,N_1585);
and U2233 (N_2233,N_1764,In_2439);
and U2234 (N_2234,N_1814,N_1888);
nand U2235 (N_2235,N_1948,N_1799);
or U2236 (N_2236,N_1946,N_1697);
and U2237 (N_2237,N_1752,N_1419);
and U2238 (N_2238,N_1873,N_1465);
or U2239 (N_2239,N_1917,N_1861);
nand U2240 (N_2240,N_1634,N_1303);
xor U2241 (N_2241,N_1854,N_1879);
or U2242 (N_2242,N_1194,N_1976);
and U2243 (N_2243,N_396,N_1761);
and U2244 (N_2244,N_1523,In_583);
nor U2245 (N_2245,N_1810,N_1842);
and U2246 (N_2246,N_1837,N_1458);
xor U2247 (N_2247,N_1841,N_1867);
nand U2248 (N_2248,In_413,N_1677);
xor U2249 (N_2249,N_1596,In_2399);
nand U2250 (N_2250,N_2013,N_2087);
or U2251 (N_2251,N_2142,N_2026);
and U2252 (N_2252,N_2214,N_2229);
nand U2253 (N_2253,N_2008,N_2213);
and U2254 (N_2254,N_2245,N_2248);
or U2255 (N_2255,N_2007,N_2084);
nand U2256 (N_2256,N_2190,N_2183);
nor U2257 (N_2257,N_2057,N_2083);
nor U2258 (N_2258,N_2135,N_2067);
or U2259 (N_2259,N_2097,N_2046);
and U2260 (N_2260,N_2092,N_2033);
xor U2261 (N_2261,N_2003,N_2212);
nand U2262 (N_2262,N_2231,N_2112);
nand U2263 (N_2263,N_2088,N_2004);
and U2264 (N_2264,N_2158,N_2078);
xor U2265 (N_2265,N_2193,N_2030);
nor U2266 (N_2266,N_2133,N_2058);
and U2267 (N_2267,N_2143,N_2093);
nor U2268 (N_2268,N_2187,N_2049);
or U2269 (N_2269,N_2232,N_2059);
xor U2270 (N_2270,N_2146,N_2230);
and U2271 (N_2271,N_2085,N_2120);
nand U2272 (N_2272,N_2042,N_2101);
nor U2273 (N_2273,N_2073,N_2186);
nand U2274 (N_2274,N_2243,N_2156);
nor U2275 (N_2275,N_2096,N_2028);
or U2276 (N_2276,N_2063,N_2237);
nor U2277 (N_2277,N_2197,N_2218);
nor U2278 (N_2278,N_2136,N_2211);
nor U2279 (N_2279,N_2148,N_2208);
xnor U2280 (N_2280,N_2216,N_2036);
or U2281 (N_2281,N_2130,N_2239);
or U2282 (N_2282,N_2098,N_2246);
nor U2283 (N_2283,N_2124,N_2094);
or U2284 (N_2284,N_2116,N_2210);
nor U2285 (N_2285,N_2020,N_2110);
nand U2286 (N_2286,N_2188,N_2189);
and U2287 (N_2287,N_2150,N_2090);
nand U2288 (N_2288,N_2200,N_2009);
xor U2289 (N_2289,N_2141,N_2226);
or U2290 (N_2290,N_2069,N_2053);
or U2291 (N_2291,N_2126,N_2076);
and U2292 (N_2292,N_2151,N_2249);
and U2293 (N_2293,N_2119,N_2192);
and U2294 (N_2294,N_2080,N_2018);
nor U2295 (N_2295,N_2244,N_2123);
or U2296 (N_2296,N_2041,N_2002);
nor U2297 (N_2297,N_2198,N_2115);
nand U2298 (N_2298,N_2086,N_2064);
xor U2299 (N_2299,N_2241,N_2223);
nand U2300 (N_2300,N_2131,N_2127);
or U2301 (N_2301,N_2164,N_2109);
xor U2302 (N_2302,N_2068,N_2048);
or U2303 (N_2303,N_2104,N_2144);
xor U2304 (N_2304,N_2196,N_2180);
and U2305 (N_2305,N_2065,N_2016);
and U2306 (N_2306,N_2015,N_2107);
and U2307 (N_2307,N_2052,N_2228);
and U2308 (N_2308,N_2176,N_2159);
nand U2309 (N_2309,N_2075,N_2105);
or U2310 (N_2310,N_2175,N_2235);
and U2311 (N_2311,N_2160,N_2155);
nand U2312 (N_2312,N_2081,N_2027);
nor U2313 (N_2313,N_2022,N_2061);
nor U2314 (N_2314,N_2163,N_2034);
and U2315 (N_2315,N_2000,N_2204);
and U2316 (N_2316,N_2103,N_2099);
nand U2317 (N_2317,N_2157,N_2082);
xnor U2318 (N_2318,N_2024,N_2201);
and U2319 (N_2319,N_2219,N_2066);
nand U2320 (N_2320,N_2031,N_2145);
and U2321 (N_2321,N_2217,N_2209);
nor U2322 (N_2322,N_2234,N_2025);
and U2323 (N_2323,N_2060,N_2170);
nor U2324 (N_2324,N_2132,N_2137);
nor U2325 (N_2325,N_2247,N_2147);
and U2326 (N_2326,N_2012,N_2173);
nand U2327 (N_2327,N_2039,N_2023);
nor U2328 (N_2328,N_2040,N_2017);
nor U2329 (N_2329,N_2113,N_2162);
and U2330 (N_2330,N_2233,N_2220);
nand U2331 (N_2331,N_2128,N_2240);
xnor U2332 (N_2332,N_2047,N_2011);
or U2333 (N_2333,N_2152,N_2054);
and U2334 (N_2334,N_2169,N_2038);
nand U2335 (N_2335,N_2079,N_2185);
xor U2336 (N_2336,N_2056,N_2014);
and U2337 (N_2337,N_2165,N_2102);
nor U2338 (N_2338,N_2074,N_2010);
nor U2339 (N_2339,N_2154,N_2117);
nor U2340 (N_2340,N_2203,N_2174);
nand U2341 (N_2341,N_2019,N_2177);
nor U2342 (N_2342,N_2227,N_2006);
or U2343 (N_2343,N_2238,N_2050);
nor U2344 (N_2344,N_2171,N_2051);
xor U2345 (N_2345,N_2055,N_2222);
xor U2346 (N_2346,N_2181,N_2100);
or U2347 (N_2347,N_2195,N_2236);
nand U2348 (N_2348,N_2125,N_2184);
nor U2349 (N_2349,N_2037,N_2089);
or U2350 (N_2350,N_2202,N_2191);
or U2351 (N_2351,N_2106,N_2178);
nor U2352 (N_2352,N_2207,N_2029);
xor U2353 (N_2353,N_2070,N_2224);
nor U2354 (N_2354,N_2153,N_2149);
xor U2355 (N_2355,N_2172,N_2122);
xor U2356 (N_2356,N_2205,N_2095);
or U2357 (N_2357,N_2182,N_2206);
and U2358 (N_2358,N_2035,N_2062);
nor U2359 (N_2359,N_2194,N_2111);
or U2360 (N_2360,N_2108,N_2001);
nand U2361 (N_2361,N_2005,N_2045);
nor U2362 (N_2362,N_2118,N_2071);
xor U2363 (N_2363,N_2225,N_2167);
xor U2364 (N_2364,N_2043,N_2114);
xor U2365 (N_2365,N_2032,N_2139);
nand U2366 (N_2366,N_2199,N_2129);
and U2367 (N_2367,N_2242,N_2168);
and U2368 (N_2368,N_2140,N_2044);
or U2369 (N_2369,N_2166,N_2215);
nand U2370 (N_2370,N_2134,N_2091);
or U2371 (N_2371,N_2072,N_2121);
nand U2372 (N_2372,N_2077,N_2138);
or U2373 (N_2373,N_2179,N_2221);
or U2374 (N_2374,N_2161,N_2021);
nor U2375 (N_2375,N_2121,N_2220);
nor U2376 (N_2376,N_2235,N_2065);
nor U2377 (N_2377,N_2176,N_2164);
and U2378 (N_2378,N_2026,N_2171);
nor U2379 (N_2379,N_2238,N_2168);
xor U2380 (N_2380,N_2182,N_2014);
nor U2381 (N_2381,N_2207,N_2185);
xor U2382 (N_2382,N_2233,N_2083);
or U2383 (N_2383,N_2010,N_2152);
xor U2384 (N_2384,N_2085,N_2046);
xnor U2385 (N_2385,N_2226,N_2222);
nand U2386 (N_2386,N_2174,N_2114);
nor U2387 (N_2387,N_2197,N_2005);
nand U2388 (N_2388,N_2033,N_2063);
nand U2389 (N_2389,N_2098,N_2047);
or U2390 (N_2390,N_2050,N_2002);
nor U2391 (N_2391,N_2045,N_2080);
xor U2392 (N_2392,N_2007,N_2052);
or U2393 (N_2393,N_2030,N_2114);
nand U2394 (N_2394,N_2054,N_2059);
nand U2395 (N_2395,N_2057,N_2228);
nor U2396 (N_2396,N_2046,N_2000);
nor U2397 (N_2397,N_2100,N_2015);
and U2398 (N_2398,N_2214,N_2056);
nor U2399 (N_2399,N_2161,N_2060);
nor U2400 (N_2400,N_2155,N_2095);
nor U2401 (N_2401,N_2231,N_2182);
nand U2402 (N_2402,N_2111,N_2081);
xor U2403 (N_2403,N_2140,N_2214);
and U2404 (N_2404,N_2206,N_2091);
nor U2405 (N_2405,N_2036,N_2103);
nor U2406 (N_2406,N_2111,N_2207);
nor U2407 (N_2407,N_2104,N_2205);
nor U2408 (N_2408,N_2187,N_2161);
or U2409 (N_2409,N_2192,N_2174);
xnor U2410 (N_2410,N_2047,N_2144);
nor U2411 (N_2411,N_2190,N_2008);
and U2412 (N_2412,N_2037,N_2013);
xnor U2413 (N_2413,N_2129,N_2016);
or U2414 (N_2414,N_2054,N_2067);
or U2415 (N_2415,N_2142,N_2068);
xnor U2416 (N_2416,N_2157,N_2186);
and U2417 (N_2417,N_2212,N_2223);
or U2418 (N_2418,N_2203,N_2171);
xnor U2419 (N_2419,N_2140,N_2194);
or U2420 (N_2420,N_2188,N_2109);
or U2421 (N_2421,N_2017,N_2112);
nor U2422 (N_2422,N_2162,N_2223);
nand U2423 (N_2423,N_2058,N_2123);
nand U2424 (N_2424,N_2193,N_2007);
and U2425 (N_2425,N_2024,N_2183);
xnor U2426 (N_2426,N_2010,N_2247);
xnor U2427 (N_2427,N_2214,N_2117);
nor U2428 (N_2428,N_2180,N_2168);
or U2429 (N_2429,N_2091,N_2205);
nor U2430 (N_2430,N_2132,N_2057);
xnor U2431 (N_2431,N_2159,N_2197);
nand U2432 (N_2432,N_2080,N_2101);
and U2433 (N_2433,N_2178,N_2172);
nor U2434 (N_2434,N_2140,N_2146);
nand U2435 (N_2435,N_2032,N_2055);
xor U2436 (N_2436,N_2069,N_2015);
or U2437 (N_2437,N_2141,N_2131);
xnor U2438 (N_2438,N_2015,N_2064);
and U2439 (N_2439,N_2089,N_2011);
and U2440 (N_2440,N_2216,N_2224);
nor U2441 (N_2441,N_2134,N_2022);
nand U2442 (N_2442,N_2170,N_2212);
or U2443 (N_2443,N_2177,N_2075);
xor U2444 (N_2444,N_2150,N_2040);
nand U2445 (N_2445,N_2244,N_2093);
xor U2446 (N_2446,N_2238,N_2230);
nor U2447 (N_2447,N_2164,N_2098);
nor U2448 (N_2448,N_2199,N_2249);
nor U2449 (N_2449,N_2023,N_2183);
nor U2450 (N_2450,N_2057,N_2031);
and U2451 (N_2451,N_2133,N_2097);
nor U2452 (N_2452,N_2087,N_2247);
xor U2453 (N_2453,N_2215,N_2220);
xnor U2454 (N_2454,N_2028,N_2151);
nor U2455 (N_2455,N_2033,N_2107);
and U2456 (N_2456,N_2015,N_2031);
or U2457 (N_2457,N_2249,N_2164);
or U2458 (N_2458,N_2223,N_2184);
nand U2459 (N_2459,N_2104,N_2003);
or U2460 (N_2460,N_2133,N_2139);
or U2461 (N_2461,N_2054,N_2096);
xnor U2462 (N_2462,N_2051,N_2148);
xnor U2463 (N_2463,N_2128,N_2080);
xnor U2464 (N_2464,N_2147,N_2089);
nand U2465 (N_2465,N_2059,N_2205);
xor U2466 (N_2466,N_2012,N_2194);
or U2467 (N_2467,N_2075,N_2011);
or U2468 (N_2468,N_2092,N_2094);
and U2469 (N_2469,N_2097,N_2028);
and U2470 (N_2470,N_2238,N_2091);
nand U2471 (N_2471,N_2152,N_2249);
nor U2472 (N_2472,N_2079,N_2033);
or U2473 (N_2473,N_2099,N_2024);
or U2474 (N_2474,N_2183,N_2139);
nand U2475 (N_2475,N_2136,N_2074);
nor U2476 (N_2476,N_2102,N_2163);
nor U2477 (N_2477,N_2065,N_2218);
and U2478 (N_2478,N_2129,N_2105);
and U2479 (N_2479,N_2012,N_2156);
xor U2480 (N_2480,N_2131,N_2145);
and U2481 (N_2481,N_2045,N_2106);
xor U2482 (N_2482,N_2205,N_2006);
or U2483 (N_2483,N_2103,N_2023);
or U2484 (N_2484,N_2176,N_2228);
and U2485 (N_2485,N_2201,N_2177);
or U2486 (N_2486,N_2126,N_2035);
or U2487 (N_2487,N_2242,N_2219);
nand U2488 (N_2488,N_2115,N_2202);
xnor U2489 (N_2489,N_2165,N_2235);
xor U2490 (N_2490,N_2135,N_2124);
xor U2491 (N_2491,N_2159,N_2028);
xor U2492 (N_2492,N_2100,N_2062);
xor U2493 (N_2493,N_2131,N_2064);
xnor U2494 (N_2494,N_2185,N_2196);
or U2495 (N_2495,N_2194,N_2134);
xnor U2496 (N_2496,N_2245,N_2167);
nand U2497 (N_2497,N_2139,N_2245);
and U2498 (N_2498,N_2054,N_2226);
nor U2499 (N_2499,N_2169,N_2027);
nor U2500 (N_2500,N_2390,N_2469);
nand U2501 (N_2501,N_2480,N_2373);
and U2502 (N_2502,N_2376,N_2445);
nand U2503 (N_2503,N_2474,N_2352);
or U2504 (N_2504,N_2328,N_2499);
or U2505 (N_2505,N_2484,N_2314);
nor U2506 (N_2506,N_2355,N_2455);
nor U2507 (N_2507,N_2354,N_2333);
xor U2508 (N_2508,N_2312,N_2387);
or U2509 (N_2509,N_2475,N_2345);
or U2510 (N_2510,N_2460,N_2407);
xor U2511 (N_2511,N_2436,N_2440);
xor U2512 (N_2512,N_2365,N_2476);
or U2513 (N_2513,N_2358,N_2256);
nor U2514 (N_2514,N_2275,N_2496);
and U2515 (N_2515,N_2270,N_2493);
and U2516 (N_2516,N_2393,N_2450);
or U2517 (N_2517,N_2367,N_2439);
nand U2518 (N_2518,N_2297,N_2250);
nand U2519 (N_2519,N_2409,N_2471);
and U2520 (N_2520,N_2265,N_2410);
xor U2521 (N_2521,N_2391,N_2428);
nor U2522 (N_2522,N_2281,N_2363);
or U2523 (N_2523,N_2336,N_2261);
xor U2524 (N_2524,N_2382,N_2285);
nor U2525 (N_2525,N_2449,N_2424);
xnor U2526 (N_2526,N_2286,N_2403);
nor U2527 (N_2527,N_2431,N_2309);
or U2528 (N_2528,N_2346,N_2421);
and U2529 (N_2529,N_2444,N_2262);
or U2530 (N_2530,N_2448,N_2263);
or U2531 (N_2531,N_2451,N_2377);
nor U2532 (N_2532,N_2260,N_2498);
and U2533 (N_2533,N_2276,N_2385);
or U2534 (N_2534,N_2413,N_2492);
nor U2535 (N_2535,N_2349,N_2402);
nand U2536 (N_2536,N_2405,N_2386);
xnor U2537 (N_2537,N_2299,N_2366);
nor U2538 (N_2538,N_2462,N_2304);
nand U2539 (N_2539,N_2441,N_2458);
nor U2540 (N_2540,N_2267,N_2378);
xor U2541 (N_2541,N_2338,N_2488);
nand U2542 (N_2542,N_2490,N_2434);
and U2543 (N_2543,N_2470,N_2326);
nor U2544 (N_2544,N_2330,N_2303);
xnor U2545 (N_2545,N_2478,N_2257);
and U2546 (N_2546,N_2271,N_2334);
xor U2547 (N_2547,N_2425,N_2381);
and U2548 (N_2548,N_2408,N_2278);
and U2549 (N_2549,N_2322,N_2273);
or U2550 (N_2550,N_2368,N_2307);
nor U2551 (N_2551,N_2310,N_2432);
or U2552 (N_2552,N_2341,N_2411);
and U2553 (N_2553,N_2362,N_2423);
nor U2554 (N_2554,N_2394,N_2292);
or U2555 (N_2555,N_2351,N_2348);
or U2556 (N_2556,N_2347,N_2427);
and U2557 (N_2557,N_2259,N_2319);
or U2558 (N_2558,N_2486,N_2400);
nor U2559 (N_2559,N_2252,N_2302);
xor U2560 (N_2560,N_2472,N_2388);
and U2561 (N_2561,N_2477,N_2456);
or U2562 (N_2562,N_2308,N_2426);
or U2563 (N_2563,N_2282,N_2331);
nand U2564 (N_2564,N_2283,N_2437);
or U2565 (N_2565,N_2277,N_2464);
nand U2566 (N_2566,N_2438,N_2318);
and U2567 (N_2567,N_2343,N_2300);
and U2568 (N_2568,N_2459,N_2274);
nor U2569 (N_2569,N_2287,N_2399);
nor U2570 (N_2570,N_2372,N_2481);
nor U2571 (N_2571,N_2266,N_2397);
or U2572 (N_2572,N_2453,N_2284);
or U2573 (N_2573,N_2418,N_2296);
nand U2574 (N_2574,N_2442,N_2433);
or U2575 (N_2575,N_2396,N_2406);
and U2576 (N_2576,N_2447,N_2494);
or U2577 (N_2577,N_2419,N_2301);
xor U2578 (N_2578,N_2268,N_2384);
nor U2579 (N_2579,N_2329,N_2251);
nand U2580 (N_2580,N_2311,N_2482);
nand U2581 (N_2581,N_2392,N_2294);
nand U2582 (N_2582,N_2272,N_2253);
nand U2583 (N_2583,N_2461,N_2356);
nor U2584 (N_2584,N_2337,N_2415);
nand U2585 (N_2585,N_2401,N_2305);
nor U2586 (N_2586,N_2374,N_2264);
xor U2587 (N_2587,N_2357,N_2457);
or U2588 (N_2588,N_2443,N_2468);
and U2589 (N_2589,N_2306,N_2254);
nand U2590 (N_2590,N_2422,N_2313);
nand U2591 (N_2591,N_2290,N_2452);
nand U2592 (N_2592,N_2317,N_2454);
nand U2593 (N_2593,N_2435,N_2340);
and U2594 (N_2594,N_2269,N_2371);
and U2595 (N_2595,N_2327,N_2350);
xnor U2596 (N_2596,N_2473,N_2417);
xor U2597 (N_2597,N_2446,N_2320);
or U2598 (N_2598,N_2295,N_2279);
nand U2599 (N_2599,N_2398,N_2342);
xnor U2600 (N_2600,N_2258,N_2332);
nand U2601 (N_2601,N_2335,N_2414);
nor U2602 (N_2602,N_2339,N_2429);
or U2603 (N_2603,N_2495,N_2420);
and U2604 (N_2604,N_2491,N_2395);
nand U2605 (N_2605,N_2465,N_2466);
and U2606 (N_2606,N_2353,N_2412);
nor U2607 (N_2607,N_2479,N_2323);
xor U2608 (N_2608,N_2370,N_2404);
nor U2609 (N_2609,N_2325,N_2293);
or U2610 (N_2610,N_2416,N_2430);
nand U2611 (N_2611,N_2463,N_2361);
and U2612 (N_2612,N_2483,N_2280);
nand U2613 (N_2613,N_2359,N_2489);
or U2614 (N_2614,N_2344,N_2291);
xor U2615 (N_2615,N_2375,N_2380);
nand U2616 (N_2616,N_2288,N_2298);
xnor U2617 (N_2617,N_2389,N_2379);
nand U2618 (N_2618,N_2383,N_2360);
xor U2619 (N_2619,N_2315,N_2289);
nor U2620 (N_2620,N_2255,N_2321);
xor U2621 (N_2621,N_2316,N_2324);
and U2622 (N_2622,N_2369,N_2497);
or U2623 (N_2623,N_2487,N_2467);
nor U2624 (N_2624,N_2485,N_2364);
or U2625 (N_2625,N_2422,N_2439);
nand U2626 (N_2626,N_2286,N_2416);
nand U2627 (N_2627,N_2335,N_2461);
or U2628 (N_2628,N_2494,N_2273);
or U2629 (N_2629,N_2265,N_2448);
and U2630 (N_2630,N_2344,N_2355);
xor U2631 (N_2631,N_2307,N_2469);
nand U2632 (N_2632,N_2477,N_2351);
nor U2633 (N_2633,N_2369,N_2424);
nor U2634 (N_2634,N_2381,N_2283);
or U2635 (N_2635,N_2491,N_2434);
xnor U2636 (N_2636,N_2289,N_2402);
nand U2637 (N_2637,N_2332,N_2397);
nand U2638 (N_2638,N_2468,N_2450);
nor U2639 (N_2639,N_2499,N_2312);
xnor U2640 (N_2640,N_2284,N_2493);
nand U2641 (N_2641,N_2448,N_2330);
nor U2642 (N_2642,N_2310,N_2495);
nand U2643 (N_2643,N_2362,N_2458);
xnor U2644 (N_2644,N_2264,N_2482);
nand U2645 (N_2645,N_2471,N_2415);
nor U2646 (N_2646,N_2324,N_2415);
and U2647 (N_2647,N_2296,N_2275);
or U2648 (N_2648,N_2350,N_2472);
xor U2649 (N_2649,N_2395,N_2442);
xnor U2650 (N_2650,N_2269,N_2475);
nand U2651 (N_2651,N_2336,N_2340);
nand U2652 (N_2652,N_2405,N_2487);
nor U2653 (N_2653,N_2364,N_2351);
and U2654 (N_2654,N_2308,N_2266);
and U2655 (N_2655,N_2446,N_2270);
or U2656 (N_2656,N_2273,N_2404);
xnor U2657 (N_2657,N_2400,N_2411);
xor U2658 (N_2658,N_2341,N_2321);
and U2659 (N_2659,N_2498,N_2461);
nand U2660 (N_2660,N_2372,N_2418);
nand U2661 (N_2661,N_2423,N_2368);
nor U2662 (N_2662,N_2362,N_2414);
xor U2663 (N_2663,N_2495,N_2474);
nor U2664 (N_2664,N_2455,N_2477);
or U2665 (N_2665,N_2274,N_2257);
nand U2666 (N_2666,N_2468,N_2315);
nand U2667 (N_2667,N_2407,N_2457);
nand U2668 (N_2668,N_2370,N_2357);
and U2669 (N_2669,N_2276,N_2258);
or U2670 (N_2670,N_2384,N_2283);
and U2671 (N_2671,N_2456,N_2276);
nand U2672 (N_2672,N_2420,N_2478);
nand U2673 (N_2673,N_2451,N_2282);
nand U2674 (N_2674,N_2300,N_2400);
nor U2675 (N_2675,N_2341,N_2400);
xnor U2676 (N_2676,N_2484,N_2478);
or U2677 (N_2677,N_2307,N_2257);
xor U2678 (N_2678,N_2374,N_2254);
xor U2679 (N_2679,N_2298,N_2354);
nand U2680 (N_2680,N_2405,N_2350);
or U2681 (N_2681,N_2349,N_2369);
and U2682 (N_2682,N_2358,N_2381);
and U2683 (N_2683,N_2449,N_2371);
and U2684 (N_2684,N_2459,N_2252);
or U2685 (N_2685,N_2372,N_2496);
or U2686 (N_2686,N_2290,N_2435);
nor U2687 (N_2687,N_2381,N_2411);
and U2688 (N_2688,N_2485,N_2492);
xor U2689 (N_2689,N_2365,N_2290);
nand U2690 (N_2690,N_2255,N_2445);
nor U2691 (N_2691,N_2437,N_2357);
nand U2692 (N_2692,N_2358,N_2456);
nand U2693 (N_2693,N_2448,N_2408);
nor U2694 (N_2694,N_2331,N_2276);
nand U2695 (N_2695,N_2460,N_2322);
nor U2696 (N_2696,N_2390,N_2389);
nor U2697 (N_2697,N_2380,N_2425);
nand U2698 (N_2698,N_2302,N_2371);
or U2699 (N_2699,N_2444,N_2339);
or U2700 (N_2700,N_2339,N_2256);
or U2701 (N_2701,N_2280,N_2365);
nor U2702 (N_2702,N_2298,N_2270);
or U2703 (N_2703,N_2485,N_2394);
nor U2704 (N_2704,N_2296,N_2449);
nor U2705 (N_2705,N_2467,N_2328);
xor U2706 (N_2706,N_2268,N_2450);
or U2707 (N_2707,N_2433,N_2290);
and U2708 (N_2708,N_2321,N_2489);
nor U2709 (N_2709,N_2281,N_2412);
nand U2710 (N_2710,N_2308,N_2298);
or U2711 (N_2711,N_2434,N_2257);
nor U2712 (N_2712,N_2275,N_2344);
nor U2713 (N_2713,N_2262,N_2381);
nand U2714 (N_2714,N_2262,N_2324);
nand U2715 (N_2715,N_2413,N_2353);
or U2716 (N_2716,N_2315,N_2260);
or U2717 (N_2717,N_2275,N_2332);
and U2718 (N_2718,N_2320,N_2415);
xnor U2719 (N_2719,N_2477,N_2330);
xor U2720 (N_2720,N_2362,N_2317);
nor U2721 (N_2721,N_2387,N_2462);
xor U2722 (N_2722,N_2302,N_2347);
xnor U2723 (N_2723,N_2413,N_2488);
nand U2724 (N_2724,N_2287,N_2430);
nor U2725 (N_2725,N_2409,N_2387);
nand U2726 (N_2726,N_2256,N_2409);
nand U2727 (N_2727,N_2460,N_2377);
nand U2728 (N_2728,N_2368,N_2382);
or U2729 (N_2729,N_2285,N_2415);
or U2730 (N_2730,N_2348,N_2340);
xor U2731 (N_2731,N_2428,N_2439);
nand U2732 (N_2732,N_2304,N_2497);
or U2733 (N_2733,N_2279,N_2350);
nor U2734 (N_2734,N_2372,N_2276);
xnor U2735 (N_2735,N_2498,N_2335);
nor U2736 (N_2736,N_2261,N_2258);
or U2737 (N_2737,N_2405,N_2435);
nor U2738 (N_2738,N_2285,N_2260);
xor U2739 (N_2739,N_2265,N_2405);
and U2740 (N_2740,N_2358,N_2331);
nor U2741 (N_2741,N_2446,N_2272);
and U2742 (N_2742,N_2434,N_2331);
nor U2743 (N_2743,N_2344,N_2294);
and U2744 (N_2744,N_2287,N_2492);
or U2745 (N_2745,N_2284,N_2402);
or U2746 (N_2746,N_2335,N_2366);
xor U2747 (N_2747,N_2400,N_2463);
xnor U2748 (N_2748,N_2495,N_2292);
and U2749 (N_2749,N_2407,N_2356);
or U2750 (N_2750,N_2747,N_2618);
and U2751 (N_2751,N_2538,N_2624);
nor U2752 (N_2752,N_2639,N_2688);
and U2753 (N_2753,N_2603,N_2622);
nand U2754 (N_2754,N_2595,N_2502);
or U2755 (N_2755,N_2581,N_2615);
xor U2756 (N_2756,N_2719,N_2686);
xnor U2757 (N_2757,N_2580,N_2633);
and U2758 (N_2758,N_2642,N_2501);
nor U2759 (N_2759,N_2535,N_2721);
nand U2760 (N_2760,N_2579,N_2628);
or U2761 (N_2761,N_2706,N_2527);
nor U2762 (N_2762,N_2729,N_2715);
nor U2763 (N_2763,N_2515,N_2740);
nand U2764 (N_2764,N_2528,N_2597);
xor U2765 (N_2765,N_2551,N_2672);
nand U2766 (N_2766,N_2649,N_2604);
nand U2767 (N_2767,N_2687,N_2522);
or U2768 (N_2768,N_2629,N_2609);
nand U2769 (N_2769,N_2608,N_2557);
or U2770 (N_2770,N_2554,N_2505);
xor U2771 (N_2771,N_2525,N_2569);
nor U2772 (N_2772,N_2722,N_2549);
or U2773 (N_2773,N_2627,N_2735);
xnor U2774 (N_2774,N_2526,N_2697);
or U2775 (N_2775,N_2613,N_2705);
nand U2776 (N_2776,N_2620,N_2713);
and U2777 (N_2777,N_2692,N_2647);
nand U2778 (N_2778,N_2651,N_2621);
nor U2779 (N_2779,N_2690,N_2572);
nor U2780 (N_2780,N_2641,N_2561);
xnor U2781 (N_2781,N_2524,N_2673);
nor U2782 (N_2782,N_2563,N_2704);
nor U2783 (N_2783,N_2521,N_2599);
nor U2784 (N_2784,N_2632,N_2625);
nor U2785 (N_2785,N_2614,N_2739);
and U2786 (N_2786,N_2733,N_2514);
nand U2787 (N_2787,N_2646,N_2589);
nand U2788 (N_2788,N_2699,N_2577);
xnor U2789 (N_2789,N_2540,N_2749);
nand U2790 (N_2790,N_2634,N_2725);
and U2791 (N_2791,N_2600,N_2737);
or U2792 (N_2792,N_2709,N_2573);
and U2793 (N_2793,N_2559,N_2567);
and U2794 (N_2794,N_2547,N_2520);
or U2795 (N_2795,N_2578,N_2689);
nor U2796 (N_2796,N_2703,N_2678);
xnor U2797 (N_2797,N_2668,N_2586);
nor U2798 (N_2798,N_2545,N_2653);
xor U2799 (N_2799,N_2698,N_2606);
and U2800 (N_2800,N_2723,N_2745);
and U2801 (N_2801,N_2548,N_2743);
and U2802 (N_2802,N_2591,N_2516);
nor U2803 (N_2803,N_2662,N_2531);
xnor U2804 (N_2804,N_2724,N_2708);
xor U2805 (N_2805,N_2523,N_2552);
or U2806 (N_2806,N_2560,N_2675);
or U2807 (N_2807,N_2718,N_2504);
nor U2808 (N_2808,N_2644,N_2663);
nor U2809 (N_2809,N_2596,N_2574);
and U2810 (N_2810,N_2558,N_2693);
nand U2811 (N_2811,N_2671,N_2710);
or U2812 (N_2812,N_2617,N_2616);
nand U2813 (N_2813,N_2717,N_2636);
and U2814 (N_2814,N_2640,N_2619);
xor U2815 (N_2815,N_2652,N_2684);
and U2816 (N_2816,N_2677,N_2533);
nor U2817 (N_2817,N_2638,N_2682);
or U2818 (N_2818,N_2681,N_2500);
and U2819 (N_2819,N_2714,N_2511);
or U2820 (N_2820,N_2680,N_2611);
and U2821 (N_2821,N_2544,N_2566);
nor U2822 (N_2822,N_2584,N_2637);
nor U2823 (N_2823,N_2601,N_2695);
or U2824 (N_2824,N_2654,N_2656);
nand U2825 (N_2825,N_2635,N_2503);
and U2826 (N_2826,N_2667,N_2562);
nand U2827 (N_2827,N_2659,N_2657);
xor U2828 (N_2828,N_2702,N_2666);
or U2829 (N_2829,N_2679,N_2720);
xnor U2830 (N_2830,N_2691,N_2534);
nor U2831 (N_2831,N_2541,N_2594);
xnor U2832 (N_2832,N_2734,N_2746);
xnor U2833 (N_2833,N_2518,N_2661);
nand U2834 (N_2834,N_2513,N_2658);
and U2835 (N_2835,N_2605,N_2727);
nand U2836 (N_2836,N_2676,N_2665);
or U2837 (N_2837,N_2542,N_2736);
xnor U2838 (N_2838,N_2593,N_2716);
nor U2839 (N_2839,N_2602,N_2701);
nor U2840 (N_2840,N_2512,N_2623);
nand U2841 (N_2841,N_2648,N_2508);
nor U2842 (N_2842,N_2738,N_2696);
xnor U2843 (N_2843,N_2732,N_2674);
nand U2844 (N_2844,N_2587,N_2546);
xor U2845 (N_2845,N_2568,N_2588);
or U2846 (N_2846,N_2685,N_2711);
nand U2847 (N_2847,N_2741,N_2694);
nor U2848 (N_2848,N_2592,N_2728);
nand U2849 (N_2849,N_2532,N_2556);
xor U2850 (N_2850,N_2598,N_2742);
nand U2851 (N_2851,N_2585,N_2645);
nor U2852 (N_2852,N_2555,N_2543);
nor U2853 (N_2853,N_2519,N_2669);
xnor U2854 (N_2854,N_2510,N_2590);
or U2855 (N_2855,N_2748,N_2630);
and U2856 (N_2856,N_2517,N_2506);
xnor U2857 (N_2857,N_2565,N_2576);
or U2858 (N_2858,N_2583,N_2564);
and U2859 (N_2859,N_2570,N_2643);
or U2860 (N_2860,N_2650,N_2553);
or U2861 (N_2861,N_2509,N_2536);
nand U2862 (N_2862,N_2610,N_2507);
and U2863 (N_2863,N_2575,N_2731);
nand U2864 (N_2864,N_2626,N_2607);
and U2865 (N_2865,N_2582,N_2683);
nor U2866 (N_2866,N_2726,N_2655);
nor U2867 (N_2867,N_2664,N_2700);
nor U2868 (N_2868,N_2631,N_2571);
nand U2869 (N_2869,N_2660,N_2530);
nor U2870 (N_2870,N_2529,N_2744);
xor U2871 (N_2871,N_2707,N_2670);
xor U2872 (N_2872,N_2537,N_2612);
or U2873 (N_2873,N_2539,N_2550);
nor U2874 (N_2874,N_2730,N_2712);
nand U2875 (N_2875,N_2566,N_2681);
nand U2876 (N_2876,N_2711,N_2603);
nor U2877 (N_2877,N_2683,N_2550);
nor U2878 (N_2878,N_2701,N_2620);
nand U2879 (N_2879,N_2725,N_2722);
xor U2880 (N_2880,N_2542,N_2682);
or U2881 (N_2881,N_2617,N_2612);
nand U2882 (N_2882,N_2583,N_2556);
nor U2883 (N_2883,N_2504,N_2603);
and U2884 (N_2884,N_2707,N_2500);
nand U2885 (N_2885,N_2511,N_2680);
nor U2886 (N_2886,N_2742,N_2531);
or U2887 (N_2887,N_2602,N_2704);
xnor U2888 (N_2888,N_2597,N_2717);
xnor U2889 (N_2889,N_2600,N_2736);
and U2890 (N_2890,N_2622,N_2716);
or U2891 (N_2891,N_2578,N_2542);
and U2892 (N_2892,N_2535,N_2657);
xor U2893 (N_2893,N_2600,N_2627);
nand U2894 (N_2894,N_2653,N_2507);
and U2895 (N_2895,N_2593,N_2530);
xnor U2896 (N_2896,N_2640,N_2515);
and U2897 (N_2897,N_2704,N_2588);
nor U2898 (N_2898,N_2702,N_2565);
and U2899 (N_2899,N_2505,N_2722);
nand U2900 (N_2900,N_2519,N_2526);
nand U2901 (N_2901,N_2633,N_2681);
nand U2902 (N_2902,N_2552,N_2608);
or U2903 (N_2903,N_2730,N_2718);
and U2904 (N_2904,N_2697,N_2520);
or U2905 (N_2905,N_2555,N_2678);
or U2906 (N_2906,N_2609,N_2637);
or U2907 (N_2907,N_2568,N_2671);
nor U2908 (N_2908,N_2598,N_2549);
xor U2909 (N_2909,N_2647,N_2657);
xnor U2910 (N_2910,N_2618,N_2592);
xnor U2911 (N_2911,N_2583,N_2522);
and U2912 (N_2912,N_2628,N_2622);
and U2913 (N_2913,N_2699,N_2646);
nand U2914 (N_2914,N_2577,N_2608);
xnor U2915 (N_2915,N_2627,N_2530);
nor U2916 (N_2916,N_2696,N_2673);
nand U2917 (N_2917,N_2660,N_2619);
and U2918 (N_2918,N_2688,N_2700);
and U2919 (N_2919,N_2655,N_2747);
xnor U2920 (N_2920,N_2598,N_2592);
nand U2921 (N_2921,N_2667,N_2508);
or U2922 (N_2922,N_2507,N_2699);
xor U2923 (N_2923,N_2646,N_2577);
nand U2924 (N_2924,N_2632,N_2692);
or U2925 (N_2925,N_2550,N_2526);
xor U2926 (N_2926,N_2696,N_2603);
or U2927 (N_2927,N_2578,N_2715);
or U2928 (N_2928,N_2530,N_2549);
nand U2929 (N_2929,N_2738,N_2735);
nand U2930 (N_2930,N_2632,N_2549);
or U2931 (N_2931,N_2506,N_2668);
xor U2932 (N_2932,N_2715,N_2529);
xor U2933 (N_2933,N_2600,N_2524);
nor U2934 (N_2934,N_2690,N_2503);
nand U2935 (N_2935,N_2706,N_2555);
or U2936 (N_2936,N_2692,N_2606);
xor U2937 (N_2937,N_2735,N_2631);
nand U2938 (N_2938,N_2532,N_2720);
nor U2939 (N_2939,N_2636,N_2673);
nor U2940 (N_2940,N_2717,N_2675);
or U2941 (N_2941,N_2728,N_2505);
and U2942 (N_2942,N_2570,N_2555);
and U2943 (N_2943,N_2588,N_2555);
nor U2944 (N_2944,N_2703,N_2611);
or U2945 (N_2945,N_2643,N_2673);
or U2946 (N_2946,N_2577,N_2706);
and U2947 (N_2947,N_2508,N_2724);
xor U2948 (N_2948,N_2572,N_2651);
nand U2949 (N_2949,N_2615,N_2509);
and U2950 (N_2950,N_2728,N_2534);
or U2951 (N_2951,N_2511,N_2638);
nand U2952 (N_2952,N_2670,N_2679);
nand U2953 (N_2953,N_2747,N_2520);
nand U2954 (N_2954,N_2529,N_2542);
or U2955 (N_2955,N_2731,N_2617);
xnor U2956 (N_2956,N_2711,N_2700);
or U2957 (N_2957,N_2528,N_2555);
or U2958 (N_2958,N_2703,N_2554);
nor U2959 (N_2959,N_2687,N_2591);
nor U2960 (N_2960,N_2743,N_2704);
xnor U2961 (N_2961,N_2582,N_2639);
and U2962 (N_2962,N_2524,N_2552);
or U2963 (N_2963,N_2539,N_2589);
nand U2964 (N_2964,N_2635,N_2671);
xnor U2965 (N_2965,N_2516,N_2691);
xnor U2966 (N_2966,N_2648,N_2545);
and U2967 (N_2967,N_2529,N_2653);
xor U2968 (N_2968,N_2519,N_2645);
or U2969 (N_2969,N_2590,N_2678);
nor U2970 (N_2970,N_2594,N_2643);
and U2971 (N_2971,N_2743,N_2533);
nor U2972 (N_2972,N_2520,N_2517);
and U2973 (N_2973,N_2579,N_2500);
or U2974 (N_2974,N_2688,N_2663);
nand U2975 (N_2975,N_2528,N_2640);
and U2976 (N_2976,N_2595,N_2631);
nand U2977 (N_2977,N_2541,N_2612);
nand U2978 (N_2978,N_2651,N_2684);
nand U2979 (N_2979,N_2599,N_2602);
and U2980 (N_2980,N_2650,N_2723);
xnor U2981 (N_2981,N_2730,N_2662);
and U2982 (N_2982,N_2506,N_2564);
xor U2983 (N_2983,N_2638,N_2698);
nand U2984 (N_2984,N_2544,N_2584);
and U2985 (N_2985,N_2736,N_2529);
or U2986 (N_2986,N_2600,N_2569);
xnor U2987 (N_2987,N_2548,N_2633);
xor U2988 (N_2988,N_2608,N_2612);
and U2989 (N_2989,N_2652,N_2659);
and U2990 (N_2990,N_2551,N_2586);
nor U2991 (N_2991,N_2669,N_2514);
nand U2992 (N_2992,N_2514,N_2506);
xnor U2993 (N_2993,N_2616,N_2545);
nand U2994 (N_2994,N_2702,N_2688);
xnor U2995 (N_2995,N_2593,N_2746);
xor U2996 (N_2996,N_2697,N_2739);
nor U2997 (N_2997,N_2682,N_2512);
xnor U2998 (N_2998,N_2551,N_2683);
nand U2999 (N_2999,N_2529,N_2686);
and U3000 (N_3000,N_2832,N_2751);
nand U3001 (N_3001,N_2861,N_2798);
nor U3002 (N_3002,N_2962,N_2789);
xor U3003 (N_3003,N_2944,N_2800);
or U3004 (N_3004,N_2872,N_2860);
nand U3005 (N_3005,N_2884,N_2986);
and U3006 (N_3006,N_2893,N_2938);
or U3007 (N_3007,N_2994,N_2768);
and U3008 (N_3008,N_2972,N_2996);
and U3009 (N_3009,N_2999,N_2912);
nor U3010 (N_3010,N_2858,N_2982);
xor U3011 (N_3011,N_2917,N_2787);
nand U3012 (N_3012,N_2937,N_2752);
or U3013 (N_3013,N_2911,N_2891);
or U3014 (N_3014,N_2920,N_2910);
nor U3015 (N_3015,N_2955,N_2969);
xnor U3016 (N_3016,N_2892,N_2881);
nor U3017 (N_3017,N_2859,N_2878);
xnor U3018 (N_3018,N_2974,N_2846);
nor U3019 (N_3019,N_2983,N_2809);
or U3020 (N_3020,N_2845,N_2890);
and U3021 (N_3021,N_2755,N_2896);
and U3022 (N_3022,N_2762,N_2791);
xnor U3023 (N_3023,N_2954,N_2781);
and U3024 (N_3024,N_2792,N_2788);
nor U3025 (N_3025,N_2810,N_2801);
nand U3026 (N_3026,N_2818,N_2807);
or U3027 (N_3027,N_2750,N_2942);
or U3028 (N_3028,N_2922,N_2841);
and U3029 (N_3029,N_2965,N_2867);
xor U3030 (N_3030,N_2831,N_2899);
xnor U3031 (N_3031,N_2772,N_2963);
nand U3032 (N_3032,N_2812,N_2855);
nand U3033 (N_3033,N_2784,N_2977);
and U3034 (N_3034,N_2829,N_2838);
nor U3035 (N_3035,N_2756,N_2853);
nand U3036 (N_3036,N_2978,N_2825);
nor U3037 (N_3037,N_2925,N_2758);
nand U3038 (N_3038,N_2946,N_2952);
and U3039 (N_3039,N_2975,N_2900);
nand U3040 (N_3040,N_2786,N_2826);
xnor U3041 (N_3041,N_2988,N_2868);
or U3042 (N_3042,N_2980,N_2927);
and U3043 (N_3043,N_2813,N_2840);
xor U3044 (N_3044,N_2847,N_2987);
xor U3045 (N_3045,N_2875,N_2779);
nand U3046 (N_3046,N_2761,N_2770);
nor U3047 (N_3047,N_2759,N_2764);
nand U3048 (N_3048,N_2997,N_2869);
xnor U3049 (N_3049,N_2828,N_2909);
nor U3050 (N_3050,N_2913,N_2834);
nor U3051 (N_3051,N_2908,N_2971);
xor U3052 (N_3052,N_2802,N_2760);
nand U3053 (N_3053,N_2928,N_2814);
and U3054 (N_3054,N_2990,N_2794);
and U3055 (N_3055,N_2961,N_2943);
or U3056 (N_3056,N_2901,N_2919);
xnor U3057 (N_3057,N_2763,N_2898);
nand U3058 (N_3058,N_2870,N_2929);
xor U3059 (N_3059,N_2803,N_2866);
or U3060 (N_3060,N_2836,N_2904);
nand U3061 (N_3061,N_2851,N_2811);
and U3062 (N_3062,N_2765,N_2777);
xor U3063 (N_3063,N_2776,N_2864);
nand U3064 (N_3064,N_2848,N_2796);
and U3065 (N_3065,N_2822,N_2985);
or U3066 (N_3066,N_2981,N_2865);
and U3067 (N_3067,N_2992,N_2854);
nor U3068 (N_3068,N_2808,N_2973);
nor U3069 (N_3069,N_2905,N_2902);
or U3070 (N_3070,N_2939,N_2766);
nor U3071 (N_3071,N_2993,N_2880);
or U3072 (N_3072,N_2856,N_2903);
xnor U3073 (N_3073,N_2767,N_2918);
xnor U3074 (N_3074,N_2976,N_2871);
or U3075 (N_3075,N_2995,N_2885);
or U3076 (N_3076,N_2849,N_2835);
xnor U3077 (N_3077,N_2979,N_2966);
and U3078 (N_3078,N_2916,N_2863);
xor U3079 (N_3079,N_2959,N_2793);
nor U3080 (N_3080,N_2876,N_2753);
and U3081 (N_3081,N_2757,N_2940);
nor U3082 (N_3082,N_2956,N_2821);
nand U3083 (N_3083,N_2921,N_2941);
and U3084 (N_3084,N_2887,N_2957);
nand U3085 (N_3085,N_2850,N_2797);
or U3086 (N_3086,N_2783,N_2931);
nor U3087 (N_3087,N_2970,N_2837);
nor U3088 (N_3088,N_2960,N_2948);
and U3089 (N_3089,N_2819,N_2895);
or U3090 (N_3090,N_2926,N_2778);
nor U3091 (N_3091,N_2806,N_2873);
or U3092 (N_3092,N_2795,N_2804);
and U3093 (N_3093,N_2799,N_2950);
xnor U3094 (N_3094,N_2894,N_2949);
and U3095 (N_3095,N_2827,N_2935);
nand U3096 (N_3096,N_2923,N_2879);
nand U3097 (N_3097,N_2889,N_2888);
or U3098 (N_3098,N_2930,N_2882);
nor U3099 (N_3099,N_2945,N_2790);
nand U3100 (N_3100,N_2886,N_2958);
nand U3101 (N_3101,N_2775,N_2843);
or U3102 (N_3102,N_2947,N_2936);
or U3103 (N_3103,N_2857,N_2915);
nand U3104 (N_3104,N_2914,N_2924);
nor U3105 (N_3105,N_2805,N_2780);
or U3106 (N_3106,N_2824,N_2816);
or U3107 (N_3107,N_2933,N_2842);
nand U3108 (N_3108,N_2967,N_2771);
nor U3109 (N_3109,N_2754,N_2830);
nand U3110 (N_3110,N_2862,N_2823);
nand U3111 (N_3111,N_2964,N_2906);
nor U3112 (N_3112,N_2951,N_2844);
nand U3113 (N_3113,N_2883,N_2897);
or U3114 (N_3114,N_2815,N_2839);
nor U3115 (N_3115,N_2782,N_2932);
nand U3116 (N_3116,N_2989,N_2785);
nor U3117 (N_3117,N_2953,N_2907);
nand U3118 (N_3118,N_2968,N_2774);
and U3119 (N_3119,N_2874,N_2984);
or U3120 (N_3120,N_2833,N_2817);
and U3121 (N_3121,N_2877,N_2852);
nor U3122 (N_3122,N_2769,N_2934);
nor U3123 (N_3123,N_2773,N_2991);
nand U3124 (N_3124,N_2820,N_2998);
nor U3125 (N_3125,N_2844,N_2974);
nand U3126 (N_3126,N_2761,N_2806);
nor U3127 (N_3127,N_2871,N_2828);
or U3128 (N_3128,N_2818,N_2795);
nand U3129 (N_3129,N_2897,N_2893);
or U3130 (N_3130,N_2872,N_2883);
nand U3131 (N_3131,N_2758,N_2764);
xnor U3132 (N_3132,N_2949,N_2877);
nor U3133 (N_3133,N_2864,N_2977);
nand U3134 (N_3134,N_2976,N_2891);
nand U3135 (N_3135,N_2964,N_2938);
nor U3136 (N_3136,N_2903,N_2797);
or U3137 (N_3137,N_2803,N_2870);
nor U3138 (N_3138,N_2803,N_2901);
or U3139 (N_3139,N_2771,N_2917);
or U3140 (N_3140,N_2971,N_2913);
nor U3141 (N_3141,N_2810,N_2775);
or U3142 (N_3142,N_2895,N_2830);
or U3143 (N_3143,N_2934,N_2898);
nand U3144 (N_3144,N_2835,N_2881);
or U3145 (N_3145,N_2821,N_2765);
or U3146 (N_3146,N_2773,N_2752);
nor U3147 (N_3147,N_2759,N_2877);
nand U3148 (N_3148,N_2995,N_2806);
nor U3149 (N_3149,N_2784,N_2802);
nand U3150 (N_3150,N_2994,N_2912);
and U3151 (N_3151,N_2855,N_2880);
or U3152 (N_3152,N_2892,N_2918);
and U3153 (N_3153,N_2921,N_2987);
nand U3154 (N_3154,N_2828,N_2851);
and U3155 (N_3155,N_2798,N_2878);
and U3156 (N_3156,N_2793,N_2978);
nor U3157 (N_3157,N_2841,N_2881);
or U3158 (N_3158,N_2790,N_2828);
and U3159 (N_3159,N_2945,N_2886);
and U3160 (N_3160,N_2806,N_2773);
and U3161 (N_3161,N_2976,N_2797);
nor U3162 (N_3162,N_2880,N_2866);
and U3163 (N_3163,N_2976,N_2905);
nor U3164 (N_3164,N_2879,N_2976);
nand U3165 (N_3165,N_2999,N_2987);
and U3166 (N_3166,N_2843,N_2938);
nor U3167 (N_3167,N_2879,N_2874);
or U3168 (N_3168,N_2816,N_2993);
nor U3169 (N_3169,N_2779,N_2790);
or U3170 (N_3170,N_2797,N_2985);
nor U3171 (N_3171,N_2798,N_2928);
or U3172 (N_3172,N_2804,N_2944);
nand U3173 (N_3173,N_2848,N_2847);
xnor U3174 (N_3174,N_2771,N_2956);
xnor U3175 (N_3175,N_2888,N_2970);
or U3176 (N_3176,N_2776,N_2995);
nor U3177 (N_3177,N_2760,N_2998);
xnor U3178 (N_3178,N_2774,N_2772);
and U3179 (N_3179,N_2888,N_2851);
and U3180 (N_3180,N_2931,N_2899);
and U3181 (N_3181,N_2858,N_2884);
and U3182 (N_3182,N_2825,N_2880);
nand U3183 (N_3183,N_2803,N_2775);
nand U3184 (N_3184,N_2797,N_2894);
or U3185 (N_3185,N_2873,N_2821);
xnor U3186 (N_3186,N_2977,N_2758);
and U3187 (N_3187,N_2918,N_2819);
nor U3188 (N_3188,N_2932,N_2924);
xnor U3189 (N_3189,N_2954,N_2784);
xnor U3190 (N_3190,N_2823,N_2854);
and U3191 (N_3191,N_2889,N_2861);
or U3192 (N_3192,N_2846,N_2786);
nand U3193 (N_3193,N_2793,N_2815);
and U3194 (N_3194,N_2859,N_2835);
nor U3195 (N_3195,N_2924,N_2935);
and U3196 (N_3196,N_2980,N_2907);
and U3197 (N_3197,N_2797,N_2858);
xor U3198 (N_3198,N_2960,N_2907);
nand U3199 (N_3199,N_2915,N_2938);
and U3200 (N_3200,N_2827,N_2982);
nor U3201 (N_3201,N_2919,N_2757);
or U3202 (N_3202,N_2954,N_2947);
and U3203 (N_3203,N_2906,N_2942);
xnor U3204 (N_3204,N_2887,N_2874);
nand U3205 (N_3205,N_2785,N_2958);
nand U3206 (N_3206,N_2985,N_2837);
nand U3207 (N_3207,N_2869,N_2965);
nand U3208 (N_3208,N_2890,N_2865);
xnor U3209 (N_3209,N_2782,N_2893);
xnor U3210 (N_3210,N_2921,N_2864);
or U3211 (N_3211,N_2918,N_2853);
nand U3212 (N_3212,N_2879,N_2961);
nor U3213 (N_3213,N_2789,N_2966);
nand U3214 (N_3214,N_2882,N_2826);
or U3215 (N_3215,N_2935,N_2971);
nand U3216 (N_3216,N_2972,N_2816);
nor U3217 (N_3217,N_2868,N_2991);
xor U3218 (N_3218,N_2937,N_2992);
nand U3219 (N_3219,N_2998,N_2906);
nand U3220 (N_3220,N_2760,N_2755);
nor U3221 (N_3221,N_2930,N_2767);
or U3222 (N_3222,N_2966,N_2802);
xnor U3223 (N_3223,N_2852,N_2808);
and U3224 (N_3224,N_2790,N_2885);
xnor U3225 (N_3225,N_2843,N_2842);
xnor U3226 (N_3226,N_2809,N_2887);
and U3227 (N_3227,N_2764,N_2878);
or U3228 (N_3228,N_2835,N_2761);
xor U3229 (N_3229,N_2857,N_2940);
or U3230 (N_3230,N_2876,N_2889);
and U3231 (N_3231,N_2982,N_2823);
xor U3232 (N_3232,N_2941,N_2938);
and U3233 (N_3233,N_2959,N_2964);
xor U3234 (N_3234,N_2839,N_2754);
or U3235 (N_3235,N_2918,N_2917);
and U3236 (N_3236,N_2863,N_2774);
or U3237 (N_3237,N_2794,N_2877);
xor U3238 (N_3238,N_2994,N_2838);
or U3239 (N_3239,N_2919,N_2881);
and U3240 (N_3240,N_2899,N_2945);
and U3241 (N_3241,N_2765,N_2752);
and U3242 (N_3242,N_2895,N_2922);
nand U3243 (N_3243,N_2939,N_2795);
nor U3244 (N_3244,N_2821,N_2755);
or U3245 (N_3245,N_2802,N_2819);
and U3246 (N_3246,N_2870,N_2776);
and U3247 (N_3247,N_2881,N_2828);
xor U3248 (N_3248,N_2927,N_2916);
xnor U3249 (N_3249,N_2871,N_2972);
nand U3250 (N_3250,N_3002,N_3005);
nor U3251 (N_3251,N_3077,N_3138);
nor U3252 (N_3252,N_3024,N_3240);
nand U3253 (N_3253,N_3091,N_3196);
nand U3254 (N_3254,N_3226,N_3137);
nand U3255 (N_3255,N_3007,N_3067);
and U3256 (N_3256,N_3117,N_3123);
and U3257 (N_3257,N_3103,N_3026);
nand U3258 (N_3258,N_3035,N_3139);
xor U3259 (N_3259,N_3092,N_3175);
nor U3260 (N_3260,N_3183,N_3159);
or U3261 (N_3261,N_3191,N_3168);
nand U3262 (N_3262,N_3048,N_3185);
nand U3263 (N_3263,N_3144,N_3225);
xnor U3264 (N_3264,N_3165,N_3058);
or U3265 (N_3265,N_3065,N_3025);
nor U3266 (N_3266,N_3131,N_3179);
nor U3267 (N_3267,N_3201,N_3006);
xor U3268 (N_3268,N_3095,N_3083);
xnor U3269 (N_3269,N_3021,N_3224);
xor U3270 (N_3270,N_3173,N_3228);
or U3271 (N_3271,N_3051,N_3190);
and U3272 (N_3272,N_3090,N_3038);
nor U3273 (N_3273,N_3081,N_3204);
nor U3274 (N_3274,N_3187,N_3116);
nand U3275 (N_3275,N_3040,N_3106);
xnor U3276 (N_3276,N_3064,N_3189);
or U3277 (N_3277,N_3218,N_3184);
nand U3278 (N_3278,N_3246,N_3219);
xor U3279 (N_3279,N_3162,N_3200);
nor U3280 (N_3280,N_3122,N_3133);
nor U3281 (N_3281,N_3163,N_3244);
nor U3282 (N_3282,N_3015,N_3094);
or U3283 (N_3283,N_3020,N_3109);
nand U3284 (N_3284,N_3205,N_3132);
nand U3285 (N_3285,N_3032,N_3172);
or U3286 (N_3286,N_3161,N_3096);
nand U3287 (N_3287,N_3030,N_3154);
or U3288 (N_3288,N_3059,N_3121);
xnor U3289 (N_3289,N_3164,N_3008);
and U3290 (N_3290,N_3014,N_3055);
and U3291 (N_3291,N_3199,N_3045);
nand U3292 (N_3292,N_3243,N_3232);
nand U3293 (N_3293,N_3241,N_3118);
nand U3294 (N_3294,N_3155,N_3156);
nand U3295 (N_3295,N_3171,N_3076);
and U3296 (N_3296,N_3247,N_3061);
nand U3297 (N_3297,N_3223,N_3198);
or U3298 (N_3298,N_3071,N_3010);
or U3299 (N_3299,N_3003,N_3146);
xnor U3300 (N_3300,N_3149,N_3042);
nand U3301 (N_3301,N_3220,N_3099);
nor U3302 (N_3302,N_3158,N_3078);
xnor U3303 (N_3303,N_3097,N_3129);
nand U3304 (N_3304,N_3239,N_3105);
or U3305 (N_3305,N_3115,N_3028);
xnor U3306 (N_3306,N_3195,N_3249);
nor U3307 (N_3307,N_3069,N_3217);
nor U3308 (N_3308,N_3233,N_3027);
xor U3309 (N_3309,N_3160,N_3011);
and U3310 (N_3310,N_3231,N_3093);
or U3311 (N_3311,N_3114,N_3018);
or U3312 (N_3312,N_3031,N_3230);
nand U3313 (N_3313,N_3192,N_3221);
or U3314 (N_3314,N_3053,N_3056);
or U3315 (N_3315,N_3029,N_3178);
and U3316 (N_3316,N_3214,N_3110);
nand U3317 (N_3317,N_3216,N_3101);
and U3318 (N_3318,N_3147,N_3148);
and U3319 (N_3319,N_3111,N_3215);
and U3320 (N_3320,N_3066,N_3124);
nand U3321 (N_3321,N_3211,N_3000);
nor U3322 (N_3322,N_3054,N_3033);
nand U3323 (N_3323,N_3227,N_3125);
or U3324 (N_3324,N_3074,N_3188);
or U3325 (N_3325,N_3229,N_3052);
xnor U3326 (N_3326,N_3100,N_3242);
and U3327 (N_3327,N_3120,N_3238);
nand U3328 (N_3328,N_3167,N_3085);
and U3329 (N_3329,N_3142,N_3210);
nand U3330 (N_3330,N_3012,N_3169);
nor U3331 (N_3331,N_3203,N_3212);
and U3332 (N_3332,N_3208,N_3235);
xnor U3333 (N_3333,N_3108,N_3022);
nor U3334 (N_3334,N_3050,N_3222);
nand U3335 (N_3335,N_3170,N_3176);
and U3336 (N_3336,N_3072,N_3174);
or U3337 (N_3337,N_3209,N_3039);
xnor U3338 (N_3338,N_3127,N_3107);
xnor U3339 (N_3339,N_3043,N_3016);
and U3340 (N_3340,N_3166,N_3062);
nor U3341 (N_3341,N_3152,N_3234);
nand U3342 (N_3342,N_3023,N_3060);
nor U3343 (N_3343,N_3143,N_3180);
nor U3344 (N_3344,N_3041,N_3136);
nand U3345 (N_3345,N_3134,N_3181);
and U3346 (N_3346,N_3151,N_3145);
and U3347 (N_3347,N_3248,N_3034);
and U3348 (N_3348,N_3186,N_3036);
or U3349 (N_3349,N_3202,N_3130);
xnor U3350 (N_3350,N_3084,N_3073);
nand U3351 (N_3351,N_3206,N_3213);
and U3352 (N_3352,N_3082,N_3098);
xor U3353 (N_3353,N_3044,N_3089);
and U3354 (N_3354,N_3126,N_3150);
nor U3355 (N_3355,N_3237,N_3070);
nor U3356 (N_3356,N_3087,N_3207);
nor U3357 (N_3357,N_3017,N_3019);
xor U3358 (N_3358,N_3088,N_3037);
or U3359 (N_3359,N_3135,N_3153);
or U3360 (N_3360,N_3057,N_3113);
and U3361 (N_3361,N_3112,N_3049);
and U3362 (N_3362,N_3177,N_3086);
and U3363 (N_3363,N_3009,N_3080);
nor U3364 (N_3364,N_3140,N_3079);
nand U3365 (N_3365,N_3013,N_3004);
and U3366 (N_3366,N_3102,N_3075);
or U3367 (N_3367,N_3001,N_3063);
nand U3368 (N_3368,N_3157,N_3047);
or U3369 (N_3369,N_3046,N_3197);
or U3370 (N_3370,N_3236,N_3104);
nand U3371 (N_3371,N_3182,N_3193);
or U3372 (N_3372,N_3068,N_3245);
and U3373 (N_3373,N_3119,N_3194);
and U3374 (N_3374,N_3128,N_3141);
or U3375 (N_3375,N_3230,N_3087);
nand U3376 (N_3376,N_3135,N_3174);
nor U3377 (N_3377,N_3064,N_3083);
xnor U3378 (N_3378,N_3137,N_3089);
xor U3379 (N_3379,N_3121,N_3187);
nand U3380 (N_3380,N_3166,N_3164);
xnor U3381 (N_3381,N_3156,N_3090);
nand U3382 (N_3382,N_3035,N_3141);
nand U3383 (N_3383,N_3179,N_3240);
nand U3384 (N_3384,N_3031,N_3246);
or U3385 (N_3385,N_3033,N_3146);
nand U3386 (N_3386,N_3129,N_3125);
and U3387 (N_3387,N_3162,N_3201);
and U3388 (N_3388,N_3095,N_3165);
nand U3389 (N_3389,N_3157,N_3159);
nor U3390 (N_3390,N_3126,N_3073);
nand U3391 (N_3391,N_3153,N_3025);
and U3392 (N_3392,N_3168,N_3209);
nor U3393 (N_3393,N_3007,N_3232);
nor U3394 (N_3394,N_3002,N_3033);
and U3395 (N_3395,N_3131,N_3147);
and U3396 (N_3396,N_3115,N_3167);
and U3397 (N_3397,N_3194,N_3176);
nand U3398 (N_3398,N_3247,N_3121);
nand U3399 (N_3399,N_3211,N_3113);
nor U3400 (N_3400,N_3093,N_3195);
nor U3401 (N_3401,N_3180,N_3130);
and U3402 (N_3402,N_3233,N_3123);
xnor U3403 (N_3403,N_3204,N_3158);
xor U3404 (N_3404,N_3168,N_3158);
and U3405 (N_3405,N_3007,N_3081);
xnor U3406 (N_3406,N_3195,N_3118);
or U3407 (N_3407,N_3197,N_3163);
nor U3408 (N_3408,N_3024,N_3103);
nand U3409 (N_3409,N_3150,N_3184);
or U3410 (N_3410,N_3199,N_3023);
or U3411 (N_3411,N_3121,N_3111);
xnor U3412 (N_3412,N_3170,N_3056);
xnor U3413 (N_3413,N_3185,N_3071);
and U3414 (N_3414,N_3237,N_3208);
nor U3415 (N_3415,N_3214,N_3239);
nor U3416 (N_3416,N_3060,N_3215);
and U3417 (N_3417,N_3190,N_3189);
or U3418 (N_3418,N_3036,N_3096);
nor U3419 (N_3419,N_3174,N_3223);
xor U3420 (N_3420,N_3079,N_3014);
xor U3421 (N_3421,N_3044,N_3066);
and U3422 (N_3422,N_3098,N_3167);
nor U3423 (N_3423,N_3242,N_3173);
and U3424 (N_3424,N_3198,N_3079);
nor U3425 (N_3425,N_3107,N_3016);
nor U3426 (N_3426,N_3239,N_3155);
nor U3427 (N_3427,N_3186,N_3224);
xor U3428 (N_3428,N_3039,N_3096);
and U3429 (N_3429,N_3194,N_3160);
nor U3430 (N_3430,N_3042,N_3236);
nor U3431 (N_3431,N_3040,N_3213);
nand U3432 (N_3432,N_3206,N_3207);
xor U3433 (N_3433,N_3186,N_3010);
nand U3434 (N_3434,N_3052,N_3145);
xor U3435 (N_3435,N_3050,N_3066);
nor U3436 (N_3436,N_3247,N_3067);
nand U3437 (N_3437,N_3011,N_3047);
and U3438 (N_3438,N_3195,N_3211);
nand U3439 (N_3439,N_3020,N_3136);
and U3440 (N_3440,N_3151,N_3137);
nand U3441 (N_3441,N_3174,N_3133);
xnor U3442 (N_3442,N_3083,N_3012);
and U3443 (N_3443,N_3156,N_3127);
and U3444 (N_3444,N_3081,N_3210);
nor U3445 (N_3445,N_3053,N_3049);
or U3446 (N_3446,N_3242,N_3215);
nor U3447 (N_3447,N_3046,N_3126);
or U3448 (N_3448,N_3210,N_3034);
nand U3449 (N_3449,N_3066,N_3215);
xor U3450 (N_3450,N_3210,N_3063);
nor U3451 (N_3451,N_3122,N_3153);
and U3452 (N_3452,N_3201,N_3088);
nor U3453 (N_3453,N_3128,N_3196);
nand U3454 (N_3454,N_3161,N_3201);
xnor U3455 (N_3455,N_3168,N_3060);
nor U3456 (N_3456,N_3008,N_3137);
and U3457 (N_3457,N_3003,N_3212);
or U3458 (N_3458,N_3040,N_3070);
and U3459 (N_3459,N_3025,N_3074);
and U3460 (N_3460,N_3008,N_3146);
or U3461 (N_3461,N_3199,N_3212);
and U3462 (N_3462,N_3117,N_3036);
and U3463 (N_3463,N_3025,N_3102);
nand U3464 (N_3464,N_3108,N_3165);
xor U3465 (N_3465,N_3235,N_3242);
and U3466 (N_3466,N_3191,N_3144);
xnor U3467 (N_3467,N_3245,N_3161);
xor U3468 (N_3468,N_3112,N_3127);
and U3469 (N_3469,N_3153,N_3220);
xnor U3470 (N_3470,N_3096,N_3166);
xor U3471 (N_3471,N_3118,N_3204);
and U3472 (N_3472,N_3201,N_3155);
xnor U3473 (N_3473,N_3180,N_3114);
nor U3474 (N_3474,N_3018,N_3209);
and U3475 (N_3475,N_3005,N_3150);
xnor U3476 (N_3476,N_3193,N_3156);
and U3477 (N_3477,N_3047,N_3153);
or U3478 (N_3478,N_3169,N_3249);
and U3479 (N_3479,N_3187,N_3243);
and U3480 (N_3480,N_3006,N_3025);
or U3481 (N_3481,N_3160,N_3249);
xor U3482 (N_3482,N_3039,N_3234);
or U3483 (N_3483,N_3233,N_3051);
nand U3484 (N_3484,N_3151,N_3212);
or U3485 (N_3485,N_3106,N_3186);
xor U3486 (N_3486,N_3164,N_3046);
or U3487 (N_3487,N_3049,N_3171);
nand U3488 (N_3488,N_3233,N_3150);
nor U3489 (N_3489,N_3120,N_3131);
and U3490 (N_3490,N_3089,N_3051);
xor U3491 (N_3491,N_3021,N_3172);
or U3492 (N_3492,N_3150,N_3165);
nor U3493 (N_3493,N_3180,N_3034);
or U3494 (N_3494,N_3144,N_3190);
nor U3495 (N_3495,N_3248,N_3002);
nand U3496 (N_3496,N_3038,N_3062);
and U3497 (N_3497,N_3131,N_3167);
or U3498 (N_3498,N_3162,N_3026);
nand U3499 (N_3499,N_3162,N_3022);
nor U3500 (N_3500,N_3298,N_3471);
nand U3501 (N_3501,N_3417,N_3337);
or U3502 (N_3502,N_3458,N_3357);
and U3503 (N_3503,N_3279,N_3489);
nor U3504 (N_3504,N_3349,N_3327);
or U3505 (N_3505,N_3455,N_3361);
nor U3506 (N_3506,N_3449,N_3414);
and U3507 (N_3507,N_3469,N_3320);
nor U3508 (N_3508,N_3391,N_3396);
xnor U3509 (N_3509,N_3368,N_3321);
xnor U3510 (N_3510,N_3313,N_3369);
and U3511 (N_3511,N_3392,N_3304);
or U3512 (N_3512,N_3460,N_3477);
and U3513 (N_3513,N_3302,N_3328);
nor U3514 (N_3514,N_3345,N_3448);
nor U3515 (N_3515,N_3370,N_3467);
xor U3516 (N_3516,N_3453,N_3277);
nand U3517 (N_3517,N_3492,N_3332);
nor U3518 (N_3518,N_3338,N_3404);
xnor U3519 (N_3519,N_3436,N_3483);
and U3520 (N_3520,N_3331,N_3284);
nor U3521 (N_3521,N_3346,N_3254);
xor U3522 (N_3522,N_3476,N_3330);
and U3523 (N_3523,N_3408,N_3275);
xor U3524 (N_3524,N_3442,N_3428);
xnor U3525 (N_3525,N_3461,N_3423);
xor U3526 (N_3526,N_3497,N_3433);
nand U3527 (N_3527,N_3441,N_3339);
and U3528 (N_3528,N_3389,N_3367);
nor U3529 (N_3529,N_3488,N_3409);
nand U3530 (N_3530,N_3253,N_3474);
xnor U3531 (N_3531,N_3486,N_3324);
nand U3532 (N_3532,N_3435,N_3491);
and U3533 (N_3533,N_3341,N_3424);
nand U3534 (N_3534,N_3494,N_3329);
or U3535 (N_3535,N_3293,N_3401);
xor U3536 (N_3536,N_3388,N_3490);
or U3537 (N_3537,N_3355,N_3358);
and U3538 (N_3538,N_3462,N_3382);
xnor U3539 (N_3539,N_3451,N_3323);
xor U3540 (N_3540,N_3271,N_3410);
or U3541 (N_3541,N_3250,N_3305);
nand U3542 (N_3542,N_3282,N_3457);
xnor U3543 (N_3543,N_3289,N_3482);
nor U3544 (N_3544,N_3257,N_3265);
nand U3545 (N_3545,N_3336,N_3485);
nor U3546 (N_3546,N_3438,N_3278);
xnor U3547 (N_3547,N_3283,N_3333);
or U3548 (N_3548,N_3466,N_3405);
and U3549 (N_3549,N_3463,N_3294);
nor U3550 (N_3550,N_3312,N_3495);
and U3551 (N_3551,N_3344,N_3267);
or U3552 (N_3552,N_3400,N_3286);
or U3553 (N_3553,N_3356,N_3398);
and U3554 (N_3554,N_3266,N_3383);
xnor U3555 (N_3555,N_3459,N_3385);
or U3556 (N_3556,N_3261,N_3372);
xor U3557 (N_3557,N_3454,N_3430);
nor U3558 (N_3558,N_3319,N_3412);
xor U3559 (N_3559,N_3413,N_3262);
nand U3560 (N_3560,N_3285,N_3465);
xnor U3561 (N_3561,N_3443,N_3363);
nor U3562 (N_3562,N_3380,N_3445);
nor U3563 (N_3563,N_3348,N_3342);
or U3564 (N_3564,N_3386,N_3468);
nor U3565 (N_3565,N_3281,N_3420);
nand U3566 (N_3566,N_3418,N_3373);
xor U3567 (N_3567,N_3411,N_3354);
nor U3568 (N_3568,N_3437,N_3446);
or U3569 (N_3569,N_3264,N_3310);
xnor U3570 (N_3570,N_3326,N_3499);
xnor U3571 (N_3571,N_3416,N_3475);
nor U3572 (N_3572,N_3447,N_3340);
nand U3573 (N_3573,N_3350,N_3307);
or U3574 (N_3574,N_3252,N_3484);
nand U3575 (N_3575,N_3360,N_3394);
and U3576 (N_3576,N_3258,N_3478);
and U3577 (N_3577,N_3255,N_3352);
nand U3578 (N_3578,N_3407,N_3292);
and U3579 (N_3579,N_3452,N_3479);
nand U3580 (N_3580,N_3316,N_3426);
nand U3581 (N_3581,N_3434,N_3395);
xor U3582 (N_3582,N_3297,N_3498);
and U3583 (N_3583,N_3300,N_3353);
or U3584 (N_3584,N_3470,N_3444);
or U3585 (N_3585,N_3377,N_3427);
and U3586 (N_3586,N_3291,N_3308);
nor U3587 (N_3587,N_3299,N_3450);
and U3588 (N_3588,N_3439,N_3472);
xnor U3589 (N_3589,N_3270,N_3493);
nand U3590 (N_3590,N_3287,N_3274);
and U3591 (N_3591,N_3306,N_3347);
and U3592 (N_3592,N_3390,N_3269);
xor U3593 (N_3593,N_3311,N_3364);
nand U3594 (N_3594,N_3318,N_3429);
nor U3595 (N_3595,N_3322,N_3276);
nand U3596 (N_3596,N_3378,N_3280);
nor U3597 (N_3597,N_3359,N_3314);
xor U3598 (N_3598,N_3425,N_3415);
or U3599 (N_3599,N_3487,N_3374);
nand U3600 (N_3600,N_3351,N_3419);
and U3601 (N_3601,N_3325,N_3422);
nor U3602 (N_3602,N_3260,N_3288);
xnor U3603 (N_3603,N_3403,N_3259);
or U3604 (N_3604,N_3397,N_3375);
nor U3605 (N_3605,N_3251,N_3481);
or U3606 (N_3606,N_3387,N_3456);
and U3607 (N_3607,N_3432,N_3379);
xnor U3608 (N_3608,N_3296,N_3473);
xor U3609 (N_3609,N_3315,N_3399);
xor U3610 (N_3610,N_3393,N_3384);
xnor U3611 (N_3611,N_3406,N_3295);
nand U3612 (N_3612,N_3273,N_3402);
or U3613 (N_3613,N_3309,N_3421);
nand U3614 (N_3614,N_3317,N_3464);
and U3615 (N_3615,N_3362,N_3381);
and U3616 (N_3616,N_3335,N_3268);
xor U3617 (N_3617,N_3334,N_3272);
xor U3618 (N_3618,N_3256,N_3376);
nor U3619 (N_3619,N_3343,N_3371);
xnor U3620 (N_3620,N_3365,N_3263);
xor U3621 (N_3621,N_3290,N_3480);
xor U3622 (N_3622,N_3431,N_3303);
nor U3623 (N_3623,N_3366,N_3301);
or U3624 (N_3624,N_3496,N_3440);
nand U3625 (N_3625,N_3296,N_3493);
and U3626 (N_3626,N_3391,N_3461);
or U3627 (N_3627,N_3322,N_3316);
nand U3628 (N_3628,N_3344,N_3476);
xnor U3629 (N_3629,N_3326,N_3306);
xnor U3630 (N_3630,N_3347,N_3314);
xnor U3631 (N_3631,N_3448,N_3337);
or U3632 (N_3632,N_3291,N_3462);
and U3633 (N_3633,N_3420,N_3264);
or U3634 (N_3634,N_3475,N_3389);
and U3635 (N_3635,N_3323,N_3491);
xnor U3636 (N_3636,N_3378,N_3308);
nor U3637 (N_3637,N_3477,N_3273);
xor U3638 (N_3638,N_3408,N_3415);
nor U3639 (N_3639,N_3417,N_3499);
and U3640 (N_3640,N_3267,N_3264);
nor U3641 (N_3641,N_3489,N_3439);
nand U3642 (N_3642,N_3350,N_3250);
xor U3643 (N_3643,N_3305,N_3466);
or U3644 (N_3644,N_3427,N_3433);
nor U3645 (N_3645,N_3499,N_3473);
nand U3646 (N_3646,N_3461,N_3469);
xor U3647 (N_3647,N_3346,N_3375);
and U3648 (N_3648,N_3425,N_3289);
and U3649 (N_3649,N_3440,N_3354);
and U3650 (N_3650,N_3292,N_3327);
xor U3651 (N_3651,N_3283,N_3270);
and U3652 (N_3652,N_3359,N_3434);
xnor U3653 (N_3653,N_3337,N_3349);
xor U3654 (N_3654,N_3424,N_3430);
nand U3655 (N_3655,N_3478,N_3331);
nor U3656 (N_3656,N_3372,N_3457);
or U3657 (N_3657,N_3305,N_3279);
xor U3658 (N_3658,N_3418,N_3396);
xnor U3659 (N_3659,N_3454,N_3276);
or U3660 (N_3660,N_3290,N_3298);
nand U3661 (N_3661,N_3392,N_3395);
nor U3662 (N_3662,N_3378,N_3261);
nor U3663 (N_3663,N_3390,N_3289);
nor U3664 (N_3664,N_3262,N_3326);
xor U3665 (N_3665,N_3363,N_3255);
and U3666 (N_3666,N_3437,N_3257);
or U3667 (N_3667,N_3414,N_3328);
nand U3668 (N_3668,N_3420,N_3251);
nor U3669 (N_3669,N_3268,N_3359);
xor U3670 (N_3670,N_3467,N_3292);
or U3671 (N_3671,N_3252,N_3478);
nor U3672 (N_3672,N_3426,N_3301);
and U3673 (N_3673,N_3303,N_3469);
nor U3674 (N_3674,N_3440,N_3364);
nor U3675 (N_3675,N_3259,N_3353);
nor U3676 (N_3676,N_3330,N_3283);
xor U3677 (N_3677,N_3294,N_3408);
or U3678 (N_3678,N_3442,N_3392);
nor U3679 (N_3679,N_3275,N_3341);
or U3680 (N_3680,N_3486,N_3400);
nand U3681 (N_3681,N_3486,N_3357);
xnor U3682 (N_3682,N_3425,N_3310);
and U3683 (N_3683,N_3410,N_3257);
nor U3684 (N_3684,N_3437,N_3495);
nand U3685 (N_3685,N_3287,N_3443);
xnor U3686 (N_3686,N_3449,N_3403);
and U3687 (N_3687,N_3404,N_3311);
nand U3688 (N_3688,N_3275,N_3478);
nor U3689 (N_3689,N_3470,N_3464);
nor U3690 (N_3690,N_3484,N_3308);
and U3691 (N_3691,N_3411,N_3468);
and U3692 (N_3692,N_3443,N_3305);
nand U3693 (N_3693,N_3498,N_3440);
nor U3694 (N_3694,N_3307,N_3341);
or U3695 (N_3695,N_3370,N_3474);
or U3696 (N_3696,N_3421,N_3401);
xnor U3697 (N_3697,N_3355,N_3323);
or U3698 (N_3698,N_3383,N_3270);
or U3699 (N_3699,N_3481,N_3420);
xnor U3700 (N_3700,N_3483,N_3273);
xnor U3701 (N_3701,N_3354,N_3297);
and U3702 (N_3702,N_3382,N_3444);
xor U3703 (N_3703,N_3430,N_3252);
and U3704 (N_3704,N_3396,N_3374);
and U3705 (N_3705,N_3478,N_3398);
and U3706 (N_3706,N_3475,N_3385);
xor U3707 (N_3707,N_3381,N_3342);
and U3708 (N_3708,N_3345,N_3404);
and U3709 (N_3709,N_3484,N_3316);
and U3710 (N_3710,N_3452,N_3475);
and U3711 (N_3711,N_3348,N_3438);
nand U3712 (N_3712,N_3399,N_3466);
xnor U3713 (N_3713,N_3326,N_3445);
nor U3714 (N_3714,N_3333,N_3285);
xnor U3715 (N_3715,N_3497,N_3317);
and U3716 (N_3716,N_3300,N_3325);
or U3717 (N_3717,N_3452,N_3293);
nor U3718 (N_3718,N_3420,N_3407);
xor U3719 (N_3719,N_3489,N_3277);
nor U3720 (N_3720,N_3407,N_3439);
nor U3721 (N_3721,N_3346,N_3454);
nor U3722 (N_3722,N_3399,N_3377);
and U3723 (N_3723,N_3394,N_3264);
nand U3724 (N_3724,N_3298,N_3330);
nand U3725 (N_3725,N_3435,N_3251);
nor U3726 (N_3726,N_3391,N_3330);
nor U3727 (N_3727,N_3484,N_3354);
nand U3728 (N_3728,N_3436,N_3412);
xor U3729 (N_3729,N_3420,N_3477);
nand U3730 (N_3730,N_3450,N_3440);
nand U3731 (N_3731,N_3480,N_3493);
nand U3732 (N_3732,N_3291,N_3489);
xor U3733 (N_3733,N_3412,N_3482);
nand U3734 (N_3734,N_3436,N_3297);
nand U3735 (N_3735,N_3484,N_3348);
and U3736 (N_3736,N_3498,N_3355);
and U3737 (N_3737,N_3369,N_3251);
xnor U3738 (N_3738,N_3459,N_3473);
nor U3739 (N_3739,N_3445,N_3349);
nor U3740 (N_3740,N_3436,N_3388);
and U3741 (N_3741,N_3474,N_3473);
and U3742 (N_3742,N_3332,N_3282);
nand U3743 (N_3743,N_3375,N_3294);
xnor U3744 (N_3744,N_3389,N_3369);
nand U3745 (N_3745,N_3367,N_3307);
or U3746 (N_3746,N_3375,N_3264);
xnor U3747 (N_3747,N_3436,N_3420);
nand U3748 (N_3748,N_3413,N_3466);
and U3749 (N_3749,N_3344,N_3272);
and U3750 (N_3750,N_3507,N_3718);
or U3751 (N_3751,N_3573,N_3599);
nor U3752 (N_3752,N_3730,N_3505);
or U3753 (N_3753,N_3729,N_3580);
and U3754 (N_3754,N_3619,N_3659);
nor U3755 (N_3755,N_3696,N_3508);
or U3756 (N_3756,N_3546,N_3702);
and U3757 (N_3757,N_3519,N_3663);
or U3758 (N_3758,N_3656,N_3723);
or U3759 (N_3759,N_3612,N_3748);
or U3760 (N_3760,N_3694,N_3568);
and U3761 (N_3761,N_3699,N_3737);
or U3762 (N_3762,N_3606,N_3570);
or U3763 (N_3763,N_3711,N_3649);
nor U3764 (N_3764,N_3608,N_3685);
nor U3765 (N_3765,N_3740,N_3677);
and U3766 (N_3766,N_3624,N_3597);
xnor U3767 (N_3767,N_3544,N_3572);
or U3768 (N_3768,N_3506,N_3549);
or U3769 (N_3769,N_3538,N_3610);
nor U3770 (N_3770,N_3578,N_3561);
nor U3771 (N_3771,N_3531,N_3741);
nor U3772 (N_3772,N_3710,N_3552);
nor U3773 (N_3773,N_3747,N_3593);
nand U3774 (N_3774,N_3524,N_3667);
nand U3775 (N_3775,N_3714,N_3703);
nor U3776 (N_3776,N_3717,N_3690);
nand U3777 (N_3777,N_3749,N_3734);
nand U3778 (N_3778,N_3707,N_3736);
nor U3779 (N_3779,N_3692,N_3536);
nand U3780 (N_3780,N_3529,N_3648);
or U3781 (N_3781,N_3512,N_3509);
nand U3782 (N_3782,N_3587,N_3735);
or U3783 (N_3783,N_3521,N_3581);
nor U3784 (N_3784,N_3591,N_3637);
nand U3785 (N_3785,N_3642,N_3674);
nor U3786 (N_3786,N_3513,N_3629);
xor U3787 (N_3787,N_3645,N_3609);
xor U3788 (N_3788,N_3716,N_3522);
and U3789 (N_3789,N_3644,N_3541);
nor U3790 (N_3790,N_3560,N_3733);
nand U3791 (N_3791,N_3725,N_3650);
or U3792 (N_3792,N_3745,N_3671);
nor U3793 (N_3793,N_3662,N_3666);
and U3794 (N_3794,N_3559,N_3547);
or U3795 (N_3795,N_3681,N_3537);
nor U3796 (N_3796,N_3626,N_3643);
or U3797 (N_3797,N_3602,N_3502);
and U3798 (N_3798,N_3646,N_3651);
xnor U3799 (N_3799,N_3500,N_3661);
nand U3800 (N_3800,N_3652,N_3676);
or U3801 (N_3801,N_3586,N_3721);
nand U3802 (N_3802,N_3670,N_3664);
nor U3803 (N_3803,N_3744,N_3742);
or U3804 (N_3804,N_3689,N_3665);
and U3805 (N_3805,N_3563,N_3514);
or U3806 (N_3806,N_3583,N_3600);
nand U3807 (N_3807,N_3558,N_3682);
nor U3808 (N_3808,N_3553,N_3620);
xor U3809 (N_3809,N_3526,N_3616);
or U3810 (N_3810,N_3595,N_3728);
and U3811 (N_3811,N_3641,N_3715);
xor U3812 (N_3812,N_3594,N_3684);
nand U3813 (N_3813,N_3518,N_3686);
and U3814 (N_3814,N_3525,N_3556);
or U3815 (N_3815,N_3625,N_3614);
or U3816 (N_3816,N_3555,N_3501);
nor U3817 (N_3817,N_3530,N_3683);
xor U3818 (N_3818,N_3564,N_3658);
or U3819 (N_3819,N_3545,N_3635);
or U3820 (N_3820,N_3638,N_3675);
nand U3821 (N_3821,N_3706,N_3569);
nand U3822 (N_3822,N_3585,N_3708);
xor U3823 (N_3823,N_3596,N_3669);
or U3824 (N_3824,N_3695,N_3539);
and U3825 (N_3825,N_3551,N_3627);
nor U3826 (N_3826,N_3727,N_3673);
nand U3827 (N_3827,N_3705,N_3542);
nand U3828 (N_3828,N_3640,N_3712);
xnor U3829 (N_3829,N_3709,N_3653);
and U3830 (N_3830,N_3618,N_3575);
or U3831 (N_3831,N_3528,N_3679);
nand U3832 (N_3832,N_3603,N_3584);
nor U3833 (N_3833,N_3668,N_3598);
nand U3834 (N_3834,N_3565,N_3510);
nor U3835 (N_3835,N_3590,N_3571);
xor U3836 (N_3836,N_3520,N_3592);
xor U3837 (N_3837,N_3632,N_3550);
nand U3838 (N_3838,N_3535,N_3722);
and U3839 (N_3839,N_3726,N_3678);
nand U3840 (N_3840,N_3713,N_3634);
or U3841 (N_3841,N_3515,N_3720);
and U3842 (N_3842,N_3697,N_3704);
or U3843 (N_3843,N_3630,N_3688);
nor U3844 (N_3844,N_3691,N_3554);
or U3845 (N_3845,N_3517,N_3576);
and U3846 (N_3846,N_3693,N_3623);
xor U3847 (N_3847,N_3613,N_3504);
and U3848 (N_3848,N_3579,N_3503);
or U3849 (N_3849,N_3562,N_3601);
or U3850 (N_3850,N_3617,N_3533);
nor U3851 (N_3851,N_3655,N_3680);
xor U3852 (N_3852,N_3574,N_3534);
and U3853 (N_3853,N_3615,N_3732);
or U3854 (N_3854,N_3639,N_3687);
nand U3855 (N_3855,N_3698,N_3700);
nor U3856 (N_3856,N_3622,N_3636);
nor U3857 (N_3857,N_3532,N_3719);
nand U3858 (N_3858,N_3605,N_3582);
xnor U3859 (N_3859,N_3746,N_3523);
or U3860 (N_3860,N_3548,N_3511);
xnor U3861 (N_3861,N_3588,N_3731);
nand U3862 (N_3862,N_3633,N_3540);
nand U3863 (N_3863,N_3628,N_3743);
xor U3864 (N_3864,N_3654,N_3566);
and U3865 (N_3865,N_3631,N_3611);
nand U3866 (N_3866,N_3607,N_3604);
and U3867 (N_3867,N_3738,N_3672);
nor U3868 (N_3868,N_3557,N_3567);
or U3869 (N_3869,N_3516,N_3577);
and U3870 (N_3870,N_3724,N_3527);
and U3871 (N_3871,N_3621,N_3739);
and U3872 (N_3872,N_3543,N_3701);
xnor U3873 (N_3873,N_3657,N_3589);
nor U3874 (N_3874,N_3660,N_3647);
nor U3875 (N_3875,N_3691,N_3599);
nor U3876 (N_3876,N_3698,N_3745);
and U3877 (N_3877,N_3557,N_3698);
nand U3878 (N_3878,N_3504,N_3581);
or U3879 (N_3879,N_3674,N_3530);
nor U3880 (N_3880,N_3602,N_3716);
and U3881 (N_3881,N_3501,N_3549);
xor U3882 (N_3882,N_3672,N_3638);
or U3883 (N_3883,N_3552,N_3608);
or U3884 (N_3884,N_3647,N_3713);
and U3885 (N_3885,N_3577,N_3520);
or U3886 (N_3886,N_3743,N_3709);
xor U3887 (N_3887,N_3712,N_3748);
or U3888 (N_3888,N_3682,N_3602);
nor U3889 (N_3889,N_3697,N_3666);
nor U3890 (N_3890,N_3510,N_3555);
nand U3891 (N_3891,N_3618,N_3679);
nand U3892 (N_3892,N_3728,N_3631);
xor U3893 (N_3893,N_3682,N_3617);
or U3894 (N_3894,N_3721,N_3576);
and U3895 (N_3895,N_3592,N_3567);
nand U3896 (N_3896,N_3674,N_3723);
or U3897 (N_3897,N_3678,N_3595);
nand U3898 (N_3898,N_3658,N_3593);
or U3899 (N_3899,N_3742,N_3698);
and U3900 (N_3900,N_3518,N_3573);
xor U3901 (N_3901,N_3650,N_3573);
nor U3902 (N_3902,N_3649,N_3733);
nand U3903 (N_3903,N_3713,N_3590);
xor U3904 (N_3904,N_3628,N_3610);
nand U3905 (N_3905,N_3616,N_3629);
nor U3906 (N_3906,N_3543,N_3740);
xor U3907 (N_3907,N_3566,N_3611);
xor U3908 (N_3908,N_3510,N_3574);
nor U3909 (N_3909,N_3686,N_3737);
nand U3910 (N_3910,N_3689,N_3505);
nand U3911 (N_3911,N_3652,N_3615);
and U3912 (N_3912,N_3504,N_3571);
xor U3913 (N_3913,N_3565,N_3563);
or U3914 (N_3914,N_3603,N_3625);
nand U3915 (N_3915,N_3522,N_3590);
nor U3916 (N_3916,N_3715,N_3622);
nand U3917 (N_3917,N_3681,N_3685);
nand U3918 (N_3918,N_3626,N_3698);
and U3919 (N_3919,N_3627,N_3706);
nand U3920 (N_3920,N_3729,N_3630);
or U3921 (N_3921,N_3572,N_3653);
nand U3922 (N_3922,N_3683,N_3650);
nand U3923 (N_3923,N_3563,N_3549);
xnor U3924 (N_3924,N_3606,N_3639);
xor U3925 (N_3925,N_3670,N_3582);
nor U3926 (N_3926,N_3717,N_3692);
nor U3927 (N_3927,N_3633,N_3571);
and U3928 (N_3928,N_3538,N_3676);
and U3929 (N_3929,N_3667,N_3689);
or U3930 (N_3930,N_3612,N_3665);
and U3931 (N_3931,N_3674,N_3697);
xor U3932 (N_3932,N_3734,N_3624);
nor U3933 (N_3933,N_3555,N_3600);
and U3934 (N_3934,N_3710,N_3519);
and U3935 (N_3935,N_3637,N_3612);
xor U3936 (N_3936,N_3741,N_3696);
nor U3937 (N_3937,N_3635,N_3630);
and U3938 (N_3938,N_3720,N_3678);
nand U3939 (N_3939,N_3516,N_3639);
or U3940 (N_3940,N_3516,N_3749);
or U3941 (N_3941,N_3744,N_3525);
or U3942 (N_3942,N_3711,N_3508);
nand U3943 (N_3943,N_3569,N_3716);
nor U3944 (N_3944,N_3631,N_3599);
and U3945 (N_3945,N_3575,N_3639);
nand U3946 (N_3946,N_3627,N_3581);
nand U3947 (N_3947,N_3691,N_3600);
xnor U3948 (N_3948,N_3625,N_3626);
nand U3949 (N_3949,N_3521,N_3568);
nand U3950 (N_3950,N_3678,N_3684);
or U3951 (N_3951,N_3653,N_3622);
nand U3952 (N_3952,N_3736,N_3574);
or U3953 (N_3953,N_3502,N_3689);
xor U3954 (N_3954,N_3503,N_3624);
nand U3955 (N_3955,N_3722,N_3747);
and U3956 (N_3956,N_3629,N_3666);
xnor U3957 (N_3957,N_3579,N_3664);
and U3958 (N_3958,N_3692,N_3743);
or U3959 (N_3959,N_3677,N_3705);
nor U3960 (N_3960,N_3609,N_3558);
nor U3961 (N_3961,N_3720,N_3558);
xor U3962 (N_3962,N_3643,N_3746);
nor U3963 (N_3963,N_3673,N_3500);
or U3964 (N_3964,N_3719,N_3604);
or U3965 (N_3965,N_3526,N_3567);
and U3966 (N_3966,N_3515,N_3696);
and U3967 (N_3967,N_3573,N_3665);
nor U3968 (N_3968,N_3691,N_3695);
nor U3969 (N_3969,N_3744,N_3584);
and U3970 (N_3970,N_3535,N_3715);
and U3971 (N_3971,N_3665,N_3513);
xnor U3972 (N_3972,N_3572,N_3666);
and U3973 (N_3973,N_3703,N_3693);
nor U3974 (N_3974,N_3667,N_3700);
nor U3975 (N_3975,N_3697,N_3550);
or U3976 (N_3976,N_3501,N_3539);
and U3977 (N_3977,N_3572,N_3602);
and U3978 (N_3978,N_3565,N_3713);
and U3979 (N_3979,N_3519,N_3581);
nor U3980 (N_3980,N_3726,N_3533);
and U3981 (N_3981,N_3547,N_3693);
and U3982 (N_3982,N_3596,N_3652);
nor U3983 (N_3983,N_3652,N_3707);
or U3984 (N_3984,N_3561,N_3634);
nor U3985 (N_3985,N_3686,N_3635);
xor U3986 (N_3986,N_3540,N_3641);
or U3987 (N_3987,N_3661,N_3719);
and U3988 (N_3988,N_3641,N_3574);
xor U3989 (N_3989,N_3737,N_3537);
nor U3990 (N_3990,N_3664,N_3540);
and U3991 (N_3991,N_3595,N_3726);
nor U3992 (N_3992,N_3539,N_3598);
nand U3993 (N_3993,N_3529,N_3689);
nor U3994 (N_3994,N_3666,N_3624);
xor U3995 (N_3995,N_3665,N_3553);
and U3996 (N_3996,N_3586,N_3626);
nand U3997 (N_3997,N_3664,N_3528);
nor U3998 (N_3998,N_3523,N_3666);
or U3999 (N_3999,N_3530,N_3724);
nand U4000 (N_4000,N_3832,N_3963);
nand U4001 (N_4001,N_3831,N_3817);
nand U4002 (N_4002,N_3935,N_3942);
nand U4003 (N_4003,N_3898,N_3985);
or U4004 (N_4004,N_3926,N_3774);
and U4005 (N_4005,N_3909,N_3953);
xor U4006 (N_4006,N_3859,N_3777);
nor U4007 (N_4007,N_3921,N_3752);
nand U4008 (N_4008,N_3839,N_3772);
and U4009 (N_4009,N_3893,N_3904);
xor U4010 (N_4010,N_3986,N_3871);
and U4011 (N_4011,N_3965,N_3932);
or U4012 (N_4012,N_3785,N_3759);
xnor U4013 (N_4013,N_3861,N_3998);
or U4014 (N_4014,N_3996,N_3790);
or U4015 (N_4015,N_3860,N_3762);
and U4016 (N_4016,N_3851,N_3823);
nor U4017 (N_4017,N_3853,N_3951);
or U4018 (N_4018,N_3810,N_3895);
nor U4019 (N_4019,N_3833,N_3882);
xnor U4020 (N_4020,N_3936,N_3783);
nand U4021 (N_4021,N_3946,N_3910);
xor U4022 (N_4022,N_3891,N_3931);
nor U4023 (N_4023,N_3906,N_3956);
nand U4024 (N_4024,N_3753,N_3940);
nor U4025 (N_4025,N_3896,N_3820);
xnor U4026 (N_4026,N_3880,N_3813);
xor U4027 (N_4027,N_3829,N_3773);
nor U4028 (N_4028,N_3868,N_3838);
and U4029 (N_4029,N_3781,N_3954);
or U4030 (N_4030,N_3750,N_3879);
or U4031 (N_4031,N_3760,N_3802);
nor U4032 (N_4032,N_3999,N_3768);
nor U4033 (N_4033,N_3903,N_3830);
nand U4034 (N_4034,N_3763,N_3855);
nand U4035 (N_4035,N_3850,N_3870);
or U4036 (N_4036,N_3801,N_3907);
xor U4037 (N_4037,N_3991,N_3885);
nor U4038 (N_4038,N_3865,N_3990);
nand U4039 (N_4039,N_3842,N_3966);
nand U4040 (N_4040,N_3983,N_3866);
nand U4041 (N_4041,N_3789,N_3794);
or U4042 (N_4042,N_3979,N_3884);
xor U4043 (N_4043,N_3755,N_3930);
nor U4044 (N_4044,N_3835,N_3765);
and U4045 (N_4045,N_3796,N_3788);
nor U4046 (N_4046,N_3771,N_3800);
nor U4047 (N_4047,N_3857,N_3797);
nand U4048 (N_4048,N_3766,N_3841);
xor U4049 (N_4049,N_3843,N_3978);
nand U4050 (N_4050,N_3920,N_3957);
or U4051 (N_4051,N_3937,N_3875);
and U4052 (N_4052,N_3892,N_3872);
xor U4053 (N_4053,N_3908,N_3812);
nand U4054 (N_4054,N_3867,N_3949);
nor U4055 (N_4055,N_3929,N_3976);
xor U4056 (N_4056,N_3913,N_3846);
xnor U4057 (N_4057,N_3798,N_3803);
xnor U4058 (N_4058,N_3925,N_3761);
xor U4059 (N_4059,N_3947,N_3992);
nand U4060 (N_4060,N_3905,N_3887);
and U4061 (N_4061,N_3852,N_3828);
and U4062 (N_4062,N_3901,N_3764);
or U4063 (N_4063,N_3894,N_3784);
nand U4064 (N_4064,N_3899,N_3944);
nor U4065 (N_4065,N_3915,N_3881);
xnor U4066 (N_4066,N_3970,N_3993);
xnor U4067 (N_4067,N_3858,N_3793);
and U4068 (N_4068,N_3757,N_3834);
or U4069 (N_4069,N_3811,N_3856);
nand U4070 (N_4070,N_3987,N_3786);
and U4071 (N_4071,N_3969,N_3988);
xnor U4072 (N_4072,N_3938,N_3818);
xor U4073 (N_4073,N_3943,N_3981);
nor U4074 (N_4074,N_3883,N_3805);
and U4075 (N_4075,N_3758,N_3847);
nor U4076 (N_4076,N_3945,N_3815);
nor U4077 (N_4077,N_3864,N_3961);
and U4078 (N_4078,N_3917,N_3977);
or U4079 (N_4079,N_3776,N_3997);
nor U4080 (N_4080,N_3756,N_3919);
or U4081 (N_4081,N_3751,N_3918);
and U4082 (N_4082,N_3827,N_3821);
and U4083 (N_4083,N_3886,N_3982);
and U4084 (N_4084,N_3955,N_3914);
nor U4085 (N_4085,N_3825,N_3989);
nor U4086 (N_4086,N_3927,N_3950);
xnor U4087 (N_4087,N_3837,N_3822);
and U4088 (N_4088,N_3964,N_3862);
and U4089 (N_4089,N_3767,N_3971);
or U4090 (N_4090,N_3775,N_3962);
or U4091 (N_4091,N_3779,N_3916);
nor U4092 (N_4092,N_3924,N_3819);
xor U4093 (N_4093,N_3911,N_3769);
nand U4094 (N_4094,N_3876,N_3877);
xor U4095 (N_4095,N_3770,N_3958);
xnor U4096 (N_4096,N_3897,N_3980);
or U4097 (N_4097,N_3791,N_3902);
nor U4098 (N_4098,N_3972,N_3848);
xor U4099 (N_4099,N_3854,N_3952);
xnor U4100 (N_4100,N_3782,N_3948);
or U4101 (N_4101,N_3869,N_3863);
nand U4102 (N_4102,N_3836,N_3994);
and U4103 (N_4103,N_3795,N_3995);
xor U4104 (N_4104,N_3941,N_3975);
nand U4105 (N_4105,N_3984,N_3890);
or U4106 (N_4106,N_3808,N_3780);
nand U4107 (N_4107,N_3778,N_3939);
or U4108 (N_4108,N_3960,N_3968);
nor U4109 (N_4109,N_3792,N_3824);
nand U4110 (N_4110,N_3809,N_3959);
nand U4111 (N_4111,N_3923,N_3799);
nand U4112 (N_4112,N_3826,N_3873);
xor U4113 (N_4113,N_3845,N_3933);
and U4114 (N_4114,N_3900,N_3844);
xor U4115 (N_4115,N_3922,N_3814);
xnor U4116 (N_4116,N_3974,N_3912);
xor U4117 (N_4117,N_3973,N_3849);
or U4118 (N_4118,N_3878,N_3934);
nor U4119 (N_4119,N_3816,N_3874);
nor U4120 (N_4120,N_3840,N_3967);
or U4121 (N_4121,N_3787,N_3928);
nor U4122 (N_4122,N_3889,N_3888);
or U4123 (N_4123,N_3806,N_3807);
nand U4124 (N_4124,N_3804,N_3754);
or U4125 (N_4125,N_3866,N_3971);
or U4126 (N_4126,N_3915,N_3961);
xor U4127 (N_4127,N_3803,N_3946);
xnor U4128 (N_4128,N_3990,N_3905);
xor U4129 (N_4129,N_3901,N_3773);
nand U4130 (N_4130,N_3929,N_3881);
and U4131 (N_4131,N_3774,N_3999);
or U4132 (N_4132,N_3972,N_3887);
and U4133 (N_4133,N_3970,N_3874);
nor U4134 (N_4134,N_3897,N_3878);
xnor U4135 (N_4135,N_3961,N_3984);
nand U4136 (N_4136,N_3834,N_3815);
xnor U4137 (N_4137,N_3980,N_3885);
xnor U4138 (N_4138,N_3765,N_3854);
or U4139 (N_4139,N_3955,N_3926);
and U4140 (N_4140,N_3944,N_3963);
or U4141 (N_4141,N_3956,N_3988);
xor U4142 (N_4142,N_3816,N_3860);
or U4143 (N_4143,N_3813,N_3961);
or U4144 (N_4144,N_3851,N_3886);
nand U4145 (N_4145,N_3806,N_3763);
nor U4146 (N_4146,N_3809,N_3885);
and U4147 (N_4147,N_3839,N_3758);
nand U4148 (N_4148,N_3818,N_3847);
xor U4149 (N_4149,N_3905,N_3798);
and U4150 (N_4150,N_3890,N_3785);
or U4151 (N_4151,N_3826,N_3783);
xor U4152 (N_4152,N_3849,N_3893);
xor U4153 (N_4153,N_3875,N_3978);
nand U4154 (N_4154,N_3910,N_3978);
and U4155 (N_4155,N_3993,N_3785);
nor U4156 (N_4156,N_3757,N_3792);
and U4157 (N_4157,N_3894,N_3838);
nor U4158 (N_4158,N_3751,N_3862);
nor U4159 (N_4159,N_3889,N_3795);
nand U4160 (N_4160,N_3857,N_3848);
nand U4161 (N_4161,N_3843,N_3891);
nor U4162 (N_4162,N_3793,N_3970);
xnor U4163 (N_4163,N_3753,N_3869);
and U4164 (N_4164,N_3868,N_3959);
or U4165 (N_4165,N_3880,N_3782);
xor U4166 (N_4166,N_3850,N_3778);
nor U4167 (N_4167,N_3766,N_3898);
nor U4168 (N_4168,N_3817,N_3850);
nand U4169 (N_4169,N_3973,N_3870);
and U4170 (N_4170,N_3865,N_3761);
xnor U4171 (N_4171,N_3766,N_3955);
nand U4172 (N_4172,N_3978,N_3998);
nand U4173 (N_4173,N_3857,N_3862);
nor U4174 (N_4174,N_3778,N_3971);
and U4175 (N_4175,N_3855,N_3888);
nor U4176 (N_4176,N_3954,N_3861);
nand U4177 (N_4177,N_3942,N_3959);
nand U4178 (N_4178,N_3788,N_3786);
nand U4179 (N_4179,N_3917,N_3842);
or U4180 (N_4180,N_3765,N_3784);
nor U4181 (N_4181,N_3875,N_3764);
or U4182 (N_4182,N_3874,N_3992);
or U4183 (N_4183,N_3834,N_3773);
and U4184 (N_4184,N_3762,N_3996);
and U4185 (N_4185,N_3967,N_3944);
nand U4186 (N_4186,N_3755,N_3884);
nor U4187 (N_4187,N_3919,N_3872);
and U4188 (N_4188,N_3801,N_3951);
and U4189 (N_4189,N_3830,N_3802);
nand U4190 (N_4190,N_3996,N_3775);
or U4191 (N_4191,N_3764,N_3921);
or U4192 (N_4192,N_3852,N_3965);
nor U4193 (N_4193,N_3921,N_3780);
or U4194 (N_4194,N_3838,N_3822);
or U4195 (N_4195,N_3764,N_3950);
xnor U4196 (N_4196,N_3882,N_3972);
xnor U4197 (N_4197,N_3905,N_3839);
nand U4198 (N_4198,N_3808,N_3829);
nand U4199 (N_4199,N_3920,N_3919);
and U4200 (N_4200,N_3856,N_3825);
nand U4201 (N_4201,N_3929,N_3954);
nand U4202 (N_4202,N_3827,N_3979);
and U4203 (N_4203,N_3893,N_3933);
and U4204 (N_4204,N_3889,N_3751);
nor U4205 (N_4205,N_3870,N_3797);
xnor U4206 (N_4206,N_3835,N_3874);
nor U4207 (N_4207,N_3948,N_3832);
nor U4208 (N_4208,N_3955,N_3814);
or U4209 (N_4209,N_3987,N_3912);
xnor U4210 (N_4210,N_3972,N_3945);
or U4211 (N_4211,N_3816,N_3948);
xor U4212 (N_4212,N_3941,N_3892);
xor U4213 (N_4213,N_3881,N_3811);
xor U4214 (N_4214,N_3982,N_3872);
nand U4215 (N_4215,N_3892,N_3861);
nand U4216 (N_4216,N_3912,N_3874);
xor U4217 (N_4217,N_3759,N_3864);
or U4218 (N_4218,N_3907,N_3774);
xnor U4219 (N_4219,N_3894,N_3878);
and U4220 (N_4220,N_3848,N_3953);
or U4221 (N_4221,N_3991,N_3884);
nor U4222 (N_4222,N_3823,N_3778);
xor U4223 (N_4223,N_3921,N_3870);
xor U4224 (N_4224,N_3994,N_3960);
or U4225 (N_4225,N_3813,N_3923);
nand U4226 (N_4226,N_3772,N_3824);
xnor U4227 (N_4227,N_3867,N_3813);
nor U4228 (N_4228,N_3914,N_3762);
xor U4229 (N_4229,N_3975,N_3807);
nor U4230 (N_4230,N_3854,N_3888);
or U4231 (N_4231,N_3911,N_3937);
and U4232 (N_4232,N_3913,N_3963);
or U4233 (N_4233,N_3809,N_3981);
and U4234 (N_4234,N_3788,N_3930);
nand U4235 (N_4235,N_3857,N_3935);
and U4236 (N_4236,N_3940,N_3806);
nand U4237 (N_4237,N_3903,N_3788);
nor U4238 (N_4238,N_3916,N_3984);
nand U4239 (N_4239,N_3987,N_3874);
and U4240 (N_4240,N_3969,N_3975);
or U4241 (N_4241,N_3880,N_3831);
xor U4242 (N_4242,N_3825,N_3870);
nor U4243 (N_4243,N_3885,N_3936);
nor U4244 (N_4244,N_3950,N_3977);
xor U4245 (N_4245,N_3927,N_3820);
or U4246 (N_4246,N_3877,N_3789);
nand U4247 (N_4247,N_3967,N_3804);
nand U4248 (N_4248,N_3861,N_3888);
and U4249 (N_4249,N_3916,N_3981);
and U4250 (N_4250,N_4238,N_4231);
or U4251 (N_4251,N_4138,N_4217);
nor U4252 (N_4252,N_4222,N_4183);
nor U4253 (N_4253,N_4076,N_4195);
xor U4254 (N_4254,N_4153,N_4111);
and U4255 (N_4255,N_4119,N_4063);
xnor U4256 (N_4256,N_4194,N_4201);
or U4257 (N_4257,N_4016,N_4139);
nor U4258 (N_4258,N_4107,N_4006);
or U4259 (N_4259,N_4077,N_4230);
nor U4260 (N_4260,N_4215,N_4037);
or U4261 (N_4261,N_4154,N_4017);
nor U4262 (N_4262,N_4212,N_4056);
and U4263 (N_4263,N_4001,N_4242);
nand U4264 (N_4264,N_4202,N_4009);
nand U4265 (N_4265,N_4027,N_4171);
nand U4266 (N_4266,N_4169,N_4047);
nand U4267 (N_4267,N_4032,N_4034);
nor U4268 (N_4268,N_4012,N_4235);
nor U4269 (N_4269,N_4136,N_4046);
nor U4270 (N_4270,N_4246,N_4224);
and U4271 (N_4271,N_4181,N_4233);
or U4272 (N_4272,N_4148,N_4244);
or U4273 (N_4273,N_4102,N_4147);
nand U4274 (N_4274,N_4226,N_4184);
nor U4275 (N_4275,N_4140,N_4072);
nand U4276 (N_4276,N_4179,N_4010);
nor U4277 (N_4277,N_4156,N_4237);
xnor U4278 (N_4278,N_4090,N_4018);
nand U4279 (N_4279,N_4143,N_4108);
nor U4280 (N_4280,N_4099,N_4022);
or U4281 (N_4281,N_4228,N_4190);
nor U4282 (N_4282,N_4101,N_4095);
nand U4283 (N_4283,N_4019,N_4053);
nor U4284 (N_4284,N_4191,N_4064);
xnor U4285 (N_4285,N_4227,N_4024);
nor U4286 (N_4286,N_4152,N_4124);
or U4287 (N_4287,N_4085,N_4091);
nor U4288 (N_4288,N_4070,N_4097);
nor U4289 (N_4289,N_4120,N_4223);
nand U4290 (N_4290,N_4177,N_4060);
nor U4291 (N_4291,N_4208,N_4051);
nor U4292 (N_4292,N_4192,N_4113);
nand U4293 (N_4293,N_4081,N_4248);
nor U4294 (N_4294,N_4245,N_4214);
nor U4295 (N_4295,N_4232,N_4132);
and U4296 (N_4296,N_4182,N_4015);
nor U4297 (N_4297,N_4155,N_4149);
nor U4298 (N_4298,N_4236,N_4062);
nor U4299 (N_4299,N_4115,N_4249);
nand U4300 (N_4300,N_4158,N_4186);
nand U4301 (N_4301,N_4104,N_4096);
or U4302 (N_4302,N_4067,N_4164);
or U4303 (N_4303,N_4100,N_4000);
xor U4304 (N_4304,N_4023,N_4160);
nand U4305 (N_4305,N_4065,N_4042);
xnor U4306 (N_4306,N_4128,N_4165);
nor U4307 (N_4307,N_4008,N_4144);
and U4308 (N_4308,N_4007,N_4030);
nand U4309 (N_4309,N_4075,N_4172);
or U4310 (N_4310,N_4157,N_4112);
nand U4311 (N_4311,N_4173,N_4218);
nor U4312 (N_4312,N_4031,N_4205);
nand U4313 (N_4313,N_4094,N_4078);
xnor U4314 (N_4314,N_4028,N_4106);
or U4315 (N_4315,N_4175,N_4011);
or U4316 (N_4316,N_4048,N_4103);
xnor U4317 (N_4317,N_4021,N_4033);
nor U4318 (N_4318,N_4145,N_4066);
nand U4319 (N_4319,N_4013,N_4130);
nand U4320 (N_4320,N_4005,N_4026);
and U4321 (N_4321,N_4040,N_4003);
nor U4322 (N_4322,N_4239,N_4197);
or U4323 (N_4323,N_4200,N_4151);
or U4324 (N_4324,N_4061,N_4054);
or U4325 (N_4325,N_4117,N_4109);
nand U4326 (N_4326,N_4123,N_4125);
nand U4327 (N_4327,N_4073,N_4088);
xnor U4328 (N_4328,N_4216,N_4220);
xor U4329 (N_4329,N_4198,N_4247);
xor U4330 (N_4330,N_4089,N_4114);
xor U4331 (N_4331,N_4059,N_4161);
or U4332 (N_4332,N_4079,N_4142);
nor U4333 (N_4333,N_4122,N_4105);
and U4334 (N_4334,N_4213,N_4038);
nand U4335 (N_4335,N_4049,N_4131);
xor U4336 (N_4336,N_4187,N_4135);
nand U4337 (N_4337,N_4168,N_4189);
nand U4338 (N_4338,N_4080,N_4203);
nor U4339 (N_4339,N_4146,N_4240);
and U4340 (N_4340,N_4166,N_4170);
xor U4341 (N_4341,N_4002,N_4129);
or U4342 (N_4342,N_4086,N_4110);
and U4343 (N_4343,N_4041,N_4225);
and U4344 (N_4344,N_4219,N_4092);
nand U4345 (N_4345,N_4084,N_4127);
and U4346 (N_4346,N_4055,N_4121);
xor U4347 (N_4347,N_4193,N_4057);
and U4348 (N_4348,N_4118,N_4176);
nor U4349 (N_4349,N_4241,N_4206);
and U4350 (N_4350,N_4185,N_4159);
and U4351 (N_4351,N_4162,N_4133);
nor U4352 (N_4352,N_4141,N_4074);
xor U4353 (N_4353,N_4116,N_4134);
nor U4354 (N_4354,N_4068,N_4050);
nand U4355 (N_4355,N_4174,N_4196);
or U4356 (N_4356,N_4083,N_4188);
or U4357 (N_4357,N_4199,N_4210);
and U4358 (N_4358,N_4087,N_4014);
xnor U4359 (N_4359,N_4082,N_4180);
and U4360 (N_4360,N_4204,N_4126);
nor U4361 (N_4361,N_4052,N_4167);
and U4362 (N_4362,N_4178,N_4229);
or U4363 (N_4363,N_4058,N_4043);
nand U4364 (N_4364,N_4234,N_4207);
and U4365 (N_4365,N_4069,N_4004);
and U4366 (N_4366,N_4044,N_4211);
nor U4367 (N_4367,N_4209,N_4071);
and U4368 (N_4368,N_4025,N_4093);
nand U4369 (N_4369,N_4029,N_4035);
xor U4370 (N_4370,N_4243,N_4045);
or U4371 (N_4371,N_4098,N_4020);
nand U4372 (N_4372,N_4150,N_4221);
nand U4373 (N_4373,N_4039,N_4163);
xor U4374 (N_4374,N_4137,N_4036);
nand U4375 (N_4375,N_4011,N_4059);
and U4376 (N_4376,N_4122,N_4069);
and U4377 (N_4377,N_4147,N_4223);
nor U4378 (N_4378,N_4009,N_4150);
and U4379 (N_4379,N_4096,N_4216);
nor U4380 (N_4380,N_4158,N_4226);
and U4381 (N_4381,N_4003,N_4222);
nor U4382 (N_4382,N_4186,N_4156);
nand U4383 (N_4383,N_4135,N_4107);
and U4384 (N_4384,N_4092,N_4240);
xnor U4385 (N_4385,N_4142,N_4151);
nand U4386 (N_4386,N_4158,N_4123);
or U4387 (N_4387,N_4118,N_4066);
xor U4388 (N_4388,N_4118,N_4012);
nor U4389 (N_4389,N_4100,N_4048);
or U4390 (N_4390,N_4077,N_4023);
nor U4391 (N_4391,N_4108,N_4216);
and U4392 (N_4392,N_4120,N_4002);
or U4393 (N_4393,N_4007,N_4231);
nand U4394 (N_4394,N_4014,N_4074);
nand U4395 (N_4395,N_4054,N_4031);
nor U4396 (N_4396,N_4044,N_4229);
xor U4397 (N_4397,N_4093,N_4026);
nand U4398 (N_4398,N_4184,N_4008);
nor U4399 (N_4399,N_4109,N_4040);
and U4400 (N_4400,N_4211,N_4225);
or U4401 (N_4401,N_4048,N_4027);
nand U4402 (N_4402,N_4097,N_4139);
nand U4403 (N_4403,N_4199,N_4160);
nand U4404 (N_4404,N_4040,N_4216);
xor U4405 (N_4405,N_4197,N_4238);
xor U4406 (N_4406,N_4182,N_4185);
nor U4407 (N_4407,N_4206,N_4161);
xnor U4408 (N_4408,N_4208,N_4059);
xor U4409 (N_4409,N_4169,N_4126);
xor U4410 (N_4410,N_4081,N_4092);
nand U4411 (N_4411,N_4234,N_4186);
or U4412 (N_4412,N_4227,N_4070);
nor U4413 (N_4413,N_4248,N_4045);
and U4414 (N_4414,N_4239,N_4040);
and U4415 (N_4415,N_4209,N_4217);
or U4416 (N_4416,N_4175,N_4087);
xor U4417 (N_4417,N_4072,N_4135);
and U4418 (N_4418,N_4211,N_4010);
or U4419 (N_4419,N_4153,N_4154);
or U4420 (N_4420,N_4014,N_4161);
xnor U4421 (N_4421,N_4143,N_4131);
nand U4422 (N_4422,N_4012,N_4236);
and U4423 (N_4423,N_4153,N_4176);
nor U4424 (N_4424,N_4017,N_4040);
nand U4425 (N_4425,N_4005,N_4144);
nand U4426 (N_4426,N_4019,N_4209);
or U4427 (N_4427,N_4028,N_4069);
nor U4428 (N_4428,N_4144,N_4052);
or U4429 (N_4429,N_4169,N_4004);
xnor U4430 (N_4430,N_4035,N_4203);
and U4431 (N_4431,N_4189,N_4243);
nor U4432 (N_4432,N_4026,N_4172);
or U4433 (N_4433,N_4200,N_4160);
nor U4434 (N_4434,N_4051,N_4001);
xor U4435 (N_4435,N_4092,N_4100);
or U4436 (N_4436,N_4205,N_4013);
or U4437 (N_4437,N_4163,N_4120);
nand U4438 (N_4438,N_4071,N_4223);
or U4439 (N_4439,N_4121,N_4203);
xnor U4440 (N_4440,N_4004,N_4141);
nor U4441 (N_4441,N_4234,N_4083);
xnor U4442 (N_4442,N_4102,N_4025);
and U4443 (N_4443,N_4237,N_4146);
and U4444 (N_4444,N_4160,N_4015);
xor U4445 (N_4445,N_4098,N_4080);
nand U4446 (N_4446,N_4243,N_4052);
or U4447 (N_4447,N_4197,N_4080);
or U4448 (N_4448,N_4038,N_4049);
and U4449 (N_4449,N_4228,N_4211);
or U4450 (N_4450,N_4207,N_4157);
and U4451 (N_4451,N_4060,N_4061);
xor U4452 (N_4452,N_4130,N_4175);
xor U4453 (N_4453,N_4157,N_4083);
or U4454 (N_4454,N_4057,N_4086);
nand U4455 (N_4455,N_4102,N_4112);
nor U4456 (N_4456,N_4020,N_4177);
or U4457 (N_4457,N_4247,N_4059);
nor U4458 (N_4458,N_4201,N_4149);
and U4459 (N_4459,N_4198,N_4036);
nand U4460 (N_4460,N_4022,N_4000);
nor U4461 (N_4461,N_4001,N_4209);
xor U4462 (N_4462,N_4229,N_4043);
nand U4463 (N_4463,N_4180,N_4000);
xnor U4464 (N_4464,N_4014,N_4102);
nor U4465 (N_4465,N_4016,N_4081);
xnor U4466 (N_4466,N_4232,N_4002);
nor U4467 (N_4467,N_4050,N_4141);
xor U4468 (N_4468,N_4052,N_4215);
xnor U4469 (N_4469,N_4014,N_4129);
or U4470 (N_4470,N_4132,N_4011);
nor U4471 (N_4471,N_4020,N_4125);
or U4472 (N_4472,N_4110,N_4109);
xor U4473 (N_4473,N_4220,N_4065);
and U4474 (N_4474,N_4152,N_4018);
and U4475 (N_4475,N_4201,N_4235);
nand U4476 (N_4476,N_4173,N_4179);
xor U4477 (N_4477,N_4111,N_4163);
nand U4478 (N_4478,N_4005,N_4135);
nor U4479 (N_4479,N_4060,N_4053);
and U4480 (N_4480,N_4024,N_4080);
nor U4481 (N_4481,N_4023,N_4249);
nor U4482 (N_4482,N_4036,N_4061);
nand U4483 (N_4483,N_4231,N_4046);
and U4484 (N_4484,N_4020,N_4192);
nor U4485 (N_4485,N_4048,N_4203);
xor U4486 (N_4486,N_4057,N_4226);
nand U4487 (N_4487,N_4112,N_4082);
and U4488 (N_4488,N_4023,N_4113);
or U4489 (N_4489,N_4037,N_4132);
nand U4490 (N_4490,N_4182,N_4140);
and U4491 (N_4491,N_4200,N_4245);
nand U4492 (N_4492,N_4199,N_4140);
nor U4493 (N_4493,N_4175,N_4241);
or U4494 (N_4494,N_4049,N_4234);
xnor U4495 (N_4495,N_4242,N_4014);
and U4496 (N_4496,N_4026,N_4163);
xnor U4497 (N_4497,N_4142,N_4082);
nor U4498 (N_4498,N_4003,N_4215);
nor U4499 (N_4499,N_4049,N_4012);
or U4500 (N_4500,N_4277,N_4406);
nor U4501 (N_4501,N_4263,N_4491);
nand U4502 (N_4502,N_4333,N_4371);
nor U4503 (N_4503,N_4419,N_4397);
xor U4504 (N_4504,N_4395,N_4387);
xor U4505 (N_4505,N_4368,N_4311);
and U4506 (N_4506,N_4355,N_4288);
nor U4507 (N_4507,N_4303,N_4280);
nor U4508 (N_4508,N_4421,N_4461);
xor U4509 (N_4509,N_4274,N_4439);
nand U4510 (N_4510,N_4443,N_4324);
nor U4511 (N_4511,N_4310,N_4262);
or U4512 (N_4512,N_4389,N_4489);
xor U4513 (N_4513,N_4320,N_4348);
xnor U4514 (N_4514,N_4334,N_4392);
and U4515 (N_4515,N_4290,N_4377);
nand U4516 (N_4516,N_4374,N_4317);
xor U4517 (N_4517,N_4420,N_4367);
nand U4518 (N_4518,N_4474,N_4437);
nor U4519 (N_4519,N_4457,N_4251);
and U4520 (N_4520,N_4449,N_4287);
or U4521 (N_4521,N_4429,N_4422);
nand U4522 (N_4522,N_4412,N_4466);
nor U4523 (N_4523,N_4292,N_4362);
and U4524 (N_4524,N_4431,N_4276);
or U4525 (N_4525,N_4430,N_4341);
or U4526 (N_4526,N_4448,N_4451);
xnor U4527 (N_4527,N_4286,N_4345);
nand U4528 (N_4528,N_4401,N_4417);
xor U4529 (N_4529,N_4464,N_4269);
and U4530 (N_4530,N_4253,N_4436);
nand U4531 (N_4531,N_4470,N_4256);
and U4532 (N_4532,N_4283,N_4325);
xor U4533 (N_4533,N_4364,N_4273);
or U4534 (N_4534,N_4354,N_4336);
xnor U4535 (N_4535,N_4279,N_4453);
nor U4536 (N_4536,N_4346,N_4440);
xnor U4537 (N_4537,N_4328,N_4265);
and U4538 (N_4538,N_4376,N_4257);
nand U4539 (N_4539,N_4472,N_4267);
and U4540 (N_4540,N_4427,N_4450);
or U4541 (N_4541,N_4275,N_4352);
and U4542 (N_4542,N_4483,N_4384);
xor U4543 (N_4543,N_4382,N_4293);
xor U4544 (N_4544,N_4441,N_4399);
nand U4545 (N_4545,N_4282,N_4281);
nand U4546 (N_4546,N_4314,N_4432);
nor U4547 (N_4547,N_4459,N_4379);
nor U4548 (N_4548,N_4497,N_4396);
nand U4549 (N_4549,N_4363,N_4468);
nor U4550 (N_4550,N_4299,N_4258);
and U4551 (N_4551,N_4447,N_4261);
nand U4552 (N_4552,N_4458,N_4360);
nand U4553 (N_4553,N_4388,N_4375);
nor U4554 (N_4554,N_4343,N_4494);
and U4555 (N_4555,N_4418,N_4271);
xnor U4556 (N_4556,N_4296,N_4347);
or U4557 (N_4557,N_4358,N_4438);
or U4558 (N_4558,N_4254,N_4498);
and U4559 (N_4559,N_4408,N_4252);
nor U4560 (N_4560,N_4465,N_4488);
and U4561 (N_4561,N_4359,N_4322);
xor U4562 (N_4562,N_4302,N_4297);
or U4563 (N_4563,N_4295,N_4460);
nor U4564 (N_4564,N_4285,N_4260);
nand U4565 (N_4565,N_4493,N_4486);
and U4566 (N_4566,N_4351,N_4411);
and U4567 (N_4567,N_4473,N_4416);
and U4568 (N_4568,N_4309,N_4381);
nor U4569 (N_4569,N_4380,N_4316);
nand U4570 (N_4570,N_4259,N_4475);
or U4571 (N_4571,N_4323,N_4394);
nand U4572 (N_4572,N_4306,N_4462);
or U4573 (N_4573,N_4312,N_4445);
nor U4574 (N_4574,N_4484,N_4423);
or U4575 (N_4575,N_4289,N_4487);
xor U4576 (N_4576,N_4383,N_4369);
nor U4577 (N_4577,N_4313,N_4272);
and U4578 (N_4578,N_4353,N_4372);
or U4579 (N_4579,N_4326,N_4403);
nor U4580 (N_4580,N_4469,N_4335);
and U4581 (N_4581,N_4329,N_4467);
and U4582 (N_4582,N_4357,N_4496);
nor U4583 (N_4583,N_4318,N_4342);
nor U4584 (N_4584,N_4327,N_4410);
xor U4585 (N_4585,N_4305,N_4331);
nor U4586 (N_4586,N_4463,N_4482);
xnor U4587 (N_4587,N_4315,N_4444);
nor U4588 (N_4588,N_4308,N_4391);
and U4589 (N_4589,N_4485,N_4378);
and U4590 (N_4590,N_4332,N_4319);
nor U4591 (N_4591,N_4393,N_4471);
or U4592 (N_4592,N_4402,N_4492);
nor U4593 (N_4593,N_4338,N_4479);
or U4594 (N_4594,N_4278,N_4407);
and U4595 (N_4595,N_4250,N_4270);
nor U4596 (N_4596,N_4495,N_4452);
or U4597 (N_4597,N_4321,N_4294);
nand U4598 (N_4598,N_4490,N_4301);
and U4599 (N_4599,N_4435,N_4291);
xnor U4600 (N_4600,N_4414,N_4300);
xor U4601 (N_4601,N_4330,N_4337);
and U4602 (N_4602,N_4454,N_4424);
nor U4603 (N_4603,N_4481,N_4339);
and U4604 (N_4604,N_4428,N_4255);
nor U4605 (N_4605,N_4370,N_4304);
nand U4606 (N_4606,N_4477,N_4268);
nand U4607 (N_4607,N_4284,N_4404);
nand U4608 (N_4608,N_4413,N_4344);
nor U4609 (N_4609,N_4425,N_4398);
or U4610 (N_4610,N_4356,N_4307);
nand U4611 (N_4611,N_4433,N_4415);
nand U4612 (N_4612,N_4390,N_4373);
and U4613 (N_4613,N_4365,N_4349);
nand U4614 (N_4614,N_4385,N_4264);
nor U4615 (N_4615,N_4499,N_4340);
xor U4616 (N_4616,N_4386,N_4476);
nand U4617 (N_4617,N_4426,N_4350);
and U4618 (N_4618,N_4446,N_4456);
or U4619 (N_4619,N_4442,N_4400);
and U4620 (N_4620,N_4405,N_4409);
or U4621 (N_4621,N_4361,N_4480);
nor U4622 (N_4622,N_4366,N_4455);
and U4623 (N_4623,N_4434,N_4478);
nor U4624 (N_4624,N_4266,N_4298);
nand U4625 (N_4625,N_4251,N_4412);
nand U4626 (N_4626,N_4293,N_4334);
nand U4627 (N_4627,N_4490,N_4402);
nand U4628 (N_4628,N_4371,N_4300);
or U4629 (N_4629,N_4293,N_4310);
or U4630 (N_4630,N_4396,N_4450);
nor U4631 (N_4631,N_4494,N_4365);
nand U4632 (N_4632,N_4429,N_4317);
and U4633 (N_4633,N_4457,N_4405);
xor U4634 (N_4634,N_4252,N_4382);
xor U4635 (N_4635,N_4309,N_4468);
xnor U4636 (N_4636,N_4368,N_4498);
nand U4637 (N_4637,N_4407,N_4305);
and U4638 (N_4638,N_4468,N_4423);
and U4639 (N_4639,N_4439,N_4387);
nor U4640 (N_4640,N_4341,N_4415);
nand U4641 (N_4641,N_4414,N_4275);
or U4642 (N_4642,N_4470,N_4489);
or U4643 (N_4643,N_4492,N_4335);
and U4644 (N_4644,N_4292,N_4430);
nand U4645 (N_4645,N_4479,N_4283);
or U4646 (N_4646,N_4471,N_4435);
and U4647 (N_4647,N_4474,N_4428);
xnor U4648 (N_4648,N_4486,N_4280);
and U4649 (N_4649,N_4312,N_4354);
nor U4650 (N_4650,N_4433,N_4341);
nor U4651 (N_4651,N_4491,N_4281);
nand U4652 (N_4652,N_4307,N_4330);
xor U4653 (N_4653,N_4490,N_4268);
nor U4654 (N_4654,N_4359,N_4262);
nand U4655 (N_4655,N_4365,N_4305);
xor U4656 (N_4656,N_4380,N_4318);
nand U4657 (N_4657,N_4292,N_4424);
and U4658 (N_4658,N_4346,N_4303);
nor U4659 (N_4659,N_4274,N_4431);
xor U4660 (N_4660,N_4412,N_4285);
or U4661 (N_4661,N_4316,N_4455);
or U4662 (N_4662,N_4316,N_4345);
nor U4663 (N_4663,N_4376,N_4458);
xnor U4664 (N_4664,N_4493,N_4302);
nor U4665 (N_4665,N_4325,N_4492);
xor U4666 (N_4666,N_4366,N_4398);
or U4667 (N_4667,N_4429,N_4340);
and U4668 (N_4668,N_4336,N_4348);
and U4669 (N_4669,N_4350,N_4408);
nor U4670 (N_4670,N_4253,N_4285);
xnor U4671 (N_4671,N_4276,N_4380);
xnor U4672 (N_4672,N_4445,N_4482);
and U4673 (N_4673,N_4281,N_4376);
nand U4674 (N_4674,N_4452,N_4449);
or U4675 (N_4675,N_4289,N_4285);
xor U4676 (N_4676,N_4407,N_4289);
nand U4677 (N_4677,N_4259,N_4418);
xnor U4678 (N_4678,N_4380,N_4429);
and U4679 (N_4679,N_4453,N_4399);
nor U4680 (N_4680,N_4285,N_4480);
or U4681 (N_4681,N_4287,N_4253);
nand U4682 (N_4682,N_4490,N_4262);
nand U4683 (N_4683,N_4412,N_4327);
and U4684 (N_4684,N_4253,N_4277);
xor U4685 (N_4685,N_4272,N_4474);
nor U4686 (N_4686,N_4363,N_4385);
xnor U4687 (N_4687,N_4253,N_4494);
or U4688 (N_4688,N_4273,N_4250);
nor U4689 (N_4689,N_4418,N_4471);
xor U4690 (N_4690,N_4480,N_4302);
nand U4691 (N_4691,N_4314,N_4455);
or U4692 (N_4692,N_4446,N_4259);
xor U4693 (N_4693,N_4317,N_4382);
xor U4694 (N_4694,N_4278,N_4370);
or U4695 (N_4695,N_4456,N_4298);
nor U4696 (N_4696,N_4317,N_4493);
nor U4697 (N_4697,N_4364,N_4420);
and U4698 (N_4698,N_4291,N_4279);
nor U4699 (N_4699,N_4304,N_4458);
nand U4700 (N_4700,N_4380,N_4432);
xnor U4701 (N_4701,N_4457,N_4277);
and U4702 (N_4702,N_4452,N_4294);
nor U4703 (N_4703,N_4399,N_4384);
nand U4704 (N_4704,N_4433,N_4295);
xnor U4705 (N_4705,N_4356,N_4495);
or U4706 (N_4706,N_4291,N_4322);
xnor U4707 (N_4707,N_4380,N_4446);
nor U4708 (N_4708,N_4324,N_4284);
and U4709 (N_4709,N_4378,N_4420);
and U4710 (N_4710,N_4339,N_4372);
nor U4711 (N_4711,N_4312,N_4250);
and U4712 (N_4712,N_4260,N_4267);
nand U4713 (N_4713,N_4267,N_4339);
nor U4714 (N_4714,N_4283,N_4298);
or U4715 (N_4715,N_4274,N_4317);
nand U4716 (N_4716,N_4484,N_4481);
or U4717 (N_4717,N_4470,N_4367);
or U4718 (N_4718,N_4431,N_4353);
nor U4719 (N_4719,N_4278,N_4477);
nor U4720 (N_4720,N_4397,N_4303);
xnor U4721 (N_4721,N_4442,N_4350);
xor U4722 (N_4722,N_4445,N_4419);
or U4723 (N_4723,N_4398,N_4447);
nor U4724 (N_4724,N_4311,N_4297);
and U4725 (N_4725,N_4441,N_4295);
and U4726 (N_4726,N_4435,N_4419);
and U4727 (N_4727,N_4280,N_4341);
nor U4728 (N_4728,N_4364,N_4407);
and U4729 (N_4729,N_4461,N_4399);
xnor U4730 (N_4730,N_4282,N_4380);
xor U4731 (N_4731,N_4488,N_4376);
nand U4732 (N_4732,N_4272,N_4479);
and U4733 (N_4733,N_4476,N_4438);
or U4734 (N_4734,N_4258,N_4375);
and U4735 (N_4735,N_4444,N_4476);
xnor U4736 (N_4736,N_4329,N_4403);
or U4737 (N_4737,N_4375,N_4406);
nand U4738 (N_4738,N_4380,N_4455);
xnor U4739 (N_4739,N_4415,N_4410);
or U4740 (N_4740,N_4424,N_4250);
and U4741 (N_4741,N_4289,N_4398);
xor U4742 (N_4742,N_4355,N_4380);
nor U4743 (N_4743,N_4405,N_4431);
nand U4744 (N_4744,N_4344,N_4338);
and U4745 (N_4745,N_4469,N_4425);
nor U4746 (N_4746,N_4484,N_4350);
nor U4747 (N_4747,N_4387,N_4415);
nand U4748 (N_4748,N_4425,N_4252);
or U4749 (N_4749,N_4287,N_4252);
xnor U4750 (N_4750,N_4684,N_4586);
nand U4751 (N_4751,N_4693,N_4533);
and U4752 (N_4752,N_4673,N_4737);
nand U4753 (N_4753,N_4590,N_4719);
nand U4754 (N_4754,N_4720,N_4568);
and U4755 (N_4755,N_4744,N_4747);
or U4756 (N_4756,N_4717,N_4553);
nor U4757 (N_4757,N_4502,N_4599);
nor U4758 (N_4758,N_4598,N_4635);
nor U4759 (N_4759,N_4594,N_4540);
nor U4760 (N_4760,N_4708,N_4709);
and U4761 (N_4761,N_4541,N_4581);
xnor U4762 (N_4762,N_4560,N_4734);
or U4763 (N_4763,N_4608,N_4703);
nor U4764 (N_4764,N_4680,N_4542);
nor U4765 (N_4765,N_4710,N_4707);
xor U4766 (N_4766,N_4668,N_4582);
nor U4767 (N_4767,N_4517,N_4531);
or U4768 (N_4768,N_4733,N_4704);
nand U4769 (N_4769,N_4624,N_4548);
nor U4770 (N_4770,N_4577,N_4549);
xnor U4771 (N_4771,N_4666,N_4551);
nand U4772 (N_4772,N_4529,N_4605);
xor U4773 (N_4773,N_4652,N_4596);
and U4774 (N_4774,N_4539,N_4735);
nand U4775 (N_4775,N_4535,N_4514);
and U4776 (N_4776,N_4524,N_4676);
or U4777 (N_4777,N_4600,N_4626);
and U4778 (N_4778,N_4623,N_4567);
xnor U4779 (N_4779,N_4730,N_4595);
nor U4780 (N_4780,N_4534,N_4593);
xnor U4781 (N_4781,N_4739,N_4715);
nor U4782 (N_4782,N_4736,N_4667);
xnor U4783 (N_4783,N_4711,N_4573);
or U4784 (N_4784,N_4543,N_4697);
nor U4785 (N_4785,N_4681,N_4616);
xor U4786 (N_4786,N_4569,N_4654);
or U4787 (N_4787,N_4724,N_4741);
and U4788 (N_4788,N_4634,N_4674);
nand U4789 (N_4789,N_4660,N_4618);
xnor U4790 (N_4790,N_4546,N_4523);
nand U4791 (N_4791,N_4562,N_4686);
and U4792 (N_4792,N_4547,N_4503);
and U4793 (N_4793,N_4658,N_4507);
or U4794 (N_4794,N_4748,N_4669);
nand U4795 (N_4795,N_4613,N_4558);
and U4796 (N_4796,N_4525,N_4550);
xor U4797 (N_4797,N_4638,N_4633);
nand U4798 (N_4798,N_4572,N_4677);
nand U4799 (N_4799,N_4530,N_4636);
nor U4800 (N_4800,N_4665,N_4500);
nand U4801 (N_4801,N_4506,N_4611);
and U4802 (N_4802,N_4504,N_4563);
nor U4803 (N_4803,N_4629,N_4725);
nand U4804 (N_4804,N_4688,N_4555);
or U4805 (N_4805,N_4589,N_4587);
nor U4806 (N_4806,N_4661,N_4682);
xor U4807 (N_4807,N_4538,N_4509);
and U4808 (N_4808,N_4726,N_4557);
or U4809 (N_4809,N_4585,N_4700);
nor U4810 (N_4810,N_4544,N_4645);
and U4811 (N_4811,N_4716,N_4640);
nand U4812 (N_4812,N_4511,N_4526);
xnor U4813 (N_4813,N_4625,N_4699);
nor U4814 (N_4814,N_4537,N_4713);
or U4815 (N_4815,N_4721,N_4631);
xnor U4816 (N_4816,N_4646,N_4678);
and U4817 (N_4817,N_4642,N_4722);
xnor U4818 (N_4818,N_4718,N_4662);
or U4819 (N_4819,N_4612,N_4643);
nor U4820 (N_4820,N_4727,N_4580);
or U4821 (N_4821,N_4628,N_4584);
xor U4822 (N_4822,N_4651,N_4692);
nand U4823 (N_4823,N_4649,N_4519);
and U4824 (N_4824,N_4655,N_4691);
nor U4825 (N_4825,N_4632,N_4728);
and U4826 (N_4826,N_4664,N_4565);
and U4827 (N_4827,N_4644,N_4556);
nor U4828 (N_4828,N_4588,N_4576);
nor U4829 (N_4829,N_4621,N_4670);
xnor U4830 (N_4830,N_4513,N_4650);
nor U4831 (N_4831,N_4657,N_4592);
and U4832 (N_4832,N_4731,N_4687);
nand U4833 (N_4833,N_4685,N_4653);
or U4834 (N_4834,N_4714,N_4749);
or U4835 (N_4835,N_4518,N_4515);
xnor U4836 (N_4836,N_4663,N_4679);
nor U4837 (N_4837,N_4604,N_4740);
xnor U4838 (N_4838,N_4610,N_4706);
xor U4839 (N_4839,N_4561,N_4723);
nor U4840 (N_4840,N_4528,N_4505);
xor U4841 (N_4841,N_4602,N_4570);
or U4842 (N_4842,N_4620,N_4702);
xnor U4843 (N_4843,N_4532,N_4579);
or U4844 (N_4844,N_4705,N_4630);
nand U4845 (N_4845,N_4641,N_4637);
xnor U4846 (N_4846,N_4571,N_4552);
nor U4847 (N_4847,N_4619,N_4745);
xnor U4848 (N_4848,N_4508,N_4564);
xnor U4849 (N_4849,N_4566,N_4574);
nand U4850 (N_4850,N_4583,N_4554);
nor U4851 (N_4851,N_4578,N_4696);
nand U4852 (N_4852,N_4656,N_4683);
nand U4853 (N_4853,N_4671,N_4520);
nand U4854 (N_4854,N_4732,N_4742);
nor U4855 (N_4855,N_4659,N_4672);
nand U4856 (N_4856,N_4575,N_4607);
nand U4857 (N_4857,N_4510,N_4738);
nor U4858 (N_4858,N_4701,N_4512);
and U4859 (N_4859,N_4545,N_4712);
nor U4860 (N_4860,N_4648,N_4746);
nor U4861 (N_4861,N_4617,N_4603);
and U4862 (N_4862,N_4527,N_4694);
nor U4863 (N_4863,N_4689,N_4647);
xor U4864 (N_4864,N_4627,N_4606);
xnor U4865 (N_4865,N_4614,N_4522);
xor U4866 (N_4866,N_4601,N_4675);
nand U4867 (N_4867,N_4516,N_4622);
nand U4868 (N_4868,N_4609,N_4591);
or U4869 (N_4869,N_4536,N_4559);
or U4870 (N_4870,N_4729,N_4597);
nand U4871 (N_4871,N_4501,N_4698);
nand U4872 (N_4872,N_4743,N_4639);
nor U4873 (N_4873,N_4521,N_4690);
nand U4874 (N_4874,N_4615,N_4695);
nor U4875 (N_4875,N_4519,N_4665);
nor U4876 (N_4876,N_4598,N_4504);
and U4877 (N_4877,N_4697,N_4674);
nand U4878 (N_4878,N_4566,N_4604);
nor U4879 (N_4879,N_4500,N_4617);
xor U4880 (N_4880,N_4549,N_4520);
xnor U4881 (N_4881,N_4710,N_4539);
and U4882 (N_4882,N_4509,N_4638);
xnor U4883 (N_4883,N_4530,N_4647);
nor U4884 (N_4884,N_4590,N_4661);
or U4885 (N_4885,N_4665,N_4511);
and U4886 (N_4886,N_4536,N_4736);
xnor U4887 (N_4887,N_4609,N_4726);
and U4888 (N_4888,N_4511,N_4519);
and U4889 (N_4889,N_4682,N_4739);
xor U4890 (N_4890,N_4504,N_4585);
nand U4891 (N_4891,N_4643,N_4668);
or U4892 (N_4892,N_4547,N_4565);
nand U4893 (N_4893,N_4575,N_4590);
or U4894 (N_4894,N_4624,N_4608);
xor U4895 (N_4895,N_4619,N_4689);
nand U4896 (N_4896,N_4641,N_4596);
or U4897 (N_4897,N_4677,N_4595);
or U4898 (N_4898,N_4548,N_4667);
nand U4899 (N_4899,N_4650,N_4645);
nand U4900 (N_4900,N_4521,N_4620);
xor U4901 (N_4901,N_4550,N_4710);
nor U4902 (N_4902,N_4738,N_4569);
xnor U4903 (N_4903,N_4711,N_4690);
or U4904 (N_4904,N_4523,N_4607);
and U4905 (N_4905,N_4678,N_4504);
nand U4906 (N_4906,N_4703,N_4696);
and U4907 (N_4907,N_4562,N_4681);
xnor U4908 (N_4908,N_4589,N_4727);
nand U4909 (N_4909,N_4602,N_4552);
and U4910 (N_4910,N_4707,N_4709);
and U4911 (N_4911,N_4574,N_4737);
nor U4912 (N_4912,N_4696,N_4653);
and U4913 (N_4913,N_4553,N_4646);
xnor U4914 (N_4914,N_4641,N_4744);
xor U4915 (N_4915,N_4696,N_4589);
nand U4916 (N_4916,N_4508,N_4565);
or U4917 (N_4917,N_4511,N_4694);
xnor U4918 (N_4918,N_4601,N_4551);
nand U4919 (N_4919,N_4648,N_4599);
nand U4920 (N_4920,N_4640,N_4550);
and U4921 (N_4921,N_4650,N_4627);
nor U4922 (N_4922,N_4733,N_4626);
and U4923 (N_4923,N_4571,N_4640);
and U4924 (N_4924,N_4549,N_4681);
or U4925 (N_4925,N_4564,N_4661);
nor U4926 (N_4926,N_4702,N_4598);
xor U4927 (N_4927,N_4613,N_4538);
and U4928 (N_4928,N_4692,N_4721);
xor U4929 (N_4929,N_4636,N_4669);
nor U4930 (N_4930,N_4724,N_4547);
or U4931 (N_4931,N_4694,N_4721);
nand U4932 (N_4932,N_4708,N_4524);
or U4933 (N_4933,N_4690,N_4519);
nand U4934 (N_4934,N_4560,N_4638);
or U4935 (N_4935,N_4573,N_4663);
or U4936 (N_4936,N_4648,N_4663);
nor U4937 (N_4937,N_4674,N_4616);
nand U4938 (N_4938,N_4716,N_4606);
xor U4939 (N_4939,N_4705,N_4729);
nor U4940 (N_4940,N_4748,N_4649);
and U4941 (N_4941,N_4595,N_4723);
xnor U4942 (N_4942,N_4534,N_4578);
xor U4943 (N_4943,N_4594,N_4601);
and U4944 (N_4944,N_4503,N_4674);
nor U4945 (N_4945,N_4738,N_4718);
xor U4946 (N_4946,N_4653,N_4525);
xnor U4947 (N_4947,N_4540,N_4734);
or U4948 (N_4948,N_4622,N_4512);
and U4949 (N_4949,N_4528,N_4715);
xnor U4950 (N_4950,N_4553,N_4580);
and U4951 (N_4951,N_4578,N_4682);
and U4952 (N_4952,N_4568,N_4749);
nor U4953 (N_4953,N_4515,N_4664);
nor U4954 (N_4954,N_4515,N_4747);
or U4955 (N_4955,N_4521,N_4596);
and U4956 (N_4956,N_4603,N_4552);
or U4957 (N_4957,N_4524,N_4593);
or U4958 (N_4958,N_4556,N_4580);
or U4959 (N_4959,N_4566,N_4551);
or U4960 (N_4960,N_4675,N_4534);
nor U4961 (N_4961,N_4621,N_4529);
xnor U4962 (N_4962,N_4716,N_4570);
and U4963 (N_4963,N_4530,N_4540);
or U4964 (N_4964,N_4584,N_4618);
and U4965 (N_4965,N_4656,N_4745);
nand U4966 (N_4966,N_4651,N_4592);
and U4967 (N_4967,N_4737,N_4682);
nand U4968 (N_4968,N_4501,N_4657);
nor U4969 (N_4969,N_4619,N_4556);
and U4970 (N_4970,N_4608,N_4660);
xnor U4971 (N_4971,N_4509,N_4629);
and U4972 (N_4972,N_4696,N_4574);
xor U4973 (N_4973,N_4556,N_4700);
xor U4974 (N_4974,N_4618,N_4524);
nand U4975 (N_4975,N_4736,N_4524);
or U4976 (N_4976,N_4647,N_4533);
nand U4977 (N_4977,N_4566,N_4658);
or U4978 (N_4978,N_4687,N_4724);
and U4979 (N_4979,N_4659,N_4719);
nand U4980 (N_4980,N_4548,N_4645);
and U4981 (N_4981,N_4673,N_4574);
xnor U4982 (N_4982,N_4718,N_4619);
nand U4983 (N_4983,N_4621,N_4595);
xnor U4984 (N_4984,N_4668,N_4749);
and U4985 (N_4985,N_4659,N_4741);
nor U4986 (N_4986,N_4533,N_4701);
or U4987 (N_4987,N_4734,N_4648);
nand U4988 (N_4988,N_4653,N_4559);
and U4989 (N_4989,N_4613,N_4589);
and U4990 (N_4990,N_4532,N_4631);
and U4991 (N_4991,N_4531,N_4707);
and U4992 (N_4992,N_4573,N_4702);
xnor U4993 (N_4993,N_4584,N_4624);
or U4994 (N_4994,N_4551,N_4558);
nand U4995 (N_4995,N_4737,N_4581);
or U4996 (N_4996,N_4747,N_4577);
and U4997 (N_4997,N_4603,N_4532);
or U4998 (N_4998,N_4517,N_4603);
or U4999 (N_4999,N_4598,N_4748);
and U5000 (N_5000,N_4967,N_4988);
nor U5001 (N_5001,N_4911,N_4809);
nor U5002 (N_5002,N_4774,N_4974);
nand U5003 (N_5003,N_4814,N_4892);
nand U5004 (N_5004,N_4796,N_4833);
and U5005 (N_5005,N_4884,N_4922);
xnor U5006 (N_5006,N_4785,N_4782);
nor U5007 (N_5007,N_4812,N_4894);
or U5008 (N_5008,N_4961,N_4835);
nor U5009 (N_5009,N_4890,N_4818);
nand U5010 (N_5010,N_4760,N_4834);
xnor U5011 (N_5011,N_4813,N_4994);
and U5012 (N_5012,N_4979,N_4925);
xnor U5013 (N_5013,N_4764,N_4982);
xnor U5014 (N_5014,N_4879,N_4829);
and U5015 (N_5015,N_4975,N_4986);
nor U5016 (N_5016,N_4940,N_4987);
nor U5017 (N_5017,N_4827,N_4870);
or U5018 (N_5018,N_4969,N_4895);
nor U5019 (N_5019,N_4877,N_4897);
nor U5020 (N_5020,N_4968,N_4807);
and U5021 (N_5021,N_4886,N_4959);
or U5022 (N_5022,N_4995,N_4946);
xnor U5023 (N_5023,N_4784,N_4871);
or U5024 (N_5024,N_4921,N_4917);
nor U5025 (N_5025,N_4849,N_4786);
or U5026 (N_5026,N_4855,N_4865);
nand U5027 (N_5027,N_4866,N_4965);
and U5028 (N_5028,N_4938,N_4878);
or U5029 (N_5029,N_4773,N_4953);
nor U5030 (N_5030,N_4904,N_4983);
xor U5031 (N_5031,N_4989,N_4758);
nand U5032 (N_5032,N_4929,N_4984);
xnor U5033 (N_5033,N_4816,N_4920);
and U5034 (N_5034,N_4950,N_4930);
nand U5035 (N_5035,N_4841,N_4873);
and U5036 (N_5036,N_4932,N_4956);
nand U5037 (N_5037,N_4781,N_4757);
or U5038 (N_5038,N_4811,N_4838);
nand U5039 (N_5039,N_4880,N_4863);
and U5040 (N_5040,N_4963,N_4952);
and U5041 (N_5041,N_4903,N_4822);
or U5042 (N_5042,N_4945,N_4859);
or U5043 (N_5043,N_4913,N_4862);
and U5044 (N_5044,N_4820,N_4875);
nor U5045 (N_5045,N_4836,N_4750);
and U5046 (N_5046,N_4957,N_4798);
and U5047 (N_5047,N_4991,N_4896);
nand U5048 (N_5048,N_4900,N_4815);
or U5049 (N_5049,N_4867,N_4847);
nand U5050 (N_5050,N_4964,N_4848);
nor U5051 (N_5051,N_4935,N_4850);
nand U5052 (N_5052,N_4891,N_4864);
xnor U5053 (N_5053,N_4936,N_4985);
nor U5054 (N_5054,N_4759,N_4810);
or U5055 (N_5055,N_4845,N_4804);
and U5056 (N_5056,N_4977,N_4797);
or U5057 (N_5057,N_4902,N_4909);
or U5058 (N_5058,N_4801,N_4844);
xor U5059 (N_5059,N_4860,N_4934);
nand U5060 (N_5060,N_4825,N_4876);
nand U5061 (N_5061,N_4944,N_4830);
nand U5062 (N_5062,N_4787,N_4996);
and U5063 (N_5063,N_4800,N_4752);
or U5064 (N_5064,N_4923,N_4916);
or U5065 (N_5065,N_4802,N_4772);
or U5066 (N_5066,N_4762,N_4771);
and U5067 (N_5067,N_4924,N_4931);
or U5068 (N_5068,N_4881,N_4861);
or U5069 (N_5069,N_4980,N_4839);
xor U5070 (N_5070,N_4793,N_4933);
and U5071 (N_5071,N_4888,N_4868);
or U5072 (N_5072,N_4978,N_4853);
xnor U5073 (N_5073,N_4778,N_4831);
or U5074 (N_5074,N_4817,N_4966);
or U5075 (N_5075,N_4779,N_4768);
xnor U5076 (N_5076,N_4790,N_4914);
or U5077 (N_5077,N_4981,N_4958);
nand U5078 (N_5078,N_4887,N_4898);
xnor U5079 (N_5079,N_4872,N_4842);
nor U5080 (N_5080,N_4908,N_4854);
nand U5081 (N_5081,N_4840,N_4949);
or U5082 (N_5082,N_4756,N_4776);
nor U5083 (N_5083,N_4972,N_4766);
nor U5084 (N_5084,N_4954,N_4795);
nor U5085 (N_5085,N_4918,N_4828);
or U5086 (N_5086,N_4928,N_4973);
and U5087 (N_5087,N_4955,N_4791);
nand U5088 (N_5088,N_4769,N_4803);
nand U5089 (N_5089,N_4885,N_4780);
xnor U5090 (N_5090,N_4927,N_4837);
nand U5091 (N_5091,N_4832,N_4754);
or U5092 (N_5092,N_4856,N_4824);
xor U5093 (N_5093,N_4788,N_4883);
nand U5094 (N_5094,N_4775,N_4857);
xnor U5095 (N_5095,N_4789,N_4767);
and U5096 (N_5096,N_4926,N_4751);
nand U5097 (N_5097,N_4947,N_4858);
nor U5098 (N_5098,N_4765,N_4970);
and U5099 (N_5099,N_4821,N_4889);
and U5100 (N_5100,N_4951,N_4819);
and U5101 (N_5101,N_4971,N_4901);
and U5102 (N_5102,N_4843,N_4794);
nand U5103 (N_5103,N_4948,N_4808);
or U5104 (N_5104,N_4937,N_4846);
nand U5105 (N_5105,N_4905,N_4806);
nor U5106 (N_5106,N_4906,N_4792);
xnor U5107 (N_5107,N_4997,N_4826);
nor U5108 (N_5108,N_4869,N_4939);
nor U5109 (N_5109,N_4874,N_4999);
and U5110 (N_5110,N_4915,N_4893);
or U5111 (N_5111,N_4976,N_4960);
and U5112 (N_5112,N_4993,N_4942);
xor U5113 (N_5113,N_4941,N_4990);
nor U5114 (N_5114,N_4777,N_4770);
or U5115 (N_5115,N_4755,N_4799);
nand U5116 (N_5116,N_4919,N_4882);
and U5117 (N_5117,N_4907,N_4992);
nor U5118 (N_5118,N_4910,N_4753);
nand U5119 (N_5119,N_4761,N_4783);
or U5120 (N_5120,N_4943,N_4852);
xor U5121 (N_5121,N_4962,N_4912);
xor U5122 (N_5122,N_4823,N_4805);
or U5123 (N_5123,N_4998,N_4763);
xor U5124 (N_5124,N_4899,N_4851);
or U5125 (N_5125,N_4910,N_4856);
and U5126 (N_5126,N_4755,N_4789);
and U5127 (N_5127,N_4959,N_4869);
and U5128 (N_5128,N_4923,N_4978);
or U5129 (N_5129,N_4796,N_4886);
and U5130 (N_5130,N_4880,N_4836);
or U5131 (N_5131,N_4959,N_4824);
nand U5132 (N_5132,N_4882,N_4832);
xor U5133 (N_5133,N_4928,N_4882);
nand U5134 (N_5134,N_4858,N_4984);
and U5135 (N_5135,N_4864,N_4784);
nand U5136 (N_5136,N_4767,N_4900);
nand U5137 (N_5137,N_4890,N_4816);
or U5138 (N_5138,N_4865,N_4934);
nor U5139 (N_5139,N_4909,N_4964);
nor U5140 (N_5140,N_4816,N_4839);
nor U5141 (N_5141,N_4940,N_4911);
and U5142 (N_5142,N_4795,N_4816);
and U5143 (N_5143,N_4891,N_4827);
and U5144 (N_5144,N_4965,N_4987);
and U5145 (N_5145,N_4833,N_4822);
and U5146 (N_5146,N_4846,N_4858);
and U5147 (N_5147,N_4761,N_4759);
nand U5148 (N_5148,N_4987,N_4784);
nor U5149 (N_5149,N_4799,N_4894);
or U5150 (N_5150,N_4768,N_4776);
or U5151 (N_5151,N_4820,N_4962);
xor U5152 (N_5152,N_4944,N_4985);
nor U5153 (N_5153,N_4806,N_4855);
nand U5154 (N_5154,N_4810,N_4907);
nor U5155 (N_5155,N_4756,N_4898);
and U5156 (N_5156,N_4889,N_4971);
or U5157 (N_5157,N_4770,N_4875);
and U5158 (N_5158,N_4818,N_4853);
or U5159 (N_5159,N_4988,N_4912);
nand U5160 (N_5160,N_4903,N_4938);
and U5161 (N_5161,N_4940,N_4950);
or U5162 (N_5162,N_4860,N_4859);
and U5163 (N_5163,N_4993,N_4808);
nand U5164 (N_5164,N_4914,N_4928);
xnor U5165 (N_5165,N_4921,N_4777);
xor U5166 (N_5166,N_4857,N_4880);
and U5167 (N_5167,N_4922,N_4880);
nor U5168 (N_5168,N_4870,N_4915);
and U5169 (N_5169,N_4956,N_4816);
and U5170 (N_5170,N_4969,N_4912);
nor U5171 (N_5171,N_4922,N_4799);
or U5172 (N_5172,N_4824,N_4989);
or U5173 (N_5173,N_4930,N_4922);
nor U5174 (N_5174,N_4934,N_4782);
xor U5175 (N_5175,N_4966,N_4860);
nor U5176 (N_5176,N_4907,N_4984);
nand U5177 (N_5177,N_4959,N_4813);
or U5178 (N_5178,N_4869,N_4821);
and U5179 (N_5179,N_4927,N_4919);
nor U5180 (N_5180,N_4960,N_4910);
xor U5181 (N_5181,N_4988,N_4797);
nor U5182 (N_5182,N_4904,N_4891);
nand U5183 (N_5183,N_4965,N_4980);
xor U5184 (N_5184,N_4822,N_4783);
xor U5185 (N_5185,N_4998,N_4788);
nand U5186 (N_5186,N_4850,N_4832);
nand U5187 (N_5187,N_4917,N_4922);
xor U5188 (N_5188,N_4786,N_4937);
and U5189 (N_5189,N_4834,N_4918);
xor U5190 (N_5190,N_4763,N_4760);
xnor U5191 (N_5191,N_4929,N_4895);
and U5192 (N_5192,N_4887,N_4829);
or U5193 (N_5193,N_4910,N_4758);
and U5194 (N_5194,N_4925,N_4908);
nor U5195 (N_5195,N_4895,N_4881);
nand U5196 (N_5196,N_4998,N_4774);
xnor U5197 (N_5197,N_4912,N_4977);
and U5198 (N_5198,N_4863,N_4967);
or U5199 (N_5199,N_4812,N_4920);
nor U5200 (N_5200,N_4771,N_4895);
xor U5201 (N_5201,N_4989,N_4785);
or U5202 (N_5202,N_4858,N_4944);
xor U5203 (N_5203,N_4959,N_4864);
xor U5204 (N_5204,N_4848,N_4854);
nand U5205 (N_5205,N_4810,N_4961);
nor U5206 (N_5206,N_4874,N_4842);
xnor U5207 (N_5207,N_4792,N_4810);
xnor U5208 (N_5208,N_4751,N_4969);
nand U5209 (N_5209,N_4840,N_4986);
xor U5210 (N_5210,N_4841,N_4954);
and U5211 (N_5211,N_4883,N_4936);
nand U5212 (N_5212,N_4873,N_4781);
xor U5213 (N_5213,N_4833,N_4948);
or U5214 (N_5214,N_4924,N_4846);
nand U5215 (N_5215,N_4871,N_4954);
nand U5216 (N_5216,N_4958,N_4920);
or U5217 (N_5217,N_4925,N_4862);
nand U5218 (N_5218,N_4782,N_4927);
and U5219 (N_5219,N_4952,N_4831);
or U5220 (N_5220,N_4923,N_4836);
xor U5221 (N_5221,N_4759,N_4790);
or U5222 (N_5222,N_4750,N_4990);
nor U5223 (N_5223,N_4807,N_4998);
nor U5224 (N_5224,N_4938,N_4797);
or U5225 (N_5225,N_4951,N_4824);
and U5226 (N_5226,N_4855,N_4781);
nor U5227 (N_5227,N_4982,N_4860);
xnor U5228 (N_5228,N_4845,N_4762);
and U5229 (N_5229,N_4951,N_4948);
nor U5230 (N_5230,N_4993,N_4881);
nor U5231 (N_5231,N_4825,N_4861);
or U5232 (N_5232,N_4757,N_4992);
or U5233 (N_5233,N_4810,N_4994);
xor U5234 (N_5234,N_4833,N_4813);
or U5235 (N_5235,N_4902,N_4764);
xnor U5236 (N_5236,N_4814,N_4757);
xor U5237 (N_5237,N_4886,N_4830);
or U5238 (N_5238,N_4782,N_4876);
nand U5239 (N_5239,N_4774,N_4833);
nor U5240 (N_5240,N_4858,N_4889);
or U5241 (N_5241,N_4868,N_4857);
nand U5242 (N_5242,N_4825,N_4881);
xnor U5243 (N_5243,N_4880,N_4911);
nand U5244 (N_5244,N_4938,N_4920);
and U5245 (N_5245,N_4828,N_4953);
or U5246 (N_5246,N_4925,N_4847);
nand U5247 (N_5247,N_4918,N_4763);
xor U5248 (N_5248,N_4777,N_4896);
and U5249 (N_5249,N_4867,N_4833);
nand U5250 (N_5250,N_5198,N_5035);
xor U5251 (N_5251,N_5082,N_5170);
and U5252 (N_5252,N_5167,N_5138);
nor U5253 (N_5253,N_5133,N_5107);
nor U5254 (N_5254,N_5234,N_5128);
nor U5255 (N_5255,N_5010,N_5227);
nor U5256 (N_5256,N_5049,N_5076);
nand U5257 (N_5257,N_5193,N_5201);
xnor U5258 (N_5258,N_5117,N_5226);
nand U5259 (N_5259,N_5143,N_5245);
and U5260 (N_5260,N_5023,N_5142);
or U5261 (N_5261,N_5194,N_5085);
and U5262 (N_5262,N_5109,N_5174);
or U5263 (N_5263,N_5052,N_5043);
xnor U5264 (N_5264,N_5209,N_5086);
or U5265 (N_5265,N_5146,N_5233);
xor U5266 (N_5266,N_5092,N_5057);
or U5267 (N_5267,N_5077,N_5215);
xor U5268 (N_5268,N_5047,N_5009);
and U5269 (N_5269,N_5243,N_5205);
or U5270 (N_5270,N_5235,N_5157);
or U5271 (N_5271,N_5025,N_5195);
xnor U5272 (N_5272,N_5229,N_5132);
xnor U5273 (N_5273,N_5131,N_5074);
and U5274 (N_5274,N_5207,N_5061);
or U5275 (N_5275,N_5248,N_5161);
xor U5276 (N_5276,N_5098,N_5064);
xor U5277 (N_5277,N_5137,N_5213);
nand U5278 (N_5278,N_5181,N_5055);
nor U5279 (N_5279,N_5091,N_5104);
nor U5280 (N_5280,N_5017,N_5134);
and U5281 (N_5281,N_5136,N_5217);
or U5282 (N_5282,N_5220,N_5225);
and U5283 (N_5283,N_5185,N_5040);
nand U5284 (N_5284,N_5176,N_5216);
or U5285 (N_5285,N_5066,N_5056);
xnor U5286 (N_5286,N_5121,N_5173);
nand U5287 (N_5287,N_5051,N_5059);
nor U5288 (N_5288,N_5200,N_5007);
xnor U5289 (N_5289,N_5154,N_5027);
and U5290 (N_5290,N_5171,N_5011);
or U5291 (N_5291,N_5046,N_5116);
or U5292 (N_5292,N_5097,N_5089);
nor U5293 (N_5293,N_5060,N_5018);
nand U5294 (N_5294,N_5165,N_5054);
nand U5295 (N_5295,N_5124,N_5189);
and U5296 (N_5296,N_5166,N_5048);
xor U5297 (N_5297,N_5041,N_5102);
or U5298 (N_5298,N_5030,N_5210);
xor U5299 (N_5299,N_5223,N_5214);
and U5300 (N_5300,N_5062,N_5184);
and U5301 (N_5301,N_5021,N_5228);
nand U5302 (N_5302,N_5212,N_5083);
nor U5303 (N_5303,N_5087,N_5172);
nand U5304 (N_5304,N_5020,N_5242);
xor U5305 (N_5305,N_5094,N_5148);
and U5306 (N_5306,N_5179,N_5079);
nor U5307 (N_5307,N_5065,N_5150);
and U5308 (N_5308,N_5140,N_5081);
nor U5309 (N_5309,N_5151,N_5152);
nor U5310 (N_5310,N_5034,N_5208);
or U5311 (N_5311,N_5203,N_5202);
xor U5312 (N_5312,N_5111,N_5036);
nand U5313 (N_5313,N_5247,N_5178);
and U5314 (N_5314,N_5113,N_5101);
xnor U5315 (N_5315,N_5069,N_5114);
xnor U5316 (N_5316,N_5053,N_5112);
nor U5317 (N_5317,N_5067,N_5110);
and U5318 (N_5318,N_5099,N_5168);
or U5319 (N_5319,N_5115,N_5045);
nand U5320 (N_5320,N_5032,N_5096);
xor U5321 (N_5321,N_5125,N_5028);
xor U5322 (N_5322,N_5003,N_5037);
xnor U5323 (N_5323,N_5177,N_5105);
or U5324 (N_5324,N_5015,N_5050);
nor U5325 (N_5325,N_5080,N_5000);
xor U5326 (N_5326,N_5163,N_5159);
xor U5327 (N_5327,N_5162,N_5070);
or U5328 (N_5328,N_5224,N_5204);
nand U5329 (N_5329,N_5218,N_5249);
or U5330 (N_5330,N_5175,N_5002);
nor U5331 (N_5331,N_5001,N_5239);
xnor U5332 (N_5332,N_5129,N_5183);
xnor U5333 (N_5333,N_5237,N_5044);
xor U5334 (N_5334,N_5240,N_5093);
nor U5335 (N_5335,N_5187,N_5068);
and U5336 (N_5336,N_5095,N_5130);
or U5337 (N_5337,N_5108,N_5197);
or U5338 (N_5338,N_5126,N_5004);
or U5339 (N_5339,N_5206,N_5075);
nand U5340 (N_5340,N_5024,N_5156);
nand U5341 (N_5341,N_5238,N_5182);
or U5342 (N_5342,N_5013,N_5190);
nand U5343 (N_5343,N_5016,N_5158);
or U5344 (N_5344,N_5244,N_5100);
and U5345 (N_5345,N_5031,N_5231);
and U5346 (N_5346,N_5122,N_5006);
nor U5347 (N_5347,N_5008,N_5120);
nor U5348 (N_5348,N_5232,N_5145);
nor U5349 (N_5349,N_5219,N_5058);
nand U5350 (N_5350,N_5236,N_5144);
nor U5351 (N_5351,N_5135,N_5127);
or U5352 (N_5352,N_5147,N_5119);
nor U5353 (N_5353,N_5063,N_5078);
xnor U5354 (N_5354,N_5196,N_5139);
or U5355 (N_5355,N_5088,N_5222);
xor U5356 (N_5356,N_5019,N_5033);
or U5357 (N_5357,N_5153,N_5039);
nand U5358 (N_5358,N_5106,N_5191);
and U5359 (N_5359,N_5160,N_5155);
xor U5360 (N_5360,N_5042,N_5123);
and U5361 (N_5361,N_5221,N_5246);
nand U5362 (N_5362,N_5073,N_5012);
nand U5363 (N_5363,N_5005,N_5072);
nand U5364 (N_5364,N_5192,N_5103);
nand U5365 (N_5365,N_5090,N_5230);
and U5366 (N_5366,N_5038,N_5118);
or U5367 (N_5367,N_5149,N_5186);
xor U5368 (N_5368,N_5199,N_5169);
nand U5369 (N_5369,N_5141,N_5029);
nand U5370 (N_5370,N_5014,N_5026);
or U5371 (N_5371,N_5084,N_5022);
and U5372 (N_5372,N_5164,N_5180);
xnor U5373 (N_5373,N_5071,N_5241);
nor U5374 (N_5374,N_5188,N_5211);
or U5375 (N_5375,N_5239,N_5230);
xnor U5376 (N_5376,N_5062,N_5080);
xor U5377 (N_5377,N_5110,N_5015);
nand U5378 (N_5378,N_5248,N_5133);
xor U5379 (N_5379,N_5180,N_5085);
nor U5380 (N_5380,N_5097,N_5056);
nor U5381 (N_5381,N_5168,N_5222);
nor U5382 (N_5382,N_5185,N_5088);
or U5383 (N_5383,N_5182,N_5243);
and U5384 (N_5384,N_5058,N_5207);
xnor U5385 (N_5385,N_5005,N_5043);
xnor U5386 (N_5386,N_5241,N_5115);
nand U5387 (N_5387,N_5035,N_5146);
or U5388 (N_5388,N_5158,N_5133);
nor U5389 (N_5389,N_5133,N_5230);
or U5390 (N_5390,N_5006,N_5038);
xor U5391 (N_5391,N_5136,N_5165);
nand U5392 (N_5392,N_5203,N_5090);
nor U5393 (N_5393,N_5233,N_5119);
nor U5394 (N_5394,N_5108,N_5063);
or U5395 (N_5395,N_5065,N_5111);
nor U5396 (N_5396,N_5169,N_5093);
xnor U5397 (N_5397,N_5011,N_5232);
or U5398 (N_5398,N_5175,N_5061);
nor U5399 (N_5399,N_5091,N_5192);
xnor U5400 (N_5400,N_5127,N_5148);
nor U5401 (N_5401,N_5025,N_5234);
nor U5402 (N_5402,N_5147,N_5042);
nor U5403 (N_5403,N_5194,N_5018);
and U5404 (N_5404,N_5126,N_5010);
and U5405 (N_5405,N_5188,N_5183);
or U5406 (N_5406,N_5032,N_5131);
nand U5407 (N_5407,N_5039,N_5116);
or U5408 (N_5408,N_5030,N_5141);
and U5409 (N_5409,N_5083,N_5026);
nand U5410 (N_5410,N_5208,N_5152);
nor U5411 (N_5411,N_5039,N_5232);
nand U5412 (N_5412,N_5171,N_5068);
and U5413 (N_5413,N_5178,N_5159);
and U5414 (N_5414,N_5023,N_5189);
or U5415 (N_5415,N_5130,N_5004);
and U5416 (N_5416,N_5193,N_5167);
and U5417 (N_5417,N_5044,N_5235);
nand U5418 (N_5418,N_5231,N_5017);
xor U5419 (N_5419,N_5166,N_5228);
and U5420 (N_5420,N_5052,N_5226);
or U5421 (N_5421,N_5072,N_5207);
nor U5422 (N_5422,N_5232,N_5072);
and U5423 (N_5423,N_5148,N_5157);
or U5424 (N_5424,N_5137,N_5205);
xnor U5425 (N_5425,N_5009,N_5225);
nor U5426 (N_5426,N_5113,N_5076);
and U5427 (N_5427,N_5180,N_5030);
nand U5428 (N_5428,N_5019,N_5059);
and U5429 (N_5429,N_5048,N_5226);
nor U5430 (N_5430,N_5073,N_5110);
nor U5431 (N_5431,N_5089,N_5144);
nand U5432 (N_5432,N_5089,N_5153);
xnor U5433 (N_5433,N_5013,N_5016);
nor U5434 (N_5434,N_5054,N_5143);
or U5435 (N_5435,N_5082,N_5141);
and U5436 (N_5436,N_5049,N_5197);
nand U5437 (N_5437,N_5188,N_5019);
nor U5438 (N_5438,N_5088,N_5216);
nand U5439 (N_5439,N_5198,N_5217);
xor U5440 (N_5440,N_5249,N_5171);
nand U5441 (N_5441,N_5065,N_5202);
or U5442 (N_5442,N_5042,N_5247);
nand U5443 (N_5443,N_5127,N_5054);
and U5444 (N_5444,N_5060,N_5233);
or U5445 (N_5445,N_5050,N_5224);
nor U5446 (N_5446,N_5136,N_5071);
or U5447 (N_5447,N_5004,N_5029);
nor U5448 (N_5448,N_5199,N_5193);
nand U5449 (N_5449,N_5167,N_5011);
and U5450 (N_5450,N_5126,N_5015);
nor U5451 (N_5451,N_5094,N_5038);
nor U5452 (N_5452,N_5190,N_5129);
xor U5453 (N_5453,N_5127,N_5205);
nor U5454 (N_5454,N_5202,N_5030);
nand U5455 (N_5455,N_5001,N_5157);
xnor U5456 (N_5456,N_5143,N_5031);
nor U5457 (N_5457,N_5030,N_5025);
nor U5458 (N_5458,N_5010,N_5206);
nor U5459 (N_5459,N_5240,N_5095);
xor U5460 (N_5460,N_5026,N_5060);
and U5461 (N_5461,N_5031,N_5208);
or U5462 (N_5462,N_5229,N_5175);
or U5463 (N_5463,N_5027,N_5129);
xnor U5464 (N_5464,N_5201,N_5054);
nand U5465 (N_5465,N_5098,N_5089);
nor U5466 (N_5466,N_5211,N_5152);
or U5467 (N_5467,N_5144,N_5181);
or U5468 (N_5468,N_5182,N_5144);
nand U5469 (N_5469,N_5114,N_5178);
or U5470 (N_5470,N_5088,N_5214);
xor U5471 (N_5471,N_5179,N_5124);
nand U5472 (N_5472,N_5098,N_5050);
or U5473 (N_5473,N_5161,N_5154);
xor U5474 (N_5474,N_5081,N_5165);
nand U5475 (N_5475,N_5021,N_5172);
and U5476 (N_5476,N_5151,N_5189);
and U5477 (N_5477,N_5246,N_5105);
xor U5478 (N_5478,N_5081,N_5152);
or U5479 (N_5479,N_5013,N_5125);
and U5480 (N_5480,N_5111,N_5092);
or U5481 (N_5481,N_5074,N_5144);
xor U5482 (N_5482,N_5196,N_5149);
and U5483 (N_5483,N_5249,N_5239);
nor U5484 (N_5484,N_5087,N_5110);
or U5485 (N_5485,N_5217,N_5111);
and U5486 (N_5486,N_5201,N_5089);
nand U5487 (N_5487,N_5061,N_5031);
and U5488 (N_5488,N_5128,N_5202);
nor U5489 (N_5489,N_5105,N_5139);
nand U5490 (N_5490,N_5101,N_5201);
and U5491 (N_5491,N_5054,N_5059);
xor U5492 (N_5492,N_5070,N_5078);
and U5493 (N_5493,N_5179,N_5058);
xor U5494 (N_5494,N_5154,N_5217);
nand U5495 (N_5495,N_5110,N_5063);
nor U5496 (N_5496,N_5198,N_5158);
or U5497 (N_5497,N_5036,N_5180);
nor U5498 (N_5498,N_5085,N_5184);
nor U5499 (N_5499,N_5151,N_5026);
nor U5500 (N_5500,N_5324,N_5265);
and U5501 (N_5501,N_5311,N_5411);
nand U5502 (N_5502,N_5337,N_5384);
nor U5503 (N_5503,N_5330,N_5454);
nor U5504 (N_5504,N_5395,N_5284);
xnor U5505 (N_5505,N_5262,N_5362);
and U5506 (N_5506,N_5427,N_5313);
xor U5507 (N_5507,N_5470,N_5278);
nand U5508 (N_5508,N_5336,N_5279);
nor U5509 (N_5509,N_5309,N_5436);
nand U5510 (N_5510,N_5486,N_5351);
or U5511 (N_5511,N_5349,N_5301);
xor U5512 (N_5512,N_5267,N_5342);
or U5513 (N_5513,N_5438,N_5251);
xnor U5514 (N_5514,N_5338,N_5302);
nor U5515 (N_5515,N_5449,N_5271);
and U5516 (N_5516,N_5442,N_5408);
nor U5517 (N_5517,N_5396,N_5425);
or U5518 (N_5518,N_5382,N_5264);
and U5519 (N_5519,N_5333,N_5319);
nor U5520 (N_5520,N_5308,N_5266);
nand U5521 (N_5521,N_5322,N_5418);
or U5522 (N_5522,N_5318,N_5364);
nor U5523 (N_5523,N_5482,N_5376);
nand U5524 (N_5524,N_5433,N_5498);
or U5525 (N_5525,N_5441,N_5355);
nand U5526 (N_5526,N_5466,N_5378);
nand U5527 (N_5527,N_5399,N_5401);
or U5528 (N_5528,N_5463,N_5276);
and U5529 (N_5529,N_5310,N_5413);
nor U5530 (N_5530,N_5306,N_5422);
and U5531 (N_5531,N_5312,N_5406);
xnor U5532 (N_5532,N_5492,N_5256);
and U5533 (N_5533,N_5494,N_5440);
xnor U5534 (N_5534,N_5457,N_5424);
and U5535 (N_5535,N_5331,N_5367);
and U5536 (N_5536,N_5260,N_5314);
nand U5537 (N_5537,N_5393,N_5426);
or U5538 (N_5538,N_5334,N_5460);
nand U5539 (N_5539,N_5476,N_5405);
and U5540 (N_5540,N_5446,N_5471);
xor U5541 (N_5541,N_5431,N_5285);
or U5542 (N_5542,N_5356,N_5277);
nand U5543 (N_5543,N_5327,N_5300);
nand U5544 (N_5544,N_5295,N_5381);
nand U5545 (N_5545,N_5432,N_5372);
xor U5546 (N_5546,N_5347,N_5430);
nand U5547 (N_5547,N_5478,N_5315);
or U5548 (N_5548,N_5400,N_5473);
nor U5549 (N_5549,N_5445,N_5451);
xor U5550 (N_5550,N_5412,N_5472);
nor U5551 (N_5551,N_5257,N_5402);
or U5552 (N_5552,N_5409,N_5496);
xnor U5553 (N_5553,N_5281,N_5495);
xnor U5554 (N_5554,N_5345,N_5350);
nor U5555 (N_5555,N_5286,N_5386);
or U5556 (N_5556,N_5272,N_5294);
nand U5557 (N_5557,N_5428,N_5283);
and U5558 (N_5558,N_5299,N_5371);
or U5559 (N_5559,N_5488,N_5484);
and U5560 (N_5560,N_5465,N_5453);
nor U5561 (N_5561,N_5250,N_5398);
and U5562 (N_5562,N_5369,N_5415);
or U5563 (N_5563,N_5291,N_5481);
nand U5564 (N_5564,N_5489,N_5417);
nor U5565 (N_5565,N_5363,N_5305);
nand U5566 (N_5566,N_5335,N_5332);
and U5567 (N_5567,N_5448,N_5435);
nor U5568 (N_5568,N_5307,N_5490);
nand U5569 (N_5569,N_5274,N_5293);
nor U5570 (N_5570,N_5447,N_5370);
xor U5571 (N_5571,N_5290,N_5353);
nor U5572 (N_5572,N_5467,N_5464);
nor U5573 (N_5573,N_5358,N_5298);
nand U5574 (N_5574,N_5258,N_5456);
and U5575 (N_5575,N_5416,N_5474);
xnor U5576 (N_5576,N_5329,N_5420);
nor U5577 (N_5577,N_5361,N_5468);
nand U5578 (N_5578,N_5374,N_5304);
xnor U5579 (N_5579,N_5317,N_5377);
nor U5580 (N_5580,N_5491,N_5387);
xor U5581 (N_5581,N_5270,N_5357);
and U5582 (N_5582,N_5388,N_5423);
xnor U5583 (N_5583,N_5323,N_5275);
and U5584 (N_5584,N_5344,N_5414);
xor U5585 (N_5585,N_5288,N_5485);
and U5586 (N_5586,N_5343,N_5380);
xnor U5587 (N_5587,N_5366,N_5254);
nor U5588 (N_5588,N_5443,N_5487);
nor U5589 (N_5589,N_5316,N_5352);
nand U5590 (N_5590,N_5469,N_5493);
or U5591 (N_5591,N_5499,N_5346);
or U5592 (N_5592,N_5391,N_5253);
or U5593 (N_5593,N_5383,N_5282);
xnor U5594 (N_5594,N_5475,N_5373);
and U5595 (N_5595,N_5297,N_5348);
or U5596 (N_5596,N_5263,N_5434);
nor U5597 (N_5597,N_5365,N_5410);
or U5598 (N_5598,N_5497,N_5479);
or U5599 (N_5599,N_5341,N_5392);
and U5600 (N_5600,N_5407,N_5403);
nand U5601 (N_5601,N_5444,N_5390);
nand U5602 (N_5602,N_5452,N_5320);
nor U5603 (N_5603,N_5268,N_5325);
xor U5604 (N_5604,N_5261,N_5439);
or U5605 (N_5605,N_5328,N_5477);
nor U5606 (N_5606,N_5269,N_5375);
and U5607 (N_5607,N_5360,N_5385);
nand U5608 (N_5608,N_5404,N_5455);
nor U5609 (N_5609,N_5397,N_5394);
or U5610 (N_5610,N_5321,N_5354);
and U5611 (N_5611,N_5480,N_5289);
nor U5612 (N_5612,N_5287,N_5461);
xor U5613 (N_5613,N_5296,N_5458);
xor U5614 (N_5614,N_5339,N_5437);
and U5615 (N_5615,N_5389,N_5368);
and U5616 (N_5616,N_5359,N_5273);
nor U5617 (N_5617,N_5429,N_5379);
and U5618 (N_5618,N_5419,N_5421);
and U5619 (N_5619,N_5459,N_5326);
nor U5620 (N_5620,N_5450,N_5462);
and U5621 (N_5621,N_5303,N_5252);
nand U5622 (N_5622,N_5255,N_5259);
or U5623 (N_5623,N_5483,N_5340);
xnor U5624 (N_5624,N_5280,N_5292);
xor U5625 (N_5625,N_5310,N_5276);
nand U5626 (N_5626,N_5416,N_5392);
nand U5627 (N_5627,N_5441,N_5254);
and U5628 (N_5628,N_5386,N_5382);
nor U5629 (N_5629,N_5380,N_5314);
and U5630 (N_5630,N_5438,N_5332);
nand U5631 (N_5631,N_5269,N_5327);
nor U5632 (N_5632,N_5457,N_5410);
or U5633 (N_5633,N_5319,N_5274);
xor U5634 (N_5634,N_5378,N_5293);
nand U5635 (N_5635,N_5389,N_5350);
and U5636 (N_5636,N_5472,N_5302);
or U5637 (N_5637,N_5454,N_5352);
and U5638 (N_5638,N_5371,N_5378);
xnor U5639 (N_5639,N_5259,N_5438);
nand U5640 (N_5640,N_5447,N_5358);
and U5641 (N_5641,N_5413,N_5458);
nand U5642 (N_5642,N_5458,N_5305);
or U5643 (N_5643,N_5461,N_5402);
nand U5644 (N_5644,N_5353,N_5314);
or U5645 (N_5645,N_5418,N_5473);
xor U5646 (N_5646,N_5267,N_5482);
nand U5647 (N_5647,N_5325,N_5427);
and U5648 (N_5648,N_5314,N_5482);
nand U5649 (N_5649,N_5308,N_5353);
and U5650 (N_5650,N_5478,N_5394);
xor U5651 (N_5651,N_5278,N_5300);
or U5652 (N_5652,N_5469,N_5377);
or U5653 (N_5653,N_5284,N_5463);
nor U5654 (N_5654,N_5282,N_5493);
nor U5655 (N_5655,N_5487,N_5372);
and U5656 (N_5656,N_5353,N_5320);
xnor U5657 (N_5657,N_5432,N_5477);
nand U5658 (N_5658,N_5255,N_5412);
or U5659 (N_5659,N_5436,N_5281);
and U5660 (N_5660,N_5437,N_5383);
and U5661 (N_5661,N_5270,N_5329);
nand U5662 (N_5662,N_5416,N_5437);
nand U5663 (N_5663,N_5426,N_5475);
xor U5664 (N_5664,N_5299,N_5262);
or U5665 (N_5665,N_5328,N_5356);
and U5666 (N_5666,N_5306,N_5488);
or U5667 (N_5667,N_5387,N_5449);
nand U5668 (N_5668,N_5464,N_5457);
and U5669 (N_5669,N_5388,N_5442);
and U5670 (N_5670,N_5469,N_5302);
nor U5671 (N_5671,N_5317,N_5366);
xnor U5672 (N_5672,N_5430,N_5405);
nor U5673 (N_5673,N_5480,N_5461);
nor U5674 (N_5674,N_5497,N_5491);
nand U5675 (N_5675,N_5260,N_5277);
xnor U5676 (N_5676,N_5329,N_5407);
nand U5677 (N_5677,N_5448,N_5370);
xor U5678 (N_5678,N_5483,N_5253);
nor U5679 (N_5679,N_5389,N_5378);
or U5680 (N_5680,N_5470,N_5261);
nand U5681 (N_5681,N_5448,N_5350);
and U5682 (N_5682,N_5281,N_5350);
nand U5683 (N_5683,N_5360,N_5437);
nand U5684 (N_5684,N_5398,N_5426);
nor U5685 (N_5685,N_5312,N_5262);
nand U5686 (N_5686,N_5288,N_5297);
xnor U5687 (N_5687,N_5293,N_5374);
nand U5688 (N_5688,N_5425,N_5402);
and U5689 (N_5689,N_5310,N_5274);
or U5690 (N_5690,N_5317,N_5277);
or U5691 (N_5691,N_5261,N_5263);
xor U5692 (N_5692,N_5268,N_5491);
and U5693 (N_5693,N_5260,N_5275);
or U5694 (N_5694,N_5258,N_5441);
nor U5695 (N_5695,N_5433,N_5304);
xor U5696 (N_5696,N_5296,N_5415);
nand U5697 (N_5697,N_5312,N_5401);
or U5698 (N_5698,N_5402,N_5449);
nand U5699 (N_5699,N_5385,N_5452);
and U5700 (N_5700,N_5497,N_5451);
and U5701 (N_5701,N_5274,N_5400);
nand U5702 (N_5702,N_5291,N_5473);
xnor U5703 (N_5703,N_5285,N_5499);
xor U5704 (N_5704,N_5401,N_5396);
or U5705 (N_5705,N_5273,N_5488);
or U5706 (N_5706,N_5368,N_5387);
nor U5707 (N_5707,N_5454,N_5396);
or U5708 (N_5708,N_5365,N_5267);
and U5709 (N_5709,N_5286,N_5289);
or U5710 (N_5710,N_5347,N_5486);
xnor U5711 (N_5711,N_5356,N_5337);
nand U5712 (N_5712,N_5374,N_5265);
xor U5713 (N_5713,N_5255,N_5338);
or U5714 (N_5714,N_5350,N_5482);
xor U5715 (N_5715,N_5498,N_5366);
nand U5716 (N_5716,N_5274,N_5288);
and U5717 (N_5717,N_5354,N_5424);
xor U5718 (N_5718,N_5333,N_5496);
xor U5719 (N_5719,N_5383,N_5499);
or U5720 (N_5720,N_5402,N_5279);
nand U5721 (N_5721,N_5267,N_5394);
nor U5722 (N_5722,N_5352,N_5432);
and U5723 (N_5723,N_5339,N_5427);
nor U5724 (N_5724,N_5492,N_5310);
nand U5725 (N_5725,N_5306,N_5469);
nor U5726 (N_5726,N_5474,N_5264);
or U5727 (N_5727,N_5258,N_5370);
nor U5728 (N_5728,N_5286,N_5353);
xnor U5729 (N_5729,N_5466,N_5483);
xnor U5730 (N_5730,N_5401,N_5280);
nand U5731 (N_5731,N_5426,N_5305);
and U5732 (N_5732,N_5478,N_5385);
nor U5733 (N_5733,N_5294,N_5251);
xor U5734 (N_5734,N_5358,N_5375);
and U5735 (N_5735,N_5327,N_5409);
xnor U5736 (N_5736,N_5308,N_5407);
and U5737 (N_5737,N_5315,N_5370);
or U5738 (N_5738,N_5282,N_5473);
or U5739 (N_5739,N_5352,N_5376);
and U5740 (N_5740,N_5479,N_5421);
xnor U5741 (N_5741,N_5348,N_5338);
xnor U5742 (N_5742,N_5464,N_5378);
nand U5743 (N_5743,N_5442,N_5425);
or U5744 (N_5744,N_5479,N_5467);
and U5745 (N_5745,N_5379,N_5272);
nand U5746 (N_5746,N_5442,N_5435);
nand U5747 (N_5747,N_5345,N_5261);
nor U5748 (N_5748,N_5442,N_5477);
xnor U5749 (N_5749,N_5430,N_5461);
nor U5750 (N_5750,N_5689,N_5676);
or U5751 (N_5751,N_5609,N_5554);
and U5752 (N_5752,N_5693,N_5647);
or U5753 (N_5753,N_5734,N_5748);
nor U5754 (N_5754,N_5532,N_5736);
or U5755 (N_5755,N_5721,N_5747);
xnor U5756 (N_5756,N_5688,N_5691);
and U5757 (N_5757,N_5615,N_5530);
xor U5758 (N_5758,N_5509,N_5616);
nand U5759 (N_5759,N_5719,N_5524);
or U5760 (N_5760,N_5670,N_5522);
and U5761 (N_5761,N_5610,N_5656);
nor U5762 (N_5762,N_5588,N_5675);
nand U5763 (N_5763,N_5646,N_5660);
nor U5764 (N_5764,N_5744,N_5537);
or U5765 (N_5765,N_5683,N_5669);
nand U5766 (N_5766,N_5644,N_5692);
xnor U5767 (N_5767,N_5504,N_5582);
or U5768 (N_5768,N_5513,N_5624);
nand U5769 (N_5769,N_5584,N_5533);
and U5770 (N_5770,N_5686,N_5722);
nand U5771 (N_5771,N_5601,N_5711);
xor U5772 (N_5772,N_5694,N_5743);
and U5773 (N_5773,N_5724,N_5506);
nand U5774 (N_5774,N_5529,N_5502);
nor U5775 (N_5775,N_5632,N_5617);
nand U5776 (N_5776,N_5710,N_5673);
nand U5777 (N_5777,N_5643,N_5668);
nand U5778 (N_5778,N_5561,N_5514);
nor U5779 (N_5779,N_5505,N_5542);
and U5780 (N_5780,N_5745,N_5574);
nand U5781 (N_5781,N_5629,N_5709);
xnor U5782 (N_5782,N_5706,N_5742);
nand U5783 (N_5783,N_5515,N_5528);
or U5784 (N_5784,N_5720,N_5550);
xor U5785 (N_5785,N_5690,N_5685);
nor U5786 (N_5786,N_5600,N_5557);
xnor U5787 (N_5787,N_5679,N_5575);
or U5788 (N_5788,N_5592,N_5746);
and U5789 (N_5789,N_5612,N_5732);
nor U5790 (N_5790,N_5671,N_5526);
and U5791 (N_5791,N_5593,N_5531);
nor U5792 (N_5792,N_5568,N_5520);
nand U5793 (N_5793,N_5687,N_5594);
xnor U5794 (N_5794,N_5635,N_5587);
nor U5795 (N_5795,N_5697,N_5651);
nand U5796 (N_5796,N_5628,N_5716);
and U5797 (N_5797,N_5738,N_5603);
nor U5798 (N_5798,N_5649,N_5645);
nor U5799 (N_5799,N_5712,N_5641);
and U5800 (N_5800,N_5549,N_5726);
nand U5801 (N_5801,N_5698,N_5637);
nor U5802 (N_5802,N_5555,N_5700);
and U5803 (N_5803,N_5604,N_5614);
nor U5804 (N_5804,N_5715,N_5562);
xnor U5805 (N_5805,N_5666,N_5541);
xnor U5806 (N_5806,N_5538,N_5563);
nor U5807 (N_5807,N_5662,N_5701);
nor U5808 (N_5808,N_5639,N_5512);
xnor U5809 (N_5809,N_5739,N_5625);
or U5810 (N_5810,N_5717,N_5525);
nor U5811 (N_5811,N_5519,N_5606);
nand U5812 (N_5812,N_5567,N_5730);
or U5813 (N_5813,N_5684,N_5579);
and U5814 (N_5814,N_5611,N_5523);
nor U5815 (N_5815,N_5544,N_5677);
xnor U5816 (N_5816,N_5503,N_5672);
or U5817 (N_5817,N_5718,N_5620);
and U5818 (N_5818,N_5626,N_5634);
or U5819 (N_5819,N_5546,N_5590);
and U5820 (N_5820,N_5652,N_5558);
and U5821 (N_5821,N_5501,N_5725);
or U5822 (N_5822,N_5545,N_5619);
xnor U5823 (N_5823,N_5569,N_5605);
nand U5824 (N_5824,N_5714,N_5566);
and U5825 (N_5825,N_5723,N_5571);
nor U5826 (N_5826,N_5681,N_5613);
nand U5827 (N_5827,N_5572,N_5729);
and U5828 (N_5828,N_5543,N_5705);
nor U5829 (N_5829,N_5713,N_5699);
xnor U5830 (N_5830,N_5680,N_5642);
nor U5831 (N_5831,N_5573,N_5648);
nor U5832 (N_5832,N_5682,N_5535);
and U5833 (N_5833,N_5508,N_5622);
or U5834 (N_5834,N_5728,N_5663);
xor U5835 (N_5835,N_5507,N_5536);
or U5836 (N_5836,N_5565,N_5581);
nor U5837 (N_5837,N_5551,N_5577);
nand U5838 (N_5838,N_5727,N_5703);
nor U5839 (N_5839,N_5560,N_5517);
xor U5840 (N_5840,N_5578,N_5657);
and U5841 (N_5841,N_5586,N_5589);
nand U5842 (N_5842,N_5638,N_5595);
xor U5843 (N_5843,N_5500,N_5598);
nor U5844 (N_5844,N_5534,N_5591);
and U5845 (N_5845,N_5731,N_5627);
and U5846 (N_5846,N_5596,N_5655);
or U5847 (N_5847,N_5602,N_5640);
and U5848 (N_5848,N_5695,N_5704);
nor U5849 (N_5849,N_5665,N_5553);
xor U5850 (N_5850,N_5678,N_5597);
xor U5851 (N_5851,N_5552,N_5631);
xnor U5852 (N_5852,N_5696,N_5608);
nor U5853 (N_5853,N_5659,N_5548);
nor U5854 (N_5854,N_5702,N_5516);
and U5855 (N_5855,N_5576,N_5607);
and U5856 (N_5856,N_5599,N_5559);
and U5857 (N_5857,N_5580,N_5667);
or U5858 (N_5858,N_5737,N_5664);
nor U5859 (N_5859,N_5564,N_5653);
or U5860 (N_5860,N_5658,N_5661);
and U5861 (N_5861,N_5510,N_5633);
nand U5862 (N_5862,N_5556,N_5636);
nor U5863 (N_5863,N_5585,N_5735);
xnor U5864 (N_5864,N_5741,N_5740);
nor U5865 (N_5865,N_5527,N_5511);
nand U5866 (N_5866,N_5630,N_5539);
and U5867 (N_5867,N_5621,N_5623);
and U5868 (N_5868,N_5708,N_5749);
nor U5869 (N_5869,N_5654,N_5733);
nand U5870 (N_5870,N_5707,N_5618);
nand U5871 (N_5871,N_5521,N_5540);
and U5872 (N_5872,N_5518,N_5570);
and U5873 (N_5873,N_5650,N_5547);
xnor U5874 (N_5874,N_5674,N_5583);
nor U5875 (N_5875,N_5500,N_5745);
xor U5876 (N_5876,N_5689,N_5647);
and U5877 (N_5877,N_5678,N_5728);
nand U5878 (N_5878,N_5714,N_5703);
or U5879 (N_5879,N_5511,N_5559);
or U5880 (N_5880,N_5518,N_5583);
nor U5881 (N_5881,N_5667,N_5725);
nand U5882 (N_5882,N_5507,N_5735);
and U5883 (N_5883,N_5527,N_5605);
nand U5884 (N_5884,N_5532,N_5618);
and U5885 (N_5885,N_5679,N_5501);
or U5886 (N_5886,N_5647,N_5529);
xor U5887 (N_5887,N_5645,N_5683);
or U5888 (N_5888,N_5717,N_5514);
nor U5889 (N_5889,N_5640,N_5679);
or U5890 (N_5890,N_5639,N_5748);
or U5891 (N_5891,N_5510,N_5531);
nand U5892 (N_5892,N_5549,N_5545);
and U5893 (N_5893,N_5546,N_5531);
and U5894 (N_5894,N_5573,N_5601);
and U5895 (N_5895,N_5630,N_5722);
xnor U5896 (N_5896,N_5523,N_5746);
nand U5897 (N_5897,N_5636,N_5502);
nand U5898 (N_5898,N_5549,N_5604);
and U5899 (N_5899,N_5623,N_5509);
or U5900 (N_5900,N_5615,N_5617);
nand U5901 (N_5901,N_5709,N_5512);
nand U5902 (N_5902,N_5573,N_5739);
nand U5903 (N_5903,N_5618,N_5637);
or U5904 (N_5904,N_5640,N_5518);
xor U5905 (N_5905,N_5715,N_5698);
nand U5906 (N_5906,N_5697,N_5535);
or U5907 (N_5907,N_5509,N_5536);
and U5908 (N_5908,N_5734,N_5537);
and U5909 (N_5909,N_5746,N_5654);
nor U5910 (N_5910,N_5620,N_5572);
and U5911 (N_5911,N_5666,N_5551);
nand U5912 (N_5912,N_5653,N_5580);
nand U5913 (N_5913,N_5612,N_5739);
nor U5914 (N_5914,N_5636,N_5571);
xnor U5915 (N_5915,N_5647,N_5739);
xnor U5916 (N_5916,N_5521,N_5732);
or U5917 (N_5917,N_5590,N_5554);
nand U5918 (N_5918,N_5676,N_5592);
nor U5919 (N_5919,N_5749,N_5679);
or U5920 (N_5920,N_5606,N_5694);
nand U5921 (N_5921,N_5572,N_5671);
nand U5922 (N_5922,N_5748,N_5733);
nand U5923 (N_5923,N_5557,N_5609);
and U5924 (N_5924,N_5695,N_5658);
or U5925 (N_5925,N_5620,N_5566);
nor U5926 (N_5926,N_5698,N_5626);
nor U5927 (N_5927,N_5644,N_5700);
nand U5928 (N_5928,N_5740,N_5701);
nor U5929 (N_5929,N_5587,N_5737);
nor U5930 (N_5930,N_5556,N_5739);
and U5931 (N_5931,N_5748,N_5552);
xor U5932 (N_5932,N_5630,N_5730);
and U5933 (N_5933,N_5526,N_5725);
and U5934 (N_5934,N_5589,N_5720);
nor U5935 (N_5935,N_5688,N_5638);
xnor U5936 (N_5936,N_5576,N_5570);
nand U5937 (N_5937,N_5716,N_5529);
and U5938 (N_5938,N_5639,N_5623);
nor U5939 (N_5939,N_5701,N_5505);
or U5940 (N_5940,N_5509,N_5621);
nor U5941 (N_5941,N_5646,N_5506);
nor U5942 (N_5942,N_5716,N_5597);
nor U5943 (N_5943,N_5732,N_5619);
nand U5944 (N_5944,N_5537,N_5664);
and U5945 (N_5945,N_5577,N_5583);
and U5946 (N_5946,N_5711,N_5657);
nand U5947 (N_5947,N_5582,N_5679);
xor U5948 (N_5948,N_5540,N_5657);
xor U5949 (N_5949,N_5721,N_5590);
nand U5950 (N_5950,N_5604,N_5722);
xor U5951 (N_5951,N_5535,N_5716);
or U5952 (N_5952,N_5576,N_5590);
and U5953 (N_5953,N_5608,N_5645);
or U5954 (N_5954,N_5582,N_5630);
nor U5955 (N_5955,N_5742,N_5667);
and U5956 (N_5956,N_5682,N_5586);
xnor U5957 (N_5957,N_5719,N_5544);
nand U5958 (N_5958,N_5617,N_5740);
xor U5959 (N_5959,N_5663,N_5647);
nor U5960 (N_5960,N_5744,N_5557);
nor U5961 (N_5961,N_5737,N_5565);
nand U5962 (N_5962,N_5739,N_5562);
xor U5963 (N_5963,N_5668,N_5649);
and U5964 (N_5964,N_5624,N_5561);
xnor U5965 (N_5965,N_5632,N_5607);
or U5966 (N_5966,N_5626,N_5621);
nor U5967 (N_5967,N_5673,N_5568);
or U5968 (N_5968,N_5640,N_5569);
nor U5969 (N_5969,N_5728,N_5721);
nand U5970 (N_5970,N_5501,N_5623);
nand U5971 (N_5971,N_5534,N_5732);
and U5972 (N_5972,N_5633,N_5506);
and U5973 (N_5973,N_5719,N_5691);
nand U5974 (N_5974,N_5655,N_5741);
nor U5975 (N_5975,N_5633,N_5557);
nand U5976 (N_5976,N_5729,N_5657);
or U5977 (N_5977,N_5677,N_5728);
xnor U5978 (N_5978,N_5649,N_5542);
nand U5979 (N_5979,N_5737,N_5698);
xor U5980 (N_5980,N_5571,N_5681);
and U5981 (N_5981,N_5501,N_5631);
nor U5982 (N_5982,N_5711,N_5732);
or U5983 (N_5983,N_5686,N_5640);
or U5984 (N_5984,N_5555,N_5640);
nand U5985 (N_5985,N_5582,N_5744);
nand U5986 (N_5986,N_5709,N_5674);
xor U5987 (N_5987,N_5600,N_5688);
nand U5988 (N_5988,N_5653,N_5659);
xor U5989 (N_5989,N_5603,N_5558);
or U5990 (N_5990,N_5616,N_5533);
xor U5991 (N_5991,N_5643,N_5650);
or U5992 (N_5992,N_5735,N_5595);
nor U5993 (N_5993,N_5708,N_5522);
xor U5994 (N_5994,N_5507,N_5563);
or U5995 (N_5995,N_5520,N_5719);
xnor U5996 (N_5996,N_5616,N_5545);
xnor U5997 (N_5997,N_5691,N_5749);
nor U5998 (N_5998,N_5521,N_5500);
or U5999 (N_5999,N_5541,N_5578);
nand U6000 (N_6000,N_5879,N_5924);
and U6001 (N_6001,N_5897,N_5829);
nand U6002 (N_6002,N_5997,N_5957);
xor U6003 (N_6003,N_5853,N_5914);
nor U6004 (N_6004,N_5968,N_5844);
nand U6005 (N_6005,N_5894,N_5971);
nor U6006 (N_6006,N_5799,N_5796);
nand U6007 (N_6007,N_5974,N_5870);
nand U6008 (N_6008,N_5977,N_5833);
or U6009 (N_6009,N_5826,N_5941);
xor U6010 (N_6010,N_5918,N_5795);
nor U6011 (N_6011,N_5842,N_5801);
nand U6012 (N_6012,N_5999,N_5965);
or U6013 (N_6013,N_5972,N_5828);
or U6014 (N_6014,N_5905,N_5910);
nand U6015 (N_6015,N_5919,N_5781);
and U6016 (N_6016,N_5979,N_5991);
xnor U6017 (N_6017,N_5989,N_5865);
nand U6018 (N_6018,N_5765,N_5818);
or U6019 (N_6019,N_5975,N_5877);
xor U6020 (N_6020,N_5978,N_5932);
and U6021 (N_6021,N_5774,N_5944);
or U6022 (N_6022,N_5767,N_5786);
xnor U6023 (N_6023,N_5792,N_5779);
or U6024 (N_6024,N_5955,N_5852);
or U6025 (N_6025,N_5831,N_5936);
or U6026 (N_6026,N_5804,N_5902);
xor U6027 (N_6027,N_5950,N_5836);
or U6028 (N_6028,N_5791,N_5811);
xor U6029 (N_6029,N_5827,N_5908);
nor U6030 (N_6030,N_5993,N_5817);
or U6031 (N_6031,N_5788,N_5954);
xor U6032 (N_6032,N_5899,N_5798);
nor U6033 (N_6033,N_5851,N_5784);
or U6034 (N_6034,N_5881,N_5874);
nor U6035 (N_6035,N_5893,N_5963);
xor U6036 (N_6036,N_5871,N_5901);
nand U6037 (N_6037,N_5906,N_5854);
or U6038 (N_6038,N_5940,N_5956);
xor U6039 (N_6039,N_5808,N_5922);
nand U6040 (N_6040,N_5835,N_5813);
nor U6041 (N_6041,N_5825,N_5807);
or U6042 (N_6042,N_5863,N_5888);
nor U6043 (N_6043,N_5953,N_5752);
xor U6044 (N_6044,N_5759,N_5770);
and U6045 (N_6045,N_5876,N_5857);
and U6046 (N_6046,N_5873,N_5911);
xor U6047 (N_6047,N_5772,N_5809);
nand U6048 (N_6048,N_5896,N_5937);
and U6049 (N_6049,N_5846,N_5959);
and U6050 (N_6050,N_5994,N_5960);
nor U6051 (N_6051,N_5751,N_5983);
nor U6052 (N_6052,N_5783,N_5938);
nor U6053 (N_6053,N_5878,N_5861);
nor U6054 (N_6054,N_5850,N_5821);
nand U6055 (N_6055,N_5787,N_5951);
xor U6056 (N_6056,N_5929,N_5889);
nor U6057 (N_6057,N_5970,N_5845);
nand U6058 (N_6058,N_5832,N_5921);
and U6059 (N_6059,N_5755,N_5952);
and U6060 (N_6060,N_5992,N_5802);
nand U6061 (N_6061,N_5907,N_5837);
xnor U6062 (N_6062,N_5756,N_5982);
nand U6063 (N_6063,N_5859,N_5909);
or U6064 (N_6064,N_5782,N_5976);
and U6065 (N_6065,N_5834,N_5875);
or U6066 (N_6066,N_5800,N_5754);
nor U6067 (N_6067,N_5814,N_5789);
nor U6068 (N_6068,N_5867,N_5840);
nand U6069 (N_6069,N_5860,N_5981);
nand U6070 (N_6070,N_5885,N_5947);
nor U6071 (N_6071,N_5778,N_5883);
xor U6072 (N_6072,N_5785,N_5912);
nand U6073 (N_6073,N_5880,N_5961);
nor U6074 (N_6074,N_5841,N_5856);
nand U6075 (N_6075,N_5904,N_5998);
or U6076 (N_6076,N_5987,N_5812);
and U6077 (N_6077,N_5933,N_5886);
or U6078 (N_6078,N_5771,N_5815);
nor U6079 (N_6079,N_5930,N_5864);
nand U6080 (N_6080,N_5882,N_5869);
nor U6081 (N_6081,N_5766,N_5934);
or U6082 (N_6082,N_5805,N_5872);
nand U6083 (N_6083,N_5797,N_5973);
nor U6084 (N_6084,N_5988,N_5920);
nand U6085 (N_6085,N_5773,N_5942);
xor U6086 (N_6086,N_5768,N_5927);
or U6087 (N_6087,N_5757,N_5923);
xnor U6088 (N_6088,N_5763,N_5892);
xor U6089 (N_6089,N_5887,N_5769);
xor U6090 (N_6090,N_5855,N_5898);
and U6091 (N_6091,N_5969,N_5945);
nand U6092 (N_6092,N_5843,N_5966);
nor U6093 (N_6093,N_5761,N_5780);
and U6094 (N_6094,N_5917,N_5986);
and U6095 (N_6095,N_5916,N_5868);
and U6096 (N_6096,N_5985,N_5946);
or U6097 (N_6097,N_5990,N_5900);
nor U6098 (N_6098,N_5758,N_5823);
xor U6099 (N_6099,N_5803,N_5884);
nand U6100 (N_6100,N_5806,N_5776);
xnor U6101 (N_6101,N_5764,N_5895);
xnor U6102 (N_6102,N_5949,N_5777);
nor U6103 (N_6103,N_5847,N_5931);
and U6104 (N_6104,N_5790,N_5943);
and U6105 (N_6105,N_5984,N_5948);
nor U6106 (N_6106,N_5794,N_5964);
nor U6107 (N_6107,N_5915,N_5939);
xnor U6108 (N_6108,N_5775,N_5824);
nand U6109 (N_6109,N_5819,N_5862);
nor U6110 (N_6110,N_5925,N_5849);
or U6111 (N_6111,N_5891,N_5996);
xor U6112 (N_6112,N_5858,N_5816);
and U6113 (N_6113,N_5967,N_5762);
nor U6114 (N_6114,N_5962,N_5820);
or U6115 (N_6115,N_5750,N_5958);
nand U6116 (N_6116,N_5839,N_5903);
xor U6117 (N_6117,N_5830,N_5935);
nor U6118 (N_6118,N_5928,N_5753);
or U6119 (N_6119,N_5793,N_5890);
xnor U6120 (N_6120,N_5848,N_5926);
and U6121 (N_6121,N_5810,N_5995);
and U6122 (N_6122,N_5913,N_5760);
or U6123 (N_6123,N_5838,N_5866);
and U6124 (N_6124,N_5980,N_5822);
nor U6125 (N_6125,N_5756,N_5988);
nor U6126 (N_6126,N_5939,N_5993);
or U6127 (N_6127,N_5942,N_5895);
xor U6128 (N_6128,N_5918,N_5780);
nand U6129 (N_6129,N_5917,N_5867);
nor U6130 (N_6130,N_5949,N_5917);
or U6131 (N_6131,N_5943,N_5863);
nor U6132 (N_6132,N_5959,N_5784);
and U6133 (N_6133,N_5838,N_5773);
and U6134 (N_6134,N_5863,N_5972);
nand U6135 (N_6135,N_5831,N_5928);
nand U6136 (N_6136,N_5940,N_5766);
and U6137 (N_6137,N_5888,N_5940);
nor U6138 (N_6138,N_5940,N_5921);
and U6139 (N_6139,N_5969,N_5902);
or U6140 (N_6140,N_5799,N_5897);
xnor U6141 (N_6141,N_5785,N_5978);
xnor U6142 (N_6142,N_5957,N_5920);
nand U6143 (N_6143,N_5804,N_5769);
and U6144 (N_6144,N_5752,N_5751);
nand U6145 (N_6145,N_5864,N_5845);
nor U6146 (N_6146,N_5950,N_5751);
and U6147 (N_6147,N_5760,N_5818);
or U6148 (N_6148,N_5834,N_5909);
nor U6149 (N_6149,N_5956,N_5941);
and U6150 (N_6150,N_5946,N_5796);
nor U6151 (N_6151,N_5898,N_5843);
xnor U6152 (N_6152,N_5821,N_5949);
xor U6153 (N_6153,N_5907,N_5815);
xor U6154 (N_6154,N_5866,N_5894);
and U6155 (N_6155,N_5826,N_5758);
nor U6156 (N_6156,N_5908,N_5950);
nor U6157 (N_6157,N_5793,N_5964);
and U6158 (N_6158,N_5797,N_5979);
and U6159 (N_6159,N_5860,N_5900);
xor U6160 (N_6160,N_5836,N_5862);
and U6161 (N_6161,N_5865,N_5958);
or U6162 (N_6162,N_5916,N_5982);
nand U6163 (N_6163,N_5803,N_5854);
and U6164 (N_6164,N_5804,N_5836);
nor U6165 (N_6165,N_5830,N_5928);
nor U6166 (N_6166,N_5865,N_5918);
or U6167 (N_6167,N_5972,N_5911);
nand U6168 (N_6168,N_5965,N_5868);
xnor U6169 (N_6169,N_5779,N_5998);
or U6170 (N_6170,N_5848,N_5781);
nor U6171 (N_6171,N_5939,N_5793);
nand U6172 (N_6172,N_5865,N_5857);
and U6173 (N_6173,N_5933,N_5907);
nand U6174 (N_6174,N_5890,N_5800);
nand U6175 (N_6175,N_5994,N_5764);
xor U6176 (N_6176,N_5813,N_5783);
nand U6177 (N_6177,N_5972,N_5851);
xor U6178 (N_6178,N_5875,N_5923);
nor U6179 (N_6179,N_5855,N_5937);
nor U6180 (N_6180,N_5992,N_5869);
and U6181 (N_6181,N_5999,N_5847);
or U6182 (N_6182,N_5973,N_5790);
and U6183 (N_6183,N_5823,N_5768);
nor U6184 (N_6184,N_5918,N_5752);
nand U6185 (N_6185,N_5816,N_5877);
nand U6186 (N_6186,N_5845,N_5760);
nor U6187 (N_6187,N_5874,N_5847);
xnor U6188 (N_6188,N_5838,N_5940);
or U6189 (N_6189,N_5827,N_5764);
nand U6190 (N_6190,N_5770,N_5894);
nor U6191 (N_6191,N_5757,N_5894);
nand U6192 (N_6192,N_5911,N_5877);
nor U6193 (N_6193,N_5773,N_5824);
xor U6194 (N_6194,N_5822,N_5962);
xor U6195 (N_6195,N_5785,N_5884);
xnor U6196 (N_6196,N_5881,N_5940);
and U6197 (N_6197,N_5994,N_5971);
nor U6198 (N_6198,N_5766,N_5926);
xor U6199 (N_6199,N_5970,N_5944);
nor U6200 (N_6200,N_5888,N_5790);
and U6201 (N_6201,N_5913,N_5873);
xor U6202 (N_6202,N_5918,N_5877);
or U6203 (N_6203,N_5873,N_5768);
and U6204 (N_6204,N_5873,N_5842);
or U6205 (N_6205,N_5799,N_5899);
nand U6206 (N_6206,N_5816,N_5818);
and U6207 (N_6207,N_5926,N_5942);
nor U6208 (N_6208,N_5904,N_5909);
xnor U6209 (N_6209,N_5776,N_5971);
nor U6210 (N_6210,N_5944,N_5812);
nand U6211 (N_6211,N_5956,N_5950);
or U6212 (N_6212,N_5984,N_5817);
and U6213 (N_6213,N_5927,N_5775);
or U6214 (N_6214,N_5814,N_5838);
nor U6215 (N_6215,N_5968,N_5940);
nand U6216 (N_6216,N_5927,N_5933);
xnor U6217 (N_6217,N_5758,N_5832);
nand U6218 (N_6218,N_5924,N_5906);
and U6219 (N_6219,N_5920,N_5991);
xor U6220 (N_6220,N_5917,N_5886);
and U6221 (N_6221,N_5930,N_5773);
xnor U6222 (N_6222,N_5832,N_5844);
xor U6223 (N_6223,N_5771,N_5809);
nand U6224 (N_6224,N_5854,N_5831);
or U6225 (N_6225,N_5765,N_5875);
nand U6226 (N_6226,N_5982,N_5978);
nor U6227 (N_6227,N_5813,N_5777);
or U6228 (N_6228,N_5853,N_5813);
nand U6229 (N_6229,N_5924,N_5890);
and U6230 (N_6230,N_5945,N_5929);
nand U6231 (N_6231,N_5783,N_5785);
xnor U6232 (N_6232,N_5795,N_5844);
or U6233 (N_6233,N_5850,N_5969);
and U6234 (N_6234,N_5934,N_5864);
nor U6235 (N_6235,N_5777,N_5895);
xnor U6236 (N_6236,N_5958,N_5861);
nand U6237 (N_6237,N_5813,N_5944);
nand U6238 (N_6238,N_5812,N_5980);
or U6239 (N_6239,N_5895,N_5981);
nor U6240 (N_6240,N_5887,N_5977);
xor U6241 (N_6241,N_5814,N_5783);
nor U6242 (N_6242,N_5922,N_5863);
or U6243 (N_6243,N_5934,N_5991);
nand U6244 (N_6244,N_5983,N_5826);
nand U6245 (N_6245,N_5829,N_5792);
xor U6246 (N_6246,N_5966,N_5886);
or U6247 (N_6247,N_5893,N_5923);
and U6248 (N_6248,N_5817,N_5937);
and U6249 (N_6249,N_5809,N_5896);
nor U6250 (N_6250,N_6098,N_6141);
nor U6251 (N_6251,N_6026,N_6158);
nand U6252 (N_6252,N_6202,N_6083);
nor U6253 (N_6253,N_6032,N_6213);
xnor U6254 (N_6254,N_6166,N_6063);
nand U6255 (N_6255,N_6087,N_6060);
or U6256 (N_6256,N_6221,N_6238);
xor U6257 (N_6257,N_6161,N_6006);
xor U6258 (N_6258,N_6105,N_6046);
nor U6259 (N_6259,N_6134,N_6013);
and U6260 (N_6260,N_6115,N_6057);
and U6261 (N_6261,N_6078,N_6004);
xor U6262 (N_6262,N_6206,N_6170);
nor U6263 (N_6263,N_6030,N_6076);
xor U6264 (N_6264,N_6073,N_6222);
xor U6265 (N_6265,N_6109,N_6233);
or U6266 (N_6266,N_6122,N_6173);
or U6267 (N_6267,N_6204,N_6018);
xor U6268 (N_6268,N_6138,N_6242);
nor U6269 (N_6269,N_6235,N_6090);
nor U6270 (N_6270,N_6248,N_6038);
or U6271 (N_6271,N_6097,N_6107);
and U6272 (N_6272,N_6217,N_6174);
nor U6273 (N_6273,N_6240,N_6000);
or U6274 (N_6274,N_6029,N_6082);
xnor U6275 (N_6275,N_6187,N_6081);
and U6276 (N_6276,N_6157,N_6111);
or U6277 (N_6277,N_6056,N_6080);
or U6278 (N_6278,N_6169,N_6216);
xor U6279 (N_6279,N_6153,N_6163);
and U6280 (N_6280,N_6031,N_6229);
nand U6281 (N_6281,N_6199,N_6086);
xnor U6282 (N_6282,N_6117,N_6092);
or U6283 (N_6283,N_6175,N_6033);
xnor U6284 (N_6284,N_6015,N_6214);
or U6285 (N_6285,N_6108,N_6225);
xnor U6286 (N_6286,N_6198,N_6064);
nand U6287 (N_6287,N_6041,N_6003);
nand U6288 (N_6288,N_6218,N_6118);
and U6289 (N_6289,N_6121,N_6024);
and U6290 (N_6290,N_6167,N_6223);
nand U6291 (N_6291,N_6051,N_6211);
xor U6292 (N_6292,N_6027,N_6234);
nand U6293 (N_6293,N_6093,N_6181);
xnor U6294 (N_6294,N_6089,N_6125);
nand U6295 (N_6295,N_6110,N_6106);
xnor U6296 (N_6296,N_6011,N_6022);
nand U6297 (N_6297,N_6205,N_6065);
nand U6298 (N_6298,N_6028,N_6120);
nor U6299 (N_6299,N_6084,N_6179);
nand U6300 (N_6300,N_6137,N_6094);
nand U6301 (N_6301,N_6140,N_6232);
xor U6302 (N_6302,N_6014,N_6001);
or U6303 (N_6303,N_6236,N_6247);
and U6304 (N_6304,N_6192,N_6085);
xor U6305 (N_6305,N_6207,N_6100);
xnor U6306 (N_6306,N_6184,N_6019);
nor U6307 (N_6307,N_6220,N_6127);
xnor U6308 (N_6308,N_6156,N_6178);
xor U6309 (N_6309,N_6188,N_6114);
and U6310 (N_6310,N_6196,N_6243);
and U6311 (N_6311,N_6165,N_6045);
nand U6312 (N_6312,N_6025,N_6058);
nor U6313 (N_6313,N_6129,N_6095);
nand U6314 (N_6314,N_6139,N_6145);
or U6315 (N_6315,N_6246,N_6249);
nand U6316 (N_6316,N_6146,N_6099);
nor U6317 (N_6317,N_6203,N_6164);
and U6318 (N_6318,N_6168,N_6171);
nor U6319 (N_6319,N_6124,N_6016);
nand U6320 (N_6320,N_6079,N_6112);
or U6321 (N_6321,N_6062,N_6017);
xnor U6322 (N_6322,N_6245,N_6002);
nand U6323 (N_6323,N_6209,N_6208);
and U6324 (N_6324,N_6008,N_6103);
or U6325 (N_6325,N_6005,N_6193);
xor U6326 (N_6326,N_6023,N_6009);
nand U6327 (N_6327,N_6050,N_6101);
xnor U6328 (N_6328,N_6162,N_6043);
nand U6329 (N_6329,N_6237,N_6066);
nand U6330 (N_6330,N_6104,N_6231);
or U6331 (N_6331,N_6177,N_6072);
nand U6332 (N_6332,N_6123,N_6075);
or U6333 (N_6333,N_6219,N_6067);
nand U6334 (N_6334,N_6091,N_6052);
xnor U6335 (N_6335,N_6061,N_6010);
nand U6336 (N_6336,N_6036,N_6034);
and U6337 (N_6337,N_6155,N_6088);
and U6338 (N_6338,N_6227,N_6241);
or U6339 (N_6339,N_6069,N_6096);
nand U6340 (N_6340,N_6176,N_6201);
or U6341 (N_6341,N_6197,N_6182);
nand U6342 (N_6342,N_6144,N_6186);
and U6343 (N_6343,N_6152,N_6131);
and U6344 (N_6344,N_6068,N_6035);
xnor U6345 (N_6345,N_6126,N_6074);
nor U6346 (N_6346,N_6055,N_6044);
and U6347 (N_6347,N_6135,N_6136);
nor U6348 (N_6348,N_6183,N_6012);
xor U6349 (N_6349,N_6116,N_6039);
or U6350 (N_6350,N_6071,N_6132);
or U6351 (N_6351,N_6150,N_6037);
and U6352 (N_6352,N_6151,N_6048);
xor U6353 (N_6353,N_6020,N_6021);
nor U6354 (N_6354,N_6226,N_6224);
and U6355 (N_6355,N_6143,N_6047);
xor U6356 (N_6356,N_6070,N_6200);
and U6357 (N_6357,N_6128,N_6228);
and U6358 (N_6358,N_6190,N_6191);
nor U6359 (N_6359,N_6077,N_6215);
nand U6360 (N_6360,N_6230,N_6049);
nor U6361 (N_6361,N_6059,N_6195);
nor U6362 (N_6362,N_6042,N_6147);
or U6363 (N_6363,N_6239,N_6210);
and U6364 (N_6364,N_6040,N_6113);
and U6365 (N_6365,N_6054,N_6172);
or U6366 (N_6366,N_6194,N_6148);
xnor U6367 (N_6367,N_6149,N_6130);
or U6368 (N_6368,N_6244,N_6185);
or U6369 (N_6369,N_6180,N_6053);
nand U6370 (N_6370,N_6159,N_6142);
or U6371 (N_6371,N_6154,N_6189);
nor U6372 (N_6372,N_6133,N_6212);
xnor U6373 (N_6373,N_6007,N_6119);
nand U6374 (N_6374,N_6160,N_6102);
and U6375 (N_6375,N_6033,N_6115);
or U6376 (N_6376,N_6113,N_6017);
or U6377 (N_6377,N_6182,N_6232);
and U6378 (N_6378,N_6036,N_6167);
and U6379 (N_6379,N_6059,N_6057);
nor U6380 (N_6380,N_6209,N_6197);
nand U6381 (N_6381,N_6065,N_6092);
nand U6382 (N_6382,N_6177,N_6082);
nor U6383 (N_6383,N_6049,N_6098);
nand U6384 (N_6384,N_6190,N_6043);
or U6385 (N_6385,N_6219,N_6095);
nand U6386 (N_6386,N_6240,N_6121);
nor U6387 (N_6387,N_6145,N_6188);
or U6388 (N_6388,N_6012,N_6149);
xor U6389 (N_6389,N_6245,N_6133);
or U6390 (N_6390,N_6056,N_6207);
nor U6391 (N_6391,N_6068,N_6173);
xor U6392 (N_6392,N_6107,N_6212);
and U6393 (N_6393,N_6018,N_6152);
nand U6394 (N_6394,N_6046,N_6180);
xnor U6395 (N_6395,N_6224,N_6027);
or U6396 (N_6396,N_6218,N_6166);
xnor U6397 (N_6397,N_6026,N_6003);
nor U6398 (N_6398,N_6139,N_6001);
nor U6399 (N_6399,N_6202,N_6221);
and U6400 (N_6400,N_6040,N_6191);
nor U6401 (N_6401,N_6123,N_6145);
and U6402 (N_6402,N_6232,N_6242);
or U6403 (N_6403,N_6054,N_6094);
nor U6404 (N_6404,N_6040,N_6041);
or U6405 (N_6405,N_6096,N_6168);
xnor U6406 (N_6406,N_6242,N_6033);
xor U6407 (N_6407,N_6212,N_6033);
xnor U6408 (N_6408,N_6185,N_6235);
xor U6409 (N_6409,N_6054,N_6177);
nor U6410 (N_6410,N_6091,N_6073);
nand U6411 (N_6411,N_6086,N_6062);
xor U6412 (N_6412,N_6232,N_6233);
or U6413 (N_6413,N_6121,N_6041);
or U6414 (N_6414,N_6147,N_6211);
nand U6415 (N_6415,N_6021,N_6065);
or U6416 (N_6416,N_6058,N_6039);
nand U6417 (N_6417,N_6063,N_6188);
nor U6418 (N_6418,N_6202,N_6084);
or U6419 (N_6419,N_6089,N_6173);
or U6420 (N_6420,N_6069,N_6191);
nor U6421 (N_6421,N_6143,N_6126);
xnor U6422 (N_6422,N_6031,N_6179);
nor U6423 (N_6423,N_6210,N_6248);
or U6424 (N_6424,N_6059,N_6110);
nor U6425 (N_6425,N_6055,N_6058);
nor U6426 (N_6426,N_6163,N_6202);
nand U6427 (N_6427,N_6116,N_6193);
xor U6428 (N_6428,N_6207,N_6249);
xor U6429 (N_6429,N_6133,N_6087);
nand U6430 (N_6430,N_6172,N_6140);
or U6431 (N_6431,N_6003,N_6066);
xnor U6432 (N_6432,N_6053,N_6198);
nand U6433 (N_6433,N_6059,N_6074);
nor U6434 (N_6434,N_6132,N_6081);
and U6435 (N_6435,N_6162,N_6183);
nand U6436 (N_6436,N_6139,N_6215);
xor U6437 (N_6437,N_6020,N_6080);
or U6438 (N_6438,N_6190,N_6161);
and U6439 (N_6439,N_6036,N_6053);
and U6440 (N_6440,N_6149,N_6242);
and U6441 (N_6441,N_6218,N_6156);
xor U6442 (N_6442,N_6063,N_6019);
nand U6443 (N_6443,N_6175,N_6017);
xor U6444 (N_6444,N_6231,N_6007);
nor U6445 (N_6445,N_6183,N_6095);
or U6446 (N_6446,N_6108,N_6110);
xnor U6447 (N_6447,N_6249,N_6042);
nand U6448 (N_6448,N_6237,N_6189);
nand U6449 (N_6449,N_6070,N_6056);
nor U6450 (N_6450,N_6185,N_6076);
nor U6451 (N_6451,N_6051,N_6068);
xnor U6452 (N_6452,N_6202,N_6152);
nand U6453 (N_6453,N_6180,N_6230);
nor U6454 (N_6454,N_6137,N_6220);
or U6455 (N_6455,N_6121,N_6016);
and U6456 (N_6456,N_6193,N_6133);
nand U6457 (N_6457,N_6235,N_6008);
nor U6458 (N_6458,N_6084,N_6134);
nor U6459 (N_6459,N_6194,N_6239);
and U6460 (N_6460,N_6141,N_6008);
nand U6461 (N_6461,N_6106,N_6135);
nor U6462 (N_6462,N_6008,N_6009);
and U6463 (N_6463,N_6133,N_6207);
or U6464 (N_6464,N_6037,N_6142);
and U6465 (N_6465,N_6244,N_6081);
and U6466 (N_6466,N_6245,N_6159);
nand U6467 (N_6467,N_6211,N_6186);
and U6468 (N_6468,N_6204,N_6217);
and U6469 (N_6469,N_6149,N_6015);
or U6470 (N_6470,N_6068,N_6165);
nor U6471 (N_6471,N_6143,N_6170);
and U6472 (N_6472,N_6228,N_6094);
and U6473 (N_6473,N_6246,N_6124);
nor U6474 (N_6474,N_6166,N_6228);
nand U6475 (N_6475,N_6144,N_6060);
or U6476 (N_6476,N_6180,N_6179);
nor U6477 (N_6477,N_6219,N_6168);
or U6478 (N_6478,N_6069,N_6168);
or U6479 (N_6479,N_6149,N_6005);
or U6480 (N_6480,N_6126,N_6075);
xnor U6481 (N_6481,N_6035,N_6017);
xnor U6482 (N_6482,N_6244,N_6111);
and U6483 (N_6483,N_6199,N_6216);
or U6484 (N_6484,N_6085,N_6146);
nor U6485 (N_6485,N_6212,N_6215);
xor U6486 (N_6486,N_6136,N_6070);
xnor U6487 (N_6487,N_6206,N_6196);
nand U6488 (N_6488,N_6055,N_6151);
and U6489 (N_6489,N_6046,N_6071);
nand U6490 (N_6490,N_6241,N_6073);
and U6491 (N_6491,N_6214,N_6201);
nor U6492 (N_6492,N_6204,N_6007);
and U6493 (N_6493,N_6192,N_6198);
nand U6494 (N_6494,N_6049,N_6032);
nor U6495 (N_6495,N_6113,N_6213);
nand U6496 (N_6496,N_6090,N_6106);
nor U6497 (N_6497,N_6023,N_6153);
xnor U6498 (N_6498,N_6050,N_6170);
nor U6499 (N_6499,N_6117,N_6001);
and U6500 (N_6500,N_6461,N_6251);
and U6501 (N_6501,N_6481,N_6367);
or U6502 (N_6502,N_6480,N_6337);
nor U6503 (N_6503,N_6347,N_6274);
and U6504 (N_6504,N_6250,N_6391);
xnor U6505 (N_6505,N_6382,N_6387);
and U6506 (N_6506,N_6309,N_6463);
or U6507 (N_6507,N_6334,N_6497);
nor U6508 (N_6508,N_6401,N_6331);
nor U6509 (N_6509,N_6451,N_6482);
and U6510 (N_6510,N_6293,N_6386);
or U6511 (N_6511,N_6414,N_6345);
or U6512 (N_6512,N_6487,N_6404);
and U6513 (N_6513,N_6266,N_6490);
xnor U6514 (N_6514,N_6454,N_6422);
nor U6515 (N_6515,N_6333,N_6253);
or U6516 (N_6516,N_6476,N_6311);
nor U6517 (N_6517,N_6296,N_6312);
or U6518 (N_6518,N_6393,N_6326);
xnor U6519 (N_6519,N_6332,N_6300);
nor U6520 (N_6520,N_6283,N_6433);
nand U6521 (N_6521,N_6389,N_6379);
nor U6522 (N_6522,N_6486,N_6460);
nand U6523 (N_6523,N_6264,N_6488);
and U6524 (N_6524,N_6479,N_6324);
nor U6525 (N_6525,N_6438,N_6304);
and U6526 (N_6526,N_6349,N_6259);
xor U6527 (N_6527,N_6318,N_6350);
xnor U6528 (N_6528,N_6355,N_6362);
nand U6529 (N_6529,N_6286,N_6342);
nor U6530 (N_6530,N_6385,N_6258);
nand U6531 (N_6531,N_6319,N_6361);
nand U6532 (N_6532,N_6366,N_6429);
nor U6533 (N_6533,N_6493,N_6364);
nor U6534 (N_6534,N_6257,N_6336);
or U6535 (N_6535,N_6464,N_6335);
nand U6536 (N_6536,N_6357,N_6498);
nand U6537 (N_6537,N_6327,N_6427);
nand U6538 (N_6538,N_6343,N_6275);
xor U6539 (N_6539,N_6282,N_6330);
or U6540 (N_6540,N_6428,N_6453);
nand U6541 (N_6541,N_6290,N_6262);
nor U6542 (N_6542,N_6284,N_6484);
and U6543 (N_6543,N_6425,N_6383);
nand U6544 (N_6544,N_6470,N_6279);
nand U6545 (N_6545,N_6281,N_6462);
and U6546 (N_6546,N_6491,N_6458);
or U6547 (N_6547,N_6365,N_6270);
or U6548 (N_6548,N_6411,N_6372);
or U6549 (N_6549,N_6340,N_6378);
or U6550 (N_6550,N_6255,N_6437);
or U6551 (N_6551,N_6374,N_6289);
nand U6552 (N_6552,N_6419,N_6441);
and U6553 (N_6553,N_6417,N_6354);
nor U6554 (N_6554,N_6444,N_6373);
and U6555 (N_6555,N_6265,N_6384);
or U6556 (N_6556,N_6256,N_6492);
nor U6557 (N_6557,N_6267,N_6371);
nor U6558 (N_6558,N_6377,N_6420);
xor U6559 (N_6559,N_6313,N_6459);
and U6560 (N_6560,N_6489,N_6329);
xnor U6561 (N_6561,N_6341,N_6485);
nand U6562 (N_6562,N_6431,N_6421);
nor U6563 (N_6563,N_6370,N_6358);
nand U6564 (N_6564,N_6439,N_6306);
nor U6565 (N_6565,N_6430,N_6314);
and U6566 (N_6566,N_6352,N_6452);
nand U6567 (N_6567,N_6418,N_6495);
and U6568 (N_6568,N_6472,N_6325);
or U6569 (N_6569,N_6400,N_6317);
xor U6570 (N_6570,N_6397,N_6473);
or U6571 (N_6571,N_6443,N_6388);
nor U6572 (N_6572,N_6432,N_6465);
and U6573 (N_6573,N_6447,N_6285);
or U6574 (N_6574,N_6315,N_6483);
nand U6575 (N_6575,N_6353,N_6398);
or U6576 (N_6576,N_6322,N_6294);
nand U6577 (N_6577,N_6269,N_6346);
or U6578 (N_6578,N_6298,N_6413);
xor U6579 (N_6579,N_6399,N_6310);
nand U6580 (N_6580,N_6499,N_6456);
nor U6581 (N_6581,N_6405,N_6457);
nor U6582 (N_6582,N_6424,N_6351);
nand U6583 (N_6583,N_6273,N_6477);
nor U6584 (N_6584,N_6423,N_6408);
or U6585 (N_6585,N_6426,N_6446);
or U6586 (N_6586,N_6407,N_6392);
and U6587 (N_6587,N_6308,N_6471);
nor U6588 (N_6588,N_6302,N_6445);
or U6589 (N_6589,N_6261,N_6301);
and U6590 (N_6590,N_6403,N_6396);
nand U6591 (N_6591,N_6494,N_6415);
nand U6592 (N_6592,N_6369,N_6468);
and U6593 (N_6593,N_6475,N_6381);
or U6594 (N_6594,N_6394,N_6410);
nand U6595 (N_6595,N_6328,N_6272);
nand U6596 (N_6596,N_6416,N_6467);
xnor U6597 (N_6597,N_6316,N_6321);
nand U6598 (N_6598,N_6278,N_6436);
nor U6599 (N_6599,N_6360,N_6406);
xnor U6600 (N_6600,N_6380,N_6252);
nand U6601 (N_6601,N_6478,N_6295);
and U6602 (N_6602,N_6450,N_6466);
or U6603 (N_6603,N_6375,N_6276);
nor U6604 (N_6604,N_6287,N_6288);
nand U6605 (N_6605,N_6292,N_6268);
xor U6606 (N_6606,N_6469,N_6435);
xnor U6607 (N_6607,N_6344,N_6320);
nand U6608 (N_6608,N_6440,N_6434);
and U6609 (N_6609,N_6356,N_6448);
xor U6610 (N_6610,N_6359,N_6280);
nand U6611 (N_6611,N_6395,N_6254);
nand U6612 (N_6612,N_6449,N_6363);
or U6613 (N_6613,N_6305,N_6303);
nand U6614 (N_6614,N_6307,N_6291);
xnor U6615 (N_6615,N_6376,N_6277);
or U6616 (N_6616,N_6455,N_6474);
xor U6617 (N_6617,N_6390,N_6402);
or U6618 (N_6618,N_6271,N_6339);
nor U6619 (N_6619,N_6299,N_6323);
nand U6620 (N_6620,N_6442,N_6368);
xnor U6621 (N_6621,N_6260,N_6338);
nand U6622 (N_6622,N_6297,N_6263);
nor U6623 (N_6623,N_6496,N_6348);
nor U6624 (N_6624,N_6412,N_6409);
xnor U6625 (N_6625,N_6341,N_6417);
and U6626 (N_6626,N_6286,N_6463);
or U6627 (N_6627,N_6305,N_6414);
nor U6628 (N_6628,N_6385,N_6266);
nor U6629 (N_6629,N_6451,N_6416);
nor U6630 (N_6630,N_6458,N_6316);
xnor U6631 (N_6631,N_6488,N_6405);
nor U6632 (N_6632,N_6466,N_6460);
nand U6633 (N_6633,N_6389,N_6424);
and U6634 (N_6634,N_6285,N_6331);
nand U6635 (N_6635,N_6299,N_6385);
nor U6636 (N_6636,N_6461,N_6495);
or U6637 (N_6637,N_6298,N_6435);
nor U6638 (N_6638,N_6392,N_6482);
xnor U6639 (N_6639,N_6405,N_6494);
nor U6640 (N_6640,N_6323,N_6434);
and U6641 (N_6641,N_6429,N_6343);
nand U6642 (N_6642,N_6346,N_6477);
nor U6643 (N_6643,N_6387,N_6447);
or U6644 (N_6644,N_6330,N_6252);
and U6645 (N_6645,N_6296,N_6289);
and U6646 (N_6646,N_6272,N_6464);
xor U6647 (N_6647,N_6441,N_6272);
and U6648 (N_6648,N_6406,N_6350);
or U6649 (N_6649,N_6421,N_6432);
xnor U6650 (N_6650,N_6274,N_6444);
xor U6651 (N_6651,N_6304,N_6454);
nand U6652 (N_6652,N_6294,N_6391);
xor U6653 (N_6653,N_6357,N_6418);
nand U6654 (N_6654,N_6464,N_6491);
nor U6655 (N_6655,N_6265,N_6420);
nand U6656 (N_6656,N_6469,N_6433);
nand U6657 (N_6657,N_6287,N_6420);
and U6658 (N_6658,N_6442,N_6285);
or U6659 (N_6659,N_6436,N_6402);
nor U6660 (N_6660,N_6277,N_6463);
xnor U6661 (N_6661,N_6358,N_6498);
nand U6662 (N_6662,N_6407,N_6368);
nor U6663 (N_6663,N_6328,N_6295);
xor U6664 (N_6664,N_6428,N_6451);
nor U6665 (N_6665,N_6349,N_6303);
and U6666 (N_6666,N_6338,N_6371);
nor U6667 (N_6667,N_6448,N_6499);
nor U6668 (N_6668,N_6443,N_6305);
or U6669 (N_6669,N_6291,N_6415);
and U6670 (N_6670,N_6491,N_6362);
nand U6671 (N_6671,N_6483,N_6463);
or U6672 (N_6672,N_6281,N_6371);
nor U6673 (N_6673,N_6454,N_6328);
and U6674 (N_6674,N_6478,N_6492);
and U6675 (N_6675,N_6434,N_6378);
xnor U6676 (N_6676,N_6292,N_6397);
nand U6677 (N_6677,N_6271,N_6319);
nand U6678 (N_6678,N_6465,N_6403);
nor U6679 (N_6679,N_6484,N_6330);
xor U6680 (N_6680,N_6274,N_6328);
nor U6681 (N_6681,N_6257,N_6278);
xnor U6682 (N_6682,N_6449,N_6473);
nand U6683 (N_6683,N_6401,N_6434);
nand U6684 (N_6684,N_6281,N_6294);
or U6685 (N_6685,N_6366,N_6465);
or U6686 (N_6686,N_6398,N_6487);
nand U6687 (N_6687,N_6475,N_6463);
xnor U6688 (N_6688,N_6297,N_6451);
xnor U6689 (N_6689,N_6497,N_6265);
and U6690 (N_6690,N_6274,N_6470);
or U6691 (N_6691,N_6360,N_6453);
and U6692 (N_6692,N_6253,N_6450);
xnor U6693 (N_6693,N_6291,N_6350);
and U6694 (N_6694,N_6401,N_6373);
nor U6695 (N_6695,N_6323,N_6268);
xnor U6696 (N_6696,N_6432,N_6401);
nand U6697 (N_6697,N_6424,N_6381);
nand U6698 (N_6698,N_6476,N_6346);
and U6699 (N_6699,N_6378,N_6306);
and U6700 (N_6700,N_6343,N_6302);
or U6701 (N_6701,N_6373,N_6316);
nand U6702 (N_6702,N_6449,N_6277);
or U6703 (N_6703,N_6428,N_6319);
nand U6704 (N_6704,N_6353,N_6347);
and U6705 (N_6705,N_6310,N_6409);
and U6706 (N_6706,N_6441,N_6444);
or U6707 (N_6707,N_6408,N_6281);
and U6708 (N_6708,N_6409,N_6260);
xnor U6709 (N_6709,N_6483,N_6393);
nand U6710 (N_6710,N_6373,N_6344);
nand U6711 (N_6711,N_6435,N_6287);
nor U6712 (N_6712,N_6387,N_6260);
nor U6713 (N_6713,N_6394,N_6291);
or U6714 (N_6714,N_6284,N_6398);
or U6715 (N_6715,N_6370,N_6431);
xor U6716 (N_6716,N_6306,N_6362);
and U6717 (N_6717,N_6250,N_6336);
nor U6718 (N_6718,N_6257,N_6342);
or U6719 (N_6719,N_6445,N_6444);
nor U6720 (N_6720,N_6281,N_6480);
xnor U6721 (N_6721,N_6324,N_6349);
xnor U6722 (N_6722,N_6366,N_6398);
nand U6723 (N_6723,N_6425,N_6366);
xor U6724 (N_6724,N_6489,N_6286);
xnor U6725 (N_6725,N_6419,N_6285);
xor U6726 (N_6726,N_6329,N_6412);
nor U6727 (N_6727,N_6439,N_6326);
nor U6728 (N_6728,N_6360,N_6457);
xnor U6729 (N_6729,N_6296,N_6299);
or U6730 (N_6730,N_6417,N_6289);
nor U6731 (N_6731,N_6408,N_6418);
and U6732 (N_6732,N_6293,N_6356);
nand U6733 (N_6733,N_6441,N_6482);
xnor U6734 (N_6734,N_6414,N_6420);
or U6735 (N_6735,N_6492,N_6439);
xnor U6736 (N_6736,N_6449,N_6491);
xnor U6737 (N_6737,N_6426,N_6429);
nor U6738 (N_6738,N_6371,N_6277);
xnor U6739 (N_6739,N_6322,N_6347);
xnor U6740 (N_6740,N_6345,N_6474);
nand U6741 (N_6741,N_6326,N_6305);
or U6742 (N_6742,N_6365,N_6386);
or U6743 (N_6743,N_6266,N_6360);
xnor U6744 (N_6744,N_6418,N_6323);
and U6745 (N_6745,N_6443,N_6454);
or U6746 (N_6746,N_6371,N_6291);
xor U6747 (N_6747,N_6365,N_6284);
nor U6748 (N_6748,N_6366,N_6381);
nor U6749 (N_6749,N_6311,N_6430);
and U6750 (N_6750,N_6582,N_6731);
or U6751 (N_6751,N_6739,N_6612);
or U6752 (N_6752,N_6562,N_6618);
nand U6753 (N_6753,N_6743,N_6736);
xor U6754 (N_6754,N_6501,N_6570);
or U6755 (N_6755,N_6599,N_6584);
nand U6756 (N_6756,N_6628,N_6633);
or U6757 (N_6757,N_6635,N_6523);
nand U6758 (N_6758,N_6590,N_6676);
nand U6759 (N_6759,N_6504,N_6620);
nand U6760 (N_6760,N_6573,N_6694);
nor U6761 (N_6761,N_6686,N_6639);
or U6762 (N_6762,N_6643,N_6671);
and U6763 (N_6763,N_6687,N_6653);
nor U6764 (N_6764,N_6536,N_6601);
xor U6765 (N_6765,N_6563,N_6626);
nor U6766 (N_6766,N_6502,N_6566);
xor U6767 (N_6767,N_6511,N_6551);
nor U6768 (N_6768,N_6592,N_6726);
nor U6769 (N_6769,N_6638,N_6652);
xor U6770 (N_6770,N_6544,N_6651);
or U6771 (N_6771,N_6611,N_6575);
xnor U6772 (N_6772,N_6520,N_6623);
or U6773 (N_6773,N_6666,N_6644);
or U6774 (N_6774,N_6588,N_6675);
xor U6775 (N_6775,N_6578,N_6598);
xnor U6776 (N_6776,N_6569,N_6669);
and U6777 (N_6777,N_6722,N_6553);
nand U6778 (N_6778,N_6572,N_6703);
nand U6779 (N_6779,N_6614,N_6568);
and U6780 (N_6780,N_6581,N_6593);
xor U6781 (N_6781,N_6571,N_6595);
and U6782 (N_6782,N_6717,N_6738);
xor U6783 (N_6783,N_6547,N_6522);
nand U6784 (N_6784,N_6613,N_6604);
nor U6785 (N_6785,N_6622,N_6559);
nor U6786 (N_6786,N_6558,N_6552);
and U6787 (N_6787,N_6707,N_6541);
and U6788 (N_6788,N_6503,N_6561);
xor U6789 (N_6789,N_6539,N_6712);
xnor U6790 (N_6790,N_6554,N_6577);
nand U6791 (N_6791,N_6699,N_6602);
and U6792 (N_6792,N_6673,N_6690);
nand U6793 (N_6793,N_6709,N_6677);
nor U6794 (N_6794,N_6745,N_6720);
nand U6795 (N_6795,N_6519,N_6701);
xnor U6796 (N_6796,N_6596,N_6579);
xor U6797 (N_6797,N_6667,N_6531);
nor U6798 (N_6798,N_6659,N_6663);
nand U6799 (N_6799,N_6637,N_6733);
nor U6800 (N_6800,N_6550,N_6606);
or U6801 (N_6801,N_6640,N_6656);
xnor U6802 (N_6802,N_6728,N_6528);
nand U6803 (N_6803,N_6715,N_6615);
and U6804 (N_6804,N_6713,N_6710);
or U6805 (N_6805,N_6723,N_6548);
nor U6806 (N_6806,N_6688,N_6509);
and U6807 (N_6807,N_6603,N_6744);
nand U6808 (N_6808,N_6698,N_6674);
nor U6809 (N_6809,N_6514,N_6672);
and U6810 (N_6810,N_6660,N_6537);
nand U6811 (N_6811,N_6585,N_6532);
nand U6812 (N_6812,N_6591,N_6624);
or U6813 (N_6813,N_6734,N_6682);
or U6814 (N_6814,N_6729,N_6625);
xnor U6815 (N_6815,N_6714,N_6629);
xnor U6816 (N_6816,N_6608,N_6505);
xor U6817 (N_6817,N_6708,N_6556);
nand U6818 (N_6818,N_6557,N_6691);
nor U6819 (N_6819,N_6576,N_6605);
nand U6820 (N_6820,N_6580,N_6518);
and U6821 (N_6821,N_6670,N_6678);
or U6822 (N_6822,N_6740,N_6661);
and U6823 (N_6823,N_6508,N_6727);
and U6824 (N_6824,N_6646,N_6711);
nor U6825 (N_6825,N_6645,N_6648);
or U6826 (N_6826,N_6642,N_6683);
nor U6827 (N_6827,N_6538,N_6695);
nor U6828 (N_6828,N_6679,N_6724);
nand U6829 (N_6829,N_6540,N_6632);
and U6830 (N_6830,N_6607,N_6680);
nand U6831 (N_6831,N_6650,N_6630);
nand U6832 (N_6832,N_6693,N_6649);
or U6833 (N_6833,N_6685,N_6749);
and U6834 (N_6834,N_6658,N_6515);
nor U6835 (N_6835,N_6735,N_6589);
xnor U6836 (N_6836,N_6730,N_6610);
xor U6837 (N_6837,N_6741,N_6600);
and U6838 (N_6838,N_6597,N_6594);
or U6839 (N_6839,N_6721,N_6748);
nor U6840 (N_6840,N_6725,N_6631);
xor U6841 (N_6841,N_6574,N_6587);
xnor U6842 (N_6842,N_6747,N_6533);
xnor U6843 (N_6843,N_6526,N_6534);
nand U6844 (N_6844,N_6527,N_6655);
nor U6845 (N_6845,N_6718,N_6545);
nand U6846 (N_6846,N_6542,N_6662);
or U6847 (N_6847,N_6529,N_6516);
nor U6848 (N_6848,N_6716,N_6546);
nand U6849 (N_6849,N_6510,N_6530);
xor U6850 (N_6850,N_6692,N_6647);
or U6851 (N_6851,N_6567,N_6746);
nand U6852 (N_6852,N_6617,N_6549);
and U6853 (N_6853,N_6697,N_6535);
xnor U6854 (N_6854,N_6513,N_6621);
or U6855 (N_6855,N_6521,N_6586);
nor U6856 (N_6856,N_6689,N_6619);
and U6857 (N_6857,N_6668,N_6719);
and U6858 (N_6858,N_6512,N_6634);
and U6859 (N_6859,N_6742,N_6565);
or U6860 (N_6860,N_6500,N_6627);
nand U6861 (N_6861,N_6665,N_6507);
nand U6862 (N_6862,N_6506,N_6702);
and U6863 (N_6863,N_6704,N_6583);
or U6864 (N_6864,N_6705,N_6616);
xor U6865 (N_6865,N_6641,N_6555);
or U6866 (N_6866,N_6525,N_6560);
nor U6867 (N_6867,N_6636,N_6684);
nor U6868 (N_6868,N_6564,N_6543);
or U6869 (N_6869,N_6681,N_6524);
xnor U6870 (N_6870,N_6737,N_6654);
or U6871 (N_6871,N_6664,N_6706);
xor U6872 (N_6872,N_6609,N_6517);
and U6873 (N_6873,N_6732,N_6657);
or U6874 (N_6874,N_6700,N_6696);
nand U6875 (N_6875,N_6727,N_6546);
xor U6876 (N_6876,N_6740,N_6621);
or U6877 (N_6877,N_6587,N_6643);
xor U6878 (N_6878,N_6616,N_6656);
or U6879 (N_6879,N_6661,N_6692);
xnor U6880 (N_6880,N_6670,N_6684);
and U6881 (N_6881,N_6704,N_6616);
xnor U6882 (N_6882,N_6684,N_6679);
nand U6883 (N_6883,N_6563,N_6651);
nor U6884 (N_6884,N_6615,N_6700);
or U6885 (N_6885,N_6569,N_6737);
nor U6886 (N_6886,N_6691,N_6588);
xnor U6887 (N_6887,N_6647,N_6680);
and U6888 (N_6888,N_6602,N_6689);
and U6889 (N_6889,N_6719,N_6653);
or U6890 (N_6890,N_6670,N_6527);
nand U6891 (N_6891,N_6582,N_6600);
or U6892 (N_6892,N_6747,N_6569);
nand U6893 (N_6893,N_6524,N_6697);
or U6894 (N_6894,N_6665,N_6560);
xnor U6895 (N_6895,N_6736,N_6707);
nor U6896 (N_6896,N_6558,N_6726);
and U6897 (N_6897,N_6555,N_6724);
or U6898 (N_6898,N_6723,N_6559);
nand U6899 (N_6899,N_6723,N_6530);
nand U6900 (N_6900,N_6704,N_6690);
nand U6901 (N_6901,N_6575,N_6522);
nand U6902 (N_6902,N_6700,N_6721);
or U6903 (N_6903,N_6700,N_6740);
xor U6904 (N_6904,N_6643,N_6695);
or U6905 (N_6905,N_6735,N_6693);
or U6906 (N_6906,N_6524,N_6511);
xor U6907 (N_6907,N_6705,N_6711);
or U6908 (N_6908,N_6717,N_6612);
or U6909 (N_6909,N_6516,N_6557);
nor U6910 (N_6910,N_6539,N_6557);
nand U6911 (N_6911,N_6646,N_6707);
nand U6912 (N_6912,N_6585,N_6741);
xor U6913 (N_6913,N_6604,N_6639);
nand U6914 (N_6914,N_6559,N_6573);
and U6915 (N_6915,N_6659,N_6706);
nor U6916 (N_6916,N_6616,N_6523);
xnor U6917 (N_6917,N_6702,N_6611);
nor U6918 (N_6918,N_6536,N_6590);
nor U6919 (N_6919,N_6599,N_6666);
nor U6920 (N_6920,N_6595,N_6736);
nand U6921 (N_6921,N_6617,N_6657);
xor U6922 (N_6922,N_6505,N_6729);
or U6923 (N_6923,N_6556,N_6639);
xnor U6924 (N_6924,N_6573,N_6625);
or U6925 (N_6925,N_6688,N_6660);
or U6926 (N_6926,N_6570,N_6571);
and U6927 (N_6927,N_6596,N_6583);
nor U6928 (N_6928,N_6541,N_6620);
xnor U6929 (N_6929,N_6542,N_6546);
or U6930 (N_6930,N_6502,N_6527);
nor U6931 (N_6931,N_6535,N_6713);
xor U6932 (N_6932,N_6676,N_6666);
nand U6933 (N_6933,N_6746,N_6503);
or U6934 (N_6934,N_6666,N_6706);
xor U6935 (N_6935,N_6747,N_6706);
or U6936 (N_6936,N_6538,N_6519);
xnor U6937 (N_6937,N_6714,N_6684);
and U6938 (N_6938,N_6609,N_6561);
and U6939 (N_6939,N_6508,N_6579);
and U6940 (N_6940,N_6694,N_6611);
nand U6941 (N_6941,N_6638,N_6579);
nand U6942 (N_6942,N_6645,N_6669);
nor U6943 (N_6943,N_6686,N_6533);
nor U6944 (N_6944,N_6739,N_6566);
xnor U6945 (N_6945,N_6653,N_6701);
and U6946 (N_6946,N_6556,N_6574);
xor U6947 (N_6947,N_6564,N_6607);
nand U6948 (N_6948,N_6655,N_6658);
or U6949 (N_6949,N_6594,N_6701);
or U6950 (N_6950,N_6537,N_6693);
xnor U6951 (N_6951,N_6700,N_6542);
nor U6952 (N_6952,N_6512,N_6591);
nand U6953 (N_6953,N_6533,N_6728);
xnor U6954 (N_6954,N_6556,N_6526);
nand U6955 (N_6955,N_6536,N_6630);
nor U6956 (N_6956,N_6654,N_6694);
xnor U6957 (N_6957,N_6560,N_6603);
nor U6958 (N_6958,N_6595,N_6650);
nand U6959 (N_6959,N_6579,N_6716);
xor U6960 (N_6960,N_6709,N_6614);
or U6961 (N_6961,N_6683,N_6556);
and U6962 (N_6962,N_6747,N_6710);
nor U6963 (N_6963,N_6627,N_6564);
xnor U6964 (N_6964,N_6629,N_6627);
nand U6965 (N_6965,N_6706,N_6675);
or U6966 (N_6966,N_6608,N_6516);
or U6967 (N_6967,N_6594,N_6643);
xor U6968 (N_6968,N_6623,N_6638);
xor U6969 (N_6969,N_6565,N_6529);
xor U6970 (N_6970,N_6699,N_6545);
nor U6971 (N_6971,N_6651,N_6652);
or U6972 (N_6972,N_6641,N_6747);
xnor U6973 (N_6973,N_6578,N_6706);
or U6974 (N_6974,N_6531,N_6555);
nor U6975 (N_6975,N_6527,N_6614);
xor U6976 (N_6976,N_6533,N_6709);
xnor U6977 (N_6977,N_6722,N_6611);
nor U6978 (N_6978,N_6529,N_6572);
nor U6979 (N_6979,N_6674,N_6731);
nand U6980 (N_6980,N_6647,N_6704);
nor U6981 (N_6981,N_6603,N_6665);
xnor U6982 (N_6982,N_6530,N_6532);
xnor U6983 (N_6983,N_6569,N_6612);
and U6984 (N_6984,N_6522,N_6549);
xor U6985 (N_6985,N_6627,N_6702);
xnor U6986 (N_6986,N_6600,N_6713);
nor U6987 (N_6987,N_6634,N_6680);
nand U6988 (N_6988,N_6587,N_6604);
nand U6989 (N_6989,N_6735,N_6606);
nor U6990 (N_6990,N_6642,N_6584);
nand U6991 (N_6991,N_6735,N_6643);
nand U6992 (N_6992,N_6539,N_6697);
and U6993 (N_6993,N_6624,N_6527);
and U6994 (N_6994,N_6737,N_6552);
nor U6995 (N_6995,N_6696,N_6746);
xor U6996 (N_6996,N_6569,N_6512);
nand U6997 (N_6997,N_6515,N_6716);
nor U6998 (N_6998,N_6563,N_6559);
nor U6999 (N_6999,N_6594,N_6705);
or U7000 (N_7000,N_6874,N_6965);
nor U7001 (N_7001,N_6920,N_6772);
xor U7002 (N_7002,N_6891,N_6930);
or U7003 (N_7003,N_6881,N_6958);
nand U7004 (N_7004,N_6990,N_6901);
nor U7005 (N_7005,N_6919,N_6816);
nand U7006 (N_7006,N_6935,N_6973);
nor U7007 (N_7007,N_6789,N_6976);
xnor U7008 (N_7008,N_6883,N_6906);
and U7009 (N_7009,N_6803,N_6888);
and U7010 (N_7010,N_6807,N_6941);
xnor U7011 (N_7011,N_6926,N_6963);
xor U7012 (N_7012,N_6895,N_6945);
nand U7013 (N_7013,N_6970,N_6819);
nand U7014 (N_7014,N_6866,N_6854);
nand U7015 (N_7015,N_6972,N_6840);
and U7016 (N_7016,N_6837,N_6823);
or U7017 (N_7017,N_6839,N_6953);
nor U7018 (N_7018,N_6910,N_6811);
xor U7019 (N_7019,N_6944,N_6787);
nand U7020 (N_7020,N_6946,N_6836);
nor U7021 (N_7021,N_6890,N_6774);
nand U7022 (N_7022,N_6848,N_6959);
nand U7023 (N_7023,N_6957,N_6824);
xnor U7024 (N_7024,N_6898,N_6755);
nand U7025 (N_7025,N_6809,N_6821);
nand U7026 (N_7026,N_6869,N_6877);
nor U7027 (N_7027,N_6750,N_6842);
xnor U7028 (N_7028,N_6796,N_6951);
or U7029 (N_7029,N_6799,N_6915);
or U7030 (N_7030,N_6790,N_6776);
nand U7031 (N_7031,N_6762,N_6923);
and U7032 (N_7032,N_6868,N_6937);
xnor U7033 (N_7033,N_6832,N_6993);
nor U7034 (N_7034,N_6801,N_6812);
and U7035 (N_7035,N_6966,N_6781);
nand U7036 (N_7036,N_6934,N_6834);
or U7037 (N_7037,N_6880,N_6788);
xnor U7038 (N_7038,N_6810,N_6798);
nand U7039 (N_7039,N_6967,N_6897);
nand U7040 (N_7040,N_6765,N_6994);
and U7041 (N_7041,N_6975,N_6918);
nor U7042 (N_7042,N_6763,N_6899);
or U7043 (N_7043,N_6845,N_6850);
nor U7044 (N_7044,N_6981,N_6949);
xor U7045 (N_7045,N_6887,N_6940);
nor U7046 (N_7046,N_6753,N_6863);
or U7047 (N_7047,N_6871,N_6779);
or U7048 (N_7048,N_6838,N_6955);
nor U7049 (N_7049,N_6815,N_6828);
or U7050 (N_7050,N_6766,N_6768);
nand U7051 (N_7051,N_6835,N_6875);
nor U7052 (N_7052,N_6947,N_6998);
nor U7053 (N_7053,N_6956,N_6980);
and U7054 (N_7054,N_6974,N_6933);
and U7055 (N_7055,N_6969,N_6769);
or U7056 (N_7056,N_6861,N_6870);
or U7057 (N_7057,N_6770,N_6939);
xor U7058 (N_7058,N_6797,N_6917);
xor U7059 (N_7059,N_6800,N_6985);
nor U7060 (N_7060,N_6978,N_6813);
nand U7061 (N_7061,N_6808,N_6833);
and U7062 (N_7062,N_6761,N_6979);
and U7063 (N_7063,N_6997,N_6847);
nand U7064 (N_7064,N_6829,N_6983);
or U7065 (N_7065,N_6977,N_6855);
and U7066 (N_7066,N_6794,N_6950);
and U7067 (N_7067,N_6989,N_6878);
or U7068 (N_7068,N_6818,N_6912);
nor U7069 (N_7069,N_6921,N_6773);
or U7070 (N_7070,N_6860,N_6913);
nor U7071 (N_7071,N_6795,N_6756);
or U7072 (N_7072,N_6914,N_6864);
nand U7073 (N_7073,N_6907,N_6889);
xor U7074 (N_7074,N_6771,N_6791);
nor U7075 (N_7075,N_6767,N_6885);
and U7076 (N_7076,N_6784,N_6826);
nand U7077 (N_7077,N_6938,N_6841);
nor U7078 (N_7078,N_6844,N_6830);
or U7079 (N_7079,N_6852,N_6988);
nor U7080 (N_7080,N_6778,N_6805);
nor U7081 (N_7081,N_6896,N_6825);
xor U7082 (N_7082,N_6793,N_6879);
nand U7083 (N_7083,N_6886,N_6857);
xnor U7084 (N_7084,N_6777,N_6752);
nand U7085 (N_7085,N_6827,N_6751);
nor U7086 (N_7086,N_6804,N_6991);
or U7087 (N_7087,N_6892,N_6822);
xnor U7088 (N_7088,N_6786,N_6916);
or U7089 (N_7089,N_6849,N_6900);
xnor U7090 (N_7090,N_6814,N_6758);
and U7091 (N_7091,N_6846,N_6936);
xnor U7092 (N_7092,N_6882,N_6931);
and U7093 (N_7093,N_6908,N_6865);
nor U7094 (N_7094,N_6909,N_6922);
nand U7095 (N_7095,N_6952,N_6785);
nand U7096 (N_7096,N_6929,N_6843);
and U7097 (N_7097,N_6902,N_6853);
nor U7098 (N_7098,N_6876,N_6859);
xnor U7099 (N_7099,N_6894,N_6925);
xnor U7100 (N_7100,N_6851,N_6995);
or U7101 (N_7101,N_6954,N_6831);
or U7102 (N_7102,N_6802,N_6928);
xnor U7103 (N_7103,N_6754,N_6856);
and U7104 (N_7104,N_6872,N_6905);
nor U7105 (N_7105,N_6971,N_6862);
nor U7106 (N_7106,N_6932,N_6911);
xor U7107 (N_7107,N_6943,N_6792);
or U7108 (N_7108,N_6817,N_6964);
nor U7109 (N_7109,N_6858,N_6782);
or U7110 (N_7110,N_6948,N_6992);
and U7111 (N_7111,N_6968,N_6759);
xnor U7112 (N_7112,N_6757,N_6996);
xnor U7113 (N_7113,N_6760,N_6806);
or U7114 (N_7114,N_6960,N_6927);
and U7115 (N_7115,N_6764,N_6904);
and U7116 (N_7116,N_6942,N_6984);
nor U7117 (N_7117,N_6903,N_6884);
xnor U7118 (N_7118,N_6867,N_6962);
and U7119 (N_7119,N_6820,N_6873);
nor U7120 (N_7120,N_6775,N_6986);
xnor U7121 (N_7121,N_6783,N_6961);
xor U7122 (N_7122,N_6982,N_6999);
nor U7123 (N_7123,N_6780,N_6924);
nand U7124 (N_7124,N_6893,N_6987);
or U7125 (N_7125,N_6964,N_6786);
nand U7126 (N_7126,N_6985,N_6838);
and U7127 (N_7127,N_6772,N_6871);
or U7128 (N_7128,N_6950,N_6771);
nand U7129 (N_7129,N_6886,N_6998);
and U7130 (N_7130,N_6789,N_6995);
and U7131 (N_7131,N_6902,N_6936);
or U7132 (N_7132,N_6951,N_6808);
nor U7133 (N_7133,N_6904,N_6865);
nor U7134 (N_7134,N_6842,N_6962);
or U7135 (N_7135,N_6861,N_6914);
nor U7136 (N_7136,N_6938,N_6909);
or U7137 (N_7137,N_6796,N_6903);
nand U7138 (N_7138,N_6783,N_6918);
nand U7139 (N_7139,N_6926,N_6828);
and U7140 (N_7140,N_6977,N_6952);
nor U7141 (N_7141,N_6841,N_6847);
or U7142 (N_7142,N_6788,N_6947);
or U7143 (N_7143,N_6807,N_6875);
nor U7144 (N_7144,N_6912,N_6881);
or U7145 (N_7145,N_6979,N_6952);
or U7146 (N_7146,N_6750,N_6988);
or U7147 (N_7147,N_6919,N_6793);
nand U7148 (N_7148,N_6913,N_6816);
nor U7149 (N_7149,N_6769,N_6986);
nor U7150 (N_7150,N_6762,N_6968);
xnor U7151 (N_7151,N_6994,N_6938);
xnor U7152 (N_7152,N_6982,N_6778);
nor U7153 (N_7153,N_6846,N_6981);
nor U7154 (N_7154,N_6792,N_6967);
or U7155 (N_7155,N_6897,N_6762);
or U7156 (N_7156,N_6828,N_6968);
nand U7157 (N_7157,N_6988,N_6992);
nor U7158 (N_7158,N_6954,N_6795);
and U7159 (N_7159,N_6903,N_6974);
nand U7160 (N_7160,N_6945,N_6862);
and U7161 (N_7161,N_6940,N_6916);
xnor U7162 (N_7162,N_6903,N_6917);
or U7163 (N_7163,N_6799,N_6809);
and U7164 (N_7164,N_6841,N_6817);
nor U7165 (N_7165,N_6878,N_6827);
or U7166 (N_7166,N_6843,N_6812);
nor U7167 (N_7167,N_6832,N_6763);
xor U7168 (N_7168,N_6960,N_6956);
or U7169 (N_7169,N_6756,N_6933);
and U7170 (N_7170,N_6915,N_6954);
or U7171 (N_7171,N_6860,N_6983);
or U7172 (N_7172,N_6948,N_6906);
xor U7173 (N_7173,N_6900,N_6919);
xor U7174 (N_7174,N_6921,N_6864);
and U7175 (N_7175,N_6774,N_6985);
and U7176 (N_7176,N_6958,N_6930);
or U7177 (N_7177,N_6967,N_6815);
or U7178 (N_7178,N_6813,N_6900);
nor U7179 (N_7179,N_6848,N_6943);
nand U7180 (N_7180,N_6970,N_6865);
or U7181 (N_7181,N_6899,N_6787);
and U7182 (N_7182,N_6796,N_6917);
or U7183 (N_7183,N_6849,N_6885);
or U7184 (N_7184,N_6868,N_6947);
nor U7185 (N_7185,N_6854,N_6898);
or U7186 (N_7186,N_6813,N_6868);
or U7187 (N_7187,N_6976,N_6823);
nor U7188 (N_7188,N_6818,N_6913);
nand U7189 (N_7189,N_6807,N_6957);
or U7190 (N_7190,N_6778,N_6852);
or U7191 (N_7191,N_6856,N_6875);
or U7192 (N_7192,N_6985,N_6781);
nand U7193 (N_7193,N_6850,N_6763);
and U7194 (N_7194,N_6956,N_6967);
and U7195 (N_7195,N_6756,N_6878);
nand U7196 (N_7196,N_6808,N_6819);
or U7197 (N_7197,N_6989,N_6948);
nand U7198 (N_7198,N_6908,N_6795);
xnor U7199 (N_7199,N_6867,N_6892);
or U7200 (N_7200,N_6845,N_6900);
nor U7201 (N_7201,N_6988,N_6760);
nor U7202 (N_7202,N_6953,N_6908);
xor U7203 (N_7203,N_6986,N_6925);
nor U7204 (N_7204,N_6925,N_6777);
or U7205 (N_7205,N_6982,N_6996);
and U7206 (N_7206,N_6988,N_6967);
xnor U7207 (N_7207,N_6891,N_6802);
nand U7208 (N_7208,N_6830,N_6914);
nand U7209 (N_7209,N_6934,N_6905);
nor U7210 (N_7210,N_6938,N_6908);
and U7211 (N_7211,N_6946,N_6757);
xnor U7212 (N_7212,N_6914,N_6788);
nor U7213 (N_7213,N_6845,N_6783);
nand U7214 (N_7214,N_6985,N_6983);
nor U7215 (N_7215,N_6830,N_6943);
nor U7216 (N_7216,N_6969,N_6838);
or U7217 (N_7217,N_6876,N_6959);
xor U7218 (N_7218,N_6937,N_6972);
nor U7219 (N_7219,N_6888,N_6786);
and U7220 (N_7220,N_6996,N_6792);
and U7221 (N_7221,N_6913,N_6970);
and U7222 (N_7222,N_6873,N_6897);
and U7223 (N_7223,N_6912,N_6838);
or U7224 (N_7224,N_6872,N_6871);
nor U7225 (N_7225,N_6808,N_6927);
xnor U7226 (N_7226,N_6780,N_6776);
and U7227 (N_7227,N_6837,N_6785);
or U7228 (N_7228,N_6835,N_6806);
nor U7229 (N_7229,N_6852,N_6810);
nand U7230 (N_7230,N_6923,N_6969);
and U7231 (N_7231,N_6817,N_6786);
nand U7232 (N_7232,N_6978,N_6802);
and U7233 (N_7233,N_6866,N_6799);
or U7234 (N_7234,N_6860,N_6890);
nor U7235 (N_7235,N_6958,N_6774);
xnor U7236 (N_7236,N_6767,N_6855);
nand U7237 (N_7237,N_6863,N_6833);
xnor U7238 (N_7238,N_6764,N_6961);
nor U7239 (N_7239,N_6792,N_6782);
nand U7240 (N_7240,N_6952,N_6770);
or U7241 (N_7241,N_6892,N_6906);
and U7242 (N_7242,N_6863,N_6898);
nand U7243 (N_7243,N_6908,N_6830);
nand U7244 (N_7244,N_6858,N_6875);
nor U7245 (N_7245,N_6844,N_6800);
and U7246 (N_7246,N_6989,N_6891);
xnor U7247 (N_7247,N_6770,N_6822);
xnor U7248 (N_7248,N_6811,N_6849);
xor U7249 (N_7249,N_6991,N_6889);
and U7250 (N_7250,N_7101,N_7096);
and U7251 (N_7251,N_7159,N_7081);
and U7252 (N_7252,N_7059,N_7086);
xor U7253 (N_7253,N_7236,N_7129);
nand U7254 (N_7254,N_7131,N_7139);
and U7255 (N_7255,N_7188,N_7073);
or U7256 (N_7256,N_7220,N_7109);
or U7257 (N_7257,N_7009,N_7244);
and U7258 (N_7258,N_7022,N_7173);
or U7259 (N_7259,N_7155,N_7175);
or U7260 (N_7260,N_7238,N_7209);
nand U7261 (N_7261,N_7006,N_7003);
xor U7262 (N_7262,N_7061,N_7121);
and U7263 (N_7263,N_7053,N_7118);
nor U7264 (N_7264,N_7093,N_7213);
nand U7265 (N_7265,N_7152,N_7240);
or U7266 (N_7266,N_7034,N_7145);
xnor U7267 (N_7267,N_7084,N_7027);
and U7268 (N_7268,N_7067,N_7219);
and U7269 (N_7269,N_7141,N_7114);
xnor U7270 (N_7270,N_7024,N_7187);
xor U7271 (N_7271,N_7211,N_7001);
nor U7272 (N_7272,N_7134,N_7070);
and U7273 (N_7273,N_7106,N_7176);
xnor U7274 (N_7274,N_7202,N_7013);
nor U7275 (N_7275,N_7012,N_7161);
nor U7276 (N_7276,N_7181,N_7063);
and U7277 (N_7277,N_7221,N_7092);
nor U7278 (N_7278,N_7052,N_7196);
or U7279 (N_7279,N_7172,N_7107);
and U7280 (N_7280,N_7130,N_7124);
xnor U7281 (N_7281,N_7040,N_7080);
nor U7282 (N_7282,N_7117,N_7064);
and U7283 (N_7283,N_7206,N_7039);
xnor U7284 (N_7284,N_7033,N_7110);
and U7285 (N_7285,N_7185,N_7143);
and U7286 (N_7286,N_7076,N_7190);
and U7287 (N_7287,N_7068,N_7007);
and U7288 (N_7288,N_7150,N_7045);
and U7289 (N_7289,N_7232,N_7186);
nand U7290 (N_7290,N_7099,N_7023);
xnor U7291 (N_7291,N_7234,N_7217);
nor U7292 (N_7292,N_7163,N_7104);
and U7293 (N_7293,N_7123,N_7216);
or U7294 (N_7294,N_7242,N_7182);
and U7295 (N_7295,N_7204,N_7002);
xnor U7296 (N_7296,N_7165,N_7066);
xor U7297 (N_7297,N_7168,N_7017);
xnor U7298 (N_7298,N_7199,N_7077);
nor U7299 (N_7299,N_7088,N_7029);
xor U7300 (N_7300,N_7249,N_7091);
nand U7301 (N_7301,N_7230,N_7098);
or U7302 (N_7302,N_7158,N_7178);
nor U7303 (N_7303,N_7011,N_7193);
xor U7304 (N_7304,N_7097,N_7184);
xor U7305 (N_7305,N_7103,N_7014);
and U7306 (N_7306,N_7164,N_7038);
nand U7307 (N_7307,N_7025,N_7237);
xor U7308 (N_7308,N_7146,N_7179);
or U7309 (N_7309,N_7136,N_7051);
nand U7310 (N_7310,N_7015,N_7054);
nor U7311 (N_7311,N_7169,N_7245);
and U7312 (N_7312,N_7167,N_7020);
nand U7313 (N_7313,N_7198,N_7194);
and U7314 (N_7314,N_7069,N_7154);
nand U7315 (N_7315,N_7083,N_7225);
or U7316 (N_7316,N_7082,N_7010);
and U7317 (N_7317,N_7115,N_7043);
nor U7318 (N_7318,N_7127,N_7113);
or U7319 (N_7319,N_7205,N_7037);
and U7320 (N_7320,N_7112,N_7031);
or U7321 (N_7321,N_7227,N_7032);
and U7322 (N_7322,N_7180,N_7128);
and U7323 (N_7323,N_7089,N_7100);
nor U7324 (N_7324,N_7079,N_7018);
xor U7325 (N_7325,N_7019,N_7229);
and U7326 (N_7326,N_7215,N_7049);
or U7327 (N_7327,N_7075,N_7153);
nand U7328 (N_7328,N_7036,N_7016);
and U7329 (N_7329,N_7138,N_7197);
or U7330 (N_7330,N_7135,N_7223);
nand U7331 (N_7331,N_7246,N_7005);
xnor U7332 (N_7332,N_7162,N_7021);
nand U7333 (N_7333,N_7208,N_7026);
or U7334 (N_7334,N_7057,N_7239);
xnor U7335 (N_7335,N_7000,N_7247);
nand U7336 (N_7336,N_7105,N_7071);
xnor U7337 (N_7337,N_7008,N_7200);
nor U7338 (N_7338,N_7144,N_7210);
nand U7339 (N_7339,N_7111,N_7214);
and U7340 (N_7340,N_7055,N_7191);
nor U7341 (N_7341,N_7235,N_7241);
or U7342 (N_7342,N_7094,N_7041);
or U7343 (N_7343,N_7030,N_7177);
or U7344 (N_7344,N_7132,N_7189);
or U7345 (N_7345,N_7090,N_7047);
nor U7346 (N_7346,N_7060,N_7170);
nor U7347 (N_7347,N_7222,N_7133);
and U7348 (N_7348,N_7224,N_7072);
and U7349 (N_7349,N_7226,N_7156);
nor U7350 (N_7350,N_7166,N_7116);
nand U7351 (N_7351,N_7085,N_7119);
nor U7352 (N_7352,N_7120,N_7192);
nor U7353 (N_7353,N_7160,N_7035);
nand U7354 (N_7354,N_7228,N_7207);
and U7355 (N_7355,N_7147,N_7126);
and U7356 (N_7356,N_7050,N_7195);
xor U7357 (N_7357,N_7183,N_7108);
and U7358 (N_7358,N_7046,N_7044);
or U7359 (N_7359,N_7142,N_7004);
and U7360 (N_7360,N_7065,N_7148);
nand U7361 (N_7361,N_7137,N_7095);
xnor U7362 (N_7362,N_7231,N_7203);
nor U7363 (N_7363,N_7074,N_7218);
and U7364 (N_7364,N_7028,N_7056);
nor U7365 (N_7365,N_7171,N_7122);
nand U7366 (N_7366,N_7243,N_7125);
or U7367 (N_7367,N_7042,N_7151);
nand U7368 (N_7368,N_7102,N_7157);
nor U7369 (N_7369,N_7140,N_7087);
and U7370 (N_7370,N_7078,N_7048);
nor U7371 (N_7371,N_7233,N_7058);
nor U7372 (N_7372,N_7212,N_7201);
nand U7373 (N_7373,N_7174,N_7149);
or U7374 (N_7374,N_7062,N_7248);
nor U7375 (N_7375,N_7131,N_7082);
nor U7376 (N_7376,N_7003,N_7134);
xnor U7377 (N_7377,N_7143,N_7151);
nor U7378 (N_7378,N_7244,N_7072);
nor U7379 (N_7379,N_7026,N_7113);
and U7380 (N_7380,N_7161,N_7183);
nand U7381 (N_7381,N_7019,N_7052);
xnor U7382 (N_7382,N_7186,N_7226);
nand U7383 (N_7383,N_7142,N_7139);
and U7384 (N_7384,N_7068,N_7187);
and U7385 (N_7385,N_7218,N_7182);
nor U7386 (N_7386,N_7215,N_7077);
nand U7387 (N_7387,N_7186,N_7140);
and U7388 (N_7388,N_7001,N_7090);
and U7389 (N_7389,N_7060,N_7112);
or U7390 (N_7390,N_7053,N_7069);
nor U7391 (N_7391,N_7226,N_7070);
and U7392 (N_7392,N_7113,N_7231);
nor U7393 (N_7393,N_7182,N_7159);
nand U7394 (N_7394,N_7205,N_7197);
and U7395 (N_7395,N_7004,N_7139);
nor U7396 (N_7396,N_7020,N_7105);
or U7397 (N_7397,N_7167,N_7010);
or U7398 (N_7398,N_7049,N_7003);
and U7399 (N_7399,N_7194,N_7021);
nor U7400 (N_7400,N_7198,N_7083);
and U7401 (N_7401,N_7141,N_7057);
or U7402 (N_7402,N_7091,N_7038);
nand U7403 (N_7403,N_7188,N_7048);
nand U7404 (N_7404,N_7191,N_7003);
nand U7405 (N_7405,N_7080,N_7113);
xor U7406 (N_7406,N_7051,N_7249);
or U7407 (N_7407,N_7234,N_7049);
xnor U7408 (N_7408,N_7126,N_7014);
and U7409 (N_7409,N_7022,N_7243);
and U7410 (N_7410,N_7160,N_7100);
or U7411 (N_7411,N_7026,N_7144);
nor U7412 (N_7412,N_7197,N_7245);
nand U7413 (N_7413,N_7164,N_7174);
nand U7414 (N_7414,N_7027,N_7068);
and U7415 (N_7415,N_7026,N_7219);
and U7416 (N_7416,N_7041,N_7055);
or U7417 (N_7417,N_7150,N_7026);
and U7418 (N_7418,N_7101,N_7161);
nand U7419 (N_7419,N_7036,N_7014);
or U7420 (N_7420,N_7145,N_7041);
nor U7421 (N_7421,N_7232,N_7175);
xor U7422 (N_7422,N_7162,N_7172);
or U7423 (N_7423,N_7078,N_7088);
or U7424 (N_7424,N_7152,N_7120);
or U7425 (N_7425,N_7137,N_7089);
nand U7426 (N_7426,N_7192,N_7018);
or U7427 (N_7427,N_7127,N_7167);
xor U7428 (N_7428,N_7093,N_7050);
nand U7429 (N_7429,N_7172,N_7085);
nor U7430 (N_7430,N_7144,N_7216);
nand U7431 (N_7431,N_7207,N_7231);
xor U7432 (N_7432,N_7093,N_7242);
nor U7433 (N_7433,N_7107,N_7085);
nor U7434 (N_7434,N_7038,N_7092);
nor U7435 (N_7435,N_7057,N_7026);
nor U7436 (N_7436,N_7228,N_7136);
or U7437 (N_7437,N_7107,N_7123);
nor U7438 (N_7438,N_7097,N_7104);
nand U7439 (N_7439,N_7052,N_7080);
or U7440 (N_7440,N_7033,N_7238);
nand U7441 (N_7441,N_7164,N_7036);
xor U7442 (N_7442,N_7229,N_7081);
and U7443 (N_7443,N_7020,N_7104);
and U7444 (N_7444,N_7007,N_7030);
or U7445 (N_7445,N_7172,N_7071);
and U7446 (N_7446,N_7124,N_7018);
and U7447 (N_7447,N_7170,N_7126);
nand U7448 (N_7448,N_7086,N_7168);
and U7449 (N_7449,N_7097,N_7231);
nand U7450 (N_7450,N_7083,N_7184);
nor U7451 (N_7451,N_7135,N_7249);
nand U7452 (N_7452,N_7009,N_7063);
or U7453 (N_7453,N_7181,N_7169);
xor U7454 (N_7454,N_7063,N_7081);
xor U7455 (N_7455,N_7112,N_7236);
nor U7456 (N_7456,N_7166,N_7018);
nand U7457 (N_7457,N_7033,N_7246);
nor U7458 (N_7458,N_7190,N_7231);
xnor U7459 (N_7459,N_7022,N_7105);
or U7460 (N_7460,N_7214,N_7168);
and U7461 (N_7461,N_7155,N_7187);
nand U7462 (N_7462,N_7165,N_7071);
nor U7463 (N_7463,N_7193,N_7033);
nor U7464 (N_7464,N_7119,N_7034);
nand U7465 (N_7465,N_7071,N_7027);
or U7466 (N_7466,N_7097,N_7090);
xor U7467 (N_7467,N_7019,N_7191);
nand U7468 (N_7468,N_7153,N_7204);
and U7469 (N_7469,N_7230,N_7190);
or U7470 (N_7470,N_7079,N_7214);
and U7471 (N_7471,N_7043,N_7247);
or U7472 (N_7472,N_7081,N_7211);
and U7473 (N_7473,N_7216,N_7006);
nand U7474 (N_7474,N_7144,N_7135);
and U7475 (N_7475,N_7067,N_7043);
nor U7476 (N_7476,N_7100,N_7073);
nor U7477 (N_7477,N_7154,N_7029);
or U7478 (N_7478,N_7090,N_7108);
nand U7479 (N_7479,N_7175,N_7219);
xnor U7480 (N_7480,N_7091,N_7005);
nand U7481 (N_7481,N_7176,N_7008);
nor U7482 (N_7482,N_7129,N_7075);
nand U7483 (N_7483,N_7058,N_7090);
xnor U7484 (N_7484,N_7015,N_7249);
nand U7485 (N_7485,N_7083,N_7079);
or U7486 (N_7486,N_7046,N_7173);
nor U7487 (N_7487,N_7008,N_7132);
xor U7488 (N_7488,N_7080,N_7165);
nand U7489 (N_7489,N_7119,N_7025);
xnor U7490 (N_7490,N_7212,N_7106);
or U7491 (N_7491,N_7054,N_7028);
nor U7492 (N_7492,N_7174,N_7218);
nand U7493 (N_7493,N_7083,N_7065);
xnor U7494 (N_7494,N_7205,N_7041);
nor U7495 (N_7495,N_7096,N_7012);
xnor U7496 (N_7496,N_7058,N_7046);
or U7497 (N_7497,N_7167,N_7021);
or U7498 (N_7498,N_7066,N_7009);
and U7499 (N_7499,N_7195,N_7225);
xnor U7500 (N_7500,N_7312,N_7291);
xnor U7501 (N_7501,N_7493,N_7424);
xor U7502 (N_7502,N_7304,N_7400);
nand U7503 (N_7503,N_7420,N_7298);
or U7504 (N_7504,N_7485,N_7314);
or U7505 (N_7505,N_7361,N_7473);
or U7506 (N_7506,N_7283,N_7385);
nand U7507 (N_7507,N_7296,N_7413);
or U7508 (N_7508,N_7459,N_7263);
and U7509 (N_7509,N_7490,N_7461);
and U7510 (N_7510,N_7332,N_7282);
nand U7511 (N_7511,N_7325,N_7345);
or U7512 (N_7512,N_7386,N_7257);
xnor U7513 (N_7513,N_7383,N_7266);
nand U7514 (N_7514,N_7430,N_7271);
or U7515 (N_7515,N_7301,N_7417);
nor U7516 (N_7516,N_7446,N_7317);
or U7517 (N_7517,N_7453,N_7255);
nand U7518 (N_7518,N_7487,N_7418);
xor U7519 (N_7519,N_7456,N_7324);
nand U7520 (N_7520,N_7256,N_7320);
xnor U7521 (N_7521,N_7449,N_7342);
nor U7522 (N_7522,N_7469,N_7399);
or U7523 (N_7523,N_7445,N_7346);
or U7524 (N_7524,N_7462,N_7463);
xor U7525 (N_7525,N_7276,N_7484);
xor U7526 (N_7526,N_7497,N_7349);
nand U7527 (N_7527,N_7269,N_7443);
nor U7528 (N_7528,N_7372,N_7362);
nand U7529 (N_7529,N_7378,N_7458);
or U7530 (N_7530,N_7308,N_7406);
and U7531 (N_7531,N_7409,N_7394);
xor U7532 (N_7532,N_7405,N_7471);
xnor U7533 (N_7533,N_7297,N_7495);
nand U7534 (N_7534,N_7415,N_7439);
or U7535 (N_7535,N_7371,N_7474);
nor U7536 (N_7536,N_7337,N_7441);
nor U7537 (N_7537,N_7381,N_7486);
xnor U7538 (N_7538,N_7335,N_7273);
nor U7539 (N_7539,N_7410,N_7328);
nor U7540 (N_7540,N_7290,N_7481);
nand U7541 (N_7541,N_7464,N_7307);
nor U7542 (N_7542,N_7465,N_7295);
or U7543 (N_7543,N_7470,N_7375);
nand U7544 (N_7544,N_7368,N_7272);
nor U7545 (N_7545,N_7259,N_7480);
nor U7546 (N_7546,N_7275,N_7476);
or U7547 (N_7547,N_7452,N_7403);
xnor U7548 (N_7548,N_7251,N_7329);
xnor U7549 (N_7549,N_7348,N_7280);
nand U7550 (N_7550,N_7398,N_7444);
xor U7551 (N_7551,N_7357,N_7448);
xnor U7552 (N_7552,N_7302,N_7350);
or U7553 (N_7553,N_7306,N_7478);
or U7554 (N_7554,N_7412,N_7419);
xnor U7555 (N_7555,N_7310,N_7451);
nand U7556 (N_7556,N_7387,N_7366);
or U7557 (N_7557,N_7479,N_7364);
and U7558 (N_7558,N_7427,N_7323);
and U7559 (N_7559,N_7391,N_7351);
nor U7560 (N_7560,N_7299,N_7475);
and U7561 (N_7561,N_7414,N_7311);
or U7562 (N_7562,N_7294,N_7267);
or U7563 (N_7563,N_7395,N_7293);
xor U7564 (N_7564,N_7286,N_7354);
or U7565 (N_7565,N_7494,N_7392);
nand U7566 (N_7566,N_7369,N_7260);
xnor U7567 (N_7567,N_7384,N_7355);
xor U7568 (N_7568,N_7379,N_7258);
nand U7569 (N_7569,N_7488,N_7316);
nor U7570 (N_7570,N_7315,N_7416);
xnor U7571 (N_7571,N_7421,N_7352);
and U7572 (N_7572,N_7277,N_7343);
or U7573 (N_7573,N_7397,N_7376);
xor U7574 (N_7574,N_7434,N_7404);
and U7575 (N_7575,N_7360,N_7336);
xor U7576 (N_7576,N_7389,N_7455);
and U7577 (N_7577,N_7344,N_7450);
nor U7578 (N_7578,N_7285,N_7252);
and U7579 (N_7579,N_7460,N_7374);
and U7580 (N_7580,N_7279,N_7401);
xnor U7581 (N_7581,N_7367,N_7334);
nand U7582 (N_7582,N_7353,N_7442);
and U7583 (N_7583,N_7466,N_7402);
and U7584 (N_7584,N_7333,N_7327);
or U7585 (N_7585,N_7278,N_7382);
nand U7586 (N_7586,N_7318,N_7390);
nand U7587 (N_7587,N_7373,N_7338);
nor U7588 (N_7588,N_7491,N_7321);
xnor U7589 (N_7589,N_7408,N_7429);
xor U7590 (N_7590,N_7426,N_7423);
nand U7591 (N_7591,N_7341,N_7477);
nor U7592 (N_7592,N_7288,N_7436);
nor U7593 (N_7593,N_7437,N_7326);
nand U7594 (N_7594,N_7287,N_7281);
nand U7595 (N_7595,N_7447,N_7431);
nand U7596 (N_7596,N_7330,N_7322);
nor U7597 (N_7597,N_7356,N_7472);
or U7598 (N_7598,N_7340,N_7411);
nand U7599 (N_7599,N_7303,N_7440);
nor U7600 (N_7600,N_7268,N_7492);
nor U7601 (N_7601,N_7380,N_7454);
nand U7602 (N_7602,N_7300,N_7347);
nor U7603 (N_7603,N_7270,N_7262);
and U7604 (N_7604,N_7407,N_7396);
nand U7605 (N_7605,N_7428,N_7489);
nor U7606 (N_7606,N_7331,N_7483);
or U7607 (N_7607,N_7496,N_7435);
or U7608 (N_7608,N_7365,N_7363);
nor U7609 (N_7609,N_7359,N_7482);
and U7610 (N_7610,N_7289,N_7425);
or U7611 (N_7611,N_7370,N_7261);
and U7612 (N_7612,N_7264,N_7250);
nor U7613 (N_7613,N_7274,N_7422);
or U7614 (N_7614,N_7254,N_7319);
or U7615 (N_7615,N_7292,N_7432);
nand U7616 (N_7616,N_7265,N_7433);
and U7617 (N_7617,N_7468,N_7457);
or U7618 (N_7618,N_7284,N_7253);
or U7619 (N_7619,N_7377,N_7339);
nor U7620 (N_7620,N_7388,N_7499);
nand U7621 (N_7621,N_7438,N_7358);
nand U7622 (N_7622,N_7467,N_7305);
and U7623 (N_7623,N_7498,N_7313);
nor U7624 (N_7624,N_7309,N_7393);
nor U7625 (N_7625,N_7261,N_7473);
or U7626 (N_7626,N_7423,N_7416);
xor U7627 (N_7627,N_7311,N_7386);
or U7628 (N_7628,N_7367,N_7337);
and U7629 (N_7629,N_7453,N_7419);
nand U7630 (N_7630,N_7278,N_7424);
and U7631 (N_7631,N_7493,N_7418);
nand U7632 (N_7632,N_7268,N_7385);
and U7633 (N_7633,N_7450,N_7471);
nand U7634 (N_7634,N_7478,N_7447);
nand U7635 (N_7635,N_7402,N_7342);
xnor U7636 (N_7636,N_7312,N_7392);
or U7637 (N_7637,N_7354,N_7448);
xnor U7638 (N_7638,N_7310,N_7492);
or U7639 (N_7639,N_7306,N_7290);
and U7640 (N_7640,N_7360,N_7477);
nand U7641 (N_7641,N_7414,N_7295);
nor U7642 (N_7642,N_7262,N_7467);
nor U7643 (N_7643,N_7390,N_7301);
or U7644 (N_7644,N_7454,N_7357);
and U7645 (N_7645,N_7466,N_7454);
nor U7646 (N_7646,N_7354,N_7397);
nand U7647 (N_7647,N_7411,N_7488);
nor U7648 (N_7648,N_7334,N_7292);
and U7649 (N_7649,N_7407,N_7456);
xnor U7650 (N_7650,N_7391,N_7316);
nand U7651 (N_7651,N_7389,N_7362);
nor U7652 (N_7652,N_7367,N_7459);
or U7653 (N_7653,N_7353,N_7289);
xor U7654 (N_7654,N_7313,N_7359);
or U7655 (N_7655,N_7264,N_7432);
or U7656 (N_7656,N_7407,N_7370);
xor U7657 (N_7657,N_7472,N_7376);
xor U7658 (N_7658,N_7280,N_7474);
nand U7659 (N_7659,N_7315,N_7384);
nor U7660 (N_7660,N_7452,N_7289);
or U7661 (N_7661,N_7331,N_7372);
or U7662 (N_7662,N_7270,N_7385);
and U7663 (N_7663,N_7307,N_7387);
nand U7664 (N_7664,N_7461,N_7335);
and U7665 (N_7665,N_7269,N_7474);
nand U7666 (N_7666,N_7460,N_7469);
or U7667 (N_7667,N_7353,N_7459);
or U7668 (N_7668,N_7495,N_7388);
xnor U7669 (N_7669,N_7322,N_7273);
nand U7670 (N_7670,N_7339,N_7412);
or U7671 (N_7671,N_7329,N_7274);
nand U7672 (N_7672,N_7263,N_7250);
or U7673 (N_7673,N_7362,N_7410);
and U7674 (N_7674,N_7253,N_7394);
nand U7675 (N_7675,N_7416,N_7397);
xor U7676 (N_7676,N_7441,N_7275);
nor U7677 (N_7677,N_7480,N_7253);
nor U7678 (N_7678,N_7453,N_7498);
nor U7679 (N_7679,N_7271,N_7282);
xnor U7680 (N_7680,N_7282,N_7278);
or U7681 (N_7681,N_7277,N_7264);
nand U7682 (N_7682,N_7264,N_7283);
nand U7683 (N_7683,N_7481,N_7370);
nor U7684 (N_7684,N_7469,N_7358);
nand U7685 (N_7685,N_7402,N_7488);
nand U7686 (N_7686,N_7401,N_7290);
nor U7687 (N_7687,N_7370,N_7415);
nand U7688 (N_7688,N_7272,N_7313);
xnor U7689 (N_7689,N_7367,N_7300);
or U7690 (N_7690,N_7409,N_7318);
xnor U7691 (N_7691,N_7275,N_7331);
xor U7692 (N_7692,N_7484,N_7482);
and U7693 (N_7693,N_7395,N_7262);
nor U7694 (N_7694,N_7302,N_7367);
xor U7695 (N_7695,N_7281,N_7354);
nand U7696 (N_7696,N_7499,N_7489);
xnor U7697 (N_7697,N_7410,N_7493);
or U7698 (N_7698,N_7480,N_7417);
nor U7699 (N_7699,N_7485,N_7295);
and U7700 (N_7700,N_7299,N_7491);
nor U7701 (N_7701,N_7378,N_7455);
and U7702 (N_7702,N_7353,N_7356);
xor U7703 (N_7703,N_7479,N_7303);
nor U7704 (N_7704,N_7455,N_7261);
nand U7705 (N_7705,N_7395,N_7302);
nand U7706 (N_7706,N_7314,N_7460);
xor U7707 (N_7707,N_7423,N_7491);
nor U7708 (N_7708,N_7341,N_7451);
xnor U7709 (N_7709,N_7296,N_7291);
and U7710 (N_7710,N_7280,N_7412);
and U7711 (N_7711,N_7288,N_7348);
and U7712 (N_7712,N_7347,N_7470);
and U7713 (N_7713,N_7284,N_7305);
and U7714 (N_7714,N_7407,N_7348);
nor U7715 (N_7715,N_7363,N_7461);
or U7716 (N_7716,N_7338,N_7465);
xnor U7717 (N_7717,N_7472,N_7296);
nand U7718 (N_7718,N_7498,N_7440);
nor U7719 (N_7719,N_7478,N_7449);
xor U7720 (N_7720,N_7307,N_7324);
xnor U7721 (N_7721,N_7296,N_7339);
or U7722 (N_7722,N_7498,N_7450);
and U7723 (N_7723,N_7419,N_7452);
nor U7724 (N_7724,N_7397,N_7454);
or U7725 (N_7725,N_7360,N_7478);
and U7726 (N_7726,N_7278,N_7457);
nor U7727 (N_7727,N_7421,N_7395);
nand U7728 (N_7728,N_7269,N_7496);
xor U7729 (N_7729,N_7403,N_7395);
and U7730 (N_7730,N_7367,N_7429);
nand U7731 (N_7731,N_7286,N_7361);
nor U7732 (N_7732,N_7326,N_7417);
xor U7733 (N_7733,N_7324,N_7349);
nand U7734 (N_7734,N_7280,N_7311);
and U7735 (N_7735,N_7416,N_7259);
nor U7736 (N_7736,N_7316,N_7492);
or U7737 (N_7737,N_7481,N_7444);
and U7738 (N_7738,N_7412,N_7458);
nor U7739 (N_7739,N_7390,N_7469);
or U7740 (N_7740,N_7427,N_7261);
or U7741 (N_7741,N_7465,N_7303);
or U7742 (N_7742,N_7274,N_7428);
nor U7743 (N_7743,N_7295,N_7301);
xor U7744 (N_7744,N_7480,N_7415);
or U7745 (N_7745,N_7462,N_7492);
xor U7746 (N_7746,N_7401,N_7275);
nor U7747 (N_7747,N_7416,N_7479);
or U7748 (N_7748,N_7286,N_7384);
or U7749 (N_7749,N_7360,N_7355);
nand U7750 (N_7750,N_7551,N_7698);
or U7751 (N_7751,N_7574,N_7713);
and U7752 (N_7752,N_7717,N_7659);
nor U7753 (N_7753,N_7516,N_7631);
or U7754 (N_7754,N_7668,N_7609);
or U7755 (N_7755,N_7563,N_7593);
nand U7756 (N_7756,N_7532,N_7710);
xor U7757 (N_7757,N_7673,N_7730);
and U7758 (N_7758,N_7575,N_7579);
nand U7759 (N_7759,N_7583,N_7678);
nor U7760 (N_7760,N_7513,N_7716);
xor U7761 (N_7761,N_7680,N_7610);
xor U7762 (N_7762,N_7547,N_7682);
nand U7763 (N_7763,N_7633,N_7656);
or U7764 (N_7764,N_7719,N_7694);
or U7765 (N_7765,N_7515,N_7505);
nor U7766 (N_7766,N_7524,N_7604);
or U7767 (N_7767,N_7556,N_7708);
nand U7768 (N_7768,N_7540,N_7500);
nand U7769 (N_7769,N_7661,N_7614);
xnor U7770 (N_7770,N_7569,N_7714);
nor U7771 (N_7771,N_7667,N_7570);
nand U7772 (N_7772,N_7620,N_7543);
xnor U7773 (N_7773,N_7587,N_7725);
nand U7774 (N_7774,N_7744,N_7566);
nand U7775 (N_7775,N_7677,N_7534);
and U7776 (N_7776,N_7572,N_7553);
nor U7777 (N_7777,N_7526,N_7726);
nand U7778 (N_7778,N_7695,N_7520);
nand U7779 (N_7779,N_7650,N_7697);
and U7780 (N_7780,N_7729,N_7724);
and U7781 (N_7781,N_7709,N_7648);
or U7782 (N_7782,N_7501,N_7676);
nor U7783 (N_7783,N_7595,N_7644);
nand U7784 (N_7784,N_7687,N_7723);
nor U7785 (N_7785,N_7601,N_7514);
or U7786 (N_7786,N_7696,N_7635);
and U7787 (N_7787,N_7689,N_7720);
or U7788 (N_7788,N_7508,N_7584);
xor U7789 (N_7789,N_7746,N_7712);
nor U7790 (N_7790,N_7627,N_7586);
and U7791 (N_7791,N_7679,N_7623);
xor U7792 (N_7792,N_7519,N_7550);
nand U7793 (N_7793,N_7743,N_7552);
nand U7794 (N_7794,N_7632,N_7548);
nor U7795 (N_7795,N_7615,N_7647);
nand U7796 (N_7796,N_7518,N_7649);
nor U7797 (N_7797,N_7666,N_7701);
nand U7798 (N_7798,N_7596,N_7704);
nor U7799 (N_7799,N_7739,N_7603);
xor U7800 (N_7800,N_7608,N_7654);
or U7801 (N_7801,N_7703,N_7693);
xnor U7802 (N_7802,N_7617,N_7692);
nand U7803 (N_7803,N_7747,N_7699);
xor U7804 (N_7804,N_7564,N_7736);
or U7805 (N_7805,N_7576,N_7545);
xnor U7806 (N_7806,N_7517,N_7625);
xnor U7807 (N_7807,N_7523,N_7504);
nand U7808 (N_7808,N_7585,N_7681);
or U7809 (N_7809,N_7662,N_7683);
xnor U7810 (N_7810,N_7742,N_7549);
or U7811 (N_7811,N_7542,N_7525);
or U7812 (N_7812,N_7581,N_7640);
nor U7813 (N_7813,N_7503,N_7691);
xnor U7814 (N_7814,N_7559,N_7598);
and U7815 (N_7815,N_7672,N_7506);
nor U7816 (N_7816,N_7619,N_7658);
nor U7817 (N_7817,N_7705,N_7621);
or U7818 (N_7818,N_7521,N_7684);
nor U7819 (N_7819,N_7711,N_7641);
or U7820 (N_7820,N_7533,N_7544);
or U7821 (N_7821,N_7655,N_7657);
and U7822 (N_7822,N_7613,N_7688);
nand U7823 (N_7823,N_7599,N_7628);
nand U7824 (N_7824,N_7580,N_7616);
nor U7825 (N_7825,N_7745,N_7642);
or U7826 (N_7826,N_7646,N_7728);
and U7827 (N_7827,N_7606,N_7541);
and U7828 (N_7828,N_7589,N_7733);
nor U7829 (N_7829,N_7555,N_7722);
nand U7830 (N_7830,N_7671,N_7735);
xor U7831 (N_7831,N_7536,N_7567);
nand U7832 (N_7832,N_7590,N_7578);
and U7833 (N_7833,N_7748,N_7690);
xor U7834 (N_7834,N_7571,N_7702);
or U7835 (N_7835,N_7664,N_7630);
and U7836 (N_7836,N_7718,N_7731);
nand U7837 (N_7837,N_7600,N_7502);
nor U7838 (N_7838,N_7741,N_7531);
xnor U7839 (N_7839,N_7685,N_7629);
or U7840 (N_7840,N_7597,N_7740);
nor U7841 (N_7841,N_7528,N_7535);
nand U7842 (N_7842,N_7622,N_7602);
nor U7843 (N_7843,N_7573,N_7611);
nor U7844 (N_7844,N_7727,N_7592);
nor U7845 (N_7845,N_7588,N_7607);
xnor U7846 (N_7846,N_7510,N_7558);
or U7847 (N_7847,N_7554,N_7591);
nor U7848 (N_7848,N_7660,N_7669);
xnor U7849 (N_7849,N_7707,N_7734);
xor U7850 (N_7850,N_7537,N_7686);
and U7851 (N_7851,N_7624,N_7560);
and U7852 (N_7852,N_7653,N_7568);
nor U7853 (N_7853,N_7651,N_7507);
and U7854 (N_7854,N_7652,N_7738);
or U7855 (N_7855,N_7582,N_7638);
nor U7856 (N_7856,N_7732,N_7715);
nor U7857 (N_7857,N_7645,N_7529);
nand U7858 (N_7858,N_7665,N_7737);
and U7859 (N_7859,N_7509,N_7561);
xor U7860 (N_7860,N_7618,N_7721);
xor U7861 (N_7861,N_7605,N_7670);
or U7862 (N_7862,N_7706,N_7749);
nor U7863 (N_7863,N_7634,N_7557);
or U7864 (N_7864,N_7522,N_7594);
xor U7865 (N_7865,N_7643,N_7562);
and U7866 (N_7866,N_7675,N_7538);
nand U7867 (N_7867,N_7512,N_7636);
and U7868 (N_7868,N_7674,N_7565);
xor U7869 (N_7869,N_7612,N_7546);
and U7870 (N_7870,N_7626,N_7663);
nor U7871 (N_7871,N_7577,N_7700);
nand U7872 (N_7872,N_7539,N_7527);
nand U7873 (N_7873,N_7511,N_7637);
nand U7874 (N_7874,N_7639,N_7530);
or U7875 (N_7875,N_7744,N_7710);
nand U7876 (N_7876,N_7579,N_7554);
or U7877 (N_7877,N_7520,N_7681);
nor U7878 (N_7878,N_7502,N_7525);
nand U7879 (N_7879,N_7740,N_7560);
and U7880 (N_7880,N_7648,N_7723);
and U7881 (N_7881,N_7640,N_7717);
and U7882 (N_7882,N_7730,N_7572);
or U7883 (N_7883,N_7714,N_7566);
xnor U7884 (N_7884,N_7513,N_7594);
nor U7885 (N_7885,N_7679,N_7660);
nand U7886 (N_7886,N_7560,N_7554);
or U7887 (N_7887,N_7629,N_7718);
nor U7888 (N_7888,N_7580,N_7558);
and U7889 (N_7889,N_7519,N_7674);
xor U7890 (N_7890,N_7646,N_7528);
xnor U7891 (N_7891,N_7519,N_7561);
xnor U7892 (N_7892,N_7692,N_7696);
nand U7893 (N_7893,N_7600,N_7733);
xor U7894 (N_7894,N_7736,N_7657);
and U7895 (N_7895,N_7523,N_7588);
nor U7896 (N_7896,N_7632,N_7531);
and U7897 (N_7897,N_7635,N_7511);
or U7898 (N_7898,N_7649,N_7633);
and U7899 (N_7899,N_7559,N_7661);
xor U7900 (N_7900,N_7659,N_7615);
xnor U7901 (N_7901,N_7534,N_7685);
nand U7902 (N_7902,N_7656,N_7545);
xnor U7903 (N_7903,N_7562,N_7688);
or U7904 (N_7904,N_7548,N_7712);
nand U7905 (N_7905,N_7650,N_7559);
and U7906 (N_7906,N_7643,N_7514);
nor U7907 (N_7907,N_7655,N_7689);
nand U7908 (N_7908,N_7575,N_7634);
and U7909 (N_7909,N_7550,N_7714);
and U7910 (N_7910,N_7555,N_7639);
xnor U7911 (N_7911,N_7512,N_7621);
nand U7912 (N_7912,N_7515,N_7616);
nand U7913 (N_7913,N_7659,N_7557);
nor U7914 (N_7914,N_7607,N_7657);
xnor U7915 (N_7915,N_7715,N_7659);
nand U7916 (N_7916,N_7676,N_7526);
nor U7917 (N_7917,N_7633,N_7556);
nor U7918 (N_7918,N_7505,N_7689);
or U7919 (N_7919,N_7503,N_7595);
nor U7920 (N_7920,N_7724,N_7590);
xnor U7921 (N_7921,N_7598,N_7551);
nand U7922 (N_7922,N_7514,N_7531);
or U7923 (N_7923,N_7715,N_7623);
and U7924 (N_7924,N_7558,N_7682);
and U7925 (N_7925,N_7675,N_7645);
nor U7926 (N_7926,N_7606,N_7593);
or U7927 (N_7927,N_7640,N_7691);
or U7928 (N_7928,N_7676,N_7699);
nand U7929 (N_7929,N_7719,N_7687);
and U7930 (N_7930,N_7673,N_7551);
nor U7931 (N_7931,N_7721,N_7515);
or U7932 (N_7932,N_7518,N_7591);
nor U7933 (N_7933,N_7715,N_7536);
or U7934 (N_7934,N_7627,N_7523);
nor U7935 (N_7935,N_7703,N_7675);
nand U7936 (N_7936,N_7680,N_7503);
xnor U7937 (N_7937,N_7538,N_7674);
and U7938 (N_7938,N_7575,N_7671);
nor U7939 (N_7939,N_7576,N_7697);
nand U7940 (N_7940,N_7579,N_7537);
nor U7941 (N_7941,N_7556,N_7737);
nand U7942 (N_7942,N_7561,N_7737);
and U7943 (N_7943,N_7635,N_7749);
nor U7944 (N_7944,N_7524,N_7620);
nand U7945 (N_7945,N_7521,N_7510);
nor U7946 (N_7946,N_7536,N_7516);
and U7947 (N_7947,N_7715,N_7647);
nand U7948 (N_7948,N_7595,N_7680);
nor U7949 (N_7949,N_7512,N_7716);
nand U7950 (N_7950,N_7732,N_7645);
nand U7951 (N_7951,N_7607,N_7701);
xor U7952 (N_7952,N_7713,N_7609);
and U7953 (N_7953,N_7729,N_7722);
xnor U7954 (N_7954,N_7556,N_7721);
or U7955 (N_7955,N_7556,N_7646);
nor U7956 (N_7956,N_7644,N_7657);
nand U7957 (N_7957,N_7727,N_7630);
nor U7958 (N_7958,N_7726,N_7511);
xnor U7959 (N_7959,N_7541,N_7577);
nor U7960 (N_7960,N_7733,N_7588);
nand U7961 (N_7961,N_7672,N_7629);
and U7962 (N_7962,N_7744,N_7657);
nor U7963 (N_7963,N_7582,N_7595);
nor U7964 (N_7964,N_7716,N_7698);
xor U7965 (N_7965,N_7573,N_7585);
nand U7966 (N_7966,N_7643,N_7704);
nand U7967 (N_7967,N_7722,N_7683);
and U7968 (N_7968,N_7512,N_7564);
xnor U7969 (N_7969,N_7549,N_7671);
and U7970 (N_7970,N_7721,N_7720);
and U7971 (N_7971,N_7727,N_7649);
xnor U7972 (N_7972,N_7658,N_7600);
xnor U7973 (N_7973,N_7522,N_7501);
nand U7974 (N_7974,N_7664,N_7627);
and U7975 (N_7975,N_7711,N_7680);
and U7976 (N_7976,N_7603,N_7579);
nor U7977 (N_7977,N_7522,N_7531);
xnor U7978 (N_7978,N_7588,N_7513);
or U7979 (N_7979,N_7563,N_7531);
or U7980 (N_7980,N_7645,N_7559);
or U7981 (N_7981,N_7703,N_7579);
and U7982 (N_7982,N_7722,N_7735);
nand U7983 (N_7983,N_7648,N_7590);
nand U7984 (N_7984,N_7722,N_7500);
or U7985 (N_7985,N_7549,N_7532);
and U7986 (N_7986,N_7727,N_7505);
nor U7987 (N_7987,N_7518,N_7555);
nand U7988 (N_7988,N_7726,N_7536);
xor U7989 (N_7989,N_7569,N_7679);
nand U7990 (N_7990,N_7652,N_7559);
nand U7991 (N_7991,N_7661,N_7601);
and U7992 (N_7992,N_7565,N_7517);
nor U7993 (N_7993,N_7725,N_7718);
xnor U7994 (N_7994,N_7568,N_7589);
and U7995 (N_7995,N_7537,N_7593);
or U7996 (N_7996,N_7629,N_7612);
xnor U7997 (N_7997,N_7606,N_7562);
or U7998 (N_7998,N_7653,N_7532);
and U7999 (N_7999,N_7592,N_7501);
nor U8000 (N_8000,N_7890,N_7962);
nor U8001 (N_8001,N_7980,N_7854);
xnor U8002 (N_8002,N_7918,N_7938);
xnor U8003 (N_8003,N_7947,N_7992);
nand U8004 (N_8004,N_7883,N_7793);
nand U8005 (N_8005,N_7973,N_7831);
and U8006 (N_8006,N_7878,N_7920);
nor U8007 (N_8007,N_7795,N_7921);
or U8008 (N_8008,N_7910,N_7950);
xnor U8009 (N_8009,N_7812,N_7750);
and U8010 (N_8010,N_7889,N_7966);
nand U8011 (N_8011,N_7948,N_7982);
nand U8012 (N_8012,N_7825,N_7909);
nor U8013 (N_8013,N_7827,N_7760);
and U8014 (N_8014,N_7850,N_7944);
xor U8015 (N_8015,N_7761,N_7993);
nor U8016 (N_8016,N_7880,N_7868);
or U8017 (N_8017,N_7971,N_7876);
nor U8018 (N_8018,N_7783,N_7939);
or U8019 (N_8019,N_7849,N_7904);
nor U8020 (N_8020,N_7914,N_7798);
xor U8021 (N_8021,N_7986,N_7835);
nand U8022 (N_8022,N_7797,N_7811);
or U8023 (N_8023,N_7927,N_7963);
xor U8024 (N_8024,N_7881,N_7861);
xor U8025 (N_8025,N_7885,N_7924);
nor U8026 (N_8026,N_7888,N_7975);
nand U8027 (N_8027,N_7900,N_7958);
nor U8028 (N_8028,N_7786,N_7829);
nor U8029 (N_8029,N_7832,N_7940);
nand U8030 (N_8030,N_7840,N_7857);
and U8031 (N_8031,N_7789,N_7942);
or U8032 (N_8032,N_7941,N_7778);
xor U8033 (N_8033,N_7870,N_7902);
or U8034 (N_8034,N_7931,N_7844);
or U8035 (N_8035,N_7926,N_7758);
and U8036 (N_8036,N_7806,N_7933);
and U8037 (N_8037,N_7837,N_7851);
or U8038 (N_8038,N_7979,N_7838);
xor U8039 (N_8039,N_7988,N_7913);
xor U8040 (N_8040,N_7893,N_7859);
and U8041 (N_8041,N_7932,N_7898);
and U8042 (N_8042,N_7807,N_7957);
xor U8043 (N_8043,N_7952,N_7802);
and U8044 (N_8044,N_7894,N_7908);
or U8045 (N_8045,N_7804,N_7946);
and U8046 (N_8046,N_7792,N_7871);
or U8047 (N_8047,N_7899,N_7998);
nor U8048 (N_8048,N_7862,N_7943);
nor U8049 (N_8049,N_7954,N_7886);
or U8050 (N_8050,N_7901,N_7949);
xor U8051 (N_8051,N_7945,N_7770);
and U8052 (N_8052,N_7964,N_7818);
xor U8053 (N_8053,N_7977,N_7803);
xnor U8054 (N_8054,N_7959,N_7858);
nand U8055 (N_8055,N_7821,N_7989);
nand U8056 (N_8056,N_7752,N_7824);
and U8057 (N_8057,N_7872,N_7784);
and U8058 (N_8058,N_7903,N_7810);
xnor U8059 (N_8059,N_7763,N_7905);
and U8060 (N_8060,N_7956,N_7777);
xor U8061 (N_8061,N_7934,N_7863);
nand U8062 (N_8062,N_7981,N_7874);
and U8063 (N_8063,N_7997,N_7765);
nand U8064 (N_8064,N_7774,N_7937);
xnor U8065 (N_8065,N_7843,N_7841);
and U8066 (N_8066,N_7855,N_7794);
nor U8067 (N_8067,N_7766,N_7995);
nor U8068 (N_8068,N_7801,N_7836);
and U8069 (N_8069,N_7891,N_7790);
or U8070 (N_8070,N_7771,N_7955);
nand U8071 (N_8071,N_7994,N_7873);
or U8072 (N_8072,N_7848,N_7936);
xnor U8073 (N_8073,N_7805,N_7974);
and U8074 (N_8074,N_7845,N_7953);
and U8075 (N_8075,N_7983,N_7895);
xor U8076 (N_8076,N_7756,N_7814);
nor U8077 (N_8077,N_7842,N_7751);
and U8078 (N_8078,N_7788,N_7864);
xnor U8079 (N_8079,N_7987,N_7985);
nor U8080 (N_8080,N_7757,N_7820);
or U8081 (N_8081,N_7907,N_7978);
and U8082 (N_8082,N_7839,N_7866);
or U8083 (N_8083,N_7767,N_7791);
nor U8084 (N_8084,N_7916,N_7867);
nand U8085 (N_8085,N_7796,N_7834);
nand U8086 (N_8086,N_7892,N_7846);
or U8087 (N_8087,N_7930,N_7815);
nor U8088 (N_8088,N_7951,N_7852);
or U8089 (N_8089,N_7877,N_7755);
nand U8090 (N_8090,N_7787,N_7999);
and U8091 (N_8091,N_7912,N_7822);
and U8092 (N_8092,N_7799,N_7928);
nand U8093 (N_8093,N_7813,N_7929);
nor U8094 (N_8094,N_7911,N_7919);
and U8095 (N_8095,N_7884,N_7967);
xnor U8096 (N_8096,N_7817,N_7800);
nor U8097 (N_8097,N_7869,N_7826);
and U8098 (N_8098,N_7976,N_7847);
and U8099 (N_8099,N_7776,N_7764);
nand U8100 (N_8100,N_7969,N_7769);
and U8101 (N_8101,N_7965,N_7970);
nor U8102 (N_8102,N_7853,N_7808);
or U8103 (N_8103,N_7753,N_7875);
nand U8104 (N_8104,N_7990,N_7925);
xor U8105 (N_8105,N_7882,N_7816);
nor U8106 (N_8106,N_7828,N_7809);
xor U8107 (N_8107,N_7780,N_7775);
xnor U8108 (N_8108,N_7860,N_7865);
and U8109 (N_8109,N_7772,N_7923);
nand U8110 (N_8110,N_7782,N_7830);
or U8111 (N_8111,N_7996,N_7984);
and U8112 (N_8112,N_7879,N_7773);
nor U8113 (N_8113,N_7915,N_7781);
xor U8114 (N_8114,N_7779,N_7906);
or U8115 (N_8115,N_7785,N_7991);
nor U8116 (N_8116,N_7972,N_7856);
nor U8117 (N_8117,N_7897,N_7935);
xor U8118 (N_8118,N_7823,N_7961);
xnor U8119 (N_8119,N_7960,N_7754);
xnor U8120 (N_8120,N_7819,N_7896);
xnor U8121 (N_8121,N_7922,N_7887);
and U8122 (N_8122,N_7762,N_7968);
and U8123 (N_8123,N_7917,N_7833);
or U8124 (N_8124,N_7759,N_7768);
and U8125 (N_8125,N_7904,N_7907);
and U8126 (N_8126,N_7993,N_7945);
and U8127 (N_8127,N_7880,N_7983);
and U8128 (N_8128,N_7774,N_7837);
xor U8129 (N_8129,N_7997,N_7942);
and U8130 (N_8130,N_7816,N_7866);
nand U8131 (N_8131,N_7871,N_7834);
xnor U8132 (N_8132,N_7796,N_7830);
nand U8133 (N_8133,N_7763,N_7827);
xnor U8134 (N_8134,N_7983,N_7966);
xnor U8135 (N_8135,N_7862,N_7882);
nand U8136 (N_8136,N_7854,N_7876);
and U8137 (N_8137,N_7834,N_7758);
xor U8138 (N_8138,N_7997,N_7798);
and U8139 (N_8139,N_7831,N_7881);
and U8140 (N_8140,N_7758,N_7990);
or U8141 (N_8141,N_7908,N_7948);
or U8142 (N_8142,N_7889,N_7808);
nand U8143 (N_8143,N_7817,N_7901);
or U8144 (N_8144,N_7962,N_7965);
nand U8145 (N_8145,N_7903,N_7973);
or U8146 (N_8146,N_7805,N_7944);
and U8147 (N_8147,N_7892,N_7883);
nor U8148 (N_8148,N_7968,N_7982);
and U8149 (N_8149,N_7827,N_7995);
and U8150 (N_8150,N_7873,N_7870);
nor U8151 (N_8151,N_7820,N_7781);
xnor U8152 (N_8152,N_7815,N_7814);
xor U8153 (N_8153,N_7782,N_7913);
and U8154 (N_8154,N_7967,N_7864);
or U8155 (N_8155,N_7915,N_7800);
nor U8156 (N_8156,N_7755,N_7787);
xnor U8157 (N_8157,N_7831,N_7972);
or U8158 (N_8158,N_7982,N_7895);
or U8159 (N_8159,N_7797,N_7824);
xor U8160 (N_8160,N_7895,N_7769);
nand U8161 (N_8161,N_7841,N_7807);
and U8162 (N_8162,N_7898,N_7882);
xor U8163 (N_8163,N_7941,N_7917);
and U8164 (N_8164,N_7755,N_7907);
nor U8165 (N_8165,N_7999,N_7969);
and U8166 (N_8166,N_7839,N_7791);
nor U8167 (N_8167,N_7914,N_7751);
xnor U8168 (N_8168,N_7785,N_7904);
and U8169 (N_8169,N_7877,N_7762);
xor U8170 (N_8170,N_7960,N_7891);
nor U8171 (N_8171,N_7995,N_7799);
nand U8172 (N_8172,N_7932,N_7956);
xnor U8173 (N_8173,N_7806,N_7795);
nand U8174 (N_8174,N_7894,N_7960);
or U8175 (N_8175,N_7969,N_7812);
nor U8176 (N_8176,N_7778,N_7914);
or U8177 (N_8177,N_7991,N_7977);
or U8178 (N_8178,N_7932,N_7849);
and U8179 (N_8179,N_7959,N_7861);
and U8180 (N_8180,N_7849,N_7804);
xor U8181 (N_8181,N_7762,N_7886);
nand U8182 (N_8182,N_7759,N_7887);
nor U8183 (N_8183,N_7999,N_7827);
and U8184 (N_8184,N_7863,N_7793);
xnor U8185 (N_8185,N_7766,N_7750);
nor U8186 (N_8186,N_7954,N_7804);
or U8187 (N_8187,N_7878,N_7823);
and U8188 (N_8188,N_7890,N_7756);
xnor U8189 (N_8189,N_7953,N_7876);
or U8190 (N_8190,N_7838,N_7848);
xnor U8191 (N_8191,N_7886,N_7775);
or U8192 (N_8192,N_7902,N_7802);
and U8193 (N_8193,N_7902,N_7916);
or U8194 (N_8194,N_7859,N_7803);
nand U8195 (N_8195,N_7788,N_7831);
xor U8196 (N_8196,N_7813,N_7806);
and U8197 (N_8197,N_7993,N_7801);
and U8198 (N_8198,N_7979,N_7998);
nor U8199 (N_8199,N_7907,N_7915);
xor U8200 (N_8200,N_7846,N_7936);
and U8201 (N_8201,N_7818,N_7848);
nor U8202 (N_8202,N_7861,N_7757);
nand U8203 (N_8203,N_7986,N_7969);
xnor U8204 (N_8204,N_7888,N_7766);
xor U8205 (N_8205,N_7982,N_7847);
nor U8206 (N_8206,N_7765,N_7876);
nor U8207 (N_8207,N_7873,N_7802);
nor U8208 (N_8208,N_7805,N_7765);
or U8209 (N_8209,N_7831,N_7948);
nor U8210 (N_8210,N_7782,N_7881);
and U8211 (N_8211,N_7895,N_7914);
or U8212 (N_8212,N_7897,N_7847);
nor U8213 (N_8213,N_7789,N_7906);
nand U8214 (N_8214,N_7915,N_7972);
nor U8215 (N_8215,N_7982,N_7913);
and U8216 (N_8216,N_7959,N_7960);
or U8217 (N_8217,N_7876,N_7945);
and U8218 (N_8218,N_7859,N_7856);
and U8219 (N_8219,N_7976,N_7923);
nor U8220 (N_8220,N_7831,N_7930);
nand U8221 (N_8221,N_7997,N_7807);
nand U8222 (N_8222,N_7822,N_7771);
nor U8223 (N_8223,N_7801,N_7986);
nand U8224 (N_8224,N_7932,N_7960);
and U8225 (N_8225,N_7896,N_7974);
xor U8226 (N_8226,N_7815,N_7834);
or U8227 (N_8227,N_7992,N_7943);
and U8228 (N_8228,N_7893,N_7790);
and U8229 (N_8229,N_7840,N_7997);
nand U8230 (N_8230,N_7940,N_7992);
nor U8231 (N_8231,N_7965,N_7752);
or U8232 (N_8232,N_7841,N_7818);
and U8233 (N_8233,N_7915,N_7750);
nand U8234 (N_8234,N_7870,N_7831);
xor U8235 (N_8235,N_7897,N_7907);
or U8236 (N_8236,N_7962,N_7924);
nand U8237 (N_8237,N_7926,N_7988);
xnor U8238 (N_8238,N_7978,N_7919);
or U8239 (N_8239,N_7924,N_7774);
nor U8240 (N_8240,N_7797,N_7891);
nand U8241 (N_8241,N_7885,N_7918);
and U8242 (N_8242,N_7763,N_7911);
or U8243 (N_8243,N_7779,N_7817);
or U8244 (N_8244,N_7816,N_7857);
nor U8245 (N_8245,N_7785,N_7761);
and U8246 (N_8246,N_7812,N_7966);
nand U8247 (N_8247,N_7965,N_7839);
and U8248 (N_8248,N_7968,N_7837);
xor U8249 (N_8249,N_7751,N_7982);
nand U8250 (N_8250,N_8158,N_8228);
and U8251 (N_8251,N_8152,N_8095);
xnor U8252 (N_8252,N_8077,N_8115);
and U8253 (N_8253,N_8070,N_8119);
or U8254 (N_8254,N_8105,N_8169);
or U8255 (N_8255,N_8054,N_8075);
nor U8256 (N_8256,N_8197,N_8028);
and U8257 (N_8257,N_8202,N_8109);
nand U8258 (N_8258,N_8160,N_8029);
and U8259 (N_8259,N_8023,N_8080);
nand U8260 (N_8260,N_8231,N_8003);
xnor U8261 (N_8261,N_8089,N_8014);
xor U8262 (N_8262,N_8235,N_8009);
or U8263 (N_8263,N_8181,N_8087);
or U8264 (N_8264,N_8011,N_8190);
or U8265 (N_8265,N_8225,N_8219);
or U8266 (N_8266,N_8198,N_8092);
nand U8267 (N_8267,N_8141,N_8108);
nand U8268 (N_8268,N_8199,N_8034);
xnor U8269 (N_8269,N_8024,N_8211);
nor U8270 (N_8270,N_8093,N_8144);
nand U8271 (N_8271,N_8037,N_8229);
nor U8272 (N_8272,N_8082,N_8010);
nor U8273 (N_8273,N_8203,N_8149);
xnor U8274 (N_8274,N_8043,N_8059);
nand U8275 (N_8275,N_8163,N_8084);
and U8276 (N_8276,N_8186,N_8142);
nor U8277 (N_8277,N_8127,N_8153);
nor U8278 (N_8278,N_8207,N_8061);
nand U8279 (N_8279,N_8122,N_8124);
nand U8280 (N_8280,N_8155,N_8137);
and U8281 (N_8281,N_8106,N_8002);
or U8282 (N_8282,N_8191,N_8143);
xor U8283 (N_8283,N_8001,N_8175);
and U8284 (N_8284,N_8019,N_8173);
and U8285 (N_8285,N_8222,N_8123);
nand U8286 (N_8286,N_8074,N_8146);
xnor U8287 (N_8287,N_8090,N_8006);
nand U8288 (N_8288,N_8136,N_8150);
xor U8289 (N_8289,N_8097,N_8147);
nor U8290 (N_8290,N_8218,N_8171);
xor U8291 (N_8291,N_8154,N_8188);
and U8292 (N_8292,N_8068,N_8110);
xnor U8293 (N_8293,N_8187,N_8226);
and U8294 (N_8294,N_8069,N_8052);
xor U8295 (N_8295,N_8102,N_8208);
and U8296 (N_8296,N_8145,N_8140);
and U8297 (N_8297,N_8193,N_8118);
or U8298 (N_8298,N_8026,N_8189);
or U8299 (N_8299,N_8081,N_8239);
xnor U8300 (N_8300,N_8030,N_8128);
and U8301 (N_8301,N_8099,N_8096);
and U8302 (N_8302,N_8020,N_8168);
or U8303 (N_8303,N_8248,N_8129);
or U8304 (N_8304,N_8174,N_8016);
nor U8305 (N_8305,N_8172,N_8088);
or U8306 (N_8306,N_8015,N_8206);
nor U8307 (N_8307,N_8053,N_8148);
nor U8308 (N_8308,N_8008,N_8067);
xor U8309 (N_8309,N_8072,N_8100);
and U8310 (N_8310,N_8164,N_8247);
nor U8311 (N_8311,N_8161,N_8103);
nor U8312 (N_8312,N_8241,N_8049);
and U8313 (N_8313,N_8117,N_8035);
nor U8314 (N_8314,N_8004,N_8033);
nor U8315 (N_8315,N_8085,N_8114);
or U8316 (N_8316,N_8138,N_8214);
or U8317 (N_8317,N_8064,N_8139);
or U8318 (N_8318,N_8063,N_8176);
and U8319 (N_8319,N_8185,N_8178);
nor U8320 (N_8320,N_8057,N_8055);
and U8321 (N_8321,N_8167,N_8132);
or U8322 (N_8322,N_8159,N_8204);
or U8323 (N_8323,N_8121,N_8047);
xor U8324 (N_8324,N_8183,N_8116);
nor U8325 (N_8325,N_8113,N_8039);
xnor U8326 (N_8326,N_8244,N_8133);
or U8327 (N_8327,N_8078,N_8220);
xor U8328 (N_8328,N_8134,N_8005);
or U8329 (N_8329,N_8111,N_8083);
or U8330 (N_8330,N_8212,N_8201);
or U8331 (N_8331,N_8021,N_8126);
nand U8332 (N_8332,N_8240,N_8194);
xor U8333 (N_8333,N_8200,N_8101);
xnor U8334 (N_8334,N_8065,N_8036);
nand U8335 (N_8335,N_8213,N_8232);
or U8336 (N_8336,N_8184,N_8062);
xor U8337 (N_8337,N_8071,N_8195);
nand U8338 (N_8338,N_8086,N_8227);
and U8339 (N_8339,N_8058,N_8156);
nor U8340 (N_8340,N_8098,N_8217);
and U8341 (N_8341,N_8162,N_8066);
nand U8342 (N_8342,N_8205,N_8215);
nor U8343 (N_8343,N_8131,N_8079);
nand U8344 (N_8344,N_8179,N_8038);
or U8345 (N_8345,N_8025,N_8040);
xor U8346 (N_8346,N_8073,N_8044);
and U8347 (N_8347,N_8042,N_8051);
nor U8348 (N_8348,N_8151,N_8233);
or U8349 (N_8349,N_8120,N_8135);
xor U8350 (N_8350,N_8107,N_8245);
and U8351 (N_8351,N_8022,N_8236);
nand U8352 (N_8352,N_8018,N_8165);
nor U8353 (N_8353,N_8041,N_8032);
or U8354 (N_8354,N_8007,N_8046);
or U8355 (N_8355,N_8013,N_8056);
or U8356 (N_8356,N_8246,N_8050);
nand U8357 (N_8357,N_8045,N_8177);
xnor U8358 (N_8358,N_8017,N_8031);
nand U8359 (N_8359,N_8104,N_8091);
and U8360 (N_8360,N_8180,N_8237);
and U8361 (N_8361,N_8112,N_8224);
or U8362 (N_8362,N_8209,N_8094);
nor U8363 (N_8363,N_8166,N_8210);
and U8364 (N_8364,N_8027,N_8238);
nor U8365 (N_8365,N_8242,N_8221);
xnor U8366 (N_8366,N_8196,N_8182);
and U8367 (N_8367,N_8130,N_8230);
and U8368 (N_8368,N_8012,N_8000);
xor U8369 (N_8369,N_8234,N_8170);
nand U8370 (N_8370,N_8048,N_8060);
nand U8371 (N_8371,N_8249,N_8223);
nand U8372 (N_8372,N_8125,N_8157);
xnor U8373 (N_8373,N_8076,N_8192);
nand U8374 (N_8374,N_8243,N_8216);
xnor U8375 (N_8375,N_8164,N_8112);
and U8376 (N_8376,N_8016,N_8171);
xnor U8377 (N_8377,N_8066,N_8240);
or U8378 (N_8378,N_8186,N_8141);
or U8379 (N_8379,N_8199,N_8184);
nand U8380 (N_8380,N_8075,N_8204);
or U8381 (N_8381,N_8047,N_8094);
nand U8382 (N_8382,N_8082,N_8079);
or U8383 (N_8383,N_8089,N_8083);
xor U8384 (N_8384,N_8016,N_8052);
xnor U8385 (N_8385,N_8027,N_8131);
or U8386 (N_8386,N_8102,N_8013);
nor U8387 (N_8387,N_8177,N_8121);
xnor U8388 (N_8388,N_8172,N_8061);
xor U8389 (N_8389,N_8119,N_8191);
xnor U8390 (N_8390,N_8207,N_8247);
xor U8391 (N_8391,N_8245,N_8092);
and U8392 (N_8392,N_8047,N_8001);
xor U8393 (N_8393,N_8028,N_8203);
xor U8394 (N_8394,N_8160,N_8101);
nand U8395 (N_8395,N_8045,N_8195);
and U8396 (N_8396,N_8056,N_8219);
xnor U8397 (N_8397,N_8082,N_8202);
and U8398 (N_8398,N_8118,N_8081);
and U8399 (N_8399,N_8033,N_8153);
xnor U8400 (N_8400,N_8157,N_8088);
and U8401 (N_8401,N_8217,N_8101);
and U8402 (N_8402,N_8081,N_8072);
nand U8403 (N_8403,N_8247,N_8008);
or U8404 (N_8404,N_8001,N_8210);
and U8405 (N_8405,N_8119,N_8208);
and U8406 (N_8406,N_8101,N_8123);
or U8407 (N_8407,N_8073,N_8177);
nor U8408 (N_8408,N_8099,N_8115);
and U8409 (N_8409,N_8018,N_8155);
xor U8410 (N_8410,N_8079,N_8027);
and U8411 (N_8411,N_8249,N_8161);
and U8412 (N_8412,N_8156,N_8208);
nor U8413 (N_8413,N_8116,N_8227);
nand U8414 (N_8414,N_8037,N_8054);
nor U8415 (N_8415,N_8024,N_8160);
and U8416 (N_8416,N_8210,N_8170);
nor U8417 (N_8417,N_8191,N_8079);
nor U8418 (N_8418,N_8229,N_8014);
xor U8419 (N_8419,N_8003,N_8065);
and U8420 (N_8420,N_8026,N_8183);
nor U8421 (N_8421,N_8188,N_8079);
nand U8422 (N_8422,N_8103,N_8058);
xor U8423 (N_8423,N_8057,N_8001);
or U8424 (N_8424,N_8173,N_8061);
or U8425 (N_8425,N_8092,N_8143);
and U8426 (N_8426,N_8164,N_8019);
and U8427 (N_8427,N_8170,N_8028);
nand U8428 (N_8428,N_8007,N_8048);
xnor U8429 (N_8429,N_8199,N_8197);
nor U8430 (N_8430,N_8190,N_8236);
nand U8431 (N_8431,N_8172,N_8233);
nand U8432 (N_8432,N_8092,N_8202);
xor U8433 (N_8433,N_8227,N_8173);
and U8434 (N_8434,N_8109,N_8208);
and U8435 (N_8435,N_8025,N_8094);
or U8436 (N_8436,N_8031,N_8171);
nand U8437 (N_8437,N_8221,N_8074);
nor U8438 (N_8438,N_8011,N_8109);
nand U8439 (N_8439,N_8212,N_8085);
nand U8440 (N_8440,N_8234,N_8035);
xor U8441 (N_8441,N_8119,N_8178);
or U8442 (N_8442,N_8131,N_8084);
xnor U8443 (N_8443,N_8015,N_8119);
nand U8444 (N_8444,N_8052,N_8058);
xor U8445 (N_8445,N_8064,N_8074);
nand U8446 (N_8446,N_8186,N_8160);
xor U8447 (N_8447,N_8236,N_8027);
nand U8448 (N_8448,N_8126,N_8103);
or U8449 (N_8449,N_8217,N_8179);
and U8450 (N_8450,N_8075,N_8019);
nor U8451 (N_8451,N_8045,N_8040);
nor U8452 (N_8452,N_8187,N_8092);
nand U8453 (N_8453,N_8004,N_8000);
or U8454 (N_8454,N_8232,N_8219);
nand U8455 (N_8455,N_8044,N_8179);
nor U8456 (N_8456,N_8156,N_8036);
or U8457 (N_8457,N_8010,N_8247);
xor U8458 (N_8458,N_8009,N_8213);
nand U8459 (N_8459,N_8131,N_8219);
nor U8460 (N_8460,N_8089,N_8060);
xor U8461 (N_8461,N_8181,N_8085);
or U8462 (N_8462,N_8187,N_8113);
xnor U8463 (N_8463,N_8034,N_8030);
xor U8464 (N_8464,N_8069,N_8238);
or U8465 (N_8465,N_8092,N_8225);
xor U8466 (N_8466,N_8239,N_8016);
nand U8467 (N_8467,N_8190,N_8089);
nand U8468 (N_8468,N_8049,N_8160);
xor U8469 (N_8469,N_8172,N_8185);
nor U8470 (N_8470,N_8090,N_8239);
or U8471 (N_8471,N_8112,N_8226);
nand U8472 (N_8472,N_8245,N_8091);
and U8473 (N_8473,N_8014,N_8049);
nor U8474 (N_8474,N_8166,N_8071);
and U8475 (N_8475,N_8248,N_8028);
nand U8476 (N_8476,N_8133,N_8152);
nand U8477 (N_8477,N_8175,N_8155);
and U8478 (N_8478,N_8164,N_8081);
and U8479 (N_8479,N_8194,N_8221);
nor U8480 (N_8480,N_8109,N_8163);
xor U8481 (N_8481,N_8133,N_8007);
or U8482 (N_8482,N_8217,N_8029);
xnor U8483 (N_8483,N_8249,N_8241);
nand U8484 (N_8484,N_8067,N_8201);
xor U8485 (N_8485,N_8192,N_8164);
nand U8486 (N_8486,N_8159,N_8162);
xnor U8487 (N_8487,N_8071,N_8223);
or U8488 (N_8488,N_8048,N_8249);
nor U8489 (N_8489,N_8059,N_8141);
nor U8490 (N_8490,N_8202,N_8043);
nor U8491 (N_8491,N_8087,N_8048);
xor U8492 (N_8492,N_8124,N_8025);
xnor U8493 (N_8493,N_8151,N_8120);
nand U8494 (N_8494,N_8192,N_8249);
nor U8495 (N_8495,N_8229,N_8054);
xnor U8496 (N_8496,N_8020,N_8233);
xor U8497 (N_8497,N_8076,N_8079);
xnor U8498 (N_8498,N_8230,N_8212);
nor U8499 (N_8499,N_8163,N_8051);
xnor U8500 (N_8500,N_8333,N_8376);
xor U8501 (N_8501,N_8288,N_8426);
xnor U8502 (N_8502,N_8457,N_8350);
nand U8503 (N_8503,N_8418,N_8352);
nand U8504 (N_8504,N_8398,N_8444);
xnor U8505 (N_8505,N_8462,N_8357);
nand U8506 (N_8506,N_8332,N_8477);
nor U8507 (N_8507,N_8468,N_8252);
xor U8508 (N_8508,N_8329,N_8292);
nor U8509 (N_8509,N_8436,N_8429);
nand U8510 (N_8510,N_8309,N_8365);
nand U8511 (N_8511,N_8262,N_8289);
and U8512 (N_8512,N_8314,N_8282);
nand U8513 (N_8513,N_8264,N_8312);
nor U8514 (N_8514,N_8318,N_8271);
xor U8515 (N_8515,N_8406,N_8498);
xor U8516 (N_8516,N_8395,N_8491);
xor U8517 (N_8517,N_8277,N_8300);
or U8518 (N_8518,N_8294,N_8308);
or U8519 (N_8519,N_8327,N_8479);
nand U8520 (N_8520,N_8290,N_8257);
nand U8521 (N_8521,N_8443,N_8409);
nand U8522 (N_8522,N_8391,N_8475);
or U8523 (N_8523,N_8484,N_8305);
and U8524 (N_8524,N_8400,N_8280);
and U8525 (N_8525,N_8354,N_8311);
and U8526 (N_8526,N_8349,N_8325);
nand U8527 (N_8527,N_8412,N_8323);
nand U8528 (N_8528,N_8270,N_8480);
nand U8529 (N_8529,N_8346,N_8483);
xnor U8530 (N_8530,N_8343,N_8416);
nand U8531 (N_8531,N_8362,N_8466);
nor U8532 (N_8532,N_8303,N_8393);
nand U8533 (N_8533,N_8404,N_8263);
and U8534 (N_8534,N_8268,N_8254);
or U8535 (N_8535,N_8432,N_8250);
xnor U8536 (N_8536,N_8298,N_8339);
xnor U8537 (N_8537,N_8451,N_8439);
or U8538 (N_8538,N_8478,N_8330);
nor U8539 (N_8539,N_8390,N_8431);
xor U8540 (N_8540,N_8403,N_8379);
nand U8541 (N_8541,N_8453,N_8369);
nor U8542 (N_8542,N_8359,N_8276);
nor U8543 (N_8543,N_8320,N_8413);
or U8544 (N_8544,N_8425,N_8299);
and U8545 (N_8545,N_8260,N_8407);
nand U8546 (N_8546,N_8341,N_8421);
and U8547 (N_8547,N_8291,N_8363);
xnor U8548 (N_8548,N_8384,N_8496);
nand U8549 (N_8549,N_8251,N_8495);
nor U8550 (N_8550,N_8415,N_8402);
and U8551 (N_8551,N_8378,N_8417);
nor U8552 (N_8552,N_8470,N_8322);
and U8553 (N_8553,N_8284,N_8437);
xnor U8554 (N_8554,N_8422,N_8319);
and U8555 (N_8555,N_8313,N_8304);
or U8556 (N_8556,N_8338,N_8489);
xnor U8557 (N_8557,N_8366,N_8360);
xor U8558 (N_8558,N_8399,N_8317);
nor U8559 (N_8559,N_8255,N_8396);
or U8560 (N_8560,N_8337,N_8445);
or U8561 (N_8561,N_8279,N_8356);
xnor U8562 (N_8562,N_8410,N_8485);
and U8563 (N_8563,N_8256,N_8328);
nand U8564 (N_8564,N_8374,N_8497);
and U8565 (N_8565,N_8316,N_8267);
nor U8566 (N_8566,N_8377,N_8287);
nor U8567 (N_8567,N_8324,N_8296);
nand U8568 (N_8568,N_8471,N_8351);
or U8569 (N_8569,N_8342,N_8430);
xnor U8570 (N_8570,N_8438,N_8419);
or U8571 (N_8571,N_8448,N_8427);
or U8572 (N_8572,N_8253,N_8394);
or U8573 (N_8573,N_8499,N_8301);
nor U8574 (N_8574,N_8482,N_8405);
or U8575 (N_8575,N_8464,N_8293);
and U8576 (N_8576,N_8435,N_8459);
nand U8577 (N_8577,N_8494,N_8307);
xor U8578 (N_8578,N_8486,N_8414);
or U8579 (N_8579,N_8297,N_8321);
and U8580 (N_8580,N_8274,N_8458);
nand U8581 (N_8581,N_8456,N_8433);
nand U8582 (N_8582,N_8392,N_8281);
nand U8583 (N_8583,N_8285,N_8434);
xor U8584 (N_8584,N_8355,N_8408);
or U8585 (N_8585,N_8420,N_8382);
or U8586 (N_8586,N_8306,N_8273);
xnor U8587 (N_8587,N_8272,N_8474);
nand U8588 (N_8588,N_8259,N_8278);
nand U8589 (N_8589,N_8455,N_8315);
and U8590 (N_8590,N_8310,N_8335);
nand U8591 (N_8591,N_8440,N_8460);
or U8592 (N_8592,N_8353,N_8467);
xor U8593 (N_8593,N_8266,N_8441);
nand U8594 (N_8594,N_8383,N_8388);
and U8595 (N_8595,N_8368,N_8386);
and U8596 (N_8596,N_8476,N_8295);
nor U8597 (N_8597,N_8442,N_8447);
or U8598 (N_8598,N_8302,N_8469);
or U8599 (N_8599,N_8450,N_8387);
or U8600 (N_8600,N_8344,N_8454);
xnor U8601 (N_8601,N_8372,N_8465);
nand U8602 (N_8602,N_8275,N_8261);
nand U8603 (N_8603,N_8401,N_8493);
or U8604 (N_8604,N_8269,N_8473);
or U8605 (N_8605,N_8487,N_8286);
nor U8606 (N_8606,N_8258,N_8283);
nor U8607 (N_8607,N_8361,N_8492);
or U8608 (N_8608,N_8364,N_8481);
or U8609 (N_8609,N_8446,N_8340);
or U8610 (N_8610,N_8428,N_8348);
or U8611 (N_8611,N_8452,N_8490);
or U8612 (N_8612,N_8381,N_8371);
nor U8613 (N_8613,N_8423,N_8331);
nand U8614 (N_8614,N_8265,N_8370);
nand U8615 (N_8615,N_8375,N_8389);
xnor U8616 (N_8616,N_8358,N_8397);
nand U8617 (N_8617,N_8347,N_8463);
xnor U8618 (N_8618,N_8373,N_8411);
xor U8619 (N_8619,N_8380,N_8472);
xnor U8620 (N_8620,N_8461,N_8385);
nor U8621 (N_8621,N_8334,N_8336);
nand U8622 (N_8622,N_8424,N_8488);
nand U8623 (N_8623,N_8345,N_8367);
or U8624 (N_8624,N_8326,N_8449);
xnor U8625 (N_8625,N_8350,N_8394);
nor U8626 (N_8626,N_8384,N_8453);
nand U8627 (N_8627,N_8288,N_8360);
or U8628 (N_8628,N_8335,N_8457);
or U8629 (N_8629,N_8450,N_8325);
and U8630 (N_8630,N_8453,N_8477);
nand U8631 (N_8631,N_8451,N_8364);
xor U8632 (N_8632,N_8365,N_8412);
or U8633 (N_8633,N_8329,N_8495);
nand U8634 (N_8634,N_8421,N_8366);
nor U8635 (N_8635,N_8457,N_8364);
and U8636 (N_8636,N_8321,N_8339);
nor U8637 (N_8637,N_8422,N_8463);
xor U8638 (N_8638,N_8269,N_8340);
xor U8639 (N_8639,N_8343,N_8405);
xnor U8640 (N_8640,N_8395,N_8465);
xor U8641 (N_8641,N_8288,N_8275);
nand U8642 (N_8642,N_8409,N_8383);
and U8643 (N_8643,N_8302,N_8317);
nor U8644 (N_8644,N_8452,N_8410);
nand U8645 (N_8645,N_8408,N_8253);
or U8646 (N_8646,N_8289,N_8317);
xor U8647 (N_8647,N_8462,N_8495);
nor U8648 (N_8648,N_8449,N_8350);
or U8649 (N_8649,N_8499,N_8252);
nor U8650 (N_8650,N_8489,N_8415);
xor U8651 (N_8651,N_8460,N_8319);
or U8652 (N_8652,N_8484,N_8286);
nand U8653 (N_8653,N_8386,N_8294);
nand U8654 (N_8654,N_8375,N_8259);
and U8655 (N_8655,N_8269,N_8358);
nand U8656 (N_8656,N_8252,N_8405);
or U8657 (N_8657,N_8372,N_8444);
nor U8658 (N_8658,N_8252,N_8489);
xor U8659 (N_8659,N_8404,N_8357);
and U8660 (N_8660,N_8348,N_8418);
nand U8661 (N_8661,N_8471,N_8475);
xnor U8662 (N_8662,N_8487,N_8462);
nand U8663 (N_8663,N_8419,N_8464);
nand U8664 (N_8664,N_8270,N_8367);
nor U8665 (N_8665,N_8392,N_8271);
nor U8666 (N_8666,N_8263,N_8327);
xnor U8667 (N_8667,N_8255,N_8288);
or U8668 (N_8668,N_8296,N_8404);
nand U8669 (N_8669,N_8285,N_8485);
or U8670 (N_8670,N_8353,N_8348);
nor U8671 (N_8671,N_8443,N_8255);
or U8672 (N_8672,N_8257,N_8273);
nand U8673 (N_8673,N_8405,N_8487);
nor U8674 (N_8674,N_8262,N_8292);
nor U8675 (N_8675,N_8318,N_8383);
and U8676 (N_8676,N_8463,N_8304);
xnor U8677 (N_8677,N_8254,N_8272);
nor U8678 (N_8678,N_8344,N_8485);
nand U8679 (N_8679,N_8268,N_8280);
nor U8680 (N_8680,N_8465,N_8323);
and U8681 (N_8681,N_8472,N_8374);
nor U8682 (N_8682,N_8310,N_8443);
xor U8683 (N_8683,N_8364,N_8380);
nand U8684 (N_8684,N_8459,N_8334);
and U8685 (N_8685,N_8334,N_8276);
xor U8686 (N_8686,N_8389,N_8475);
xor U8687 (N_8687,N_8293,N_8269);
xnor U8688 (N_8688,N_8262,N_8297);
or U8689 (N_8689,N_8408,N_8391);
or U8690 (N_8690,N_8323,N_8263);
nor U8691 (N_8691,N_8399,N_8308);
xnor U8692 (N_8692,N_8385,N_8267);
nor U8693 (N_8693,N_8471,N_8277);
nand U8694 (N_8694,N_8468,N_8331);
nand U8695 (N_8695,N_8322,N_8434);
nand U8696 (N_8696,N_8275,N_8348);
xnor U8697 (N_8697,N_8396,N_8389);
and U8698 (N_8698,N_8487,N_8348);
xor U8699 (N_8699,N_8306,N_8403);
nand U8700 (N_8700,N_8250,N_8357);
or U8701 (N_8701,N_8477,N_8417);
nor U8702 (N_8702,N_8302,N_8367);
or U8703 (N_8703,N_8341,N_8290);
and U8704 (N_8704,N_8291,N_8295);
or U8705 (N_8705,N_8333,N_8339);
and U8706 (N_8706,N_8370,N_8384);
or U8707 (N_8707,N_8496,N_8294);
xor U8708 (N_8708,N_8314,N_8360);
xnor U8709 (N_8709,N_8472,N_8409);
nand U8710 (N_8710,N_8364,N_8494);
nor U8711 (N_8711,N_8336,N_8252);
xor U8712 (N_8712,N_8254,N_8473);
nand U8713 (N_8713,N_8462,N_8490);
or U8714 (N_8714,N_8421,N_8430);
xnor U8715 (N_8715,N_8279,N_8326);
nor U8716 (N_8716,N_8469,N_8398);
or U8717 (N_8717,N_8335,N_8313);
xnor U8718 (N_8718,N_8380,N_8268);
nand U8719 (N_8719,N_8453,N_8376);
nor U8720 (N_8720,N_8330,N_8326);
or U8721 (N_8721,N_8467,N_8450);
nor U8722 (N_8722,N_8416,N_8497);
and U8723 (N_8723,N_8405,N_8304);
xnor U8724 (N_8724,N_8477,N_8357);
or U8725 (N_8725,N_8427,N_8495);
and U8726 (N_8726,N_8464,N_8292);
nand U8727 (N_8727,N_8345,N_8464);
and U8728 (N_8728,N_8282,N_8268);
or U8729 (N_8729,N_8262,N_8466);
and U8730 (N_8730,N_8261,N_8381);
nand U8731 (N_8731,N_8262,N_8489);
nor U8732 (N_8732,N_8302,N_8426);
or U8733 (N_8733,N_8301,N_8381);
nor U8734 (N_8734,N_8364,N_8498);
and U8735 (N_8735,N_8402,N_8294);
or U8736 (N_8736,N_8420,N_8349);
or U8737 (N_8737,N_8370,N_8488);
and U8738 (N_8738,N_8425,N_8380);
nor U8739 (N_8739,N_8296,N_8337);
or U8740 (N_8740,N_8494,N_8381);
or U8741 (N_8741,N_8398,N_8250);
xnor U8742 (N_8742,N_8446,N_8468);
or U8743 (N_8743,N_8461,N_8288);
nor U8744 (N_8744,N_8274,N_8463);
or U8745 (N_8745,N_8324,N_8334);
or U8746 (N_8746,N_8390,N_8474);
nor U8747 (N_8747,N_8418,N_8475);
nand U8748 (N_8748,N_8358,N_8283);
nand U8749 (N_8749,N_8303,N_8442);
nand U8750 (N_8750,N_8667,N_8707);
or U8751 (N_8751,N_8551,N_8749);
or U8752 (N_8752,N_8654,N_8606);
nand U8753 (N_8753,N_8748,N_8669);
and U8754 (N_8754,N_8611,N_8735);
xnor U8755 (N_8755,N_8536,N_8695);
or U8756 (N_8756,N_8648,N_8603);
xor U8757 (N_8757,N_8513,N_8670);
nor U8758 (N_8758,N_8562,N_8689);
nor U8759 (N_8759,N_8715,N_8526);
and U8760 (N_8760,N_8702,N_8737);
nand U8761 (N_8761,N_8601,N_8580);
xnor U8762 (N_8762,N_8607,N_8691);
and U8763 (N_8763,N_8539,N_8547);
and U8764 (N_8764,N_8560,N_8509);
nor U8765 (N_8765,N_8527,N_8506);
nor U8766 (N_8766,N_8525,N_8598);
or U8767 (N_8767,N_8716,N_8535);
nor U8768 (N_8768,N_8596,N_8550);
or U8769 (N_8769,N_8665,N_8576);
nand U8770 (N_8770,N_8555,N_8587);
xnor U8771 (N_8771,N_8676,N_8677);
and U8772 (N_8772,N_8714,N_8668);
nor U8773 (N_8773,N_8659,N_8679);
or U8774 (N_8774,N_8522,N_8646);
nor U8775 (N_8775,N_8593,N_8719);
nor U8776 (N_8776,N_8616,N_8556);
and U8777 (N_8777,N_8652,N_8618);
or U8778 (N_8778,N_8684,N_8635);
nor U8779 (N_8779,N_8696,N_8521);
nor U8780 (N_8780,N_8740,N_8730);
and U8781 (N_8781,N_8733,N_8586);
and U8782 (N_8782,N_8704,N_8626);
nand U8783 (N_8783,N_8741,N_8682);
nor U8784 (N_8784,N_8542,N_8680);
nor U8785 (N_8785,N_8502,N_8701);
xnor U8786 (N_8786,N_8615,N_8627);
nor U8787 (N_8787,N_8747,N_8583);
or U8788 (N_8788,N_8540,N_8674);
xnor U8789 (N_8789,N_8655,N_8608);
or U8790 (N_8790,N_8563,N_8514);
nor U8791 (N_8791,N_8657,N_8686);
nand U8792 (N_8792,N_8564,N_8683);
nor U8793 (N_8793,N_8561,N_8675);
nand U8794 (N_8794,N_8636,N_8722);
nor U8795 (N_8795,N_8694,N_8570);
nand U8796 (N_8796,N_8738,N_8575);
nand U8797 (N_8797,N_8569,N_8666);
and U8798 (N_8798,N_8545,N_8508);
xnor U8799 (N_8799,N_8571,N_8544);
xor U8800 (N_8800,N_8706,N_8724);
and U8801 (N_8801,N_8632,N_8644);
nand U8802 (N_8802,N_8692,N_8661);
nand U8803 (N_8803,N_8725,N_8531);
nor U8804 (N_8804,N_8731,N_8621);
nand U8805 (N_8805,N_8612,N_8543);
and U8806 (N_8806,N_8577,N_8662);
and U8807 (N_8807,N_8515,N_8519);
and U8808 (N_8808,N_8663,N_8595);
xor U8809 (N_8809,N_8638,N_8639);
nand U8810 (N_8810,N_8641,N_8688);
or U8811 (N_8811,N_8708,N_8697);
and U8812 (N_8812,N_8610,N_8501);
nor U8813 (N_8813,N_8524,N_8734);
and U8814 (N_8814,N_8567,N_8712);
nand U8815 (N_8815,N_8673,N_8718);
or U8816 (N_8816,N_8705,N_8507);
and U8817 (N_8817,N_8637,N_8510);
nor U8818 (N_8818,N_8541,N_8711);
nor U8819 (N_8819,N_8728,N_8709);
or U8820 (N_8820,N_8744,N_8518);
nor U8821 (N_8821,N_8630,N_8572);
and U8822 (N_8822,N_8671,N_8651);
or U8823 (N_8823,N_8642,N_8614);
nor U8824 (N_8824,N_8631,N_8720);
nand U8825 (N_8825,N_8681,N_8605);
nor U8826 (N_8826,N_8678,N_8504);
and U8827 (N_8827,N_8745,N_8685);
nor U8828 (N_8828,N_8529,N_8710);
or U8829 (N_8829,N_8578,N_8589);
or U8830 (N_8830,N_8619,N_8546);
xnor U8831 (N_8831,N_8698,N_8559);
or U8832 (N_8832,N_8623,N_8643);
nand U8833 (N_8833,N_8574,N_8602);
nor U8834 (N_8834,N_8594,N_8537);
nand U8835 (N_8835,N_8558,N_8505);
xnor U8836 (N_8836,N_8512,N_8520);
or U8837 (N_8837,N_8628,N_8653);
nor U8838 (N_8838,N_8503,N_8511);
nor U8839 (N_8839,N_8729,N_8528);
nand U8840 (N_8840,N_8742,N_8664);
nor U8841 (N_8841,N_8597,N_8693);
and U8842 (N_8842,N_8534,N_8703);
nand U8843 (N_8843,N_8532,N_8656);
nor U8844 (N_8844,N_8746,N_8565);
xor U8845 (N_8845,N_8568,N_8516);
nor U8846 (N_8846,N_8650,N_8647);
xor U8847 (N_8847,N_8581,N_8717);
xor U8848 (N_8848,N_8588,N_8736);
xnor U8849 (N_8849,N_8645,N_8660);
nor U8850 (N_8850,N_8634,N_8523);
nor U8851 (N_8851,N_8573,N_8739);
and U8852 (N_8852,N_8591,N_8533);
or U8853 (N_8853,N_8723,N_8590);
or U8854 (N_8854,N_8585,N_8557);
and U8855 (N_8855,N_8584,N_8599);
and U8856 (N_8856,N_8592,N_8649);
nor U8857 (N_8857,N_8553,N_8604);
nor U8858 (N_8858,N_8530,N_8699);
and U8859 (N_8859,N_8713,N_8500);
and U8860 (N_8860,N_8554,N_8566);
nand U8861 (N_8861,N_8624,N_8549);
or U8862 (N_8862,N_8517,N_8579);
xor U8863 (N_8863,N_8629,N_8617);
nand U8864 (N_8864,N_8672,N_8600);
xnor U8865 (N_8865,N_8743,N_8613);
xor U8866 (N_8866,N_8721,N_8609);
xnor U8867 (N_8867,N_8625,N_8552);
nand U8868 (N_8868,N_8726,N_8633);
or U8869 (N_8869,N_8727,N_8658);
or U8870 (N_8870,N_8700,N_8538);
xnor U8871 (N_8871,N_8732,N_8687);
xor U8872 (N_8872,N_8582,N_8620);
nand U8873 (N_8873,N_8548,N_8622);
xor U8874 (N_8874,N_8690,N_8640);
xnor U8875 (N_8875,N_8579,N_8654);
or U8876 (N_8876,N_8593,N_8509);
nor U8877 (N_8877,N_8721,N_8669);
or U8878 (N_8878,N_8521,N_8674);
nand U8879 (N_8879,N_8500,N_8617);
or U8880 (N_8880,N_8534,N_8723);
xnor U8881 (N_8881,N_8590,N_8732);
or U8882 (N_8882,N_8518,N_8676);
xor U8883 (N_8883,N_8621,N_8671);
nand U8884 (N_8884,N_8622,N_8700);
xnor U8885 (N_8885,N_8726,N_8542);
nand U8886 (N_8886,N_8520,N_8684);
xnor U8887 (N_8887,N_8501,N_8582);
or U8888 (N_8888,N_8574,N_8672);
nand U8889 (N_8889,N_8697,N_8514);
nand U8890 (N_8890,N_8623,N_8589);
and U8891 (N_8891,N_8688,N_8606);
nand U8892 (N_8892,N_8734,N_8638);
and U8893 (N_8893,N_8554,N_8623);
or U8894 (N_8894,N_8628,N_8616);
and U8895 (N_8895,N_8749,N_8699);
and U8896 (N_8896,N_8532,N_8643);
and U8897 (N_8897,N_8689,N_8631);
nor U8898 (N_8898,N_8732,N_8737);
xnor U8899 (N_8899,N_8633,N_8638);
and U8900 (N_8900,N_8535,N_8625);
nor U8901 (N_8901,N_8707,N_8597);
xor U8902 (N_8902,N_8547,N_8712);
xnor U8903 (N_8903,N_8705,N_8637);
nand U8904 (N_8904,N_8745,N_8606);
nand U8905 (N_8905,N_8740,N_8525);
nor U8906 (N_8906,N_8641,N_8592);
nor U8907 (N_8907,N_8541,N_8617);
and U8908 (N_8908,N_8694,N_8583);
xnor U8909 (N_8909,N_8506,N_8702);
nor U8910 (N_8910,N_8644,N_8532);
nor U8911 (N_8911,N_8575,N_8660);
nor U8912 (N_8912,N_8511,N_8662);
or U8913 (N_8913,N_8698,N_8544);
and U8914 (N_8914,N_8739,N_8731);
nor U8915 (N_8915,N_8503,N_8654);
nand U8916 (N_8916,N_8724,N_8558);
or U8917 (N_8917,N_8704,N_8678);
nor U8918 (N_8918,N_8579,N_8588);
nand U8919 (N_8919,N_8595,N_8599);
and U8920 (N_8920,N_8587,N_8665);
nand U8921 (N_8921,N_8608,N_8529);
xor U8922 (N_8922,N_8713,N_8550);
or U8923 (N_8923,N_8551,N_8546);
xnor U8924 (N_8924,N_8593,N_8609);
xnor U8925 (N_8925,N_8716,N_8649);
nor U8926 (N_8926,N_8597,N_8596);
or U8927 (N_8927,N_8698,N_8601);
nand U8928 (N_8928,N_8625,N_8514);
and U8929 (N_8929,N_8683,N_8671);
and U8930 (N_8930,N_8517,N_8574);
nor U8931 (N_8931,N_8526,N_8529);
and U8932 (N_8932,N_8692,N_8608);
or U8933 (N_8933,N_8748,N_8550);
nor U8934 (N_8934,N_8558,N_8537);
or U8935 (N_8935,N_8678,N_8520);
nor U8936 (N_8936,N_8734,N_8666);
xor U8937 (N_8937,N_8594,N_8550);
xor U8938 (N_8938,N_8713,N_8663);
or U8939 (N_8939,N_8672,N_8526);
nand U8940 (N_8940,N_8502,N_8501);
xor U8941 (N_8941,N_8602,N_8735);
xnor U8942 (N_8942,N_8632,N_8564);
nor U8943 (N_8943,N_8512,N_8566);
xor U8944 (N_8944,N_8617,N_8693);
nand U8945 (N_8945,N_8511,N_8676);
xor U8946 (N_8946,N_8601,N_8662);
nor U8947 (N_8947,N_8735,N_8696);
or U8948 (N_8948,N_8531,N_8518);
nor U8949 (N_8949,N_8693,N_8677);
or U8950 (N_8950,N_8587,N_8647);
xnor U8951 (N_8951,N_8544,N_8604);
nand U8952 (N_8952,N_8689,N_8704);
nor U8953 (N_8953,N_8538,N_8701);
nand U8954 (N_8954,N_8500,N_8506);
xor U8955 (N_8955,N_8639,N_8528);
nand U8956 (N_8956,N_8707,N_8720);
or U8957 (N_8957,N_8665,N_8551);
nor U8958 (N_8958,N_8539,N_8530);
and U8959 (N_8959,N_8723,N_8713);
or U8960 (N_8960,N_8711,N_8656);
or U8961 (N_8961,N_8680,N_8717);
xor U8962 (N_8962,N_8652,N_8641);
xnor U8963 (N_8963,N_8687,N_8698);
nor U8964 (N_8964,N_8552,N_8569);
or U8965 (N_8965,N_8527,N_8626);
and U8966 (N_8966,N_8640,N_8744);
nand U8967 (N_8967,N_8598,N_8653);
nand U8968 (N_8968,N_8509,N_8609);
and U8969 (N_8969,N_8602,N_8748);
xor U8970 (N_8970,N_8633,N_8692);
nor U8971 (N_8971,N_8655,N_8695);
and U8972 (N_8972,N_8671,N_8733);
xnor U8973 (N_8973,N_8509,N_8550);
or U8974 (N_8974,N_8672,N_8512);
and U8975 (N_8975,N_8587,N_8576);
xnor U8976 (N_8976,N_8727,N_8640);
and U8977 (N_8977,N_8508,N_8709);
nor U8978 (N_8978,N_8582,N_8694);
nand U8979 (N_8979,N_8667,N_8621);
or U8980 (N_8980,N_8655,N_8657);
or U8981 (N_8981,N_8636,N_8502);
nand U8982 (N_8982,N_8596,N_8729);
or U8983 (N_8983,N_8685,N_8601);
nor U8984 (N_8984,N_8524,N_8733);
nand U8985 (N_8985,N_8584,N_8524);
nor U8986 (N_8986,N_8709,N_8555);
or U8987 (N_8987,N_8509,N_8740);
nor U8988 (N_8988,N_8670,N_8700);
xor U8989 (N_8989,N_8562,N_8512);
nand U8990 (N_8990,N_8614,N_8651);
xnor U8991 (N_8991,N_8555,N_8702);
xnor U8992 (N_8992,N_8623,N_8596);
or U8993 (N_8993,N_8635,N_8627);
nor U8994 (N_8994,N_8614,N_8568);
nor U8995 (N_8995,N_8629,N_8726);
and U8996 (N_8996,N_8557,N_8595);
or U8997 (N_8997,N_8646,N_8717);
and U8998 (N_8998,N_8695,N_8631);
nor U8999 (N_8999,N_8576,N_8586);
or U9000 (N_9000,N_8930,N_8994);
nand U9001 (N_9001,N_8950,N_8821);
or U9002 (N_9002,N_8845,N_8935);
nand U9003 (N_9003,N_8823,N_8954);
nor U9004 (N_9004,N_8805,N_8840);
and U9005 (N_9005,N_8989,N_8797);
nor U9006 (N_9006,N_8960,N_8892);
nor U9007 (N_9007,N_8976,N_8906);
nor U9008 (N_9008,N_8854,N_8880);
and U9009 (N_9009,N_8763,N_8876);
xnor U9010 (N_9010,N_8977,N_8924);
nor U9011 (N_9011,N_8953,N_8990);
or U9012 (N_9012,N_8865,N_8882);
xor U9013 (N_9013,N_8921,N_8828);
nand U9014 (N_9014,N_8959,N_8972);
or U9015 (N_9015,N_8804,N_8956);
xor U9016 (N_9016,N_8957,N_8941);
and U9017 (N_9017,N_8914,N_8759);
and U9018 (N_9018,N_8864,N_8982);
and U9019 (N_9019,N_8755,N_8827);
or U9020 (N_9020,N_8775,N_8904);
xnor U9021 (N_9021,N_8800,N_8975);
or U9022 (N_9022,N_8971,N_8945);
nand U9023 (N_9023,N_8838,N_8907);
or U9024 (N_9024,N_8753,N_8936);
or U9025 (N_9025,N_8983,N_8781);
nor U9026 (N_9026,N_8862,N_8872);
or U9027 (N_9027,N_8911,N_8883);
nor U9028 (N_9028,N_8861,N_8832);
and U9029 (N_9029,N_8961,N_8929);
xor U9030 (N_9030,N_8813,N_8810);
xor U9031 (N_9031,N_8939,N_8844);
xnor U9032 (N_9032,N_8942,N_8839);
xor U9033 (N_9033,N_8836,N_8875);
nand U9034 (N_9034,N_8870,N_8949);
and U9035 (N_9035,N_8760,N_8984);
xnor U9036 (N_9036,N_8969,N_8850);
nand U9037 (N_9037,N_8996,N_8997);
or U9038 (N_9038,N_8947,N_8770);
and U9039 (N_9039,N_8852,N_8963);
xnor U9040 (N_9040,N_8894,N_8807);
nand U9041 (N_9041,N_8931,N_8798);
or U9042 (N_9042,N_8768,N_8979);
nand U9043 (N_9043,N_8974,N_8999);
xor U9044 (N_9044,N_8968,N_8920);
nand U9045 (N_9045,N_8783,N_8928);
nand U9046 (N_9046,N_8913,N_8857);
nand U9047 (N_9047,N_8750,N_8767);
xnor U9048 (N_9048,N_8752,N_8884);
nor U9049 (N_9049,N_8843,N_8816);
nor U9050 (N_9050,N_8833,N_8849);
xor U9051 (N_9051,N_8866,N_8938);
nor U9052 (N_9052,N_8903,N_8937);
nor U9053 (N_9053,N_8815,N_8782);
and U9054 (N_9054,N_8902,N_8881);
and U9055 (N_9055,N_8991,N_8985);
nand U9056 (N_9056,N_8958,N_8898);
nand U9057 (N_9057,N_8812,N_8764);
and U9058 (N_9058,N_8923,N_8784);
nor U9059 (N_9059,N_8918,N_8809);
nor U9060 (N_9060,N_8793,N_8966);
or U9061 (N_9061,N_8915,N_8889);
or U9062 (N_9062,N_8774,N_8912);
or U9063 (N_9063,N_8825,N_8905);
or U9064 (N_9064,N_8869,N_8758);
nand U9065 (N_9065,N_8826,N_8834);
or U9066 (N_9066,N_8967,N_8873);
nand U9067 (N_9067,N_8830,N_8853);
nand U9068 (N_9068,N_8796,N_8814);
and U9069 (N_9069,N_8871,N_8818);
xor U9070 (N_9070,N_8980,N_8932);
xnor U9071 (N_9071,N_8856,N_8841);
and U9072 (N_9072,N_8788,N_8981);
xnor U9073 (N_9073,N_8791,N_8754);
or U9074 (N_9074,N_8820,N_8801);
nand U9075 (N_9075,N_8792,N_8926);
nand U9076 (N_9076,N_8837,N_8842);
nor U9077 (N_9077,N_8891,N_8851);
nand U9078 (N_9078,N_8927,N_8925);
nand U9079 (N_9079,N_8806,N_8900);
nand U9080 (N_9080,N_8785,N_8822);
nand U9081 (N_9081,N_8934,N_8799);
nand U9082 (N_9082,N_8794,N_8893);
nor U9083 (N_9083,N_8772,N_8895);
or U9084 (N_9084,N_8751,N_8786);
xnor U9085 (N_9085,N_8878,N_8901);
or U9086 (N_9086,N_8922,N_8847);
nand U9087 (N_9087,N_8917,N_8916);
nand U9088 (N_9088,N_8993,N_8855);
xor U9089 (N_9089,N_8859,N_8773);
or U9090 (N_9090,N_8899,N_8987);
xor U9091 (N_9091,N_8795,N_8766);
nand U9092 (N_9092,N_8973,N_8765);
nor U9093 (N_9093,N_8896,N_8831);
nor U9094 (N_9094,N_8874,N_8777);
nand U9095 (N_9095,N_8860,N_8819);
and U9096 (N_9096,N_8919,N_8867);
xor U9097 (N_9097,N_8978,N_8848);
and U9098 (N_9098,N_8756,N_8944);
xnor U9099 (N_9099,N_8955,N_8965);
nor U9100 (N_9100,N_8824,N_8962);
or U9101 (N_9101,N_8811,N_8803);
or U9102 (N_9102,N_8877,N_8780);
or U9103 (N_9103,N_8890,N_8808);
xor U9104 (N_9104,N_8943,N_8886);
or U9105 (N_9105,N_8789,N_8771);
nand U9106 (N_9106,N_8817,N_8802);
and U9107 (N_9107,N_8908,N_8995);
xor U9108 (N_9108,N_8779,N_8946);
or U9109 (N_9109,N_8952,N_8879);
and U9110 (N_9110,N_8885,N_8868);
xor U9111 (N_9111,N_8863,N_8762);
xor U9112 (N_9112,N_8988,N_8888);
xnor U9113 (N_9113,N_8769,N_8846);
nand U9114 (N_9114,N_8790,N_8829);
or U9115 (N_9115,N_8778,N_8761);
xor U9116 (N_9116,N_8970,N_8897);
and U9117 (N_9117,N_8998,N_8964);
or U9118 (N_9118,N_8933,N_8787);
or U9119 (N_9119,N_8948,N_8835);
nand U9120 (N_9120,N_8992,N_8940);
and U9121 (N_9121,N_8910,N_8951);
or U9122 (N_9122,N_8858,N_8986);
and U9123 (N_9123,N_8887,N_8757);
xor U9124 (N_9124,N_8909,N_8776);
nand U9125 (N_9125,N_8780,N_8888);
and U9126 (N_9126,N_8963,N_8895);
or U9127 (N_9127,N_8780,N_8795);
or U9128 (N_9128,N_8886,N_8996);
nand U9129 (N_9129,N_8825,N_8967);
xor U9130 (N_9130,N_8951,N_8776);
nand U9131 (N_9131,N_8774,N_8893);
or U9132 (N_9132,N_8898,N_8863);
and U9133 (N_9133,N_8915,N_8855);
and U9134 (N_9134,N_8781,N_8783);
nor U9135 (N_9135,N_8780,N_8926);
or U9136 (N_9136,N_8963,N_8986);
xor U9137 (N_9137,N_8974,N_8903);
nand U9138 (N_9138,N_8798,N_8796);
nor U9139 (N_9139,N_8916,N_8883);
nor U9140 (N_9140,N_8995,N_8952);
and U9141 (N_9141,N_8768,N_8945);
xnor U9142 (N_9142,N_8923,N_8758);
or U9143 (N_9143,N_8791,N_8985);
nand U9144 (N_9144,N_8939,N_8836);
xnor U9145 (N_9145,N_8944,N_8984);
nor U9146 (N_9146,N_8837,N_8861);
nor U9147 (N_9147,N_8893,N_8797);
nor U9148 (N_9148,N_8825,N_8783);
xnor U9149 (N_9149,N_8998,N_8896);
nand U9150 (N_9150,N_8823,N_8965);
xnor U9151 (N_9151,N_8963,N_8752);
and U9152 (N_9152,N_8941,N_8969);
and U9153 (N_9153,N_8756,N_8793);
or U9154 (N_9154,N_8797,N_8943);
nand U9155 (N_9155,N_8896,N_8786);
or U9156 (N_9156,N_8801,N_8935);
xnor U9157 (N_9157,N_8924,N_8925);
and U9158 (N_9158,N_8835,N_8863);
nand U9159 (N_9159,N_8780,N_8800);
and U9160 (N_9160,N_8860,N_8924);
xnor U9161 (N_9161,N_8902,N_8982);
and U9162 (N_9162,N_8916,N_8980);
or U9163 (N_9163,N_8909,N_8993);
nand U9164 (N_9164,N_8832,N_8877);
nor U9165 (N_9165,N_8840,N_8998);
and U9166 (N_9166,N_8853,N_8951);
and U9167 (N_9167,N_8799,N_8914);
and U9168 (N_9168,N_8762,N_8900);
nand U9169 (N_9169,N_8762,N_8766);
nand U9170 (N_9170,N_8998,N_8933);
and U9171 (N_9171,N_8959,N_8793);
xnor U9172 (N_9172,N_8783,N_8977);
nand U9173 (N_9173,N_8842,N_8828);
nor U9174 (N_9174,N_8862,N_8784);
nand U9175 (N_9175,N_8769,N_8758);
and U9176 (N_9176,N_8828,N_8762);
and U9177 (N_9177,N_8990,N_8955);
and U9178 (N_9178,N_8770,N_8956);
or U9179 (N_9179,N_8820,N_8960);
or U9180 (N_9180,N_8901,N_8896);
nand U9181 (N_9181,N_8827,N_8907);
nor U9182 (N_9182,N_8851,N_8752);
or U9183 (N_9183,N_8993,N_8754);
or U9184 (N_9184,N_8825,N_8764);
or U9185 (N_9185,N_8975,N_8919);
and U9186 (N_9186,N_8978,N_8855);
xnor U9187 (N_9187,N_8856,N_8796);
and U9188 (N_9188,N_8916,N_8902);
nand U9189 (N_9189,N_8868,N_8963);
and U9190 (N_9190,N_8752,N_8750);
and U9191 (N_9191,N_8801,N_8872);
xnor U9192 (N_9192,N_8891,N_8952);
and U9193 (N_9193,N_8863,N_8899);
nor U9194 (N_9194,N_8857,N_8882);
nor U9195 (N_9195,N_8994,N_8979);
xor U9196 (N_9196,N_8859,N_8871);
xnor U9197 (N_9197,N_8950,N_8777);
and U9198 (N_9198,N_8965,N_8960);
and U9199 (N_9199,N_8921,N_8773);
nand U9200 (N_9200,N_8805,N_8834);
nor U9201 (N_9201,N_8921,N_8780);
nand U9202 (N_9202,N_8844,N_8881);
or U9203 (N_9203,N_8886,N_8948);
nor U9204 (N_9204,N_8817,N_8857);
nor U9205 (N_9205,N_8854,N_8945);
or U9206 (N_9206,N_8794,N_8945);
and U9207 (N_9207,N_8916,N_8855);
nor U9208 (N_9208,N_8895,N_8791);
xor U9209 (N_9209,N_8912,N_8901);
and U9210 (N_9210,N_8971,N_8835);
nand U9211 (N_9211,N_8913,N_8887);
xnor U9212 (N_9212,N_8968,N_8980);
nand U9213 (N_9213,N_8795,N_8797);
or U9214 (N_9214,N_8887,N_8958);
nor U9215 (N_9215,N_8930,N_8751);
or U9216 (N_9216,N_8968,N_8801);
or U9217 (N_9217,N_8981,N_8842);
xor U9218 (N_9218,N_8835,N_8775);
nor U9219 (N_9219,N_8778,N_8858);
xor U9220 (N_9220,N_8958,N_8939);
xnor U9221 (N_9221,N_8796,N_8809);
or U9222 (N_9222,N_8899,N_8976);
nor U9223 (N_9223,N_8983,N_8868);
nor U9224 (N_9224,N_8877,N_8923);
xnor U9225 (N_9225,N_8807,N_8831);
or U9226 (N_9226,N_8791,N_8908);
nand U9227 (N_9227,N_8947,N_8763);
xnor U9228 (N_9228,N_8929,N_8936);
nor U9229 (N_9229,N_8909,N_8923);
nand U9230 (N_9230,N_8773,N_8904);
xnor U9231 (N_9231,N_8847,N_8894);
and U9232 (N_9232,N_8939,N_8877);
nor U9233 (N_9233,N_8916,N_8904);
and U9234 (N_9234,N_8998,N_8893);
nand U9235 (N_9235,N_8863,N_8827);
nor U9236 (N_9236,N_8964,N_8961);
xnor U9237 (N_9237,N_8882,N_8778);
xnor U9238 (N_9238,N_8890,N_8920);
or U9239 (N_9239,N_8899,N_8769);
and U9240 (N_9240,N_8979,N_8810);
nand U9241 (N_9241,N_8771,N_8752);
nor U9242 (N_9242,N_8892,N_8757);
xor U9243 (N_9243,N_8897,N_8787);
nand U9244 (N_9244,N_8958,N_8991);
or U9245 (N_9245,N_8863,N_8959);
nand U9246 (N_9246,N_8925,N_8803);
and U9247 (N_9247,N_8769,N_8771);
or U9248 (N_9248,N_8916,N_8919);
nand U9249 (N_9249,N_8788,N_8772);
nand U9250 (N_9250,N_9217,N_9098);
nor U9251 (N_9251,N_9172,N_9035);
xor U9252 (N_9252,N_9016,N_9184);
or U9253 (N_9253,N_9227,N_9128);
and U9254 (N_9254,N_9198,N_9244);
and U9255 (N_9255,N_9183,N_9045);
or U9256 (N_9256,N_9024,N_9041);
xnor U9257 (N_9257,N_9054,N_9179);
and U9258 (N_9258,N_9146,N_9211);
nand U9259 (N_9259,N_9019,N_9004);
and U9260 (N_9260,N_9005,N_9206);
nor U9261 (N_9261,N_9010,N_9207);
nor U9262 (N_9262,N_9104,N_9247);
nand U9263 (N_9263,N_9190,N_9007);
xnor U9264 (N_9264,N_9018,N_9163);
or U9265 (N_9265,N_9075,N_9080);
nor U9266 (N_9266,N_9222,N_9088);
nor U9267 (N_9267,N_9173,N_9218);
xor U9268 (N_9268,N_9047,N_9021);
and U9269 (N_9269,N_9103,N_9000);
xor U9270 (N_9270,N_9236,N_9029);
xor U9271 (N_9271,N_9090,N_9112);
and U9272 (N_9272,N_9028,N_9056);
nand U9273 (N_9273,N_9052,N_9081);
nor U9274 (N_9274,N_9209,N_9229);
xor U9275 (N_9275,N_9203,N_9109);
xnor U9276 (N_9276,N_9065,N_9210);
and U9277 (N_9277,N_9117,N_9133);
xnor U9278 (N_9278,N_9115,N_9219);
nand U9279 (N_9279,N_9138,N_9027);
xor U9280 (N_9280,N_9061,N_9097);
or U9281 (N_9281,N_9102,N_9144);
and U9282 (N_9282,N_9132,N_9046);
nand U9283 (N_9283,N_9188,N_9225);
and U9284 (N_9284,N_9038,N_9053);
xor U9285 (N_9285,N_9074,N_9023);
xor U9286 (N_9286,N_9230,N_9226);
nor U9287 (N_9287,N_9240,N_9224);
xnor U9288 (N_9288,N_9161,N_9170);
xor U9289 (N_9289,N_9189,N_9212);
xnor U9290 (N_9290,N_9011,N_9214);
nand U9291 (N_9291,N_9122,N_9145);
or U9292 (N_9292,N_9022,N_9095);
nand U9293 (N_9293,N_9114,N_9020);
nand U9294 (N_9294,N_9037,N_9237);
nor U9295 (N_9295,N_9082,N_9094);
or U9296 (N_9296,N_9157,N_9185);
nand U9297 (N_9297,N_9208,N_9153);
nor U9298 (N_9298,N_9249,N_9036);
or U9299 (N_9299,N_9195,N_9130);
xor U9300 (N_9300,N_9014,N_9213);
nor U9301 (N_9301,N_9160,N_9220);
nand U9302 (N_9302,N_9026,N_9239);
nand U9303 (N_9303,N_9142,N_9223);
or U9304 (N_9304,N_9033,N_9025);
nor U9305 (N_9305,N_9246,N_9121);
and U9306 (N_9306,N_9205,N_9241);
and U9307 (N_9307,N_9156,N_9136);
and U9308 (N_9308,N_9200,N_9048);
and U9309 (N_9309,N_9221,N_9155);
nand U9310 (N_9310,N_9069,N_9238);
xnor U9311 (N_9311,N_9182,N_9072);
nand U9312 (N_9312,N_9196,N_9140);
xnor U9313 (N_9313,N_9042,N_9154);
xnor U9314 (N_9314,N_9086,N_9181);
xor U9315 (N_9315,N_9168,N_9034);
or U9316 (N_9316,N_9204,N_9079);
xor U9317 (N_9317,N_9076,N_9191);
nand U9318 (N_9318,N_9158,N_9091);
nand U9319 (N_9319,N_9044,N_9073);
nor U9320 (N_9320,N_9127,N_9177);
nand U9321 (N_9321,N_9137,N_9039);
nand U9322 (N_9322,N_9233,N_9078);
and U9323 (N_9323,N_9167,N_9118);
nor U9324 (N_9324,N_9031,N_9101);
xnor U9325 (N_9325,N_9096,N_9231);
xnor U9326 (N_9326,N_9180,N_9099);
and U9327 (N_9327,N_9120,N_9067);
nand U9328 (N_9328,N_9192,N_9202);
and U9329 (N_9329,N_9009,N_9171);
xor U9330 (N_9330,N_9070,N_9235);
xor U9331 (N_9331,N_9123,N_9175);
xor U9332 (N_9332,N_9057,N_9068);
nand U9333 (N_9333,N_9150,N_9242);
and U9334 (N_9334,N_9148,N_9124);
or U9335 (N_9335,N_9113,N_9234);
xor U9336 (N_9336,N_9201,N_9092);
or U9337 (N_9337,N_9077,N_9126);
and U9338 (N_9338,N_9194,N_9060);
or U9339 (N_9339,N_9129,N_9216);
nor U9340 (N_9340,N_9131,N_9110);
and U9341 (N_9341,N_9051,N_9066);
or U9342 (N_9342,N_9165,N_9166);
and U9343 (N_9343,N_9050,N_9199);
nor U9344 (N_9344,N_9119,N_9186);
nand U9345 (N_9345,N_9087,N_9063);
or U9346 (N_9346,N_9149,N_9107);
nand U9347 (N_9347,N_9002,N_9159);
xor U9348 (N_9348,N_9135,N_9058);
nor U9349 (N_9349,N_9169,N_9108);
xnor U9350 (N_9350,N_9100,N_9049);
or U9351 (N_9351,N_9105,N_9071);
xor U9352 (N_9352,N_9125,N_9012);
nor U9353 (N_9353,N_9040,N_9083);
nor U9354 (N_9354,N_9228,N_9187);
xor U9355 (N_9355,N_9008,N_9151);
xor U9356 (N_9356,N_9085,N_9141);
nor U9357 (N_9357,N_9043,N_9059);
and U9358 (N_9358,N_9084,N_9116);
nor U9359 (N_9359,N_9062,N_9197);
nand U9360 (N_9360,N_9001,N_9015);
nand U9361 (N_9361,N_9174,N_9193);
and U9362 (N_9362,N_9176,N_9017);
or U9363 (N_9363,N_9147,N_9055);
and U9364 (N_9364,N_9248,N_9106);
nand U9365 (N_9365,N_9162,N_9089);
nor U9366 (N_9366,N_9003,N_9143);
nand U9367 (N_9367,N_9064,N_9030);
xnor U9368 (N_9368,N_9093,N_9013);
or U9369 (N_9369,N_9245,N_9111);
nand U9370 (N_9370,N_9243,N_9164);
nand U9371 (N_9371,N_9232,N_9152);
or U9372 (N_9372,N_9006,N_9134);
xor U9373 (N_9373,N_9139,N_9215);
xnor U9374 (N_9374,N_9178,N_9032);
and U9375 (N_9375,N_9175,N_9195);
or U9376 (N_9376,N_9016,N_9027);
nor U9377 (N_9377,N_9030,N_9180);
and U9378 (N_9378,N_9178,N_9096);
and U9379 (N_9379,N_9219,N_9104);
and U9380 (N_9380,N_9168,N_9187);
or U9381 (N_9381,N_9019,N_9132);
or U9382 (N_9382,N_9085,N_9025);
and U9383 (N_9383,N_9017,N_9226);
xor U9384 (N_9384,N_9184,N_9234);
and U9385 (N_9385,N_9180,N_9185);
or U9386 (N_9386,N_9162,N_9017);
nor U9387 (N_9387,N_9220,N_9198);
xor U9388 (N_9388,N_9237,N_9246);
nor U9389 (N_9389,N_9048,N_9083);
or U9390 (N_9390,N_9202,N_9015);
nor U9391 (N_9391,N_9028,N_9200);
and U9392 (N_9392,N_9052,N_9011);
or U9393 (N_9393,N_9184,N_9195);
nor U9394 (N_9394,N_9008,N_9084);
xnor U9395 (N_9395,N_9032,N_9048);
nor U9396 (N_9396,N_9223,N_9048);
nor U9397 (N_9397,N_9073,N_9088);
xor U9398 (N_9398,N_9117,N_9181);
nand U9399 (N_9399,N_9125,N_9141);
and U9400 (N_9400,N_9245,N_9099);
nand U9401 (N_9401,N_9107,N_9227);
nor U9402 (N_9402,N_9173,N_9058);
or U9403 (N_9403,N_9180,N_9199);
nand U9404 (N_9404,N_9235,N_9011);
nand U9405 (N_9405,N_9183,N_9153);
nor U9406 (N_9406,N_9187,N_9227);
xnor U9407 (N_9407,N_9218,N_9001);
xnor U9408 (N_9408,N_9091,N_9184);
and U9409 (N_9409,N_9033,N_9101);
xnor U9410 (N_9410,N_9208,N_9119);
or U9411 (N_9411,N_9095,N_9077);
or U9412 (N_9412,N_9049,N_9198);
or U9413 (N_9413,N_9200,N_9166);
xnor U9414 (N_9414,N_9206,N_9059);
nand U9415 (N_9415,N_9023,N_9060);
nor U9416 (N_9416,N_9139,N_9054);
nor U9417 (N_9417,N_9222,N_9048);
xor U9418 (N_9418,N_9108,N_9161);
or U9419 (N_9419,N_9168,N_9060);
or U9420 (N_9420,N_9047,N_9066);
and U9421 (N_9421,N_9100,N_9195);
xnor U9422 (N_9422,N_9017,N_9127);
nand U9423 (N_9423,N_9234,N_9157);
and U9424 (N_9424,N_9227,N_9136);
or U9425 (N_9425,N_9162,N_9026);
xnor U9426 (N_9426,N_9102,N_9081);
nand U9427 (N_9427,N_9162,N_9139);
and U9428 (N_9428,N_9170,N_9049);
and U9429 (N_9429,N_9115,N_9059);
nand U9430 (N_9430,N_9062,N_9188);
or U9431 (N_9431,N_9105,N_9099);
and U9432 (N_9432,N_9066,N_9168);
nor U9433 (N_9433,N_9202,N_9165);
nor U9434 (N_9434,N_9003,N_9051);
and U9435 (N_9435,N_9196,N_9070);
nand U9436 (N_9436,N_9226,N_9196);
nand U9437 (N_9437,N_9214,N_9098);
nand U9438 (N_9438,N_9237,N_9192);
nand U9439 (N_9439,N_9000,N_9099);
xnor U9440 (N_9440,N_9210,N_9134);
xor U9441 (N_9441,N_9184,N_9192);
nor U9442 (N_9442,N_9188,N_9056);
or U9443 (N_9443,N_9064,N_9063);
xnor U9444 (N_9444,N_9101,N_9074);
xor U9445 (N_9445,N_9128,N_9202);
xnor U9446 (N_9446,N_9039,N_9101);
nor U9447 (N_9447,N_9249,N_9093);
nand U9448 (N_9448,N_9096,N_9134);
or U9449 (N_9449,N_9033,N_9201);
or U9450 (N_9450,N_9130,N_9104);
nor U9451 (N_9451,N_9180,N_9214);
or U9452 (N_9452,N_9111,N_9109);
nor U9453 (N_9453,N_9028,N_9089);
and U9454 (N_9454,N_9018,N_9244);
or U9455 (N_9455,N_9186,N_9076);
nand U9456 (N_9456,N_9047,N_9092);
xnor U9457 (N_9457,N_9165,N_9057);
nor U9458 (N_9458,N_9231,N_9152);
xor U9459 (N_9459,N_9204,N_9033);
or U9460 (N_9460,N_9110,N_9038);
nor U9461 (N_9461,N_9178,N_9196);
xnor U9462 (N_9462,N_9181,N_9091);
or U9463 (N_9463,N_9249,N_9174);
or U9464 (N_9464,N_9040,N_9110);
xor U9465 (N_9465,N_9210,N_9129);
nand U9466 (N_9466,N_9222,N_9046);
nand U9467 (N_9467,N_9218,N_9174);
and U9468 (N_9468,N_9054,N_9154);
and U9469 (N_9469,N_9154,N_9224);
xnor U9470 (N_9470,N_9033,N_9245);
or U9471 (N_9471,N_9117,N_9147);
or U9472 (N_9472,N_9241,N_9245);
xor U9473 (N_9473,N_9140,N_9039);
nor U9474 (N_9474,N_9159,N_9065);
nor U9475 (N_9475,N_9153,N_9237);
nand U9476 (N_9476,N_9114,N_9187);
nor U9477 (N_9477,N_9230,N_9161);
nor U9478 (N_9478,N_9053,N_9173);
nand U9479 (N_9479,N_9082,N_9194);
and U9480 (N_9480,N_9159,N_9168);
xor U9481 (N_9481,N_9178,N_9018);
or U9482 (N_9482,N_9090,N_9085);
nand U9483 (N_9483,N_9117,N_9151);
and U9484 (N_9484,N_9225,N_9194);
nor U9485 (N_9485,N_9142,N_9071);
nor U9486 (N_9486,N_9059,N_9133);
and U9487 (N_9487,N_9050,N_9083);
nand U9488 (N_9488,N_9143,N_9203);
xor U9489 (N_9489,N_9151,N_9245);
nor U9490 (N_9490,N_9068,N_9110);
nand U9491 (N_9491,N_9021,N_9046);
nor U9492 (N_9492,N_9108,N_9114);
or U9493 (N_9493,N_9098,N_9055);
nand U9494 (N_9494,N_9119,N_9086);
xor U9495 (N_9495,N_9141,N_9154);
and U9496 (N_9496,N_9040,N_9154);
nor U9497 (N_9497,N_9089,N_9246);
and U9498 (N_9498,N_9014,N_9106);
or U9499 (N_9499,N_9042,N_9209);
and U9500 (N_9500,N_9267,N_9347);
nor U9501 (N_9501,N_9300,N_9315);
nand U9502 (N_9502,N_9454,N_9406);
and U9503 (N_9503,N_9327,N_9426);
nor U9504 (N_9504,N_9298,N_9316);
xor U9505 (N_9505,N_9464,N_9466);
nand U9506 (N_9506,N_9254,N_9442);
nor U9507 (N_9507,N_9287,N_9306);
xnor U9508 (N_9508,N_9278,N_9284);
and U9509 (N_9509,N_9294,N_9429);
xnor U9510 (N_9510,N_9331,N_9388);
and U9511 (N_9511,N_9394,N_9486);
or U9512 (N_9512,N_9310,N_9261);
or U9513 (N_9513,N_9418,N_9414);
xor U9514 (N_9514,N_9283,N_9461);
nand U9515 (N_9515,N_9422,N_9367);
and U9516 (N_9516,N_9373,N_9441);
and U9517 (N_9517,N_9258,N_9489);
or U9518 (N_9518,N_9274,N_9385);
or U9519 (N_9519,N_9391,N_9271);
or U9520 (N_9520,N_9337,N_9308);
or U9521 (N_9521,N_9400,N_9313);
nor U9522 (N_9522,N_9380,N_9393);
nand U9523 (N_9523,N_9288,N_9372);
nand U9524 (N_9524,N_9481,N_9438);
and U9525 (N_9525,N_9496,N_9265);
nor U9526 (N_9526,N_9378,N_9477);
and U9527 (N_9527,N_9399,N_9455);
xor U9528 (N_9528,N_9324,N_9450);
xnor U9529 (N_9529,N_9432,N_9362);
and U9530 (N_9530,N_9404,N_9302);
and U9531 (N_9531,N_9390,N_9498);
or U9532 (N_9532,N_9431,N_9439);
nor U9533 (N_9533,N_9251,N_9350);
nor U9534 (N_9534,N_9255,N_9451);
and U9535 (N_9535,N_9387,N_9475);
xor U9536 (N_9536,N_9275,N_9412);
nor U9537 (N_9537,N_9428,N_9482);
nor U9538 (N_9538,N_9370,N_9292);
or U9539 (N_9539,N_9334,N_9289);
xnor U9540 (N_9540,N_9460,N_9487);
or U9541 (N_9541,N_9329,N_9479);
or U9542 (N_9542,N_9382,N_9330);
and U9543 (N_9543,N_9250,N_9325);
xor U9544 (N_9544,N_9398,N_9446);
nand U9545 (N_9545,N_9447,N_9457);
and U9546 (N_9546,N_9467,N_9342);
and U9547 (N_9547,N_9354,N_9358);
nor U9548 (N_9548,N_9369,N_9341);
nor U9549 (N_9549,N_9279,N_9491);
nand U9550 (N_9550,N_9492,N_9345);
or U9551 (N_9551,N_9305,N_9304);
or U9552 (N_9552,N_9332,N_9335);
nand U9553 (N_9553,N_9386,N_9407);
nor U9554 (N_9554,N_9485,N_9408);
and U9555 (N_9555,N_9360,N_9262);
xor U9556 (N_9556,N_9290,N_9417);
and U9557 (N_9557,N_9413,N_9272);
xor U9558 (N_9558,N_9469,N_9449);
nand U9559 (N_9559,N_9493,N_9352);
nor U9560 (N_9560,N_9495,N_9427);
nand U9561 (N_9561,N_9395,N_9420);
xor U9562 (N_9562,N_9494,N_9276);
or U9563 (N_9563,N_9397,N_9319);
nor U9564 (N_9564,N_9293,N_9269);
and U9565 (N_9565,N_9266,N_9452);
or U9566 (N_9566,N_9340,N_9356);
nand U9567 (N_9567,N_9314,N_9322);
and U9568 (N_9568,N_9389,N_9480);
nor U9569 (N_9569,N_9458,N_9366);
or U9570 (N_9570,N_9383,N_9415);
nor U9571 (N_9571,N_9270,N_9476);
nand U9572 (N_9572,N_9472,N_9361);
or U9573 (N_9573,N_9423,N_9291);
or U9574 (N_9574,N_9473,N_9484);
or U9575 (N_9575,N_9280,N_9321);
or U9576 (N_9576,N_9421,N_9277);
and U9577 (N_9577,N_9435,N_9375);
nor U9578 (N_9578,N_9433,N_9497);
and U9579 (N_9579,N_9470,N_9499);
nor U9580 (N_9580,N_9405,N_9410);
nand U9581 (N_9581,N_9465,N_9301);
or U9582 (N_9582,N_9323,N_9403);
xnor U9583 (N_9583,N_9328,N_9474);
and U9584 (N_9584,N_9320,N_9309);
and U9585 (N_9585,N_9368,N_9462);
or U9586 (N_9586,N_9411,N_9295);
xnor U9587 (N_9587,N_9379,N_9351);
nand U9588 (N_9588,N_9416,N_9299);
or U9589 (N_9589,N_9285,N_9263);
nand U9590 (N_9590,N_9338,N_9456);
and U9591 (N_9591,N_9376,N_9318);
nor U9592 (N_9592,N_9443,N_9448);
or U9593 (N_9593,N_9268,N_9381);
or U9594 (N_9594,N_9374,N_9333);
xor U9595 (N_9595,N_9286,N_9483);
or U9596 (N_9596,N_9281,N_9359);
and U9597 (N_9597,N_9257,N_9478);
xnor U9598 (N_9598,N_9419,N_9409);
nor U9599 (N_9599,N_9311,N_9307);
and U9600 (N_9600,N_9363,N_9273);
and U9601 (N_9601,N_9471,N_9396);
xnor U9602 (N_9602,N_9326,N_9440);
and U9603 (N_9603,N_9459,N_9430);
nor U9604 (N_9604,N_9364,N_9444);
or U9605 (N_9605,N_9346,N_9317);
and U9606 (N_9606,N_9348,N_9425);
or U9607 (N_9607,N_9463,N_9377);
or U9608 (N_9608,N_9424,N_9392);
nor U9609 (N_9609,N_9353,N_9445);
and U9610 (N_9610,N_9488,N_9264);
nand U9611 (N_9611,N_9384,N_9339);
nand U9612 (N_9612,N_9490,N_9312);
nand U9613 (N_9613,N_9252,N_9401);
xnor U9614 (N_9614,N_9365,N_9343);
xor U9615 (N_9615,N_9256,N_9349);
nand U9616 (N_9616,N_9296,N_9253);
xor U9617 (N_9617,N_9436,N_9336);
nor U9618 (N_9618,N_9344,N_9453);
and U9619 (N_9619,N_9303,N_9371);
nor U9620 (N_9620,N_9260,N_9357);
or U9621 (N_9621,N_9437,N_9402);
or U9622 (N_9622,N_9259,N_9434);
nand U9623 (N_9623,N_9297,N_9282);
or U9624 (N_9624,N_9468,N_9355);
or U9625 (N_9625,N_9287,N_9439);
xnor U9626 (N_9626,N_9463,N_9403);
and U9627 (N_9627,N_9497,N_9421);
or U9628 (N_9628,N_9328,N_9319);
xor U9629 (N_9629,N_9291,N_9432);
and U9630 (N_9630,N_9252,N_9467);
xor U9631 (N_9631,N_9457,N_9357);
xnor U9632 (N_9632,N_9371,N_9391);
nor U9633 (N_9633,N_9400,N_9357);
nor U9634 (N_9634,N_9468,N_9269);
nand U9635 (N_9635,N_9456,N_9434);
nor U9636 (N_9636,N_9320,N_9254);
or U9637 (N_9637,N_9321,N_9371);
and U9638 (N_9638,N_9347,N_9436);
xor U9639 (N_9639,N_9364,N_9345);
nand U9640 (N_9640,N_9436,N_9458);
and U9641 (N_9641,N_9449,N_9497);
or U9642 (N_9642,N_9426,N_9473);
nor U9643 (N_9643,N_9290,N_9382);
or U9644 (N_9644,N_9270,N_9281);
nor U9645 (N_9645,N_9360,N_9425);
xnor U9646 (N_9646,N_9285,N_9489);
or U9647 (N_9647,N_9384,N_9393);
nand U9648 (N_9648,N_9449,N_9415);
nor U9649 (N_9649,N_9265,N_9361);
nor U9650 (N_9650,N_9472,N_9409);
xor U9651 (N_9651,N_9356,N_9386);
or U9652 (N_9652,N_9295,N_9499);
nand U9653 (N_9653,N_9415,N_9283);
xor U9654 (N_9654,N_9337,N_9360);
nor U9655 (N_9655,N_9456,N_9496);
or U9656 (N_9656,N_9418,N_9387);
and U9657 (N_9657,N_9358,N_9465);
nor U9658 (N_9658,N_9459,N_9355);
and U9659 (N_9659,N_9494,N_9417);
nand U9660 (N_9660,N_9384,N_9268);
or U9661 (N_9661,N_9304,N_9427);
nand U9662 (N_9662,N_9258,N_9291);
xnor U9663 (N_9663,N_9498,N_9313);
xnor U9664 (N_9664,N_9427,N_9361);
and U9665 (N_9665,N_9273,N_9476);
and U9666 (N_9666,N_9488,N_9252);
or U9667 (N_9667,N_9472,N_9391);
nand U9668 (N_9668,N_9459,N_9299);
nand U9669 (N_9669,N_9301,N_9289);
and U9670 (N_9670,N_9329,N_9411);
xor U9671 (N_9671,N_9422,N_9411);
and U9672 (N_9672,N_9393,N_9449);
xor U9673 (N_9673,N_9448,N_9254);
nand U9674 (N_9674,N_9478,N_9400);
nand U9675 (N_9675,N_9402,N_9279);
nand U9676 (N_9676,N_9489,N_9358);
xor U9677 (N_9677,N_9462,N_9478);
or U9678 (N_9678,N_9327,N_9421);
nand U9679 (N_9679,N_9485,N_9279);
or U9680 (N_9680,N_9255,N_9479);
xnor U9681 (N_9681,N_9373,N_9350);
or U9682 (N_9682,N_9424,N_9404);
xnor U9683 (N_9683,N_9254,N_9421);
and U9684 (N_9684,N_9480,N_9367);
and U9685 (N_9685,N_9469,N_9413);
or U9686 (N_9686,N_9376,N_9498);
nand U9687 (N_9687,N_9319,N_9392);
nand U9688 (N_9688,N_9474,N_9337);
or U9689 (N_9689,N_9276,N_9257);
or U9690 (N_9690,N_9409,N_9482);
or U9691 (N_9691,N_9367,N_9260);
nand U9692 (N_9692,N_9303,N_9467);
nor U9693 (N_9693,N_9332,N_9420);
and U9694 (N_9694,N_9395,N_9411);
and U9695 (N_9695,N_9335,N_9481);
nor U9696 (N_9696,N_9456,N_9376);
xor U9697 (N_9697,N_9405,N_9413);
nor U9698 (N_9698,N_9464,N_9471);
or U9699 (N_9699,N_9436,N_9281);
and U9700 (N_9700,N_9331,N_9256);
nor U9701 (N_9701,N_9433,N_9393);
and U9702 (N_9702,N_9285,N_9252);
or U9703 (N_9703,N_9479,N_9253);
nand U9704 (N_9704,N_9291,N_9377);
xnor U9705 (N_9705,N_9462,N_9372);
nor U9706 (N_9706,N_9442,N_9423);
nor U9707 (N_9707,N_9267,N_9268);
xor U9708 (N_9708,N_9372,N_9440);
nand U9709 (N_9709,N_9483,N_9300);
and U9710 (N_9710,N_9395,N_9457);
xor U9711 (N_9711,N_9353,N_9379);
and U9712 (N_9712,N_9294,N_9495);
or U9713 (N_9713,N_9473,N_9392);
or U9714 (N_9714,N_9432,N_9301);
and U9715 (N_9715,N_9283,N_9442);
nand U9716 (N_9716,N_9339,N_9402);
nand U9717 (N_9717,N_9307,N_9326);
nand U9718 (N_9718,N_9271,N_9416);
and U9719 (N_9719,N_9341,N_9467);
xor U9720 (N_9720,N_9320,N_9390);
nand U9721 (N_9721,N_9370,N_9256);
xor U9722 (N_9722,N_9395,N_9362);
or U9723 (N_9723,N_9391,N_9301);
nor U9724 (N_9724,N_9456,N_9323);
nand U9725 (N_9725,N_9307,N_9460);
xnor U9726 (N_9726,N_9294,N_9460);
or U9727 (N_9727,N_9289,N_9446);
and U9728 (N_9728,N_9445,N_9262);
xnor U9729 (N_9729,N_9257,N_9432);
and U9730 (N_9730,N_9261,N_9375);
xnor U9731 (N_9731,N_9468,N_9327);
nor U9732 (N_9732,N_9371,N_9287);
or U9733 (N_9733,N_9462,N_9255);
xnor U9734 (N_9734,N_9377,N_9497);
nor U9735 (N_9735,N_9277,N_9385);
nor U9736 (N_9736,N_9358,N_9381);
or U9737 (N_9737,N_9421,N_9375);
nor U9738 (N_9738,N_9280,N_9357);
or U9739 (N_9739,N_9382,N_9457);
or U9740 (N_9740,N_9377,N_9367);
nand U9741 (N_9741,N_9440,N_9355);
nand U9742 (N_9742,N_9312,N_9327);
nand U9743 (N_9743,N_9468,N_9367);
nor U9744 (N_9744,N_9306,N_9470);
nor U9745 (N_9745,N_9411,N_9293);
and U9746 (N_9746,N_9385,N_9478);
or U9747 (N_9747,N_9313,N_9357);
nor U9748 (N_9748,N_9451,N_9468);
nand U9749 (N_9749,N_9309,N_9377);
and U9750 (N_9750,N_9556,N_9577);
or U9751 (N_9751,N_9502,N_9567);
and U9752 (N_9752,N_9658,N_9620);
xor U9753 (N_9753,N_9696,N_9723);
nor U9754 (N_9754,N_9548,N_9511);
xor U9755 (N_9755,N_9640,N_9619);
xor U9756 (N_9756,N_9503,N_9552);
xor U9757 (N_9757,N_9614,N_9598);
xnor U9758 (N_9758,N_9516,N_9508);
and U9759 (N_9759,N_9607,N_9547);
xor U9760 (N_9760,N_9505,N_9527);
nor U9761 (N_9761,N_9674,N_9671);
nor U9762 (N_9762,N_9659,N_9745);
xor U9763 (N_9763,N_9690,N_9717);
or U9764 (N_9764,N_9626,N_9738);
and U9765 (N_9765,N_9629,N_9689);
nor U9766 (N_9766,N_9722,N_9656);
xnor U9767 (N_9767,N_9720,N_9563);
xor U9768 (N_9768,N_9681,N_9682);
xor U9769 (N_9769,N_9729,N_9582);
nand U9770 (N_9770,N_9538,N_9521);
and U9771 (N_9771,N_9572,N_9518);
xnor U9772 (N_9772,N_9710,N_9686);
xor U9773 (N_9773,N_9721,N_9712);
xnor U9774 (N_9774,N_9550,N_9597);
nand U9775 (N_9775,N_9676,N_9741);
nor U9776 (N_9776,N_9529,N_9535);
nand U9777 (N_9777,N_9517,N_9665);
or U9778 (N_9778,N_9675,N_9501);
and U9779 (N_9779,N_9705,N_9513);
nand U9780 (N_9780,N_9641,N_9555);
or U9781 (N_9781,N_9673,N_9525);
xor U9782 (N_9782,N_9726,N_9559);
nand U9783 (N_9783,N_9624,N_9747);
xor U9784 (N_9784,N_9585,N_9684);
nand U9785 (N_9785,N_9638,N_9546);
nand U9786 (N_9786,N_9730,N_9584);
xor U9787 (N_9787,N_9688,N_9603);
xor U9788 (N_9788,N_9699,N_9522);
or U9789 (N_9789,N_9691,N_9731);
nand U9790 (N_9790,N_9743,N_9561);
or U9791 (N_9791,N_9703,N_9683);
or U9792 (N_9792,N_9570,N_9576);
nor U9793 (N_9793,N_9617,N_9541);
and U9794 (N_9794,N_9558,N_9672);
xor U9795 (N_9795,N_9540,N_9718);
xor U9796 (N_9796,N_9532,N_9605);
xor U9797 (N_9797,N_9588,N_9654);
and U9798 (N_9798,N_9666,N_9647);
nor U9799 (N_9799,N_9661,N_9519);
xor U9800 (N_9800,N_9560,N_9589);
xor U9801 (N_9801,N_9510,N_9677);
and U9802 (N_9802,N_9644,N_9500);
xnor U9803 (N_9803,N_9531,N_9571);
and U9804 (N_9804,N_9643,N_9714);
xor U9805 (N_9805,N_9711,N_9615);
or U9806 (N_9806,N_9507,N_9627);
xnor U9807 (N_9807,N_9634,N_9549);
or U9808 (N_9808,N_9612,N_9574);
or U9809 (N_9809,N_9590,N_9581);
xnor U9810 (N_9810,N_9602,N_9650);
nor U9811 (N_9811,N_9704,N_9740);
xnor U9812 (N_9812,N_9606,N_9685);
nand U9813 (N_9813,N_9551,N_9653);
or U9814 (N_9814,N_9706,N_9664);
nand U9815 (N_9815,N_9655,N_9600);
xor U9816 (N_9816,N_9568,N_9749);
and U9817 (N_9817,N_9663,N_9724);
or U9818 (N_9818,N_9744,N_9630);
or U9819 (N_9819,N_9520,N_9524);
nor U9820 (N_9820,N_9586,N_9575);
or U9821 (N_9821,N_9700,N_9573);
and U9822 (N_9822,N_9725,N_9680);
nor U9823 (N_9823,N_9735,N_9732);
nor U9824 (N_9824,N_9526,N_9679);
and U9825 (N_9825,N_9727,N_9622);
nor U9826 (N_9826,N_9702,N_9534);
and U9827 (N_9827,N_9748,N_9639);
nand U9828 (N_9828,N_9746,N_9569);
xor U9829 (N_9829,N_9695,N_9609);
nor U9830 (N_9830,N_9557,N_9737);
xor U9831 (N_9831,N_9633,N_9566);
xor U9832 (N_9832,N_9583,N_9565);
nor U9833 (N_9833,N_9707,N_9539);
or U9834 (N_9834,N_9578,N_9596);
nor U9835 (N_9835,N_9636,N_9530);
or U9836 (N_9836,N_9719,N_9545);
xnor U9837 (N_9837,N_9713,N_9514);
xnor U9838 (N_9838,N_9536,N_9708);
xnor U9839 (N_9839,N_9594,N_9554);
and U9840 (N_9840,N_9506,N_9604);
xnor U9841 (N_9841,N_9593,N_9562);
nor U9842 (N_9842,N_9693,N_9504);
nor U9843 (N_9843,N_9736,N_9657);
nor U9844 (N_9844,N_9608,N_9698);
xor U9845 (N_9845,N_9742,N_9591);
nand U9846 (N_9846,N_9625,N_9646);
nand U9847 (N_9847,N_9543,N_9579);
nor U9848 (N_9848,N_9660,N_9635);
xor U9849 (N_9849,N_9715,N_9697);
nor U9850 (N_9850,N_9610,N_9595);
xor U9851 (N_9851,N_9599,N_9533);
nand U9852 (N_9852,N_9716,N_9515);
nor U9853 (N_9853,N_9616,N_9728);
and U9854 (N_9854,N_9523,N_9662);
nor U9855 (N_9855,N_9537,N_9528);
nand U9856 (N_9856,N_9637,N_9669);
xnor U9857 (N_9857,N_9652,N_9694);
nand U9858 (N_9858,N_9734,N_9544);
and U9859 (N_9859,N_9668,N_9628);
or U9860 (N_9860,N_9667,N_9632);
or U9861 (N_9861,N_9509,N_9613);
or U9862 (N_9862,N_9587,N_9618);
and U9863 (N_9863,N_9642,N_9512);
nand U9864 (N_9864,N_9580,N_9649);
xnor U9865 (N_9865,N_9701,N_9733);
or U9866 (N_9866,N_9564,N_9670);
xnor U9867 (N_9867,N_9542,N_9601);
and U9868 (N_9868,N_9553,N_9651);
nor U9869 (N_9869,N_9592,N_9648);
nor U9870 (N_9870,N_9645,N_9687);
or U9871 (N_9871,N_9739,N_9621);
or U9872 (N_9872,N_9709,N_9611);
nor U9873 (N_9873,N_9631,N_9678);
xnor U9874 (N_9874,N_9623,N_9692);
xnor U9875 (N_9875,N_9577,N_9728);
nand U9876 (N_9876,N_9706,N_9508);
or U9877 (N_9877,N_9580,N_9598);
and U9878 (N_9878,N_9545,N_9633);
and U9879 (N_9879,N_9510,N_9563);
or U9880 (N_9880,N_9516,N_9616);
and U9881 (N_9881,N_9572,N_9691);
nand U9882 (N_9882,N_9507,N_9508);
nor U9883 (N_9883,N_9533,N_9694);
and U9884 (N_9884,N_9607,N_9577);
nand U9885 (N_9885,N_9630,N_9738);
or U9886 (N_9886,N_9518,N_9721);
xnor U9887 (N_9887,N_9603,N_9710);
nor U9888 (N_9888,N_9683,N_9500);
and U9889 (N_9889,N_9646,N_9620);
nand U9890 (N_9890,N_9574,N_9576);
and U9891 (N_9891,N_9686,N_9716);
or U9892 (N_9892,N_9516,N_9514);
nor U9893 (N_9893,N_9614,N_9595);
or U9894 (N_9894,N_9606,N_9628);
xor U9895 (N_9895,N_9596,N_9726);
nor U9896 (N_9896,N_9736,N_9733);
xor U9897 (N_9897,N_9573,N_9541);
nand U9898 (N_9898,N_9704,N_9663);
or U9899 (N_9899,N_9590,N_9583);
xor U9900 (N_9900,N_9599,N_9711);
nand U9901 (N_9901,N_9571,N_9735);
nand U9902 (N_9902,N_9625,N_9612);
or U9903 (N_9903,N_9545,N_9565);
xor U9904 (N_9904,N_9742,N_9637);
xnor U9905 (N_9905,N_9539,N_9500);
nand U9906 (N_9906,N_9749,N_9702);
and U9907 (N_9907,N_9539,N_9589);
xnor U9908 (N_9908,N_9740,N_9657);
or U9909 (N_9909,N_9519,N_9720);
nand U9910 (N_9910,N_9615,N_9713);
or U9911 (N_9911,N_9621,N_9748);
xnor U9912 (N_9912,N_9545,N_9577);
xnor U9913 (N_9913,N_9643,N_9502);
nor U9914 (N_9914,N_9516,N_9662);
or U9915 (N_9915,N_9541,N_9511);
nor U9916 (N_9916,N_9696,N_9746);
or U9917 (N_9917,N_9633,N_9735);
nor U9918 (N_9918,N_9681,N_9512);
xnor U9919 (N_9919,N_9564,N_9551);
and U9920 (N_9920,N_9548,N_9745);
xnor U9921 (N_9921,N_9556,N_9658);
nor U9922 (N_9922,N_9549,N_9513);
nand U9923 (N_9923,N_9572,N_9667);
xnor U9924 (N_9924,N_9665,N_9593);
or U9925 (N_9925,N_9547,N_9500);
and U9926 (N_9926,N_9548,N_9718);
nand U9927 (N_9927,N_9570,N_9712);
nand U9928 (N_9928,N_9741,N_9726);
or U9929 (N_9929,N_9605,N_9730);
or U9930 (N_9930,N_9684,N_9698);
nand U9931 (N_9931,N_9506,N_9695);
or U9932 (N_9932,N_9644,N_9610);
or U9933 (N_9933,N_9698,N_9723);
or U9934 (N_9934,N_9712,N_9724);
nor U9935 (N_9935,N_9655,N_9523);
nand U9936 (N_9936,N_9565,N_9581);
xnor U9937 (N_9937,N_9612,N_9547);
nor U9938 (N_9938,N_9697,N_9560);
nor U9939 (N_9939,N_9522,N_9713);
and U9940 (N_9940,N_9559,N_9619);
nand U9941 (N_9941,N_9631,N_9656);
or U9942 (N_9942,N_9601,N_9734);
and U9943 (N_9943,N_9531,N_9687);
and U9944 (N_9944,N_9542,N_9670);
xnor U9945 (N_9945,N_9642,N_9600);
or U9946 (N_9946,N_9747,N_9628);
and U9947 (N_9947,N_9737,N_9748);
nand U9948 (N_9948,N_9548,N_9516);
xnor U9949 (N_9949,N_9743,N_9687);
nand U9950 (N_9950,N_9638,N_9639);
xnor U9951 (N_9951,N_9715,N_9507);
and U9952 (N_9952,N_9620,N_9512);
and U9953 (N_9953,N_9509,N_9523);
nand U9954 (N_9954,N_9652,N_9659);
nor U9955 (N_9955,N_9518,N_9571);
and U9956 (N_9956,N_9505,N_9678);
and U9957 (N_9957,N_9586,N_9520);
and U9958 (N_9958,N_9530,N_9659);
and U9959 (N_9959,N_9574,N_9598);
or U9960 (N_9960,N_9684,N_9563);
and U9961 (N_9961,N_9636,N_9645);
and U9962 (N_9962,N_9720,N_9696);
nand U9963 (N_9963,N_9661,N_9690);
and U9964 (N_9964,N_9500,N_9595);
or U9965 (N_9965,N_9510,N_9749);
nor U9966 (N_9966,N_9720,N_9611);
or U9967 (N_9967,N_9541,N_9591);
nor U9968 (N_9968,N_9564,N_9588);
and U9969 (N_9969,N_9576,N_9612);
or U9970 (N_9970,N_9626,N_9610);
nand U9971 (N_9971,N_9623,N_9706);
and U9972 (N_9972,N_9585,N_9694);
and U9973 (N_9973,N_9625,N_9585);
and U9974 (N_9974,N_9740,N_9501);
nand U9975 (N_9975,N_9668,N_9639);
nor U9976 (N_9976,N_9630,N_9583);
nand U9977 (N_9977,N_9712,N_9537);
or U9978 (N_9978,N_9665,N_9722);
or U9979 (N_9979,N_9627,N_9567);
nand U9980 (N_9980,N_9745,N_9592);
and U9981 (N_9981,N_9651,N_9557);
and U9982 (N_9982,N_9692,N_9533);
nand U9983 (N_9983,N_9662,N_9672);
and U9984 (N_9984,N_9690,N_9612);
or U9985 (N_9985,N_9737,N_9746);
nor U9986 (N_9986,N_9541,N_9685);
and U9987 (N_9987,N_9500,N_9527);
nor U9988 (N_9988,N_9561,N_9689);
nand U9989 (N_9989,N_9506,N_9599);
nor U9990 (N_9990,N_9683,N_9586);
and U9991 (N_9991,N_9724,N_9538);
nor U9992 (N_9992,N_9732,N_9515);
xnor U9993 (N_9993,N_9724,N_9547);
and U9994 (N_9994,N_9637,N_9630);
and U9995 (N_9995,N_9667,N_9505);
nor U9996 (N_9996,N_9723,N_9652);
and U9997 (N_9997,N_9612,N_9541);
or U9998 (N_9998,N_9562,N_9514);
and U9999 (N_9999,N_9573,N_9691);
xnor U10000 (N_10000,N_9944,N_9979);
or U10001 (N_10001,N_9913,N_9846);
xor U10002 (N_10002,N_9828,N_9884);
xnor U10003 (N_10003,N_9922,N_9782);
and U10004 (N_10004,N_9916,N_9761);
and U10005 (N_10005,N_9926,N_9938);
nor U10006 (N_10006,N_9790,N_9854);
nor U10007 (N_10007,N_9806,N_9811);
nand U10008 (N_10008,N_9779,N_9927);
xor U10009 (N_10009,N_9934,N_9982);
nand U10010 (N_10010,N_9925,N_9805);
and U10011 (N_10011,N_9835,N_9977);
nand U10012 (N_10012,N_9980,N_9851);
and U10013 (N_10013,N_9885,N_9853);
or U10014 (N_10014,N_9917,N_9996);
and U10015 (N_10015,N_9904,N_9825);
nor U10016 (N_10016,N_9882,N_9914);
nor U10017 (N_10017,N_9787,N_9892);
nand U10018 (N_10018,N_9896,N_9831);
or U10019 (N_10019,N_9860,N_9819);
nor U10020 (N_10020,N_9883,N_9997);
and U10021 (N_10021,N_9942,N_9918);
xnor U10022 (N_10022,N_9903,N_9875);
and U10023 (N_10023,N_9893,N_9798);
xor U10024 (N_10024,N_9850,N_9866);
and U10025 (N_10025,N_9836,N_9778);
and U10026 (N_10026,N_9911,N_9908);
and U10027 (N_10027,N_9858,N_9847);
xor U10028 (N_10028,N_9784,N_9877);
nor U10029 (N_10029,N_9848,N_9767);
xor U10030 (N_10030,N_9766,N_9910);
nand U10031 (N_10031,N_9786,N_9834);
nand U10032 (N_10032,N_9861,N_9753);
nor U10033 (N_10033,N_9750,N_9960);
or U10034 (N_10034,N_9824,N_9890);
and U10035 (N_10035,N_9775,N_9762);
and U10036 (N_10036,N_9953,N_9765);
xnor U10037 (N_10037,N_9985,N_9958);
nor U10038 (N_10038,N_9952,N_9795);
xnor U10039 (N_10039,N_9933,N_9951);
and U10040 (N_10040,N_9921,N_9948);
or U10041 (N_10041,N_9919,N_9876);
nor U10042 (N_10042,N_9788,N_9974);
and U10043 (N_10043,N_9895,N_9844);
and U10044 (N_10044,N_9832,N_9769);
nor U10045 (N_10045,N_9969,N_9807);
or U10046 (N_10046,N_9907,N_9965);
xnor U10047 (N_10047,N_9801,N_9770);
or U10048 (N_10048,N_9783,N_9880);
and U10049 (N_10049,N_9781,N_9868);
nand U10050 (N_10050,N_9773,N_9812);
and U10051 (N_10051,N_9931,N_9827);
nor U10052 (N_10052,N_9891,N_9864);
or U10053 (N_10053,N_9772,N_9794);
xor U10054 (N_10054,N_9940,N_9838);
nand U10055 (N_10055,N_9791,N_9929);
and U10056 (N_10056,N_9818,N_9930);
and U10057 (N_10057,N_9785,N_9870);
or U10058 (N_10058,N_9898,N_9797);
and U10059 (N_10059,N_9966,N_9839);
and U10060 (N_10060,N_9852,N_9962);
nor U10061 (N_10061,N_9842,N_9751);
nand U10062 (N_10062,N_9774,N_9970);
nand U10063 (N_10063,N_9889,N_9792);
or U10064 (N_10064,N_9820,N_9999);
nand U10065 (N_10065,N_9862,N_9961);
and U10066 (N_10066,N_9768,N_9814);
nor U10067 (N_10067,N_9793,N_9803);
and U10068 (N_10068,N_9950,N_9764);
or U10069 (N_10069,N_9856,N_9989);
xor U10070 (N_10070,N_9777,N_9990);
nor U10071 (N_10071,N_9984,N_9986);
xor U10072 (N_10072,N_9995,N_9888);
and U10073 (N_10073,N_9956,N_9758);
or U10074 (N_10074,N_9945,N_9867);
and U10075 (N_10075,N_9859,N_9992);
and U10076 (N_10076,N_9967,N_9849);
nand U10077 (N_10077,N_9954,N_9817);
xnor U10078 (N_10078,N_9897,N_9988);
xor U10079 (N_10079,N_9972,N_9809);
nand U10080 (N_10080,N_9802,N_9915);
or U10081 (N_10081,N_9959,N_9833);
and U10082 (N_10082,N_9998,N_9909);
and U10083 (N_10083,N_9936,N_9789);
and U10084 (N_10084,N_9928,N_9826);
xnor U10085 (N_10085,N_9899,N_9804);
xnor U10086 (N_10086,N_9901,N_9976);
and U10087 (N_10087,N_9957,N_9874);
and U10088 (N_10088,N_9799,N_9872);
or U10089 (N_10089,N_9973,N_9756);
xor U10090 (N_10090,N_9810,N_9993);
and U10091 (N_10091,N_9943,N_9947);
and U10092 (N_10092,N_9902,N_9887);
nand U10093 (N_10093,N_9808,N_9763);
and U10094 (N_10094,N_9780,N_9813);
and U10095 (N_10095,N_9881,N_9939);
nand U10096 (N_10096,N_9857,N_9923);
and U10097 (N_10097,N_9983,N_9987);
or U10098 (N_10098,N_9946,N_9776);
and U10099 (N_10099,N_9841,N_9955);
or U10100 (N_10100,N_9771,N_9941);
and U10101 (N_10101,N_9843,N_9886);
and U10102 (N_10102,N_9800,N_9815);
nand U10103 (N_10103,N_9855,N_9963);
xor U10104 (N_10104,N_9906,N_9816);
and U10105 (N_10105,N_9871,N_9878);
nand U10106 (N_10106,N_9937,N_9935);
xor U10107 (N_10107,N_9759,N_9981);
nor U10108 (N_10108,N_9863,N_9829);
and U10109 (N_10109,N_9757,N_9971);
or U10110 (N_10110,N_9754,N_9840);
xor U10111 (N_10111,N_9879,N_9873);
nand U10112 (N_10112,N_9964,N_9752);
nand U10113 (N_10113,N_9905,N_9865);
xnor U10114 (N_10114,N_9920,N_9755);
nor U10115 (N_10115,N_9912,N_9830);
or U10116 (N_10116,N_9894,N_9900);
or U10117 (N_10117,N_9924,N_9978);
nand U10118 (N_10118,N_9845,N_9822);
or U10119 (N_10119,N_9821,N_9991);
or U10120 (N_10120,N_9760,N_9994);
or U10121 (N_10121,N_9869,N_9823);
nor U10122 (N_10122,N_9796,N_9968);
nand U10123 (N_10123,N_9837,N_9932);
xor U10124 (N_10124,N_9975,N_9949);
or U10125 (N_10125,N_9997,N_9769);
xnor U10126 (N_10126,N_9920,N_9776);
or U10127 (N_10127,N_9925,N_9982);
nand U10128 (N_10128,N_9854,N_9948);
or U10129 (N_10129,N_9924,N_9853);
xnor U10130 (N_10130,N_9859,N_9864);
nand U10131 (N_10131,N_9982,N_9774);
nand U10132 (N_10132,N_9850,N_9878);
or U10133 (N_10133,N_9869,N_9962);
nor U10134 (N_10134,N_9817,N_9916);
nor U10135 (N_10135,N_9832,N_9822);
or U10136 (N_10136,N_9842,N_9863);
nand U10137 (N_10137,N_9802,N_9852);
nand U10138 (N_10138,N_9772,N_9766);
xnor U10139 (N_10139,N_9882,N_9913);
xnor U10140 (N_10140,N_9764,N_9880);
nor U10141 (N_10141,N_9960,N_9917);
and U10142 (N_10142,N_9967,N_9962);
or U10143 (N_10143,N_9817,N_9828);
nand U10144 (N_10144,N_9756,N_9791);
nor U10145 (N_10145,N_9806,N_9895);
nand U10146 (N_10146,N_9992,N_9783);
and U10147 (N_10147,N_9910,N_9821);
and U10148 (N_10148,N_9888,N_9838);
xor U10149 (N_10149,N_9936,N_9906);
nor U10150 (N_10150,N_9834,N_9893);
nand U10151 (N_10151,N_9907,N_9824);
xnor U10152 (N_10152,N_9934,N_9806);
or U10153 (N_10153,N_9891,N_9803);
or U10154 (N_10154,N_9780,N_9830);
and U10155 (N_10155,N_9851,N_9979);
nand U10156 (N_10156,N_9952,N_9983);
nand U10157 (N_10157,N_9992,N_9961);
nor U10158 (N_10158,N_9968,N_9847);
nand U10159 (N_10159,N_9955,N_9910);
nand U10160 (N_10160,N_9989,N_9837);
or U10161 (N_10161,N_9795,N_9943);
or U10162 (N_10162,N_9841,N_9894);
or U10163 (N_10163,N_9827,N_9829);
and U10164 (N_10164,N_9989,N_9833);
and U10165 (N_10165,N_9909,N_9857);
xnor U10166 (N_10166,N_9950,N_9918);
nor U10167 (N_10167,N_9951,N_9939);
nand U10168 (N_10168,N_9870,N_9986);
xor U10169 (N_10169,N_9779,N_9775);
xnor U10170 (N_10170,N_9800,N_9762);
nor U10171 (N_10171,N_9867,N_9879);
xor U10172 (N_10172,N_9982,N_9967);
or U10173 (N_10173,N_9949,N_9942);
nand U10174 (N_10174,N_9979,N_9798);
or U10175 (N_10175,N_9814,N_9767);
or U10176 (N_10176,N_9925,N_9783);
xor U10177 (N_10177,N_9907,N_9986);
and U10178 (N_10178,N_9909,N_9828);
nand U10179 (N_10179,N_9782,N_9998);
nor U10180 (N_10180,N_9924,N_9994);
nand U10181 (N_10181,N_9798,N_9939);
nor U10182 (N_10182,N_9995,N_9913);
xnor U10183 (N_10183,N_9781,N_9775);
xor U10184 (N_10184,N_9832,N_9908);
nand U10185 (N_10185,N_9926,N_9911);
nand U10186 (N_10186,N_9985,N_9801);
nor U10187 (N_10187,N_9925,N_9881);
or U10188 (N_10188,N_9809,N_9962);
nand U10189 (N_10189,N_9968,N_9815);
nand U10190 (N_10190,N_9806,N_9815);
or U10191 (N_10191,N_9878,N_9797);
xor U10192 (N_10192,N_9862,N_9938);
xor U10193 (N_10193,N_9911,N_9958);
or U10194 (N_10194,N_9834,N_9947);
nand U10195 (N_10195,N_9897,N_9976);
and U10196 (N_10196,N_9856,N_9789);
or U10197 (N_10197,N_9884,N_9898);
xnor U10198 (N_10198,N_9951,N_9902);
xnor U10199 (N_10199,N_9761,N_9818);
nand U10200 (N_10200,N_9854,N_9819);
nor U10201 (N_10201,N_9753,N_9915);
xnor U10202 (N_10202,N_9973,N_9958);
and U10203 (N_10203,N_9923,N_9948);
and U10204 (N_10204,N_9985,N_9858);
nor U10205 (N_10205,N_9845,N_9902);
and U10206 (N_10206,N_9813,N_9781);
and U10207 (N_10207,N_9861,N_9869);
xnor U10208 (N_10208,N_9757,N_9865);
nor U10209 (N_10209,N_9984,N_9804);
xnor U10210 (N_10210,N_9964,N_9882);
xnor U10211 (N_10211,N_9863,N_9839);
nand U10212 (N_10212,N_9918,N_9915);
nor U10213 (N_10213,N_9890,N_9860);
and U10214 (N_10214,N_9813,N_9856);
and U10215 (N_10215,N_9778,N_9980);
xor U10216 (N_10216,N_9932,N_9770);
or U10217 (N_10217,N_9953,N_9908);
or U10218 (N_10218,N_9896,N_9972);
nor U10219 (N_10219,N_9963,N_9889);
or U10220 (N_10220,N_9765,N_9792);
and U10221 (N_10221,N_9773,N_9879);
nand U10222 (N_10222,N_9935,N_9917);
xnor U10223 (N_10223,N_9783,N_9958);
nand U10224 (N_10224,N_9783,N_9841);
and U10225 (N_10225,N_9833,N_9880);
nor U10226 (N_10226,N_9949,N_9965);
and U10227 (N_10227,N_9842,N_9811);
and U10228 (N_10228,N_9797,N_9838);
xnor U10229 (N_10229,N_9861,N_9769);
nor U10230 (N_10230,N_9773,N_9751);
nor U10231 (N_10231,N_9945,N_9920);
and U10232 (N_10232,N_9849,N_9933);
xnor U10233 (N_10233,N_9928,N_9981);
xnor U10234 (N_10234,N_9980,N_9837);
or U10235 (N_10235,N_9782,N_9798);
nor U10236 (N_10236,N_9961,N_9927);
or U10237 (N_10237,N_9915,N_9966);
xnor U10238 (N_10238,N_9989,N_9901);
and U10239 (N_10239,N_9963,N_9915);
nor U10240 (N_10240,N_9753,N_9908);
and U10241 (N_10241,N_9943,N_9904);
nor U10242 (N_10242,N_9997,N_9831);
or U10243 (N_10243,N_9768,N_9818);
or U10244 (N_10244,N_9899,N_9904);
or U10245 (N_10245,N_9915,N_9855);
and U10246 (N_10246,N_9839,N_9773);
and U10247 (N_10247,N_9897,N_9941);
or U10248 (N_10248,N_9805,N_9752);
and U10249 (N_10249,N_9842,N_9999);
nor U10250 (N_10250,N_10123,N_10086);
nor U10251 (N_10251,N_10110,N_10227);
nor U10252 (N_10252,N_10025,N_10095);
nor U10253 (N_10253,N_10157,N_10220);
xor U10254 (N_10254,N_10001,N_10104);
xor U10255 (N_10255,N_10239,N_10152);
xnor U10256 (N_10256,N_10049,N_10207);
nor U10257 (N_10257,N_10184,N_10174);
nand U10258 (N_10258,N_10097,N_10083);
or U10259 (N_10259,N_10158,N_10117);
or U10260 (N_10260,N_10208,N_10091);
nand U10261 (N_10261,N_10010,N_10004);
and U10262 (N_10262,N_10132,N_10163);
nand U10263 (N_10263,N_10186,N_10214);
nor U10264 (N_10264,N_10199,N_10216);
or U10265 (N_10265,N_10231,N_10213);
and U10266 (N_10266,N_10074,N_10180);
xnor U10267 (N_10267,N_10242,N_10176);
or U10268 (N_10268,N_10022,N_10177);
nand U10269 (N_10269,N_10203,N_10169);
xnor U10270 (N_10270,N_10032,N_10234);
nand U10271 (N_10271,N_10218,N_10012);
and U10272 (N_10272,N_10081,N_10172);
or U10273 (N_10273,N_10089,N_10046);
and U10274 (N_10274,N_10047,N_10087);
and U10275 (N_10275,N_10000,N_10175);
or U10276 (N_10276,N_10206,N_10210);
xor U10277 (N_10277,N_10135,N_10136);
nor U10278 (N_10278,N_10201,N_10181);
xnor U10279 (N_10279,N_10171,N_10112);
nor U10280 (N_10280,N_10064,N_10063);
nor U10281 (N_10281,N_10071,N_10014);
and U10282 (N_10282,N_10228,N_10246);
nor U10283 (N_10283,N_10031,N_10125);
xor U10284 (N_10284,N_10072,N_10209);
xor U10285 (N_10285,N_10044,N_10215);
or U10286 (N_10286,N_10098,N_10153);
nor U10287 (N_10287,N_10198,N_10235);
nor U10288 (N_10288,N_10017,N_10193);
nor U10289 (N_10289,N_10043,N_10232);
nand U10290 (N_10290,N_10173,N_10102);
nand U10291 (N_10291,N_10062,N_10093);
xor U10292 (N_10292,N_10058,N_10129);
and U10293 (N_10293,N_10223,N_10142);
nor U10294 (N_10294,N_10050,N_10160);
nand U10295 (N_10295,N_10077,N_10080);
or U10296 (N_10296,N_10109,N_10008);
nor U10297 (N_10297,N_10204,N_10196);
and U10298 (N_10298,N_10108,N_10154);
nor U10299 (N_10299,N_10066,N_10055);
nor U10300 (N_10300,N_10159,N_10090);
xnor U10301 (N_10301,N_10145,N_10121);
or U10302 (N_10302,N_10187,N_10028);
nor U10303 (N_10303,N_10144,N_10229);
nand U10304 (N_10304,N_10226,N_10131);
nand U10305 (N_10305,N_10059,N_10076);
xor U10306 (N_10306,N_10057,N_10079);
nand U10307 (N_10307,N_10065,N_10202);
nand U10308 (N_10308,N_10221,N_10027);
and U10309 (N_10309,N_10245,N_10197);
nand U10310 (N_10310,N_10007,N_10069);
xnor U10311 (N_10311,N_10238,N_10224);
xor U10312 (N_10312,N_10101,N_10016);
xnor U10313 (N_10313,N_10040,N_10155);
nand U10314 (N_10314,N_10191,N_10013);
or U10315 (N_10315,N_10192,N_10051);
and U10316 (N_10316,N_10118,N_10088);
or U10317 (N_10317,N_10230,N_10190);
nor U10318 (N_10318,N_10060,N_10100);
nand U10319 (N_10319,N_10185,N_10240);
or U10320 (N_10320,N_10021,N_10078);
nor U10321 (N_10321,N_10130,N_10164);
nand U10322 (N_10322,N_10225,N_10105);
xor U10323 (N_10323,N_10212,N_10011);
nor U10324 (N_10324,N_10096,N_10033);
or U10325 (N_10325,N_10085,N_10084);
xor U10326 (N_10326,N_10026,N_10143);
nor U10327 (N_10327,N_10030,N_10237);
xnor U10328 (N_10328,N_10124,N_10120);
or U10329 (N_10329,N_10183,N_10222);
and U10330 (N_10330,N_10140,N_10119);
and U10331 (N_10331,N_10205,N_10166);
or U10332 (N_10332,N_10149,N_10094);
and U10333 (N_10333,N_10106,N_10002);
nor U10334 (N_10334,N_10148,N_10075);
xor U10335 (N_10335,N_10038,N_10217);
xnor U10336 (N_10336,N_10006,N_10248);
xor U10337 (N_10337,N_10182,N_10041);
nor U10338 (N_10338,N_10162,N_10053);
or U10339 (N_10339,N_10167,N_10116);
xnor U10340 (N_10340,N_10115,N_10194);
nand U10341 (N_10341,N_10133,N_10039);
or U10342 (N_10342,N_10211,N_10054);
nor U10343 (N_10343,N_10082,N_10092);
or U10344 (N_10344,N_10029,N_10139);
nand U10345 (N_10345,N_10052,N_10018);
nand U10346 (N_10346,N_10137,N_10019);
nand U10347 (N_10347,N_10127,N_10107);
and U10348 (N_10348,N_10128,N_10015);
nor U10349 (N_10349,N_10151,N_10141);
nor U10350 (N_10350,N_10168,N_10073);
nor U10351 (N_10351,N_10122,N_10161);
nand U10352 (N_10352,N_10219,N_10236);
xnor U10353 (N_10353,N_10111,N_10189);
or U10354 (N_10354,N_10003,N_10146);
nor U10355 (N_10355,N_10247,N_10179);
or U10356 (N_10356,N_10070,N_10147);
xor U10357 (N_10357,N_10243,N_10241);
or U10358 (N_10358,N_10048,N_10165);
nand U10359 (N_10359,N_10178,N_10099);
and U10360 (N_10360,N_10037,N_10023);
nor U10361 (N_10361,N_10188,N_10035);
xor U10362 (N_10362,N_10134,N_10024);
xor U10363 (N_10363,N_10067,N_10061);
or U10364 (N_10364,N_10113,N_10009);
nor U10365 (N_10365,N_10244,N_10233);
nor U10366 (N_10366,N_10150,N_10249);
xnor U10367 (N_10367,N_10103,N_10200);
and U10368 (N_10368,N_10195,N_10036);
xnor U10369 (N_10369,N_10126,N_10068);
nor U10370 (N_10370,N_10156,N_10138);
or U10371 (N_10371,N_10045,N_10056);
nor U10372 (N_10372,N_10114,N_10034);
nand U10373 (N_10373,N_10020,N_10170);
or U10374 (N_10374,N_10042,N_10005);
or U10375 (N_10375,N_10057,N_10068);
xor U10376 (N_10376,N_10126,N_10164);
nor U10377 (N_10377,N_10133,N_10155);
nand U10378 (N_10378,N_10083,N_10090);
nor U10379 (N_10379,N_10065,N_10226);
nor U10380 (N_10380,N_10218,N_10190);
nor U10381 (N_10381,N_10195,N_10135);
or U10382 (N_10382,N_10110,N_10099);
nand U10383 (N_10383,N_10063,N_10088);
and U10384 (N_10384,N_10030,N_10121);
and U10385 (N_10385,N_10205,N_10069);
nor U10386 (N_10386,N_10132,N_10235);
nor U10387 (N_10387,N_10058,N_10207);
nor U10388 (N_10388,N_10229,N_10097);
or U10389 (N_10389,N_10195,N_10063);
or U10390 (N_10390,N_10150,N_10011);
and U10391 (N_10391,N_10220,N_10140);
or U10392 (N_10392,N_10016,N_10127);
or U10393 (N_10393,N_10078,N_10068);
and U10394 (N_10394,N_10005,N_10108);
xor U10395 (N_10395,N_10231,N_10101);
or U10396 (N_10396,N_10171,N_10124);
or U10397 (N_10397,N_10224,N_10089);
nor U10398 (N_10398,N_10120,N_10171);
nand U10399 (N_10399,N_10120,N_10008);
or U10400 (N_10400,N_10141,N_10037);
or U10401 (N_10401,N_10118,N_10164);
nor U10402 (N_10402,N_10219,N_10177);
nor U10403 (N_10403,N_10104,N_10241);
or U10404 (N_10404,N_10069,N_10190);
and U10405 (N_10405,N_10107,N_10137);
nor U10406 (N_10406,N_10033,N_10124);
nor U10407 (N_10407,N_10229,N_10150);
nand U10408 (N_10408,N_10158,N_10154);
xor U10409 (N_10409,N_10244,N_10045);
xor U10410 (N_10410,N_10148,N_10228);
xor U10411 (N_10411,N_10020,N_10157);
nor U10412 (N_10412,N_10000,N_10077);
and U10413 (N_10413,N_10201,N_10113);
nand U10414 (N_10414,N_10062,N_10211);
nor U10415 (N_10415,N_10117,N_10200);
and U10416 (N_10416,N_10211,N_10014);
or U10417 (N_10417,N_10208,N_10128);
nor U10418 (N_10418,N_10081,N_10184);
or U10419 (N_10419,N_10034,N_10010);
or U10420 (N_10420,N_10102,N_10175);
xnor U10421 (N_10421,N_10177,N_10069);
nand U10422 (N_10422,N_10088,N_10053);
or U10423 (N_10423,N_10052,N_10024);
nand U10424 (N_10424,N_10022,N_10140);
or U10425 (N_10425,N_10158,N_10138);
and U10426 (N_10426,N_10220,N_10110);
and U10427 (N_10427,N_10201,N_10147);
nand U10428 (N_10428,N_10023,N_10016);
and U10429 (N_10429,N_10187,N_10108);
and U10430 (N_10430,N_10234,N_10196);
xnor U10431 (N_10431,N_10084,N_10019);
nor U10432 (N_10432,N_10195,N_10144);
xnor U10433 (N_10433,N_10131,N_10133);
xnor U10434 (N_10434,N_10065,N_10035);
nand U10435 (N_10435,N_10205,N_10222);
and U10436 (N_10436,N_10078,N_10097);
and U10437 (N_10437,N_10010,N_10089);
and U10438 (N_10438,N_10118,N_10144);
and U10439 (N_10439,N_10204,N_10085);
and U10440 (N_10440,N_10053,N_10118);
nor U10441 (N_10441,N_10220,N_10136);
nor U10442 (N_10442,N_10149,N_10232);
or U10443 (N_10443,N_10049,N_10133);
and U10444 (N_10444,N_10089,N_10085);
and U10445 (N_10445,N_10082,N_10166);
nand U10446 (N_10446,N_10041,N_10145);
xor U10447 (N_10447,N_10084,N_10043);
and U10448 (N_10448,N_10226,N_10108);
and U10449 (N_10449,N_10204,N_10000);
xor U10450 (N_10450,N_10170,N_10024);
or U10451 (N_10451,N_10091,N_10198);
and U10452 (N_10452,N_10098,N_10231);
nand U10453 (N_10453,N_10221,N_10019);
or U10454 (N_10454,N_10137,N_10007);
and U10455 (N_10455,N_10109,N_10212);
nand U10456 (N_10456,N_10218,N_10198);
nor U10457 (N_10457,N_10160,N_10070);
nand U10458 (N_10458,N_10192,N_10103);
or U10459 (N_10459,N_10039,N_10112);
or U10460 (N_10460,N_10184,N_10088);
nand U10461 (N_10461,N_10108,N_10025);
nand U10462 (N_10462,N_10191,N_10198);
nand U10463 (N_10463,N_10088,N_10176);
nor U10464 (N_10464,N_10042,N_10037);
and U10465 (N_10465,N_10065,N_10124);
nor U10466 (N_10466,N_10187,N_10091);
nand U10467 (N_10467,N_10223,N_10106);
nand U10468 (N_10468,N_10150,N_10216);
or U10469 (N_10469,N_10020,N_10016);
nand U10470 (N_10470,N_10080,N_10170);
and U10471 (N_10471,N_10177,N_10151);
nand U10472 (N_10472,N_10119,N_10042);
or U10473 (N_10473,N_10157,N_10244);
xnor U10474 (N_10474,N_10023,N_10211);
or U10475 (N_10475,N_10166,N_10091);
nor U10476 (N_10476,N_10092,N_10035);
and U10477 (N_10477,N_10228,N_10113);
xnor U10478 (N_10478,N_10179,N_10151);
nand U10479 (N_10479,N_10054,N_10139);
nand U10480 (N_10480,N_10039,N_10183);
nor U10481 (N_10481,N_10194,N_10242);
nand U10482 (N_10482,N_10230,N_10044);
or U10483 (N_10483,N_10096,N_10225);
nand U10484 (N_10484,N_10210,N_10040);
nor U10485 (N_10485,N_10112,N_10094);
and U10486 (N_10486,N_10040,N_10079);
xnor U10487 (N_10487,N_10080,N_10127);
or U10488 (N_10488,N_10212,N_10034);
or U10489 (N_10489,N_10085,N_10190);
nor U10490 (N_10490,N_10046,N_10224);
xor U10491 (N_10491,N_10209,N_10026);
nor U10492 (N_10492,N_10106,N_10022);
or U10493 (N_10493,N_10151,N_10196);
nor U10494 (N_10494,N_10146,N_10223);
nand U10495 (N_10495,N_10017,N_10024);
nor U10496 (N_10496,N_10042,N_10150);
nand U10497 (N_10497,N_10119,N_10028);
nor U10498 (N_10498,N_10141,N_10180);
nand U10499 (N_10499,N_10115,N_10140);
and U10500 (N_10500,N_10406,N_10260);
and U10501 (N_10501,N_10469,N_10320);
and U10502 (N_10502,N_10428,N_10474);
or U10503 (N_10503,N_10454,N_10340);
nor U10504 (N_10504,N_10316,N_10280);
xor U10505 (N_10505,N_10481,N_10263);
nand U10506 (N_10506,N_10321,N_10420);
nor U10507 (N_10507,N_10453,N_10480);
nor U10508 (N_10508,N_10387,N_10265);
nor U10509 (N_10509,N_10254,N_10276);
or U10510 (N_10510,N_10369,N_10336);
and U10511 (N_10511,N_10315,N_10410);
xor U10512 (N_10512,N_10436,N_10365);
nor U10513 (N_10513,N_10490,N_10413);
or U10514 (N_10514,N_10465,N_10430);
nand U10515 (N_10515,N_10298,N_10251);
and U10516 (N_10516,N_10479,N_10455);
nand U10517 (N_10517,N_10429,N_10373);
and U10518 (N_10518,N_10417,N_10293);
xor U10519 (N_10519,N_10271,N_10422);
nand U10520 (N_10520,N_10297,N_10288);
nand U10521 (N_10521,N_10414,N_10359);
nand U10522 (N_10522,N_10355,N_10326);
xor U10523 (N_10523,N_10356,N_10366);
or U10524 (N_10524,N_10312,N_10468);
or U10525 (N_10525,N_10341,N_10449);
and U10526 (N_10526,N_10456,N_10331);
nand U10527 (N_10527,N_10437,N_10444);
nor U10528 (N_10528,N_10302,N_10471);
nor U10529 (N_10529,N_10448,N_10400);
nor U10530 (N_10530,N_10475,N_10394);
or U10531 (N_10531,N_10305,N_10269);
and U10532 (N_10532,N_10277,N_10289);
xor U10533 (N_10533,N_10270,N_10342);
nand U10534 (N_10534,N_10252,N_10311);
nand U10535 (N_10535,N_10499,N_10376);
nor U10536 (N_10536,N_10425,N_10268);
and U10537 (N_10537,N_10409,N_10397);
nor U10538 (N_10538,N_10353,N_10339);
or U10539 (N_10539,N_10354,N_10446);
nand U10540 (N_10540,N_10282,N_10367);
or U10541 (N_10541,N_10404,N_10364);
xnor U10542 (N_10542,N_10303,N_10427);
or U10543 (N_10543,N_10418,N_10439);
nor U10544 (N_10544,N_10402,N_10330);
xor U10545 (N_10545,N_10485,N_10424);
or U10546 (N_10546,N_10493,N_10374);
nand U10547 (N_10547,N_10274,N_10348);
nand U10548 (N_10548,N_10283,N_10349);
nand U10549 (N_10549,N_10377,N_10256);
nand U10550 (N_10550,N_10435,N_10396);
xnor U10551 (N_10551,N_10467,N_10415);
nand U10552 (N_10552,N_10419,N_10257);
or U10553 (N_10553,N_10441,N_10284);
and U10554 (N_10554,N_10497,N_10307);
nor U10555 (N_10555,N_10447,N_10466);
nor U10556 (N_10556,N_10488,N_10266);
xnor U10557 (N_10557,N_10345,N_10462);
or U10558 (N_10558,N_10389,N_10478);
nor U10559 (N_10559,N_10262,N_10328);
nand U10560 (N_10560,N_10433,N_10292);
nor U10561 (N_10561,N_10484,N_10346);
nand U10562 (N_10562,N_10318,N_10395);
and U10563 (N_10563,N_10451,N_10379);
or U10564 (N_10564,N_10391,N_10421);
nor U10565 (N_10565,N_10335,N_10370);
and U10566 (N_10566,N_10290,N_10368);
xnor U10567 (N_10567,N_10495,N_10399);
or U10568 (N_10568,N_10332,N_10489);
nand U10569 (N_10569,N_10412,N_10386);
xor U10570 (N_10570,N_10426,N_10445);
xnor U10571 (N_10571,N_10472,N_10294);
or U10572 (N_10572,N_10486,N_10382);
and U10573 (N_10573,N_10329,N_10295);
or U10574 (N_10574,N_10411,N_10333);
and U10575 (N_10575,N_10264,N_10498);
nor U10576 (N_10576,N_10487,N_10250);
or U10577 (N_10577,N_10423,N_10258);
and U10578 (N_10578,N_10310,N_10325);
and U10579 (N_10579,N_10494,N_10492);
xnor U10580 (N_10580,N_10287,N_10363);
and U10581 (N_10581,N_10253,N_10408);
and U10582 (N_10582,N_10458,N_10324);
xnor U10583 (N_10583,N_10309,N_10375);
nand U10584 (N_10584,N_10463,N_10272);
or U10585 (N_10585,N_10344,N_10390);
nand U10586 (N_10586,N_10319,N_10362);
nor U10587 (N_10587,N_10432,N_10281);
or U10588 (N_10588,N_10491,N_10300);
nand U10589 (N_10589,N_10357,N_10464);
nor U10590 (N_10590,N_10440,N_10306);
xnor U10591 (N_10591,N_10322,N_10378);
nand U10592 (N_10592,N_10476,N_10459);
nand U10593 (N_10593,N_10380,N_10361);
or U10594 (N_10594,N_10317,N_10347);
nor U10595 (N_10595,N_10442,N_10461);
nand U10596 (N_10596,N_10473,N_10381);
and U10597 (N_10597,N_10261,N_10351);
or U10598 (N_10598,N_10275,N_10477);
nand U10599 (N_10599,N_10313,N_10267);
and U10600 (N_10600,N_10450,N_10443);
nand U10601 (N_10601,N_10301,N_10278);
or U10602 (N_10602,N_10405,N_10383);
nor U10603 (N_10603,N_10327,N_10401);
and U10604 (N_10604,N_10279,N_10460);
and U10605 (N_10605,N_10323,N_10338);
or U10606 (N_10606,N_10403,N_10398);
nand U10607 (N_10607,N_10452,N_10334);
and U10608 (N_10608,N_10388,N_10352);
nand U10609 (N_10609,N_10285,N_10286);
nor U10610 (N_10610,N_10392,N_10314);
xnor U10611 (N_10611,N_10431,N_10371);
and U10612 (N_10612,N_10291,N_10343);
nor U10613 (N_10613,N_10416,N_10337);
nor U10614 (N_10614,N_10296,N_10259);
xnor U10615 (N_10615,N_10255,N_10434);
xor U10616 (N_10616,N_10483,N_10358);
xnor U10617 (N_10617,N_10470,N_10273);
xnor U10618 (N_10618,N_10308,N_10385);
or U10619 (N_10619,N_10299,N_10482);
and U10620 (N_10620,N_10360,N_10407);
nand U10621 (N_10621,N_10457,N_10384);
and U10622 (N_10622,N_10438,N_10393);
and U10623 (N_10623,N_10496,N_10372);
nand U10624 (N_10624,N_10304,N_10350);
nand U10625 (N_10625,N_10274,N_10464);
nor U10626 (N_10626,N_10497,N_10297);
nor U10627 (N_10627,N_10286,N_10406);
or U10628 (N_10628,N_10485,N_10291);
nor U10629 (N_10629,N_10361,N_10328);
and U10630 (N_10630,N_10320,N_10395);
or U10631 (N_10631,N_10277,N_10408);
nor U10632 (N_10632,N_10310,N_10252);
xor U10633 (N_10633,N_10445,N_10344);
and U10634 (N_10634,N_10465,N_10254);
xor U10635 (N_10635,N_10271,N_10335);
xor U10636 (N_10636,N_10463,N_10283);
and U10637 (N_10637,N_10455,N_10314);
nor U10638 (N_10638,N_10374,N_10415);
and U10639 (N_10639,N_10448,N_10451);
nor U10640 (N_10640,N_10378,N_10340);
xnor U10641 (N_10641,N_10357,N_10375);
nand U10642 (N_10642,N_10266,N_10451);
nand U10643 (N_10643,N_10336,N_10450);
xor U10644 (N_10644,N_10268,N_10269);
nand U10645 (N_10645,N_10308,N_10253);
or U10646 (N_10646,N_10311,N_10323);
and U10647 (N_10647,N_10338,N_10437);
or U10648 (N_10648,N_10433,N_10475);
or U10649 (N_10649,N_10491,N_10476);
nor U10650 (N_10650,N_10434,N_10290);
and U10651 (N_10651,N_10279,N_10258);
xor U10652 (N_10652,N_10321,N_10408);
or U10653 (N_10653,N_10349,N_10352);
xor U10654 (N_10654,N_10322,N_10464);
xor U10655 (N_10655,N_10344,N_10306);
or U10656 (N_10656,N_10259,N_10314);
and U10657 (N_10657,N_10304,N_10371);
and U10658 (N_10658,N_10404,N_10311);
xnor U10659 (N_10659,N_10439,N_10370);
and U10660 (N_10660,N_10333,N_10256);
nor U10661 (N_10661,N_10378,N_10373);
or U10662 (N_10662,N_10456,N_10264);
and U10663 (N_10663,N_10409,N_10355);
and U10664 (N_10664,N_10253,N_10421);
nand U10665 (N_10665,N_10352,N_10255);
nor U10666 (N_10666,N_10273,N_10266);
xnor U10667 (N_10667,N_10400,N_10376);
nand U10668 (N_10668,N_10433,N_10319);
or U10669 (N_10669,N_10379,N_10258);
and U10670 (N_10670,N_10446,N_10494);
and U10671 (N_10671,N_10365,N_10268);
xnor U10672 (N_10672,N_10488,N_10267);
or U10673 (N_10673,N_10310,N_10385);
nand U10674 (N_10674,N_10337,N_10356);
nor U10675 (N_10675,N_10455,N_10295);
or U10676 (N_10676,N_10368,N_10275);
nand U10677 (N_10677,N_10278,N_10450);
and U10678 (N_10678,N_10357,N_10383);
or U10679 (N_10679,N_10293,N_10384);
and U10680 (N_10680,N_10428,N_10264);
xor U10681 (N_10681,N_10386,N_10318);
nor U10682 (N_10682,N_10269,N_10346);
xor U10683 (N_10683,N_10298,N_10318);
xor U10684 (N_10684,N_10456,N_10380);
or U10685 (N_10685,N_10268,N_10374);
and U10686 (N_10686,N_10303,N_10316);
and U10687 (N_10687,N_10488,N_10327);
xnor U10688 (N_10688,N_10383,N_10271);
nand U10689 (N_10689,N_10280,N_10434);
nand U10690 (N_10690,N_10323,N_10294);
nor U10691 (N_10691,N_10450,N_10407);
or U10692 (N_10692,N_10329,N_10452);
and U10693 (N_10693,N_10301,N_10298);
and U10694 (N_10694,N_10413,N_10482);
or U10695 (N_10695,N_10489,N_10322);
or U10696 (N_10696,N_10350,N_10393);
or U10697 (N_10697,N_10463,N_10318);
nor U10698 (N_10698,N_10446,N_10426);
xnor U10699 (N_10699,N_10306,N_10335);
nor U10700 (N_10700,N_10410,N_10469);
nor U10701 (N_10701,N_10278,N_10311);
xor U10702 (N_10702,N_10479,N_10373);
nor U10703 (N_10703,N_10490,N_10465);
nor U10704 (N_10704,N_10482,N_10289);
and U10705 (N_10705,N_10291,N_10292);
nand U10706 (N_10706,N_10483,N_10408);
nor U10707 (N_10707,N_10343,N_10460);
nor U10708 (N_10708,N_10341,N_10477);
nor U10709 (N_10709,N_10436,N_10328);
xor U10710 (N_10710,N_10346,N_10470);
xor U10711 (N_10711,N_10344,N_10489);
and U10712 (N_10712,N_10442,N_10351);
and U10713 (N_10713,N_10333,N_10267);
and U10714 (N_10714,N_10281,N_10388);
or U10715 (N_10715,N_10459,N_10392);
and U10716 (N_10716,N_10290,N_10483);
nand U10717 (N_10717,N_10275,N_10258);
nor U10718 (N_10718,N_10483,N_10383);
xor U10719 (N_10719,N_10262,N_10313);
nor U10720 (N_10720,N_10449,N_10422);
nor U10721 (N_10721,N_10385,N_10362);
nor U10722 (N_10722,N_10397,N_10399);
nor U10723 (N_10723,N_10362,N_10426);
nor U10724 (N_10724,N_10397,N_10404);
xnor U10725 (N_10725,N_10305,N_10404);
or U10726 (N_10726,N_10267,N_10373);
or U10727 (N_10727,N_10422,N_10303);
xnor U10728 (N_10728,N_10287,N_10337);
nor U10729 (N_10729,N_10447,N_10269);
nor U10730 (N_10730,N_10302,N_10288);
xnor U10731 (N_10731,N_10251,N_10277);
or U10732 (N_10732,N_10286,N_10293);
or U10733 (N_10733,N_10435,N_10263);
nor U10734 (N_10734,N_10363,N_10493);
nand U10735 (N_10735,N_10454,N_10327);
or U10736 (N_10736,N_10327,N_10441);
and U10737 (N_10737,N_10313,N_10311);
xor U10738 (N_10738,N_10362,N_10434);
nand U10739 (N_10739,N_10358,N_10473);
xnor U10740 (N_10740,N_10499,N_10266);
and U10741 (N_10741,N_10265,N_10434);
nand U10742 (N_10742,N_10287,N_10256);
nor U10743 (N_10743,N_10469,N_10486);
nand U10744 (N_10744,N_10372,N_10405);
or U10745 (N_10745,N_10405,N_10440);
or U10746 (N_10746,N_10291,N_10324);
nand U10747 (N_10747,N_10414,N_10365);
nor U10748 (N_10748,N_10262,N_10351);
nor U10749 (N_10749,N_10364,N_10460);
and U10750 (N_10750,N_10554,N_10652);
and U10751 (N_10751,N_10706,N_10571);
nor U10752 (N_10752,N_10542,N_10532);
nor U10753 (N_10753,N_10665,N_10608);
nand U10754 (N_10754,N_10610,N_10513);
nand U10755 (N_10755,N_10628,N_10606);
nor U10756 (N_10756,N_10619,N_10732);
nor U10757 (N_10757,N_10599,N_10587);
nand U10758 (N_10758,N_10714,N_10537);
or U10759 (N_10759,N_10602,N_10689);
nand U10760 (N_10760,N_10720,N_10640);
or U10761 (N_10761,N_10617,N_10684);
xor U10762 (N_10762,N_10647,N_10746);
and U10763 (N_10763,N_10516,N_10653);
and U10764 (N_10764,N_10518,N_10627);
nor U10765 (N_10765,N_10728,N_10590);
nand U10766 (N_10766,N_10658,N_10510);
nor U10767 (N_10767,N_10543,N_10578);
or U10768 (N_10768,N_10663,N_10611);
nand U10769 (N_10769,N_10701,N_10592);
and U10770 (N_10770,N_10702,N_10557);
and U10771 (N_10771,N_10668,N_10679);
nor U10772 (N_10772,N_10614,N_10678);
nand U10773 (N_10773,N_10531,N_10675);
nand U10774 (N_10774,N_10593,N_10646);
nor U10775 (N_10775,N_10584,N_10677);
xor U10776 (N_10776,N_10664,N_10545);
xnor U10777 (N_10777,N_10736,N_10735);
nand U10778 (N_10778,N_10695,N_10504);
xnor U10779 (N_10779,N_10580,N_10572);
nor U10780 (N_10780,N_10670,N_10568);
nor U10781 (N_10781,N_10582,N_10644);
nand U10782 (N_10782,N_10625,N_10723);
and U10783 (N_10783,N_10729,N_10639);
nand U10784 (N_10784,N_10512,N_10747);
or U10785 (N_10785,N_10630,N_10620);
or U10786 (N_10786,N_10713,N_10674);
nor U10787 (N_10787,N_10509,N_10603);
and U10788 (N_10788,N_10525,N_10740);
nor U10789 (N_10789,N_10563,N_10676);
and U10790 (N_10790,N_10685,N_10618);
nand U10791 (N_10791,N_10503,N_10704);
xnor U10792 (N_10792,N_10624,N_10528);
or U10793 (N_10793,N_10654,N_10694);
or U10794 (N_10794,N_10530,N_10561);
or U10795 (N_10795,N_10607,N_10520);
and U10796 (N_10796,N_10626,N_10691);
xnor U10797 (N_10797,N_10718,N_10648);
xor U10798 (N_10798,N_10583,N_10562);
nor U10799 (N_10799,N_10687,N_10589);
and U10800 (N_10800,N_10699,N_10502);
or U10801 (N_10801,N_10641,N_10739);
nand U10802 (N_10802,N_10629,N_10743);
xor U10803 (N_10803,N_10662,N_10514);
and U10804 (N_10804,N_10634,N_10598);
nand U10805 (N_10805,N_10635,N_10656);
xor U10806 (N_10806,N_10738,N_10637);
or U10807 (N_10807,N_10552,N_10730);
xnor U10808 (N_10808,N_10579,N_10632);
and U10809 (N_10809,N_10708,N_10696);
or U10810 (N_10810,N_10534,N_10650);
nand U10811 (N_10811,N_10574,N_10550);
xor U10812 (N_10812,N_10709,N_10597);
and U10813 (N_10813,N_10529,N_10712);
xor U10814 (N_10814,N_10683,N_10621);
and U10815 (N_10815,N_10507,N_10692);
nor U10816 (N_10816,N_10749,N_10601);
nand U10817 (N_10817,N_10524,N_10671);
nor U10818 (N_10818,N_10716,N_10538);
nand U10819 (N_10819,N_10551,N_10501);
or U10820 (N_10820,N_10613,N_10560);
and U10821 (N_10821,N_10705,N_10657);
nor U10822 (N_10822,N_10585,N_10576);
and U10823 (N_10823,N_10544,N_10703);
xnor U10824 (N_10824,N_10500,N_10748);
xnor U10825 (N_10825,N_10725,N_10737);
or U10826 (N_10826,N_10661,N_10731);
nand U10827 (N_10827,N_10605,N_10609);
and U10828 (N_10828,N_10570,N_10642);
nor U10829 (N_10829,N_10744,N_10558);
and U10830 (N_10830,N_10564,N_10721);
or U10831 (N_10831,N_10719,N_10588);
and U10832 (N_10832,N_10565,N_10660);
nand U10833 (N_10833,N_10717,N_10726);
xor U10834 (N_10834,N_10710,N_10681);
or U10835 (N_10835,N_10535,N_10536);
nor U10836 (N_10836,N_10577,N_10553);
nor U10837 (N_10837,N_10734,N_10548);
and U10838 (N_10838,N_10547,N_10690);
nand U10839 (N_10839,N_10526,N_10700);
or U10840 (N_10840,N_10616,N_10511);
xnor U10841 (N_10841,N_10659,N_10615);
nor U10842 (N_10842,N_10680,N_10688);
xnor U10843 (N_10843,N_10612,N_10643);
xor U10844 (N_10844,N_10569,N_10581);
or U10845 (N_10845,N_10586,N_10693);
nor U10846 (N_10846,N_10655,N_10669);
xnor U10847 (N_10847,N_10645,N_10521);
nor U10848 (N_10848,N_10711,N_10631);
or U10849 (N_10849,N_10636,N_10672);
or U10850 (N_10850,N_10724,N_10697);
or U10851 (N_10851,N_10549,N_10519);
and U10852 (N_10852,N_10686,N_10666);
and U10853 (N_10853,N_10600,N_10517);
nand U10854 (N_10854,N_10596,N_10566);
or U10855 (N_10855,N_10595,N_10604);
and U10856 (N_10856,N_10523,N_10522);
nor U10857 (N_10857,N_10567,N_10673);
nand U10858 (N_10858,N_10559,N_10707);
nand U10859 (N_10859,N_10742,N_10594);
or U10860 (N_10860,N_10556,N_10527);
and U10861 (N_10861,N_10508,N_10733);
nand U10862 (N_10862,N_10540,N_10533);
or U10863 (N_10863,N_10722,N_10575);
xnor U10864 (N_10864,N_10715,N_10623);
nor U10865 (N_10865,N_10539,N_10505);
nor U10866 (N_10866,N_10741,N_10745);
and U10867 (N_10867,N_10682,N_10633);
nand U10868 (N_10868,N_10515,N_10573);
nor U10869 (N_10869,N_10649,N_10506);
nand U10870 (N_10870,N_10651,N_10555);
and U10871 (N_10871,N_10622,N_10546);
xor U10872 (N_10872,N_10541,N_10698);
or U10873 (N_10873,N_10727,N_10667);
and U10874 (N_10874,N_10638,N_10591);
xnor U10875 (N_10875,N_10610,N_10578);
xor U10876 (N_10876,N_10512,N_10705);
nor U10877 (N_10877,N_10683,N_10556);
nand U10878 (N_10878,N_10672,N_10559);
nor U10879 (N_10879,N_10678,N_10674);
and U10880 (N_10880,N_10611,N_10664);
or U10881 (N_10881,N_10577,N_10645);
nor U10882 (N_10882,N_10669,N_10611);
or U10883 (N_10883,N_10508,N_10588);
nand U10884 (N_10884,N_10743,N_10522);
xor U10885 (N_10885,N_10511,N_10591);
nor U10886 (N_10886,N_10581,N_10628);
nor U10887 (N_10887,N_10629,N_10514);
nor U10888 (N_10888,N_10685,N_10724);
nor U10889 (N_10889,N_10597,N_10580);
and U10890 (N_10890,N_10718,N_10652);
xnor U10891 (N_10891,N_10652,N_10661);
or U10892 (N_10892,N_10587,N_10682);
and U10893 (N_10893,N_10681,N_10532);
nand U10894 (N_10894,N_10547,N_10503);
and U10895 (N_10895,N_10528,N_10662);
and U10896 (N_10896,N_10726,N_10716);
nor U10897 (N_10897,N_10696,N_10615);
and U10898 (N_10898,N_10552,N_10591);
nor U10899 (N_10899,N_10678,N_10554);
nor U10900 (N_10900,N_10628,N_10549);
nor U10901 (N_10901,N_10650,N_10586);
nor U10902 (N_10902,N_10602,N_10597);
nand U10903 (N_10903,N_10605,N_10579);
xnor U10904 (N_10904,N_10653,N_10581);
nand U10905 (N_10905,N_10522,N_10624);
xor U10906 (N_10906,N_10666,N_10603);
nor U10907 (N_10907,N_10726,N_10586);
and U10908 (N_10908,N_10539,N_10547);
or U10909 (N_10909,N_10553,N_10590);
and U10910 (N_10910,N_10640,N_10556);
or U10911 (N_10911,N_10657,N_10644);
xnor U10912 (N_10912,N_10624,N_10715);
nand U10913 (N_10913,N_10730,N_10689);
nor U10914 (N_10914,N_10517,N_10513);
nand U10915 (N_10915,N_10511,N_10513);
and U10916 (N_10916,N_10512,N_10573);
xnor U10917 (N_10917,N_10725,N_10598);
nor U10918 (N_10918,N_10715,N_10565);
or U10919 (N_10919,N_10709,N_10608);
and U10920 (N_10920,N_10686,N_10659);
xor U10921 (N_10921,N_10633,N_10599);
nand U10922 (N_10922,N_10584,N_10560);
or U10923 (N_10923,N_10509,N_10519);
nor U10924 (N_10924,N_10672,N_10538);
nor U10925 (N_10925,N_10647,N_10648);
or U10926 (N_10926,N_10661,N_10686);
or U10927 (N_10927,N_10740,N_10549);
xor U10928 (N_10928,N_10622,N_10606);
xor U10929 (N_10929,N_10593,N_10651);
xor U10930 (N_10930,N_10590,N_10609);
or U10931 (N_10931,N_10571,N_10646);
and U10932 (N_10932,N_10705,N_10621);
nor U10933 (N_10933,N_10506,N_10568);
and U10934 (N_10934,N_10635,N_10741);
or U10935 (N_10935,N_10554,N_10510);
xor U10936 (N_10936,N_10660,N_10537);
and U10937 (N_10937,N_10682,N_10659);
or U10938 (N_10938,N_10593,N_10550);
nor U10939 (N_10939,N_10542,N_10688);
xor U10940 (N_10940,N_10693,N_10687);
nand U10941 (N_10941,N_10547,N_10532);
and U10942 (N_10942,N_10579,N_10633);
xor U10943 (N_10943,N_10554,N_10649);
nor U10944 (N_10944,N_10519,N_10561);
nor U10945 (N_10945,N_10609,N_10604);
or U10946 (N_10946,N_10594,N_10527);
xor U10947 (N_10947,N_10535,N_10587);
nand U10948 (N_10948,N_10727,N_10589);
xnor U10949 (N_10949,N_10601,N_10525);
nor U10950 (N_10950,N_10727,N_10641);
xor U10951 (N_10951,N_10691,N_10593);
or U10952 (N_10952,N_10509,N_10540);
nor U10953 (N_10953,N_10551,N_10645);
or U10954 (N_10954,N_10537,N_10711);
and U10955 (N_10955,N_10741,N_10500);
or U10956 (N_10956,N_10503,N_10689);
xor U10957 (N_10957,N_10638,N_10648);
or U10958 (N_10958,N_10608,N_10586);
nand U10959 (N_10959,N_10525,N_10747);
xor U10960 (N_10960,N_10592,N_10713);
or U10961 (N_10961,N_10594,N_10562);
or U10962 (N_10962,N_10644,N_10687);
nor U10963 (N_10963,N_10575,N_10645);
nor U10964 (N_10964,N_10571,N_10620);
nor U10965 (N_10965,N_10590,N_10679);
xor U10966 (N_10966,N_10523,N_10660);
nand U10967 (N_10967,N_10600,N_10513);
xor U10968 (N_10968,N_10675,N_10737);
and U10969 (N_10969,N_10535,N_10633);
xnor U10970 (N_10970,N_10609,N_10696);
nor U10971 (N_10971,N_10722,N_10669);
or U10972 (N_10972,N_10673,N_10624);
xnor U10973 (N_10973,N_10511,N_10572);
nor U10974 (N_10974,N_10664,N_10728);
or U10975 (N_10975,N_10688,N_10702);
nand U10976 (N_10976,N_10589,N_10717);
and U10977 (N_10977,N_10697,N_10620);
and U10978 (N_10978,N_10630,N_10624);
and U10979 (N_10979,N_10689,N_10659);
and U10980 (N_10980,N_10642,N_10646);
xor U10981 (N_10981,N_10619,N_10585);
and U10982 (N_10982,N_10652,N_10665);
nor U10983 (N_10983,N_10714,N_10511);
xor U10984 (N_10984,N_10572,N_10724);
and U10985 (N_10985,N_10644,N_10515);
and U10986 (N_10986,N_10728,N_10627);
nor U10987 (N_10987,N_10629,N_10699);
xor U10988 (N_10988,N_10581,N_10544);
nor U10989 (N_10989,N_10605,N_10547);
nor U10990 (N_10990,N_10745,N_10744);
nor U10991 (N_10991,N_10506,N_10685);
nor U10992 (N_10992,N_10548,N_10635);
and U10993 (N_10993,N_10538,N_10549);
and U10994 (N_10994,N_10534,N_10595);
or U10995 (N_10995,N_10647,N_10722);
and U10996 (N_10996,N_10743,N_10649);
nor U10997 (N_10997,N_10710,N_10612);
or U10998 (N_10998,N_10615,N_10581);
nor U10999 (N_10999,N_10734,N_10528);
and U11000 (N_11000,N_10881,N_10794);
nand U11001 (N_11001,N_10854,N_10954);
nor U11002 (N_11002,N_10896,N_10962);
nand U11003 (N_11003,N_10792,N_10762);
nor U11004 (N_11004,N_10936,N_10877);
or U11005 (N_11005,N_10917,N_10947);
nand U11006 (N_11006,N_10949,N_10829);
xnor U11007 (N_11007,N_10933,N_10946);
or U11008 (N_11008,N_10822,N_10959);
and U11009 (N_11009,N_10860,N_10826);
and U11010 (N_11010,N_10913,N_10892);
nor U11011 (N_11011,N_10978,N_10943);
xor U11012 (N_11012,N_10890,N_10845);
and U11013 (N_11013,N_10793,N_10920);
nor U11014 (N_11014,N_10931,N_10873);
or U11015 (N_11015,N_10850,N_10998);
nor U11016 (N_11016,N_10895,N_10758);
xnor U11017 (N_11017,N_10889,N_10825);
xnor U11018 (N_11018,N_10948,N_10904);
nand U11019 (N_11019,N_10790,N_10884);
nand U11020 (N_11020,N_10880,N_10862);
or U11021 (N_11021,N_10966,N_10769);
and U11022 (N_11022,N_10839,N_10777);
nand U11023 (N_11023,N_10971,N_10874);
xor U11024 (N_11024,N_10765,N_10926);
xnor U11025 (N_11025,N_10914,N_10941);
xor U11026 (N_11026,N_10784,N_10972);
nand U11027 (N_11027,N_10841,N_10887);
or U11028 (N_11028,N_10870,N_10852);
or U11029 (N_11029,N_10849,N_10940);
nor U11030 (N_11030,N_10879,N_10886);
nor U11031 (N_11031,N_10857,N_10897);
nand U11032 (N_11032,N_10844,N_10900);
nor U11033 (N_11033,N_10859,N_10950);
or U11034 (N_11034,N_10967,N_10867);
nand U11035 (N_11035,N_10778,N_10970);
nand U11036 (N_11036,N_10842,N_10754);
or U11037 (N_11037,N_10816,N_10922);
xor U11038 (N_11038,N_10830,N_10837);
or U11039 (N_11039,N_10773,N_10770);
or U11040 (N_11040,N_10819,N_10969);
nand U11041 (N_11041,N_10851,N_10760);
nor U11042 (N_11042,N_10802,N_10958);
and U11043 (N_11043,N_10985,N_10963);
nor U11044 (N_11044,N_10811,N_10994);
and U11045 (N_11045,N_10975,N_10891);
xnor U11046 (N_11046,N_10813,N_10983);
nand U11047 (N_11047,N_10903,N_10810);
xnor U11048 (N_11048,N_10861,N_10821);
xnor U11049 (N_11049,N_10905,N_10751);
xor U11050 (N_11050,N_10907,N_10836);
or U11051 (N_11051,N_10757,N_10952);
nand U11052 (N_11052,N_10981,N_10753);
nor U11053 (N_11053,N_10806,N_10800);
and U11054 (N_11054,N_10803,N_10853);
xnor U11055 (N_11055,N_10894,N_10768);
nand U11056 (N_11056,N_10875,N_10902);
xor U11057 (N_11057,N_10766,N_10865);
and U11058 (N_11058,N_10910,N_10866);
nor U11059 (N_11059,N_10820,N_10782);
and U11060 (N_11060,N_10957,N_10964);
and U11061 (N_11061,N_10937,N_10997);
or U11062 (N_11062,N_10763,N_10847);
or U11063 (N_11063,N_10840,N_10797);
and U11064 (N_11064,N_10786,N_10974);
xnor U11065 (N_11065,N_10814,N_10955);
nand U11066 (N_11066,N_10973,N_10961);
nor U11067 (N_11067,N_10752,N_10930);
and U11068 (N_11068,N_10883,N_10750);
or U11069 (N_11069,N_10918,N_10838);
or U11070 (N_11070,N_10855,N_10827);
xnor U11071 (N_11071,N_10796,N_10858);
xor U11072 (N_11072,N_10869,N_10764);
nand U11073 (N_11073,N_10927,N_10756);
and U11074 (N_11074,N_10771,N_10992);
nor U11075 (N_11075,N_10824,N_10808);
or U11076 (N_11076,N_10901,N_10831);
nor U11077 (N_11077,N_10779,N_10988);
and U11078 (N_11078,N_10834,N_10801);
or U11079 (N_11079,N_10888,N_10864);
nor U11080 (N_11080,N_10939,N_10965);
or U11081 (N_11081,N_10921,N_10899);
xor U11082 (N_11082,N_10893,N_10906);
or U11083 (N_11083,N_10916,N_10924);
nor U11084 (N_11084,N_10987,N_10791);
xor U11085 (N_11085,N_10795,N_10925);
or U11086 (N_11086,N_10909,N_10938);
or U11087 (N_11087,N_10799,N_10761);
nand U11088 (N_11088,N_10772,N_10809);
xnor U11089 (N_11089,N_10928,N_10929);
nand U11090 (N_11090,N_10977,N_10976);
and U11091 (N_11091,N_10817,N_10812);
or U11092 (N_11092,N_10856,N_10908);
nand U11093 (N_11093,N_10953,N_10984);
xor U11094 (N_11094,N_10815,N_10934);
or U11095 (N_11095,N_10876,N_10923);
or U11096 (N_11096,N_10807,N_10911);
nand U11097 (N_11097,N_10878,N_10781);
and U11098 (N_11098,N_10805,N_10833);
nor U11099 (N_11099,N_10995,N_10956);
nand U11100 (N_11100,N_10789,N_10755);
or U11101 (N_11101,N_10775,N_10783);
xnor U11102 (N_11102,N_10871,N_10898);
xnor U11103 (N_11103,N_10882,N_10787);
nor U11104 (N_11104,N_10776,N_10863);
xnor U11105 (N_11105,N_10990,N_10986);
and U11106 (N_11106,N_10804,N_10935);
nor U11107 (N_11107,N_10991,N_10980);
and U11108 (N_11108,N_10996,N_10872);
and U11109 (N_11109,N_10912,N_10848);
nor U11110 (N_11110,N_10835,N_10785);
or U11111 (N_11111,N_10828,N_10885);
nor U11112 (N_11112,N_10942,N_10774);
xnor U11113 (N_11113,N_10982,N_10951);
nor U11114 (N_11114,N_10989,N_10818);
xor U11115 (N_11115,N_10999,N_10932);
or U11116 (N_11116,N_10868,N_10919);
xnor U11117 (N_11117,N_10915,N_10788);
or U11118 (N_11118,N_10968,N_10780);
and U11119 (N_11119,N_10960,N_10979);
and U11120 (N_11120,N_10832,N_10823);
and U11121 (N_11121,N_10759,N_10767);
nand U11122 (N_11122,N_10944,N_10798);
nand U11123 (N_11123,N_10993,N_10945);
xnor U11124 (N_11124,N_10846,N_10843);
and U11125 (N_11125,N_10768,N_10906);
xnor U11126 (N_11126,N_10943,N_10936);
and U11127 (N_11127,N_10832,N_10841);
or U11128 (N_11128,N_10869,N_10997);
or U11129 (N_11129,N_10895,N_10984);
xnor U11130 (N_11130,N_10873,N_10970);
xor U11131 (N_11131,N_10986,N_10887);
nand U11132 (N_11132,N_10849,N_10897);
and U11133 (N_11133,N_10781,N_10901);
nand U11134 (N_11134,N_10888,N_10919);
xnor U11135 (N_11135,N_10823,N_10879);
nor U11136 (N_11136,N_10766,N_10925);
xnor U11137 (N_11137,N_10982,N_10816);
and U11138 (N_11138,N_10897,N_10881);
or U11139 (N_11139,N_10894,N_10904);
nor U11140 (N_11140,N_10936,N_10871);
or U11141 (N_11141,N_10872,N_10975);
xnor U11142 (N_11142,N_10817,N_10768);
and U11143 (N_11143,N_10810,N_10984);
or U11144 (N_11144,N_10945,N_10997);
or U11145 (N_11145,N_10819,N_10897);
and U11146 (N_11146,N_10793,N_10869);
xnor U11147 (N_11147,N_10798,N_10843);
nor U11148 (N_11148,N_10751,N_10798);
nand U11149 (N_11149,N_10891,N_10912);
or U11150 (N_11150,N_10917,N_10836);
nand U11151 (N_11151,N_10863,N_10814);
nor U11152 (N_11152,N_10967,N_10794);
nand U11153 (N_11153,N_10839,N_10934);
nand U11154 (N_11154,N_10777,N_10794);
nor U11155 (N_11155,N_10962,N_10853);
and U11156 (N_11156,N_10854,N_10924);
xor U11157 (N_11157,N_10772,N_10995);
or U11158 (N_11158,N_10892,N_10881);
nand U11159 (N_11159,N_10788,N_10882);
xnor U11160 (N_11160,N_10965,N_10926);
and U11161 (N_11161,N_10902,N_10849);
nor U11162 (N_11162,N_10755,N_10832);
nor U11163 (N_11163,N_10988,N_10751);
and U11164 (N_11164,N_10973,N_10928);
xnor U11165 (N_11165,N_10762,N_10805);
nor U11166 (N_11166,N_10990,N_10927);
xor U11167 (N_11167,N_10944,N_10786);
or U11168 (N_11168,N_10809,N_10752);
xor U11169 (N_11169,N_10910,N_10796);
nor U11170 (N_11170,N_10870,N_10768);
nor U11171 (N_11171,N_10852,N_10864);
xor U11172 (N_11172,N_10756,N_10879);
or U11173 (N_11173,N_10801,N_10918);
nor U11174 (N_11174,N_10996,N_10895);
xor U11175 (N_11175,N_10857,N_10800);
and U11176 (N_11176,N_10848,N_10763);
or U11177 (N_11177,N_10847,N_10907);
and U11178 (N_11178,N_10757,N_10901);
or U11179 (N_11179,N_10819,N_10866);
and U11180 (N_11180,N_10995,N_10969);
nand U11181 (N_11181,N_10873,N_10781);
xor U11182 (N_11182,N_10770,N_10870);
nor U11183 (N_11183,N_10977,N_10863);
nor U11184 (N_11184,N_10827,N_10864);
xnor U11185 (N_11185,N_10877,N_10993);
or U11186 (N_11186,N_10990,N_10829);
or U11187 (N_11187,N_10776,N_10864);
nor U11188 (N_11188,N_10917,N_10940);
and U11189 (N_11189,N_10871,N_10887);
xor U11190 (N_11190,N_10868,N_10832);
nand U11191 (N_11191,N_10984,N_10891);
or U11192 (N_11192,N_10953,N_10877);
and U11193 (N_11193,N_10857,N_10828);
and U11194 (N_11194,N_10931,N_10851);
xor U11195 (N_11195,N_10991,N_10909);
nand U11196 (N_11196,N_10988,N_10827);
and U11197 (N_11197,N_10925,N_10880);
nand U11198 (N_11198,N_10826,N_10955);
xor U11199 (N_11199,N_10888,N_10818);
nor U11200 (N_11200,N_10861,N_10769);
xor U11201 (N_11201,N_10900,N_10888);
or U11202 (N_11202,N_10949,N_10792);
nand U11203 (N_11203,N_10807,N_10904);
and U11204 (N_11204,N_10847,N_10829);
or U11205 (N_11205,N_10768,N_10991);
nor U11206 (N_11206,N_10945,N_10835);
or U11207 (N_11207,N_10979,N_10992);
or U11208 (N_11208,N_10950,N_10873);
xor U11209 (N_11209,N_10782,N_10948);
nand U11210 (N_11210,N_10986,N_10781);
and U11211 (N_11211,N_10754,N_10782);
and U11212 (N_11212,N_10780,N_10758);
and U11213 (N_11213,N_10952,N_10940);
nor U11214 (N_11214,N_10780,N_10914);
and U11215 (N_11215,N_10773,N_10880);
xnor U11216 (N_11216,N_10860,N_10963);
nor U11217 (N_11217,N_10965,N_10770);
or U11218 (N_11218,N_10985,N_10752);
nor U11219 (N_11219,N_10801,N_10764);
and U11220 (N_11220,N_10869,N_10941);
and U11221 (N_11221,N_10888,N_10763);
xor U11222 (N_11222,N_10877,N_10797);
xnor U11223 (N_11223,N_10985,N_10822);
xnor U11224 (N_11224,N_10942,N_10908);
xnor U11225 (N_11225,N_10795,N_10950);
and U11226 (N_11226,N_10835,N_10858);
or U11227 (N_11227,N_10899,N_10803);
xnor U11228 (N_11228,N_10862,N_10870);
xor U11229 (N_11229,N_10897,N_10951);
nand U11230 (N_11230,N_10863,N_10942);
nand U11231 (N_11231,N_10889,N_10892);
xor U11232 (N_11232,N_10762,N_10876);
or U11233 (N_11233,N_10902,N_10893);
or U11234 (N_11234,N_10834,N_10896);
nor U11235 (N_11235,N_10907,N_10909);
xnor U11236 (N_11236,N_10796,N_10760);
nand U11237 (N_11237,N_10876,N_10777);
and U11238 (N_11238,N_10937,N_10946);
and U11239 (N_11239,N_10787,N_10876);
xor U11240 (N_11240,N_10970,N_10972);
and U11241 (N_11241,N_10782,N_10943);
xor U11242 (N_11242,N_10954,N_10893);
or U11243 (N_11243,N_10794,N_10773);
or U11244 (N_11244,N_10845,N_10842);
and U11245 (N_11245,N_10918,N_10839);
xor U11246 (N_11246,N_10919,N_10971);
nor U11247 (N_11247,N_10829,N_10885);
and U11248 (N_11248,N_10899,N_10839);
and U11249 (N_11249,N_10908,N_10891);
nand U11250 (N_11250,N_11223,N_11138);
nor U11251 (N_11251,N_11193,N_11143);
and U11252 (N_11252,N_11000,N_11236);
or U11253 (N_11253,N_11038,N_11210);
nor U11254 (N_11254,N_11001,N_11114);
xnor U11255 (N_11255,N_11002,N_11183);
nand U11256 (N_11256,N_11207,N_11046);
xor U11257 (N_11257,N_11135,N_11106);
nor U11258 (N_11258,N_11028,N_11240);
xor U11259 (N_11259,N_11241,N_11045);
nand U11260 (N_11260,N_11129,N_11168);
and U11261 (N_11261,N_11147,N_11057);
xnor U11262 (N_11262,N_11111,N_11093);
xnor U11263 (N_11263,N_11101,N_11026);
xor U11264 (N_11264,N_11072,N_11204);
xnor U11265 (N_11265,N_11234,N_11062);
xor U11266 (N_11266,N_11044,N_11120);
and U11267 (N_11267,N_11095,N_11167);
and U11268 (N_11268,N_11119,N_11176);
xor U11269 (N_11269,N_11148,N_11018);
nand U11270 (N_11270,N_11125,N_11209);
or U11271 (N_11271,N_11079,N_11075);
xor U11272 (N_11272,N_11034,N_11212);
nor U11273 (N_11273,N_11071,N_11218);
nand U11274 (N_11274,N_11011,N_11203);
nor U11275 (N_11275,N_11144,N_11151);
or U11276 (N_11276,N_11134,N_11246);
nor U11277 (N_11277,N_11105,N_11030);
nor U11278 (N_11278,N_11098,N_11088);
nor U11279 (N_11279,N_11213,N_11050);
and U11280 (N_11280,N_11237,N_11006);
and U11281 (N_11281,N_11199,N_11021);
nor U11282 (N_11282,N_11235,N_11163);
nor U11283 (N_11283,N_11007,N_11200);
and U11284 (N_11284,N_11003,N_11153);
nand U11285 (N_11285,N_11226,N_11152);
nand U11286 (N_11286,N_11103,N_11113);
nand U11287 (N_11287,N_11159,N_11078);
nor U11288 (N_11288,N_11086,N_11208);
nand U11289 (N_11289,N_11109,N_11197);
xor U11290 (N_11290,N_11162,N_11224);
and U11291 (N_11291,N_11054,N_11025);
and U11292 (N_11292,N_11172,N_11191);
or U11293 (N_11293,N_11137,N_11222);
xnor U11294 (N_11294,N_11139,N_11177);
or U11295 (N_11295,N_11067,N_11126);
nand U11296 (N_11296,N_11090,N_11189);
and U11297 (N_11297,N_11190,N_11037);
and U11298 (N_11298,N_11042,N_11115);
nand U11299 (N_11299,N_11085,N_11205);
xor U11300 (N_11300,N_11158,N_11082);
or U11301 (N_11301,N_11013,N_11225);
nand U11302 (N_11302,N_11108,N_11080);
nand U11303 (N_11303,N_11227,N_11027);
and U11304 (N_11304,N_11121,N_11211);
and U11305 (N_11305,N_11175,N_11130);
and U11306 (N_11306,N_11228,N_11160);
nor U11307 (N_11307,N_11060,N_11084);
nand U11308 (N_11308,N_11039,N_11171);
nand U11309 (N_11309,N_11174,N_11049);
xnor U11310 (N_11310,N_11068,N_11184);
and U11311 (N_11311,N_11052,N_11077);
or U11312 (N_11312,N_11219,N_11186);
nor U11313 (N_11313,N_11179,N_11102);
xor U11314 (N_11314,N_11055,N_11248);
nor U11315 (N_11315,N_11117,N_11024);
nor U11316 (N_11316,N_11194,N_11047);
nor U11317 (N_11317,N_11136,N_11201);
and U11318 (N_11318,N_11048,N_11074);
nor U11319 (N_11319,N_11229,N_11061);
nor U11320 (N_11320,N_11231,N_11112);
or U11321 (N_11321,N_11032,N_11036);
and U11322 (N_11322,N_11009,N_11244);
nand U11323 (N_11323,N_11118,N_11022);
and U11324 (N_11324,N_11107,N_11065);
or U11325 (N_11325,N_11169,N_11249);
xnor U11326 (N_11326,N_11041,N_11012);
nor U11327 (N_11327,N_11170,N_11245);
nor U11328 (N_11328,N_11202,N_11031);
nand U11329 (N_11329,N_11097,N_11239);
xnor U11330 (N_11330,N_11164,N_11221);
xnor U11331 (N_11331,N_11188,N_11166);
xor U11332 (N_11332,N_11220,N_11215);
xnor U11333 (N_11333,N_11232,N_11216);
nand U11334 (N_11334,N_11096,N_11073);
xor U11335 (N_11335,N_11247,N_11142);
nor U11336 (N_11336,N_11092,N_11059);
or U11337 (N_11337,N_11217,N_11081);
nand U11338 (N_11338,N_11141,N_11015);
nand U11339 (N_11339,N_11178,N_11035);
or U11340 (N_11340,N_11242,N_11127);
nand U11341 (N_11341,N_11233,N_11058);
xnor U11342 (N_11342,N_11033,N_11091);
and U11343 (N_11343,N_11198,N_11070);
nand U11344 (N_11344,N_11110,N_11182);
xnor U11345 (N_11345,N_11150,N_11100);
xnor U11346 (N_11346,N_11243,N_11083);
nand U11347 (N_11347,N_11195,N_11131);
and U11348 (N_11348,N_11149,N_11023);
and U11349 (N_11349,N_11017,N_11066);
nand U11350 (N_11350,N_11155,N_11192);
nand U11351 (N_11351,N_11056,N_11128);
nor U11352 (N_11352,N_11206,N_11099);
and U11353 (N_11353,N_11094,N_11187);
and U11354 (N_11354,N_11087,N_11064);
and U11355 (N_11355,N_11063,N_11069);
xnor U11356 (N_11356,N_11019,N_11076);
nand U11357 (N_11357,N_11145,N_11230);
nand U11358 (N_11358,N_11005,N_11053);
and U11359 (N_11359,N_11161,N_11156);
xnor U11360 (N_11360,N_11185,N_11180);
and U11361 (N_11361,N_11008,N_11123);
nor U11362 (N_11362,N_11165,N_11004);
and U11363 (N_11363,N_11116,N_11010);
xnor U11364 (N_11364,N_11089,N_11133);
nand U11365 (N_11365,N_11043,N_11181);
or U11366 (N_11366,N_11238,N_11029);
xor U11367 (N_11367,N_11173,N_11196);
xor U11368 (N_11368,N_11140,N_11124);
or U11369 (N_11369,N_11014,N_11051);
or U11370 (N_11370,N_11020,N_11122);
and U11371 (N_11371,N_11016,N_11104);
nor U11372 (N_11372,N_11040,N_11146);
nor U11373 (N_11373,N_11214,N_11154);
or U11374 (N_11374,N_11157,N_11132);
or U11375 (N_11375,N_11149,N_11032);
or U11376 (N_11376,N_11146,N_11030);
xnor U11377 (N_11377,N_11175,N_11086);
xnor U11378 (N_11378,N_11144,N_11173);
xor U11379 (N_11379,N_11157,N_11142);
nor U11380 (N_11380,N_11015,N_11173);
nor U11381 (N_11381,N_11082,N_11220);
xor U11382 (N_11382,N_11031,N_11231);
xnor U11383 (N_11383,N_11210,N_11244);
or U11384 (N_11384,N_11175,N_11080);
xnor U11385 (N_11385,N_11187,N_11080);
and U11386 (N_11386,N_11173,N_11241);
nand U11387 (N_11387,N_11232,N_11075);
nand U11388 (N_11388,N_11125,N_11158);
xor U11389 (N_11389,N_11126,N_11009);
xnor U11390 (N_11390,N_11089,N_11222);
nand U11391 (N_11391,N_11070,N_11109);
and U11392 (N_11392,N_11143,N_11058);
nand U11393 (N_11393,N_11046,N_11023);
nand U11394 (N_11394,N_11189,N_11249);
nand U11395 (N_11395,N_11079,N_11193);
and U11396 (N_11396,N_11161,N_11045);
nor U11397 (N_11397,N_11128,N_11130);
xor U11398 (N_11398,N_11214,N_11036);
and U11399 (N_11399,N_11152,N_11039);
or U11400 (N_11400,N_11221,N_11030);
nor U11401 (N_11401,N_11115,N_11160);
nand U11402 (N_11402,N_11227,N_11088);
xnor U11403 (N_11403,N_11052,N_11144);
xnor U11404 (N_11404,N_11112,N_11061);
xor U11405 (N_11405,N_11066,N_11096);
nand U11406 (N_11406,N_11129,N_11149);
nor U11407 (N_11407,N_11130,N_11197);
nand U11408 (N_11408,N_11036,N_11169);
xnor U11409 (N_11409,N_11131,N_11219);
and U11410 (N_11410,N_11107,N_11028);
nand U11411 (N_11411,N_11211,N_11238);
nand U11412 (N_11412,N_11155,N_11112);
nand U11413 (N_11413,N_11228,N_11126);
nor U11414 (N_11414,N_11216,N_11080);
nand U11415 (N_11415,N_11130,N_11042);
nand U11416 (N_11416,N_11143,N_11180);
and U11417 (N_11417,N_11096,N_11189);
or U11418 (N_11418,N_11158,N_11195);
nor U11419 (N_11419,N_11101,N_11139);
xor U11420 (N_11420,N_11212,N_11201);
or U11421 (N_11421,N_11247,N_11170);
or U11422 (N_11422,N_11080,N_11090);
and U11423 (N_11423,N_11023,N_11218);
xnor U11424 (N_11424,N_11138,N_11038);
xor U11425 (N_11425,N_11218,N_11030);
nor U11426 (N_11426,N_11152,N_11041);
nor U11427 (N_11427,N_11047,N_11069);
and U11428 (N_11428,N_11059,N_11235);
nand U11429 (N_11429,N_11091,N_11029);
nor U11430 (N_11430,N_11209,N_11193);
nand U11431 (N_11431,N_11163,N_11069);
nand U11432 (N_11432,N_11071,N_11126);
nand U11433 (N_11433,N_11157,N_11208);
nor U11434 (N_11434,N_11098,N_11123);
xor U11435 (N_11435,N_11031,N_11131);
nand U11436 (N_11436,N_11220,N_11186);
or U11437 (N_11437,N_11171,N_11036);
nand U11438 (N_11438,N_11101,N_11035);
or U11439 (N_11439,N_11200,N_11242);
nand U11440 (N_11440,N_11176,N_11223);
or U11441 (N_11441,N_11089,N_11163);
or U11442 (N_11442,N_11001,N_11045);
nor U11443 (N_11443,N_11071,N_11099);
and U11444 (N_11444,N_11175,N_11169);
nor U11445 (N_11445,N_11225,N_11114);
xor U11446 (N_11446,N_11014,N_11171);
xor U11447 (N_11447,N_11073,N_11024);
and U11448 (N_11448,N_11183,N_11101);
xnor U11449 (N_11449,N_11027,N_11084);
or U11450 (N_11450,N_11047,N_11113);
and U11451 (N_11451,N_11110,N_11061);
nand U11452 (N_11452,N_11014,N_11186);
nor U11453 (N_11453,N_11153,N_11218);
or U11454 (N_11454,N_11122,N_11246);
nand U11455 (N_11455,N_11118,N_11171);
or U11456 (N_11456,N_11052,N_11128);
nand U11457 (N_11457,N_11091,N_11022);
or U11458 (N_11458,N_11232,N_11163);
or U11459 (N_11459,N_11055,N_11053);
xnor U11460 (N_11460,N_11218,N_11183);
or U11461 (N_11461,N_11047,N_11167);
xnor U11462 (N_11462,N_11016,N_11105);
nand U11463 (N_11463,N_11217,N_11029);
xnor U11464 (N_11464,N_11210,N_11097);
nor U11465 (N_11465,N_11200,N_11089);
nand U11466 (N_11466,N_11040,N_11241);
nor U11467 (N_11467,N_11121,N_11200);
and U11468 (N_11468,N_11242,N_11216);
xnor U11469 (N_11469,N_11183,N_11217);
xnor U11470 (N_11470,N_11101,N_11042);
nand U11471 (N_11471,N_11217,N_11244);
or U11472 (N_11472,N_11097,N_11187);
nand U11473 (N_11473,N_11162,N_11121);
nor U11474 (N_11474,N_11222,N_11086);
nand U11475 (N_11475,N_11074,N_11093);
nor U11476 (N_11476,N_11026,N_11243);
xor U11477 (N_11477,N_11091,N_11131);
nor U11478 (N_11478,N_11009,N_11003);
nand U11479 (N_11479,N_11165,N_11143);
and U11480 (N_11480,N_11135,N_11178);
or U11481 (N_11481,N_11008,N_11067);
nand U11482 (N_11482,N_11134,N_11234);
nand U11483 (N_11483,N_11014,N_11129);
nand U11484 (N_11484,N_11216,N_11206);
nor U11485 (N_11485,N_11202,N_11234);
nand U11486 (N_11486,N_11060,N_11070);
or U11487 (N_11487,N_11011,N_11127);
xor U11488 (N_11488,N_11030,N_11188);
or U11489 (N_11489,N_11158,N_11193);
xor U11490 (N_11490,N_11211,N_11093);
and U11491 (N_11491,N_11081,N_11045);
nand U11492 (N_11492,N_11005,N_11088);
and U11493 (N_11493,N_11133,N_11064);
xnor U11494 (N_11494,N_11117,N_11246);
xor U11495 (N_11495,N_11104,N_11217);
or U11496 (N_11496,N_11151,N_11046);
nor U11497 (N_11497,N_11034,N_11118);
xnor U11498 (N_11498,N_11183,N_11233);
nand U11499 (N_11499,N_11179,N_11205);
or U11500 (N_11500,N_11433,N_11380);
xnor U11501 (N_11501,N_11352,N_11441);
or U11502 (N_11502,N_11260,N_11421);
nand U11503 (N_11503,N_11342,N_11474);
and U11504 (N_11504,N_11486,N_11489);
xnor U11505 (N_11505,N_11458,N_11387);
nor U11506 (N_11506,N_11481,N_11468);
and U11507 (N_11507,N_11268,N_11417);
or U11508 (N_11508,N_11425,N_11343);
or U11509 (N_11509,N_11294,N_11412);
or U11510 (N_11510,N_11375,N_11404);
nand U11511 (N_11511,N_11272,N_11482);
nand U11512 (N_11512,N_11393,N_11477);
xor U11513 (N_11513,N_11469,N_11357);
nor U11514 (N_11514,N_11490,N_11324);
and U11515 (N_11515,N_11478,N_11471);
or U11516 (N_11516,N_11407,N_11367);
or U11517 (N_11517,N_11312,N_11472);
or U11518 (N_11518,N_11399,N_11310);
and U11519 (N_11519,N_11303,N_11498);
nand U11520 (N_11520,N_11492,N_11320);
and U11521 (N_11521,N_11276,N_11374);
or U11522 (N_11522,N_11302,N_11361);
or U11523 (N_11523,N_11423,N_11385);
nand U11524 (N_11524,N_11456,N_11292);
or U11525 (N_11525,N_11463,N_11484);
and U11526 (N_11526,N_11304,N_11392);
or U11527 (N_11527,N_11327,N_11345);
and U11528 (N_11528,N_11325,N_11265);
nor U11529 (N_11529,N_11358,N_11460);
nor U11530 (N_11530,N_11445,N_11452);
or U11531 (N_11531,N_11283,N_11255);
nand U11532 (N_11532,N_11400,N_11443);
nand U11533 (N_11533,N_11317,N_11410);
and U11534 (N_11534,N_11328,N_11348);
nand U11535 (N_11535,N_11363,N_11279);
or U11536 (N_11536,N_11377,N_11473);
and U11537 (N_11537,N_11493,N_11497);
nand U11538 (N_11538,N_11290,N_11395);
or U11539 (N_11539,N_11495,N_11251);
nor U11540 (N_11540,N_11259,N_11419);
and U11541 (N_11541,N_11379,N_11288);
nand U11542 (N_11542,N_11281,N_11470);
nor U11543 (N_11543,N_11381,N_11416);
or U11544 (N_11544,N_11293,N_11346);
nor U11545 (N_11545,N_11262,N_11261);
or U11546 (N_11546,N_11275,N_11439);
nand U11547 (N_11547,N_11326,N_11321);
or U11548 (N_11548,N_11313,N_11355);
and U11549 (N_11549,N_11431,N_11284);
or U11550 (N_11550,N_11384,N_11306);
nand U11551 (N_11551,N_11333,N_11368);
xor U11552 (N_11552,N_11397,N_11365);
xnor U11553 (N_11553,N_11285,N_11301);
and U11554 (N_11554,N_11323,N_11453);
nor U11555 (N_11555,N_11450,N_11273);
and U11556 (N_11556,N_11447,N_11388);
nand U11557 (N_11557,N_11252,N_11315);
or U11558 (N_11558,N_11394,N_11319);
nand U11559 (N_11559,N_11396,N_11370);
nand U11560 (N_11560,N_11341,N_11455);
xnor U11561 (N_11561,N_11349,N_11257);
nor U11562 (N_11562,N_11408,N_11295);
nand U11563 (N_11563,N_11389,N_11267);
nor U11564 (N_11564,N_11274,N_11369);
nor U11565 (N_11565,N_11351,N_11464);
nand U11566 (N_11566,N_11411,N_11483);
and U11567 (N_11567,N_11364,N_11401);
nand U11568 (N_11568,N_11308,N_11434);
or U11569 (N_11569,N_11436,N_11475);
xnor U11570 (N_11570,N_11496,N_11253);
xnor U11571 (N_11571,N_11428,N_11413);
and U11572 (N_11572,N_11378,N_11376);
or U11573 (N_11573,N_11422,N_11296);
nand U11574 (N_11574,N_11430,N_11494);
xnor U11575 (N_11575,N_11485,N_11332);
xnor U11576 (N_11576,N_11347,N_11476);
xor U11577 (N_11577,N_11353,N_11479);
and U11578 (N_11578,N_11289,N_11491);
or U11579 (N_11579,N_11286,N_11318);
or U11580 (N_11580,N_11454,N_11264);
nor U11581 (N_11581,N_11311,N_11403);
and U11582 (N_11582,N_11287,N_11373);
or U11583 (N_11583,N_11465,N_11405);
xnor U11584 (N_11584,N_11444,N_11258);
nand U11585 (N_11585,N_11386,N_11338);
nand U11586 (N_11586,N_11330,N_11406);
xor U11587 (N_11587,N_11309,N_11339);
or U11588 (N_11588,N_11440,N_11442);
nand U11589 (N_11589,N_11427,N_11305);
nor U11590 (N_11590,N_11329,N_11383);
nand U11591 (N_11591,N_11266,N_11402);
or U11592 (N_11592,N_11340,N_11270);
nand U11593 (N_11593,N_11344,N_11390);
or U11594 (N_11594,N_11446,N_11414);
nor U11595 (N_11595,N_11278,N_11356);
nor U11596 (N_11596,N_11398,N_11371);
or U11597 (N_11597,N_11300,N_11331);
or U11598 (N_11598,N_11466,N_11337);
and U11599 (N_11599,N_11280,N_11437);
or U11600 (N_11600,N_11409,N_11256);
nand U11601 (N_11601,N_11282,N_11366);
nor U11602 (N_11602,N_11354,N_11435);
or U11603 (N_11603,N_11487,N_11336);
xnor U11604 (N_11604,N_11499,N_11415);
or U11605 (N_11605,N_11271,N_11254);
and U11606 (N_11606,N_11480,N_11307);
or U11607 (N_11607,N_11350,N_11359);
and U11608 (N_11608,N_11438,N_11277);
nand U11609 (N_11609,N_11297,N_11314);
nor U11610 (N_11610,N_11372,N_11462);
or U11611 (N_11611,N_11457,N_11459);
nand U11612 (N_11612,N_11420,N_11426);
or U11613 (N_11613,N_11432,N_11488);
xor U11614 (N_11614,N_11448,N_11316);
or U11615 (N_11615,N_11291,N_11461);
and U11616 (N_11616,N_11263,N_11449);
xor U11617 (N_11617,N_11429,N_11424);
xnor U11618 (N_11618,N_11269,N_11334);
nor U11619 (N_11619,N_11250,N_11451);
or U11620 (N_11620,N_11418,N_11322);
xnor U11621 (N_11621,N_11391,N_11362);
and U11622 (N_11622,N_11382,N_11299);
nor U11623 (N_11623,N_11335,N_11298);
or U11624 (N_11624,N_11467,N_11360);
xnor U11625 (N_11625,N_11335,N_11385);
xor U11626 (N_11626,N_11279,N_11372);
and U11627 (N_11627,N_11475,N_11442);
nor U11628 (N_11628,N_11346,N_11492);
nor U11629 (N_11629,N_11453,N_11484);
or U11630 (N_11630,N_11298,N_11364);
xnor U11631 (N_11631,N_11387,N_11279);
nand U11632 (N_11632,N_11376,N_11415);
nor U11633 (N_11633,N_11304,N_11311);
nor U11634 (N_11634,N_11454,N_11416);
xor U11635 (N_11635,N_11336,N_11298);
or U11636 (N_11636,N_11261,N_11376);
or U11637 (N_11637,N_11333,N_11311);
or U11638 (N_11638,N_11417,N_11494);
and U11639 (N_11639,N_11420,N_11458);
or U11640 (N_11640,N_11447,N_11334);
and U11641 (N_11641,N_11452,N_11344);
and U11642 (N_11642,N_11361,N_11468);
xor U11643 (N_11643,N_11486,N_11336);
xor U11644 (N_11644,N_11370,N_11454);
nor U11645 (N_11645,N_11494,N_11294);
or U11646 (N_11646,N_11426,N_11356);
nor U11647 (N_11647,N_11440,N_11425);
nand U11648 (N_11648,N_11479,N_11497);
xor U11649 (N_11649,N_11357,N_11254);
xnor U11650 (N_11650,N_11435,N_11449);
nor U11651 (N_11651,N_11316,N_11484);
and U11652 (N_11652,N_11394,N_11430);
or U11653 (N_11653,N_11414,N_11265);
and U11654 (N_11654,N_11492,N_11285);
or U11655 (N_11655,N_11425,N_11429);
and U11656 (N_11656,N_11376,N_11267);
or U11657 (N_11657,N_11323,N_11311);
xnor U11658 (N_11658,N_11404,N_11303);
nor U11659 (N_11659,N_11300,N_11466);
xor U11660 (N_11660,N_11450,N_11434);
nor U11661 (N_11661,N_11455,N_11447);
and U11662 (N_11662,N_11449,N_11317);
or U11663 (N_11663,N_11434,N_11359);
and U11664 (N_11664,N_11358,N_11307);
xnor U11665 (N_11665,N_11285,N_11372);
xor U11666 (N_11666,N_11428,N_11363);
and U11667 (N_11667,N_11416,N_11483);
and U11668 (N_11668,N_11441,N_11486);
nand U11669 (N_11669,N_11395,N_11408);
and U11670 (N_11670,N_11415,N_11482);
xor U11671 (N_11671,N_11477,N_11362);
or U11672 (N_11672,N_11397,N_11375);
and U11673 (N_11673,N_11393,N_11269);
xor U11674 (N_11674,N_11404,N_11357);
nor U11675 (N_11675,N_11256,N_11267);
nand U11676 (N_11676,N_11414,N_11447);
xnor U11677 (N_11677,N_11480,N_11300);
xnor U11678 (N_11678,N_11452,N_11314);
or U11679 (N_11679,N_11408,N_11454);
xnor U11680 (N_11680,N_11499,N_11481);
nand U11681 (N_11681,N_11361,N_11301);
or U11682 (N_11682,N_11427,N_11316);
xor U11683 (N_11683,N_11282,N_11477);
or U11684 (N_11684,N_11361,N_11469);
xor U11685 (N_11685,N_11463,N_11475);
nor U11686 (N_11686,N_11378,N_11253);
nor U11687 (N_11687,N_11373,N_11296);
nand U11688 (N_11688,N_11279,N_11350);
and U11689 (N_11689,N_11308,N_11440);
xnor U11690 (N_11690,N_11413,N_11400);
xor U11691 (N_11691,N_11378,N_11331);
or U11692 (N_11692,N_11333,N_11428);
or U11693 (N_11693,N_11358,N_11278);
xor U11694 (N_11694,N_11446,N_11309);
nor U11695 (N_11695,N_11440,N_11465);
or U11696 (N_11696,N_11433,N_11374);
and U11697 (N_11697,N_11275,N_11488);
xnor U11698 (N_11698,N_11263,N_11327);
nand U11699 (N_11699,N_11315,N_11351);
nand U11700 (N_11700,N_11275,N_11443);
nand U11701 (N_11701,N_11384,N_11307);
nor U11702 (N_11702,N_11477,N_11442);
xor U11703 (N_11703,N_11391,N_11329);
xor U11704 (N_11704,N_11327,N_11389);
xor U11705 (N_11705,N_11407,N_11419);
and U11706 (N_11706,N_11380,N_11359);
nor U11707 (N_11707,N_11258,N_11472);
or U11708 (N_11708,N_11446,N_11397);
nor U11709 (N_11709,N_11286,N_11469);
or U11710 (N_11710,N_11454,N_11262);
and U11711 (N_11711,N_11405,N_11404);
xor U11712 (N_11712,N_11370,N_11430);
nor U11713 (N_11713,N_11464,N_11431);
nor U11714 (N_11714,N_11358,N_11426);
or U11715 (N_11715,N_11482,N_11369);
and U11716 (N_11716,N_11302,N_11458);
and U11717 (N_11717,N_11464,N_11403);
nand U11718 (N_11718,N_11293,N_11480);
or U11719 (N_11719,N_11348,N_11252);
nor U11720 (N_11720,N_11294,N_11468);
xor U11721 (N_11721,N_11481,N_11448);
xnor U11722 (N_11722,N_11316,N_11463);
xor U11723 (N_11723,N_11435,N_11397);
nand U11724 (N_11724,N_11267,N_11384);
and U11725 (N_11725,N_11363,N_11383);
and U11726 (N_11726,N_11448,N_11257);
nand U11727 (N_11727,N_11411,N_11336);
xor U11728 (N_11728,N_11377,N_11318);
nor U11729 (N_11729,N_11341,N_11449);
and U11730 (N_11730,N_11315,N_11477);
or U11731 (N_11731,N_11269,N_11490);
xnor U11732 (N_11732,N_11311,N_11301);
nand U11733 (N_11733,N_11271,N_11354);
nor U11734 (N_11734,N_11276,N_11492);
xor U11735 (N_11735,N_11380,N_11332);
or U11736 (N_11736,N_11451,N_11370);
nor U11737 (N_11737,N_11411,N_11361);
nor U11738 (N_11738,N_11405,N_11302);
and U11739 (N_11739,N_11354,N_11251);
and U11740 (N_11740,N_11253,N_11293);
and U11741 (N_11741,N_11402,N_11313);
or U11742 (N_11742,N_11476,N_11286);
nand U11743 (N_11743,N_11297,N_11313);
nand U11744 (N_11744,N_11337,N_11491);
nand U11745 (N_11745,N_11254,N_11312);
and U11746 (N_11746,N_11344,N_11341);
and U11747 (N_11747,N_11434,N_11494);
nand U11748 (N_11748,N_11455,N_11420);
nand U11749 (N_11749,N_11290,N_11265);
nor U11750 (N_11750,N_11735,N_11518);
and U11751 (N_11751,N_11733,N_11720);
nand U11752 (N_11752,N_11551,N_11749);
and U11753 (N_11753,N_11724,N_11536);
and U11754 (N_11754,N_11538,N_11646);
nand U11755 (N_11755,N_11700,N_11615);
or U11756 (N_11756,N_11734,N_11689);
and U11757 (N_11757,N_11731,N_11699);
nor U11758 (N_11758,N_11544,N_11514);
or U11759 (N_11759,N_11533,N_11708);
and U11760 (N_11760,N_11509,N_11523);
nor U11761 (N_11761,N_11541,N_11529);
and U11762 (N_11762,N_11578,N_11637);
nand U11763 (N_11763,N_11717,N_11694);
xnor U11764 (N_11764,N_11555,N_11569);
and U11765 (N_11765,N_11547,N_11704);
and U11766 (N_11766,N_11613,N_11664);
xor U11767 (N_11767,N_11622,N_11573);
xnor U11768 (N_11768,N_11586,N_11617);
or U11769 (N_11769,N_11603,N_11675);
nand U11770 (N_11770,N_11517,N_11621);
and U11771 (N_11771,N_11527,N_11552);
or U11772 (N_11772,N_11743,N_11680);
nand U11773 (N_11773,N_11587,N_11530);
nand U11774 (N_11774,N_11737,N_11686);
nand U11775 (N_11775,N_11625,N_11643);
nand U11776 (N_11776,N_11607,N_11581);
or U11777 (N_11777,N_11685,N_11719);
nor U11778 (N_11778,N_11744,N_11508);
nor U11779 (N_11779,N_11515,N_11653);
xnor U11780 (N_11780,N_11666,N_11672);
nor U11781 (N_11781,N_11549,N_11504);
nor U11782 (N_11782,N_11542,N_11678);
nor U11783 (N_11783,N_11559,N_11725);
and U11784 (N_11784,N_11568,N_11683);
and U11785 (N_11785,N_11526,N_11674);
xor U11786 (N_11786,N_11532,N_11682);
nor U11787 (N_11787,N_11701,N_11618);
nor U11788 (N_11788,N_11679,N_11612);
xnor U11789 (N_11789,N_11534,N_11535);
nor U11790 (N_11790,N_11567,N_11747);
xnor U11791 (N_11791,N_11673,N_11563);
nor U11792 (N_11792,N_11654,N_11626);
xor U11793 (N_11793,N_11642,N_11669);
and U11794 (N_11794,N_11597,N_11740);
nand U11795 (N_11795,N_11553,N_11606);
xor U11796 (N_11796,N_11600,N_11506);
or U11797 (N_11797,N_11565,N_11690);
nor U11798 (N_11798,N_11714,N_11732);
nor U11799 (N_11799,N_11507,N_11636);
and U11800 (N_11800,N_11648,N_11630);
nand U11801 (N_11801,N_11608,N_11710);
xor U11802 (N_11802,N_11566,N_11705);
and U11803 (N_11803,N_11539,N_11665);
nor U11804 (N_11804,N_11645,N_11579);
or U11805 (N_11805,N_11564,N_11575);
nand U11806 (N_11806,N_11592,N_11543);
nor U11807 (N_11807,N_11571,N_11545);
or U11808 (N_11808,N_11531,N_11659);
nand U11809 (N_11809,N_11623,N_11624);
nor U11810 (N_11810,N_11687,N_11519);
and U11811 (N_11811,N_11677,N_11512);
xor U11812 (N_11812,N_11745,N_11524);
and U11813 (N_11813,N_11639,N_11616);
nand U11814 (N_11814,N_11596,N_11729);
and U11815 (N_11815,N_11620,N_11604);
nor U11816 (N_11816,N_11660,N_11663);
nor U11817 (N_11817,N_11667,N_11510);
nor U11818 (N_11818,N_11649,N_11550);
nor U11819 (N_11819,N_11580,N_11684);
nand U11820 (N_11820,N_11501,N_11525);
nor U11821 (N_11821,N_11676,N_11562);
or U11822 (N_11822,N_11528,N_11582);
and U11823 (N_11823,N_11556,N_11650);
nor U11824 (N_11824,N_11598,N_11560);
and U11825 (N_11825,N_11726,N_11632);
nor U11826 (N_11826,N_11634,N_11748);
nand U11827 (N_11827,N_11697,N_11671);
or U11828 (N_11828,N_11712,N_11576);
and U11829 (N_11829,N_11554,N_11703);
nand U11830 (N_11830,N_11584,N_11670);
nand U11831 (N_11831,N_11537,N_11591);
nand U11832 (N_11832,N_11658,N_11691);
nor U11833 (N_11833,N_11656,N_11721);
xor U11834 (N_11834,N_11513,N_11692);
or U11835 (N_11835,N_11502,N_11594);
nor U11836 (N_11836,N_11601,N_11570);
nor U11837 (N_11837,N_11695,N_11651);
nand U11838 (N_11838,N_11681,N_11593);
or U11839 (N_11839,N_11709,N_11500);
xnor U11840 (N_11840,N_11698,N_11718);
nand U11841 (N_11841,N_11711,N_11572);
or U11842 (N_11842,N_11561,N_11589);
xnor U11843 (N_11843,N_11611,N_11557);
nor U11844 (N_11844,N_11657,N_11610);
and U11845 (N_11845,N_11595,N_11574);
or U11846 (N_11846,N_11590,N_11702);
nand U11847 (N_11847,N_11738,N_11605);
nand U11848 (N_11848,N_11521,N_11707);
nor U11849 (N_11849,N_11614,N_11722);
nor U11850 (N_11850,N_11736,N_11585);
nand U11851 (N_11851,N_11540,N_11548);
xnor U11852 (N_11852,N_11742,N_11602);
nor U11853 (N_11853,N_11588,N_11713);
xor U11854 (N_11854,N_11696,N_11520);
nor U11855 (N_11855,N_11688,N_11629);
and U11856 (N_11856,N_11640,N_11716);
xnor U11857 (N_11857,N_11728,N_11638);
nor U11858 (N_11858,N_11693,N_11635);
or U11859 (N_11859,N_11641,N_11583);
and U11860 (N_11860,N_11746,N_11730);
nor U11861 (N_11861,N_11727,N_11662);
xor U11862 (N_11862,N_11516,N_11609);
nor U11863 (N_11863,N_11661,N_11644);
and U11864 (N_11864,N_11723,N_11652);
and U11865 (N_11865,N_11505,N_11706);
and U11866 (N_11866,N_11558,N_11577);
xnor U11867 (N_11867,N_11633,N_11628);
nand U11868 (N_11868,N_11599,N_11619);
or U11869 (N_11869,N_11546,N_11511);
nor U11870 (N_11870,N_11668,N_11627);
nand U11871 (N_11871,N_11739,N_11631);
nor U11872 (N_11872,N_11522,N_11647);
nor U11873 (N_11873,N_11655,N_11715);
xor U11874 (N_11874,N_11503,N_11741);
nor U11875 (N_11875,N_11554,N_11714);
nor U11876 (N_11876,N_11519,N_11666);
xor U11877 (N_11877,N_11545,N_11636);
xor U11878 (N_11878,N_11734,N_11627);
or U11879 (N_11879,N_11690,N_11714);
and U11880 (N_11880,N_11737,N_11536);
and U11881 (N_11881,N_11527,N_11674);
or U11882 (N_11882,N_11519,N_11538);
xnor U11883 (N_11883,N_11718,N_11630);
nor U11884 (N_11884,N_11531,N_11564);
xnor U11885 (N_11885,N_11646,N_11708);
or U11886 (N_11886,N_11507,N_11586);
nor U11887 (N_11887,N_11564,N_11580);
xor U11888 (N_11888,N_11635,N_11580);
and U11889 (N_11889,N_11697,N_11662);
and U11890 (N_11890,N_11744,N_11728);
nor U11891 (N_11891,N_11575,N_11510);
and U11892 (N_11892,N_11572,N_11582);
nand U11893 (N_11893,N_11613,N_11687);
nor U11894 (N_11894,N_11675,N_11614);
xor U11895 (N_11895,N_11545,N_11556);
and U11896 (N_11896,N_11706,N_11541);
nand U11897 (N_11897,N_11541,N_11547);
xnor U11898 (N_11898,N_11608,N_11736);
and U11899 (N_11899,N_11629,N_11696);
or U11900 (N_11900,N_11657,N_11668);
xnor U11901 (N_11901,N_11532,N_11626);
nor U11902 (N_11902,N_11640,N_11517);
and U11903 (N_11903,N_11570,N_11600);
nand U11904 (N_11904,N_11737,N_11544);
or U11905 (N_11905,N_11544,N_11602);
xnor U11906 (N_11906,N_11560,N_11554);
nor U11907 (N_11907,N_11605,N_11640);
and U11908 (N_11908,N_11727,N_11578);
nor U11909 (N_11909,N_11581,N_11512);
and U11910 (N_11910,N_11503,N_11556);
xor U11911 (N_11911,N_11688,N_11630);
xnor U11912 (N_11912,N_11529,N_11692);
nand U11913 (N_11913,N_11662,N_11576);
nor U11914 (N_11914,N_11684,N_11623);
or U11915 (N_11915,N_11670,N_11518);
nand U11916 (N_11916,N_11696,N_11740);
or U11917 (N_11917,N_11629,N_11611);
nand U11918 (N_11918,N_11616,N_11641);
xor U11919 (N_11919,N_11718,N_11578);
nand U11920 (N_11920,N_11715,N_11520);
or U11921 (N_11921,N_11648,N_11611);
xor U11922 (N_11922,N_11590,N_11500);
or U11923 (N_11923,N_11580,N_11555);
or U11924 (N_11924,N_11535,N_11566);
xor U11925 (N_11925,N_11640,N_11731);
nor U11926 (N_11926,N_11575,N_11603);
nand U11927 (N_11927,N_11664,N_11591);
or U11928 (N_11928,N_11636,N_11599);
and U11929 (N_11929,N_11539,N_11537);
and U11930 (N_11930,N_11719,N_11623);
or U11931 (N_11931,N_11650,N_11745);
or U11932 (N_11932,N_11513,N_11609);
nor U11933 (N_11933,N_11687,N_11502);
nor U11934 (N_11934,N_11720,N_11607);
xnor U11935 (N_11935,N_11727,N_11643);
nor U11936 (N_11936,N_11506,N_11515);
and U11937 (N_11937,N_11656,N_11629);
and U11938 (N_11938,N_11536,N_11681);
or U11939 (N_11939,N_11646,N_11649);
nand U11940 (N_11940,N_11610,N_11749);
nand U11941 (N_11941,N_11547,N_11743);
nor U11942 (N_11942,N_11613,N_11525);
nor U11943 (N_11943,N_11719,N_11588);
nor U11944 (N_11944,N_11697,N_11547);
and U11945 (N_11945,N_11741,N_11749);
and U11946 (N_11946,N_11573,N_11720);
nor U11947 (N_11947,N_11608,N_11552);
xnor U11948 (N_11948,N_11715,N_11697);
nand U11949 (N_11949,N_11567,N_11568);
or U11950 (N_11950,N_11519,N_11516);
nand U11951 (N_11951,N_11583,N_11598);
nand U11952 (N_11952,N_11682,N_11533);
and U11953 (N_11953,N_11658,N_11569);
xnor U11954 (N_11954,N_11648,N_11536);
or U11955 (N_11955,N_11735,N_11714);
nor U11956 (N_11956,N_11668,N_11590);
and U11957 (N_11957,N_11728,N_11583);
and U11958 (N_11958,N_11604,N_11627);
or U11959 (N_11959,N_11505,N_11569);
xnor U11960 (N_11960,N_11594,N_11685);
or U11961 (N_11961,N_11720,N_11600);
nor U11962 (N_11962,N_11674,N_11513);
or U11963 (N_11963,N_11602,N_11540);
or U11964 (N_11964,N_11604,N_11602);
or U11965 (N_11965,N_11744,N_11543);
or U11966 (N_11966,N_11612,N_11649);
or U11967 (N_11967,N_11683,N_11534);
nor U11968 (N_11968,N_11590,N_11605);
xnor U11969 (N_11969,N_11604,N_11623);
nand U11970 (N_11970,N_11578,N_11674);
xnor U11971 (N_11971,N_11710,N_11624);
xor U11972 (N_11972,N_11699,N_11611);
nor U11973 (N_11973,N_11631,N_11658);
xor U11974 (N_11974,N_11513,N_11650);
or U11975 (N_11975,N_11674,N_11701);
xor U11976 (N_11976,N_11615,N_11588);
xor U11977 (N_11977,N_11599,N_11561);
and U11978 (N_11978,N_11651,N_11504);
nand U11979 (N_11979,N_11740,N_11572);
nor U11980 (N_11980,N_11509,N_11525);
nor U11981 (N_11981,N_11627,N_11597);
or U11982 (N_11982,N_11592,N_11586);
xnor U11983 (N_11983,N_11521,N_11675);
nor U11984 (N_11984,N_11717,N_11500);
xor U11985 (N_11985,N_11582,N_11658);
nand U11986 (N_11986,N_11544,N_11523);
or U11987 (N_11987,N_11665,N_11520);
xnor U11988 (N_11988,N_11546,N_11674);
and U11989 (N_11989,N_11589,N_11566);
and U11990 (N_11990,N_11652,N_11510);
or U11991 (N_11991,N_11735,N_11542);
and U11992 (N_11992,N_11579,N_11664);
nand U11993 (N_11993,N_11716,N_11643);
xor U11994 (N_11994,N_11544,N_11669);
and U11995 (N_11995,N_11633,N_11666);
xnor U11996 (N_11996,N_11633,N_11630);
nor U11997 (N_11997,N_11742,N_11705);
nand U11998 (N_11998,N_11673,N_11735);
nor U11999 (N_11999,N_11657,N_11721);
and U12000 (N_12000,N_11782,N_11837);
nand U12001 (N_12001,N_11868,N_11791);
xor U12002 (N_12002,N_11917,N_11806);
nor U12003 (N_12003,N_11983,N_11894);
nor U12004 (N_12004,N_11967,N_11816);
or U12005 (N_12005,N_11803,N_11956);
nor U12006 (N_12006,N_11990,N_11788);
and U12007 (N_12007,N_11986,N_11857);
and U12008 (N_12008,N_11954,N_11909);
or U12009 (N_12009,N_11766,N_11854);
and U12010 (N_12010,N_11943,N_11913);
or U12011 (N_12011,N_11940,N_11760);
or U12012 (N_12012,N_11807,N_11959);
nor U12013 (N_12013,N_11982,N_11910);
xor U12014 (N_12014,N_11793,N_11865);
nor U12015 (N_12015,N_11796,N_11885);
nand U12016 (N_12016,N_11897,N_11970);
xnor U12017 (N_12017,N_11753,N_11921);
or U12018 (N_12018,N_11767,N_11955);
xnor U12019 (N_12019,N_11991,N_11972);
or U12020 (N_12020,N_11929,N_11805);
and U12021 (N_12021,N_11935,N_11808);
nand U12022 (N_12022,N_11864,N_11814);
nor U12023 (N_12023,N_11930,N_11876);
nand U12024 (N_12024,N_11751,N_11764);
or U12025 (N_12025,N_11965,N_11998);
nand U12026 (N_12026,N_11984,N_11755);
xor U12027 (N_12027,N_11780,N_11877);
xnor U12028 (N_12028,N_11922,N_11896);
or U12029 (N_12029,N_11810,N_11925);
or U12030 (N_12030,N_11999,N_11989);
or U12031 (N_12031,N_11895,N_11971);
or U12032 (N_12032,N_11939,N_11825);
nand U12033 (N_12033,N_11773,N_11919);
xnor U12034 (N_12034,N_11833,N_11846);
or U12035 (N_12035,N_11996,N_11976);
xnor U12036 (N_12036,N_11756,N_11867);
and U12037 (N_12037,N_11856,N_11951);
nand U12038 (N_12038,N_11884,N_11878);
nand U12039 (N_12039,N_11941,N_11928);
xnor U12040 (N_12040,N_11774,N_11916);
or U12041 (N_12041,N_11824,N_11750);
or U12042 (N_12042,N_11900,N_11823);
and U12043 (N_12043,N_11860,N_11995);
or U12044 (N_12044,N_11792,N_11781);
xnor U12045 (N_12045,N_11934,N_11835);
nor U12046 (N_12046,N_11847,N_11786);
nor U12047 (N_12047,N_11849,N_11830);
or U12048 (N_12048,N_11875,N_11890);
xnor U12049 (N_12049,N_11777,N_11831);
or U12050 (N_12050,N_11827,N_11820);
nand U12051 (N_12051,N_11889,N_11992);
xnor U12052 (N_12052,N_11765,N_11985);
nor U12053 (N_12053,N_11947,N_11794);
nor U12054 (N_12054,N_11839,N_11844);
xor U12055 (N_12055,N_11855,N_11845);
xnor U12056 (N_12056,N_11953,N_11871);
xor U12057 (N_12057,N_11759,N_11787);
and U12058 (N_12058,N_11872,N_11969);
nor U12059 (N_12059,N_11933,N_11988);
nand U12060 (N_12060,N_11838,N_11874);
nand U12061 (N_12061,N_11906,N_11901);
nand U12062 (N_12062,N_11804,N_11822);
or U12063 (N_12063,N_11932,N_11973);
and U12064 (N_12064,N_11752,N_11904);
or U12065 (N_12065,N_11945,N_11800);
nor U12066 (N_12066,N_11873,N_11938);
or U12067 (N_12067,N_11836,N_11776);
or U12068 (N_12068,N_11797,N_11802);
and U12069 (N_12069,N_11757,N_11961);
nor U12070 (N_12070,N_11888,N_11966);
xor U12071 (N_12071,N_11798,N_11936);
nor U12072 (N_12072,N_11908,N_11819);
and U12073 (N_12073,N_11975,N_11758);
or U12074 (N_12074,N_11881,N_11974);
xor U12075 (N_12075,N_11812,N_11911);
nand U12076 (N_12076,N_11914,N_11891);
and U12077 (N_12077,N_11903,N_11958);
nor U12078 (N_12078,N_11858,N_11851);
nor U12079 (N_12079,N_11769,N_11841);
and U12080 (N_12080,N_11987,N_11946);
xor U12081 (N_12081,N_11840,N_11862);
and U12082 (N_12082,N_11863,N_11815);
nand U12083 (N_12083,N_11772,N_11784);
xor U12084 (N_12084,N_11892,N_11866);
or U12085 (N_12085,N_11937,N_11801);
xnor U12086 (N_12086,N_11942,N_11981);
nor U12087 (N_12087,N_11869,N_11926);
nand U12088 (N_12088,N_11950,N_11918);
nor U12089 (N_12089,N_11994,N_11795);
nand U12090 (N_12090,N_11962,N_11754);
xor U12091 (N_12091,N_11993,N_11809);
or U12092 (N_12092,N_11898,N_11915);
nor U12093 (N_12093,N_11924,N_11770);
nand U12094 (N_12094,N_11887,N_11775);
xor U12095 (N_12095,N_11850,N_11880);
or U12096 (N_12096,N_11963,N_11978);
xnor U12097 (N_12097,N_11960,N_11861);
nand U12098 (N_12098,N_11859,N_11902);
xor U12099 (N_12099,N_11848,N_11785);
nor U12100 (N_12100,N_11979,N_11944);
nor U12101 (N_12101,N_11927,N_11879);
nor U12102 (N_12102,N_11842,N_11852);
or U12103 (N_12103,N_11843,N_11952);
or U12104 (N_12104,N_11826,N_11893);
and U12105 (N_12105,N_11907,N_11968);
xor U12106 (N_12106,N_11870,N_11771);
xor U12107 (N_12107,N_11763,N_11923);
nor U12108 (N_12108,N_11828,N_11980);
xnor U12109 (N_12109,N_11905,N_11949);
xor U12110 (N_12110,N_11899,N_11997);
nand U12111 (N_12111,N_11778,N_11957);
and U12112 (N_12112,N_11761,N_11948);
nor U12113 (N_12113,N_11799,N_11811);
and U12114 (N_12114,N_11768,N_11783);
nand U12115 (N_12115,N_11813,N_11883);
nor U12116 (N_12116,N_11834,N_11964);
nand U12117 (N_12117,N_11886,N_11818);
or U12118 (N_12118,N_11829,N_11779);
nor U12119 (N_12119,N_11931,N_11920);
and U12120 (N_12120,N_11882,N_11832);
or U12121 (N_12121,N_11762,N_11912);
nor U12122 (N_12122,N_11853,N_11790);
nor U12123 (N_12123,N_11977,N_11817);
and U12124 (N_12124,N_11821,N_11789);
and U12125 (N_12125,N_11896,N_11843);
nand U12126 (N_12126,N_11965,N_11890);
and U12127 (N_12127,N_11890,N_11994);
xnor U12128 (N_12128,N_11843,N_11902);
xor U12129 (N_12129,N_11978,N_11831);
nand U12130 (N_12130,N_11987,N_11956);
and U12131 (N_12131,N_11807,N_11980);
nand U12132 (N_12132,N_11891,N_11878);
and U12133 (N_12133,N_11907,N_11870);
nand U12134 (N_12134,N_11823,N_11763);
or U12135 (N_12135,N_11760,N_11827);
or U12136 (N_12136,N_11923,N_11788);
or U12137 (N_12137,N_11807,N_11844);
nor U12138 (N_12138,N_11889,N_11753);
xor U12139 (N_12139,N_11999,N_11911);
nand U12140 (N_12140,N_11812,N_11750);
nor U12141 (N_12141,N_11949,N_11934);
nand U12142 (N_12142,N_11997,N_11874);
or U12143 (N_12143,N_11898,N_11999);
xor U12144 (N_12144,N_11961,N_11824);
and U12145 (N_12145,N_11972,N_11797);
or U12146 (N_12146,N_11994,N_11985);
or U12147 (N_12147,N_11918,N_11986);
and U12148 (N_12148,N_11810,N_11821);
xor U12149 (N_12149,N_11949,N_11939);
nand U12150 (N_12150,N_11926,N_11867);
and U12151 (N_12151,N_11896,N_11965);
nor U12152 (N_12152,N_11829,N_11992);
nand U12153 (N_12153,N_11998,N_11932);
or U12154 (N_12154,N_11928,N_11824);
nand U12155 (N_12155,N_11969,N_11795);
xor U12156 (N_12156,N_11956,N_11783);
nand U12157 (N_12157,N_11782,N_11829);
xor U12158 (N_12158,N_11834,N_11909);
or U12159 (N_12159,N_11792,N_11944);
or U12160 (N_12160,N_11833,N_11781);
and U12161 (N_12161,N_11978,N_11905);
and U12162 (N_12162,N_11816,N_11785);
xor U12163 (N_12163,N_11998,N_11988);
and U12164 (N_12164,N_11938,N_11998);
nand U12165 (N_12165,N_11940,N_11865);
nand U12166 (N_12166,N_11884,N_11871);
xnor U12167 (N_12167,N_11969,N_11805);
and U12168 (N_12168,N_11820,N_11783);
nand U12169 (N_12169,N_11923,N_11881);
xnor U12170 (N_12170,N_11907,N_11928);
or U12171 (N_12171,N_11924,N_11962);
xor U12172 (N_12172,N_11801,N_11999);
nand U12173 (N_12173,N_11787,N_11958);
xnor U12174 (N_12174,N_11867,N_11911);
nor U12175 (N_12175,N_11898,N_11899);
or U12176 (N_12176,N_11913,N_11778);
nor U12177 (N_12177,N_11929,N_11980);
nor U12178 (N_12178,N_11910,N_11761);
xor U12179 (N_12179,N_11870,N_11866);
and U12180 (N_12180,N_11939,N_11919);
nand U12181 (N_12181,N_11982,N_11913);
nand U12182 (N_12182,N_11990,N_11951);
or U12183 (N_12183,N_11844,N_11867);
or U12184 (N_12184,N_11862,N_11916);
or U12185 (N_12185,N_11928,N_11829);
xnor U12186 (N_12186,N_11967,N_11887);
and U12187 (N_12187,N_11859,N_11825);
xor U12188 (N_12188,N_11813,N_11854);
xor U12189 (N_12189,N_11831,N_11865);
nand U12190 (N_12190,N_11761,N_11836);
nor U12191 (N_12191,N_11904,N_11922);
nand U12192 (N_12192,N_11946,N_11849);
and U12193 (N_12193,N_11997,N_11952);
and U12194 (N_12194,N_11896,N_11892);
xnor U12195 (N_12195,N_11810,N_11853);
xnor U12196 (N_12196,N_11769,N_11891);
xnor U12197 (N_12197,N_11884,N_11897);
and U12198 (N_12198,N_11893,N_11945);
nand U12199 (N_12199,N_11894,N_11848);
xnor U12200 (N_12200,N_11856,N_11913);
nor U12201 (N_12201,N_11776,N_11970);
nand U12202 (N_12202,N_11869,N_11771);
and U12203 (N_12203,N_11923,N_11928);
nor U12204 (N_12204,N_11805,N_11760);
or U12205 (N_12205,N_11812,N_11795);
or U12206 (N_12206,N_11913,N_11758);
nand U12207 (N_12207,N_11835,N_11873);
or U12208 (N_12208,N_11951,N_11978);
nand U12209 (N_12209,N_11904,N_11841);
and U12210 (N_12210,N_11948,N_11951);
nand U12211 (N_12211,N_11767,N_11980);
nor U12212 (N_12212,N_11909,N_11875);
nor U12213 (N_12213,N_11922,N_11769);
nand U12214 (N_12214,N_11797,N_11937);
nor U12215 (N_12215,N_11874,N_11804);
xor U12216 (N_12216,N_11925,N_11877);
nand U12217 (N_12217,N_11955,N_11853);
nand U12218 (N_12218,N_11879,N_11988);
nand U12219 (N_12219,N_11845,N_11853);
nand U12220 (N_12220,N_11806,N_11908);
nand U12221 (N_12221,N_11911,N_11929);
or U12222 (N_12222,N_11876,N_11823);
and U12223 (N_12223,N_11909,N_11904);
nor U12224 (N_12224,N_11921,N_11825);
nand U12225 (N_12225,N_11857,N_11917);
nor U12226 (N_12226,N_11984,N_11871);
xor U12227 (N_12227,N_11789,N_11973);
nor U12228 (N_12228,N_11968,N_11803);
nand U12229 (N_12229,N_11807,N_11875);
or U12230 (N_12230,N_11851,N_11934);
xor U12231 (N_12231,N_11912,N_11807);
xnor U12232 (N_12232,N_11876,N_11971);
nor U12233 (N_12233,N_11856,N_11800);
and U12234 (N_12234,N_11930,N_11977);
nor U12235 (N_12235,N_11770,N_11869);
nor U12236 (N_12236,N_11932,N_11888);
xor U12237 (N_12237,N_11937,N_11932);
nand U12238 (N_12238,N_11807,N_11866);
or U12239 (N_12239,N_11819,N_11954);
nand U12240 (N_12240,N_11843,N_11873);
nor U12241 (N_12241,N_11951,N_11782);
nor U12242 (N_12242,N_11964,N_11777);
nor U12243 (N_12243,N_11969,N_11830);
and U12244 (N_12244,N_11783,N_11799);
or U12245 (N_12245,N_11896,N_11800);
nand U12246 (N_12246,N_11950,N_11817);
nor U12247 (N_12247,N_11978,N_11853);
xnor U12248 (N_12248,N_11843,N_11799);
and U12249 (N_12249,N_11818,N_11985);
or U12250 (N_12250,N_12153,N_12051);
nor U12251 (N_12251,N_12031,N_12045);
nor U12252 (N_12252,N_12210,N_12213);
and U12253 (N_12253,N_12234,N_12196);
and U12254 (N_12254,N_12131,N_12172);
nand U12255 (N_12255,N_12165,N_12025);
and U12256 (N_12256,N_12109,N_12097);
or U12257 (N_12257,N_12104,N_12102);
nand U12258 (N_12258,N_12168,N_12059);
nand U12259 (N_12259,N_12065,N_12143);
nor U12260 (N_12260,N_12159,N_12164);
nand U12261 (N_12261,N_12005,N_12001);
nor U12262 (N_12262,N_12007,N_12145);
nor U12263 (N_12263,N_12207,N_12082);
and U12264 (N_12264,N_12119,N_12042);
nor U12265 (N_12265,N_12011,N_12003);
or U12266 (N_12266,N_12105,N_12053);
and U12267 (N_12267,N_12130,N_12189);
or U12268 (N_12268,N_12066,N_12044);
nand U12269 (N_12269,N_12106,N_12112);
nor U12270 (N_12270,N_12133,N_12089);
and U12271 (N_12271,N_12081,N_12160);
or U12272 (N_12272,N_12030,N_12014);
nor U12273 (N_12273,N_12010,N_12077);
nand U12274 (N_12274,N_12099,N_12079);
or U12275 (N_12275,N_12046,N_12058);
and U12276 (N_12276,N_12080,N_12071);
and U12277 (N_12277,N_12166,N_12035);
xor U12278 (N_12278,N_12138,N_12220);
nand U12279 (N_12279,N_12236,N_12180);
nor U12280 (N_12280,N_12027,N_12154);
xor U12281 (N_12281,N_12094,N_12199);
nor U12282 (N_12282,N_12039,N_12101);
and U12283 (N_12283,N_12016,N_12232);
or U12284 (N_12284,N_12052,N_12125);
xnor U12285 (N_12285,N_12040,N_12090);
nand U12286 (N_12286,N_12239,N_12151);
xor U12287 (N_12287,N_12198,N_12224);
nor U12288 (N_12288,N_12201,N_12078);
nor U12289 (N_12289,N_12150,N_12216);
and U12290 (N_12290,N_12017,N_12068);
nand U12291 (N_12291,N_12074,N_12032);
or U12292 (N_12292,N_12048,N_12121);
and U12293 (N_12293,N_12137,N_12136);
xor U12294 (N_12294,N_12120,N_12229);
nand U12295 (N_12295,N_12200,N_12211);
xnor U12296 (N_12296,N_12194,N_12186);
nor U12297 (N_12297,N_12061,N_12047);
nor U12298 (N_12298,N_12233,N_12206);
xor U12299 (N_12299,N_12100,N_12161);
or U12300 (N_12300,N_12242,N_12113);
nand U12301 (N_12301,N_12029,N_12069);
nand U12302 (N_12302,N_12240,N_12221);
nor U12303 (N_12303,N_12009,N_12249);
xor U12304 (N_12304,N_12086,N_12049);
nand U12305 (N_12305,N_12050,N_12245);
and U12306 (N_12306,N_12013,N_12162);
xnor U12307 (N_12307,N_12054,N_12037);
xnor U12308 (N_12308,N_12181,N_12212);
nor U12309 (N_12309,N_12067,N_12070);
nand U12310 (N_12310,N_12190,N_12148);
nand U12311 (N_12311,N_12149,N_12177);
nor U12312 (N_12312,N_12191,N_12020);
and U12313 (N_12313,N_12188,N_12183);
nand U12314 (N_12314,N_12171,N_12083);
nand U12315 (N_12315,N_12055,N_12036);
nor U12316 (N_12316,N_12169,N_12021);
and U12317 (N_12317,N_12176,N_12111);
or U12318 (N_12318,N_12202,N_12006);
and U12319 (N_12319,N_12060,N_12144);
or U12320 (N_12320,N_12095,N_12056);
xnor U12321 (N_12321,N_12062,N_12000);
and U12322 (N_12322,N_12085,N_12231);
nand U12323 (N_12323,N_12114,N_12122);
or U12324 (N_12324,N_12117,N_12129);
and U12325 (N_12325,N_12063,N_12033);
or U12326 (N_12326,N_12127,N_12026);
and U12327 (N_12327,N_12185,N_12023);
nor U12328 (N_12328,N_12015,N_12038);
nor U12329 (N_12329,N_12248,N_12241);
nand U12330 (N_12330,N_12091,N_12088);
nand U12331 (N_12331,N_12197,N_12237);
nor U12332 (N_12332,N_12178,N_12064);
nand U12333 (N_12333,N_12115,N_12012);
nand U12334 (N_12334,N_12041,N_12173);
and U12335 (N_12335,N_12128,N_12187);
nor U12336 (N_12336,N_12141,N_12184);
nand U12337 (N_12337,N_12209,N_12002);
and U12338 (N_12338,N_12142,N_12019);
xor U12339 (N_12339,N_12155,N_12226);
nand U12340 (N_12340,N_12163,N_12135);
and U12341 (N_12341,N_12116,N_12072);
xor U12342 (N_12342,N_12246,N_12156);
xnor U12343 (N_12343,N_12228,N_12247);
nor U12344 (N_12344,N_12238,N_12139);
nor U12345 (N_12345,N_12107,N_12075);
nand U12346 (N_12346,N_12208,N_12092);
and U12347 (N_12347,N_12084,N_12024);
xnor U12348 (N_12348,N_12235,N_12118);
nand U12349 (N_12349,N_12087,N_12195);
xnor U12350 (N_12350,N_12175,N_12057);
and U12351 (N_12351,N_12158,N_12152);
or U12352 (N_12352,N_12179,N_12146);
nand U12353 (N_12353,N_12222,N_12157);
xor U12354 (N_12354,N_12096,N_12182);
xor U12355 (N_12355,N_12132,N_12147);
nor U12356 (N_12356,N_12110,N_12205);
nor U12357 (N_12357,N_12093,N_12170);
and U12358 (N_12358,N_12218,N_12124);
nor U12359 (N_12359,N_12243,N_12022);
and U12360 (N_12360,N_12227,N_12225);
nor U12361 (N_12361,N_12004,N_12167);
nor U12362 (N_12362,N_12203,N_12103);
xor U12363 (N_12363,N_12043,N_12008);
xor U12364 (N_12364,N_12076,N_12028);
and U12365 (N_12365,N_12140,N_12223);
xnor U12366 (N_12366,N_12215,N_12230);
xnor U12367 (N_12367,N_12204,N_12174);
xnor U12368 (N_12368,N_12018,N_12034);
xor U12369 (N_12369,N_12193,N_12108);
and U12370 (N_12370,N_12073,N_12123);
xor U12371 (N_12371,N_12217,N_12126);
nor U12372 (N_12372,N_12219,N_12244);
and U12373 (N_12373,N_12098,N_12134);
and U12374 (N_12374,N_12192,N_12214);
xnor U12375 (N_12375,N_12216,N_12185);
nor U12376 (N_12376,N_12107,N_12133);
nor U12377 (N_12377,N_12003,N_12216);
and U12378 (N_12378,N_12213,N_12098);
nand U12379 (N_12379,N_12059,N_12057);
and U12380 (N_12380,N_12148,N_12140);
nand U12381 (N_12381,N_12035,N_12213);
nor U12382 (N_12382,N_12246,N_12222);
or U12383 (N_12383,N_12165,N_12133);
or U12384 (N_12384,N_12046,N_12065);
nand U12385 (N_12385,N_12073,N_12234);
or U12386 (N_12386,N_12047,N_12185);
xor U12387 (N_12387,N_12218,N_12117);
xor U12388 (N_12388,N_12151,N_12145);
xor U12389 (N_12389,N_12194,N_12214);
nor U12390 (N_12390,N_12166,N_12009);
or U12391 (N_12391,N_12163,N_12238);
nand U12392 (N_12392,N_12057,N_12050);
xor U12393 (N_12393,N_12105,N_12008);
or U12394 (N_12394,N_12243,N_12188);
nor U12395 (N_12395,N_12095,N_12029);
xnor U12396 (N_12396,N_12061,N_12086);
nor U12397 (N_12397,N_12200,N_12217);
nor U12398 (N_12398,N_12138,N_12083);
nand U12399 (N_12399,N_12218,N_12018);
nand U12400 (N_12400,N_12173,N_12080);
nor U12401 (N_12401,N_12064,N_12226);
nor U12402 (N_12402,N_12109,N_12238);
nand U12403 (N_12403,N_12032,N_12211);
and U12404 (N_12404,N_12119,N_12039);
or U12405 (N_12405,N_12058,N_12120);
and U12406 (N_12406,N_12070,N_12169);
xor U12407 (N_12407,N_12112,N_12084);
xnor U12408 (N_12408,N_12051,N_12176);
xnor U12409 (N_12409,N_12153,N_12029);
nor U12410 (N_12410,N_12079,N_12159);
and U12411 (N_12411,N_12184,N_12134);
and U12412 (N_12412,N_12188,N_12236);
or U12413 (N_12413,N_12087,N_12109);
xor U12414 (N_12414,N_12183,N_12046);
nand U12415 (N_12415,N_12179,N_12175);
or U12416 (N_12416,N_12184,N_12132);
xnor U12417 (N_12417,N_12153,N_12243);
nand U12418 (N_12418,N_12216,N_12231);
or U12419 (N_12419,N_12207,N_12223);
xnor U12420 (N_12420,N_12009,N_12097);
nand U12421 (N_12421,N_12138,N_12203);
nand U12422 (N_12422,N_12236,N_12167);
nor U12423 (N_12423,N_12140,N_12050);
nor U12424 (N_12424,N_12034,N_12212);
nand U12425 (N_12425,N_12204,N_12167);
xnor U12426 (N_12426,N_12199,N_12067);
or U12427 (N_12427,N_12014,N_12005);
nand U12428 (N_12428,N_12010,N_12098);
nor U12429 (N_12429,N_12215,N_12127);
xnor U12430 (N_12430,N_12115,N_12060);
nor U12431 (N_12431,N_12051,N_12207);
and U12432 (N_12432,N_12192,N_12143);
nor U12433 (N_12433,N_12023,N_12132);
or U12434 (N_12434,N_12030,N_12231);
and U12435 (N_12435,N_12239,N_12145);
nand U12436 (N_12436,N_12151,N_12034);
xor U12437 (N_12437,N_12215,N_12070);
and U12438 (N_12438,N_12187,N_12081);
or U12439 (N_12439,N_12212,N_12225);
nand U12440 (N_12440,N_12249,N_12232);
and U12441 (N_12441,N_12098,N_12231);
xnor U12442 (N_12442,N_12168,N_12083);
nor U12443 (N_12443,N_12212,N_12075);
or U12444 (N_12444,N_12013,N_12194);
nor U12445 (N_12445,N_12174,N_12111);
nand U12446 (N_12446,N_12106,N_12103);
and U12447 (N_12447,N_12103,N_12102);
and U12448 (N_12448,N_12121,N_12068);
and U12449 (N_12449,N_12228,N_12083);
and U12450 (N_12450,N_12220,N_12224);
or U12451 (N_12451,N_12093,N_12001);
nor U12452 (N_12452,N_12140,N_12110);
and U12453 (N_12453,N_12179,N_12211);
nor U12454 (N_12454,N_12214,N_12096);
and U12455 (N_12455,N_12109,N_12128);
nor U12456 (N_12456,N_12012,N_12184);
and U12457 (N_12457,N_12165,N_12122);
nor U12458 (N_12458,N_12006,N_12112);
or U12459 (N_12459,N_12050,N_12083);
or U12460 (N_12460,N_12063,N_12062);
nor U12461 (N_12461,N_12012,N_12238);
xnor U12462 (N_12462,N_12053,N_12069);
and U12463 (N_12463,N_12239,N_12079);
xor U12464 (N_12464,N_12108,N_12103);
or U12465 (N_12465,N_12157,N_12176);
nor U12466 (N_12466,N_12131,N_12225);
nor U12467 (N_12467,N_12010,N_12153);
xor U12468 (N_12468,N_12107,N_12228);
and U12469 (N_12469,N_12001,N_12149);
and U12470 (N_12470,N_12056,N_12032);
xor U12471 (N_12471,N_12131,N_12185);
and U12472 (N_12472,N_12128,N_12003);
nor U12473 (N_12473,N_12225,N_12142);
nor U12474 (N_12474,N_12133,N_12238);
nand U12475 (N_12475,N_12108,N_12225);
and U12476 (N_12476,N_12183,N_12117);
nor U12477 (N_12477,N_12185,N_12056);
nor U12478 (N_12478,N_12015,N_12045);
nor U12479 (N_12479,N_12173,N_12012);
nor U12480 (N_12480,N_12201,N_12220);
nand U12481 (N_12481,N_12095,N_12164);
and U12482 (N_12482,N_12181,N_12174);
nand U12483 (N_12483,N_12014,N_12122);
and U12484 (N_12484,N_12068,N_12160);
or U12485 (N_12485,N_12231,N_12088);
and U12486 (N_12486,N_12161,N_12087);
and U12487 (N_12487,N_12064,N_12207);
xor U12488 (N_12488,N_12094,N_12215);
or U12489 (N_12489,N_12104,N_12230);
nand U12490 (N_12490,N_12219,N_12186);
and U12491 (N_12491,N_12000,N_12197);
or U12492 (N_12492,N_12229,N_12060);
xor U12493 (N_12493,N_12077,N_12200);
xnor U12494 (N_12494,N_12216,N_12099);
and U12495 (N_12495,N_12006,N_12111);
and U12496 (N_12496,N_12078,N_12142);
or U12497 (N_12497,N_12170,N_12033);
nand U12498 (N_12498,N_12010,N_12029);
xor U12499 (N_12499,N_12101,N_12113);
xnor U12500 (N_12500,N_12406,N_12404);
and U12501 (N_12501,N_12457,N_12364);
and U12502 (N_12502,N_12488,N_12382);
nand U12503 (N_12503,N_12346,N_12367);
and U12504 (N_12504,N_12428,N_12442);
nand U12505 (N_12505,N_12268,N_12374);
and U12506 (N_12506,N_12474,N_12286);
and U12507 (N_12507,N_12468,N_12267);
xnor U12508 (N_12508,N_12424,N_12335);
xnor U12509 (N_12509,N_12459,N_12252);
xor U12510 (N_12510,N_12461,N_12472);
and U12511 (N_12511,N_12271,N_12299);
nor U12512 (N_12512,N_12295,N_12453);
or U12513 (N_12513,N_12279,N_12395);
or U12514 (N_12514,N_12273,N_12314);
xnor U12515 (N_12515,N_12381,N_12417);
xnor U12516 (N_12516,N_12334,N_12376);
nand U12517 (N_12517,N_12465,N_12401);
nor U12518 (N_12518,N_12470,N_12433);
xnor U12519 (N_12519,N_12276,N_12300);
and U12520 (N_12520,N_12455,N_12384);
and U12521 (N_12521,N_12407,N_12400);
nand U12522 (N_12522,N_12307,N_12264);
nand U12523 (N_12523,N_12362,N_12421);
xor U12524 (N_12524,N_12265,N_12415);
xnor U12525 (N_12525,N_12414,N_12298);
nand U12526 (N_12526,N_12356,N_12423);
xnor U12527 (N_12527,N_12481,N_12399);
nor U12528 (N_12528,N_12388,N_12447);
nor U12529 (N_12529,N_12479,N_12283);
or U12530 (N_12530,N_12427,N_12498);
or U12531 (N_12531,N_12332,N_12445);
xor U12532 (N_12532,N_12471,N_12326);
and U12533 (N_12533,N_12359,N_12483);
xnor U12534 (N_12534,N_12458,N_12385);
or U12535 (N_12535,N_12444,N_12360);
and U12536 (N_12536,N_12262,N_12439);
xor U12537 (N_12537,N_12310,N_12338);
xnor U12538 (N_12538,N_12348,N_12491);
or U12539 (N_12539,N_12318,N_12402);
and U12540 (N_12540,N_12292,N_12410);
and U12541 (N_12541,N_12323,N_12416);
and U12542 (N_12542,N_12301,N_12496);
and U12543 (N_12543,N_12393,N_12293);
and U12544 (N_12544,N_12419,N_12475);
nor U12545 (N_12545,N_12351,N_12324);
or U12546 (N_12546,N_12313,N_12492);
xnor U12547 (N_12547,N_12303,N_12386);
and U12548 (N_12548,N_12391,N_12254);
nor U12549 (N_12549,N_12263,N_12463);
xor U12550 (N_12550,N_12389,N_12284);
and U12551 (N_12551,N_12256,N_12305);
or U12552 (N_12552,N_12336,N_12451);
and U12553 (N_12553,N_12450,N_12343);
xnor U12554 (N_12554,N_12409,N_12490);
nand U12555 (N_12555,N_12390,N_12280);
and U12556 (N_12556,N_12432,N_12473);
and U12557 (N_12557,N_12350,N_12380);
xor U12558 (N_12558,N_12339,N_12426);
nor U12559 (N_12559,N_12365,N_12394);
nand U12560 (N_12560,N_12377,N_12287);
nand U12561 (N_12561,N_12486,N_12291);
and U12562 (N_12562,N_12311,N_12438);
nor U12563 (N_12563,N_12282,N_12422);
nor U12564 (N_12564,N_12317,N_12255);
or U12565 (N_12565,N_12330,N_12460);
nor U12566 (N_12566,N_12328,N_12289);
nor U12567 (N_12567,N_12495,N_12297);
xor U12568 (N_12568,N_12315,N_12448);
and U12569 (N_12569,N_12352,N_12322);
nand U12570 (N_12570,N_12369,N_12354);
xnor U12571 (N_12571,N_12397,N_12331);
xnor U12572 (N_12572,N_12452,N_12420);
xnor U12573 (N_12573,N_12251,N_12418);
or U12574 (N_12574,N_12342,N_12278);
or U12575 (N_12575,N_12411,N_12368);
or U12576 (N_12576,N_12319,N_12366);
or U12577 (N_12577,N_12304,N_12499);
xnor U12578 (N_12578,N_12329,N_12456);
and U12579 (N_12579,N_12378,N_12436);
nand U12580 (N_12580,N_12259,N_12408);
nor U12581 (N_12581,N_12261,N_12434);
or U12582 (N_12582,N_12478,N_12269);
xor U12583 (N_12583,N_12341,N_12435);
or U12584 (N_12584,N_12405,N_12253);
xor U12585 (N_12585,N_12441,N_12464);
nand U12586 (N_12586,N_12285,N_12327);
nor U12587 (N_12587,N_12355,N_12412);
nand U12588 (N_12588,N_12489,N_12446);
and U12589 (N_12589,N_12379,N_12403);
xnor U12590 (N_12590,N_12466,N_12443);
xnor U12591 (N_12591,N_12270,N_12302);
xnor U12592 (N_12592,N_12308,N_12467);
nor U12593 (N_12593,N_12437,N_12425);
xor U12594 (N_12594,N_12361,N_12371);
and U12595 (N_12595,N_12449,N_12396);
xor U12596 (N_12596,N_12387,N_12347);
nor U12597 (N_12597,N_12373,N_12430);
nand U12598 (N_12598,N_12375,N_12275);
and U12599 (N_12599,N_12257,N_12272);
nand U12600 (N_12600,N_12358,N_12316);
xnor U12601 (N_12601,N_12333,N_12266);
nor U12602 (N_12602,N_12260,N_12487);
nand U12603 (N_12603,N_12494,N_12288);
nor U12604 (N_12604,N_12296,N_12349);
and U12605 (N_12605,N_12462,N_12370);
and U12606 (N_12606,N_12306,N_12482);
nor U12607 (N_12607,N_12383,N_12476);
nor U12608 (N_12608,N_12290,N_12312);
nand U12609 (N_12609,N_12294,N_12363);
nand U12610 (N_12610,N_12320,N_12440);
or U12611 (N_12611,N_12484,N_12258);
nand U12612 (N_12612,N_12493,N_12485);
nor U12613 (N_12613,N_12372,N_12454);
nor U12614 (N_12614,N_12480,N_12274);
xnor U12615 (N_12615,N_12309,N_12277);
nand U12616 (N_12616,N_12321,N_12497);
nor U12617 (N_12617,N_12477,N_12357);
nor U12618 (N_12618,N_12281,N_12325);
or U12619 (N_12619,N_12344,N_12398);
xnor U12620 (N_12620,N_12413,N_12340);
nand U12621 (N_12621,N_12392,N_12250);
xnor U12622 (N_12622,N_12337,N_12469);
xnor U12623 (N_12623,N_12353,N_12431);
nand U12624 (N_12624,N_12429,N_12345);
nor U12625 (N_12625,N_12458,N_12419);
nand U12626 (N_12626,N_12443,N_12379);
xor U12627 (N_12627,N_12375,N_12268);
nor U12628 (N_12628,N_12250,N_12316);
nand U12629 (N_12629,N_12489,N_12420);
nor U12630 (N_12630,N_12446,N_12326);
and U12631 (N_12631,N_12469,N_12298);
nor U12632 (N_12632,N_12451,N_12397);
nand U12633 (N_12633,N_12345,N_12417);
nand U12634 (N_12634,N_12413,N_12380);
nand U12635 (N_12635,N_12458,N_12360);
xor U12636 (N_12636,N_12327,N_12404);
xnor U12637 (N_12637,N_12272,N_12462);
nand U12638 (N_12638,N_12276,N_12497);
xor U12639 (N_12639,N_12491,N_12276);
nor U12640 (N_12640,N_12319,N_12387);
or U12641 (N_12641,N_12267,N_12470);
xor U12642 (N_12642,N_12276,N_12412);
nor U12643 (N_12643,N_12369,N_12294);
xnor U12644 (N_12644,N_12479,N_12439);
nand U12645 (N_12645,N_12312,N_12491);
nor U12646 (N_12646,N_12277,N_12254);
nor U12647 (N_12647,N_12261,N_12353);
xor U12648 (N_12648,N_12360,N_12374);
xor U12649 (N_12649,N_12420,N_12377);
nand U12650 (N_12650,N_12257,N_12268);
or U12651 (N_12651,N_12304,N_12496);
nand U12652 (N_12652,N_12341,N_12466);
nand U12653 (N_12653,N_12404,N_12347);
nor U12654 (N_12654,N_12338,N_12407);
nor U12655 (N_12655,N_12414,N_12293);
nand U12656 (N_12656,N_12478,N_12459);
nand U12657 (N_12657,N_12337,N_12400);
or U12658 (N_12658,N_12323,N_12316);
nand U12659 (N_12659,N_12399,N_12498);
nand U12660 (N_12660,N_12384,N_12318);
xnor U12661 (N_12661,N_12367,N_12305);
and U12662 (N_12662,N_12251,N_12391);
nand U12663 (N_12663,N_12428,N_12302);
xor U12664 (N_12664,N_12423,N_12257);
or U12665 (N_12665,N_12260,N_12297);
nand U12666 (N_12666,N_12419,N_12345);
xor U12667 (N_12667,N_12365,N_12264);
nor U12668 (N_12668,N_12418,N_12444);
nand U12669 (N_12669,N_12355,N_12312);
or U12670 (N_12670,N_12376,N_12439);
or U12671 (N_12671,N_12319,N_12285);
nor U12672 (N_12672,N_12495,N_12467);
and U12673 (N_12673,N_12251,N_12348);
nor U12674 (N_12674,N_12396,N_12402);
nor U12675 (N_12675,N_12332,N_12454);
xor U12676 (N_12676,N_12339,N_12286);
nor U12677 (N_12677,N_12252,N_12287);
and U12678 (N_12678,N_12380,N_12491);
nor U12679 (N_12679,N_12417,N_12360);
nor U12680 (N_12680,N_12480,N_12315);
nor U12681 (N_12681,N_12320,N_12497);
xnor U12682 (N_12682,N_12333,N_12454);
nand U12683 (N_12683,N_12493,N_12328);
nor U12684 (N_12684,N_12484,N_12492);
nor U12685 (N_12685,N_12353,N_12256);
xnor U12686 (N_12686,N_12370,N_12363);
nor U12687 (N_12687,N_12462,N_12383);
and U12688 (N_12688,N_12463,N_12474);
nor U12689 (N_12689,N_12443,N_12339);
or U12690 (N_12690,N_12382,N_12296);
nand U12691 (N_12691,N_12470,N_12421);
or U12692 (N_12692,N_12483,N_12468);
xnor U12693 (N_12693,N_12455,N_12411);
nor U12694 (N_12694,N_12333,N_12282);
or U12695 (N_12695,N_12343,N_12477);
nand U12696 (N_12696,N_12321,N_12335);
nand U12697 (N_12697,N_12427,N_12475);
nor U12698 (N_12698,N_12376,N_12436);
or U12699 (N_12699,N_12462,N_12420);
nor U12700 (N_12700,N_12309,N_12356);
or U12701 (N_12701,N_12453,N_12325);
nand U12702 (N_12702,N_12477,N_12472);
and U12703 (N_12703,N_12381,N_12465);
or U12704 (N_12704,N_12353,N_12373);
xnor U12705 (N_12705,N_12300,N_12360);
xor U12706 (N_12706,N_12252,N_12469);
nor U12707 (N_12707,N_12495,N_12300);
nor U12708 (N_12708,N_12282,N_12370);
nand U12709 (N_12709,N_12372,N_12358);
nor U12710 (N_12710,N_12395,N_12439);
nor U12711 (N_12711,N_12315,N_12357);
or U12712 (N_12712,N_12255,N_12379);
nor U12713 (N_12713,N_12498,N_12266);
xnor U12714 (N_12714,N_12269,N_12340);
and U12715 (N_12715,N_12363,N_12499);
nand U12716 (N_12716,N_12285,N_12377);
nor U12717 (N_12717,N_12394,N_12488);
nor U12718 (N_12718,N_12256,N_12395);
nor U12719 (N_12719,N_12343,N_12255);
xnor U12720 (N_12720,N_12269,N_12414);
nand U12721 (N_12721,N_12446,N_12385);
and U12722 (N_12722,N_12466,N_12439);
xnor U12723 (N_12723,N_12289,N_12424);
or U12724 (N_12724,N_12410,N_12294);
or U12725 (N_12725,N_12323,N_12427);
or U12726 (N_12726,N_12297,N_12338);
and U12727 (N_12727,N_12251,N_12395);
and U12728 (N_12728,N_12427,N_12259);
nand U12729 (N_12729,N_12455,N_12495);
and U12730 (N_12730,N_12466,N_12477);
nor U12731 (N_12731,N_12342,N_12396);
nor U12732 (N_12732,N_12310,N_12355);
and U12733 (N_12733,N_12343,N_12349);
nor U12734 (N_12734,N_12334,N_12488);
xor U12735 (N_12735,N_12377,N_12307);
or U12736 (N_12736,N_12325,N_12351);
nand U12737 (N_12737,N_12400,N_12284);
nor U12738 (N_12738,N_12332,N_12399);
nor U12739 (N_12739,N_12328,N_12422);
or U12740 (N_12740,N_12479,N_12399);
or U12741 (N_12741,N_12469,N_12428);
or U12742 (N_12742,N_12452,N_12372);
xor U12743 (N_12743,N_12371,N_12457);
nand U12744 (N_12744,N_12396,N_12439);
nand U12745 (N_12745,N_12480,N_12376);
nor U12746 (N_12746,N_12446,N_12269);
nor U12747 (N_12747,N_12455,N_12450);
nand U12748 (N_12748,N_12306,N_12266);
and U12749 (N_12749,N_12266,N_12441);
and U12750 (N_12750,N_12748,N_12720);
nor U12751 (N_12751,N_12522,N_12578);
nor U12752 (N_12752,N_12699,N_12541);
nor U12753 (N_12753,N_12671,N_12561);
and U12754 (N_12754,N_12690,N_12563);
xor U12755 (N_12755,N_12652,N_12695);
nor U12756 (N_12756,N_12548,N_12634);
and U12757 (N_12757,N_12656,N_12509);
nand U12758 (N_12758,N_12620,N_12661);
and U12759 (N_12759,N_12609,N_12705);
nand U12760 (N_12760,N_12507,N_12594);
xnor U12761 (N_12761,N_12738,N_12730);
or U12762 (N_12762,N_12542,N_12693);
or U12763 (N_12763,N_12736,N_12668);
or U12764 (N_12764,N_12623,N_12581);
nand U12765 (N_12765,N_12743,N_12707);
and U12766 (N_12766,N_12729,N_12544);
and U12767 (N_12767,N_12501,N_12567);
nand U12768 (N_12768,N_12659,N_12747);
and U12769 (N_12769,N_12517,N_12545);
nor U12770 (N_12770,N_12641,N_12624);
or U12771 (N_12771,N_12639,N_12665);
nor U12772 (N_12772,N_12513,N_12653);
xnor U12773 (N_12773,N_12512,N_12734);
xnor U12774 (N_12774,N_12583,N_12564);
xor U12775 (N_12775,N_12691,N_12602);
and U12776 (N_12776,N_12536,N_12711);
or U12777 (N_12777,N_12534,N_12685);
nand U12778 (N_12778,N_12560,N_12651);
nor U12779 (N_12779,N_12603,N_12704);
or U12780 (N_12780,N_12526,N_12584);
nand U12781 (N_12781,N_12604,N_12638);
nor U12782 (N_12782,N_12601,N_12592);
nor U12783 (N_12783,N_12682,N_12529);
xnor U12784 (N_12784,N_12537,N_12657);
or U12785 (N_12785,N_12527,N_12577);
or U12786 (N_12786,N_12713,N_12669);
nor U12787 (N_12787,N_12532,N_12687);
nor U12788 (N_12788,N_12709,N_12549);
nand U12789 (N_12789,N_12675,N_12551);
xor U12790 (N_12790,N_12640,N_12539);
and U12791 (N_12791,N_12573,N_12686);
and U12792 (N_12792,N_12703,N_12684);
and U12793 (N_12793,N_12618,N_12519);
nand U12794 (N_12794,N_12621,N_12658);
and U12795 (N_12795,N_12540,N_12698);
and U12796 (N_12796,N_12700,N_12596);
and U12797 (N_12797,N_12617,N_12511);
and U12798 (N_12798,N_12721,N_12586);
nand U12799 (N_12799,N_12673,N_12531);
nor U12800 (N_12800,N_12628,N_12506);
xnor U12801 (N_12801,N_12666,N_12708);
or U12802 (N_12802,N_12735,N_12633);
or U12803 (N_12803,N_12579,N_12515);
nor U12804 (N_12804,N_12535,N_12547);
or U12805 (N_12805,N_12622,N_12590);
nor U12806 (N_12806,N_12554,N_12546);
nand U12807 (N_12807,N_12557,N_12599);
xnor U12808 (N_12808,N_12631,N_12614);
xor U12809 (N_12809,N_12716,N_12740);
and U12810 (N_12810,N_12739,N_12676);
nand U12811 (N_12811,N_12728,N_12732);
nor U12812 (N_12812,N_12642,N_12677);
nand U12813 (N_12813,N_12606,N_12649);
nand U12814 (N_12814,N_12663,N_12683);
or U12815 (N_12815,N_12608,N_12570);
nand U12816 (N_12816,N_12742,N_12524);
nor U12817 (N_12817,N_12615,N_12654);
and U12818 (N_12818,N_12645,N_12520);
nand U12819 (N_12819,N_12710,N_12530);
and U12820 (N_12820,N_12562,N_12627);
and U12821 (N_12821,N_12714,N_12538);
nor U12822 (N_12822,N_12701,N_12533);
and U12823 (N_12823,N_12702,N_12587);
nor U12824 (N_12824,N_12575,N_12625);
nand U12825 (N_12825,N_12613,N_12607);
xnor U12826 (N_12826,N_12737,N_12543);
nand U12827 (N_12827,N_12508,N_12616);
nand U12828 (N_12828,N_12574,N_12523);
and U12829 (N_12829,N_12678,N_12552);
xor U12830 (N_12830,N_12612,N_12745);
and U12831 (N_12831,N_12582,N_12502);
nor U12832 (N_12832,N_12636,N_12670);
nand U12833 (N_12833,N_12718,N_12746);
and U12834 (N_12834,N_12588,N_12528);
or U12835 (N_12835,N_12696,N_12689);
xor U12836 (N_12836,N_12725,N_12568);
nor U12837 (N_12837,N_12741,N_12648);
or U12838 (N_12838,N_12647,N_12637);
nor U12839 (N_12839,N_12723,N_12722);
xnor U12840 (N_12840,N_12632,N_12580);
nand U12841 (N_12841,N_12667,N_12510);
xnor U12842 (N_12842,N_12680,N_12674);
nand U12843 (N_12843,N_12679,N_12555);
nor U12844 (N_12844,N_12559,N_12697);
nand U12845 (N_12845,N_12727,N_12731);
and U12846 (N_12846,N_12565,N_12712);
nand U12847 (N_12847,N_12514,N_12719);
and U12848 (N_12848,N_12672,N_12593);
nor U12849 (N_12849,N_12503,N_12566);
or U12850 (N_12850,N_12585,N_12646);
xnor U12851 (N_12851,N_12619,N_12629);
or U12852 (N_12852,N_12611,N_12600);
or U12853 (N_12853,N_12610,N_12595);
and U12854 (N_12854,N_12605,N_12525);
and U12855 (N_12855,N_12589,N_12558);
or U12856 (N_12856,N_12597,N_12505);
or U12857 (N_12857,N_12744,N_12660);
and U12858 (N_12858,N_12717,N_12626);
nand U12859 (N_12859,N_12644,N_12733);
nor U12860 (N_12860,N_12504,N_12521);
and U12861 (N_12861,N_12692,N_12664);
xnor U12862 (N_12862,N_12518,N_12681);
or U12863 (N_12863,N_12694,N_12500);
xor U12864 (N_12864,N_12550,N_12715);
or U12865 (N_12865,N_12630,N_12662);
and U12866 (N_12866,N_12572,N_12598);
nand U12867 (N_12867,N_12724,N_12553);
xnor U12868 (N_12868,N_12516,N_12556);
nor U12869 (N_12869,N_12749,N_12655);
and U12870 (N_12870,N_12706,N_12591);
nor U12871 (N_12871,N_12635,N_12569);
nor U12872 (N_12872,N_12576,N_12643);
and U12873 (N_12873,N_12726,N_12650);
or U12874 (N_12874,N_12571,N_12688);
and U12875 (N_12875,N_12646,N_12656);
nor U12876 (N_12876,N_12518,N_12579);
xor U12877 (N_12877,N_12678,N_12740);
xnor U12878 (N_12878,N_12688,N_12586);
nand U12879 (N_12879,N_12544,N_12548);
nor U12880 (N_12880,N_12654,N_12527);
xnor U12881 (N_12881,N_12671,N_12690);
nor U12882 (N_12882,N_12513,N_12657);
or U12883 (N_12883,N_12733,N_12666);
nand U12884 (N_12884,N_12662,N_12599);
or U12885 (N_12885,N_12594,N_12606);
nand U12886 (N_12886,N_12710,N_12641);
xnor U12887 (N_12887,N_12664,N_12535);
nand U12888 (N_12888,N_12599,N_12742);
and U12889 (N_12889,N_12583,N_12688);
or U12890 (N_12890,N_12564,N_12577);
or U12891 (N_12891,N_12519,N_12737);
or U12892 (N_12892,N_12730,N_12533);
nand U12893 (N_12893,N_12645,N_12669);
xor U12894 (N_12894,N_12518,N_12712);
nand U12895 (N_12895,N_12714,N_12707);
or U12896 (N_12896,N_12732,N_12623);
and U12897 (N_12897,N_12586,N_12653);
or U12898 (N_12898,N_12708,N_12716);
nor U12899 (N_12899,N_12728,N_12646);
nand U12900 (N_12900,N_12516,N_12737);
nand U12901 (N_12901,N_12731,N_12625);
xor U12902 (N_12902,N_12720,N_12735);
or U12903 (N_12903,N_12722,N_12670);
or U12904 (N_12904,N_12593,N_12513);
nor U12905 (N_12905,N_12677,N_12735);
or U12906 (N_12906,N_12624,N_12570);
or U12907 (N_12907,N_12650,N_12701);
or U12908 (N_12908,N_12667,N_12737);
and U12909 (N_12909,N_12527,N_12737);
or U12910 (N_12910,N_12744,N_12560);
nor U12911 (N_12911,N_12559,N_12714);
or U12912 (N_12912,N_12619,N_12652);
or U12913 (N_12913,N_12646,N_12558);
nand U12914 (N_12914,N_12663,N_12643);
nand U12915 (N_12915,N_12507,N_12634);
xor U12916 (N_12916,N_12502,N_12720);
and U12917 (N_12917,N_12722,N_12622);
nor U12918 (N_12918,N_12549,N_12531);
nand U12919 (N_12919,N_12643,N_12599);
or U12920 (N_12920,N_12737,N_12701);
and U12921 (N_12921,N_12732,N_12562);
xor U12922 (N_12922,N_12571,N_12552);
xnor U12923 (N_12923,N_12727,N_12682);
nor U12924 (N_12924,N_12587,N_12514);
xor U12925 (N_12925,N_12646,N_12575);
and U12926 (N_12926,N_12561,N_12727);
and U12927 (N_12927,N_12559,N_12700);
nand U12928 (N_12928,N_12667,N_12517);
nor U12929 (N_12929,N_12547,N_12603);
nand U12930 (N_12930,N_12687,N_12615);
or U12931 (N_12931,N_12531,N_12715);
nand U12932 (N_12932,N_12721,N_12747);
nand U12933 (N_12933,N_12656,N_12745);
nand U12934 (N_12934,N_12715,N_12615);
nand U12935 (N_12935,N_12563,N_12632);
nand U12936 (N_12936,N_12586,N_12659);
xnor U12937 (N_12937,N_12688,N_12600);
nand U12938 (N_12938,N_12730,N_12607);
or U12939 (N_12939,N_12638,N_12675);
nand U12940 (N_12940,N_12584,N_12626);
and U12941 (N_12941,N_12721,N_12546);
nor U12942 (N_12942,N_12572,N_12530);
or U12943 (N_12943,N_12541,N_12674);
nor U12944 (N_12944,N_12503,N_12658);
or U12945 (N_12945,N_12603,N_12513);
and U12946 (N_12946,N_12689,N_12579);
nand U12947 (N_12947,N_12558,N_12665);
or U12948 (N_12948,N_12647,N_12661);
and U12949 (N_12949,N_12587,N_12730);
or U12950 (N_12950,N_12689,N_12576);
nand U12951 (N_12951,N_12706,N_12589);
nor U12952 (N_12952,N_12747,N_12574);
and U12953 (N_12953,N_12557,N_12692);
nor U12954 (N_12954,N_12605,N_12746);
and U12955 (N_12955,N_12527,N_12530);
nand U12956 (N_12956,N_12616,N_12658);
xnor U12957 (N_12957,N_12641,N_12608);
nor U12958 (N_12958,N_12535,N_12744);
nand U12959 (N_12959,N_12531,N_12650);
nor U12960 (N_12960,N_12670,N_12669);
and U12961 (N_12961,N_12713,N_12715);
or U12962 (N_12962,N_12533,N_12700);
nand U12963 (N_12963,N_12535,N_12584);
nor U12964 (N_12964,N_12712,N_12592);
and U12965 (N_12965,N_12688,N_12741);
xnor U12966 (N_12966,N_12637,N_12620);
nor U12967 (N_12967,N_12741,N_12595);
xnor U12968 (N_12968,N_12748,N_12533);
nor U12969 (N_12969,N_12616,N_12653);
nand U12970 (N_12970,N_12649,N_12693);
nand U12971 (N_12971,N_12606,N_12602);
nand U12972 (N_12972,N_12641,N_12698);
and U12973 (N_12973,N_12522,N_12567);
nand U12974 (N_12974,N_12518,N_12697);
or U12975 (N_12975,N_12561,N_12591);
xnor U12976 (N_12976,N_12558,N_12563);
nand U12977 (N_12977,N_12590,N_12585);
or U12978 (N_12978,N_12526,N_12540);
or U12979 (N_12979,N_12582,N_12642);
or U12980 (N_12980,N_12650,N_12674);
nor U12981 (N_12981,N_12744,N_12649);
and U12982 (N_12982,N_12578,N_12707);
nor U12983 (N_12983,N_12590,N_12704);
nor U12984 (N_12984,N_12512,N_12622);
and U12985 (N_12985,N_12543,N_12562);
nor U12986 (N_12986,N_12580,N_12719);
nor U12987 (N_12987,N_12611,N_12715);
and U12988 (N_12988,N_12622,N_12665);
nand U12989 (N_12989,N_12638,N_12506);
nand U12990 (N_12990,N_12636,N_12639);
xnor U12991 (N_12991,N_12535,N_12688);
nor U12992 (N_12992,N_12660,N_12618);
nand U12993 (N_12993,N_12705,N_12531);
xor U12994 (N_12994,N_12729,N_12501);
and U12995 (N_12995,N_12531,N_12618);
nor U12996 (N_12996,N_12638,N_12627);
and U12997 (N_12997,N_12641,N_12509);
nand U12998 (N_12998,N_12526,N_12664);
xor U12999 (N_12999,N_12544,N_12705);
nor U13000 (N_13000,N_12962,N_12757);
or U13001 (N_13001,N_12980,N_12914);
and U13002 (N_13002,N_12779,N_12798);
or U13003 (N_13003,N_12760,N_12926);
xnor U13004 (N_13004,N_12984,N_12953);
nand U13005 (N_13005,N_12911,N_12781);
and U13006 (N_13006,N_12761,N_12865);
xor U13007 (N_13007,N_12884,N_12994);
or U13008 (N_13008,N_12968,N_12908);
nor U13009 (N_13009,N_12906,N_12848);
and U13010 (N_13010,N_12912,N_12769);
nand U13011 (N_13011,N_12810,N_12859);
nand U13012 (N_13012,N_12857,N_12837);
or U13013 (N_13013,N_12896,N_12839);
xnor U13014 (N_13014,N_12782,N_12990);
nand U13015 (N_13015,N_12972,N_12802);
nand U13016 (N_13016,N_12875,N_12961);
nand U13017 (N_13017,N_12868,N_12890);
nand U13018 (N_13018,N_12936,N_12835);
nand U13019 (N_13019,N_12882,N_12995);
or U13020 (N_13020,N_12907,N_12955);
and U13021 (N_13021,N_12895,N_12966);
xor U13022 (N_13022,N_12776,N_12864);
xnor U13023 (N_13023,N_12822,N_12755);
nor U13024 (N_13024,N_12963,N_12965);
xnor U13025 (N_13025,N_12910,N_12897);
nor U13026 (N_13026,N_12973,N_12762);
or U13027 (N_13027,N_12836,N_12945);
nand U13028 (N_13028,N_12949,N_12944);
or U13029 (N_13029,N_12916,N_12795);
or U13030 (N_13030,N_12918,N_12983);
or U13031 (N_13031,N_12797,N_12816);
or U13032 (N_13032,N_12904,N_12826);
and U13033 (N_13033,N_12866,N_12964);
nand U13034 (N_13034,N_12909,N_12880);
and U13035 (N_13035,N_12778,N_12811);
nor U13036 (N_13036,N_12869,N_12981);
xor U13037 (N_13037,N_12969,N_12812);
and U13038 (N_13038,N_12931,N_12929);
xor U13039 (N_13039,N_12758,N_12878);
nand U13040 (N_13040,N_12818,N_12899);
and U13041 (N_13041,N_12967,N_12947);
xnor U13042 (N_13042,N_12893,N_12825);
or U13043 (N_13043,N_12791,N_12856);
nand U13044 (N_13044,N_12838,N_12996);
or U13045 (N_13045,N_12752,N_12765);
nor U13046 (N_13046,N_12861,N_12808);
xnor U13047 (N_13047,N_12974,N_12928);
xnor U13048 (N_13048,N_12937,N_12844);
nand U13049 (N_13049,N_12793,N_12922);
nand U13050 (N_13050,N_12913,N_12886);
or U13051 (N_13051,N_12954,N_12794);
or U13052 (N_13052,N_12942,N_12842);
xnor U13053 (N_13053,N_12847,N_12923);
xnor U13054 (N_13054,N_12946,N_12823);
nand U13055 (N_13055,N_12924,N_12959);
or U13056 (N_13056,N_12932,N_12796);
xnor U13057 (N_13057,N_12786,N_12809);
and U13058 (N_13058,N_12903,N_12885);
xor U13059 (N_13059,N_12766,N_12831);
nor U13060 (N_13060,N_12921,N_12957);
or U13061 (N_13061,N_12971,N_12871);
and U13062 (N_13062,N_12833,N_12905);
or U13063 (N_13063,N_12827,N_12925);
and U13064 (N_13064,N_12817,N_12845);
xnor U13065 (N_13065,N_12862,N_12813);
or U13066 (N_13066,N_12768,N_12783);
nor U13067 (N_13067,N_12920,N_12876);
xor U13068 (N_13068,N_12854,N_12881);
nor U13069 (N_13069,N_12997,N_12832);
nor U13070 (N_13070,N_12933,N_12767);
or U13071 (N_13071,N_12902,N_12787);
and U13072 (N_13072,N_12982,N_12850);
and U13073 (N_13073,N_12919,N_12999);
nor U13074 (N_13074,N_12840,N_12800);
nand U13075 (N_13075,N_12804,N_12849);
nand U13076 (N_13076,N_12846,N_12777);
and U13077 (N_13077,N_12891,N_12759);
and U13078 (N_13078,N_12887,N_12750);
and U13079 (N_13079,N_12770,N_12774);
or U13080 (N_13080,N_12943,N_12824);
nand U13081 (N_13081,N_12977,N_12883);
xnor U13082 (N_13082,N_12851,N_12948);
xnor U13083 (N_13083,N_12940,N_12958);
and U13084 (N_13084,N_12879,N_12898);
xor U13085 (N_13085,N_12775,N_12976);
or U13086 (N_13086,N_12772,N_12780);
and U13087 (N_13087,N_12989,N_12935);
nor U13088 (N_13088,N_12754,N_12892);
and U13089 (N_13089,N_12763,N_12987);
xnor U13090 (N_13090,N_12820,N_12814);
or U13091 (N_13091,N_12877,N_12756);
and U13092 (N_13092,N_12792,N_12801);
or U13093 (N_13093,N_12979,N_12998);
nand U13094 (N_13094,N_12789,N_12852);
xor U13095 (N_13095,N_12753,N_12830);
and U13096 (N_13096,N_12855,N_12901);
nor U13097 (N_13097,N_12819,N_12889);
nand U13098 (N_13098,N_12764,N_12874);
nand U13099 (N_13099,N_12785,N_12970);
xor U13100 (N_13100,N_12915,N_12828);
nor U13101 (N_13101,N_12960,N_12951);
xnor U13102 (N_13102,N_12985,N_12934);
or U13103 (N_13103,N_12978,N_12784);
xor U13104 (N_13104,N_12805,N_12806);
and U13105 (N_13105,N_12788,N_12941);
nor U13106 (N_13106,N_12803,N_12930);
nor U13107 (N_13107,N_12860,N_12843);
and U13108 (N_13108,N_12867,N_12900);
nor U13109 (N_13109,N_12986,N_12975);
xor U13110 (N_13110,N_12821,N_12815);
xor U13111 (N_13111,N_12956,N_12888);
and U13112 (N_13112,N_12952,N_12988);
or U13113 (N_13113,N_12992,N_12858);
and U13114 (N_13114,N_12939,N_12917);
xnor U13115 (N_13115,N_12773,N_12894);
or U13116 (N_13116,N_12771,N_12807);
nand U13117 (N_13117,N_12938,N_12790);
nand U13118 (N_13118,N_12950,N_12834);
nand U13119 (N_13119,N_12870,N_12829);
nor U13120 (N_13120,N_12991,N_12751);
and U13121 (N_13121,N_12863,N_12873);
and U13122 (N_13122,N_12872,N_12799);
nor U13123 (N_13123,N_12841,N_12853);
and U13124 (N_13124,N_12993,N_12927);
xnor U13125 (N_13125,N_12753,N_12943);
and U13126 (N_13126,N_12782,N_12796);
and U13127 (N_13127,N_12804,N_12879);
nand U13128 (N_13128,N_12855,N_12768);
and U13129 (N_13129,N_12797,N_12999);
and U13130 (N_13130,N_12815,N_12840);
nand U13131 (N_13131,N_12982,N_12974);
and U13132 (N_13132,N_12778,N_12909);
and U13133 (N_13133,N_12816,N_12971);
or U13134 (N_13134,N_12905,N_12901);
or U13135 (N_13135,N_12822,N_12799);
or U13136 (N_13136,N_12840,N_12863);
and U13137 (N_13137,N_12931,N_12758);
xor U13138 (N_13138,N_12841,N_12918);
nand U13139 (N_13139,N_12895,N_12879);
xnor U13140 (N_13140,N_12929,N_12855);
and U13141 (N_13141,N_12786,N_12817);
or U13142 (N_13142,N_12916,N_12857);
and U13143 (N_13143,N_12886,N_12752);
nand U13144 (N_13144,N_12875,N_12920);
nor U13145 (N_13145,N_12809,N_12988);
or U13146 (N_13146,N_12972,N_12765);
or U13147 (N_13147,N_12782,N_12907);
nand U13148 (N_13148,N_12871,N_12960);
or U13149 (N_13149,N_12892,N_12987);
nor U13150 (N_13150,N_12822,N_12837);
xnor U13151 (N_13151,N_12779,N_12846);
and U13152 (N_13152,N_12888,N_12893);
nand U13153 (N_13153,N_12860,N_12768);
nor U13154 (N_13154,N_12995,N_12758);
or U13155 (N_13155,N_12835,N_12820);
nor U13156 (N_13156,N_12806,N_12993);
nor U13157 (N_13157,N_12830,N_12984);
nand U13158 (N_13158,N_12869,N_12843);
and U13159 (N_13159,N_12853,N_12983);
nor U13160 (N_13160,N_12916,N_12975);
and U13161 (N_13161,N_12930,N_12937);
and U13162 (N_13162,N_12886,N_12986);
xnor U13163 (N_13163,N_12971,N_12968);
or U13164 (N_13164,N_12775,N_12834);
or U13165 (N_13165,N_12821,N_12870);
or U13166 (N_13166,N_12845,N_12782);
and U13167 (N_13167,N_12928,N_12962);
and U13168 (N_13168,N_12848,N_12841);
nor U13169 (N_13169,N_12965,N_12806);
xnor U13170 (N_13170,N_12872,N_12999);
xor U13171 (N_13171,N_12877,N_12908);
or U13172 (N_13172,N_12767,N_12856);
nor U13173 (N_13173,N_12864,N_12943);
and U13174 (N_13174,N_12931,N_12971);
or U13175 (N_13175,N_12861,N_12788);
or U13176 (N_13176,N_12960,N_12879);
and U13177 (N_13177,N_12979,N_12792);
nand U13178 (N_13178,N_12904,N_12759);
nor U13179 (N_13179,N_12996,N_12914);
or U13180 (N_13180,N_12938,N_12912);
nand U13181 (N_13181,N_12989,N_12992);
nor U13182 (N_13182,N_12884,N_12873);
or U13183 (N_13183,N_12804,N_12963);
nand U13184 (N_13184,N_12829,N_12978);
or U13185 (N_13185,N_12972,N_12868);
xor U13186 (N_13186,N_12982,N_12951);
or U13187 (N_13187,N_12874,N_12780);
or U13188 (N_13188,N_12765,N_12866);
or U13189 (N_13189,N_12992,N_12789);
nor U13190 (N_13190,N_12925,N_12878);
xor U13191 (N_13191,N_12877,N_12917);
nor U13192 (N_13192,N_12765,N_12863);
and U13193 (N_13193,N_12868,N_12816);
nor U13194 (N_13194,N_12992,N_12980);
or U13195 (N_13195,N_12894,N_12919);
xnor U13196 (N_13196,N_12775,N_12996);
and U13197 (N_13197,N_12913,N_12762);
xor U13198 (N_13198,N_12832,N_12961);
xnor U13199 (N_13199,N_12957,N_12906);
or U13200 (N_13200,N_12838,N_12995);
and U13201 (N_13201,N_12840,N_12771);
nand U13202 (N_13202,N_12768,N_12927);
and U13203 (N_13203,N_12757,N_12822);
nor U13204 (N_13204,N_12812,N_12890);
xnor U13205 (N_13205,N_12907,N_12821);
nand U13206 (N_13206,N_12993,N_12981);
nor U13207 (N_13207,N_12882,N_12999);
and U13208 (N_13208,N_12826,N_12997);
nand U13209 (N_13209,N_12985,N_12881);
nor U13210 (N_13210,N_12911,N_12750);
and U13211 (N_13211,N_12772,N_12900);
nand U13212 (N_13212,N_12963,N_12932);
xor U13213 (N_13213,N_12829,N_12876);
xor U13214 (N_13214,N_12766,N_12911);
or U13215 (N_13215,N_12782,N_12944);
nand U13216 (N_13216,N_12808,N_12882);
xnor U13217 (N_13217,N_12775,N_12935);
nor U13218 (N_13218,N_12790,N_12948);
xnor U13219 (N_13219,N_12800,N_12775);
nand U13220 (N_13220,N_12987,N_12907);
xnor U13221 (N_13221,N_12994,N_12868);
nor U13222 (N_13222,N_12792,N_12762);
and U13223 (N_13223,N_12842,N_12928);
xnor U13224 (N_13224,N_12947,N_12797);
and U13225 (N_13225,N_12819,N_12916);
nor U13226 (N_13226,N_12858,N_12929);
nand U13227 (N_13227,N_12985,N_12789);
or U13228 (N_13228,N_12800,N_12998);
and U13229 (N_13229,N_12927,N_12819);
nor U13230 (N_13230,N_12815,N_12826);
nor U13231 (N_13231,N_12959,N_12833);
or U13232 (N_13232,N_12759,N_12967);
or U13233 (N_13233,N_12932,N_12921);
and U13234 (N_13234,N_12803,N_12905);
nand U13235 (N_13235,N_12870,N_12830);
and U13236 (N_13236,N_12963,N_12872);
or U13237 (N_13237,N_12924,N_12976);
nand U13238 (N_13238,N_12791,N_12752);
and U13239 (N_13239,N_12838,N_12990);
and U13240 (N_13240,N_12974,N_12807);
or U13241 (N_13241,N_12845,N_12959);
or U13242 (N_13242,N_12959,N_12806);
nand U13243 (N_13243,N_12853,N_12940);
nor U13244 (N_13244,N_12989,N_12813);
xor U13245 (N_13245,N_12965,N_12927);
nor U13246 (N_13246,N_12802,N_12787);
xnor U13247 (N_13247,N_12897,N_12825);
and U13248 (N_13248,N_12893,N_12967);
and U13249 (N_13249,N_12896,N_12755);
nand U13250 (N_13250,N_13035,N_13205);
nand U13251 (N_13251,N_13113,N_13057);
xor U13252 (N_13252,N_13081,N_13123);
nor U13253 (N_13253,N_13046,N_13031);
nor U13254 (N_13254,N_13236,N_13196);
or U13255 (N_13255,N_13029,N_13103);
or U13256 (N_13256,N_13239,N_13222);
nor U13257 (N_13257,N_13030,N_13091);
and U13258 (N_13258,N_13013,N_13096);
xor U13259 (N_13259,N_13130,N_13005);
nand U13260 (N_13260,N_13137,N_13145);
and U13261 (N_13261,N_13061,N_13182);
and U13262 (N_13262,N_13125,N_13008);
and U13263 (N_13263,N_13127,N_13120);
nor U13264 (N_13264,N_13178,N_13167);
and U13265 (N_13265,N_13230,N_13242);
nor U13266 (N_13266,N_13060,N_13179);
or U13267 (N_13267,N_13184,N_13101);
xor U13268 (N_13268,N_13105,N_13162);
or U13269 (N_13269,N_13075,N_13163);
nor U13270 (N_13270,N_13050,N_13233);
nand U13271 (N_13271,N_13033,N_13164);
nor U13272 (N_13272,N_13210,N_13224);
nand U13273 (N_13273,N_13128,N_13016);
nor U13274 (N_13274,N_13002,N_13149);
nor U13275 (N_13275,N_13191,N_13022);
nand U13276 (N_13276,N_13017,N_13122);
xnor U13277 (N_13277,N_13068,N_13218);
xor U13278 (N_13278,N_13148,N_13121);
or U13279 (N_13279,N_13048,N_13047);
and U13280 (N_13280,N_13161,N_13221);
nor U13281 (N_13281,N_13241,N_13194);
nand U13282 (N_13282,N_13216,N_13229);
nand U13283 (N_13283,N_13012,N_13098);
xor U13284 (N_13284,N_13054,N_13213);
nand U13285 (N_13285,N_13069,N_13155);
or U13286 (N_13286,N_13104,N_13131);
nor U13287 (N_13287,N_13073,N_13010);
nor U13288 (N_13288,N_13040,N_13110);
nor U13289 (N_13289,N_13052,N_13011);
nand U13290 (N_13290,N_13151,N_13154);
or U13291 (N_13291,N_13107,N_13070);
or U13292 (N_13292,N_13144,N_13238);
xor U13293 (N_13293,N_13193,N_13201);
xnor U13294 (N_13294,N_13206,N_13181);
nor U13295 (N_13295,N_13166,N_13077);
nand U13296 (N_13296,N_13001,N_13109);
or U13297 (N_13297,N_13247,N_13244);
nand U13298 (N_13298,N_13100,N_13039);
xnor U13299 (N_13299,N_13134,N_13102);
nand U13300 (N_13300,N_13049,N_13097);
xor U13301 (N_13301,N_13095,N_13099);
and U13302 (N_13302,N_13062,N_13129);
or U13303 (N_13303,N_13043,N_13118);
xor U13304 (N_13304,N_13237,N_13170);
or U13305 (N_13305,N_13115,N_13108);
and U13306 (N_13306,N_13158,N_13117);
nor U13307 (N_13307,N_13092,N_13018);
and U13308 (N_13308,N_13225,N_13183);
nor U13309 (N_13309,N_13177,N_13165);
nor U13310 (N_13310,N_13228,N_13037);
nand U13311 (N_13311,N_13156,N_13245);
or U13312 (N_13312,N_13126,N_13231);
nand U13313 (N_13313,N_13169,N_13024);
nand U13314 (N_13314,N_13084,N_13203);
or U13315 (N_13315,N_13195,N_13093);
or U13316 (N_13316,N_13065,N_13019);
nand U13317 (N_13317,N_13212,N_13157);
xor U13318 (N_13318,N_13078,N_13058);
nor U13319 (N_13319,N_13153,N_13133);
nor U13320 (N_13320,N_13168,N_13023);
nand U13321 (N_13321,N_13186,N_13176);
nand U13322 (N_13322,N_13066,N_13044);
xnor U13323 (N_13323,N_13234,N_13038);
and U13324 (N_13324,N_13006,N_13055);
xor U13325 (N_13325,N_13146,N_13042);
and U13326 (N_13326,N_13056,N_13159);
nand U13327 (N_13327,N_13000,N_13059);
and U13328 (N_13328,N_13076,N_13209);
xor U13329 (N_13329,N_13180,N_13207);
nor U13330 (N_13330,N_13211,N_13027);
xor U13331 (N_13331,N_13175,N_13135);
nand U13332 (N_13332,N_13020,N_13140);
and U13333 (N_13333,N_13032,N_13172);
nor U13334 (N_13334,N_13124,N_13051);
and U13335 (N_13335,N_13025,N_13246);
nor U13336 (N_13336,N_13111,N_13174);
nor U13337 (N_13337,N_13160,N_13226);
and U13338 (N_13338,N_13173,N_13026);
and U13339 (N_13339,N_13188,N_13119);
xor U13340 (N_13340,N_13009,N_13243);
nand U13341 (N_13341,N_13014,N_13190);
xor U13342 (N_13342,N_13034,N_13217);
or U13343 (N_13343,N_13132,N_13202);
or U13344 (N_13344,N_13094,N_13083);
xnor U13345 (N_13345,N_13041,N_13114);
nor U13346 (N_13346,N_13197,N_13204);
nand U13347 (N_13347,N_13189,N_13219);
or U13348 (N_13348,N_13064,N_13199);
xnor U13349 (N_13349,N_13086,N_13067);
xnor U13350 (N_13350,N_13232,N_13071);
or U13351 (N_13351,N_13089,N_13004);
xor U13352 (N_13352,N_13249,N_13080);
xor U13353 (N_13353,N_13053,N_13036);
xnor U13354 (N_13354,N_13141,N_13198);
or U13355 (N_13355,N_13015,N_13138);
xnor U13356 (N_13356,N_13116,N_13074);
nor U13357 (N_13357,N_13223,N_13087);
xor U13358 (N_13358,N_13028,N_13021);
xnor U13359 (N_13359,N_13106,N_13200);
or U13360 (N_13360,N_13227,N_13045);
xor U13361 (N_13361,N_13152,N_13139);
and U13362 (N_13362,N_13240,N_13142);
nor U13363 (N_13363,N_13192,N_13143);
and U13364 (N_13364,N_13085,N_13187);
and U13365 (N_13365,N_13215,N_13208);
nor U13366 (N_13366,N_13185,N_13248);
or U13367 (N_13367,N_13063,N_13082);
and U13368 (N_13368,N_13007,N_13112);
nand U13369 (N_13369,N_13220,N_13171);
xor U13370 (N_13370,N_13072,N_13003);
nor U13371 (N_13371,N_13150,N_13079);
nor U13372 (N_13372,N_13136,N_13090);
and U13373 (N_13373,N_13235,N_13214);
nor U13374 (N_13374,N_13088,N_13147);
nor U13375 (N_13375,N_13247,N_13207);
or U13376 (N_13376,N_13219,N_13073);
nor U13377 (N_13377,N_13034,N_13182);
and U13378 (N_13378,N_13044,N_13014);
or U13379 (N_13379,N_13144,N_13006);
nand U13380 (N_13380,N_13097,N_13084);
and U13381 (N_13381,N_13197,N_13099);
nand U13382 (N_13382,N_13220,N_13132);
nor U13383 (N_13383,N_13029,N_13171);
or U13384 (N_13384,N_13132,N_13179);
nand U13385 (N_13385,N_13225,N_13133);
xnor U13386 (N_13386,N_13104,N_13187);
and U13387 (N_13387,N_13056,N_13000);
or U13388 (N_13388,N_13010,N_13124);
or U13389 (N_13389,N_13207,N_13027);
or U13390 (N_13390,N_13123,N_13026);
or U13391 (N_13391,N_13181,N_13060);
nor U13392 (N_13392,N_13119,N_13220);
xor U13393 (N_13393,N_13187,N_13114);
nand U13394 (N_13394,N_13143,N_13019);
nor U13395 (N_13395,N_13209,N_13152);
nor U13396 (N_13396,N_13119,N_13137);
nand U13397 (N_13397,N_13068,N_13072);
nand U13398 (N_13398,N_13129,N_13090);
nand U13399 (N_13399,N_13115,N_13127);
and U13400 (N_13400,N_13162,N_13051);
nand U13401 (N_13401,N_13004,N_13105);
nor U13402 (N_13402,N_13107,N_13026);
nor U13403 (N_13403,N_13226,N_13219);
xnor U13404 (N_13404,N_13199,N_13127);
nand U13405 (N_13405,N_13155,N_13088);
nor U13406 (N_13406,N_13038,N_13136);
nor U13407 (N_13407,N_13245,N_13004);
xor U13408 (N_13408,N_13075,N_13021);
xnor U13409 (N_13409,N_13034,N_13152);
xor U13410 (N_13410,N_13190,N_13247);
or U13411 (N_13411,N_13244,N_13240);
nand U13412 (N_13412,N_13081,N_13143);
and U13413 (N_13413,N_13238,N_13087);
nand U13414 (N_13414,N_13217,N_13197);
and U13415 (N_13415,N_13187,N_13086);
xnor U13416 (N_13416,N_13081,N_13045);
xnor U13417 (N_13417,N_13014,N_13076);
xor U13418 (N_13418,N_13244,N_13051);
nor U13419 (N_13419,N_13107,N_13035);
and U13420 (N_13420,N_13008,N_13098);
nor U13421 (N_13421,N_13225,N_13244);
or U13422 (N_13422,N_13192,N_13091);
nand U13423 (N_13423,N_13237,N_13078);
nor U13424 (N_13424,N_13221,N_13100);
nor U13425 (N_13425,N_13121,N_13209);
and U13426 (N_13426,N_13055,N_13134);
nor U13427 (N_13427,N_13064,N_13229);
xor U13428 (N_13428,N_13238,N_13124);
and U13429 (N_13429,N_13070,N_13016);
xnor U13430 (N_13430,N_13122,N_13209);
xor U13431 (N_13431,N_13241,N_13108);
or U13432 (N_13432,N_13111,N_13011);
nand U13433 (N_13433,N_13156,N_13149);
xnor U13434 (N_13434,N_13072,N_13248);
and U13435 (N_13435,N_13183,N_13164);
and U13436 (N_13436,N_13172,N_13042);
or U13437 (N_13437,N_13191,N_13086);
xnor U13438 (N_13438,N_13244,N_13154);
and U13439 (N_13439,N_13113,N_13238);
xor U13440 (N_13440,N_13059,N_13091);
and U13441 (N_13441,N_13107,N_13089);
xor U13442 (N_13442,N_13068,N_13040);
and U13443 (N_13443,N_13248,N_13195);
or U13444 (N_13444,N_13080,N_13068);
nand U13445 (N_13445,N_13195,N_13011);
nand U13446 (N_13446,N_13107,N_13209);
and U13447 (N_13447,N_13187,N_13010);
nor U13448 (N_13448,N_13008,N_13080);
nor U13449 (N_13449,N_13211,N_13136);
nand U13450 (N_13450,N_13060,N_13049);
nor U13451 (N_13451,N_13213,N_13067);
nor U13452 (N_13452,N_13133,N_13042);
or U13453 (N_13453,N_13111,N_13140);
and U13454 (N_13454,N_13134,N_13026);
nand U13455 (N_13455,N_13175,N_13120);
xnor U13456 (N_13456,N_13037,N_13188);
and U13457 (N_13457,N_13041,N_13025);
nor U13458 (N_13458,N_13220,N_13043);
nand U13459 (N_13459,N_13143,N_13012);
nor U13460 (N_13460,N_13042,N_13219);
or U13461 (N_13461,N_13049,N_13239);
nand U13462 (N_13462,N_13049,N_13041);
or U13463 (N_13463,N_13101,N_13197);
or U13464 (N_13464,N_13111,N_13073);
xnor U13465 (N_13465,N_13138,N_13182);
and U13466 (N_13466,N_13099,N_13006);
and U13467 (N_13467,N_13149,N_13205);
xnor U13468 (N_13468,N_13017,N_13246);
and U13469 (N_13469,N_13053,N_13110);
and U13470 (N_13470,N_13137,N_13083);
xor U13471 (N_13471,N_13068,N_13125);
nor U13472 (N_13472,N_13102,N_13238);
nor U13473 (N_13473,N_13057,N_13078);
xnor U13474 (N_13474,N_13230,N_13243);
nand U13475 (N_13475,N_13114,N_13030);
nor U13476 (N_13476,N_13221,N_13145);
and U13477 (N_13477,N_13158,N_13232);
or U13478 (N_13478,N_13049,N_13023);
and U13479 (N_13479,N_13218,N_13114);
nor U13480 (N_13480,N_13156,N_13039);
xnor U13481 (N_13481,N_13077,N_13144);
nand U13482 (N_13482,N_13101,N_13077);
nand U13483 (N_13483,N_13144,N_13009);
nand U13484 (N_13484,N_13137,N_13243);
or U13485 (N_13485,N_13156,N_13053);
nor U13486 (N_13486,N_13246,N_13103);
nor U13487 (N_13487,N_13115,N_13024);
nand U13488 (N_13488,N_13056,N_13031);
nor U13489 (N_13489,N_13139,N_13186);
and U13490 (N_13490,N_13115,N_13063);
nand U13491 (N_13491,N_13175,N_13101);
and U13492 (N_13492,N_13157,N_13021);
and U13493 (N_13493,N_13027,N_13109);
nor U13494 (N_13494,N_13117,N_13067);
nor U13495 (N_13495,N_13074,N_13034);
nor U13496 (N_13496,N_13218,N_13147);
or U13497 (N_13497,N_13128,N_13083);
nand U13498 (N_13498,N_13164,N_13016);
and U13499 (N_13499,N_13232,N_13244);
nand U13500 (N_13500,N_13317,N_13499);
nand U13501 (N_13501,N_13301,N_13411);
and U13502 (N_13502,N_13388,N_13367);
and U13503 (N_13503,N_13310,N_13266);
or U13504 (N_13504,N_13382,N_13346);
and U13505 (N_13505,N_13291,N_13490);
xor U13506 (N_13506,N_13289,N_13304);
xnor U13507 (N_13507,N_13326,N_13274);
and U13508 (N_13508,N_13394,N_13488);
nor U13509 (N_13509,N_13416,N_13484);
or U13510 (N_13510,N_13327,N_13283);
nor U13511 (N_13511,N_13448,N_13487);
nand U13512 (N_13512,N_13443,N_13267);
nor U13513 (N_13513,N_13480,N_13251);
nor U13514 (N_13514,N_13427,N_13425);
xnor U13515 (N_13515,N_13282,N_13264);
xnor U13516 (N_13516,N_13308,N_13329);
or U13517 (N_13517,N_13356,N_13358);
nand U13518 (N_13518,N_13284,N_13397);
xor U13519 (N_13519,N_13258,N_13254);
xnor U13520 (N_13520,N_13319,N_13297);
or U13521 (N_13521,N_13440,N_13331);
nor U13522 (N_13522,N_13479,N_13260);
nand U13523 (N_13523,N_13300,N_13442);
xor U13524 (N_13524,N_13432,N_13469);
or U13525 (N_13525,N_13369,N_13379);
and U13526 (N_13526,N_13276,N_13475);
nand U13527 (N_13527,N_13390,N_13293);
nand U13528 (N_13528,N_13497,N_13426);
and U13529 (N_13529,N_13337,N_13383);
and U13530 (N_13530,N_13295,N_13363);
nand U13531 (N_13531,N_13465,N_13328);
or U13532 (N_13532,N_13320,N_13457);
xnor U13533 (N_13533,N_13306,N_13341);
or U13534 (N_13534,N_13431,N_13271);
and U13535 (N_13535,N_13384,N_13471);
or U13536 (N_13536,N_13424,N_13262);
nand U13537 (N_13537,N_13372,N_13287);
or U13538 (N_13538,N_13419,N_13491);
or U13539 (N_13539,N_13374,N_13313);
or U13540 (N_13540,N_13463,N_13415);
and U13541 (N_13541,N_13389,N_13458);
or U13542 (N_13542,N_13376,N_13268);
nand U13543 (N_13543,N_13477,N_13391);
nand U13544 (N_13544,N_13470,N_13429);
and U13545 (N_13545,N_13273,N_13485);
nor U13546 (N_13546,N_13279,N_13395);
or U13547 (N_13547,N_13323,N_13335);
nor U13548 (N_13548,N_13349,N_13343);
xor U13549 (N_13549,N_13298,N_13478);
and U13550 (N_13550,N_13338,N_13474);
and U13551 (N_13551,N_13422,N_13322);
nor U13552 (N_13552,N_13467,N_13406);
nand U13553 (N_13553,N_13378,N_13494);
and U13554 (N_13554,N_13350,N_13353);
or U13555 (N_13555,N_13370,N_13386);
xor U13556 (N_13556,N_13340,N_13348);
nand U13557 (N_13557,N_13318,N_13399);
or U13558 (N_13558,N_13272,N_13421);
nor U13559 (N_13559,N_13309,N_13437);
or U13560 (N_13560,N_13347,N_13364);
or U13561 (N_13561,N_13352,N_13316);
or U13562 (N_13562,N_13269,N_13430);
and U13563 (N_13563,N_13486,N_13441);
and U13564 (N_13564,N_13459,N_13359);
or U13565 (N_13565,N_13489,N_13250);
nor U13566 (N_13566,N_13344,N_13396);
nand U13567 (N_13567,N_13299,N_13366);
nand U13568 (N_13568,N_13407,N_13314);
nor U13569 (N_13569,N_13259,N_13288);
nor U13570 (N_13570,N_13414,N_13373);
nor U13571 (N_13571,N_13368,N_13290);
nand U13572 (N_13572,N_13434,N_13498);
and U13573 (N_13573,N_13265,N_13307);
or U13574 (N_13574,N_13454,N_13462);
and U13575 (N_13575,N_13452,N_13481);
and U13576 (N_13576,N_13357,N_13446);
and U13577 (N_13577,N_13493,N_13361);
xnor U13578 (N_13578,N_13375,N_13355);
nand U13579 (N_13579,N_13455,N_13345);
and U13580 (N_13580,N_13296,N_13403);
or U13581 (N_13581,N_13263,N_13377);
nand U13582 (N_13582,N_13435,N_13385);
nand U13583 (N_13583,N_13275,N_13354);
xor U13584 (N_13584,N_13408,N_13286);
and U13585 (N_13585,N_13444,N_13476);
xnor U13586 (N_13586,N_13339,N_13410);
nor U13587 (N_13587,N_13257,N_13402);
or U13588 (N_13588,N_13285,N_13492);
nor U13589 (N_13589,N_13302,N_13417);
or U13590 (N_13590,N_13398,N_13393);
nand U13591 (N_13591,N_13445,N_13447);
nor U13592 (N_13592,N_13253,N_13495);
xnor U13593 (N_13593,N_13433,N_13256);
xnor U13594 (N_13594,N_13336,N_13381);
or U13595 (N_13595,N_13333,N_13428);
nand U13596 (N_13596,N_13461,N_13371);
nand U13597 (N_13597,N_13451,N_13281);
xnor U13598 (N_13598,N_13292,N_13401);
or U13599 (N_13599,N_13466,N_13362);
nor U13600 (N_13600,N_13412,N_13473);
or U13601 (N_13601,N_13472,N_13305);
xnor U13602 (N_13602,N_13360,N_13332);
nand U13603 (N_13603,N_13409,N_13423);
nand U13604 (N_13604,N_13468,N_13325);
nand U13605 (N_13605,N_13464,N_13453);
or U13606 (N_13606,N_13436,N_13438);
nor U13607 (N_13607,N_13255,N_13413);
or U13608 (N_13608,N_13330,N_13270);
or U13609 (N_13609,N_13280,N_13439);
nand U13610 (N_13610,N_13261,N_13387);
xnor U13611 (N_13611,N_13483,N_13334);
or U13612 (N_13612,N_13482,N_13342);
and U13613 (N_13613,N_13303,N_13400);
xnor U13614 (N_13614,N_13312,N_13380);
xor U13615 (N_13615,N_13456,N_13496);
or U13616 (N_13616,N_13324,N_13404);
nor U13617 (N_13617,N_13405,N_13392);
or U13618 (N_13618,N_13449,N_13321);
and U13619 (N_13619,N_13311,N_13315);
nand U13620 (N_13620,N_13460,N_13365);
or U13621 (N_13621,N_13278,N_13294);
or U13622 (N_13622,N_13420,N_13450);
nor U13623 (N_13623,N_13277,N_13351);
nor U13624 (N_13624,N_13418,N_13252);
and U13625 (N_13625,N_13367,N_13472);
and U13626 (N_13626,N_13351,N_13393);
and U13627 (N_13627,N_13413,N_13335);
nand U13628 (N_13628,N_13252,N_13499);
xnor U13629 (N_13629,N_13282,N_13291);
nand U13630 (N_13630,N_13283,N_13256);
nand U13631 (N_13631,N_13300,N_13486);
and U13632 (N_13632,N_13270,N_13485);
and U13633 (N_13633,N_13457,N_13425);
xor U13634 (N_13634,N_13355,N_13274);
nor U13635 (N_13635,N_13327,N_13267);
nand U13636 (N_13636,N_13388,N_13466);
nand U13637 (N_13637,N_13461,N_13495);
nand U13638 (N_13638,N_13362,N_13288);
and U13639 (N_13639,N_13378,N_13325);
or U13640 (N_13640,N_13495,N_13283);
nand U13641 (N_13641,N_13384,N_13392);
and U13642 (N_13642,N_13475,N_13285);
or U13643 (N_13643,N_13304,N_13478);
and U13644 (N_13644,N_13394,N_13342);
nor U13645 (N_13645,N_13361,N_13452);
nand U13646 (N_13646,N_13412,N_13344);
or U13647 (N_13647,N_13413,N_13496);
or U13648 (N_13648,N_13383,N_13490);
xor U13649 (N_13649,N_13386,N_13348);
xor U13650 (N_13650,N_13329,N_13317);
nand U13651 (N_13651,N_13329,N_13388);
xor U13652 (N_13652,N_13478,N_13278);
nand U13653 (N_13653,N_13411,N_13392);
nor U13654 (N_13654,N_13385,N_13383);
or U13655 (N_13655,N_13289,N_13374);
and U13656 (N_13656,N_13256,N_13378);
nand U13657 (N_13657,N_13496,N_13321);
or U13658 (N_13658,N_13451,N_13397);
and U13659 (N_13659,N_13280,N_13436);
and U13660 (N_13660,N_13256,N_13297);
nor U13661 (N_13661,N_13341,N_13255);
or U13662 (N_13662,N_13341,N_13254);
and U13663 (N_13663,N_13355,N_13303);
or U13664 (N_13664,N_13267,N_13382);
and U13665 (N_13665,N_13443,N_13405);
xor U13666 (N_13666,N_13499,N_13368);
xor U13667 (N_13667,N_13308,N_13317);
and U13668 (N_13668,N_13333,N_13404);
and U13669 (N_13669,N_13466,N_13351);
or U13670 (N_13670,N_13308,N_13409);
nand U13671 (N_13671,N_13492,N_13281);
or U13672 (N_13672,N_13422,N_13347);
xor U13673 (N_13673,N_13318,N_13394);
or U13674 (N_13674,N_13354,N_13258);
nor U13675 (N_13675,N_13334,N_13380);
nand U13676 (N_13676,N_13251,N_13427);
nand U13677 (N_13677,N_13389,N_13415);
xor U13678 (N_13678,N_13432,N_13483);
and U13679 (N_13679,N_13296,N_13432);
or U13680 (N_13680,N_13255,N_13250);
nand U13681 (N_13681,N_13367,N_13354);
xor U13682 (N_13682,N_13411,N_13340);
nor U13683 (N_13683,N_13311,N_13483);
nor U13684 (N_13684,N_13320,N_13295);
or U13685 (N_13685,N_13446,N_13268);
nand U13686 (N_13686,N_13372,N_13361);
or U13687 (N_13687,N_13466,N_13276);
xor U13688 (N_13688,N_13298,N_13383);
xor U13689 (N_13689,N_13378,N_13391);
and U13690 (N_13690,N_13306,N_13261);
xor U13691 (N_13691,N_13323,N_13434);
nand U13692 (N_13692,N_13443,N_13276);
nand U13693 (N_13693,N_13466,N_13296);
or U13694 (N_13694,N_13467,N_13332);
and U13695 (N_13695,N_13282,N_13253);
or U13696 (N_13696,N_13337,N_13353);
nand U13697 (N_13697,N_13305,N_13448);
or U13698 (N_13698,N_13426,N_13341);
xor U13699 (N_13699,N_13466,N_13391);
xnor U13700 (N_13700,N_13280,N_13373);
xor U13701 (N_13701,N_13305,N_13317);
nand U13702 (N_13702,N_13329,N_13495);
and U13703 (N_13703,N_13321,N_13272);
xor U13704 (N_13704,N_13386,N_13399);
nor U13705 (N_13705,N_13489,N_13468);
and U13706 (N_13706,N_13407,N_13301);
nand U13707 (N_13707,N_13436,N_13343);
xor U13708 (N_13708,N_13378,N_13277);
and U13709 (N_13709,N_13470,N_13288);
and U13710 (N_13710,N_13393,N_13392);
or U13711 (N_13711,N_13390,N_13369);
and U13712 (N_13712,N_13392,N_13472);
nor U13713 (N_13713,N_13410,N_13320);
or U13714 (N_13714,N_13287,N_13308);
nand U13715 (N_13715,N_13436,N_13465);
xor U13716 (N_13716,N_13386,N_13403);
nor U13717 (N_13717,N_13369,N_13422);
and U13718 (N_13718,N_13384,N_13462);
nor U13719 (N_13719,N_13261,N_13379);
and U13720 (N_13720,N_13493,N_13356);
or U13721 (N_13721,N_13342,N_13456);
nand U13722 (N_13722,N_13434,N_13389);
nor U13723 (N_13723,N_13319,N_13289);
or U13724 (N_13724,N_13492,N_13407);
or U13725 (N_13725,N_13355,N_13338);
nor U13726 (N_13726,N_13458,N_13251);
or U13727 (N_13727,N_13419,N_13362);
nand U13728 (N_13728,N_13316,N_13317);
or U13729 (N_13729,N_13466,N_13344);
xor U13730 (N_13730,N_13342,N_13483);
nor U13731 (N_13731,N_13328,N_13482);
and U13732 (N_13732,N_13319,N_13461);
or U13733 (N_13733,N_13393,N_13329);
and U13734 (N_13734,N_13262,N_13423);
nand U13735 (N_13735,N_13256,N_13326);
or U13736 (N_13736,N_13290,N_13491);
or U13737 (N_13737,N_13461,N_13321);
nand U13738 (N_13738,N_13326,N_13387);
and U13739 (N_13739,N_13320,N_13348);
nor U13740 (N_13740,N_13388,N_13427);
and U13741 (N_13741,N_13455,N_13307);
nand U13742 (N_13742,N_13484,N_13322);
nand U13743 (N_13743,N_13385,N_13261);
nand U13744 (N_13744,N_13478,N_13344);
nand U13745 (N_13745,N_13372,N_13343);
or U13746 (N_13746,N_13479,N_13398);
nand U13747 (N_13747,N_13333,N_13396);
xnor U13748 (N_13748,N_13437,N_13488);
nand U13749 (N_13749,N_13442,N_13477);
and U13750 (N_13750,N_13523,N_13735);
nor U13751 (N_13751,N_13619,N_13697);
xnor U13752 (N_13752,N_13514,N_13685);
and U13753 (N_13753,N_13694,N_13666);
xnor U13754 (N_13754,N_13642,N_13670);
and U13755 (N_13755,N_13576,N_13547);
nand U13756 (N_13756,N_13597,N_13638);
and U13757 (N_13757,N_13627,N_13655);
and U13758 (N_13758,N_13601,N_13609);
or U13759 (N_13759,N_13636,N_13543);
xnor U13760 (N_13760,N_13553,N_13663);
or U13761 (N_13761,N_13503,N_13709);
or U13762 (N_13762,N_13667,N_13527);
nand U13763 (N_13763,N_13644,N_13589);
nor U13764 (N_13764,N_13530,N_13749);
or U13765 (N_13765,N_13593,N_13725);
nor U13766 (N_13766,N_13595,N_13511);
nand U13767 (N_13767,N_13508,N_13538);
and U13768 (N_13768,N_13591,N_13632);
and U13769 (N_13769,N_13654,N_13677);
nor U13770 (N_13770,N_13738,N_13552);
nor U13771 (N_13771,N_13696,N_13698);
and U13772 (N_13772,N_13599,N_13711);
xor U13773 (N_13773,N_13580,N_13611);
xor U13774 (N_13774,N_13742,N_13545);
nor U13775 (N_13775,N_13639,N_13641);
nand U13776 (N_13776,N_13645,N_13557);
nor U13777 (N_13777,N_13505,N_13544);
xnor U13778 (N_13778,N_13731,N_13526);
or U13779 (N_13779,N_13693,N_13634);
nand U13780 (N_13780,N_13512,N_13703);
or U13781 (N_13781,N_13626,N_13586);
nand U13782 (N_13782,N_13722,N_13567);
xnor U13783 (N_13783,N_13525,N_13743);
xnor U13784 (N_13784,N_13571,N_13578);
nor U13785 (N_13785,N_13603,N_13605);
nor U13786 (N_13786,N_13748,N_13649);
nor U13787 (N_13787,N_13695,N_13665);
or U13788 (N_13788,N_13551,N_13513);
nor U13789 (N_13789,N_13614,N_13729);
xor U13790 (N_13790,N_13646,N_13708);
or U13791 (N_13791,N_13653,N_13561);
nand U13792 (N_13792,N_13688,N_13741);
or U13793 (N_13793,N_13621,N_13707);
nand U13794 (N_13794,N_13562,N_13504);
nor U13795 (N_13795,N_13723,N_13628);
nand U13796 (N_13796,N_13579,N_13592);
or U13797 (N_13797,N_13712,N_13509);
or U13798 (N_13798,N_13684,N_13582);
nand U13799 (N_13799,N_13568,N_13705);
nand U13800 (N_13800,N_13662,N_13651);
xor U13801 (N_13801,N_13532,N_13733);
and U13802 (N_13802,N_13515,N_13726);
nor U13803 (N_13803,N_13602,N_13518);
nor U13804 (N_13804,N_13629,N_13550);
or U13805 (N_13805,N_13507,N_13565);
xnor U13806 (N_13806,N_13554,N_13531);
nor U13807 (N_13807,N_13572,N_13623);
nor U13808 (N_13808,N_13637,N_13574);
nor U13809 (N_13809,N_13540,N_13613);
or U13810 (N_13810,N_13690,N_13564);
or U13811 (N_13811,N_13702,N_13717);
or U13812 (N_13812,N_13687,N_13546);
xnor U13813 (N_13813,N_13535,N_13672);
xnor U13814 (N_13814,N_13700,N_13630);
xor U13815 (N_13815,N_13747,N_13529);
and U13816 (N_13816,N_13563,N_13519);
nor U13817 (N_13817,N_13541,N_13676);
or U13818 (N_13818,N_13724,N_13617);
and U13819 (N_13819,N_13622,N_13596);
or U13820 (N_13820,N_13674,N_13657);
xor U13821 (N_13821,N_13739,N_13701);
xor U13822 (N_13822,N_13668,N_13522);
or U13823 (N_13823,N_13732,N_13631);
and U13824 (N_13824,N_13692,N_13615);
or U13825 (N_13825,N_13587,N_13521);
and U13826 (N_13826,N_13608,N_13656);
and U13827 (N_13827,N_13502,N_13664);
and U13828 (N_13828,N_13682,N_13585);
nor U13829 (N_13829,N_13607,N_13710);
or U13830 (N_13830,N_13620,N_13549);
and U13831 (N_13831,N_13577,N_13612);
xor U13832 (N_13832,N_13746,N_13689);
nor U13833 (N_13833,N_13618,N_13647);
nor U13834 (N_13834,N_13575,N_13673);
nand U13835 (N_13835,N_13536,N_13660);
or U13836 (N_13836,N_13730,N_13658);
or U13837 (N_13837,N_13686,N_13624);
nor U13838 (N_13838,N_13643,N_13734);
or U13839 (N_13839,N_13610,N_13745);
and U13840 (N_13840,N_13669,N_13716);
or U13841 (N_13841,N_13566,N_13555);
nor U13842 (N_13842,N_13594,N_13537);
xor U13843 (N_13843,N_13583,N_13652);
or U13844 (N_13844,N_13625,N_13661);
or U13845 (N_13845,N_13727,N_13501);
xnor U13846 (N_13846,N_13539,N_13606);
and U13847 (N_13847,N_13715,N_13560);
xnor U13848 (N_13848,N_13534,N_13720);
xnor U13849 (N_13849,N_13581,N_13604);
nand U13850 (N_13850,N_13570,N_13650);
xnor U13851 (N_13851,N_13680,N_13516);
nor U13852 (N_13852,N_13648,N_13744);
or U13853 (N_13853,N_13713,N_13584);
xor U13854 (N_13854,N_13728,N_13548);
xor U13855 (N_13855,N_13737,N_13506);
nand U13856 (N_13856,N_13691,N_13600);
or U13857 (N_13857,N_13699,N_13500);
or U13858 (N_13858,N_13520,N_13714);
or U13859 (N_13859,N_13569,N_13659);
nor U13860 (N_13860,N_13524,N_13598);
and U13861 (N_13861,N_13740,N_13671);
and U13862 (N_13862,N_13556,N_13542);
nand U13863 (N_13863,N_13588,N_13706);
or U13864 (N_13864,N_13718,N_13719);
or U13865 (N_13865,N_13510,N_13633);
nand U13866 (N_13866,N_13640,N_13616);
nor U13867 (N_13867,N_13528,N_13573);
and U13868 (N_13868,N_13704,N_13736);
and U13869 (N_13869,N_13558,N_13679);
or U13870 (N_13870,N_13683,N_13533);
xnor U13871 (N_13871,N_13590,N_13635);
and U13872 (N_13872,N_13675,N_13559);
nand U13873 (N_13873,N_13678,N_13721);
and U13874 (N_13874,N_13681,N_13517);
or U13875 (N_13875,N_13650,N_13589);
or U13876 (N_13876,N_13644,N_13525);
and U13877 (N_13877,N_13597,N_13647);
xnor U13878 (N_13878,N_13643,N_13629);
xor U13879 (N_13879,N_13696,N_13675);
and U13880 (N_13880,N_13561,N_13735);
nand U13881 (N_13881,N_13553,N_13706);
and U13882 (N_13882,N_13686,N_13667);
or U13883 (N_13883,N_13584,N_13643);
nor U13884 (N_13884,N_13668,N_13638);
and U13885 (N_13885,N_13733,N_13743);
xor U13886 (N_13886,N_13638,N_13573);
or U13887 (N_13887,N_13674,N_13512);
nand U13888 (N_13888,N_13657,N_13503);
xnor U13889 (N_13889,N_13595,N_13656);
nor U13890 (N_13890,N_13548,N_13738);
or U13891 (N_13891,N_13598,N_13552);
nand U13892 (N_13892,N_13669,N_13652);
xnor U13893 (N_13893,N_13730,N_13578);
xnor U13894 (N_13894,N_13559,N_13508);
or U13895 (N_13895,N_13599,N_13600);
and U13896 (N_13896,N_13648,N_13605);
or U13897 (N_13897,N_13555,N_13650);
and U13898 (N_13898,N_13719,N_13715);
and U13899 (N_13899,N_13715,N_13559);
and U13900 (N_13900,N_13590,N_13503);
or U13901 (N_13901,N_13521,N_13620);
or U13902 (N_13902,N_13727,N_13557);
or U13903 (N_13903,N_13606,N_13535);
and U13904 (N_13904,N_13697,N_13507);
or U13905 (N_13905,N_13526,N_13519);
xor U13906 (N_13906,N_13723,N_13742);
nand U13907 (N_13907,N_13695,N_13521);
and U13908 (N_13908,N_13730,N_13688);
nor U13909 (N_13909,N_13617,N_13723);
or U13910 (N_13910,N_13522,N_13693);
and U13911 (N_13911,N_13652,N_13687);
or U13912 (N_13912,N_13671,N_13655);
xnor U13913 (N_13913,N_13593,N_13517);
xnor U13914 (N_13914,N_13524,N_13653);
and U13915 (N_13915,N_13657,N_13714);
xnor U13916 (N_13916,N_13708,N_13681);
and U13917 (N_13917,N_13560,N_13672);
xor U13918 (N_13918,N_13596,N_13690);
nor U13919 (N_13919,N_13596,N_13550);
nand U13920 (N_13920,N_13561,N_13703);
or U13921 (N_13921,N_13703,N_13705);
and U13922 (N_13922,N_13537,N_13728);
nor U13923 (N_13923,N_13546,N_13560);
or U13924 (N_13924,N_13732,N_13668);
nand U13925 (N_13925,N_13673,N_13612);
or U13926 (N_13926,N_13604,N_13611);
nand U13927 (N_13927,N_13639,N_13714);
nand U13928 (N_13928,N_13618,N_13747);
and U13929 (N_13929,N_13596,N_13667);
or U13930 (N_13930,N_13687,N_13507);
and U13931 (N_13931,N_13616,N_13577);
nand U13932 (N_13932,N_13561,N_13529);
nor U13933 (N_13933,N_13543,N_13678);
nand U13934 (N_13934,N_13603,N_13667);
or U13935 (N_13935,N_13739,N_13696);
nor U13936 (N_13936,N_13550,N_13567);
nor U13937 (N_13937,N_13718,N_13529);
xor U13938 (N_13938,N_13596,N_13577);
nand U13939 (N_13939,N_13600,N_13703);
nor U13940 (N_13940,N_13743,N_13529);
nand U13941 (N_13941,N_13542,N_13746);
or U13942 (N_13942,N_13743,N_13520);
or U13943 (N_13943,N_13670,N_13679);
nand U13944 (N_13944,N_13685,N_13626);
nor U13945 (N_13945,N_13582,N_13533);
nor U13946 (N_13946,N_13645,N_13582);
xor U13947 (N_13947,N_13659,N_13522);
nand U13948 (N_13948,N_13601,N_13661);
nor U13949 (N_13949,N_13651,N_13501);
or U13950 (N_13950,N_13555,N_13631);
nand U13951 (N_13951,N_13686,N_13571);
and U13952 (N_13952,N_13711,N_13665);
or U13953 (N_13953,N_13500,N_13720);
and U13954 (N_13954,N_13713,N_13686);
xnor U13955 (N_13955,N_13704,N_13526);
and U13956 (N_13956,N_13709,N_13552);
or U13957 (N_13957,N_13547,N_13601);
or U13958 (N_13958,N_13506,N_13667);
and U13959 (N_13959,N_13663,N_13651);
nand U13960 (N_13960,N_13642,N_13719);
nand U13961 (N_13961,N_13503,N_13644);
or U13962 (N_13962,N_13730,N_13541);
nand U13963 (N_13963,N_13746,N_13743);
and U13964 (N_13964,N_13539,N_13572);
nor U13965 (N_13965,N_13646,N_13727);
xor U13966 (N_13966,N_13513,N_13705);
nand U13967 (N_13967,N_13665,N_13636);
nor U13968 (N_13968,N_13509,N_13729);
and U13969 (N_13969,N_13651,N_13673);
nand U13970 (N_13970,N_13611,N_13747);
or U13971 (N_13971,N_13613,N_13726);
and U13972 (N_13972,N_13562,N_13604);
and U13973 (N_13973,N_13522,N_13517);
nand U13974 (N_13974,N_13656,N_13674);
nor U13975 (N_13975,N_13646,N_13734);
xor U13976 (N_13976,N_13737,N_13710);
xnor U13977 (N_13977,N_13673,N_13611);
and U13978 (N_13978,N_13539,N_13598);
xnor U13979 (N_13979,N_13745,N_13727);
xnor U13980 (N_13980,N_13741,N_13532);
nor U13981 (N_13981,N_13570,N_13744);
or U13982 (N_13982,N_13563,N_13702);
and U13983 (N_13983,N_13540,N_13589);
nor U13984 (N_13984,N_13745,N_13616);
nand U13985 (N_13985,N_13567,N_13736);
nor U13986 (N_13986,N_13626,N_13610);
or U13987 (N_13987,N_13700,N_13726);
xnor U13988 (N_13988,N_13714,N_13617);
nor U13989 (N_13989,N_13510,N_13702);
xor U13990 (N_13990,N_13631,N_13626);
xor U13991 (N_13991,N_13657,N_13646);
nor U13992 (N_13992,N_13671,N_13587);
and U13993 (N_13993,N_13652,N_13654);
or U13994 (N_13994,N_13637,N_13515);
or U13995 (N_13995,N_13660,N_13539);
nand U13996 (N_13996,N_13701,N_13643);
nand U13997 (N_13997,N_13719,N_13703);
and U13998 (N_13998,N_13721,N_13578);
or U13999 (N_13999,N_13701,N_13583);
xor U14000 (N_14000,N_13934,N_13955);
nand U14001 (N_14001,N_13973,N_13835);
and U14002 (N_14002,N_13849,N_13996);
xnor U14003 (N_14003,N_13923,N_13952);
nand U14004 (N_14004,N_13853,N_13788);
xor U14005 (N_14005,N_13886,N_13761);
or U14006 (N_14006,N_13990,N_13994);
xnor U14007 (N_14007,N_13960,N_13899);
and U14008 (N_14008,N_13961,N_13829);
nand U14009 (N_14009,N_13792,N_13757);
and U14010 (N_14010,N_13765,N_13917);
nor U14011 (N_14011,N_13755,N_13863);
nand U14012 (N_14012,N_13866,N_13876);
or U14013 (N_14013,N_13779,N_13971);
nand U14014 (N_14014,N_13776,N_13869);
or U14015 (N_14015,N_13847,N_13772);
or U14016 (N_14016,N_13967,N_13893);
and U14017 (N_14017,N_13770,N_13984);
xnor U14018 (N_14018,N_13995,N_13965);
and U14019 (N_14019,N_13766,N_13904);
nor U14020 (N_14020,N_13762,N_13824);
or U14021 (N_14021,N_13812,N_13848);
xor U14022 (N_14022,N_13936,N_13997);
nand U14023 (N_14023,N_13796,N_13868);
nor U14024 (N_14024,N_13999,N_13875);
and U14025 (N_14025,N_13873,N_13989);
xor U14026 (N_14026,N_13887,N_13938);
nor U14027 (N_14027,N_13906,N_13845);
xor U14028 (N_14028,N_13833,N_13787);
or U14029 (N_14029,N_13902,N_13985);
nand U14030 (N_14030,N_13993,N_13974);
xor U14031 (N_14031,N_13806,N_13756);
nand U14032 (N_14032,N_13856,N_13920);
xor U14033 (N_14033,N_13850,N_13861);
or U14034 (N_14034,N_13924,N_13977);
nand U14035 (N_14035,N_13872,N_13794);
nand U14036 (N_14036,N_13910,N_13839);
nor U14037 (N_14037,N_13947,N_13752);
or U14038 (N_14038,N_13981,N_13817);
nand U14039 (N_14039,N_13793,N_13771);
xnor U14040 (N_14040,N_13805,N_13807);
nor U14041 (N_14041,N_13828,N_13908);
nand U14042 (N_14042,N_13836,N_13754);
xor U14043 (N_14043,N_13922,N_13918);
nor U14044 (N_14044,N_13825,N_13851);
xnor U14045 (N_14045,N_13940,N_13804);
nand U14046 (N_14046,N_13956,N_13950);
and U14047 (N_14047,N_13857,N_13919);
nor U14048 (N_14048,N_13798,N_13820);
xnor U14049 (N_14049,N_13890,N_13927);
and U14050 (N_14050,N_13987,N_13784);
or U14051 (N_14051,N_13946,N_13903);
nand U14052 (N_14052,N_13888,N_13852);
or U14053 (N_14053,N_13943,N_13885);
or U14054 (N_14054,N_13978,N_13858);
and U14055 (N_14055,N_13799,N_13813);
nor U14056 (N_14056,N_13895,N_13912);
nor U14057 (N_14057,N_13891,N_13992);
nand U14058 (N_14058,N_13838,N_13972);
xnor U14059 (N_14059,N_13878,N_13864);
nor U14060 (N_14060,N_13773,N_13941);
xor U14061 (N_14061,N_13871,N_13818);
and U14062 (N_14062,N_13951,N_13968);
and U14063 (N_14063,N_13859,N_13827);
and U14064 (N_14064,N_13803,N_13763);
nor U14065 (N_14065,N_13898,N_13998);
xor U14066 (N_14066,N_13877,N_13775);
or U14067 (N_14067,N_13892,N_13790);
or U14068 (N_14068,N_13831,N_13783);
or U14069 (N_14069,N_13800,N_13778);
nor U14070 (N_14070,N_13764,N_13916);
nand U14071 (N_14071,N_13808,N_13907);
nor U14072 (N_14072,N_13911,N_13809);
nor U14073 (N_14073,N_13982,N_13976);
nor U14074 (N_14074,N_13867,N_13840);
xnor U14075 (N_14075,N_13959,N_13963);
and U14076 (N_14076,N_13983,N_13780);
nand U14077 (N_14077,N_13789,N_13930);
xnor U14078 (N_14078,N_13944,N_13901);
or U14079 (N_14079,N_13913,N_13921);
and U14080 (N_14080,N_13884,N_13969);
nor U14081 (N_14081,N_13966,N_13882);
or U14082 (N_14082,N_13929,N_13782);
or U14083 (N_14083,N_13914,N_13957);
xnor U14084 (N_14084,N_13988,N_13958);
and U14085 (N_14085,N_13881,N_13862);
nor U14086 (N_14086,N_13844,N_13964);
or U14087 (N_14087,N_13865,N_13953);
or U14088 (N_14088,N_13925,N_13874);
nor U14089 (N_14089,N_13843,N_13880);
nand U14090 (N_14090,N_13774,N_13785);
nor U14091 (N_14091,N_13948,N_13889);
or U14092 (N_14092,N_13980,N_13854);
xnor U14093 (N_14093,N_13819,N_13933);
xnor U14094 (N_14094,N_13786,N_13797);
nand U14095 (N_14095,N_13768,N_13928);
nor U14096 (N_14096,N_13962,N_13896);
nor U14097 (N_14097,N_13935,N_13769);
xnor U14098 (N_14098,N_13970,N_13814);
nand U14099 (N_14099,N_13897,N_13759);
or U14100 (N_14100,N_13801,N_13846);
or U14101 (N_14101,N_13791,N_13810);
or U14102 (N_14102,N_13870,N_13894);
nor U14103 (N_14103,N_13823,N_13781);
nor U14104 (N_14104,N_13860,N_13931);
xnor U14105 (N_14105,N_13777,N_13841);
xnor U14106 (N_14106,N_13937,N_13816);
or U14107 (N_14107,N_13945,N_13767);
nor U14108 (N_14108,N_13883,N_13900);
nand U14109 (N_14109,N_13909,N_13954);
nand U14110 (N_14110,N_13815,N_13842);
nand U14111 (N_14111,N_13979,N_13822);
xor U14112 (N_14112,N_13986,N_13932);
and U14113 (N_14113,N_13802,N_13832);
and U14114 (N_14114,N_13942,N_13821);
nor U14115 (N_14115,N_13905,N_13991);
nor U14116 (N_14116,N_13926,N_13915);
nand U14117 (N_14117,N_13826,N_13975);
nand U14118 (N_14118,N_13830,N_13939);
xor U14119 (N_14119,N_13795,N_13855);
or U14120 (N_14120,N_13811,N_13834);
nor U14121 (N_14121,N_13751,N_13949);
xor U14122 (N_14122,N_13758,N_13837);
or U14123 (N_14123,N_13753,N_13760);
nand U14124 (N_14124,N_13750,N_13879);
or U14125 (N_14125,N_13824,N_13852);
and U14126 (N_14126,N_13786,N_13992);
nor U14127 (N_14127,N_13906,N_13865);
nor U14128 (N_14128,N_13801,N_13756);
nor U14129 (N_14129,N_13866,N_13753);
and U14130 (N_14130,N_13942,N_13886);
and U14131 (N_14131,N_13965,N_13830);
nand U14132 (N_14132,N_13913,N_13783);
or U14133 (N_14133,N_13964,N_13816);
nand U14134 (N_14134,N_13976,N_13885);
nand U14135 (N_14135,N_13878,N_13920);
xor U14136 (N_14136,N_13762,N_13879);
or U14137 (N_14137,N_13828,N_13776);
xnor U14138 (N_14138,N_13759,N_13892);
nand U14139 (N_14139,N_13997,N_13831);
nor U14140 (N_14140,N_13841,N_13933);
and U14141 (N_14141,N_13976,N_13990);
nand U14142 (N_14142,N_13751,N_13839);
and U14143 (N_14143,N_13963,N_13793);
xor U14144 (N_14144,N_13851,N_13984);
nor U14145 (N_14145,N_13990,N_13796);
nor U14146 (N_14146,N_13787,N_13797);
and U14147 (N_14147,N_13758,N_13783);
xor U14148 (N_14148,N_13882,N_13965);
nor U14149 (N_14149,N_13874,N_13858);
xor U14150 (N_14150,N_13818,N_13833);
nor U14151 (N_14151,N_13930,N_13845);
nand U14152 (N_14152,N_13758,N_13796);
nor U14153 (N_14153,N_13771,N_13813);
or U14154 (N_14154,N_13814,N_13832);
nor U14155 (N_14155,N_13810,N_13930);
xnor U14156 (N_14156,N_13804,N_13986);
xnor U14157 (N_14157,N_13989,N_13805);
or U14158 (N_14158,N_13962,N_13939);
or U14159 (N_14159,N_13896,N_13868);
xnor U14160 (N_14160,N_13862,N_13807);
nand U14161 (N_14161,N_13956,N_13869);
xnor U14162 (N_14162,N_13864,N_13915);
or U14163 (N_14163,N_13899,N_13873);
or U14164 (N_14164,N_13902,N_13915);
and U14165 (N_14165,N_13951,N_13852);
nor U14166 (N_14166,N_13932,N_13765);
and U14167 (N_14167,N_13939,N_13941);
or U14168 (N_14168,N_13996,N_13862);
nand U14169 (N_14169,N_13763,N_13950);
and U14170 (N_14170,N_13985,N_13967);
nor U14171 (N_14171,N_13816,N_13998);
nor U14172 (N_14172,N_13796,N_13926);
and U14173 (N_14173,N_13892,N_13765);
xor U14174 (N_14174,N_13902,N_13756);
nor U14175 (N_14175,N_13850,N_13783);
nand U14176 (N_14176,N_13878,N_13831);
xnor U14177 (N_14177,N_13821,N_13991);
and U14178 (N_14178,N_13828,N_13844);
nand U14179 (N_14179,N_13929,N_13888);
nand U14180 (N_14180,N_13949,N_13998);
nand U14181 (N_14181,N_13976,N_13924);
xor U14182 (N_14182,N_13926,N_13887);
xnor U14183 (N_14183,N_13910,N_13797);
and U14184 (N_14184,N_13971,N_13942);
or U14185 (N_14185,N_13759,N_13867);
or U14186 (N_14186,N_13855,N_13843);
nor U14187 (N_14187,N_13806,N_13851);
and U14188 (N_14188,N_13815,N_13938);
nor U14189 (N_14189,N_13991,N_13938);
and U14190 (N_14190,N_13905,N_13759);
or U14191 (N_14191,N_13878,N_13932);
or U14192 (N_14192,N_13753,N_13800);
xnor U14193 (N_14193,N_13940,N_13884);
xor U14194 (N_14194,N_13967,N_13754);
and U14195 (N_14195,N_13899,N_13967);
xor U14196 (N_14196,N_13943,N_13776);
xor U14197 (N_14197,N_13935,N_13995);
xnor U14198 (N_14198,N_13769,N_13899);
xnor U14199 (N_14199,N_13812,N_13971);
and U14200 (N_14200,N_13808,N_13990);
xor U14201 (N_14201,N_13949,N_13778);
nand U14202 (N_14202,N_13857,N_13964);
nor U14203 (N_14203,N_13891,N_13876);
and U14204 (N_14204,N_13856,N_13776);
and U14205 (N_14205,N_13856,N_13969);
and U14206 (N_14206,N_13763,N_13962);
nand U14207 (N_14207,N_13919,N_13896);
xnor U14208 (N_14208,N_13930,N_13948);
or U14209 (N_14209,N_13907,N_13830);
or U14210 (N_14210,N_13965,N_13864);
nor U14211 (N_14211,N_13940,N_13851);
nand U14212 (N_14212,N_13762,N_13798);
xnor U14213 (N_14213,N_13957,N_13792);
and U14214 (N_14214,N_13979,N_13886);
and U14215 (N_14215,N_13898,N_13874);
or U14216 (N_14216,N_13942,N_13957);
or U14217 (N_14217,N_13883,N_13921);
nor U14218 (N_14218,N_13895,N_13817);
nand U14219 (N_14219,N_13944,N_13946);
xnor U14220 (N_14220,N_13851,N_13818);
and U14221 (N_14221,N_13926,N_13968);
nor U14222 (N_14222,N_13890,N_13933);
and U14223 (N_14223,N_13897,N_13905);
and U14224 (N_14224,N_13795,N_13754);
and U14225 (N_14225,N_13808,N_13860);
nor U14226 (N_14226,N_13843,N_13863);
or U14227 (N_14227,N_13899,N_13767);
nor U14228 (N_14228,N_13809,N_13771);
and U14229 (N_14229,N_13801,N_13932);
xnor U14230 (N_14230,N_13916,N_13813);
nor U14231 (N_14231,N_13840,N_13857);
or U14232 (N_14232,N_13953,N_13896);
xor U14233 (N_14233,N_13817,N_13980);
nor U14234 (N_14234,N_13838,N_13753);
nand U14235 (N_14235,N_13789,N_13924);
and U14236 (N_14236,N_13810,N_13989);
xor U14237 (N_14237,N_13779,N_13947);
xnor U14238 (N_14238,N_13916,N_13781);
and U14239 (N_14239,N_13800,N_13755);
nand U14240 (N_14240,N_13815,N_13865);
nand U14241 (N_14241,N_13761,N_13921);
nand U14242 (N_14242,N_13864,N_13794);
xnor U14243 (N_14243,N_13984,N_13756);
nand U14244 (N_14244,N_13830,N_13792);
nor U14245 (N_14245,N_13808,N_13937);
nand U14246 (N_14246,N_13821,N_13977);
xnor U14247 (N_14247,N_13849,N_13814);
or U14248 (N_14248,N_13752,N_13764);
xnor U14249 (N_14249,N_13847,N_13766);
and U14250 (N_14250,N_14139,N_14099);
and U14251 (N_14251,N_14238,N_14243);
nor U14252 (N_14252,N_14098,N_14244);
or U14253 (N_14253,N_14031,N_14202);
and U14254 (N_14254,N_14229,N_14095);
xor U14255 (N_14255,N_14072,N_14221);
xnor U14256 (N_14256,N_14154,N_14125);
xnor U14257 (N_14257,N_14005,N_14194);
or U14258 (N_14258,N_14132,N_14135);
xor U14259 (N_14259,N_14228,N_14220);
or U14260 (N_14260,N_14199,N_14163);
nand U14261 (N_14261,N_14114,N_14054);
nor U14262 (N_14262,N_14060,N_14235);
nor U14263 (N_14263,N_14128,N_14211);
nand U14264 (N_14264,N_14152,N_14166);
nand U14265 (N_14265,N_14171,N_14102);
or U14266 (N_14266,N_14115,N_14119);
nor U14267 (N_14267,N_14028,N_14067);
nor U14268 (N_14268,N_14144,N_14065);
or U14269 (N_14269,N_14037,N_14107);
nand U14270 (N_14270,N_14232,N_14162);
nand U14271 (N_14271,N_14129,N_14160);
nand U14272 (N_14272,N_14070,N_14140);
or U14273 (N_14273,N_14161,N_14069);
nor U14274 (N_14274,N_14094,N_14055);
xor U14275 (N_14275,N_14155,N_14145);
nand U14276 (N_14276,N_14214,N_14230);
or U14277 (N_14277,N_14193,N_14225);
nor U14278 (N_14278,N_14105,N_14175);
or U14279 (N_14279,N_14173,N_14180);
and U14280 (N_14280,N_14071,N_14036);
nor U14281 (N_14281,N_14052,N_14158);
or U14282 (N_14282,N_14127,N_14130);
nor U14283 (N_14283,N_14233,N_14026);
nand U14284 (N_14284,N_14078,N_14149);
or U14285 (N_14285,N_14117,N_14020);
or U14286 (N_14286,N_14062,N_14208);
nand U14287 (N_14287,N_14148,N_14027);
and U14288 (N_14288,N_14190,N_14196);
xor U14289 (N_14289,N_14041,N_14172);
or U14290 (N_14290,N_14147,N_14164);
nor U14291 (N_14291,N_14137,N_14116);
or U14292 (N_14292,N_14122,N_14092);
nor U14293 (N_14293,N_14080,N_14151);
nand U14294 (N_14294,N_14030,N_14146);
xnor U14295 (N_14295,N_14111,N_14168);
nor U14296 (N_14296,N_14059,N_14006);
xor U14297 (N_14297,N_14010,N_14112);
and U14298 (N_14298,N_14003,N_14035);
or U14299 (N_14299,N_14204,N_14106);
and U14300 (N_14300,N_14017,N_14206);
or U14301 (N_14301,N_14091,N_14187);
or U14302 (N_14302,N_14231,N_14077);
xor U14303 (N_14303,N_14002,N_14234);
or U14304 (N_14304,N_14224,N_14183);
nand U14305 (N_14305,N_14047,N_14042);
xor U14306 (N_14306,N_14058,N_14200);
and U14307 (N_14307,N_14131,N_14014);
nand U14308 (N_14308,N_14113,N_14218);
nand U14309 (N_14309,N_14073,N_14210);
nand U14310 (N_14310,N_14046,N_14012);
xor U14311 (N_14311,N_14185,N_14179);
nor U14312 (N_14312,N_14097,N_14089);
and U14313 (N_14313,N_14188,N_14079);
xor U14314 (N_14314,N_14150,N_14240);
nand U14315 (N_14315,N_14086,N_14248);
or U14316 (N_14316,N_14011,N_14242);
nor U14317 (N_14317,N_14241,N_14057);
or U14318 (N_14318,N_14038,N_14217);
nand U14319 (N_14319,N_14050,N_14159);
and U14320 (N_14320,N_14249,N_14063);
or U14321 (N_14321,N_14195,N_14236);
nand U14322 (N_14322,N_14124,N_14021);
xnor U14323 (N_14323,N_14133,N_14045);
and U14324 (N_14324,N_14100,N_14090);
xnor U14325 (N_14325,N_14096,N_14083);
nand U14326 (N_14326,N_14239,N_14165);
nand U14327 (N_14327,N_14212,N_14025);
xnor U14328 (N_14328,N_14121,N_14215);
xor U14329 (N_14329,N_14024,N_14075);
xnor U14330 (N_14330,N_14081,N_14222);
nor U14331 (N_14331,N_14134,N_14049);
and U14332 (N_14332,N_14040,N_14033);
nand U14333 (N_14333,N_14143,N_14109);
and U14334 (N_14334,N_14167,N_14141);
nor U14335 (N_14335,N_14213,N_14108);
xor U14336 (N_14336,N_14104,N_14018);
nor U14337 (N_14337,N_14123,N_14064);
or U14338 (N_14338,N_14247,N_14181);
or U14339 (N_14339,N_14170,N_14227);
xor U14340 (N_14340,N_14156,N_14074);
nand U14341 (N_14341,N_14082,N_14189);
and U14342 (N_14342,N_14023,N_14001);
nand U14343 (N_14343,N_14007,N_14015);
nand U14344 (N_14344,N_14142,N_14000);
xnor U14345 (N_14345,N_14085,N_14066);
and U14346 (N_14346,N_14068,N_14245);
nor U14347 (N_14347,N_14192,N_14186);
nand U14348 (N_14348,N_14219,N_14084);
nor U14349 (N_14349,N_14076,N_14205);
xnor U14350 (N_14350,N_14157,N_14174);
nand U14351 (N_14351,N_14044,N_14184);
nand U14352 (N_14352,N_14203,N_14237);
nor U14353 (N_14353,N_14032,N_14103);
nand U14354 (N_14354,N_14087,N_14138);
and U14355 (N_14355,N_14008,N_14177);
xor U14356 (N_14356,N_14153,N_14207);
nor U14357 (N_14357,N_14056,N_14101);
or U14358 (N_14358,N_14136,N_14191);
or U14359 (N_14359,N_14004,N_14053);
nand U14360 (N_14360,N_14034,N_14110);
nand U14361 (N_14361,N_14013,N_14201);
nor U14362 (N_14362,N_14016,N_14061);
and U14363 (N_14363,N_14022,N_14019);
nor U14364 (N_14364,N_14216,N_14223);
xnor U14365 (N_14365,N_14198,N_14009);
nand U14366 (N_14366,N_14169,N_14176);
xor U14367 (N_14367,N_14093,N_14051);
xnor U14368 (N_14368,N_14209,N_14048);
nor U14369 (N_14369,N_14039,N_14178);
and U14370 (N_14370,N_14029,N_14120);
nor U14371 (N_14371,N_14246,N_14118);
nor U14372 (N_14372,N_14043,N_14226);
nor U14373 (N_14373,N_14088,N_14182);
and U14374 (N_14374,N_14126,N_14197);
nor U14375 (N_14375,N_14046,N_14155);
nand U14376 (N_14376,N_14159,N_14057);
nor U14377 (N_14377,N_14179,N_14121);
or U14378 (N_14378,N_14125,N_14126);
xor U14379 (N_14379,N_14183,N_14221);
xor U14380 (N_14380,N_14050,N_14044);
xor U14381 (N_14381,N_14048,N_14024);
xnor U14382 (N_14382,N_14034,N_14184);
nand U14383 (N_14383,N_14085,N_14056);
nand U14384 (N_14384,N_14125,N_14173);
or U14385 (N_14385,N_14101,N_14032);
nand U14386 (N_14386,N_14047,N_14249);
and U14387 (N_14387,N_14115,N_14054);
nor U14388 (N_14388,N_14034,N_14005);
and U14389 (N_14389,N_14046,N_14222);
xor U14390 (N_14390,N_14181,N_14219);
xor U14391 (N_14391,N_14158,N_14126);
nor U14392 (N_14392,N_14068,N_14088);
nand U14393 (N_14393,N_14124,N_14241);
nor U14394 (N_14394,N_14190,N_14049);
and U14395 (N_14395,N_14163,N_14241);
and U14396 (N_14396,N_14102,N_14123);
xnor U14397 (N_14397,N_14028,N_14242);
and U14398 (N_14398,N_14175,N_14145);
and U14399 (N_14399,N_14117,N_14110);
xor U14400 (N_14400,N_14222,N_14079);
or U14401 (N_14401,N_14051,N_14075);
and U14402 (N_14402,N_14021,N_14029);
or U14403 (N_14403,N_14246,N_14050);
nor U14404 (N_14404,N_14221,N_14214);
and U14405 (N_14405,N_14095,N_14208);
and U14406 (N_14406,N_14166,N_14218);
nor U14407 (N_14407,N_14038,N_14077);
xnor U14408 (N_14408,N_14013,N_14134);
or U14409 (N_14409,N_14092,N_14033);
and U14410 (N_14410,N_14054,N_14157);
nor U14411 (N_14411,N_14119,N_14122);
or U14412 (N_14412,N_14037,N_14171);
xnor U14413 (N_14413,N_14080,N_14225);
nand U14414 (N_14414,N_14067,N_14152);
nand U14415 (N_14415,N_14132,N_14051);
nand U14416 (N_14416,N_14212,N_14245);
nor U14417 (N_14417,N_14135,N_14048);
nor U14418 (N_14418,N_14127,N_14192);
or U14419 (N_14419,N_14237,N_14157);
or U14420 (N_14420,N_14011,N_14176);
xnor U14421 (N_14421,N_14218,N_14212);
nor U14422 (N_14422,N_14166,N_14244);
xor U14423 (N_14423,N_14025,N_14007);
and U14424 (N_14424,N_14082,N_14047);
nand U14425 (N_14425,N_14225,N_14142);
xnor U14426 (N_14426,N_14000,N_14138);
nor U14427 (N_14427,N_14095,N_14188);
nand U14428 (N_14428,N_14113,N_14109);
xor U14429 (N_14429,N_14164,N_14014);
and U14430 (N_14430,N_14046,N_14028);
or U14431 (N_14431,N_14139,N_14079);
or U14432 (N_14432,N_14233,N_14110);
nor U14433 (N_14433,N_14150,N_14164);
nor U14434 (N_14434,N_14198,N_14039);
xor U14435 (N_14435,N_14011,N_14102);
nand U14436 (N_14436,N_14085,N_14213);
or U14437 (N_14437,N_14069,N_14143);
xor U14438 (N_14438,N_14001,N_14203);
xor U14439 (N_14439,N_14032,N_14094);
xor U14440 (N_14440,N_14095,N_14245);
or U14441 (N_14441,N_14166,N_14228);
nand U14442 (N_14442,N_14066,N_14065);
nor U14443 (N_14443,N_14176,N_14122);
nor U14444 (N_14444,N_14184,N_14130);
xor U14445 (N_14445,N_14186,N_14002);
nor U14446 (N_14446,N_14132,N_14054);
nor U14447 (N_14447,N_14185,N_14171);
and U14448 (N_14448,N_14022,N_14142);
and U14449 (N_14449,N_14078,N_14226);
and U14450 (N_14450,N_14012,N_14133);
nor U14451 (N_14451,N_14172,N_14077);
nand U14452 (N_14452,N_14206,N_14000);
nand U14453 (N_14453,N_14198,N_14048);
xor U14454 (N_14454,N_14148,N_14211);
xnor U14455 (N_14455,N_14092,N_14126);
nor U14456 (N_14456,N_14021,N_14046);
xnor U14457 (N_14457,N_14180,N_14030);
nand U14458 (N_14458,N_14198,N_14104);
nor U14459 (N_14459,N_14165,N_14039);
and U14460 (N_14460,N_14043,N_14206);
nand U14461 (N_14461,N_14147,N_14178);
or U14462 (N_14462,N_14104,N_14138);
and U14463 (N_14463,N_14072,N_14203);
xnor U14464 (N_14464,N_14221,N_14023);
nand U14465 (N_14465,N_14178,N_14015);
or U14466 (N_14466,N_14098,N_14011);
or U14467 (N_14467,N_14000,N_14018);
or U14468 (N_14468,N_14004,N_14118);
nor U14469 (N_14469,N_14137,N_14017);
xor U14470 (N_14470,N_14150,N_14158);
and U14471 (N_14471,N_14128,N_14222);
or U14472 (N_14472,N_14231,N_14172);
or U14473 (N_14473,N_14053,N_14040);
nand U14474 (N_14474,N_14026,N_14192);
and U14475 (N_14475,N_14041,N_14117);
xnor U14476 (N_14476,N_14245,N_14173);
and U14477 (N_14477,N_14220,N_14105);
xnor U14478 (N_14478,N_14158,N_14154);
nand U14479 (N_14479,N_14230,N_14118);
nand U14480 (N_14480,N_14022,N_14144);
nand U14481 (N_14481,N_14188,N_14125);
nor U14482 (N_14482,N_14241,N_14205);
nor U14483 (N_14483,N_14202,N_14199);
xor U14484 (N_14484,N_14170,N_14241);
and U14485 (N_14485,N_14004,N_14181);
nand U14486 (N_14486,N_14087,N_14219);
nor U14487 (N_14487,N_14053,N_14110);
xor U14488 (N_14488,N_14225,N_14222);
xor U14489 (N_14489,N_14001,N_14173);
and U14490 (N_14490,N_14047,N_14100);
nand U14491 (N_14491,N_14063,N_14170);
or U14492 (N_14492,N_14195,N_14049);
nor U14493 (N_14493,N_14168,N_14038);
or U14494 (N_14494,N_14055,N_14023);
or U14495 (N_14495,N_14243,N_14023);
or U14496 (N_14496,N_14248,N_14113);
or U14497 (N_14497,N_14241,N_14190);
xnor U14498 (N_14498,N_14050,N_14055);
nand U14499 (N_14499,N_14165,N_14093);
xor U14500 (N_14500,N_14437,N_14469);
and U14501 (N_14501,N_14253,N_14497);
nand U14502 (N_14502,N_14498,N_14301);
nor U14503 (N_14503,N_14269,N_14405);
and U14504 (N_14504,N_14390,N_14463);
or U14505 (N_14505,N_14316,N_14255);
and U14506 (N_14506,N_14388,N_14318);
and U14507 (N_14507,N_14371,N_14491);
and U14508 (N_14508,N_14477,N_14314);
or U14509 (N_14509,N_14328,N_14288);
xor U14510 (N_14510,N_14449,N_14471);
xnor U14511 (N_14511,N_14387,N_14458);
nand U14512 (N_14512,N_14347,N_14321);
xor U14513 (N_14513,N_14459,N_14258);
and U14514 (N_14514,N_14310,N_14369);
nor U14515 (N_14515,N_14373,N_14335);
or U14516 (N_14516,N_14480,N_14453);
or U14517 (N_14517,N_14394,N_14260);
nor U14518 (N_14518,N_14429,N_14364);
and U14519 (N_14519,N_14476,N_14393);
nand U14520 (N_14520,N_14489,N_14250);
nor U14521 (N_14521,N_14434,N_14262);
xnor U14522 (N_14522,N_14326,N_14462);
nor U14523 (N_14523,N_14486,N_14276);
or U14524 (N_14524,N_14415,N_14270);
xnor U14525 (N_14525,N_14365,N_14465);
xor U14526 (N_14526,N_14304,N_14281);
nand U14527 (N_14527,N_14431,N_14425);
nand U14528 (N_14528,N_14495,N_14340);
xnor U14529 (N_14529,N_14263,N_14291);
and U14530 (N_14530,N_14423,N_14299);
or U14531 (N_14531,N_14422,N_14282);
or U14532 (N_14532,N_14385,N_14322);
nand U14533 (N_14533,N_14327,N_14363);
and U14534 (N_14534,N_14349,N_14320);
nand U14535 (N_14535,N_14444,N_14417);
nor U14536 (N_14536,N_14350,N_14351);
nand U14537 (N_14537,N_14284,N_14311);
or U14538 (N_14538,N_14474,N_14278);
xnor U14539 (N_14539,N_14428,N_14353);
or U14540 (N_14540,N_14323,N_14479);
xor U14541 (N_14541,N_14460,N_14435);
or U14542 (N_14542,N_14357,N_14448);
and U14543 (N_14543,N_14294,N_14443);
nand U14544 (N_14544,N_14419,N_14391);
or U14545 (N_14545,N_14345,N_14483);
xor U14546 (N_14546,N_14467,N_14493);
or U14547 (N_14547,N_14332,N_14398);
nor U14548 (N_14548,N_14403,N_14378);
nor U14549 (N_14549,N_14468,N_14348);
nand U14550 (N_14550,N_14426,N_14482);
xnor U14551 (N_14551,N_14374,N_14300);
or U14552 (N_14552,N_14439,N_14334);
or U14553 (N_14553,N_14370,N_14265);
nor U14554 (N_14554,N_14317,N_14380);
and U14555 (N_14555,N_14379,N_14271);
nand U14556 (N_14556,N_14275,N_14416);
or U14557 (N_14557,N_14445,N_14251);
nor U14558 (N_14558,N_14470,N_14306);
nand U14559 (N_14559,N_14257,N_14484);
nor U14560 (N_14560,N_14293,N_14466);
and U14561 (N_14561,N_14381,N_14494);
nor U14562 (N_14562,N_14341,N_14324);
nand U14563 (N_14563,N_14396,N_14404);
xor U14564 (N_14564,N_14481,N_14277);
or U14565 (N_14565,N_14325,N_14384);
nor U14566 (N_14566,N_14464,N_14264);
nand U14567 (N_14567,N_14475,N_14267);
nor U14568 (N_14568,N_14287,N_14478);
and U14569 (N_14569,N_14329,N_14360);
nor U14570 (N_14570,N_14289,N_14452);
xor U14571 (N_14571,N_14490,N_14272);
and U14572 (N_14572,N_14400,N_14331);
xnor U14573 (N_14573,N_14410,N_14280);
xnor U14574 (N_14574,N_14342,N_14254);
nor U14575 (N_14575,N_14411,N_14307);
or U14576 (N_14576,N_14420,N_14496);
xor U14577 (N_14577,N_14424,N_14485);
nor U14578 (N_14578,N_14408,N_14285);
nand U14579 (N_14579,N_14436,N_14389);
or U14580 (N_14580,N_14338,N_14418);
or U14581 (N_14581,N_14312,N_14358);
nor U14582 (N_14582,N_14414,N_14252);
xnor U14583 (N_14583,N_14412,N_14386);
and U14584 (N_14584,N_14382,N_14315);
or U14585 (N_14585,N_14366,N_14383);
and U14586 (N_14586,N_14456,N_14308);
nor U14587 (N_14587,N_14455,N_14295);
nand U14588 (N_14588,N_14401,N_14397);
xnor U14589 (N_14589,N_14313,N_14451);
and U14590 (N_14590,N_14256,N_14377);
nor U14591 (N_14591,N_14261,N_14395);
or U14592 (N_14592,N_14268,N_14362);
xnor U14593 (N_14593,N_14336,N_14339);
nor U14594 (N_14594,N_14488,N_14427);
xnor U14595 (N_14595,N_14487,N_14359);
nand U14596 (N_14596,N_14392,N_14266);
or U14597 (N_14597,N_14450,N_14290);
or U14598 (N_14598,N_14457,N_14333);
nand U14599 (N_14599,N_14279,N_14283);
or U14600 (N_14600,N_14376,N_14472);
and U14601 (N_14601,N_14407,N_14343);
and U14602 (N_14602,N_14344,N_14302);
nand U14603 (N_14603,N_14402,N_14454);
nand U14604 (N_14604,N_14372,N_14368);
nor U14605 (N_14605,N_14356,N_14305);
or U14606 (N_14606,N_14319,N_14413);
nand U14607 (N_14607,N_14499,N_14375);
xor U14608 (N_14608,N_14421,N_14367);
nor U14609 (N_14609,N_14442,N_14286);
xnor U14610 (N_14610,N_14297,N_14352);
or U14611 (N_14611,N_14274,N_14303);
nor U14612 (N_14612,N_14473,N_14406);
or U14613 (N_14613,N_14461,N_14441);
or U14614 (N_14614,N_14409,N_14273);
and U14615 (N_14615,N_14440,N_14354);
or U14616 (N_14616,N_14298,N_14330);
nor U14617 (N_14617,N_14346,N_14433);
or U14618 (N_14618,N_14447,N_14337);
nor U14619 (N_14619,N_14355,N_14309);
xor U14620 (N_14620,N_14296,N_14432);
nand U14621 (N_14621,N_14438,N_14430);
nor U14622 (N_14622,N_14259,N_14446);
nand U14623 (N_14623,N_14361,N_14292);
or U14624 (N_14624,N_14492,N_14399);
nand U14625 (N_14625,N_14477,N_14256);
and U14626 (N_14626,N_14379,N_14474);
nor U14627 (N_14627,N_14312,N_14325);
nor U14628 (N_14628,N_14335,N_14405);
or U14629 (N_14629,N_14472,N_14343);
or U14630 (N_14630,N_14371,N_14362);
nor U14631 (N_14631,N_14392,N_14298);
xor U14632 (N_14632,N_14424,N_14456);
or U14633 (N_14633,N_14355,N_14482);
or U14634 (N_14634,N_14306,N_14331);
xor U14635 (N_14635,N_14464,N_14434);
nor U14636 (N_14636,N_14286,N_14296);
nand U14637 (N_14637,N_14257,N_14494);
and U14638 (N_14638,N_14345,N_14338);
and U14639 (N_14639,N_14357,N_14340);
nor U14640 (N_14640,N_14436,N_14446);
and U14641 (N_14641,N_14371,N_14287);
and U14642 (N_14642,N_14276,N_14385);
or U14643 (N_14643,N_14386,N_14489);
and U14644 (N_14644,N_14292,N_14291);
and U14645 (N_14645,N_14296,N_14320);
nand U14646 (N_14646,N_14399,N_14256);
xnor U14647 (N_14647,N_14396,N_14338);
nand U14648 (N_14648,N_14330,N_14272);
nand U14649 (N_14649,N_14367,N_14460);
nand U14650 (N_14650,N_14287,N_14452);
or U14651 (N_14651,N_14423,N_14375);
xnor U14652 (N_14652,N_14409,N_14454);
nand U14653 (N_14653,N_14427,N_14482);
or U14654 (N_14654,N_14370,N_14336);
and U14655 (N_14655,N_14437,N_14460);
nand U14656 (N_14656,N_14494,N_14302);
or U14657 (N_14657,N_14330,N_14388);
nand U14658 (N_14658,N_14316,N_14477);
or U14659 (N_14659,N_14358,N_14466);
nor U14660 (N_14660,N_14357,N_14281);
nand U14661 (N_14661,N_14408,N_14437);
or U14662 (N_14662,N_14264,N_14304);
nor U14663 (N_14663,N_14282,N_14376);
or U14664 (N_14664,N_14462,N_14320);
and U14665 (N_14665,N_14314,N_14319);
nor U14666 (N_14666,N_14330,N_14493);
nand U14667 (N_14667,N_14466,N_14334);
xnor U14668 (N_14668,N_14386,N_14314);
xor U14669 (N_14669,N_14461,N_14398);
xnor U14670 (N_14670,N_14325,N_14382);
nor U14671 (N_14671,N_14467,N_14354);
xor U14672 (N_14672,N_14416,N_14496);
and U14673 (N_14673,N_14448,N_14466);
nor U14674 (N_14674,N_14348,N_14420);
nand U14675 (N_14675,N_14341,N_14442);
nand U14676 (N_14676,N_14450,N_14405);
nor U14677 (N_14677,N_14405,N_14288);
and U14678 (N_14678,N_14456,N_14306);
or U14679 (N_14679,N_14318,N_14333);
xor U14680 (N_14680,N_14277,N_14403);
and U14681 (N_14681,N_14295,N_14405);
nand U14682 (N_14682,N_14270,N_14334);
xnor U14683 (N_14683,N_14263,N_14423);
or U14684 (N_14684,N_14397,N_14361);
nand U14685 (N_14685,N_14306,N_14485);
and U14686 (N_14686,N_14449,N_14400);
or U14687 (N_14687,N_14286,N_14448);
nand U14688 (N_14688,N_14293,N_14370);
nor U14689 (N_14689,N_14264,N_14267);
or U14690 (N_14690,N_14322,N_14497);
nand U14691 (N_14691,N_14360,N_14445);
and U14692 (N_14692,N_14400,N_14470);
or U14693 (N_14693,N_14427,N_14257);
nand U14694 (N_14694,N_14439,N_14283);
xor U14695 (N_14695,N_14289,N_14401);
nand U14696 (N_14696,N_14438,N_14402);
or U14697 (N_14697,N_14265,N_14467);
nand U14698 (N_14698,N_14337,N_14473);
or U14699 (N_14699,N_14300,N_14355);
xor U14700 (N_14700,N_14492,N_14385);
nand U14701 (N_14701,N_14403,N_14343);
nand U14702 (N_14702,N_14498,N_14291);
xnor U14703 (N_14703,N_14419,N_14353);
xnor U14704 (N_14704,N_14445,N_14472);
xnor U14705 (N_14705,N_14393,N_14354);
nor U14706 (N_14706,N_14496,N_14483);
nand U14707 (N_14707,N_14473,N_14296);
nand U14708 (N_14708,N_14277,N_14480);
nor U14709 (N_14709,N_14386,N_14301);
nor U14710 (N_14710,N_14424,N_14389);
xor U14711 (N_14711,N_14480,N_14410);
nand U14712 (N_14712,N_14453,N_14384);
or U14713 (N_14713,N_14432,N_14328);
xnor U14714 (N_14714,N_14279,N_14273);
nor U14715 (N_14715,N_14481,N_14437);
or U14716 (N_14716,N_14383,N_14317);
and U14717 (N_14717,N_14298,N_14426);
nand U14718 (N_14718,N_14374,N_14306);
xnor U14719 (N_14719,N_14389,N_14490);
nand U14720 (N_14720,N_14271,N_14397);
or U14721 (N_14721,N_14340,N_14435);
or U14722 (N_14722,N_14284,N_14362);
and U14723 (N_14723,N_14401,N_14308);
and U14724 (N_14724,N_14489,N_14283);
xnor U14725 (N_14725,N_14371,N_14338);
nand U14726 (N_14726,N_14311,N_14382);
or U14727 (N_14727,N_14323,N_14494);
xor U14728 (N_14728,N_14362,N_14311);
and U14729 (N_14729,N_14490,N_14378);
and U14730 (N_14730,N_14435,N_14384);
or U14731 (N_14731,N_14315,N_14397);
and U14732 (N_14732,N_14460,N_14296);
nor U14733 (N_14733,N_14496,N_14466);
nor U14734 (N_14734,N_14444,N_14433);
nor U14735 (N_14735,N_14400,N_14316);
or U14736 (N_14736,N_14277,N_14484);
xnor U14737 (N_14737,N_14315,N_14258);
nand U14738 (N_14738,N_14456,N_14392);
or U14739 (N_14739,N_14280,N_14341);
and U14740 (N_14740,N_14444,N_14413);
or U14741 (N_14741,N_14450,N_14348);
and U14742 (N_14742,N_14337,N_14292);
nor U14743 (N_14743,N_14253,N_14278);
xnor U14744 (N_14744,N_14467,N_14433);
or U14745 (N_14745,N_14337,N_14396);
or U14746 (N_14746,N_14256,N_14360);
or U14747 (N_14747,N_14297,N_14423);
and U14748 (N_14748,N_14346,N_14439);
nor U14749 (N_14749,N_14488,N_14444);
nor U14750 (N_14750,N_14555,N_14578);
or U14751 (N_14751,N_14592,N_14542);
and U14752 (N_14752,N_14516,N_14728);
nor U14753 (N_14753,N_14504,N_14727);
or U14754 (N_14754,N_14673,N_14573);
and U14755 (N_14755,N_14609,N_14572);
nor U14756 (N_14756,N_14713,N_14567);
xnor U14757 (N_14757,N_14629,N_14621);
and U14758 (N_14758,N_14503,N_14682);
xnor U14759 (N_14759,N_14588,N_14672);
nor U14760 (N_14760,N_14571,N_14749);
nand U14761 (N_14761,N_14723,N_14512);
xor U14762 (N_14762,N_14530,N_14557);
or U14763 (N_14763,N_14584,N_14586);
or U14764 (N_14764,N_14513,N_14604);
or U14765 (N_14765,N_14535,N_14714);
or U14766 (N_14766,N_14694,N_14501);
or U14767 (N_14767,N_14618,N_14687);
nand U14768 (N_14768,N_14511,N_14660);
nand U14769 (N_14769,N_14551,N_14640);
and U14770 (N_14770,N_14547,N_14539);
or U14771 (N_14771,N_14734,N_14684);
or U14772 (N_14772,N_14722,N_14689);
or U14773 (N_14773,N_14680,N_14560);
and U14774 (N_14774,N_14667,N_14664);
or U14775 (N_14775,N_14634,N_14706);
nor U14776 (N_14776,N_14681,N_14608);
and U14777 (N_14777,N_14517,N_14577);
nor U14778 (N_14778,N_14653,N_14668);
nor U14779 (N_14779,N_14692,N_14576);
and U14780 (N_14780,N_14614,N_14651);
and U14781 (N_14781,N_14597,N_14671);
xor U14782 (N_14782,N_14690,N_14704);
xor U14783 (N_14783,N_14659,N_14748);
and U14784 (N_14784,N_14502,N_14627);
or U14785 (N_14785,N_14566,N_14615);
nor U14786 (N_14786,N_14505,N_14719);
nand U14787 (N_14787,N_14601,N_14738);
nand U14788 (N_14788,N_14685,N_14626);
and U14789 (N_14789,N_14725,N_14670);
xnor U14790 (N_14790,N_14645,N_14563);
xor U14791 (N_14791,N_14549,N_14648);
or U14792 (N_14792,N_14695,N_14736);
xnor U14793 (N_14793,N_14533,N_14708);
nor U14794 (N_14794,N_14663,N_14662);
or U14795 (N_14795,N_14699,N_14523);
xnor U14796 (N_14796,N_14590,N_14657);
and U14797 (N_14797,N_14729,N_14558);
or U14798 (N_14798,N_14531,N_14637);
nand U14799 (N_14799,N_14631,N_14639);
and U14800 (N_14800,N_14677,N_14652);
xor U14801 (N_14801,N_14532,N_14745);
nor U14802 (N_14802,N_14617,N_14600);
nand U14803 (N_14803,N_14747,N_14596);
nor U14804 (N_14804,N_14715,N_14550);
or U14805 (N_14805,N_14683,N_14678);
and U14806 (N_14806,N_14553,N_14595);
or U14807 (N_14807,N_14654,N_14698);
nor U14808 (N_14808,N_14515,N_14666);
xnor U14809 (N_14809,N_14733,N_14693);
nor U14810 (N_14810,N_14613,N_14633);
xor U14811 (N_14811,N_14579,N_14741);
and U14812 (N_14812,N_14552,N_14538);
nand U14813 (N_14813,N_14575,N_14674);
xnor U14814 (N_14814,N_14743,N_14730);
xnor U14815 (N_14815,N_14508,N_14564);
xnor U14816 (N_14816,N_14679,N_14691);
nor U14817 (N_14817,N_14703,N_14655);
and U14818 (N_14818,N_14589,N_14688);
xor U14819 (N_14819,N_14528,N_14628);
nor U14820 (N_14820,N_14610,N_14712);
nand U14821 (N_14821,N_14746,N_14620);
xnor U14822 (N_14822,N_14509,N_14506);
or U14823 (N_14823,N_14650,N_14570);
xnor U14824 (N_14824,N_14602,N_14642);
and U14825 (N_14825,N_14581,N_14603);
nor U14826 (N_14826,N_14636,N_14519);
or U14827 (N_14827,N_14546,N_14540);
or U14828 (N_14828,N_14669,N_14565);
or U14829 (N_14829,N_14643,N_14739);
or U14830 (N_14830,N_14559,N_14641);
nor U14831 (N_14831,N_14740,N_14510);
nor U14832 (N_14832,N_14527,N_14574);
nor U14833 (N_14833,N_14534,N_14526);
or U14834 (N_14834,N_14721,N_14720);
or U14835 (N_14835,N_14541,N_14735);
nand U14836 (N_14836,N_14521,N_14624);
or U14837 (N_14837,N_14545,N_14561);
xnor U14838 (N_14838,N_14710,N_14543);
and U14839 (N_14839,N_14500,N_14724);
and U14840 (N_14840,N_14726,N_14705);
xor U14841 (N_14841,N_14709,N_14537);
or U14842 (N_14842,N_14644,N_14718);
nand U14843 (N_14843,N_14732,N_14562);
and U14844 (N_14844,N_14568,N_14591);
xnor U14845 (N_14845,N_14611,N_14737);
xnor U14846 (N_14846,N_14522,N_14606);
and U14847 (N_14847,N_14594,N_14585);
nor U14848 (N_14848,N_14625,N_14507);
nand U14849 (N_14849,N_14605,N_14707);
nand U14850 (N_14850,N_14587,N_14514);
nor U14851 (N_14851,N_14696,N_14665);
nor U14852 (N_14852,N_14520,N_14716);
nor U14853 (N_14853,N_14607,N_14548);
or U14854 (N_14854,N_14697,N_14518);
or U14855 (N_14855,N_14638,N_14676);
and U14856 (N_14856,N_14661,N_14711);
or U14857 (N_14857,N_14529,N_14612);
nor U14858 (N_14858,N_14646,N_14525);
and U14859 (N_14859,N_14742,N_14675);
nor U14860 (N_14860,N_14658,N_14554);
xor U14861 (N_14861,N_14619,N_14524);
nor U14862 (N_14862,N_14536,N_14582);
and U14863 (N_14863,N_14701,N_14744);
and U14864 (N_14864,N_14686,N_14700);
nand U14865 (N_14865,N_14635,N_14616);
xor U14866 (N_14866,N_14569,N_14656);
nand U14867 (N_14867,N_14702,N_14731);
xnor U14868 (N_14868,N_14717,N_14630);
nor U14869 (N_14869,N_14598,N_14583);
or U14870 (N_14870,N_14599,N_14593);
nand U14871 (N_14871,N_14649,N_14622);
or U14872 (N_14872,N_14647,N_14544);
nand U14873 (N_14873,N_14556,N_14632);
xnor U14874 (N_14874,N_14623,N_14580);
xnor U14875 (N_14875,N_14656,N_14578);
or U14876 (N_14876,N_14510,N_14506);
xnor U14877 (N_14877,N_14729,N_14687);
and U14878 (N_14878,N_14622,N_14512);
xnor U14879 (N_14879,N_14571,N_14527);
nor U14880 (N_14880,N_14523,N_14675);
and U14881 (N_14881,N_14706,N_14667);
nand U14882 (N_14882,N_14584,N_14574);
nor U14883 (N_14883,N_14559,N_14744);
and U14884 (N_14884,N_14726,N_14656);
nand U14885 (N_14885,N_14743,N_14610);
xor U14886 (N_14886,N_14633,N_14734);
xnor U14887 (N_14887,N_14514,N_14532);
xnor U14888 (N_14888,N_14617,N_14643);
nand U14889 (N_14889,N_14621,N_14502);
nor U14890 (N_14890,N_14667,N_14552);
or U14891 (N_14891,N_14552,N_14558);
nand U14892 (N_14892,N_14662,N_14542);
xor U14893 (N_14893,N_14537,N_14604);
nor U14894 (N_14894,N_14579,N_14744);
nand U14895 (N_14895,N_14747,N_14608);
xnor U14896 (N_14896,N_14600,N_14737);
and U14897 (N_14897,N_14611,N_14585);
nor U14898 (N_14898,N_14672,N_14595);
xnor U14899 (N_14899,N_14548,N_14554);
and U14900 (N_14900,N_14555,N_14536);
xor U14901 (N_14901,N_14576,N_14663);
xnor U14902 (N_14902,N_14710,N_14738);
nor U14903 (N_14903,N_14698,N_14733);
nor U14904 (N_14904,N_14682,N_14667);
and U14905 (N_14905,N_14629,N_14535);
nand U14906 (N_14906,N_14589,N_14539);
or U14907 (N_14907,N_14721,N_14516);
nand U14908 (N_14908,N_14541,N_14660);
and U14909 (N_14909,N_14662,N_14681);
nand U14910 (N_14910,N_14726,N_14635);
and U14911 (N_14911,N_14586,N_14560);
nor U14912 (N_14912,N_14707,N_14726);
xor U14913 (N_14913,N_14575,N_14580);
xor U14914 (N_14914,N_14651,N_14661);
and U14915 (N_14915,N_14675,N_14541);
nand U14916 (N_14916,N_14612,N_14715);
and U14917 (N_14917,N_14512,N_14655);
and U14918 (N_14918,N_14649,N_14697);
or U14919 (N_14919,N_14512,N_14600);
nand U14920 (N_14920,N_14501,N_14606);
and U14921 (N_14921,N_14707,N_14599);
nand U14922 (N_14922,N_14508,N_14509);
nand U14923 (N_14923,N_14684,N_14699);
and U14924 (N_14924,N_14585,N_14661);
nand U14925 (N_14925,N_14575,N_14641);
and U14926 (N_14926,N_14552,N_14733);
and U14927 (N_14927,N_14587,N_14547);
nand U14928 (N_14928,N_14531,N_14570);
or U14929 (N_14929,N_14733,N_14539);
or U14930 (N_14930,N_14632,N_14749);
nand U14931 (N_14931,N_14645,N_14602);
and U14932 (N_14932,N_14731,N_14568);
nand U14933 (N_14933,N_14676,N_14717);
or U14934 (N_14934,N_14599,N_14552);
nand U14935 (N_14935,N_14604,N_14607);
nand U14936 (N_14936,N_14578,N_14544);
nand U14937 (N_14937,N_14652,N_14573);
and U14938 (N_14938,N_14508,N_14684);
nand U14939 (N_14939,N_14747,N_14743);
nand U14940 (N_14940,N_14557,N_14743);
xor U14941 (N_14941,N_14744,N_14594);
nor U14942 (N_14942,N_14747,N_14526);
nor U14943 (N_14943,N_14710,N_14745);
and U14944 (N_14944,N_14536,N_14714);
xnor U14945 (N_14945,N_14747,N_14563);
nand U14946 (N_14946,N_14549,N_14628);
or U14947 (N_14947,N_14740,N_14592);
nand U14948 (N_14948,N_14590,N_14705);
nor U14949 (N_14949,N_14587,N_14646);
and U14950 (N_14950,N_14640,N_14509);
nor U14951 (N_14951,N_14683,N_14747);
or U14952 (N_14952,N_14503,N_14660);
and U14953 (N_14953,N_14689,N_14694);
xor U14954 (N_14954,N_14506,N_14738);
nor U14955 (N_14955,N_14558,N_14699);
nand U14956 (N_14956,N_14578,N_14708);
or U14957 (N_14957,N_14515,N_14614);
nand U14958 (N_14958,N_14671,N_14507);
xnor U14959 (N_14959,N_14741,N_14504);
nor U14960 (N_14960,N_14527,N_14655);
and U14961 (N_14961,N_14652,N_14508);
xor U14962 (N_14962,N_14629,N_14717);
xnor U14963 (N_14963,N_14651,N_14658);
or U14964 (N_14964,N_14734,N_14685);
and U14965 (N_14965,N_14623,N_14507);
xnor U14966 (N_14966,N_14683,N_14595);
nor U14967 (N_14967,N_14560,N_14584);
nand U14968 (N_14968,N_14640,N_14501);
nor U14969 (N_14969,N_14578,N_14688);
or U14970 (N_14970,N_14730,N_14672);
nor U14971 (N_14971,N_14605,N_14625);
and U14972 (N_14972,N_14555,N_14695);
xor U14973 (N_14973,N_14514,N_14598);
and U14974 (N_14974,N_14634,N_14677);
xor U14975 (N_14975,N_14514,N_14636);
and U14976 (N_14976,N_14608,N_14549);
or U14977 (N_14977,N_14501,N_14713);
nand U14978 (N_14978,N_14694,N_14541);
and U14979 (N_14979,N_14608,N_14589);
xnor U14980 (N_14980,N_14678,N_14500);
or U14981 (N_14981,N_14741,N_14744);
and U14982 (N_14982,N_14561,N_14701);
nor U14983 (N_14983,N_14640,N_14645);
nand U14984 (N_14984,N_14534,N_14662);
nor U14985 (N_14985,N_14730,N_14506);
nand U14986 (N_14986,N_14536,N_14745);
or U14987 (N_14987,N_14516,N_14537);
nand U14988 (N_14988,N_14746,N_14735);
and U14989 (N_14989,N_14706,N_14635);
nor U14990 (N_14990,N_14539,N_14629);
nand U14991 (N_14991,N_14696,N_14635);
and U14992 (N_14992,N_14660,N_14602);
nor U14993 (N_14993,N_14690,N_14603);
nand U14994 (N_14994,N_14614,N_14691);
and U14995 (N_14995,N_14505,N_14571);
or U14996 (N_14996,N_14663,N_14680);
and U14997 (N_14997,N_14645,N_14619);
xnor U14998 (N_14998,N_14709,N_14561);
and U14999 (N_14999,N_14558,N_14531);
or U15000 (N_15000,N_14940,N_14857);
and U15001 (N_15001,N_14859,N_14822);
and U15002 (N_15002,N_14867,N_14829);
nand U15003 (N_15003,N_14891,N_14938);
or U15004 (N_15004,N_14875,N_14912);
nor U15005 (N_15005,N_14848,N_14953);
and U15006 (N_15006,N_14942,N_14936);
xnor U15007 (N_15007,N_14853,N_14753);
nand U15008 (N_15008,N_14947,N_14902);
nand U15009 (N_15009,N_14966,N_14894);
xnor U15010 (N_15010,N_14901,N_14830);
nor U15011 (N_15011,N_14866,N_14849);
or U15012 (N_15012,N_14910,N_14771);
or U15013 (N_15013,N_14917,N_14943);
nor U15014 (N_15014,N_14808,N_14871);
nand U15015 (N_15015,N_14925,N_14772);
nor U15016 (N_15016,N_14990,N_14759);
nor U15017 (N_15017,N_14958,N_14838);
xor U15018 (N_15018,N_14956,N_14979);
nor U15019 (N_15019,N_14995,N_14915);
nor U15020 (N_15020,N_14881,N_14946);
or U15021 (N_15021,N_14898,N_14879);
xnor U15022 (N_15022,N_14914,N_14831);
nor U15023 (N_15023,N_14991,N_14810);
or U15024 (N_15024,N_14981,N_14975);
and U15025 (N_15025,N_14844,N_14922);
nand U15026 (N_15026,N_14951,N_14937);
and U15027 (N_15027,N_14983,N_14763);
nor U15028 (N_15028,N_14978,N_14919);
and U15029 (N_15029,N_14842,N_14862);
xor U15030 (N_15030,N_14781,N_14839);
nand U15031 (N_15031,N_14920,N_14778);
and U15032 (N_15032,N_14854,N_14820);
or U15033 (N_15033,N_14803,N_14788);
xnor U15034 (N_15034,N_14861,N_14836);
nor U15035 (N_15035,N_14976,N_14782);
and U15036 (N_15036,N_14800,N_14784);
and U15037 (N_15037,N_14897,N_14965);
xnor U15038 (N_15038,N_14806,N_14904);
xor U15039 (N_15039,N_14931,N_14868);
xnor U15040 (N_15040,N_14935,N_14865);
nand U15041 (N_15041,N_14939,N_14837);
nand U15042 (N_15042,N_14864,N_14930);
nor U15043 (N_15043,N_14851,N_14863);
or U15044 (N_15044,N_14928,N_14877);
and U15045 (N_15045,N_14841,N_14885);
nand U15046 (N_15046,N_14852,N_14994);
and U15047 (N_15047,N_14923,N_14908);
xnor U15048 (N_15048,N_14815,N_14789);
nand U15049 (N_15049,N_14796,N_14809);
and U15050 (N_15050,N_14798,N_14819);
and U15051 (N_15051,N_14890,N_14766);
nor U15052 (N_15052,N_14969,N_14832);
xor U15053 (N_15053,N_14869,N_14764);
nand U15054 (N_15054,N_14821,N_14855);
nand U15055 (N_15055,N_14909,N_14964);
nor U15056 (N_15056,N_14840,N_14932);
xnor U15057 (N_15057,N_14785,N_14952);
or U15058 (N_15058,N_14760,N_14955);
nor U15059 (N_15059,N_14774,N_14751);
nor U15060 (N_15060,N_14845,N_14835);
and U15061 (N_15061,N_14959,N_14802);
and U15062 (N_15062,N_14828,N_14780);
nand U15063 (N_15063,N_14754,N_14783);
nor U15064 (N_15064,N_14860,N_14913);
nand U15065 (N_15065,N_14977,N_14755);
nand U15066 (N_15066,N_14999,N_14768);
and U15067 (N_15067,N_14758,N_14813);
nand U15068 (N_15068,N_14816,N_14756);
or U15069 (N_15069,N_14957,N_14906);
or U15070 (N_15070,N_14961,N_14945);
and U15071 (N_15071,N_14903,N_14907);
or U15072 (N_15072,N_14769,N_14792);
and U15073 (N_15073,N_14791,N_14992);
xor U15074 (N_15074,N_14807,N_14944);
or U15075 (N_15075,N_14765,N_14997);
nor U15076 (N_15076,N_14797,N_14874);
nor U15077 (N_15077,N_14776,N_14817);
xnor U15078 (N_15078,N_14982,N_14886);
nor U15079 (N_15079,N_14876,N_14972);
or U15080 (N_15080,N_14998,N_14762);
nor U15081 (N_15081,N_14980,N_14811);
xnor U15082 (N_15082,N_14916,N_14752);
and U15083 (N_15083,N_14927,N_14777);
nor U15084 (N_15084,N_14880,N_14775);
or U15085 (N_15085,N_14899,N_14962);
and U15086 (N_15086,N_14770,N_14787);
or U15087 (N_15087,N_14826,N_14889);
nor U15088 (N_15088,N_14818,N_14924);
xnor U15089 (N_15089,N_14850,N_14761);
nand U15090 (N_15090,N_14887,N_14793);
and U15091 (N_15091,N_14773,N_14827);
and U15092 (N_15092,N_14960,N_14896);
nand U15093 (N_15093,N_14888,N_14989);
xor U15094 (N_15094,N_14954,N_14921);
or U15095 (N_15095,N_14934,N_14790);
nand U15096 (N_15096,N_14950,N_14941);
xor U15097 (N_15097,N_14892,N_14825);
nor U15098 (N_15098,N_14987,N_14967);
nor U15099 (N_15099,N_14804,N_14929);
or U15100 (N_15100,N_14801,N_14973);
and U15101 (N_15101,N_14872,N_14949);
or U15102 (N_15102,N_14799,N_14750);
nand U15103 (N_15103,N_14843,N_14779);
nor U15104 (N_15104,N_14858,N_14882);
and U15105 (N_15105,N_14996,N_14905);
and U15106 (N_15106,N_14833,N_14878);
nand U15107 (N_15107,N_14963,N_14911);
and U15108 (N_15108,N_14846,N_14974);
xnor U15109 (N_15109,N_14971,N_14984);
xnor U15110 (N_15110,N_14895,N_14823);
and U15111 (N_15111,N_14786,N_14993);
nand U15112 (N_15112,N_14795,N_14767);
nor U15113 (N_15113,N_14933,N_14970);
nor U15114 (N_15114,N_14794,N_14900);
nand U15115 (N_15115,N_14926,N_14883);
xnor U15116 (N_15116,N_14948,N_14870);
nand U15117 (N_15117,N_14847,N_14834);
nor U15118 (N_15118,N_14873,N_14968);
and U15119 (N_15119,N_14812,N_14918);
and U15120 (N_15120,N_14985,N_14988);
or U15121 (N_15121,N_14893,N_14884);
nor U15122 (N_15122,N_14986,N_14824);
or U15123 (N_15123,N_14757,N_14814);
xor U15124 (N_15124,N_14856,N_14805);
xor U15125 (N_15125,N_14796,N_14862);
or U15126 (N_15126,N_14847,N_14770);
xnor U15127 (N_15127,N_14975,N_14841);
nand U15128 (N_15128,N_14930,N_14908);
nor U15129 (N_15129,N_14753,N_14857);
nand U15130 (N_15130,N_14832,N_14865);
or U15131 (N_15131,N_14951,N_14874);
nor U15132 (N_15132,N_14775,N_14827);
or U15133 (N_15133,N_14894,N_14823);
or U15134 (N_15134,N_14977,N_14817);
or U15135 (N_15135,N_14989,N_14907);
nand U15136 (N_15136,N_14805,N_14862);
and U15137 (N_15137,N_14980,N_14988);
nor U15138 (N_15138,N_14996,N_14852);
nand U15139 (N_15139,N_14874,N_14888);
nor U15140 (N_15140,N_14800,N_14928);
xor U15141 (N_15141,N_14819,N_14880);
nand U15142 (N_15142,N_14928,N_14756);
nor U15143 (N_15143,N_14851,N_14945);
nor U15144 (N_15144,N_14788,N_14837);
and U15145 (N_15145,N_14792,N_14875);
nand U15146 (N_15146,N_14954,N_14788);
or U15147 (N_15147,N_14842,N_14902);
and U15148 (N_15148,N_14764,N_14973);
nand U15149 (N_15149,N_14774,N_14898);
nor U15150 (N_15150,N_14784,N_14951);
nand U15151 (N_15151,N_14775,N_14879);
nor U15152 (N_15152,N_14995,N_14827);
nand U15153 (N_15153,N_14767,N_14922);
nor U15154 (N_15154,N_14998,N_14983);
nand U15155 (N_15155,N_14912,N_14792);
nor U15156 (N_15156,N_14815,N_14996);
xnor U15157 (N_15157,N_14882,N_14936);
nor U15158 (N_15158,N_14759,N_14806);
xor U15159 (N_15159,N_14899,N_14818);
or U15160 (N_15160,N_14945,N_14873);
nand U15161 (N_15161,N_14812,N_14884);
nand U15162 (N_15162,N_14795,N_14876);
xor U15163 (N_15163,N_14785,N_14775);
xor U15164 (N_15164,N_14777,N_14881);
and U15165 (N_15165,N_14785,N_14809);
or U15166 (N_15166,N_14950,N_14861);
nor U15167 (N_15167,N_14928,N_14875);
nand U15168 (N_15168,N_14985,N_14830);
and U15169 (N_15169,N_14934,N_14958);
or U15170 (N_15170,N_14989,N_14867);
and U15171 (N_15171,N_14865,N_14875);
nor U15172 (N_15172,N_14919,N_14984);
nand U15173 (N_15173,N_14795,N_14787);
and U15174 (N_15174,N_14790,N_14969);
nor U15175 (N_15175,N_14993,N_14988);
xnor U15176 (N_15176,N_14799,N_14881);
nand U15177 (N_15177,N_14907,N_14762);
xnor U15178 (N_15178,N_14880,N_14785);
nand U15179 (N_15179,N_14945,N_14902);
nor U15180 (N_15180,N_14771,N_14986);
and U15181 (N_15181,N_14800,N_14802);
nor U15182 (N_15182,N_14771,N_14935);
or U15183 (N_15183,N_14761,N_14775);
or U15184 (N_15184,N_14965,N_14899);
or U15185 (N_15185,N_14999,N_14896);
nand U15186 (N_15186,N_14918,N_14832);
xor U15187 (N_15187,N_14784,N_14990);
or U15188 (N_15188,N_14906,N_14965);
nor U15189 (N_15189,N_14967,N_14832);
xnor U15190 (N_15190,N_14753,N_14831);
and U15191 (N_15191,N_14975,N_14988);
nor U15192 (N_15192,N_14878,N_14909);
and U15193 (N_15193,N_14934,N_14788);
nor U15194 (N_15194,N_14903,N_14925);
xor U15195 (N_15195,N_14974,N_14822);
nor U15196 (N_15196,N_14801,N_14857);
nand U15197 (N_15197,N_14830,N_14898);
and U15198 (N_15198,N_14888,N_14791);
and U15199 (N_15199,N_14831,N_14830);
nand U15200 (N_15200,N_14784,N_14843);
nor U15201 (N_15201,N_14965,N_14818);
nand U15202 (N_15202,N_14882,N_14794);
and U15203 (N_15203,N_14834,N_14872);
or U15204 (N_15204,N_14830,N_14964);
xnor U15205 (N_15205,N_14942,N_14967);
nand U15206 (N_15206,N_14973,N_14996);
nand U15207 (N_15207,N_14785,N_14776);
and U15208 (N_15208,N_14845,N_14910);
nand U15209 (N_15209,N_14799,N_14991);
and U15210 (N_15210,N_14782,N_14859);
or U15211 (N_15211,N_14860,N_14937);
xnor U15212 (N_15212,N_14790,N_14919);
nor U15213 (N_15213,N_14787,N_14958);
nand U15214 (N_15214,N_14950,N_14891);
and U15215 (N_15215,N_14955,N_14966);
nor U15216 (N_15216,N_14989,N_14988);
xnor U15217 (N_15217,N_14930,N_14757);
and U15218 (N_15218,N_14752,N_14816);
nor U15219 (N_15219,N_14866,N_14846);
and U15220 (N_15220,N_14897,N_14762);
and U15221 (N_15221,N_14796,N_14761);
nor U15222 (N_15222,N_14965,N_14755);
and U15223 (N_15223,N_14925,N_14845);
xnor U15224 (N_15224,N_14916,N_14918);
and U15225 (N_15225,N_14811,N_14840);
nand U15226 (N_15226,N_14854,N_14838);
and U15227 (N_15227,N_14897,N_14920);
xnor U15228 (N_15228,N_14863,N_14886);
nand U15229 (N_15229,N_14998,N_14846);
nand U15230 (N_15230,N_14797,N_14925);
and U15231 (N_15231,N_14752,N_14784);
or U15232 (N_15232,N_14785,N_14959);
nand U15233 (N_15233,N_14777,N_14914);
xor U15234 (N_15234,N_14943,N_14783);
and U15235 (N_15235,N_14859,N_14951);
nor U15236 (N_15236,N_14968,N_14949);
nand U15237 (N_15237,N_14810,N_14917);
nand U15238 (N_15238,N_14998,N_14814);
xnor U15239 (N_15239,N_14999,N_14914);
xnor U15240 (N_15240,N_14893,N_14830);
and U15241 (N_15241,N_14997,N_14952);
xnor U15242 (N_15242,N_14951,N_14963);
xnor U15243 (N_15243,N_14765,N_14918);
and U15244 (N_15244,N_14958,N_14967);
nor U15245 (N_15245,N_14775,N_14808);
nor U15246 (N_15246,N_14761,N_14985);
and U15247 (N_15247,N_14846,N_14835);
nand U15248 (N_15248,N_14776,N_14790);
nand U15249 (N_15249,N_14985,N_14856);
and U15250 (N_15250,N_15199,N_15152);
or U15251 (N_15251,N_15114,N_15121);
nor U15252 (N_15252,N_15232,N_15053);
and U15253 (N_15253,N_15040,N_15016);
or U15254 (N_15254,N_15192,N_15158);
and U15255 (N_15255,N_15137,N_15205);
nand U15256 (N_15256,N_15212,N_15106);
nand U15257 (N_15257,N_15020,N_15044);
and U15258 (N_15258,N_15018,N_15248);
or U15259 (N_15259,N_15078,N_15000);
and U15260 (N_15260,N_15034,N_15170);
xnor U15261 (N_15261,N_15140,N_15014);
nor U15262 (N_15262,N_15227,N_15083);
nor U15263 (N_15263,N_15097,N_15071);
nand U15264 (N_15264,N_15146,N_15214);
nor U15265 (N_15265,N_15190,N_15105);
nor U15266 (N_15266,N_15150,N_15165);
nor U15267 (N_15267,N_15052,N_15160);
or U15268 (N_15268,N_15029,N_15135);
xor U15269 (N_15269,N_15045,N_15129);
nand U15270 (N_15270,N_15100,N_15118);
or U15271 (N_15271,N_15002,N_15225);
and U15272 (N_15272,N_15042,N_15008);
nor U15273 (N_15273,N_15245,N_15148);
or U15274 (N_15274,N_15130,N_15082);
xnor U15275 (N_15275,N_15172,N_15126);
nand U15276 (N_15276,N_15079,N_15171);
or U15277 (N_15277,N_15019,N_15133);
xor U15278 (N_15278,N_15055,N_15164);
nor U15279 (N_15279,N_15237,N_15182);
xor U15280 (N_15280,N_15151,N_15033);
nand U15281 (N_15281,N_15176,N_15023);
or U15282 (N_15282,N_15069,N_15175);
nor U15283 (N_15283,N_15244,N_15234);
nor U15284 (N_15284,N_15087,N_15235);
nand U15285 (N_15285,N_15063,N_15039);
or U15286 (N_15286,N_15025,N_15162);
and U15287 (N_15287,N_15228,N_15073);
and U15288 (N_15288,N_15021,N_15186);
or U15289 (N_15289,N_15099,N_15120);
and U15290 (N_15290,N_15085,N_15179);
nand U15291 (N_15291,N_15098,N_15153);
xor U15292 (N_15292,N_15065,N_15167);
or U15293 (N_15293,N_15015,N_15088);
and U15294 (N_15294,N_15115,N_15022);
xnor U15295 (N_15295,N_15229,N_15193);
nand U15296 (N_15296,N_15231,N_15183);
or U15297 (N_15297,N_15166,N_15138);
nor U15298 (N_15298,N_15038,N_15030);
and U15299 (N_15299,N_15059,N_15122);
nand U15300 (N_15300,N_15013,N_15060);
nand U15301 (N_15301,N_15050,N_15178);
nand U15302 (N_15302,N_15075,N_15216);
nor U15303 (N_15303,N_15057,N_15090);
or U15304 (N_15304,N_15037,N_15219);
and U15305 (N_15305,N_15224,N_15070);
nor U15306 (N_15306,N_15031,N_15111);
or U15307 (N_15307,N_15236,N_15058);
nand U15308 (N_15308,N_15210,N_15157);
nand U15309 (N_15309,N_15064,N_15154);
nor U15310 (N_15310,N_15139,N_15201);
and U15311 (N_15311,N_15102,N_15095);
or U15312 (N_15312,N_15046,N_15032);
or U15313 (N_15313,N_15094,N_15009);
nand U15314 (N_15314,N_15027,N_15001);
xnor U15315 (N_15315,N_15221,N_15180);
nor U15316 (N_15316,N_15084,N_15074);
nor U15317 (N_15317,N_15132,N_15024);
or U15318 (N_15318,N_15198,N_15127);
nand U15319 (N_15319,N_15003,N_15195);
nand U15320 (N_15320,N_15169,N_15143);
nand U15321 (N_15321,N_15086,N_15215);
and U15322 (N_15322,N_15041,N_15207);
and U15323 (N_15323,N_15246,N_15124);
nor U15324 (N_15324,N_15134,N_15247);
nand U15325 (N_15325,N_15197,N_15222);
nor U15326 (N_15326,N_15068,N_15131);
xnor U15327 (N_15327,N_15108,N_15107);
xnor U15328 (N_15328,N_15017,N_15076);
and U15329 (N_15329,N_15010,N_15213);
nand U15330 (N_15330,N_15238,N_15209);
nor U15331 (N_15331,N_15243,N_15174);
or U15332 (N_15332,N_15067,N_15123);
nor U15333 (N_15333,N_15220,N_15204);
or U15334 (N_15334,N_15110,N_15241);
nand U15335 (N_15335,N_15056,N_15049);
nand U15336 (N_15336,N_15149,N_15144);
xnor U15337 (N_15337,N_15233,N_15091);
and U15338 (N_15338,N_15217,N_15249);
nor U15339 (N_15339,N_15206,N_15047);
nand U15340 (N_15340,N_15177,N_15125);
and U15341 (N_15341,N_15109,N_15163);
nor U15342 (N_15342,N_15189,N_15136);
and U15343 (N_15343,N_15141,N_15203);
nor U15344 (N_15344,N_15240,N_15066);
and U15345 (N_15345,N_15155,N_15101);
or U15346 (N_15346,N_15043,N_15128);
and U15347 (N_15347,N_15242,N_15072);
nor U15348 (N_15348,N_15187,N_15226);
nor U15349 (N_15349,N_15185,N_15112);
or U15350 (N_15350,N_15051,N_15035);
nor U15351 (N_15351,N_15156,N_15184);
nor U15352 (N_15352,N_15080,N_15119);
xnor U15353 (N_15353,N_15061,N_15006);
or U15354 (N_15354,N_15092,N_15191);
xor U15355 (N_15355,N_15048,N_15096);
nand U15356 (N_15356,N_15007,N_15103);
nor U15357 (N_15357,N_15036,N_15054);
nor U15358 (N_15358,N_15011,N_15196);
and U15359 (N_15359,N_15028,N_15089);
and U15360 (N_15360,N_15113,N_15081);
and U15361 (N_15361,N_15093,N_15004);
and U15362 (N_15362,N_15026,N_15062);
nor U15363 (N_15363,N_15211,N_15218);
nand U15364 (N_15364,N_15077,N_15188);
or U15365 (N_15365,N_15147,N_15168);
xor U15366 (N_15366,N_15173,N_15194);
and U15367 (N_15367,N_15181,N_15159);
and U15368 (N_15368,N_15005,N_15142);
nand U15369 (N_15369,N_15145,N_15117);
and U15370 (N_15370,N_15104,N_15239);
nor U15371 (N_15371,N_15223,N_15202);
and U15372 (N_15372,N_15208,N_15012);
xnor U15373 (N_15373,N_15230,N_15200);
and U15374 (N_15374,N_15161,N_15116);
nand U15375 (N_15375,N_15122,N_15233);
nand U15376 (N_15376,N_15129,N_15004);
nand U15377 (N_15377,N_15054,N_15083);
xor U15378 (N_15378,N_15100,N_15219);
nor U15379 (N_15379,N_15119,N_15205);
nand U15380 (N_15380,N_15237,N_15162);
nand U15381 (N_15381,N_15070,N_15113);
or U15382 (N_15382,N_15001,N_15140);
nand U15383 (N_15383,N_15077,N_15160);
and U15384 (N_15384,N_15031,N_15223);
nor U15385 (N_15385,N_15171,N_15226);
xnor U15386 (N_15386,N_15235,N_15034);
nand U15387 (N_15387,N_15216,N_15135);
nor U15388 (N_15388,N_15249,N_15071);
or U15389 (N_15389,N_15047,N_15097);
nor U15390 (N_15390,N_15116,N_15155);
and U15391 (N_15391,N_15084,N_15243);
or U15392 (N_15392,N_15044,N_15218);
and U15393 (N_15393,N_15242,N_15123);
xnor U15394 (N_15394,N_15167,N_15133);
nand U15395 (N_15395,N_15122,N_15014);
and U15396 (N_15396,N_15092,N_15043);
nor U15397 (N_15397,N_15080,N_15148);
and U15398 (N_15398,N_15176,N_15147);
nor U15399 (N_15399,N_15020,N_15032);
xor U15400 (N_15400,N_15040,N_15091);
nand U15401 (N_15401,N_15023,N_15083);
and U15402 (N_15402,N_15153,N_15172);
or U15403 (N_15403,N_15015,N_15155);
and U15404 (N_15404,N_15003,N_15184);
or U15405 (N_15405,N_15210,N_15182);
nand U15406 (N_15406,N_15046,N_15067);
or U15407 (N_15407,N_15197,N_15070);
xnor U15408 (N_15408,N_15106,N_15002);
nand U15409 (N_15409,N_15159,N_15102);
nand U15410 (N_15410,N_15114,N_15130);
or U15411 (N_15411,N_15031,N_15109);
and U15412 (N_15412,N_15142,N_15220);
nand U15413 (N_15413,N_15122,N_15225);
nand U15414 (N_15414,N_15018,N_15079);
nand U15415 (N_15415,N_15056,N_15174);
and U15416 (N_15416,N_15075,N_15226);
xor U15417 (N_15417,N_15063,N_15203);
or U15418 (N_15418,N_15076,N_15000);
nor U15419 (N_15419,N_15223,N_15124);
or U15420 (N_15420,N_15137,N_15193);
xor U15421 (N_15421,N_15007,N_15234);
xor U15422 (N_15422,N_15178,N_15136);
and U15423 (N_15423,N_15166,N_15112);
or U15424 (N_15424,N_15057,N_15016);
or U15425 (N_15425,N_15049,N_15045);
nand U15426 (N_15426,N_15203,N_15220);
xor U15427 (N_15427,N_15206,N_15092);
or U15428 (N_15428,N_15107,N_15135);
nand U15429 (N_15429,N_15204,N_15158);
nand U15430 (N_15430,N_15107,N_15104);
nor U15431 (N_15431,N_15088,N_15044);
and U15432 (N_15432,N_15000,N_15115);
nor U15433 (N_15433,N_15123,N_15165);
nor U15434 (N_15434,N_15155,N_15012);
nand U15435 (N_15435,N_15090,N_15140);
or U15436 (N_15436,N_15157,N_15035);
nand U15437 (N_15437,N_15042,N_15145);
xor U15438 (N_15438,N_15241,N_15196);
nand U15439 (N_15439,N_15020,N_15023);
nor U15440 (N_15440,N_15007,N_15061);
and U15441 (N_15441,N_15145,N_15147);
nor U15442 (N_15442,N_15070,N_15016);
and U15443 (N_15443,N_15217,N_15239);
xor U15444 (N_15444,N_15044,N_15069);
nand U15445 (N_15445,N_15117,N_15088);
and U15446 (N_15446,N_15216,N_15154);
and U15447 (N_15447,N_15127,N_15248);
or U15448 (N_15448,N_15061,N_15108);
nor U15449 (N_15449,N_15037,N_15166);
nor U15450 (N_15450,N_15022,N_15066);
nand U15451 (N_15451,N_15121,N_15162);
or U15452 (N_15452,N_15244,N_15196);
nor U15453 (N_15453,N_15035,N_15093);
nor U15454 (N_15454,N_15066,N_15001);
and U15455 (N_15455,N_15162,N_15192);
nand U15456 (N_15456,N_15212,N_15102);
nand U15457 (N_15457,N_15025,N_15096);
nand U15458 (N_15458,N_15227,N_15110);
or U15459 (N_15459,N_15018,N_15031);
xnor U15460 (N_15460,N_15196,N_15208);
nand U15461 (N_15461,N_15054,N_15221);
or U15462 (N_15462,N_15215,N_15216);
nor U15463 (N_15463,N_15092,N_15132);
xor U15464 (N_15464,N_15070,N_15163);
nand U15465 (N_15465,N_15105,N_15045);
xor U15466 (N_15466,N_15022,N_15026);
nor U15467 (N_15467,N_15133,N_15142);
xor U15468 (N_15468,N_15243,N_15247);
and U15469 (N_15469,N_15086,N_15118);
nand U15470 (N_15470,N_15108,N_15003);
and U15471 (N_15471,N_15152,N_15120);
or U15472 (N_15472,N_15007,N_15169);
nand U15473 (N_15473,N_15046,N_15135);
xor U15474 (N_15474,N_15124,N_15098);
nand U15475 (N_15475,N_15049,N_15035);
or U15476 (N_15476,N_15131,N_15011);
nand U15477 (N_15477,N_15195,N_15013);
xor U15478 (N_15478,N_15135,N_15033);
or U15479 (N_15479,N_15158,N_15188);
nor U15480 (N_15480,N_15158,N_15146);
nand U15481 (N_15481,N_15092,N_15157);
or U15482 (N_15482,N_15246,N_15059);
nand U15483 (N_15483,N_15000,N_15177);
xor U15484 (N_15484,N_15188,N_15038);
xor U15485 (N_15485,N_15182,N_15130);
nand U15486 (N_15486,N_15140,N_15167);
xor U15487 (N_15487,N_15114,N_15035);
or U15488 (N_15488,N_15128,N_15194);
nor U15489 (N_15489,N_15105,N_15083);
xnor U15490 (N_15490,N_15044,N_15054);
nand U15491 (N_15491,N_15139,N_15092);
or U15492 (N_15492,N_15027,N_15095);
nor U15493 (N_15493,N_15001,N_15170);
nor U15494 (N_15494,N_15243,N_15222);
and U15495 (N_15495,N_15006,N_15014);
nor U15496 (N_15496,N_15092,N_15080);
or U15497 (N_15497,N_15204,N_15071);
and U15498 (N_15498,N_15126,N_15174);
xor U15499 (N_15499,N_15093,N_15073);
nand U15500 (N_15500,N_15338,N_15474);
nor U15501 (N_15501,N_15326,N_15453);
and U15502 (N_15502,N_15467,N_15476);
and U15503 (N_15503,N_15321,N_15360);
or U15504 (N_15504,N_15300,N_15442);
or U15505 (N_15505,N_15469,N_15389);
nor U15506 (N_15506,N_15373,N_15434);
or U15507 (N_15507,N_15271,N_15475);
nand U15508 (N_15508,N_15319,N_15375);
and U15509 (N_15509,N_15286,N_15262);
xnor U15510 (N_15510,N_15293,N_15345);
nor U15511 (N_15511,N_15334,N_15455);
nor U15512 (N_15512,N_15427,N_15342);
nand U15513 (N_15513,N_15330,N_15487);
nor U15514 (N_15514,N_15327,N_15371);
nand U15515 (N_15515,N_15409,N_15298);
and U15516 (N_15516,N_15329,N_15279);
and U15517 (N_15517,N_15464,N_15269);
nor U15518 (N_15518,N_15378,N_15454);
nor U15519 (N_15519,N_15395,N_15380);
nor U15520 (N_15520,N_15341,N_15420);
nor U15521 (N_15521,N_15445,N_15307);
nor U15522 (N_15522,N_15351,N_15408);
xnor U15523 (N_15523,N_15382,N_15448);
nor U15524 (N_15524,N_15496,N_15481);
or U15525 (N_15525,N_15361,N_15335);
nand U15526 (N_15526,N_15486,N_15302);
and U15527 (N_15527,N_15406,N_15374);
and U15528 (N_15528,N_15449,N_15436);
nand U15529 (N_15529,N_15272,N_15352);
nand U15530 (N_15530,N_15437,N_15290);
and U15531 (N_15531,N_15421,N_15441);
nor U15532 (N_15532,N_15337,N_15461);
or U15533 (N_15533,N_15462,N_15386);
or U15534 (N_15534,N_15383,N_15359);
and U15535 (N_15535,N_15425,N_15484);
nor U15536 (N_15536,N_15365,N_15324);
nand U15537 (N_15537,N_15430,N_15491);
and U15538 (N_15538,N_15276,N_15438);
or U15539 (N_15539,N_15277,N_15299);
nor U15540 (N_15540,N_15312,N_15424);
and U15541 (N_15541,N_15384,N_15363);
xnor U15542 (N_15542,N_15468,N_15369);
xnor U15543 (N_15543,N_15344,N_15499);
and U15544 (N_15544,N_15465,N_15282);
nor U15545 (N_15545,N_15364,N_15419);
or U15546 (N_15546,N_15372,N_15405);
xnor U15547 (N_15547,N_15291,N_15447);
xor U15548 (N_15548,N_15376,N_15393);
or U15549 (N_15549,N_15452,N_15460);
nand U15550 (N_15550,N_15265,N_15317);
nor U15551 (N_15551,N_15422,N_15349);
nor U15552 (N_15552,N_15332,N_15309);
and U15553 (N_15553,N_15331,N_15398);
or U15554 (N_15554,N_15478,N_15489);
xor U15555 (N_15555,N_15370,N_15367);
or U15556 (N_15556,N_15350,N_15274);
nor U15557 (N_15557,N_15368,N_15259);
or U15558 (N_15558,N_15253,N_15325);
xor U15559 (N_15559,N_15417,N_15250);
and U15560 (N_15560,N_15252,N_15428);
nand U15561 (N_15561,N_15366,N_15463);
nand U15562 (N_15562,N_15261,N_15308);
or U15563 (N_15563,N_15459,N_15355);
nand U15564 (N_15564,N_15358,N_15268);
nand U15565 (N_15565,N_15381,N_15314);
and U15566 (N_15566,N_15257,N_15347);
or U15567 (N_15567,N_15295,N_15429);
nand U15568 (N_15568,N_15494,N_15396);
xor U15569 (N_15569,N_15305,N_15480);
nand U15570 (N_15570,N_15426,N_15343);
xor U15571 (N_15571,N_15362,N_15391);
or U15572 (N_15572,N_15266,N_15403);
or U15573 (N_15573,N_15256,N_15336);
and U15574 (N_15574,N_15456,N_15485);
xnor U15575 (N_15575,N_15412,N_15303);
nand U15576 (N_15576,N_15353,N_15328);
nand U15577 (N_15577,N_15415,N_15388);
nor U15578 (N_15578,N_15411,N_15320);
xor U15579 (N_15579,N_15444,N_15400);
nor U15580 (N_15580,N_15280,N_15488);
or U15581 (N_15581,N_15479,N_15397);
and U15582 (N_15582,N_15493,N_15385);
or U15583 (N_15583,N_15323,N_15440);
nand U15584 (N_15584,N_15414,N_15258);
nand U15585 (N_15585,N_15313,N_15289);
and U15586 (N_15586,N_15275,N_15316);
or U15587 (N_15587,N_15435,N_15311);
xor U15588 (N_15588,N_15340,N_15285);
nor U15589 (N_15589,N_15315,N_15354);
and U15590 (N_15590,N_15357,N_15318);
nand U15591 (N_15591,N_15482,N_15457);
xnor U15592 (N_15592,N_15387,N_15281);
xnor U15593 (N_15593,N_15470,N_15423);
or U15594 (N_15594,N_15399,N_15377);
nor U15595 (N_15595,N_15339,N_15304);
xor U15596 (N_15596,N_15483,N_15410);
xnor U15597 (N_15597,N_15495,N_15283);
nor U15598 (N_15598,N_15413,N_15401);
nor U15599 (N_15599,N_15255,N_15477);
or U15600 (N_15600,N_15287,N_15294);
and U15601 (N_15601,N_15458,N_15322);
nand U15602 (N_15602,N_15292,N_15267);
or U15603 (N_15603,N_15450,N_15270);
or U15604 (N_15604,N_15379,N_15392);
nand U15605 (N_15605,N_15404,N_15284);
and U15606 (N_15606,N_15264,N_15490);
and U15607 (N_15607,N_15418,N_15296);
or U15608 (N_15608,N_15433,N_15492);
nand U15609 (N_15609,N_15443,N_15390);
xnor U15610 (N_15610,N_15446,N_15356);
and U15611 (N_15611,N_15278,N_15451);
nand U15612 (N_15612,N_15497,N_15297);
and U15613 (N_15613,N_15306,N_15333);
nor U15614 (N_15614,N_15471,N_15263);
and U15615 (N_15615,N_15432,N_15407);
nor U15616 (N_15616,N_15498,N_15348);
nor U15617 (N_15617,N_15431,N_15466);
xnor U15618 (N_15618,N_15251,N_15301);
xnor U15619 (N_15619,N_15472,N_15439);
or U15620 (N_15620,N_15394,N_15288);
and U15621 (N_15621,N_15254,N_15260);
and U15622 (N_15622,N_15402,N_15346);
and U15623 (N_15623,N_15273,N_15310);
and U15624 (N_15624,N_15416,N_15473);
nor U15625 (N_15625,N_15328,N_15263);
nand U15626 (N_15626,N_15359,N_15261);
xnor U15627 (N_15627,N_15383,N_15301);
or U15628 (N_15628,N_15476,N_15437);
xnor U15629 (N_15629,N_15495,N_15420);
nand U15630 (N_15630,N_15458,N_15476);
xnor U15631 (N_15631,N_15489,N_15327);
xor U15632 (N_15632,N_15498,N_15303);
or U15633 (N_15633,N_15360,N_15482);
and U15634 (N_15634,N_15424,N_15317);
nand U15635 (N_15635,N_15493,N_15405);
nor U15636 (N_15636,N_15331,N_15269);
nand U15637 (N_15637,N_15263,N_15289);
or U15638 (N_15638,N_15298,N_15437);
nor U15639 (N_15639,N_15301,N_15350);
and U15640 (N_15640,N_15347,N_15359);
or U15641 (N_15641,N_15264,N_15407);
and U15642 (N_15642,N_15312,N_15465);
xor U15643 (N_15643,N_15319,N_15279);
nand U15644 (N_15644,N_15391,N_15438);
xnor U15645 (N_15645,N_15270,N_15435);
xnor U15646 (N_15646,N_15386,N_15301);
and U15647 (N_15647,N_15445,N_15391);
or U15648 (N_15648,N_15396,N_15456);
xor U15649 (N_15649,N_15407,N_15473);
nand U15650 (N_15650,N_15447,N_15278);
nand U15651 (N_15651,N_15418,N_15309);
xnor U15652 (N_15652,N_15372,N_15439);
or U15653 (N_15653,N_15367,N_15403);
or U15654 (N_15654,N_15318,N_15282);
and U15655 (N_15655,N_15468,N_15367);
and U15656 (N_15656,N_15436,N_15419);
or U15657 (N_15657,N_15402,N_15425);
nand U15658 (N_15658,N_15272,N_15489);
or U15659 (N_15659,N_15260,N_15308);
and U15660 (N_15660,N_15467,N_15444);
nand U15661 (N_15661,N_15271,N_15305);
or U15662 (N_15662,N_15328,N_15338);
xor U15663 (N_15663,N_15387,N_15486);
nor U15664 (N_15664,N_15419,N_15352);
and U15665 (N_15665,N_15374,N_15282);
nand U15666 (N_15666,N_15496,N_15480);
nand U15667 (N_15667,N_15253,N_15371);
nand U15668 (N_15668,N_15369,N_15385);
nor U15669 (N_15669,N_15379,N_15334);
nand U15670 (N_15670,N_15328,N_15295);
and U15671 (N_15671,N_15404,N_15459);
or U15672 (N_15672,N_15334,N_15436);
xor U15673 (N_15673,N_15347,N_15491);
nor U15674 (N_15674,N_15407,N_15396);
nand U15675 (N_15675,N_15318,N_15364);
and U15676 (N_15676,N_15320,N_15291);
and U15677 (N_15677,N_15262,N_15443);
and U15678 (N_15678,N_15464,N_15427);
nand U15679 (N_15679,N_15470,N_15497);
nor U15680 (N_15680,N_15488,N_15342);
or U15681 (N_15681,N_15471,N_15342);
and U15682 (N_15682,N_15343,N_15433);
nor U15683 (N_15683,N_15454,N_15401);
or U15684 (N_15684,N_15386,N_15454);
or U15685 (N_15685,N_15360,N_15309);
or U15686 (N_15686,N_15401,N_15311);
xor U15687 (N_15687,N_15333,N_15301);
nand U15688 (N_15688,N_15276,N_15433);
xnor U15689 (N_15689,N_15275,N_15396);
nor U15690 (N_15690,N_15301,N_15332);
and U15691 (N_15691,N_15333,N_15481);
nor U15692 (N_15692,N_15311,N_15443);
or U15693 (N_15693,N_15405,N_15391);
xnor U15694 (N_15694,N_15314,N_15486);
and U15695 (N_15695,N_15445,N_15388);
nand U15696 (N_15696,N_15480,N_15404);
or U15697 (N_15697,N_15346,N_15470);
or U15698 (N_15698,N_15359,N_15443);
and U15699 (N_15699,N_15329,N_15272);
and U15700 (N_15700,N_15253,N_15485);
nor U15701 (N_15701,N_15417,N_15445);
or U15702 (N_15702,N_15328,N_15324);
nor U15703 (N_15703,N_15257,N_15298);
xor U15704 (N_15704,N_15308,N_15435);
or U15705 (N_15705,N_15379,N_15322);
nor U15706 (N_15706,N_15425,N_15407);
or U15707 (N_15707,N_15331,N_15424);
xor U15708 (N_15708,N_15276,N_15344);
nor U15709 (N_15709,N_15443,N_15487);
xor U15710 (N_15710,N_15348,N_15379);
or U15711 (N_15711,N_15390,N_15468);
nand U15712 (N_15712,N_15379,N_15436);
nand U15713 (N_15713,N_15415,N_15389);
nand U15714 (N_15714,N_15256,N_15282);
xor U15715 (N_15715,N_15267,N_15349);
xor U15716 (N_15716,N_15278,N_15397);
and U15717 (N_15717,N_15250,N_15458);
nand U15718 (N_15718,N_15400,N_15262);
nor U15719 (N_15719,N_15263,N_15462);
nand U15720 (N_15720,N_15284,N_15273);
and U15721 (N_15721,N_15399,N_15467);
nand U15722 (N_15722,N_15316,N_15455);
or U15723 (N_15723,N_15480,N_15487);
and U15724 (N_15724,N_15376,N_15301);
xor U15725 (N_15725,N_15261,N_15274);
nand U15726 (N_15726,N_15380,N_15332);
or U15727 (N_15727,N_15393,N_15272);
or U15728 (N_15728,N_15344,N_15268);
nor U15729 (N_15729,N_15388,N_15403);
nand U15730 (N_15730,N_15454,N_15337);
xnor U15731 (N_15731,N_15426,N_15465);
nand U15732 (N_15732,N_15374,N_15277);
nand U15733 (N_15733,N_15439,N_15316);
nand U15734 (N_15734,N_15347,N_15258);
or U15735 (N_15735,N_15483,N_15367);
nor U15736 (N_15736,N_15444,N_15317);
nor U15737 (N_15737,N_15431,N_15496);
and U15738 (N_15738,N_15293,N_15464);
nand U15739 (N_15739,N_15311,N_15305);
and U15740 (N_15740,N_15322,N_15256);
xnor U15741 (N_15741,N_15282,N_15440);
and U15742 (N_15742,N_15375,N_15282);
nand U15743 (N_15743,N_15340,N_15423);
or U15744 (N_15744,N_15483,N_15450);
and U15745 (N_15745,N_15309,N_15400);
or U15746 (N_15746,N_15395,N_15333);
nor U15747 (N_15747,N_15414,N_15436);
or U15748 (N_15748,N_15362,N_15329);
or U15749 (N_15749,N_15455,N_15352);
or U15750 (N_15750,N_15577,N_15726);
nor U15751 (N_15751,N_15561,N_15510);
and U15752 (N_15752,N_15715,N_15656);
nand U15753 (N_15753,N_15595,N_15523);
nand U15754 (N_15754,N_15695,N_15692);
xor U15755 (N_15755,N_15526,N_15742);
and U15756 (N_15756,N_15628,N_15673);
and U15757 (N_15757,N_15560,N_15596);
and U15758 (N_15758,N_15698,N_15505);
nor U15759 (N_15759,N_15747,N_15566);
xnor U15760 (N_15760,N_15559,N_15614);
and U15761 (N_15761,N_15545,N_15705);
or U15762 (N_15762,N_15640,N_15589);
xnor U15763 (N_15763,N_15534,N_15645);
nor U15764 (N_15764,N_15603,N_15696);
nor U15765 (N_15765,N_15624,N_15634);
xnor U15766 (N_15766,N_15736,N_15513);
or U15767 (N_15767,N_15604,N_15611);
nand U15768 (N_15768,N_15518,N_15649);
xnor U15769 (N_15769,N_15722,N_15608);
nand U15770 (N_15770,N_15740,N_15519);
or U15771 (N_15771,N_15536,N_15667);
xnor U15772 (N_15772,N_15691,N_15514);
and U15773 (N_15773,N_15570,N_15633);
nor U15774 (N_15774,N_15659,N_15728);
xor U15775 (N_15775,N_15627,N_15675);
nor U15776 (N_15776,N_15732,N_15527);
nor U15777 (N_15777,N_15708,N_15565);
xnor U15778 (N_15778,N_15644,N_15503);
xor U15779 (N_15779,N_15632,N_15672);
nor U15780 (N_15780,N_15593,N_15583);
nor U15781 (N_15781,N_15552,N_15701);
nor U15782 (N_15782,N_15509,N_15525);
nor U15783 (N_15783,N_15576,N_15548);
nor U15784 (N_15784,N_15630,N_15662);
or U15785 (N_15785,N_15617,N_15504);
nor U15786 (N_15786,N_15746,N_15569);
nor U15787 (N_15787,N_15506,N_15616);
or U15788 (N_15788,N_15606,N_15626);
or U15789 (N_15789,N_15739,N_15658);
and U15790 (N_15790,N_15621,N_15674);
or U15791 (N_15791,N_15597,N_15605);
and U15792 (N_15792,N_15648,N_15592);
and U15793 (N_15793,N_15719,N_15524);
xnor U15794 (N_15794,N_15749,N_15613);
or U15795 (N_15795,N_15680,N_15584);
and U15796 (N_15796,N_15643,N_15546);
xnor U15797 (N_15797,N_15620,N_15538);
xnor U15798 (N_15798,N_15501,N_15636);
xor U15799 (N_15799,N_15718,N_15600);
and U15800 (N_15800,N_15684,N_15744);
and U15801 (N_15801,N_15530,N_15661);
or U15802 (N_15802,N_15664,N_15670);
and U15803 (N_15803,N_15688,N_15712);
nor U15804 (N_15804,N_15727,N_15725);
xor U15805 (N_15805,N_15591,N_15567);
and U15806 (N_15806,N_15623,N_15553);
nand U15807 (N_15807,N_15544,N_15689);
or U15808 (N_15808,N_15535,N_15533);
xnor U15809 (N_15809,N_15655,N_15599);
xnor U15810 (N_15810,N_15682,N_15709);
nand U15811 (N_15811,N_15653,N_15657);
nand U15812 (N_15812,N_15685,N_15641);
nand U15813 (N_15813,N_15511,N_15529);
xnor U15814 (N_15814,N_15517,N_15502);
nor U15815 (N_15815,N_15637,N_15532);
nor U15816 (N_15816,N_15598,N_15550);
nand U15817 (N_15817,N_15619,N_15687);
xnor U15818 (N_15818,N_15690,N_15723);
and U15819 (N_15819,N_15607,N_15717);
nand U15820 (N_15820,N_15683,N_15706);
or U15821 (N_15821,N_15587,N_15639);
nand U15822 (N_15822,N_15555,N_15549);
xnor U15823 (N_15823,N_15515,N_15573);
or U15824 (N_15824,N_15729,N_15651);
nor U15825 (N_15825,N_15730,N_15563);
nand U15826 (N_15826,N_15699,N_15716);
xor U15827 (N_15827,N_15542,N_15528);
nor U15828 (N_15828,N_15676,N_15590);
or U15829 (N_15829,N_15671,N_15520);
nor U15830 (N_15830,N_15582,N_15713);
and U15831 (N_15831,N_15694,N_15721);
nor U15832 (N_15832,N_15541,N_15660);
xnor U15833 (N_15833,N_15646,N_15678);
and U15834 (N_15834,N_15700,N_15724);
nand U15835 (N_15835,N_15558,N_15586);
nand U15836 (N_15836,N_15642,N_15602);
or U15837 (N_15837,N_15562,N_15625);
and U15838 (N_15838,N_15697,N_15663);
and U15839 (N_15839,N_15512,N_15737);
xnor U15840 (N_15840,N_15652,N_15635);
and U15841 (N_15841,N_15572,N_15669);
and U15842 (N_15842,N_15571,N_15703);
nand U15843 (N_15843,N_15609,N_15745);
and U15844 (N_15844,N_15588,N_15508);
or U15845 (N_15845,N_15734,N_15551);
xnor U15846 (N_15846,N_15579,N_15522);
nor U15847 (N_15847,N_15638,N_15539);
nor U15848 (N_15848,N_15557,N_15650);
nor U15849 (N_15849,N_15629,N_15547);
xor U15850 (N_15850,N_15578,N_15720);
nor U15851 (N_15851,N_15540,N_15580);
xnor U15852 (N_15852,N_15615,N_15601);
nand U15853 (N_15853,N_15679,N_15585);
or U15854 (N_15854,N_15707,N_15516);
nand U15855 (N_15855,N_15738,N_15735);
or U15856 (N_15856,N_15686,N_15647);
and U15857 (N_15857,N_15710,N_15564);
xor U15858 (N_15858,N_15568,N_15631);
xor U15859 (N_15859,N_15677,N_15556);
xnor U15860 (N_15860,N_15654,N_15612);
xor U15861 (N_15861,N_15711,N_15554);
and U15862 (N_15862,N_15521,N_15575);
and U15863 (N_15863,N_15704,N_15543);
and U15864 (N_15864,N_15714,N_15741);
nor U15865 (N_15865,N_15702,N_15743);
or U15866 (N_15866,N_15731,N_15693);
and U15867 (N_15867,N_15622,N_15610);
nand U15868 (N_15868,N_15500,N_15537);
nand U15869 (N_15869,N_15665,N_15733);
nor U15870 (N_15870,N_15618,N_15666);
nor U15871 (N_15871,N_15581,N_15668);
nor U15872 (N_15872,N_15507,N_15594);
and U15873 (N_15873,N_15681,N_15531);
or U15874 (N_15874,N_15748,N_15574);
or U15875 (N_15875,N_15691,N_15611);
nand U15876 (N_15876,N_15623,N_15668);
xnor U15877 (N_15877,N_15534,N_15518);
nor U15878 (N_15878,N_15541,N_15652);
xor U15879 (N_15879,N_15548,N_15607);
or U15880 (N_15880,N_15595,N_15579);
nand U15881 (N_15881,N_15526,N_15738);
xor U15882 (N_15882,N_15570,N_15593);
and U15883 (N_15883,N_15531,N_15732);
or U15884 (N_15884,N_15577,N_15554);
nand U15885 (N_15885,N_15566,N_15564);
or U15886 (N_15886,N_15727,N_15559);
and U15887 (N_15887,N_15667,N_15601);
xor U15888 (N_15888,N_15672,N_15667);
xor U15889 (N_15889,N_15540,N_15732);
or U15890 (N_15890,N_15681,N_15698);
and U15891 (N_15891,N_15747,N_15512);
or U15892 (N_15892,N_15691,N_15549);
or U15893 (N_15893,N_15592,N_15636);
nand U15894 (N_15894,N_15580,N_15624);
and U15895 (N_15895,N_15580,N_15745);
xnor U15896 (N_15896,N_15568,N_15538);
and U15897 (N_15897,N_15607,N_15591);
or U15898 (N_15898,N_15615,N_15594);
xor U15899 (N_15899,N_15547,N_15661);
nand U15900 (N_15900,N_15709,N_15678);
xor U15901 (N_15901,N_15658,N_15670);
xor U15902 (N_15902,N_15572,N_15571);
nand U15903 (N_15903,N_15747,N_15706);
or U15904 (N_15904,N_15673,N_15687);
or U15905 (N_15905,N_15669,N_15713);
and U15906 (N_15906,N_15718,N_15643);
nand U15907 (N_15907,N_15595,N_15584);
or U15908 (N_15908,N_15626,N_15600);
or U15909 (N_15909,N_15730,N_15569);
nand U15910 (N_15910,N_15720,N_15595);
nand U15911 (N_15911,N_15572,N_15516);
or U15912 (N_15912,N_15616,N_15613);
nand U15913 (N_15913,N_15641,N_15623);
and U15914 (N_15914,N_15605,N_15501);
and U15915 (N_15915,N_15658,N_15702);
and U15916 (N_15916,N_15583,N_15670);
nor U15917 (N_15917,N_15706,N_15578);
nor U15918 (N_15918,N_15554,N_15683);
nor U15919 (N_15919,N_15641,N_15512);
nor U15920 (N_15920,N_15715,N_15653);
nand U15921 (N_15921,N_15575,N_15525);
nand U15922 (N_15922,N_15575,N_15667);
nand U15923 (N_15923,N_15605,N_15682);
xor U15924 (N_15924,N_15546,N_15647);
xnor U15925 (N_15925,N_15538,N_15666);
and U15926 (N_15926,N_15518,N_15702);
nor U15927 (N_15927,N_15578,N_15708);
nor U15928 (N_15928,N_15730,N_15528);
or U15929 (N_15929,N_15699,N_15568);
nor U15930 (N_15930,N_15619,N_15722);
nand U15931 (N_15931,N_15728,N_15562);
and U15932 (N_15932,N_15747,N_15515);
or U15933 (N_15933,N_15563,N_15725);
and U15934 (N_15934,N_15560,N_15670);
nor U15935 (N_15935,N_15705,N_15723);
nor U15936 (N_15936,N_15662,N_15505);
nand U15937 (N_15937,N_15715,N_15604);
nand U15938 (N_15938,N_15712,N_15727);
or U15939 (N_15939,N_15655,N_15624);
nand U15940 (N_15940,N_15632,N_15710);
or U15941 (N_15941,N_15735,N_15602);
xor U15942 (N_15942,N_15630,N_15713);
nand U15943 (N_15943,N_15661,N_15548);
nor U15944 (N_15944,N_15619,N_15723);
xor U15945 (N_15945,N_15618,N_15745);
nand U15946 (N_15946,N_15597,N_15624);
xnor U15947 (N_15947,N_15558,N_15591);
nor U15948 (N_15948,N_15736,N_15679);
and U15949 (N_15949,N_15610,N_15535);
or U15950 (N_15950,N_15670,N_15739);
and U15951 (N_15951,N_15595,N_15589);
nand U15952 (N_15952,N_15541,N_15592);
nand U15953 (N_15953,N_15647,N_15563);
or U15954 (N_15954,N_15622,N_15687);
nor U15955 (N_15955,N_15653,N_15587);
or U15956 (N_15956,N_15647,N_15672);
or U15957 (N_15957,N_15743,N_15682);
nor U15958 (N_15958,N_15549,N_15723);
nand U15959 (N_15959,N_15640,N_15538);
xor U15960 (N_15960,N_15570,N_15691);
xnor U15961 (N_15961,N_15537,N_15642);
xor U15962 (N_15962,N_15701,N_15539);
xor U15963 (N_15963,N_15505,N_15528);
or U15964 (N_15964,N_15724,N_15675);
nand U15965 (N_15965,N_15747,N_15655);
and U15966 (N_15966,N_15661,N_15743);
nor U15967 (N_15967,N_15657,N_15586);
nor U15968 (N_15968,N_15702,N_15622);
nor U15969 (N_15969,N_15710,N_15706);
and U15970 (N_15970,N_15668,N_15554);
xnor U15971 (N_15971,N_15637,N_15571);
nand U15972 (N_15972,N_15571,N_15589);
and U15973 (N_15973,N_15719,N_15628);
and U15974 (N_15974,N_15724,N_15641);
nor U15975 (N_15975,N_15520,N_15628);
xor U15976 (N_15976,N_15568,N_15662);
and U15977 (N_15977,N_15502,N_15503);
nand U15978 (N_15978,N_15740,N_15603);
xnor U15979 (N_15979,N_15717,N_15691);
and U15980 (N_15980,N_15541,N_15702);
nand U15981 (N_15981,N_15663,N_15527);
nand U15982 (N_15982,N_15650,N_15655);
and U15983 (N_15983,N_15697,N_15510);
xnor U15984 (N_15984,N_15512,N_15637);
or U15985 (N_15985,N_15562,N_15660);
and U15986 (N_15986,N_15606,N_15543);
nor U15987 (N_15987,N_15693,N_15681);
xnor U15988 (N_15988,N_15640,N_15587);
nor U15989 (N_15989,N_15743,N_15667);
or U15990 (N_15990,N_15579,N_15698);
xor U15991 (N_15991,N_15556,N_15568);
nand U15992 (N_15992,N_15513,N_15568);
xnor U15993 (N_15993,N_15659,N_15718);
and U15994 (N_15994,N_15675,N_15585);
xor U15995 (N_15995,N_15654,N_15633);
nor U15996 (N_15996,N_15602,N_15514);
and U15997 (N_15997,N_15628,N_15511);
nand U15998 (N_15998,N_15740,N_15555);
or U15999 (N_15999,N_15662,N_15669);
nand U16000 (N_16000,N_15837,N_15765);
and U16001 (N_16001,N_15873,N_15846);
xnor U16002 (N_16002,N_15754,N_15912);
xor U16003 (N_16003,N_15920,N_15780);
and U16004 (N_16004,N_15889,N_15982);
nor U16005 (N_16005,N_15805,N_15966);
and U16006 (N_16006,N_15813,N_15833);
nand U16007 (N_16007,N_15849,N_15932);
or U16008 (N_16008,N_15862,N_15801);
or U16009 (N_16009,N_15838,N_15914);
nand U16010 (N_16010,N_15972,N_15760);
nand U16011 (N_16011,N_15941,N_15935);
nor U16012 (N_16012,N_15855,N_15767);
xor U16013 (N_16013,N_15939,N_15943);
nor U16014 (N_16014,N_15953,N_15825);
xor U16015 (N_16015,N_15913,N_15870);
or U16016 (N_16016,N_15836,N_15865);
nor U16017 (N_16017,N_15869,N_15860);
and U16018 (N_16018,N_15844,N_15950);
nor U16019 (N_16019,N_15830,N_15887);
and U16020 (N_16020,N_15979,N_15964);
and U16021 (N_16021,N_15973,N_15917);
and U16022 (N_16022,N_15909,N_15867);
and U16023 (N_16023,N_15751,N_15930);
and U16024 (N_16024,N_15794,N_15821);
xor U16025 (N_16025,N_15775,N_15814);
and U16026 (N_16026,N_15901,N_15880);
nand U16027 (N_16027,N_15802,N_15940);
or U16028 (N_16028,N_15835,N_15808);
nor U16029 (N_16029,N_15905,N_15904);
nand U16030 (N_16030,N_15759,N_15993);
xor U16031 (N_16031,N_15876,N_15755);
nor U16032 (N_16032,N_15809,N_15826);
or U16033 (N_16033,N_15792,N_15992);
nor U16034 (N_16034,N_15753,N_15965);
or U16035 (N_16035,N_15791,N_15827);
xor U16036 (N_16036,N_15881,N_15858);
xnor U16037 (N_16037,N_15757,N_15763);
nand U16038 (N_16038,N_15817,N_15895);
and U16039 (N_16039,N_15848,N_15758);
or U16040 (N_16040,N_15863,N_15978);
and U16041 (N_16041,N_15946,N_15888);
xnor U16042 (N_16042,N_15958,N_15828);
nand U16043 (N_16043,N_15971,N_15892);
or U16044 (N_16044,N_15975,N_15985);
xnor U16045 (N_16045,N_15877,N_15991);
nor U16046 (N_16046,N_15852,N_15756);
and U16047 (N_16047,N_15918,N_15994);
xor U16048 (N_16048,N_15797,N_15879);
and U16049 (N_16049,N_15776,N_15786);
xor U16050 (N_16050,N_15771,N_15782);
and U16051 (N_16051,N_15926,N_15810);
nor U16052 (N_16052,N_15896,N_15948);
or U16053 (N_16053,N_15960,N_15954);
nand U16054 (N_16054,N_15764,N_15842);
or U16055 (N_16055,N_15929,N_15777);
or U16056 (N_16056,N_15807,N_15798);
xor U16057 (N_16057,N_15897,N_15822);
and U16058 (N_16058,N_15785,N_15853);
or U16059 (N_16059,N_15894,N_15968);
xnor U16060 (N_16060,N_15871,N_15937);
or U16061 (N_16061,N_15772,N_15902);
and U16062 (N_16062,N_15882,N_15866);
and U16063 (N_16063,N_15883,N_15967);
nor U16064 (N_16064,N_15773,N_15944);
or U16065 (N_16065,N_15885,N_15899);
nor U16066 (N_16066,N_15996,N_15959);
nor U16067 (N_16067,N_15750,N_15784);
nor U16068 (N_16068,N_15951,N_15819);
or U16069 (N_16069,N_15795,N_15911);
nor U16070 (N_16070,N_15970,N_15816);
nor U16071 (N_16071,N_15980,N_15924);
nor U16072 (N_16072,N_15793,N_15768);
xnor U16073 (N_16073,N_15872,N_15952);
xor U16074 (N_16074,N_15987,N_15977);
nor U16075 (N_16075,N_15942,N_15840);
nand U16076 (N_16076,N_15799,N_15997);
or U16077 (N_16077,N_15824,N_15803);
nor U16078 (N_16078,N_15878,N_15936);
xor U16079 (N_16079,N_15823,N_15857);
nor U16080 (N_16080,N_15990,N_15778);
nand U16081 (N_16081,N_15783,N_15986);
and U16082 (N_16082,N_15752,N_15963);
xor U16083 (N_16083,N_15893,N_15834);
nor U16084 (N_16084,N_15974,N_15850);
or U16085 (N_16085,N_15845,N_15875);
or U16086 (N_16086,N_15999,N_15998);
or U16087 (N_16087,N_15961,N_15770);
nor U16088 (N_16088,N_15787,N_15923);
or U16089 (N_16089,N_15956,N_15934);
xor U16090 (N_16090,N_15839,N_15864);
nor U16091 (N_16091,N_15938,N_15910);
nor U16092 (N_16092,N_15890,N_15800);
and U16093 (N_16093,N_15829,N_15925);
and U16094 (N_16094,N_15891,N_15989);
or U16095 (N_16095,N_15811,N_15957);
xnor U16096 (N_16096,N_15774,N_15818);
xnor U16097 (N_16097,N_15898,N_15928);
nor U16098 (N_16098,N_15841,N_15812);
nor U16099 (N_16099,N_15900,N_15804);
xor U16100 (N_16100,N_15922,N_15886);
and U16101 (N_16101,N_15796,N_15945);
xor U16102 (N_16102,N_15907,N_15859);
nor U16103 (N_16103,N_15995,N_15927);
and U16104 (N_16104,N_15781,N_15919);
or U16105 (N_16105,N_15984,N_15779);
xnor U16106 (N_16106,N_15868,N_15788);
and U16107 (N_16107,N_15847,N_15988);
nor U16108 (N_16108,N_15806,N_15851);
xor U16109 (N_16109,N_15761,N_15962);
nor U16110 (N_16110,N_15769,N_15884);
or U16111 (N_16111,N_15931,N_15908);
and U16112 (N_16112,N_15861,N_15915);
xnor U16113 (N_16113,N_15947,N_15832);
xnor U16114 (N_16114,N_15933,N_15921);
nand U16115 (N_16115,N_15983,N_15762);
xor U16116 (N_16116,N_15906,N_15969);
xnor U16117 (N_16117,N_15903,N_15981);
and U16118 (N_16118,N_15976,N_15843);
nand U16119 (N_16119,N_15874,N_15790);
nor U16120 (N_16120,N_15815,N_15831);
or U16121 (N_16121,N_15916,N_15820);
or U16122 (N_16122,N_15856,N_15949);
and U16123 (N_16123,N_15854,N_15955);
xor U16124 (N_16124,N_15766,N_15789);
xnor U16125 (N_16125,N_15892,N_15845);
or U16126 (N_16126,N_15867,N_15858);
xnor U16127 (N_16127,N_15768,N_15846);
nand U16128 (N_16128,N_15871,N_15880);
or U16129 (N_16129,N_15849,N_15997);
xnor U16130 (N_16130,N_15830,N_15778);
nand U16131 (N_16131,N_15819,N_15815);
nor U16132 (N_16132,N_15882,N_15976);
nand U16133 (N_16133,N_15758,N_15762);
nand U16134 (N_16134,N_15966,N_15884);
nand U16135 (N_16135,N_15829,N_15833);
nor U16136 (N_16136,N_15790,N_15882);
nor U16137 (N_16137,N_15827,N_15988);
nor U16138 (N_16138,N_15836,N_15846);
nand U16139 (N_16139,N_15820,N_15940);
and U16140 (N_16140,N_15967,N_15878);
nand U16141 (N_16141,N_15886,N_15994);
nor U16142 (N_16142,N_15916,N_15755);
nand U16143 (N_16143,N_15921,N_15785);
and U16144 (N_16144,N_15891,N_15866);
and U16145 (N_16145,N_15969,N_15767);
nor U16146 (N_16146,N_15866,N_15999);
or U16147 (N_16147,N_15990,N_15829);
and U16148 (N_16148,N_15910,N_15952);
nand U16149 (N_16149,N_15999,N_15782);
or U16150 (N_16150,N_15752,N_15912);
and U16151 (N_16151,N_15752,N_15823);
xnor U16152 (N_16152,N_15937,N_15991);
nand U16153 (N_16153,N_15769,N_15936);
xnor U16154 (N_16154,N_15857,N_15769);
nor U16155 (N_16155,N_15864,N_15913);
nor U16156 (N_16156,N_15929,N_15916);
nand U16157 (N_16157,N_15783,N_15905);
xnor U16158 (N_16158,N_15822,N_15962);
and U16159 (N_16159,N_15922,N_15767);
or U16160 (N_16160,N_15925,N_15903);
nor U16161 (N_16161,N_15951,N_15833);
and U16162 (N_16162,N_15773,N_15904);
or U16163 (N_16163,N_15904,N_15802);
xnor U16164 (N_16164,N_15989,N_15898);
nor U16165 (N_16165,N_15784,N_15812);
nor U16166 (N_16166,N_15943,N_15888);
and U16167 (N_16167,N_15766,N_15843);
xor U16168 (N_16168,N_15884,N_15887);
xnor U16169 (N_16169,N_15775,N_15970);
nor U16170 (N_16170,N_15788,N_15960);
xnor U16171 (N_16171,N_15776,N_15817);
or U16172 (N_16172,N_15811,N_15834);
xnor U16173 (N_16173,N_15780,N_15983);
and U16174 (N_16174,N_15823,N_15829);
or U16175 (N_16175,N_15784,N_15789);
nor U16176 (N_16176,N_15817,N_15752);
and U16177 (N_16177,N_15893,N_15820);
and U16178 (N_16178,N_15757,N_15844);
nand U16179 (N_16179,N_15793,N_15860);
or U16180 (N_16180,N_15827,N_15817);
xor U16181 (N_16181,N_15788,N_15834);
and U16182 (N_16182,N_15950,N_15871);
and U16183 (N_16183,N_15989,N_15851);
and U16184 (N_16184,N_15885,N_15973);
nand U16185 (N_16185,N_15925,N_15935);
xor U16186 (N_16186,N_15787,N_15842);
and U16187 (N_16187,N_15926,N_15769);
and U16188 (N_16188,N_15904,N_15804);
and U16189 (N_16189,N_15963,N_15914);
and U16190 (N_16190,N_15945,N_15940);
xor U16191 (N_16191,N_15821,N_15918);
or U16192 (N_16192,N_15897,N_15796);
and U16193 (N_16193,N_15885,N_15910);
and U16194 (N_16194,N_15801,N_15917);
or U16195 (N_16195,N_15857,N_15906);
and U16196 (N_16196,N_15934,N_15962);
or U16197 (N_16197,N_15958,N_15825);
nand U16198 (N_16198,N_15958,N_15966);
or U16199 (N_16199,N_15774,N_15867);
xor U16200 (N_16200,N_15822,N_15913);
nand U16201 (N_16201,N_15945,N_15987);
and U16202 (N_16202,N_15940,N_15773);
and U16203 (N_16203,N_15824,N_15861);
nand U16204 (N_16204,N_15976,N_15771);
and U16205 (N_16205,N_15954,N_15969);
nand U16206 (N_16206,N_15803,N_15887);
nand U16207 (N_16207,N_15759,N_15767);
and U16208 (N_16208,N_15812,N_15818);
nor U16209 (N_16209,N_15890,N_15756);
xnor U16210 (N_16210,N_15936,N_15932);
xor U16211 (N_16211,N_15790,N_15911);
nand U16212 (N_16212,N_15841,N_15977);
or U16213 (N_16213,N_15815,N_15997);
nand U16214 (N_16214,N_15917,N_15954);
and U16215 (N_16215,N_15823,N_15989);
nor U16216 (N_16216,N_15781,N_15929);
or U16217 (N_16217,N_15942,N_15820);
and U16218 (N_16218,N_15766,N_15904);
nand U16219 (N_16219,N_15972,N_15934);
xor U16220 (N_16220,N_15861,N_15878);
xnor U16221 (N_16221,N_15917,N_15906);
and U16222 (N_16222,N_15832,N_15935);
xor U16223 (N_16223,N_15872,N_15909);
and U16224 (N_16224,N_15974,N_15771);
nand U16225 (N_16225,N_15972,N_15921);
xnor U16226 (N_16226,N_15959,N_15947);
or U16227 (N_16227,N_15879,N_15844);
nor U16228 (N_16228,N_15832,N_15920);
or U16229 (N_16229,N_15816,N_15990);
xor U16230 (N_16230,N_15958,N_15905);
nand U16231 (N_16231,N_15997,N_15831);
and U16232 (N_16232,N_15968,N_15942);
nand U16233 (N_16233,N_15840,N_15900);
and U16234 (N_16234,N_15986,N_15965);
nor U16235 (N_16235,N_15939,N_15793);
nor U16236 (N_16236,N_15916,N_15927);
or U16237 (N_16237,N_15826,N_15996);
and U16238 (N_16238,N_15774,N_15937);
nand U16239 (N_16239,N_15780,N_15837);
nor U16240 (N_16240,N_15832,N_15946);
or U16241 (N_16241,N_15943,N_15914);
and U16242 (N_16242,N_15937,N_15777);
or U16243 (N_16243,N_15967,N_15995);
xnor U16244 (N_16244,N_15792,N_15899);
and U16245 (N_16245,N_15838,N_15807);
and U16246 (N_16246,N_15946,N_15917);
nand U16247 (N_16247,N_15868,N_15942);
and U16248 (N_16248,N_15804,N_15945);
or U16249 (N_16249,N_15906,N_15980);
or U16250 (N_16250,N_16156,N_16068);
nand U16251 (N_16251,N_16109,N_16143);
nor U16252 (N_16252,N_16102,N_16215);
or U16253 (N_16253,N_16036,N_16010);
or U16254 (N_16254,N_16058,N_16065);
or U16255 (N_16255,N_16218,N_16248);
xor U16256 (N_16256,N_16179,N_16008);
and U16257 (N_16257,N_16096,N_16124);
xnor U16258 (N_16258,N_16025,N_16024);
nand U16259 (N_16259,N_16000,N_16116);
nor U16260 (N_16260,N_16055,N_16052);
nor U16261 (N_16261,N_16163,N_16177);
nand U16262 (N_16262,N_16149,N_16095);
nand U16263 (N_16263,N_16172,N_16031);
and U16264 (N_16264,N_16233,N_16082);
nand U16265 (N_16265,N_16141,N_16127);
nor U16266 (N_16266,N_16070,N_16249);
and U16267 (N_16267,N_16171,N_16075);
and U16268 (N_16268,N_16184,N_16023);
nor U16269 (N_16269,N_16079,N_16067);
nor U16270 (N_16270,N_16132,N_16076);
or U16271 (N_16271,N_16244,N_16115);
or U16272 (N_16272,N_16080,N_16073);
nor U16273 (N_16273,N_16247,N_16018);
or U16274 (N_16274,N_16122,N_16016);
nor U16275 (N_16275,N_16190,N_16084);
and U16276 (N_16276,N_16140,N_16155);
or U16277 (N_16277,N_16027,N_16134);
or U16278 (N_16278,N_16221,N_16187);
and U16279 (N_16279,N_16212,N_16197);
and U16280 (N_16280,N_16222,N_16108);
xor U16281 (N_16281,N_16118,N_16189);
and U16282 (N_16282,N_16151,N_16200);
and U16283 (N_16283,N_16205,N_16195);
nand U16284 (N_16284,N_16167,N_16128);
or U16285 (N_16285,N_16029,N_16064);
or U16286 (N_16286,N_16093,N_16208);
nand U16287 (N_16287,N_16182,N_16135);
nand U16288 (N_16288,N_16107,N_16060);
nor U16289 (N_16289,N_16214,N_16130);
xor U16290 (N_16290,N_16168,N_16110);
nand U16291 (N_16291,N_16230,N_16239);
and U16292 (N_16292,N_16077,N_16012);
or U16293 (N_16293,N_16224,N_16150);
nand U16294 (N_16294,N_16198,N_16097);
xor U16295 (N_16295,N_16098,N_16015);
xnor U16296 (N_16296,N_16234,N_16046);
and U16297 (N_16297,N_16061,N_16086);
nand U16298 (N_16298,N_16188,N_16051);
nor U16299 (N_16299,N_16009,N_16074);
xor U16300 (N_16300,N_16039,N_16229);
or U16301 (N_16301,N_16170,N_16088);
xnor U16302 (N_16302,N_16069,N_16017);
nor U16303 (N_16303,N_16120,N_16131);
and U16304 (N_16304,N_16216,N_16196);
nand U16305 (N_16305,N_16228,N_16178);
or U16306 (N_16306,N_16014,N_16106);
or U16307 (N_16307,N_16174,N_16210);
xor U16308 (N_16308,N_16139,N_16213);
nand U16309 (N_16309,N_16243,N_16087);
or U16310 (N_16310,N_16091,N_16043);
or U16311 (N_16311,N_16137,N_16111);
nor U16312 (N_16312,N_16022,N_16162);
xor U16313 (N_16313,N_16083,N_16063);
nand U16314 (N_16314,N_16226,N_16159);
nand U16315 (N_16315,N_16147,N_16032);
and U16316 (N_16316,N_16125,N_16021);
nor U16317 (N_16317,N_16099,N_16081);
or U16318 (N_16318,N_16037,N_16053);
nor U16319 (N_16319,N_16185,N_16072);
nor U16320 (N_16320,N_16001,N_16047);
nor U16321 (N_16321,N_16209,N_16059);
xor U16322 (N_16322,N_16113,N_16042);
nor U16323 (N_16323,N_16175,N_16048);
and U16324 (N_16324,N_16003,N_16136);
xnor U16325 (N_16325,N_16237,N_16238);
and U16326 (N_16326,N_16211,N_16105);
and U16327 (N_16327,N_16103,N_16219);
and U16328 (N_16328,N_16246,N_16236);
xnor U16329 (N_16329,N_16166,N_16038);
and U16330 (N_16330,N_16245,N_16004);
nor U16331 (N_16331,N_16192,N_16202);
nand U16332 (N_16332,N_16041,N_16206);
or U16333 (N_16333,N_16158,N_16207);
xor U16334 (N_16334,N_16153,N_16176);
and U16335 (N_16335,N_16092,N_16054);
nor U16336 (N_16336,N_16089,N_16049);
and U16337 (N_16337,N_16181,N_16071);
xnor U16338 (N_16338,N_16006,N_16066);
and U16339 (N_16339,N_16028,N_16242);
and U16340 (N_16340,N_16056,N_16144);
xor U16341 (N_16341,N_16121,N_16160);
and U16342 (N_16342,N_16005,N_16138);
xor U16343 (N_16343,N_16191,N_16146);
nand U16344 (N_16344,N_16078,N_16157);
nor U16345 (N_16345,N_16044,N_16152);
xnor U16346 (N_16346,N_16045,N_16193);
nor U16347 (N_16347,N_16035,N_16094);
nor U16348 (N_16348,N_16057,N_16235);
nor U16349 (N_16349,N_16030,N_16104);
or U16350 (N_16350,N_16040,N_16164);
nand U16351 (N_16351,N_16148,N_16180);
or U16352 (N_16352,N_16241,N_16050);
nor U16353 (N_16353,N_16123,N_16165);
xor U16354 (N_16354,N_16154,N_16126);
nor U16355 (N_16355,N_16231,N_16062);
or U16356 (N_16356,N_16090,N_16101);
xnor U16357 (N_16357,N_16114,N_16227);
nor U16358 (N_16358,N_16129,N_16033);
and U16359 (N_16359,N_16199,N_16085);
nor U16360 (N_16360,N_16020,N_16026);
or U16361 (N_16361,N_16161,N_16183);
or U16362 (N_16362,N_16201,N_16220);
and U16363 (N_16363,N_16204,N_16186);
xnor U16364 (N_16364,N_16203,N_16173);
nand U16365 (N_16365,N_16240,N_16007);
and U16366 (N_16366,N_16225,N_16019);
nand U16367 (N_16367,N_16217,N_16112);
nor U16368 (N_16368,N_16002,N_16223);
xor U16369 (N_16369,N_16100,N_16119);
and U16370 (N_16370,N_16145,N_16034);
xor U16371 (N_16371,N_16194,N_16232);
xor U16372 (N_16372,N_16133,N_16169);
nand U16373 (N_16373,N_16142,N_16013);
nor U16374 (N_16374,N_16117,N_16011);
xor U16375 (N_16375,N_16028,N_16085);
or U16376 (N_16376,N_16084,N_16060);
nor U16377 (N_16377,N_16024,N_16089);
nand U16378 (N_16378,N_16119,N_16123);
nor U16379 (N_16379,N_16005,N_16033);
and U16380 (N_16380,N_16248,N_16181);
nor U16381 (N_16381,N_16216,N_16025);
nand U16382 (N_16382,N_16125,N_16212);
and U16383 (N_16383,N_16066,N_16187);
nand U16384 (N_16384,N_16049,N_16182);
nor U16385 (N_16385,N_16218,N_16063);
or U16386 (N_16386,N_16194,N_16089);
xor U16387 (N_16387,N_16035,N_16127);
xor U16388 (N_16388,N_16006,N_16011);
nor U16389 (N_16389,N_16067,N_16017);
nand U16390 (N_16390,N_16113,N_16174);
nor U16391 (N_16391,N_16146,N_16000);
xnor U16392 (N_16392,N_16175,N_16179);
and U16393 (N_16393,N_16183,N_16094);
and U16394 (N_16394,N_16110,N_16120);
or U16395 (N_16395,N_16072,N_16157);
xor U16396 (N_16396,N_16224,N_16107);
xor U16397 (N_16397,N_16131,N_16172);
xor U16398 (N_16398,N_16050,N_16207);
or U16399 (N_16399,N_16016,N_16152);
nand U16400 (N_16400,N_16162,N_16094);
and U16401 (N_16401,N_16038,N_16164);
nor U16402 (N_16402,N_16183,N_16182);
and U16403 (N_16403,N_16162,N_16206);
and U16404 (N_16404,N_16048,N_16197);
nor U16405 (N_16405,N_16032,N_16229);
xnor U16406 (N_16406,N_16045,N_16043);
or U16407 (N_16407,N_16197,N_16118);
xor U16408 (N_16408,N_16140,N_16053);
or U16409 (N_16409,N_16130,N_16172);
or U16410 (N_16410,N_16221,N_16159);
or U16411 (N_16411,N_16108,N_16037);
or U16412 (N_16412,N_16191,N_16027);
xnor U16413 (N_16413,N_16094,N_16123);
and U16414 (N_16414,N_16079,N_16021);
nor U16415 (N_16415,N_16238,N_16014);
or U16416 (N_16416,N_16052,N_16131);
or U16417 (N_16417,N_16232,N_16033);
nor U16418 (N_16418,N_16188,N_16111);
and U16419 (N_16419,N_16084,N_16069);
nor U16420 (N_16420,N_16164,N_16031);
nand U16421 (N_16421,N_16204,N_16061);
xnor U16422 (N_16422,N_16145,N_16020);
nor U16423 (N_16423,N_16199,N_16058);
nor U16424 (N_16424,N_16016,N_16153);
nor U16425 (N_16425,N_16081,N_16173);
and U16426 (N_16426,N_16074,N_16021);
nor U16427 (N_16427,N_16239,N_16027);
nor U16428 (N_16428,N_16146,N_16031);
or U16429 (N_16429,N_16071,N_16009);
or U16430 (N_16430,N_16193,N_16242);
and U16431 (N_16431,N_16059,N_16194);
or U16432 (N_16432,N_16216,N_16064);
xnor U16433 (N_16433,N_16155,N_16228);
or U16434 (N_16434,N_16160,N_16216);
and U16435 (N_16435,N_16031,N_16070);
and U16436 (N_16436,N_16172,N_16105);
or U16437 (N_16437,N_16034,N_16065);
nor U16438 (N_16438,N_16217,N_16110);
nand U16439 (N_16439,N_16161,N_16191);
or U16440 (N_16440,N_16187,N_16003);
nor U16441 (N_16441,N_16113,N_16013);
or U16442 (N_16442,N_16248,N_16019);
and U16443 (N_16443,N_16060,N_16158);
xor U16444 (N_16444,N_16068,N_16234);
nor U16445 (N_16445,N_16089,N_16129);
nand U16446 (N_16446,N_16046,N_16185);
nand U16447 (N_16447,N_16036,N_16134);
nor U16448 (N_16448,N_16093,N_16070);
nor U16449 (N_16449,N_16186,N_16000);
nand U16450 (N_16450,N_16140,N_16031);
and U16451 (N_16451,N_16158,N_16189);
and U16452 (N_16452,N_16068,N_16010);
nor U16453 (N_16453,N_16030,N_16084);
nand U16454 (N_16454,N_16181,N_16236);
xnor U16455 (N_16455,N_16171,N_16061);
nor U16456 (N_16456,N_16044,N_16213);
or U16457 (N_16457,N_16110,N_16245);
or U16458 (N_16458,N_16009,N_16209);
or U16459 (N_16459,N_16223,N_16238);
nand U16460 (N_16460,N_16197,N_16162);
or U16461 (N_16461,N_16146,N_16015);
and U16462 (N_16462,N_16179,N_16193);
and U16463 (N_16463,N_16196,N_16184);
xnor U16464 (N_16464,N_16161,N_16195);
and U16465 (N_16465,N_16119,N_16217);
nand U16466 (N_16466,N_16092,N_16129);
nor U16467 (N_16467,N_16245,N_16178);
or U16468 (N_16468,N_16247,N_16151);
xor U16469 (N_16469,N_16002,N_16032);
xor U16470 (N_16470,N_16030,N_16055);
or U16471 (N_16471,N_16205,N_16135);
xnor U16472 (N_16472,N_16228,N_16028);
or U16473 (N_16473,N_16145,N_16032);
and U16474 (N_16474,N_16176,N_16229);
nor U16475 (N_16475,N_16208,N_16175);
xnor U16476 (N_16476,N_16172,N_16041);
xnor U16477 (N_16477,N_16211,N_16197);
nand U16478 (N_16478,N_16131,N_16104);
nor U16479 (N_16479,N_16025,N_16189);
and U16480 (N_16480,N_16125,N_16186);
nand U16481 (N_16481,N_16167,N_16136);
nand U16482 (N_16482,N_16092,N_16235);
and U16483 (N_16483,N_16138,N_16011);
nand U16484 (N_16484,N_16231,N_16134);
nand U16485 (N_16485,N_16196,N_16193);
nor U16486 (N_16486,N_16055,N_16085);
xnor U16487 (N_16487,N_16128,N_16154);
xor U16488 (N_16488,N_16158,N_16067);
nor U16489 (N_16489,N_16069,N_16235);
or U16490 (N_16490,N_16130,N_16081);
or U16491 (N_16491,N_16230,N_16077);
or U16492 (N_16492,N_16098,N_16161);
and U16493 (N_16493,N_16165,N_16152);
xor U16494 (N_16494,N_16137,N_16246);
xnor U16495 (N_16495,N_16121,N_16074);
nor U16496 (N_16496,N_16111,N_16232);
or U16497 (N_16497,N_16113,N_16198);
nand U16498 (N_16498,N_16057,N_16219);
or U16499 (N_16499,N_16120,N_16182);
or U16500 (N_16500,N_16415,N_16394);
xnor U16501 (N_16501,N_16419,N_16347);
xnor U16502 (N_16502,N_16448,N_16316);
xnor U16503 (N_16503,N_16432,N_16405);
and U16504 (N_16504,N_16371,N_16367);
nor U16505 (N_16505,N_16327,N_16404);
nor U16506 (N_16506,N_16429,N_16477);
or U16507 (N_16507,N_16296,N_16331);
nor U16508 (N_16508,N_16355,N_16459);
xor U16509 (N_16509,N_16271,N_16441);
or U16510 (N_16510,N_16471,N_16254);
xor U16511 (N_16511,N_16291,N_16286);
xor U16512 (N_16512,N_16413,N_16285);
nor U16513 (N_16513,N_16489,N_16259);
xor U16514 (N_16514,N_16359,N_16378);
or U16515 (N_16515,N_16304,N_16434);
nor U16516 (N_16516,N_16388,N_16332);
nor U16517 (N_16517,N_16444,N_16476);
nand U16518 (N_16518,N_16402,N_16290);
nand U16519 (N_16519,N_16351,N_16474);
nand U16520 (N_16520,N_16426,N_16464);
xnor U16521 (N_16521,N_16467,N_16310);
or U16522 (N_16522,N_16366,N_16462);
or U16523 (N_16523,N_16491,N_16443);
or U16524 (N_16524,N_16365,N_16297);
nand U16525 (N_16525,N_16346,N_16356);
nor U16526 (N_16526,N_16401,N_16496);
nand U16527 (N_16527,N_16260,N_16452);
nor U16528 (N_16528,N_16383,N_16454);
nand U16529 (N_16529,N_16447,N_16412);
xor U16530 (N_16530,N_16435,N_16488);
nand U16531 (N_16531,N_16267,N_16486);
and U16532 (N_16532,N_16280,N_16484);
or U16533 (N_16533,N_16340,N_16362);
nor U16534 (N_16534,N_16320,N_16495);
or U16535 (N_16535,N_16470,N_16431);
nor U16536 (N_16536,N_16334,N_16483);
xnor U16537 (N_16537,N_16276,N_16348);
and U16538 (N_16538,N_16408,N_16480);
nand U16539 (N_16539,N_16257,N_16380);
nor U16540 (N_16540,N_16322,N_16328);
or U16541 (N_16541,N_16299,N_16256);
and U16542 (N_16542,N_16410,N_16397);
nand U16543 (N_16543,N_16363,N_16494);
nor U16544 (N_16544,N_16293,N_16272);
and U16545 (N_16545,N_16400,N_16427);
and U16546 (N_16546,N_16455,N_16349);
nor U16547 (N_16547,N_16330,N_16391);
and U16548 (N_16548,N_16460,N_16468);
or U16549 (N_16549,N_16485,N_16430);
and U16550 (N_16550,N_16321,N_16329);
xnor U16551 (N_16551,N_16399,N_16403);
nand U16552 (N_16552,N_16385,N_16428);
xor U16553 (N_16553,N_16255,N_16281);
and U16554 (N_16554,N_16418,N_16301);
or U16555 (N_16555,N_16481,N_16446);
or U16556 (N_16556,N_16354,N_16456);
nor U16557 (N_16557,N_16306,N_16416);
and U16558 (N_16558,N_16252,N_16466);
and U16559 (N_16559,N_16279,N_16294);
xor U16560 (N_16560,N_16493,N_16406);
nor U16561 (N_16561,N_16326,N_16323);
and U16562 (N_16562,N_16478,N_16337);
or U16563 (N_16563,N_16398,N_16386);
nand U16564 (N_16564,N_16372,N_16437);
nand U16565 (N_16565,N_16390,N_16449);
xnor U16566 (N_16566,N_16445,N_16357);
and U16567 (N_16567,N_16369,N_16439);
nand U16568 (N_16568,N_16475,N_16490);
nand U16569 (N_16569,N_16453,N_16457);
xnor U16570 (N_16570,N_16283,N_16343);
or U16571 (N_16571,N_16381,N_16287);
nand U16572 (N_16572,N_16451,N_16289);
nor U16573 (N_16573,N_16324,N_16487);
nand U16574 (N_16574,N_16463,N_16497);
xnor U16575 (N_16575,N_16325,N_16423);
or U16576 (N_16576,N_16374,N_16303);
and U16577 (N_16577,N_16305,N_16339);
xor U16578 (N_16578,N_16414,N_16472);
and U16579 (N_16579,N_16282,N_16433);
nand U16580 (N_16580,N_16436,N_16275);
nand U16581 (N_16581,N_16368,N_16269);
and U16582 (N_16582,N_16264,N_16440);
and U16583 (N_16583,N_16342,N_16450);
nand U16584 (N_16584,N_16392,N_16387);
and U16585 (N_16585,N_16319,N_16265);
nand U16586 (N_16586,N_16268,N_16379);
and U16587 (N_16587,N_16376,N_16407);
and U16588 (N_16588,N_16458,N_16424);
and U16589 (N_16589,N_16396,N_16422);
and U16590 (N_16590,N_16270,N_16312);
and U16591 (N_16591,N_16375,N_16314);
xnor U16592 (N_16592,N_16498,N_16262);
nand U16593 (N_16593,N_16482,N_16350);
or U16594 (N_16594,N_16352,N_16266);
xnor U16595 (N_16595,N_16382,N_16461);
xnor U16596 (N_16596,N_16344,N_16336);
or U16597 (N_16597,N_16317,N_16420);
nand U16598 (N_16598,N_16295,N_16499);
nor U16599 (N_16599,N_16341,N_16370);
xnor U16600 (N_16600,N_16309,N_16345);
xnor U16601 (N_16601,N_16438,N_16273);
xnor U16602 (N_16602,N_16421,N_16395);
nor U16603 (N_16603,N_16313,N_16250);
nor U16604 (N_16604,N_16417,N_16358);
nor U16605 (N_16605,N_16469,N_16318);
or U16606 (N_16606,N_16298,N_16251);
nor U16607 (N_16607,N_16278,N_16384);
and U16608 (N_16608,N_16307,N_16360);
nor U16609 (N_16609,N_16333,N_16253);
xnor U16610 (N_16610,N_16389,N_16261);
nor U16611 (N_16611,N_16393,N_16300);
and U16612 (N_16612,N_16274,N_16361);
or U16613 (N_16613,N_16473,N_16353);
and U16614 (N_16614,N_16364,N_16277);
nand U16615 (N_16615,N_16409,N_16442);
nand U16616 (N_16616,N_16258,N_16338);
and U16617 (N_16617,N_16315,N_16492);
nor U16618 (N_16618,N_16425,N_16288);
or U16619 (N_16619,N_16335,N_16373);
nor U16620 (N_16620,N_16292,N_16479);
xnor U16621 (N_16621,N_16308,N_16263);
xor U16622 (N_16622,N_16377,N_16311);
nor U16623 (N_16623,N_16465,N_16411);
xor U16624 (N_16624,N_16284,N_16302);
nor U16625 (N_16625,N_16300,N_16346);
and U16626 (N_16626,N_16434,N_16468);
or U16627 (N_16627,N_16277,N_16333);
or U16628 (N_16628,N_16456,N_16334);
nand U16629 (N_16629,N_16311,N_16426);
nor U16630 (N_16630,N_16300,N_16410);
nor U16631 (N_16631,N_16290,N_16358);
nand U16632 (N_16632,N_16253,N_16423);
nand U16633 (N_16633,N_16445,N_16434);
xnor U16634 (N_16634,N_16285,N_16480);
nor U16635 (N_16635,N_16360,N_16291);
or U16636 (N_16636,N_16446,N_16467);
and U16637 (N_16637,N_16370,N_16291);
nand U16638 (N_16638,N_16375,N_16470);
or U16639 (N_16639,N_16361,N_16416);
and U16640 (N_16640,N_16484,N_16436);
and U16641 (N_16641,N_16380,N_16463);
nand U16642 (N_16642,N_16358,N_16316);
or U16643 (N_16643,N_16285,N_16272);
xnor U16644 (N_16644,N_16345,N_16437);
or U16645 (N_16645,N_16319,N_16392);
nand U16646 (N_16646,N_16274,N_16429);
nor U16647 (N_16647,N_16253,N_16460);
xor U16648 (N_16648,N_16283,N_16448);
xor U16649 (N_16649,N_16318,N_16304);
nand U16650 (N_16650,N_16447,N_16352);
xnor U16651 (N_16651,N_16308,N_16487);
nor U16652 (N_16652,N_16413,N_16287);
xnor U16653 (N_16653,N_16369,N_16289);
and U16654 (N_16654,N_16489,N_16309);
or U16655 (N_16655,N_16389,N_16423);
xnor U16656 (N_16656,N_16252,N_16490);
nand U16657 (N_16657,N_16306,N_16412);
nand U16658 (N_16658,N_16346,N_16291);
nor U16659 (N_16659,N_16454,N_16470);
and U16660 (N_16660,N_16252,N_16365);
and U16661 (N_16661,N_16308,N_16312);
nor U16662 (N_16662,N_16469,N_16378);
xnor U16663 (N_16663,N_16441,N_16362);
or U16664 (N_16664,N_16416,N_16490);
nor U16665 (N_16665,N_16265,N_16407);
xor U16666 (N_16666,N_16445,N_16333);
nor U16667 (N_16667,N_16439,N_16345);
xnor U16668 (N_16668,N_16251,N_16401);
nand U16669 (N_16669,N_16374,N_16270);
nor U16670 (N_16670,N_16311,N_16314);
and U16671 (N_16671,N_16398,N_16341);
nand U16672 (N_16672,N_16259,N_16414);
or U16673 (N_16673,N_16419,N_16445);
xnor U16674 (N_16674,N_16428,N_16404);
nor U16675 (N_16675,N_16445,N_16364);
xnor U16676 (N_16676,N_16423,N_16391);
or U16677 (N_16677,N_16377,N_16380);
and U16678 (N_16678,N_16458,N_16438);
and U16679 (N_16679,N_16441,N_16436);
nand U16680 (N_16680,N_16483,N_16485);
nand U16681 (N_16681,N_16395,N_16423);
or U16682 (N_16682,N_16285,N_16281);
nor U16683 (N_16683,N_16263,N_16304);
or U16684 (N_16684,N_16378,N_16467);
or U16685 (N_16685,N_16371,N_16339);
or U16686 (N_16686,N_16267,N_16373);
or U16687 (N_16687,N_16333,N_16426);
nand U16688 (N_16688,N_16453,N_16317);
nand U16689 (N_16689,N_16271,N_16474);
nor U16690 (N_16690,N_16325,N_16482);
and U16691 (N_16691,N_16471,N_16381);
or U16692 (N_16692,N_16391,N_16377);
nor U16693 (N_16693,N_16391,N_16424);
and U16694 (N_16694,N_16462,N_16377);
xor U16695 (N_16695,N_16314,N_16481);
nand U16696 (N_16696,N_16447,N_16252);
or U16697 (N_16697,N_16259,N_16297);
nor U16698 (N_16698,N_16381,N_16483);
and U16699 (N_16699,N_16437,N_16359);
xnor U16700 (N_16700,N_16349,N_16378);
or U16701 (N_16701,N_16358,N_16476);
nor U16702 (N_16702,N_16478,N_16372);
or U16703 (N_16703,N_16492,N_16462);
and U16704 (N_16704,N_16317,N_16398);
and U16705 (N_16705,N_16367,N_16379);
or U16706 (N_16706,N_16280,N_16322);
or U16707 (N_16707,N_16407,N_16349);
xor U16708 (N_16708,N_16488,N_16273);
xnor U16709 (N_16709,N_16434,N_16408);
or U16710 (N_16710,N_16356,N_16306);
nor U16711 (N_16711,N_16475,N_16251);
xnor U16712 (N_16712,N_16445,N_16325);
nand U16713 (N_16713,N_16258,N_16490);
nand U16714 (N_16714,N_16420,N_16377);
or U16715 (N_16715,N_16269,N_16404);
and U16716 (N_16716,N_16447,N_16418);
nor U16717 (N_16717,N_16442,N_16438);
xor U16718 (N_16718,N_16250,N_16268);
nor U16719 (N_16719,N_16299,N_16287);
and U16720 (N_16720,N_16277,N_16412);
or U16721 (N_16721,N_16332,N_16462);
xor U16722 (N_16722,N_16430,N_16495);
and U16723 (N_16723,N_16494,N_16322);
or U16724 (N_16724,N_16349,N_16479);
or U16725 (N_16725,N_16308,N_16379);
xor U16726 (N_16726,N_16350,N_16287);
nor U16727 (N_16727,N_16374,N_16320);
xor U16728 (N_16728,N_16294,N_16391);
and U16729 (N_16729,N_16313,N_16328);
and U16730 (N_16730,N_16317,N_16328);
and U16731 (N_16731,N_16412,N_16301);
nand U16732 (N_16732,N_16490,N_16474);
or U16733 (N_16733,N_16335,N_16459);
and U16734 (N_16734,N_16387,N_16403);
nand U16735 (N_16735,N_16255,N_16302);
and U16736 (N_16736,N_16358,N_16402);
nand U16737 (N_16737,N_16417,N_16315);
nand U16738 (N_16738,N_16382,N_16410);
xor U16739 (N_16739,N_16258,N_16411);
nor U16740 (N_16740,N_16297,N_16449);
nand U16741 (N_16741,N_16277,N_16362);
nor U16742 (N_16742,N_16332,N_16351);
xnor U16743 (N_16743,N_16294,N_16342);
and U16744 (N_16744,N_16281,N_16466);
xnor U16745 (N_16745,N_16421,N_16489);
or U16746 (N_16746,N_16296,N_16421);
nand U16747 (N_16747,N_16370,N_16479);
nand U16748 (N_16748,N_16364,N_16475);
or U16749 (N_16749,N_16361,N_16465);
xnor U16750 (N_16750,N_16682,N_16737);
xor U16751 (N_16751,N_16647,N_16531);
xnor U16752 (N_16752,N_16590,N_16689);
or U16753 (N_16753,N_16518,N_16563);
xor U16754 (N_16754,N_16610,N_16627);
or U16755 (N_16755,N_16556,N_16738);
xnor U16756 (N_16756,N_16527,N_16658);
or U16757 (N_16757,N_16708,N_16637);
xor U16758 (N_16758,N_16500,N_16698);
or U16759 (N_16759,N_16670,N_16572);
or U16760 (N_16760,N_16690,N_16558);
xnor U16761 (N_16761,N_16722,N_16633);
and U16762 (N_16762,N_16528,N_16509);
nor U16763 (N_16763,N_16706,N_16697);
and U16764 (N_16764,N_16721,N_16602);
nand U16765 (N_16765,N_16606,N_16516);
xnor U16766 (N_16766,N_16517,N_16554);
xnor U16767 (N_16767,N_16648,N_16741);
or U16768 (N_16768,N_16545,N_16515);
nor U16769 (N_16769,N_16657,N_16594);
nor U16770 (N_16770,N_16629,N_16621);
and U16771 (N_16771,N_16560,N_16653);
or U16772 (N_16772,N_16506,N_16639);
or U16773 (N_16773,N_16593,N_16681);
nand U16774 (N_16774,N_16641,N_16605);
and U16775 (N_16775,N_16703,N_16587);
or U16776 (N_16776,N_16573,N_16619);
xor U16777 (N_16777,N_16732,N_16678);
nor U16778 (N_16778,N_16643,N_16581);
xnor U16779 (N_16779,N_16552,N_16588);
xor U16780 (N_16780,N_16569,N_16513);
or U16781 (N_16781,N_16592,N_16507);
xnor U16782 (N_16782,N_16720,N_16561);
or U16783 (N_16783,N_16622,N_16655);
xnor U16784 (N_16784,N_16532,N_16617);
xor U16785 (N_16785,N_16626,N_16656);
xor U16786 (N_16786,N_16747,N_16564);
or U16787 (N_16787,N_16618,N_16667);
xnor U16788 (N_16788,N_16715,N_16686);
or U16789 (N_16789,N_16623,N_16733);
nor U16790 (N_16790,N_16728,N_16677);
nor U16791 (N_16791,N_16505,N_16694);
nor U16792 (N_16792,N_16669,N_16688);
nand U16793 (N_16793,N_16702,N_16729);
and U16794 (N_16794,N_16589,N_16585);
or U16795 (N_16795,N_16540,N_16603);
nor U16796 (N_16796,N_16608,N_16710);
nand U16797 (N_16797,N_16601,N_16612);
and U16798 (N_16798,N_16744,N_16638);
nor U16799 (N_16799,N_16568,N_16665);
nor U16800 (N_16800,N_16685,N_16511);
and U16801 (N_16801,N_16575,N_16673);
and U16802 (N_16802,N_16695,N_16628);
or U16803 (N_16803,N_16544,N_16577);
and U16804 (N_16804,N_16548,N_16700);
or U16805 (N_16805,N_16514,N_16731);
nand U16806 (N_16806,N_16701,N_16550);
nand U16807 (N_16807,N_16562,N_16620);
and U16808 (N_16808,N_16671,N_16523);
and U16809 (N_16809,N_16662,N_16726);
and U16810 (N_16810,N_16539,N_16598);
nor U16811 (N_16811,N_16586,N_16565);
nand U16812 (N_16812,N_16557,N_16743);
nor U16813 (N_16813,N_16675,N_16680);
and U16814 (N_16814,N_16534,N_16616);
nor U16815 (N_16815,N_16745,N_16709);
nand U16816 (N_16816,N_16704,N_16659);
and U16817 (N_16817,N_16654,N_16674);
xor U16818 (N_16818,N_16696,N_16748);
nand U16819 (N_16819,N_16624,N_16734);
xnor U16820 (N_16820,N_16679,N_16526);
and U16821 (N_16821,N_16595,N_16566);
xnor U16822 (N_16822,N_16735,N_16555);
nor U16823 (N_16823,N_16636,N_16521);
and U16824 (N_16824,N_16645,N_16611);
nor U16825 (N_16825,N_16668,N_16630);
or U16826 (N_16826,N_16533,N_16672);
xnor U16827 (N_16827,N_16600,N_16583);
or U16828 (N_16828,N_16504,N_16553);
xnor U16829 (N_16829,N_16749,N_16683);
and U16830 (N_16830,N_16537,N_16512);
or U16831 (N_16831,N_16713,N_16651);
xor U16832 (N_16832,N_16525,N_16604);
nor U16833 (N_16833,N_16584,N_16520);
nand U16834 (N_16834,N_16736,N_16609);
xnor U16835 (N_16835,N_16541,N_16723);
nor U16836 (N_16836,N_16660,N_16615);
nand U16837 (N_16837,N_16714,N_16576);
or U16838 (N_16838,N_16663,N_16724);
nor U16839 (N_16839,N_16613,N_16591);
xnor U16840 (N_16840,N_16530,N_16502);
nor U16841 (N_16841,N_16538,N_16635);
or U16842 (N_16842,N_16640,N_16524);
nand U16843 (N_16843,N_16559,N_16634);
xor U16844 (N_16844,N_16644,N_16571);
or U16845 (N_16845,N_16543,N_16546);
nor U16846 (N_16846,N_16666,N_16535);
or U16847 (N_16847,N_16607,N_16632);
and U16848 (N_16848,N_16684,N_16578);
nand U16849 (N_16849,N_16661,N_16580);
nand U16850 (N_16850,N_16676,N_16508);
xor U16851 (N_16851,N_16707,N_16740);
nand U16852 (N_16852,N_16579,N_16650);
and U16853 (N_16853,N_16746,N_16742);
nand U16854 (N_16854,N_16716,N_16529);
xor U16855 (N_16855,N_16711,N_16717);
nand U16856 (N_16856,N_16705,N_16567);
nand U16857 (N_16857,N_16582,N_16719);
and U16858 (N_16858,N_16625,N_16739);
nor U16859 (N_16859,N_16692,N_16712);
xor U16860 (N_16860,N_16642,N_16503);
nor U16861 (N_16861,N_16501,N_16551);
or U16862 (N_16862,N_16631,N_16646);
xnor U16863 (N_16863,N_16718,N_16693);
nand U16864 (N_16864,N_16597,N_16510);
and U16865 (N_16865,N_16649,N_16664);
nand U16866 (N_16866,N_16730,N_16599);
xor U16867 (N_16867,N_16687,N_16547);
nor U16868 (N_16868,N_16699,N_16691);
and U16869 (N_16869,N_16519,N_16570);
nor U16870 (N_16870,N_16596,N_16574);
and U16871 (N_16871,N_16652,N_16536);
and U16872 (N_16872,N_16725,N_16727);
nand U16873 (N_16873,N_16542,N_16614);
xnor U16874 (N_16874,N_16549,N_16522);
and U16875 (N_16875,N_16707,N_16553);
xnor U16876 (N_16876,N_16727,N_16513);
nor U16877 (N_16877,N_16732,N_16715);
nand U16878 (N_16878,N_16528,N_16548);
or U16879 (N_16879,N_16635,N_16518);
nand U16880 (N_16880,N_16701,N_16706);
nand U16881 (N_16881,N_16526,N_16682);
xor U16882 (N_16882,N_16553,N_16509);
xnor U16883 (N_16883,N_16731,N_16632);
nor U16884 (N_16884,N_16507,N_16591);
nand U16885 (N_16885,N_16685,N_16714);
and U16886 (N_16886,N_16655,N_16528);
xor U16887 (N_16887,N_16520,N_16588);
or U16888 (N_16888,N_16653,N_16728);
xnor U16889 (N_16889,N_16559,N_16700);
xnor U16890 (N_16890,N_16612,N_16686);
and U16891 (N_16891,N_16707,N_16706);
xnor U16892 (N_16892,N_16718,N_16566);
or U16893 (N_16893,N_16632,N_16692);
nand U16894 (N_16894,N_16735,N_16581);
xor U16895 (N_16895,N_16727,N_16519);
and U16896 (N_16896,N_16712,N_16727);
or U16897 (N_16897,N_16522,N_16635);
nor U16898 (N_16898,N_16542,N_16738);
and U16899 (N_16899,N_16685,N_16524);
or U16900 (N_16900,N_16545,N_16680);
nand U16901 (N_16901,N_16675,N_16621);
and U16902 (N_16902,N_16668,N_16724);
or U16903 (N_16903,N_16735,N_16633);
or U16904 (N_16904,N_16625,N_16727);
nor U16905 (N_16905,N_16507,N_16679);
nand U16906 (N_16906,N_16625,N_16598);
or U16907 (N_16907,N_16530,N_16587);
xor U16908 (N_16908,N_16702,N_16565);
nand U16909 (N_16909,N_16705,N_16532);
nor U16910 (N_16910,N_16726,N_16746);
nor U16911 (N_16911,N_16636,N_16559);
and U16912 (N_16912,N_16632,N_16740);
nor U16913 (N_16913,N_16608,N_16548);
nand U16914 (N_16914,N_16657,N_16562);
nor U16915 (N_16915,N_16580,N_16543);
or U16916 (N_16916,N_16623,N_16567);
nor U16917 (N_16917,N_16563,N_16510);
xnor U16918 (N_16918,N_16686,N_16571);
nor U16919 (N_16919,N_16610,N_16520);
nor U16920 (N_16920,N_16515,N_16575);
or U16921 (N_16921,N_16679,N_16738);
xor U16922 (N_16922,N_16657,N_16746);
nand U16923 (N_16923,N_16573,N_16533);
xnor U16924 (N_16924,N_16669,N_16513);
xor U16925 (N_16925,N_16549,N_16733);
xor U16926 (N_16926,N_16536,N_16712);
nor U16927 (N_16927,N_16688,N_16746);
nor U16928 (N_16928,N_16551,N_16744);
xnor U16929 (N_16929,N_16596,N_16655);
nor U16930 (N_16930,N_16570,N_16549);
xor U16931 (N_16931,N_16658,N_16503);
and U16932 (N_16932,N_16669,N_16654);
or U16933 (N_16933,N_16530,N_16548);
nor U16934 (N_16934,N_16519,N_16704);
nor U16935 (N_16935,N_16649,N_16545);
nor U16936 (N_16936,N_16505,N_16597);
nor U16937 (N_16937,N_16638,N_16531);
and U16938 (N_16938,N_16710,N_16574);
xor U16939 (N_16939,N_16685,N_16600);
nor U16940 (N_16940,N_16642,N_16628);
and U16941 (N_16941,N_16722,N_16564);
xnor U16942 (N_16942,N_16613,N_16565);
xor U16943 (N_16943,N_16575,N_16603);
nand U16944 (N_16944,N_16720,N_16738);
or U16945 (N_16945,N_16660,N_16534);
xnor U16946 (N_16946,N_16569,N_16521);
or U16947 (N_16947,N_16738,N_16739);
or U16948 (N_16948,N_16585,N_16668);
xnor U16949 (N_16949,N_16531,N_16708);
or U16950 (N_16950,N_16534,N_16608);
or U16951 (N_16951,N_16544,N_16519);
xnor U16952 (N_16952,N_16532,N_16606);
and U16953 (N_16953,N_16738,N_16570);
and U16954 (N_16954,N_16500,N_16512);
or U16955 (N_16955,N_16594,N_16743);
xor U16956 (N_16956,N_16713,N_16578);
nand U16957 (N_16957,N_16743,N_16739);
and U16958 (N_16958,N_16595,N_16527);
nor U16959 (N_16959,N_16618,N_16670);
nand U16960 (N_16960,N_16630,N_16734);
nor U16961 (N_16961,N_16742,N_16618);
and U16962 (N_16962,N_16680,N_16718);
and U16963 (N_16963,N_16748,N_16544);
or U16964 (N_16964,N_16512,N_16646);
nor U16965 (N_16965,N_16707,N_16579);
xor U16966 (N_16966,N_16651,N_16643);
nand U16967 (N_16967,N_16698,N_16511);
nand U16968 (N_16968,N_16619,N_16598);
xnor U16969 (N_16969,N_16652,N_16701);
nor U16970 (N_16970,N_16703,N_16720);
xor U16971 (N_16971,N_16551,N_16519);
or U16972 (N_16972,N_16626,N_16645);
nor U16973 (N_16973,N_16651,N_16500);
xor U16974 (N_16974,N_16684,N_16547);
xor U16975 (N_16975,N_16691,N_16594);
xor U16976 (N_16976,N_16629,N_16545);
and U16977 (N_16977,N_16501,N_16723);
nor U16978 (N_16978,N_16547,N_16659);
or U16979 (N_16979,N_16530,N_16737);
or U16980 (N_16980,N_16536,N_16545);
nand U16981 (N_16981,N_16632,N_16701);
and U16982 (N_16982,N_16524,N_16714);
nor U16983 (N_16983,N_16655,N_16660);
and U16984 (N_16984,N_16610,N_16592);
nand U16985 (N_16985,N_16742,N_16516);
xor U16986 (N_16986,N_16599,N_16674);
nor U16987 (N_16987,N_16634,N_16670);
and U16988 (N_16988,N_16712,N_16608);
nand U16989 (N_16989,N_16704,N_16646);
and U16990 (N_16990,N_16695,N_16713);
and U16991 (N_16991,N_16527,N_16744);
or U16992 (N_16992,N_16715,N_16565);
and U16993 (N_16993,N_16522,N_16515);
nand U16994 (N_16994,N_16669,N_16711);
or U16995 (N_16995,N_16560,N_16727);
nor U16996 (N_16996,N_16528,N_16570);
and U16997 (N_16997,N_16599,N_16611);
or U16998 (N_16998,N_16551,N_16578);
and U16999 (N_16999,N_16585,N_16587);
nor U17000 (N_17000,N_16952,N_16812);
and U17001 (N_17001,N_16754,N_16924);
or U17002 (N_17002,N_16753,N_16811);
nor U17003 (N_17003,N_16760,N_16759);
or U17004 (N_17004,N_16987,N_16884);
and U17005 (N_17005,N_16932,N_16938);
or U17006 (N_17006,N_16757,N_16794);
xor U17007 (N_17007,N_16756,N_16770);
and U17008 (N_17008,N_16970,N_16935);
or U17009 (N_17009,N_16795,N_16777);
and U17010 (N_17010,N_16804,N_16984);
nor U17011 (N_17011,N_16820,N_16921);
xor U17012 (N_17012,N_16983,N_16990);
or U17013 (N_17013,N_16805,N_16891);
xnor U17014 (N_17014,N_16871,N_16818);
nand U17015 (N_17015,N_16946,N_16807);
nand U17016 (N_17016,N_16962,N_16918);
or U17017 (N_17017,N_16815,N_16890);
or U17018 (N_17018,N_16874,N_16919);
nand U17019 (N_17019,N_16776,N_16982);
nand U17020 (N_17020,N_16904,N_16894);
and U17021 (N_17021,N_16929,N_16862);
nor U17022 (N_17022,N_16945,N_16841);
and U17023 (N_17023,N_16901,N_16974);
nor U17024 (N_17024,N_16802,N_16986);
nand U17025 (N_17025,N_16917,N_16792);
nor U17026 (N_17026,N_16840,N_16790);
nor U17027 (N_17027,N_16806,N_16902);
nor U17028 (N_17028,N_16782,N_16893);
or U17029 (N_17029,N_16796,N_16784);
and U17030 (N_17030,N_16980,N_16922);
xor U17031 (N_17031,N_16763,N_16783);
nor U17032 (N_17032,N_16819,N_16781);
xnor U17033 (N_17033,N_16766,N_16858);
or U17034 (N_17034,N_16772,N_16857);
nor U17035 (N_17035,N_16875,N_16839);
nand U17036 (N_17036,N_16971,N_16863);
or U17037 (N_17037,N_16798,N_16752);
nand U17038 (N_17038,N_16957,N_16856);
and U17039 (N_17039,N_16954,N_16851);
nor U17040 (N_17040,N_16955,N_16979);
or U17041 (N_17041,N_16934,N_16859);
xnor U17042 (N_17042,N_16750,N_16809);
or U17043 (N_17043,N_16906,N_16849);
xor U17044 (N_17044,N_16976,N_16799);
nand U17045 (N_17045,N_16883,N_16900);
nand U17046 (N_17046,N_16992,N_16993);
or U17047 (N_17047,N_16847,N_16880);
and U17048 (N_17048,N_16865,N_16771);
nor U17049 (N_17049,N_16755,N_16899);
xor U17050 (N_17050,N_16835,N_16953);
xnor U17051 (N_17051,N_16867,N_16967);
and U17052 (N_17052,N_16853,N_16872);
and U17053 (N_17053,N_16780,N_16787);
xor U17054 (N_17054,N_16824,N_16758);
nor U17055 (N_17055,N_16948,N_16958);
nor U17056 (N_17056,N_16868,N_16977);
nand U17057 (N_17057,N_16789,N_16791);
nor U17058 (N_17058,N_16827,N_16965);
xor U17059 (N_17059,N_16870,N_16836);
and U17060 (N_17060,N_16936,N_16838);
nand U17061 (N_17061,N_16779,N_16844);
or U17062 (N_17062,N_16930,N_16828);
nand U17063 (N_17063,N_16774,N_16920);
nand U17064 (N_17064,N_16832,N_16994);
nor U17065 (N_17065,N_16928,N_16778);
nor U17066 (N_17066,N_16769,N_16843);
and U17067 (N_17067,N_16816,N_16751);
xor U17068 (N_17068,N_16941,N_16773);
or U17069 (N_17069,N_16999,N_16950);
nor U17070 (N_17070,N_16991,N_16956);
nor U17071 (N_17071,N_16972,N_16923);
nand U17072 (N_17072,N_16892,N_16940);
xor U17073 (N_17073,N_16925,N_16885);
xor U17074 (N_17074,N_16997,N_16960);
and U17075 (N_17075,N_16937,N_16852);
xor U17076 (N_17076,N_16810,N_16912);
or U17077 (N_17077,N_16842,N_16829);
xor U17078 (N_17078,N_16886,N_16927);
or U17079 (N_17079,N_16998,N_16989);
nand U17080 (N_17080,N_16985,N_16854);
nand U17081 (N_17081,N_16830,N_16931);
or U17082 (N_17082,N_16968,N_16889);
and U17083 (N_17083,N_16887,N_16995);
nand U17084 (N_17084,N_16939,N_16978);
nand U17085 (N_17085,N_16966,N_16821);
or U17086 (N_17086,N_16882,N_16833);
nor U17087 (N_17087,N_16813,N_16848);
xor U17088 (N_17088,N_16866,N_16808);
or U17089 (N_17089,N_16762,N_16944);
nand U17090 (N_17090,N_16873,N_16926);
and U17091 (N_17091,N_16896,N_16767);
nand U17092 (N_17092,N_16814,N_16909);
xor U17093 (N_17093,N_16911,N_16914);
and U17094 (N_17094,N_16803,N_16895);
nor U17095 (N_17095,N_16969,N_16786);
xor U17096 (N_17096,N_16765,N_16975);
nor U17097 (N_17097,N_16988,N_16837);
nor U17098 (N_17098,N_16761,N_16823);
nor U17099 (N_17099,N_16801,N_16996);
nor U17100 (N_17100,N_16916,N_16826);
or U17101 (N_17101,N_16905,N_16961);
or U17102 (N_17102,N_16973,N_16959);
nand U17103 (N_17103,N_16933,N_16764);
nor U17104 (N_17104,N_16915,N_16860);
nor U17105 (N_17105,N_16788,N_16817);
and U17106 (N_17106,N_16768,N_16864);
nor U17107 (N_17107,N_16850,N_16878);
xnor U17108 (N_17108,N_16881,N_16845);
xor U17109 (N_17109,N_16793,N_16981);
or U17110 (N_17110,N_16910,N_16907);
or U17111 (N_17111,N_16951,N_16879);
or U17112 (N_17112,N_16855,N_16831);
nor U17113 (N_17113,N_16897,N_16775);
xnor U17114 (N_17114,N_16947,N_16834);
and U17115 (N_17115,N_16908,N_16800);
xor U17116 (N_17116,N_16822,N_16913);
nand U17117 (N_17117,N_16876,N_16942);
or U17118 (N_17118,N_16785,N_16898);
or U17119 (N_17119,N_16943,N_16846);
nand U17120 (N_17120,N_16825,N_16888);
nor U17121 (N_17121,N_16869,N_16903);
nand U17122 (N_17122,N_16949,N_16963);
nand U17123 (N_17123,N_16797,N_16861);
and U17124 (N_17124,N_16877,N_16964);
and U17125 (N_17125,N_16826,N_16932);
and U17126 (N_17126,N_16926,N_16877);
or U17127 (N_17127,N_16969,N_16847);
xor U17128 (N_17128,N_16956,N_16845);
nor U17129 (N_17129,N_16914,N_16859);
and U17130 (N_17130,N_16802,N_16932);
or U17131 (N_17131,N_16856,N_16795);
xnor U17132 (N_17132,N_16890,N_16807);
and U17133 (N_17133,N_16765,N_16901);
nor U17134 (N_17134,N_16839,N_16970);
or U17135 (N_17135,N_16760,N_16812);
nand U17136 (N_17136,N_16940,N_16797);
nor U17137 (N_17137,N_16815,N_16814);
and U17138 (N_17138,N_16757,N_16927);
nand U17139 (N_17139,N_16838,N_16998);
and U17140 (N_17140,N_16877,N_16912);
or U17141 (N_17141,N_16984,N_16845);
or U17142 (N_17142,N_16987,N_16919);
or U17143 (N_17143,N_16984,N_16862);
and U17144 (N_17144,N_16867,N_16991);
xor U17145 (N_17145,N_16870,N_16758);
or U17146 (N_17146,N_16989,N_16912);
and U17147 (N_17147,N_16873,N_16918);
or U17148 (N_17148,N_16834,N_16815);
nand U17149 (N_17149,N_16831,N_16784);
xor U17150 (N_17150,N_16872,N_16866);
nor U17151 (N_17151,N_16788,N_16779);
or U17152 (N_17152,N_16818,N_16909);
or U17153 (N_17153,N_16861,N_16859);
xnor U17154 (N_17154,N_16967,N_16802);
xor U17155 (N_17155,N_16962,N_16968);
nand U17156 (N_17156,N_16799,N_16825);
xnor U17157 (N_17157,N_16789,N_16857);
or U17158 (N_17158,N_16995,N_16914);
and U17159 (N_17159,N_16776,N_16775);
and U17160 (N_17160,N_16862,N_16754);
or U17161 (N_17161,N_16926,N_16927);
or U17162 (N_17162,N_16837,N_16846);
nor U17163 (N_17163,N_16897,N_16981);
nor U17164 (N_17164,N_16894,N_16832);
nor U17165 (N_17165,N_16923,N_16909);
nand U17166 (N_17166,N_16772,N_16927);
nand U17167 (N_17167,N_16786,N_16964);
or U17168 (N_17168,N_16877,N_16884);
nand U17169 (N_17169,N_16754,N_16968);
xnor U17170 (N_17170,N_16949,N_16931);
or U17171 (N_17171,N_16846,N_16933);
and U17172 (N_17172,N_16942,N_16924);
nor U17173 (N_17173,N_16993,N_16785);
and U17174 (N_17174,N_16943,N_16823);
nand U17175 (N_17175,N_16916,N_16966);
nor U17176 (N_17176,N_16972,N_16988);
xor U17177 (N_17177,N_16834,N_16812);
and U17178 (N_17178,N_16885,N_16820);
nor U17179 (N_17179,N_16818,N_16907);
nand U17180 (N_17180,N_16826,N_16792);
or U17181 (N_17181,N_16750,N_16998);
or U17182 (N_17182,N_16810,N_16965);
or U17183 (N_17183,N_16891,N_16832);
or U17184 (N_17184,N_16973,N_16993);
and U17185 (N_17185,N_16985,N_16870);
and U17186 (N_17186,N_16778,N_16957);
nand U17187 (N_17187,N_16807,N_16881);
xor U17188 (N_17188,N_16839,N_16770);
nand U17189 (N_17189,N_16751,N_16766);
nor U17190 (N_17190,N_16996,N_16953);
and U17191 (N_17191,N_16764,N_16863);
and U17192 (N_17192,N_16917,N_16808);
nand U17193 (N_17193,N_16779,N_16928);
xor U17194 (N_17194,N_16984,N_16931);
and U17195 (N_17195,N_16832,N_16834);
or U17196 (N_17196,N_16931,N_16973);
or U17197 (N_17197,N_16881,N_16764);
xor U17198 (N_17198,N_16928,N_16984);
nor U17199 (N_17199,N_16804,N_16776);
and U17200 (N_17200,N_16767,N_16917);
nand U17201 (N_17201,N_16984,N_16958);
nand U17202 (N_17202,N_16972,N_16940);
nor U17203 (N_17203,N_16815,N_16842);
nand U17204 (N_17204,N_16819,N_16876);
xnor U17205 (N_17205,N_16799,N_16772);
xor U17206 (N_17206,N_16886,N_16815);
and U17207 (N_17207,N_16989,N_16949);
nand U17208 (N_17208,N_16807,N_16935);
or U17209 (N_17209,N_16893,N_16910);
and U17210 (N_17210,N_16865,N_16943);
and U17211 (N_17211,N_16949,N_16788);
xor U17212 (N_17212,N_16910,N_16835);
and U17213 (N_17213,N_16840,N_16938);
nor U17214 (N_17214,N_16981,N_16972);
and U17215 (N_17215,N_16904,N_16944);
nor U17216 (N_17216,N_16955,N_16947);
nand U17217 (N_17217,N_16858,N_16898);
xnor U17218 (N_17218,N_16897,N_16886);
and U17219 (N_17219,N_16919,N_16822);
and U17220 (N_17220,N_16795,N_16940);
nor U17221 (N_17221,N_16941,N_16906);
xnor U17222 (N_17222,N_16877,N_16854);
or U17223 (N_17223,N_16853,N_16969);
nor U17224 (N_17224,N_16949,N_16972);
and U17225 (N_17225,N_16813,N_16971);
nand U17226 (N_17226,N_16823,N_16830);
or U17227 (N_17227,N_16812,N_16808);
nor U17228 (N_17228,N_16926,N_16841);
xnor U17229 (N_17229,N_16946,N_16804);
and U17230 (N_17230,N_16760,N_16888);
and U17231 (N_17231,N_16789,N_16801);
and U17232 (N_17232,N_16873,N_16854);
and U17233 (N_17233,N_16766,N_16925);
or U17234 (N_17234,N_16832,N_16933);
nand U17235 (N_17235,N_16885,N_16824);
nor U17236 (N_17236,N_16843,N_16793);
nand U17237 (N_17237,N_16779,N_16948);
xor U17238 (N_17238,N_16919,N_16979);
nor U17239 (N_17239,N_16990,N_16936);
and U17240 (N_17240,N_16960,N_16872);
or U17241 (N_17241,N_16967,N_16943);
xor U17242 (N_17242,N_16777,N_16753);
and U17243 (N_17243,N_16803,N_16766);
or U17244 (N_17244,N_16886,N_16768);
and U17245 (N_17245,N_16812,N_16782);
xor U17246 (N_17246,N_16855,N_16760);
nor U17247 (N_17247,N_16837,N_16818);
xor U17248 (N_17248,N_16778,N_16767);
and U17249 (N_17249,N_16822,N_16786);
and U17250 (N_17250,N_17044,N_17097);
xor U17251 (N_17251,N_17100,N_17043);
xor U17252 (N_17252,N_17048,N_17211);
and U17253 (N_17253,N_17248,N_17012);
nand U17254 (N_17254,N_17239,N_17139);
nand U17255 (N_17255,N_17172,N_17050);
nor U17256 (N_17256,N_17168,N_17030);
nand U17257 (N_17257,N_17124,N_17166);
and U17258 (N_17258,N_17042,N_17242);
xnor U17259 (N_17259,N_17001,N_17197);
nand U17260 (N_17260,N_17026,N_17105);
or U17261 (N_17261,N_17108,N_17155);
and U17262 (N_17262,N_17249,N_17020);
or U17263 (N_17263,N_17226,N_17063);
and U17264 (N_17264,N_17013,N_17143);
or U17265 (N_17265,N_17083,N_17223);
xnor U17266 (N_17266,N_17192,N_17060);
or U17267 (N_17267,N_17099,N_17126);
xnor U17268 (N_17268,N_17089,N_17128);
or U17269 (N_17269,N_17092,N_17245);
xor U17270 (N_17270,N_17146,N_17008);
or U17271 (N_17271,N_17036,N_17062);
nor U17272 (N_17272,N_17070,N_17171);
or U17273 (N_17273,N_17104,N_17164);
xnor U17274 (N_17274,N_17022,N_17232);
or U17275 (N_17275,N_17169,N_17150);
xnor U17276 (N_17276,N_17210,N_17002);
nand U17277 (N_17277,N_17194,N_17034);
xnor U17278 (N_17278,N_17113,N_17198);
nand U17279 (N_17279,N_17084,N_17080);
nor U17280 (N_17280,N_17233,N_17147);
nor U17281 (N_17281,N_17118,N_17010);
xnor U17282 (N_17282,N_17090,N_17195);
nand U17283 (N_17283,N_17074,N_17185);
nor U17284 (N_17284,N_17246,N_17240);
and U17285 (N_17285,N_17173,N_17047);
nor U17286 (N_17286,N_17186,N_17072);
or U17287 (N_17287,N_17157,N_17087);
nand U17288 (N_17288,N_17029,N_17017);
nor U17289 (N_17289,N_17170,N_17051);
or U17290 (N_17290,N_17193,N_17218);
or U17291 (N_17291,N_17156,N_17243);
nand U17292 (N_17292,N_17069,N_17144);
and U17293 (N_17293,N_17085,N_17160);
nand U17294 (N_17294,N_17183,N_17054);
and U17295 (N_17295,N_17141,N_17111);
or U17296 (N_17296,N_17096,N_17041);
and U17297 (N_17297,N_17123,N_17209);
xnor U17298 (N_17298,N_17163,N_17122);
or U17299 (N_17299,N_17015,N_17021);
xor U17300 (N_17300,N_17009,N_17102);
xnor U17301 (N_17301,N_17007,N_17101);
and U17302 (N_17302,N_17154,N_17119);
xnor U17303 (N_17303,N_17133,N_17247);
xnor U17304 (N_17304,N_17236,N_17035);
and U17305 (N_17305,N_17130,N_17215);
nor U17306 (N_17306,N_17153,N_17094);
or U17307 (N_17307,N_17073,N_17220);
nand U17308 (N_17308,N_17049,N_17027);
nor U17309 (N_17309,N_17106,N_17206);
or U17310 (N_17310,N_17179,N_17158);
or U17311 (N_17311,N_17114,N_17011);
xnor U17312 (N_17312,N_17037,N_17018);
and U17313 (N_17313,N_17225,N_17212);
or U17314 (N_17314,N_17071,N_17189);
xor U17315 (N_17315,N_17109,N_17076);
xor U17316 (N_17316,N_17196,N_17159);
nor U17317 (N_17317,N_17187,N_17107);
nand U17318 (N_17318,N_17019,N_17091);
and U17319 (N_17319,N_17142,N_17213);
nand U17320 (N_17320,N_17135,N_17238);
nand U17321 (N_17321,N_17059,N_17184);
nand U17322 (N_17322,N_17165,N_17006);
and U17323 (N_17323,N_17204,N_17134);
nand U17324 (N_17324,N_17103,N_17237);
xor U17325 (N_17325,N_17057,N_17003);
or U17326 (N_17326,N_17038,N_17161);
nor U17327 (N_17327,N_17132,N_17061);
xnor U17328 (N_17328,N_17167,N_17046);
nand U17329 (N_17329,N_17053,N_17202);
xor U17330 (N_17330,N_17031,N_17177);
xnor U17331 (N_17331,N_17228,N_17203);
xor U17332 (N_17332,N_17088,N_17222);
or U17333 (N_17333,N_17199,N_17244);
nor U17334 (N_17334,N_17033,N_17188);
or U17335 (N_17335,N_17040,N_17205);
and U17336 (N_17336,N_17200,N_17140);
xnor U17337 (N_17337,N_17058,N_17067);
and U17338 (N_17338,N_17235,N_17023);
nor U17339 (N_17339,N_17208,N_17162);
nor U17340 (N_17340,N_17241,N_17191);
or U17341 (N_17341,N_17078,N_17115);
and U17342 (N_17342,N_17217,N_17056);
or U17343 (N_17343,N_17224,N_17148);
and U17344 (N_17344,N_17175,N_17025);
or U17345 (N_17345,N_17221,N_17068);
xor U17346 (N_17346,N_17112,N_17230);
xor U17347 (N_17347,N_17137,N_17231);
xor U17348 (N_17348,N_17064,N_17181);
nor U17349 (N_17349,N_17229,N_17045);
and U17350 (N_17350,N_17075,N_17086);
nand U17351 (N_17351,N_17000,N_17121);
xor U17352 (N_17352,N_17093,N_17120);
nor U17353 (N_17353,N_17201,N_17065);
and U17354 (N_17354,N_17176,N_17117);
nor U17355 (N_17355,N_17174,N_17190);
and U17356 (N_17356,N_17028,N_17219);
or U17357 (N_17357,N_17145,N_17095);
or U17358 (N_17358,N_17138,N_17180);
or U17359 (N_17359,N_17024,N_17005);
and U17360 (N_17360,N_17016,N_17178);
and U17361 (N_17361,N_17077,N_17136);
and U17362 (N_17362,N_17149,N_17039);
nand U17363 (N_17363,N_17098,N_17004);
xor U17364 (N_17364,N_17227,N_17079);
nor U17365 (N_17365,N_17129,N_17127);
or U17366 (N_17366,N_17207,N_17066);
and U17367 (N_17367,N_17234,N_17152);
nand U17368 (N_17368,N_17014,N_17131);
nor U17369 (N_17369,N_17125,N_17082);
nand U17370 (N_17370,N_17214,N_17055);
xor U17371 (N_17371,N_17151,N_17182);
or U17372 (N_17372,N_17110,N_17116);
and U17373 (N_17373,N_17081,N_17032);
nand U17374 (N_17374,N_17052,N_17216);
or U17375 (N_17375,N_17019,N_17186);
and U17376 (N_17376,N_17165,N_17114);
nand U17377 (N_17377,N_17120,N_17000);
or U17378 (N_17378,N_17177,N_17149);
nor U17379 (N_17379,N_17084,N_17112);
nor U17380 (N_17380,N_17153,N_17029);
nand U17381 (N_17381,N_17215,N_17072);
and U17382 (N_17382,N_17151,N_17200);
xor U17383 (N_17383,N_17121,N_17226);
nor U17384 (N_17384,N_17026,N_17111);
nor U17385 (N_17385,N_17186,N_17090);
xnor U17386 (N_17386,N_17240,N_17245);
and U17387 (N_17387,N_17044,N_17160);
or U17388 (N_17388,N_17194,N_17109);
nor U17389 (N_17389,N_17012,N_17071);
nor U17390 (N_17390,N_17188,N_17110);
xnor U17391 (N_17391,N_17214,N_17016);
or U17392 (N_17392,N_17078,N_17042);
nor U17393 (N_17393,N_17009,N_17061);
nand U17394 (N_17394,N_17161,N_17072);
xor U17395 (N_17395,N_17149,N_17170);
nor U17396 (N_17396,N_17114,N_17236);
and U17397 (N_17397,N_17241,N_17129);
nor U17398 (N_17398,N_17003,N_17114);
xnor U17399 (N_17399,N_17186,N_17160);
xor U17400 (N_17400,N_17162,N_17041);
xor U17401 (N_17401,N_17123,N_17227);
nand U17402 (N_17402,N_17230,N_17156);
and U17403 (N_17403,N_17228,N_17166);
nor U17404 (N_17404,N_17101,N_17105);
or U17405 (N_17405,N_17136,N_17133);
or U17406 (N_17406,N_17003,N_17036);
xor U17407 (N_17407,N_17238,N_17242);
nor U17408 (N_17408,N_17099,N_17115);
or U17409 (N_17409,N_17103,N_17092);
and U17410 (N_17410,N_17186,N_17022);
or U17411 (N_17411,N_17194,N_17214);
or U17412 (N_17412,N_17138,N_17079);
or U17413 (N_17413,N_17034,N_17126);
xor U17414 (N_17414,N_17175,N_17218);
nand U17415 (N_17415,N_17053,N_17167);
nand U17416 (N_17416,N_17198,N_17191);
nor U17417 (N_17417,N_17130,N_17061);
nand U17418 (N_17418,N_17212,N_17106);
nor U17419 (N_17419,N_17183,N_17159);
or U17420 (N_17420,N_17177,N_17087);
nor U17421 (N_17421,N_17126,N_17238);
nor U17422 (N_17422,N_17235,N_17009);
nand U17423 (N_17423,N_17185,N_17060);
nor U17424 (N_17424,N_17169,N_17125);
nor U17425 (N_17425,N_17054,N_17035);
nand U17426 (N_17426,N_17233,N_17057);
nor U17427 (N_17427,N_17099,N_17133);
nor U17428 (N_17428,N_17197,N_17151);
xnor U17429 (N_17429,N_17242,N_17231);
or U17430 (N_17430,N_17142,N_17191);
and U17431 (N_17431,N_17075,N_17221);
or U17432 (N_17432,N_17074,N_17057);
xnor U17433 (N_17433,N_17056,N_17097);
xnor U17434 (N_17434,N_17132,N_17017);
nand U17435 (N_17435,N_17193,N_17081);
nor U17436 (N_17436,N_17031,N_17095);
and U17437 (N_17437,N_17196,N_17009);
nor U17438 (N_17438,N_17044,N_17231);
and U17439 (N_17439,N_17063,N_17085);
and U17440 (N_17440,N_17135,N_17145);
nor U17441 (N_17441,N_17108,N_17012);
nand U17442 (N_17442,N_17235,N_17006);
xor U17443 (N_17443,N_17021,N_17198);
and U17444 (N_17444,N_17134,N_17005);
nor U17445 (N_17445,N_17058,N_17174);
or U17446 (N_17446,N_17037,N_17080);
xnor U17447 (N_17447,N_17082,N_17109);
or U17448 (N_17448,N_17143,N_17115);
and U17449 (N_17449,N_17203,N_17224);
xor U17450 (N_17450,N_17177,N_17174);
nor U17451 (N_17451,N_17114,N_17082);
and U17452 (N_17452,N_17020,N_17036);
nand U17453 (N_17453,N_17173,N_17006);
xnor U17454 (N_17454,N_17183,N_17150);
and U17455 (N_17455,N_17193,N_17129);
or U17456 (N_17456,N_17022,N_17062);
nor U17457 (N_17457,N_17005,N_17128);
or U17458 (N_17458,N_17113,N_17083);
nor U17459 (N_17459,N_17178,N_17234);
nor U17460 (N_17460,N_17021,N_17105);
nor U17461 (N_17461,N_17030,N_17236);
xnor U17462 (N_17462,N_17037,N_17009);
nand U17463 (N_17463,N_17188,N_17196);
nand U17464 (N_17464,N_17000,N_17192);
nand U17465 (N_17465,N_17198,N_17112);
and U17466 (N_17466,N_17184,N_17149);
nor U17467 (N_17467,N_17174,N_17134);
or U17468 (N_17468,N_17209,N_17158);
xnor U17469 (N_17469,N_17036,N_17052);
or U17470 (N_17470,N_17143,N_17006);
or U17471 (N_17471,N_17012,N_17162);
and U17472 (N_17472,N_17084,N_17179);
xor U17473 (N_17473,N_17051,N_17202);
or U17474 (N_17474,N_17117,N_17228);
and U17475 (N_17475,N_17050,N_17175);
or U17476 (N_17476,N_17158,N_17208);
and U17477 (N_17477,N_17010,N_17237);
nand U17478 (N_17478,N_17000,N_17143);
nand U17479 (N_17479,N_17118,N_17083);
nand U17480 (N_17480,N_17146,N_17248);
or U17481 (N_17481,N_17084,N_17215);
nor U17482 (N_17482,N_17105,N_17188);
nand U17483 (N_17483,N_17138,N_17122);
xor U17484 (N_17484,N_17223,N_17015);
nand U17485 (N_17485,N_17093,N_17209);
or U17486 (N_17486,N_17053,N_17035);
xor U17487 (N_17487,N_17163,N_17010);
or U17488 (N_17488,N_17054,N_17064);
or U17489 (N_17489,N_17171,N_17000);
xnor U17490 (N_17490,N_17162,N_17001);
nand U17491 (N_17491,N_17239,N_17054);
nor U17492 (N_17492,N_17033,N_17035);
or U17493 (N_17493,N_17002,N_17044);
nor U17494 (N_17494,N_17206,N_17226);
nor U17495 (N_17495,N_17094,N_17174);
nor U17496 (N_17496,N_17036,N_17035);
nor U17497 (N_17497,N_17190,N_17069);
or U17498 (N_17498,N_17158,N_17165);
xnor U17499 (N_17499,N_17242,N_17033);
nand U17500 (N_17500,N_17352,N_17440);
or U17501 (N_17501,N_17483,N_17273);
nand U17502 (N_17502,N_17299,N_17328);
or U17503 (N_17503,N_17388,N_17366);
nor U17504 (N_17504,N_17356,N_17472);
and U17505 (N_17505,N_17396,N_17331);
xor U17506 (N_17506,N_17435,N_17494);
xnor U17507 (N_17507,N_17432,N_17278);
or U17508 (N_17508,N_17397,N_17363);
xor U17509 (N_17509,N_17270,N_17297);
or U17510 (N_17510,N_17377,N_17464);
and U17511 (N_17511,N_17284,N_17251);
nor U17512 (N_17512,N_17332,N_17371);
or U17513 (N_17513,N_17376,N_17365);
nand U17514 (N_17514,N_17350,N_17436);
or U17515 (N_17515,N_17475,N_17311);
nand U17516 (N_17516,N_17468,N_17323);
nand U17517 (N_17517,N_17335,N_17391);
nand U17518 (N_17518,N_17266,N_17459);
nand U17519 (N_17519,N_17439,N_17267);
or U17520 (N_17520,N_17380,N_17361);
nor U17521 (N_17521,N_17362,N_17470);
xor U17522 (N_17522,N_17334,N_17455);
nor U17523 (N_17523,N_17408,N_17423);
nor U17524 (N_17524,N_17340,N_17256);
xor U17525 (N_17525,N_17449,N_17451);
or U17526 (N_17526,N_17281,N_17422);
nor U17527 (N_17527,N_17419,N_17447);
xnor U17528 (N_17528,N_17466,N_17289);
and U17529 (N_17529,N_17326,N_17387);
xnor U17530 (N_17530,N_17305,N_17402);
nor U17531 (N_17531,N_17330,N_17292);
xnor U17532 (N_17532,N_17403,N_17275);
nor U17533 (N_17533,N_17320,N_17401);
xnor U17534 (N_17534,N_17265,N_17486);
and U17535 (N_17535,N_17429,N_17287);
nand U17536 (N_17536,N_17476,N_17347);
nor U17537 (N_17537,N_17339,N_17382);
nand U17538 (N_17538,N_17279,N_17498);
or U17539 (N_17539,N_17469,N_17414);
nor U17540 (N_17540,N_17488,N_17303);
nor U17541 (N_17541,N_17316,N_17379);
nor U17542 (N_17542,N_17445,N_17345);
or U17543 (N_17543,N_17282,N_17415);
nand U17544 (N_17544,N_17269,N_17487);
xor U17545 (N_17545,N_17395,N_17253);
nand U17546 (N_17546,N_17479,N_17437);
and U17547 (N_17547,N_17369,N_17288);
xnor U17548 (N_17548,N_17480,N_17342);
nor U17549 (N_17549,N_17489,N_17460);
nand U17550 (N_17550,N_17400,N_17322);
nand U17551 (N_17551,N_17291,N_17448);
and U17552 (N_17552,N_17338,N_17484);
nor U17553 (N_17553,N_17306,N_17497);
or U17554 (N_17554,N_17370,N_17444);
nand U17555 (N_17555,N_17280,N_17274);
nor U17556 (N_17556,N_17478,N_17321);
or U17557 (N_17557,N_17485,N_17420);
or U17558 (N_17558,N_17416,N_17304);
or U17559 (N_17559,N_17375,N_17433);
and U17560 (N_17560,N_17329,N_17394);
xnor U17561 (N_17561,N_17294,N_17398);
and U17562 (N_17562,N_17424,N_17268);
nand U17563 (N_17563,N_17337,N_17277);
xnor U17564 (N_17564,N_17264,N_17404);
and U17565 (N_17565,N_17298,N_17290);
and U17566 (N_17566,N_17271,N_17384);
nor U17567 (N_17567,N_17427,N_17250);
xor U17568 (N_17568,N_17430,N_17410);
or U17569 (N_17569,N_17390,N_17252);
xor U17570 (N_17570,N_17428,N_17411);
or U17571 (N_17571,N_17367,N_17358);
or U17572 (N_17572,N_17481,N_17255);
nand U17573 (N_17573,N_17496,N_17454);
nor U17574 (N_17574,N_17319,N_17354);
nand U17575 (N_17575,N_17386,N_17450);
nor U17576 (N_17576,N_17359,N_17431);
xor U17577 (N_17577,N_17452,N_17308);
or U17578 (N_17578,N_17353,N_17467);
and U17579 (N_17579,N_17457,N_17344);
nand U17580 (N_17580,N_17442,N_17399);
nand U17581 (N_17581,N_17262,N_17458);
nor U17582 (N_17582,N_17407,N_17461);
and U17583 (N_17583,N_17381,N_17336);
nor U17584 (N_17584,N_17315,N_17364);
xnor U17585 (N_17585,N_17272,N_17492);
and U17586 (N_17586,N_17453,N_17409);
nand U17587 (N_17587,N_17283,N_17434);
nor U17588 (N_17588,N_17499,N_17446);
or U17589 (N_17589,N_17441,N_17293);
or U17590 (N_17590,N_17327,N_17261);
or U17591 (N_17591,N_17301,N_17417);
nor U17592 (N_17592,N_17257,N_17413);
xnor U17593 (N_17593,N_17285,N_17490);
nor U17594 (N_17594,N_17438,N_17351);
xor U17595 (N_17595,N_17405,N_17260);
or U17596 (N_17596,N_17296,N_17312);
nor U17597 (N_17597,N_17421,N_17286);
or U17598 (N_17598,N_17463,N_17462);
nor U17599 (N_17599,N_17374,N_17300);
xor U17600 (N_17600,N_17426,N_17343);
and U17601 (N_17601,N_17493,N_17324);
nor U17602 (N_17602,N_17333,N_17372);
nand U17603 (N_17603,N_17310,N_17309);
nor U17604 (N_17604,N_17276,N_17357);
and U17605 (N_17605,N_17385,N_17317);
and U17606 (N_17606,N_17491,N_17393);
xnor U17607 (N_17607,N_17482,N_17474);
and U17608 (N_17608,N_17325,N_17477);
or U17609 (N_17609,N_17425,N_17313);
and U17610 (N_17610,N_17389,N_17346);
or U17611 (N_17611,N_17318,N_17368);
and U17612 (N_17612,N_17254,N_17406);
and U17613 (N_17613,N_17263,N_17443);
xnor U17614 (N_17614,N_17341,N_17258);
and U17615 (N_17615,N_17392,N_17302);
xor U17616 (N_17616,N_17471,N_17418);
xnor U17617 (N_17617,N_17314,N_17378);
nand U17618 (N_17618,N_17349,N_17307);
or U17619 (N_17619,N_17373,N_17259);
or U17620 (N_17620,N_17383,N_17355);
and U17621 (N_17621,N_17412,N_17348);
nand U17622 (N_17622,N_17295,N_17465);
nor U17623 (N_17623,N_17473,N_17360);
and U17624 (N_17624,N_17456,N_17495);
nor U17625 (N_17625,N_17266,N_17355);
and U17626 (N_17626,N_17378,N_17498);
and U17627 (N_17627,N_17298,N_17312);
xor U17628 (N_17628,N_17403,N_17260);
nor U17629 (N_17629,N_17355,N_17407);
or U17630 (N_17630,N_17321,N_17434);
nand U17631 (N_17631,N_17320,N_17395);
nor U17632 (N_17632,N_17323,N_17298);
and U17633 (N_17633,N_17404,N_17445);
and U17634 (N_17634,N_17387,N_17385);
and U17635 (N_17635,N_17309,N_17406);
nor U17636 (N_17636,N_17483,N_17264);
and U17637 (N_17637,N_17410,N_17369);
xor U17638 (N_17638,N_17310,N_17344);
nand U17639 (N_17639,N_17418,N_17348);
and U17640 (N_17640,N_17299,N_17493);
nor U17641 (N_17641,N_17296,N_17413);
nor U17642 (N_17642,N_17260,N_17399);
and U17643 (N_17643,N_17344,N_17277);
xor U17644 (N_17644,N_17318,N_17314);
xor U17645 (N_17645,N_17276,N_17376);
and U17646 (N_17646,N_17453,N_17455);
nor U17647 (N_17647,N_17290,N_17345);
xnor U17648 (N_17648,N_17322,N_17382);
nor U17649 (N_17649,N_17257,N_17394);
and U17650 (N_17650,N_17318,N_17411);
nand U17651 (N_17651,N_17336,N_17441);
nand U17652 (N_17652,N_17309,N_17340);
or U17653 (N_17653,N_17463,N_17460);
and U17654 (N_17654,N_17405,N_17358);
nor U17655 (N_17655,N_17273,N_17410);
nor U17656 (N_17656,N_17363,N_17315);
and U17657 (N_17657,N_17479,N_17419);
nor U17658 (N_17658,N_17394,N_17265);
or U17659 (N_17659,N_17472,N_17312);
or U17660 (N_17660,N_17423,N_17456);
nand U17661 (N_17661,N_17495,N_17499);
and U17662 (N_17662,N_17311,N_17496);
or U17663 (N_17663,N_17496,N_17295);
and U17664 (N_17664,N_17334,N_17362);
xnor U17665 (N_17665,N_17254,N_17368);
and U17666 (N_17666,N_17385,N_17312);
nand U17667 (N_17667,N_17295,N_17443);
xor U17668 (N_17668,N_17322,N_17411);
xor U17669 (N_17669,N_17333,N_17352);
nor U17670 (N_17670,N_17448,N_17373);
and U17671 (N_17671,N_17421,N_17261);
or U17672 (N_17672,N_17393,N_17496);
xnor U17673 (N_17673,N_17281,N_17416);
and U17674 (N_17674,N_17406,N_17427);
nor U17675 (N_17675,N_17404,N_17332);
and U17676 (N_17676,N_17468,N_17266);
nor U17677 (N_17677,N_17462,N_17262);
xnor U17678 (N_17678,N_17419,N_17388);
nor U17679 (N_17679,N_17381,N_17493);
nand U17680 (N_17680,N_17263,N_17336);
xor U17681 (N_17681,N_17339,N_17461);
and U17682 (N_17682,N_17442,N_17429);
xor U17683 (N_17683,N_17401,N_17304);
xnor U17684 (N_17684,N_17290,N_17418);
and U17685 (N_17685,N_17301,N_17360);
nor U17686 (N_17686,N_17265,N_17462);
xor U17687 (N_17687,N_17415,N_17251);
or U17688 (N_17688,N_17419,N_17327);
nor U17689 (N_17689,N_17252,N_17351);
nor U17690 (N_17690,N_17384,N_17372);
nor U17691 (N_17691,N_17357,N_17340);
or U17692 (N_17692,N_17421,N_17293);
and U17693 (N_17693,N_17358,N_17491);
nand U17694 (N_17694,N_17281,N_17357);
xnor U17695 (N_17695,N_17397,N_17382);
nand U17696 (N_17696,N_17475,N_17377);
nand U17697 (N_17697,N_17394,N_17461);
nand U17698 (N_17698,N_17396,N_17261);
nand U17699 (N_17699,N_17375,N_17490);
nand U17700 (N_17700,N_17490,N_17282);
nor U17701 (N_17701,N_17331,N_17369);
and U17702 (N_17702,N_17351,N_17488);
xnor U17703 (N_17703,N_17430,N_17318);
nand U17704 (N_17704,N_17371,N_17358);
nor U17705 (N_17705,N_17314,N_17345);
xor U17706 (N_17706,N_17444,N_17461);
and U17707 (N_17707,N_17318,N_17441);
xnor U17708 (N_17708,N_17296,N_17355);
and U17709 (N_17709,N_17464,N_17349);
or U17710 (N_17710,N_17426,N_17258);
xnor U17711 (N_17711,N_17310,N_17422);
nor U17712 (N_17712,N_17427,N_17349);
and U17713 (N_17713,N_17468,N_17486);
nand U17714 (N_17714,N_17306,N_17262);
xnor U17715 (N_17715,N_17463,N_17351);
and U17716 (N_17716,N_17403,N_17485);
nand U17717 (N_17717,N_17445,N_17399);
and U17718 (N_17718,N_17315,N_17449);
or U17719 (N_17719,N_17352,N_17490);
xnor U17720 (N_17720,N_17365,N_17380);
xnor U17721 (N_17721,N_17364,N_17395);
nand U17722 (N_17722,N_17289,N_17465);
nor U17723 (N_17723,N_17250,N_17415);
nand U17724 (N_17724,N_17488,N_17367);
nand U17725 (N_17725,N_17426,N_17337);
xnor U17726 (N_17726,N_17406,N_17310);
nand U17727 (N_17727,N_17262,N_17333);
nor U17728 (N_17728,N_17295,N_17360);
xor U17729 (N_17729,N_17365,N_17268);
xnor U17730 (N_17730,N_17340,N_17264);
nor U17731 (N_17731,N_17312,N_17323);
nand U17732 (N_17732,N_17280,N_17384);
and U17733 (N_17733,N_17461,N_17295);
nand U17734 (N_17734,N_17421,N_17325);
and U17735 (N_17735,N_17448,N_17419);
nor U17736 (N_17736,N_17430,N_17454);
xor U17737 (N_17737,N_17451,N_17420);
xor U17738 (N_17738,N_17327,N_17257);
and U17739 (N_17739,N_17323,N_17345);
nand U17740 (N_17740,N_17386,N_17375);
nor U17741 (N_17741,N_17462,N_17397);
nor U17742 (N_17742,N_17271,N_17396);
and U17743 (N_17743,N_17415,N_17266);
nand U17744 (N_17744,N_17392,N_17335);
and U17745 (N_17745,N_17398,N_17298);
xor U17746 (N_17746,N_17460,N_17413);
xor U17747 (N_17747,N_17463,N_17425);
or U17748 (N_17748,N_17384,N_17432);
or U17749 (N_17749,N_17262,N_17275);
nor U17750 (N_17750,N_17535,N_17665);
nor U17751 (N_17751,N_17676,N_17719);
or U17752 (N_17752,N_17557,N_17522);
xor U17753 (N_17753,N_17650,N_17574);
or U17754 (N_17754,N_17662,N_17661);
and U17755 (N_17755,N_17521,N_17698);
nand U17756 (N_17756,N_17524,N_17612);
nand U17757 (N_17757,N_17552,N_17634);
nand U17758 (N_17758,N_17556,N_17692);
nand U17759 (N_17759,N_17605,N_17613);
and U17760 (N_17760,N_17617,N_17562);
nor U17761 (N_17761,N_17614,N_17673);
nand U17762 (N_17762,N_17685,N_17563);
xnor U17763 (N_17763,N_17532,N_17677);
nor U17764 (N_17764,N_17620,N_17606);
or U17765 (N_17765,N_17514,N_17508);
and U17766 (N_17766,N_17599,N_17529);
or U17767 (N_17767,N_17587,N_17538);
or U17768 (N_17768,N_17633,N_17517);
xor U17769 (N_17769,N_17659,N_17667);
or U17770 (N_17770,N_17509,N_17630);
nor U17771 (N_17771,N_17624,N_17635);
nor U17772 (N_17772,N_17717,N_17656);
nand U17773 (N_17773,N_17678,N_17669);
nor U17774 (N_17774,N_17530,N_17578);
xor U17775 (N_17775,N_17705,N_17622);
xnor U17776 (N_17776,N_17603,N_17520);
or U17777 (N_17777,N_17636,N_17734);
nor U17778 (N_17778,N_17646,N_17727);
xnor U17779 (N_17779,N_17592,N_17593);
xnor U17780 (N_17780,N_17604,N_17644);
xnor U17781 (N_17781,N_17648,N_17699);
nor U17782 (N_17782,N_17567,N_17642);
and U17783 (N_17783,N_17637,N_17658);
or U17784 (N_17784,N_17742,N_17697);
and U17785 (N_17785,N_17684,N_17700);
or U17786 (N_17786,N_17576,N_17581);
nor U17787 (N_17787,N_17626,N_17501);
nor U17788 (N_17788,N_17741,N_17591);
and U17789 (N_17789,N_17730,N_17610);
nand U17790 (N_17790,N_17660,N_17531);
xnor U17791 (N_17791,N_17570,N_17694);
or U17792 (N_17792,N_17670,N_17598);
nand U17793 (N_17793,N_17554,N_17731);
xor U17794 (N_17794,N_17527,N_17681);
nor U17795 (N_17795,N_17549,N_17643);
nand U17796 (N_17796,N_17687,N_17680);
nor U17797 (N_17797,N_17537,N_17629);
and U17798 (N_17798,N_17722,N_17615);
or U17799 (N_17799,N_17573,N_17735);
xor U17800 (N_17800,N_17739,N_17523);
nand U17801 (N_17801,N_17690,N_17616);
xnor U17802 (N_17802,N_17663,N_17723);
xnor U17803 (N_17803,N_17547,N_17512);
or U17804 (N_17804,N_17540,N_17707);
and U17805 (N_17805,N_17748,N_17714);
or U17806 (N_17806,N_17647,N_17601);
or U17807 (N_17807,N_17544,N_17541);
nand U17808 (N_17808,N_17589,N_17596);
and U17809 (N_17809,N_17619,N_17546);
xor U17810 (N_17810,N_17608,N_17548);
xor U17811 (N_17811,N_17513,N_17590);
and U17812 (N_17812,N_17693,N_17696);
nor U17813 (N_17813,N_17747,N_17568);
or U17814 (N_17814,N_17724,N_17565);
and U17815 (N_17815,N_17738,N_17701);
and U17816 (N_17816,N_17721,N_17510);
or U17817 (N_17817,N_17618,N_17718);
xor U17818 (N_17818,N_17516,N_17505);
nor U17819 (N_17819,N_17611,N_17609);
or U17820 (N_17820,N_17720,N_17628);
xnor U17821 (N_17821,N_17621,N_17594);
xor U17822 (N_17822,N_17526,N_17695);
and U17823 (N_17823,N_17586,N_17506);
nor U17824 (N_17824,N_17525,N_17746);
xor U17825 (N_17825,N_17625,N_17715);
and U17826 (N_17826,N_17645,N_17623);
nand U17827 (N_17827,N_17649,N_17518);
nor U17828 (N_17828,N_17671,N_17745);
nand U17829 (N_17829,N_17500,N_17712);
and U17830 (N_17830,N_17551,N_17713);
nand U17831 (N_17831,N_17640,N_17706);
or U17832 (N_17832,N_17564,N_17654);
and U17833 (N_17833,N_17675,N_17580);
nor U17834 (N_17834,N_17653,N_17632);
or U17835 (N_17835,N_17511,N_17691);
nor U17836 (N_17836,N_17566,N_17588);
or U17837 (N_17837,N_17543,N_17726);
nor U17838 (N_17838,N_17703,N_17553);
xnor U17839 (N_17839,N_17539,N_17711);
or U17840 (N_17840,N_17716,N_17584);
xor U17841 (N_17841,N_17582,N_17561);
xor U17842 (N_17842,N_17569,N_17736);
or U17843 (N_17843,N_17641,N_17668);
nor U17844 (N_17844,N_17631,N_17627);
nand U17845 (N_17845,N_17725,N_17536);
nand U17846 (N_17846,N_17550,N_17585);
and U17847 (N_17847,N_17704,N_17729);
nand U17848 (N_17848,N_17728,N_17710);
and U17849 (N_17849,N_17558,N_17749);
nor U17850 (N_17850,N_17639,N_17733);
or U17851 (N_17851,N_17519,N_17672);
nor U17852 (N_17852,N_17575,N_17708);
and U17853 (N_17853,N_17740,N_17602);
xor U17854 (N_17854,N_17515,N_17683);
nand U17855 (N_17855,N_17674,N_17595);
xnor U17856 (N_17856,N_17600,N_17664);
nand U17857 (N_17857,N_17709,N_17534);
nor U17858 (N_17858,N_17533,N_17655);
and U17859 (N_17859,N_17666,N_17689);
and U17860 (N_17860,N_17583,N_17560);
or U17861 (N_17861,N_17504,N_17743);
xnor U17862 (N_17862,N_17732,N_17572);
xnor U17863 (N_17863,N_17651,N_17577);
nand U17864 (N_17864,N_17542,N_17652);
nor U17865 (N_17865,N_17744,N_17507);
xnor U17866 (N_17866,N_17737,N_17555);
xnor U17867 (N_17867,N_17502,N_17597);
nor U17868 (N_17868,N_17571,N_17686);
nand U17869 (N_17869,N_17688,N_17679);
xor U17870 (N_17870,N_17682,N_17638);
or U17871 (N_17871,N_17528,N_17545);
nand U17872 (N_17872,N_17607,N_17579);
and U17873 (N_17873,N_17702,N_17559);
xnor U17874 (N_17874,N_17503,N_17657);
xnor U17875 (N_17875,N_17676,N_17635);
xor U17876 (N_17876,N_17592,N_17746);
xnor U17877 (N_17877,N_17672,N_17611);
nand U17878 (N_17878,N_17608,N_17624);
nand U17879 (N_17879,N_17501,N_17684);
nand U17880 (N_17880,N_17640,N_17607);
nor U17881 (N_17881,N_17701,N_17687);
xor U17882 (N_17882,N_17717,N_17601);
and U17883 (N_17883,N_17720,N_17687);
xor U17884 (N_17884,N_17674,N_17543);
xor U17885 (N_17885,N_17564,N_17578);
and U17886 (N_17886,N_17733,N_17504);
xor U17887 (N_17887,N_17638,N_17557);
nor U17888 (N_17888,N_17541,N_17585);
xnor U17889 (N_17889,N_17624,N_17570);
or U17890 (N_17890,N_17594,N_17501);
nand U17891 (N_17891,N_17593,N_17516);
or U17892 (N_17892,N_17632,N_17621);
and U17893 (N_17893,N_17567,N_17722);
nor U17894 (N_17894,N_17598,N_17619);
or U17895 (N_17895,N_17739,N_17544);
nor U17896 (N_17896,N_17524,N_17651);
nor U17897 (N_17897,N_17523,N_17582);
or U17898 (N_17898,N_17644,N_17704);
and U17899 (N_17899,N_17587,N_17549);
nor U17900 (N_17900,N_17664,N_17682);
nor U17901 (N_17901,N_17667,N_17717);
or U17902 (N_17902,N_17691,N_17519);
and U17903 (N_17903,N_17720,N_17527);
or U17904 (N_17904,N_17621,N_17602);
or U17905 (N_17905,N_17519,N_17720);
nor U17906 (N_17906,N_17514,N_17650);
nor U17907 (N_17907,N_17527,N_17703);
or U17908 (N_17908,N_17730,N_17622);
nor U17909 (N_17909,N_17545,N_17574);
xor U17910 (N_17910,N_17626,N_17673);
nand U17911 (N_17911,N_17567,N_17585);
or U17912 (N_17912,N_17576,N_17542);
nor U17913 (N_17913,N_17605,N_17746);
or U17914 (N_17914,N_17547,N_17593);
and U17915 (N_17915,N_17635,N_17550);
and U17916 (N_17916,N_17658,N_17570);
or U17917 (N_17917,N_17532,N_17739);
nor U17918 (N_17918,N_17529,N_17676);
nor U17919 (N_17919,N_17555,N_17514);
or U17920 (N_17920,N_17695,N_17647);
and U17921 (N_17921,N_17538,N_17517);
or U17922 (N_17922,N_17566,N_17676);
xor U17923 (N_17923,N_17639,N_17645);
and U17924 (N_17924,N_17631,N_17522);
and U17925 (N_17925,N_17653,N_17510);
or U17926 (N_17926,N_17686,N_17507);
and U17927 (N_17927,N_17631,N_17584);
nor U17928 (N_17928,N_17554,N_17508);
xor U17929 (N_17929,N_17593,N_17623);
nand U17930 (N_17930,N_17626,N_17714);
and U17931 (N_17931,N_17576,N_17523);
nand U17932 (N_17932,N_17701,N_17514);
nor U17933 (N_17933,N_17532,N_17560);
or U17934 (N_17934,N_17532,N_17680);
nand U17935 (N_17935,N_17724,N_17645);
or U17936 (N_17936,N_17735,N_17625);
nor U17937 (N_17937,N_17602,N_17508);
nor U17938 (N_17938,N_17697,N_17662);
nor U17939 (N_17939,N_17513,N_17562);
nand U17940 (N_17940,N_17665,N_17699);
nand U17941 (N_17941,N_17535,N_17600);
and U17942 (N_17942,N_17586,N_17532);
or U17943 (N_17943,N_17692,N_17673);
or U17944 (N_17944,N_17662,N_17682);
or U17945 (N_17945,N_17605,N_17660);
nand U17946 (N_17946,N_17711,N_17733);
or U17947 (N_17947,N_17588,N_17675);
xor U17948 (N_17948,N_17742,N_17699);
nand U17949 (N_17949,N_17743,N_17650);
and U17950 (N_17950,N_17707,N_17747);
nand U17951 (N_17951,N_17518,N_17617);
nor U17952 (N_17952,N_17705,N_17536);
or U17953 (N_17953,N_17617,N_17642);
xor U17954 (N_17954,N_17562,N_17540);
and U17955 (N_17955,N_17640,N_17627);
and U17956 (N_17956,N_17545,N_17521);
or U17957 (N_17957,N_17674,N_17732);
xnor U17958 (N_17958,N_17580,N_17665);
nor U17959 (N_17959,N_17558,N_17560);
nand U17960 (N_17960,N_17510,N_17562);
nor U17961 (N_17961,N_17627,N_17562);
nand U17962 (N_17962,N_17749,N_17676);
nor U17963 (N_17963,N_17736,N_17600);
xor U17964 (N_17964,N_17708,N_17590);
and U17965 (N_17965,N_17686,N_17688);
nand U17966 (N_17966,N_17613,N_17586);
xnor U17967 (N_17967,N_17563,N_17721);
nor U17968 (N_17968,N_17600,N_17646);
and U17969 (N_17969,N_17506,N_17730);
or U17970 (N_17970,N_17590,N_17575);
xor U17971 (N_17971,N_17515,N_17642);
nor U17972 (N_17972,N_17734,N_17747);
nand U17973 (N_17973,N_17733,N_17586);
xor U17974 (N_17974,N_17732,N_17535);
nand U17975 (N_17975,N_17705,N_17564);
xnor U17976 (N_17976,N_17679,N_17582);
and U17977 (N_17977,N_17713,N_17607);
nand U17978 (N_17978,N_17741,N_17509);
xnor U17979 (N_17979,N_17599,N_17605);
xor U17980 (N_17980,N_17570,N_17717);
and U17981 (N_17981,N_17652,N_17574);
nor U17982 (N_17982,N_17528,N_17717);
and U17983 (N_17983,N_17628,N_17749);
or U17984 (N_17984,N_17587,N_17699);
nand U17985 (N_17985,N_17545,N_17529);
xor U17986 (N_17986,N_17633,N_17748);
and U17987 (N_17987,N_17510,N_17565);
or U17988 (N_17988,N_17509,N_17546);
xor U17989 (N_17989,N_17743,N_17569);
xnor U17990 (N_17990,N_17567,N_17575);
nand U17991 (N_17991,N_17583,N_17585);
or U17992 (N_17992,N_17710,N_17619);
nor U17993 (N_17993,N_17749,N_17710);
and U17994 (N_17994,N_17522,N_17569);
nand U17995 (N_17995,N_17690,N_17568);
or U17996 (N_17996,N_17688,N_17596);
nor U17997 (N_17997,N_17556,N_17514);
or U17998 (N_17998,N_17709,N_17746);
nand U17999 (N_17999,N_17685,N_17717);
nand U18000 (N_18000,N_17751,N_17837);
nand U18001 (N_18001,N_17933,N_17826);
xor U18002 (N_18002,N_17990,N_17970);
nor U18003 (N_18003,N_17938,N_17960);
and U18004 (N_18004,N_17906,N_17770);
or U18005 (N_18005,N_17803,N_17758);
nor U18006 (N_18006,N_17936,N_17772);
xor U18007 (N_18007,N_17877,N_17842);
nand U18008 (N_18008,N_17783,N_17871);
xnor U18009 (N_18009,N_17829,N_17808);
xor U18010 (N_18010,N_17855,N_17827);
or U18011 (N_18011,N_17781,N_17780);
nor U18012 (N_18012,N_17908,N_17879);
nand U18013 (N_18013,N_17997,N_17895);
nand U18014 (N_18014,N_17915,N_17948);
nor U18015 (N_18015,N_17801,N_17995);
nand U18016 (N_18016,N_17755,N_17993);
nor U18017 (N_18017,N_17784,N_17986);
xor U18018 (N_18018,N_17853,N_17882);
nand U18019 (N_18019,N_17901,N_17893);
nor U18020 (N_18020,N_17898,N_17917);
and U18021 (N_18021,N_17896,N_17905);
nor U18022 (N_18022,N_17765,N_17954);
nand U18023 (N_18023,N_17762,N_17813);
nand U18024 (N_18024,N_17787,N_17932);
nand U18025 (N_18025,N_17806,N_17891);
nand U18026 (N_18026,N_17814,N_17923);
nand U18027 (N_18027,N_17909,N_17867);
nor U18028 (N_18028,N_17976,N_17897);
and U18029 (N_18029,N_17860,N_17825);
nor U18030 (N_18030,N_17779,N_17956);
xor U18031 (N_18031,N_17939,N_17988);
xnor U18032 (N_18032,N_17963,N_17778);
and U18033 (N_18033,N_17822,N_17768);
xor U18034 (N_18034,N_17964,N_17916);
or U18035 (N_18035,N_17987,N_17759);
and U18036 (N_18036,N_17969,N_17982);
nor U18037 (N_18037,N_17953,N_17880);
and U18038 (N_18038,N_17972,N_17856);
xor U18039 (N_18039,N_17873,N_17782);
and U18040 (N_18040,N_17830,N_17919);
and U18041 (N_18041,N_17999,N_17753);
nor U18042 (N_18042,N_17810,N_17984);
nor U18043 (N_18043,N_17818,N_17869);
nor U18044 (N_18044,N_17854,N_17796);
nand U18045 (N_18045,N_17764,N_17838);
nand U18046 (N_18046,N_17973,N_17942);
nand U18047 (N_18047,N_17754,N_17921);
and U18048 (N_18048,N_17811,N_17851);
nor U18049 (N_18049,N_17892,N_17950);
or U18050 (N_18050,N_17831,N_17777);
nand U18051 (N_18051,N_17760,N_17868);
xor U18052 (N_18052,N_17859,N_17983);
nand U18053 (N_18053,N_17996,N_17857);
nor U18054 (N_18054,N_17752,N_17918);
nand U18055 (N_18055,N_17925,N_17807);
xnor U18056 (N_18056,N_17816,N_17815);
nand U18057 (N_18057,N_17889,N_17903);
xnor U18058 (N_18058,N_17791,N_17914);
and U18059 (N_18059,N_17788,N_17794);
and U18060 (N_18060,N_17978,N_17797);
and U18061 (N_18061,N_17949,N_17817);
nand U18062 (N_18062,N_17989,N_17907);
and U18063 (N_18063,N_17894,N_17836);
and U18064 (N_18064,N_17945,N_17971);
or U18065 (N_18065,N_17861,N_17863);
or U18066 (N_18066,N_17958,N_17910);
nand U18067 (N_18067,N_17902,N_17841);
or U18068 (N_18068,N_17930,N_17756);
nand U18069 (N_18069,N_17773,N_17750);
or U18070 (N_18070,N_17800,N_17952);
xnor U18071 (N_18071,N_17965,N_17876);
and U18072 (N_18072,N_17994,N_17844);
and U18073 (N_18073,N_17824,N_17883);
nor U18074 (N_18074,N_17967,N_17771);
nand U18075 (N_18075,N_17828,N_17944);
xnor U18076 (N_18076,N_17946,N_17798);
or U18077 (N_18077,N_17874,N_17819);
and U18078 (N_18078,N_17820,N_17795);
xor U18079 (N_18079,N_17899,N_17900);
or U18080 (N_18080,N_17941,N_17786);
nand U18081 (N_18081,N_17924,N_17955);
and U18082 (N_18082,N_17920,N_17943);
xnor U18083 (N_18083,N_17872,N_17913);
and U18084 (N_18084,N_17966,N_17864);
xor U18085 (N_18085,N_17878,N_17929);
and U18086 (N_18086,N_17974,N_17804);
nor U18087 (N_18087,N_17885,N_17852);
and U18088 (N_18088,N_17775,N_17928);
nand U18089 (N_18089,N_17833,N_17843);
xnor U18090 (N_18090,N_17934,N_17846);
or U18091 (N_18091,N_17850,N_17866);
nor U18092 (N_18092,N_17935,N_17792);
nor U18093 (N_18093,N_17961,N_17858);
and U18094 (N_18094,N_17769,N_17927);
and U18095 (N_18095,N_17881,N_17937);
nor U18096 (N_18096,N_17805,N_17870);
or U18097 (N_18097,N_17847,N_17849);
nand U18098 (N_18098,N_17862,N_17979);
xnor U18099 (N_18099,N_17912,N_17980);
nand U18100 (N_18100,N_17834,N_17975);
or U18101 (N_18101,N_17940,N_17985);
and U18102 (N_18102,N_17931,N_17904);
nand U18103 (N_18103,N_17761,N_17790);
or U18104 (N_18104,N_17951,N_17835);
xnor U18105 (N_18105,N_17812,N_17959);
nand U18106 (N_18106,N_17785,N_17888);
nor U18107 (N_18107,N_17763,N_17981);
and U18108 (N_18108,N_17793,N_17799);
xnor U18109 (N_18109,N_17922,N_17968);
or U18110 (N_18110,N_17992,N_17998);
nand U18111 (N_18111,N_17802,N_17789);
xor U18112 (N_18112,N_17962,N_17911);
xor U18113 (N_18113,N_17821,N_17848);
and U18114 (N_18114,N_17887,N_17947);
nor U18115 (N_18115,N_17845,N_17890);
xnor U18116 (N_18116,N_17774,N_17957);
or U18117 (N_18117,N_17832,N_17875);
or U18118 (N_18118,N_17886,N_17977);
nor U18119 (N_18119,N_17766,N_17865);
nand U18120 (N_18120,N_17823,N_17884);
xnor U18121 (N_18121,N_17767,N_17809);
or U18122 (N_18122,N_17840,N_17926);
or U18123 (N_18123,N_17991,N_17776);
xnor U18124 (N_18124,N_17839,N_17757);
and U18125 (N_18125,N_17888,N_17828);
and U18126 (N_18126,N_17828,N_17883);
xnor U18127 (N_18127,N_17966,N_17924);
nor U18128 (N_18128,N_17951,N_17796);
or U18129 (N_18129,N_17765,N_17788);
xor U18130 (N_18130,N_17782,N_17952);
or U18131 (N_18131,N_17835,N_17883);
nor U18132 (N_18132,N_17908,N_17780);
nand U18133 (N_18133,N_17933,N_17878);
nor U18134 (N_18134,N_17888,N_17869);
xnor U18135 (N_18135,N_17979,N_17965);
nor U18136 (N_18136,N_17890,N_17773);
xnor U18137 (N_18137,N_17802,N_17817);
and U18138 (N_18138,N_17966,N_17965);
nand U18139 (N_18139,N_17793,N_17819);
xor U18140 (N_18140,N_17875,N_17822);
or U18141 (N_18141,N_17807,N_17926);
nand U18142 (N_18142,N_17816,N_17976);
xnor U18143 (N_18143,N_17873,N_17856);
xor U18144 (N_18144,N_17778,N_17991);
nand U18145 (N_18145,N_17912,N_17891);
or U18146 (N_18146,N_17920,N_17791);
or U18147 (N_18147,N_17825,N_17798);
nand U18148 (N_18148,N_17908,N_17934);
or U18149 (N_18149,N_17885,N_17778);
or U18150 (N_18150,N_17908,N_17830);
and U18151 (N_18151,N_17991,N_17980);
nor U18152 (N_18152,N_17865,N_17811);
and U18153 (N_18153,N_17848,N_17950);
xnor U18154 (N_18154,N_17898,N_17886);
or U18155 (N_18155,N_17812,N_17927);
and U18156 (N_18156,N_17912,N_17803);
nand U18157 (N_18157,N_17789,N_17965);
nand U18158 (N_18158,N_17906,N_17814);
xnor U18159 (N_18159,N_17771,N_17916);
xor U18160 (N_18160,N_17771,N_17828);
and U18161 (N_18161,N_17757,N_17750);
nand U18162 (N_18162,N_17833,N_17905);
xnor U18163 (N_18163,N_17914,N_17812);
xor U18164 (N_18164,N_17997,N_17890);
xnor U18165 (N_18165,N_17787,N_17901);
xor U18166 (N_18166,N_17999,N_17947);
nor U18167 (N_18167,N_17920,N_17760);
and U18168 (N_18168,N_17902,N_17915);
nor U18169 (N_18169,N_17760,N_17924);
nand U18170 (N_18170,N_17897,N_17875);
xor U18171 (N_18171,N_17786,N_17940);
nor U18172 (N_18172,N_17943,N_17966);
or U18173 (N_18173,N_17902,N_17816);
nor U18174 (N_18174,N_17985,N_17784);
nor U18175 (N_18175,N_17920,N_17803);
nand U18176 (N_18176,N_17965,N_17985);
and U18177 (N_18177,N_17805,N_17773);
and U18178 (N_18178,N_17814,N_17762);
nand U18179 (N_18179,N_17954,N_17852);
or U18180 (N_18180,N_17751,N_17888);
or U18181 (N_18181,N_17957,N_17993);
xnor U18182 (N_18182,N_17827,N_17917);
xnor U18183 (N_18183,N_17854,N_17887);
and U18184 (N_18184,N_17862,N_17991);
or U18185 (N_18185,N_17900,N_17995);
xor U18186 (N_18186,N_17965,N_17779);
or U18187 (N_18187,N_17878,N_17966);
or U18188 (N_18188,N_17837,N_17817);
or U18189 (N_18189,N_17770,N_17981);
nor U18190 (N_18190,N_17798,N_17994);
or U18191 (N_18191,N_17967,N_17784);
nand U18192 (N_18192,N_17902,N_17961);
or U18193 (N_18193,N_17858,N_17918);
nand U18194 (N_18194,N_17991,N_17937);
and U18195 (N_18195,N_17982,N_17930);
xnor U18196 (N_18196,N_17933,N_17864);
nand U18197 (N_18197,N_17959,N_17969);
xor U18198 (N_18198,N_17844,N_17802);
nor U18199 (N_18199,N_17753,N_17918);
or U18200 (N_18200,N_17982,N_17997);
nor U18201 (N_18201,N_17896,N_17774);
nand U18202 (N_18202,N_17759,N_17959);
or U18203 (N_18203,N_17769,N_17905);
or U18204 (N_18204,N_17773,N_17885);
and U18205 (N_18205,N_17880,N_17944);
nand U18206 (N_18206,N_17858,N_17841);
nand U18207 (N_18207,N_17972,N_17897);
or U18208 (N_18208,N_17881,N_17803);
and U18209 (N_18209,N_17985,N_17773);
nand U18210 (N_18210,N_17801,N_17871);
nor U18211 (N_18211,N_17930,N_17900);
or U18212 (N_18212,N_17870,N_17895);
and U18213 (N_18213,N_17750,N_17896);
or U18214 (N_18214,N_17897,N_17851);
nand U18215 (N_18215,N_17893,N_17784);
nand U18216 (N_18216,N_17980,N_17754);
or U18217 (N_18217,N_17774,N_17811);
nand U18218 (N_18218,N_17907,N_17895);
and U18219 (N_18219,N_17838,N_17999);
or U18220 (N_18220,N_17857,N_17990);
nand U18221 (N_18221,N_17901,N_17824);
and U18222 (N_18222,N_17926,N_17928);
nand U18223 (N_18223,N_17869,N_17929);
nand U18224 (N_18224,N_17906,N_17956);
nand U18225 (N_18225,N_17972,N_17782);
nor U18226 (N_18226,N_17836,N_17754);
nor U18227 (N_18227,N_17863,N_17834);
and U18228 (N_18228,N_17901,N_17981);
nand U18229 (N_18229,N_17896,N_17887);
or U18230 (N_18230,N_17813,N_17945);
nor U18231 (N_18231,N_17753,N_17944);
xor U18232 (N_18232,N_17920,N_17973);
or U18233 (N_18233,N_17864,N_17856);
and U18234 (N_18234,N_17903,N_17802);
and U18235 (N_18235,N_17904,N_17775);
xor U18236 (N_18236,N_17806,N_17885);
or U18237 (N_18237,N_17823,N_17851);
xor U18238 (N_18238,N_17850,N_17942);
xor U18239 (N_18239,N_17823,N_17803);
nor U18240 (N_18240,N_17994,N_17762);
and U18241 (N_18241,N_17944,N_17910);
or U18242 (N_18242,N_17938,N_17881);
or U18243 (N_18243,N_17930,N_17892);
and U18244 (N_18244,N_17798,N_17765);
xor U18245 (N_18245,N_17916,N_17766);
or U18246 (N_18246,N_17961,N_17769);
nor U18247 (N_18247,N_17819,N_17837);
nand U18248 (N_18248,N_17922,N_17980);
nor U18249 (N_18249,N_17920,N_17832);
nor U18250 (N_18250,N_18012,N_18196);
nand U18251 (N_18251,N_18040,N_18140);
xnor U18252 (N_18252,N_18179,N_18124);
and U18253 (N_18253,N_18072,N_18200);
nand U18254 (N_18254,N_18038,N_18095);
nor U18255 (N_18255,N_18067,N_18089);
xnor U18256 (N_18256,N_18151,N_18071);
nand U18257 (N_18257,N_18086,N_18016);
nand U18258 (N_18258,N_18119,N_18125);
nor U18259 (N_18259,N_18034,N_18215);
or U18260 (N_18260,N_18002,N_18000);
or U18261 (N_18261,N_18050,N_18005);
and U18262 (N_18262,N_18139,N_18168);
or U18263 (N_18263,N_18047,N_18195);
xnor U18264 (N_18264,N_18141,N_18004);
xnor U18265 (N_18265,N_18030,N_18156);
or U18266 (N_18266,N_18134,N_18246);
xnor U18267 (N_18267,N_18148,N_18221);
nand U18268 (N_18268,N_18041,N_18234);
xor U18269 (N_18269,N_18094,N_18075);
or U18270 (N_18270,N_18073,N_18060);
xor U18271 (N_18271,N_18091,N_18155);
and U18272 (N_18272,N_18013,N_18216);
and U18273 (N_18273,N_18142,N_18157);
nor U18274 (N_18274,N_18035,N_18115);
xnor U18275 (N_18275,N_18102,N_18009);
or U18276 (N_18276,N_18088,N_18045);
nor U18277 (N_18277,N_18061,N_18146);
and U18278 (N_18278,N_18058,N_18093);
nand U18279 (N_18279,N_18036,N_18027);
and U18280 (N_18280,N_18068,N_18190);
or U18281 (N_18281,N_18025,N_18007);
or U18282 (N_18282,N_18042,N_18219);
nand U18283 (N_18283,N_18112,N_18165);
or U18284 (N_18284,N_18224,N_18017);
or U18285 (N_18285,N_18123,N_18066);
or U18286 (N_18286,N_18121,N_18113);
nand U18287 (N_18287,N_18023,N_18233);
nand U18288 (N_18288,N_18210,N_18178);
xnor U18289 (N_18289,N_18046,N_18109);
and U18290 (N_18290,N_18001,N_18057);
xor U18291 (N_18291,N_18161,N_18191);
and U18292 (N_18292,N_18080,N_18163);
xor U18293 (N_18293,N_18018,N_18127);
or U18294 (N_18294,N_18096,N_18237);
or U18295 (N_18295,N_18218,N_18082);
nand U18296 (N_18296,N_18211,N_18172);
or U18297 (N_18297,N_18169,N_18240);
and U18298 (N_18298,N_18160,N_18201);
nand U18299 (N_18299,N_18049,N_18227);
nor U18300 (N_18300,N_18092,N_18166);
nor U18301 (N_18301,N_18232,N_18114);
and U18302 (N_18302,N_18105,N_18128);
and U18303 (N_18303,N_18126,N_18100);
nor U18304 (N_18304,N_18177,N_18226);
and U18305 (N_18305,N_18242,N_18174);
and U18306 (N_18306,N_18020,N_18063);
nand U18307 (N_18307,N_18241,N_18173);
nand U18308 (N_18308,N_18011,N_18175);
or U18309 (N_18309,N_18158,N_18108);
nand U18310 (N_18310,N_18006,N_18078);
nor U18311 (N_18311,N_18182,N_18199);
nand U18312 (N_18312,N_18135,N_18239);
nor U18313 (N_18313,N_18243,N_18079);
nand U18314 (N_18314,N_18164,N_18137);
or U18315 (N_18315,N_18205,N_18244);
nand U18316 (N_18316,N_18081,N_18110);
xnor U18317 (N_18317,N_18010,N_18170);
nand U18318 (N_18318,N_18107,N_18145);
or U18319 (N_18319,N_18220,N_18162);
or U18320 (N_18320,N_18024,N_18031);
nor U18321 (N_18321,N_18076,N_18209);
nand U18322 (N_18322,N_18090,N_18097);
nand U18323 (N_18323,N_18055,N_18192);
or U18324 (N_18324,N_18197,N_18133);
and U18325 (N_18325,N_18118,N_18064);
nor U18326 (N_18326,N_18202,N_18003);
and U18327 (N_18327,N_18039,N_18033);
and U18328 (N_18328,N_18144,N_18225);
or U18329 (N_18329,N_18249,N_18153);
or U18330 (N_18330,N_18150,N_18152);
and U18331 (N_18331,N_18059,N_18099);
nor U18332 (N_18332,N_18069,N_18203);
xnor U18333 (N_18333,N_18213,N_18181);
and U18334 (N_18334,N_18223,N_18183);
and U18335 (N_18335,N_18014,N_18212);
nand U18336 (N_18336,N_18070,N_18062);
xnor U18337 (N_18337,N_18180,N_18029);
xor U18338 (N_18338,N_18106,N_18189);
or U18339 (N_18339,N_18214,N_18098);
and U18340 (N_18340,N_18056,N_18245);
xnor U18341 (N_18341,N_18228,N_18132);
nand U18342 (N_18342,N_18044,N_18217);
nand U18343 (N_18343,N_18103,N_18037);
xor U18344 (N_18344,N_18208,N_18207);
and U18345 (N_18345,N_18206,N_18026);
or U18346 (N_18346,N_18028,N_18111);
and U18347 (N_18347,N_18147,N_18087);
and U18348 (N_18348,N_18065,N_18101);
nor U18349 (N_18349,N_18131,N_18188);
xnor U18350 (N_18350,N_18015,N_18231);
and U18351 (N_18351,N_18167,N_18008);
nor U18352 (N_18352,N_18053,N_18194);
xor U18353 (N_18353,N_18122,N_18186);
and U18354 (N_18354,N_18229,N_18198);
nand U18355 (N_18355,N_18022,N_18193);
nand U18356 (N_18356,N_18138,N_18236);
nor U18357 (N_18357,N_18247,N_18104);
nor U18358 (N_18358,N_18230,N_18074);
xor U18359 (N_18359,N_18136,N_18159);
or U18360 (N_18360,N_18129,N_18143);
nand U18361 (N_18361,N_18083,N_18248);
or U18362 (N_18362,N_18120,N_18019);
or U18363 (N_18363,N_18130,N_18185);
or U18364 (N_18364,N_18222,N_18043);
or U18365 (N_18365,N_18054,N_18021);
nand U18366 (N_18366,N_18187,N_18176);
and U18367 (N_18367,N_18117,N_18184);
nand U18368 (N_18368,N_18051,N_18154);
nand U18369 (N_18369,N_18116,N_18032);
or U18370 (N_18370,N_18085,N_18048);
nor U18371 (N_18371,N_18204,N_18238);
and U18372 (N_18372,N_18149,N_18084);
or U18373 (N_18373,N_18052,N_18171);
xnor U18374 (N_18374,N_18077,N_18235);
nor U18375 (N_18375,N_18206,N_18176);
and U18376 (N_18376,N_18116,N_18209);
xnor U18377 (N_18377,N_18176,N_18217);
or U18378 (N_18378,N_18199,N_18045);
xor U18379 (N_18379,N_18038,N_18033);
or U18380 (N_18380,N_18185,N_18087);
nand U18381 (N_18381,N_18017,N_18161);
xnor U18382 (N_18382,N_18020,N_18249);
or U18383 (N_18383,N_18014,N_18198);
and U18384 (N_18384,N_18007,N_18144);
or U18385 (N_18385,N_18183,N_18184);
nand U18386 (N_18386,N_18140,N_18193);
nand U18387 (N_18387,N_18119,N_18188);
nand U18388 (N_18388,N_18153,N_18236);
nand U18389 (N_18389,N_18124,N_18209);
and U18390 (N_18390,N_18002,N_18075);
nor U18391 (N_18391,N_18083,N_18203);
nor U18392 (N_18392,N_18069,N_18032);
and U18393 (N_18393,N_18152,N_18189);
nand U18394 (N_18394,N_18020,N_18072);
xnor U18395 (N_18395,N_18241,N_18008);
xnor U18396 (N_18396,N_18117,N_18239);
or U18397 (N_18397,N_18079,N_18242);
xnor U18398 (N_18398,N_18176,N_18169);
nand U18399 (N_18399,N_18094,N_18072);
nand U18400 (N_18400,N_18191,N_18195);
nand U18401 (N_18401,N_18155,N_18104);
xnor U18402 (N_18402,N_18094,N_18015);
or U18403 (N_18403,N_18176,N_18077);
and U18404 (N_18404,N_18097,N_18075);
nor U18405 (N_18405,N_18018,N_18238);
and U18406 (N_18406,N_18017,N_18133);
nand U18407 (N_18407,N_18156,N_18132);
nor U18408 (N_18408,N_18095,N_18099);
nor U18409 (N_18409,N_18126,N_18073);
xor U18410 (N_18410,N_18162,N_18133);
and U18411 (N_18411,N_18040,N_18061);
and U18412 (N_18412,N_18227,N_18043);
nand U18413 (N_18413,N_18025,N_18060);
and U18414 (N_18414,N_18154,N_18155);
nor U18415 (N_18415,N_18067,N_18027);
nor U18416 (N_18416,N_18054,N_18084);
or U18417 (N_18417,N_18084,N_18219);
nor U18418 (N_18418,N_18203,N_18089);
nor U18419 (N_18419,N_18233,N_18111);
nand U18420 (N_18420,N_18197,N_18035);
and U18421 (N_18421,N_18023,N_18090);
nand U18422 (N_18422,N_18004,N_18046);
nand U18423 (N_18423,N_18046,N_18138);
nor U18424 (N_18424,N_18138,N_18245);
xor U18425 (N_18425,N_18153,N_18089);
nor U18426 (N_18426,N_18148,N_18134);
or U18427 (N_18427,N_18107,N_18126);
and U18428 (N_18428,N_18241,N_18233);
nand U18429 (N_18429,N_18041,N_18160);
nor U18430 (N_18430,N_18002,N_18046);
nor U18431 (N_18431,N_18114,N_18053);
xnor U18432 (N_18432,N_18007,N_18032);
and U18433 (N_18433,N_18245,N_18221);
and U18434 (N_18434,N_18135,N_18130);
nor U18435 (N_18435,N_18026,N_18100);
xor U18436 (N_18436,N_18143,N_18207);
or U18437 (N_18437,N_18029,N_18227);
nand U18438 (N_18438,N_18175,N_18117);
xor U18439 (N_18439,N_18002,N_18006);
nor U18440 (N_18440,N_18090,N_18249);
and U18441 (N_18441,N_18191,N_18023);
and U18442 (N_18442,N_18072,N_18170);
nand U18443 (N_18443,N_18107,N_18061);
or U18444 (N_18444,N_18074,N_18011);
or U18445 (N_18445,N_18113,N_18212);
and U18446 (N_18446,N_18092,N_18086);
nor U18447 (N_18447,N_18204,N_18226);
or U18448 (N_18448,N_18067,N_18229);
and U18449 (N_18449,N_18198,N_18040);
and U18450 (N_18450,N_18112,N_18022);
nor U18451 (N_18451,N_18003,N_18072);
and U18452 (N_18452,N_18163,N_18189);
or U18453 (N_18453,N_18026,N_18034);
nand U18454 (N_18454,N_18198,N_18179);
and U18455 (N_18455,N_18093,N_18183);
nor U18456 (N_18456,N_18116,N_18026);
and U18457 (N_18457,N_18127,N_18238);
nor U18458 (N_18458,N_18041,N_18173);
xor U18459 (N_18459,N_18214,N_18231);
or U18460 (N_18460,N_18098,N_18097);
xor U18461 (N_18461,N_18130,N_18190);
nor U18462 (N_18462,N_18034,N_18188);
nor U18463 (N_18463,N_18084,N_18014);
and U18464 (N_18464,N_18217,N_18204);
or U18465 (N_18465,N_18071,N_18073);
or U18466 (N_18466,N_18244,N_18139);
nand U18467 (N_18467,N_18084,N_18080);
or U18468 (N_18468,N_18014,N_18147);
and U18469 (N_18469,N_18191,N_18122);
and U18470 (N_18470,N_18004,N_18081);
xor U18471 (N_18471,N_18213,N_18149);
or U18472 (N_18472,N_18199,N_18087);
nor U18473 (N_18473,N_18149,N_18079);
or U18474 (N_18474,N_18062,N_18232);
and U18475 (N_18475,N_18126,N_18059);
nand U18476 (N_18476,N_18032,N_18067);
and U18477 (N_18477,N_18082,N_18041);
nand U18478 (N_18478,N_18120,N_18247);
and U18479 (N_18479,N_18086,N_18159);
or U18480 (N_18480,N_18035,N_18133);
nor U18481 (N_18481,N_18156,N_18179);
nand U18482 (N_18482,N_18208,N_18113);
or U18483 (N_18483,N_18094,N_18091);
xnor U18484 (N_18484,N_18080,N_18172);
nand U18485 (N_18485,N_18179,N_18006);
nor U18486 (N_18486,N_18203,N_18041);
or U18487 (N_18487,N_18044,N_18109);
or U18488 (N_18488,N_18193,N_18030);
nor U18489 (N_18489,N_18209,N_18166);
nand U18490 (N_18490,N_18215,N_18117);
xnor U18491 (N_18491,N_18190,N_18020);
nand U18492 (N_18492,N_18242,N_18134);
xnor U18493 (N_18493,N_18109,N_18048);
xor U18494 (N_18494,N_18081,N_18078);
nand U18495 (N_18495,N_18044,N_18243);
xnor U18496 (N_18496,N_18162,N_18219);
nand U18497 (N_18497,N_18192,N_18239);
and U18498 (N_18498,N_18162,N_18232);
and U18499 (N_18499,N_18016,N_18200);
and U18500 (N_18500,N_18358,N_18487);
and U18501 (N_18501,N_18496,N_18267);
or U18502 (N_18502,N_18284,N_18339);
nor U18503 (N_18503,N_18326,N_18415);
or U18504 (N_18504,N_18497,N_18413);
nor U18505 (N_18505,N_18256,N_18430);
xor U18506 (N_18506,N_18416,N_18417);
nor U18507 (N_18507,N_18436,N_18325);
or U18508 (N_18508,N_18404,N_18359);
nand U18509 (N_18509,N_18376,N_18384);
xor U18510 (N_18510,N_18274,N_18362);
and U18511 (N_18511,N_18289,N_18288);
and U18512 (N_18512,N_18466,N_18319);
xnor U18513 (N_18513,N_18484,N_18476);
nor U18514 (N_18514,N_18489,N_18382);
xor U18515 (N_18515,N_18486,N_18491);
nor U18516 (N_18516,N_18409,N_18258);
and U18517 (N_18517,N_18260,N_18440);
nor U18518 (N_18518,N_18381,N_18403);
or U18519 (N_18519,N_18266,N_18261);
or U18520 (N_18520,N_18482,N_18311);
or U18521 (N_18521,N_18451,N_18493);
and U18522 (N_18522,N_18407,N_18360);
nor U18523 (N_18523,N_18469,N_18297);
xor U18524 (N_18524,N_18460,N_18471);
and U18525 (N_18525,N_18342,N_18270);
and U18526 (N_18526,N_18324,N_18265);
xnor U18527 (N_18527,N_18328,N_18456);
or U18528 (N_18528,N_18470,N_18463);
nand U18529 (N_18529,N_18299,N_18278);
nor U18530 (N_18530,N_18405,N_18457);
and U18531 (N_18531,N_18475,N_18301);
and U18532 (N_18532,N_18309,N_18313);
and U18533 (N_18533,N_18315,N_18250);
nor U18534 (N_18534,N_18492,N_18353);
nor U18535 (N_18535,N_18485,N_18383);
nand U18536 (N_18536,N_18488,N_18408);
nor U18537 (N_18537,N_18448,N_18426);
nand U18538 (N_18538,N_18418,N_18435);
xnor U18539 (N_18539,N_18346,N_18264);
and U18540 (N_18540,N_18402,N_18386);
or U18541 (N_18541,N_18272,N_18356);
xnor U18542 (N_18542,N_18401,N_18442);
or U18543 (N_18543,N_18262,N_18318);
xor U18544 (N_18544,N_18352,N_18411);
nand U18545 (N_18545,N_18254,N_18429);
or U18546 (N_18546,N_18290,N_18255);
nand U18547 (N_18547,N_18479,N_18434);
xnor U18548 (N_18548,N_18349,N_18465);
xnor U18549 (N_18549,N_18433,N_18388);
nand U18550 (N_18550,N_18375,N_18277);
nor U18551 (N_18551,N_18312,N_18444);
or U18552 (N_18552,N_18344,N_18459);
xnor U18553 (N_18553,N_18354,N_18276);
and U18554 (N_18554,N_18423,N_18377);
xor U18555 (N_18555,N_18387,N_18334);
nor U18556 (N_18556,N_18296,N_18287);
and U18557 (N_18557,N_18347,N_18425);
or U18558 (N_18558,N_18410,N_18464);
xor U18559 (N_18559,N_18281,N_18490);
xor U18560 (N_18560,N_18333,N_18330);
xnor U18561 (N_18561,N_18379,N_18253);
and U18562 (N_18562,N_18365,N_18472);
nand U18563 (N_18563,N_18302,N_18291);
or U18564 (N_18564,N_18378,N_18268);
and U18565 (N_18565,N_18280,N_18391);
xor U18566 (N_18566,N_18380,N_18259);
xnor U18567 (N_18567,N_18398,N_18419);
xor U18568 (N_18568,N_18480,N_18364);
and U18569 (N_18569,N_18420,N_18498);
nor U18570 (N_18570,N_18340,N_18283);
nor U18571 (N_18571,N_18390,N_18366);
nand U18572 (N_18572,N_18298,N_18369);
or U18573 (N_18573,N_18371,N_18368);
or U18574 (N_18574,N_18337,N_18343);
xnor U18575 (N_18575,N_18447,N_18305);
nand U18576 (N_18576,N_18495,N_18316);
nor U18577 (N_18577,N_18428,N_18449);
or U18578 (N_18578,N_18361,N_18292);
nand U18579 (N_18579,N_18374,N_18452);
nand U18580 (N_18580,N_18461,N_18396);
nand U18581 (N_18581,N_18443,N_18373);
nor U18582 (N_18582,N_18300,N_18348);
nor U18583 (N_18583,N_18307,N_18450);
nand U18584 (N_18584,N_18252,N_18345);
and U18585 (N_18585,N_18439,N_18320);
or U18586 (N_18586,N_18453,N_18412);
nand U18587 (N_18587,N_18427,N_18329);
nor U18588 (N_18588,N_18474,N_18458);
nor U18589 (N_18589,N_18257,N_18494);
nor U18590 (N_18590,N_18269,N_18392);
and U18591 (N_18591,N_18441,N_18400);
and U18592 (N_18592,N_18273,N_18473);
and U18593 (N_18593,N_18338,N_18357);
nand U18594 (N_18594,N_18414,N_18306);
nor U18595 (N_18595,N_18483,N_18394);
nor U18596 (N_18596,N_18295,N_18437);
nor U18597 (N_18597,N_18455,N_18421);
and U18598 (N_18598,N_18341,N_18308);
nor U18599 (N_18599,N_18336,N_18335);
xnor U18600 (N_18600,N_18293,N_18355);
nand U18601 (N_18601,N_18323,N_18454);
nand U18602 (N_18602,N_18331,N_18351);
and U18603 (N_18603,N_18395,N_18317);
xor U18604 (N_18604,N_18431,N_18468);
xor U18605 (N_18605,N_18251,N_18406);
nor U18606 (N_18606,N_18310,N_18399);
xor U18607 (N_18607,N_18322,N_18422);
nor U18608 (N_18608,N_18350,N_18314);
nor U18609 (N_18609,N_18424,N_18499);
or U18610 (N_18610,N_18321,N_18478);
xnor U18611 (N_18611,N_18389,N_18332);
or U18612 (N_18612,N_18385,N_18363);
xnor U18613 (N_18613,N_18367,N_18393);
xor U18614 (N_18614,N_18477,N_18467);
or U18615 (N_18615,N_18263,N_18304);
and U18616 (N_18616,N_18327,N_18285);
nor U18617 (N_18617,N_18294,N_18303);
nand U18618 (N_18618,N_18446,N_18438);
and U18619 (N_18619,N_18279,N_18370);
nand U18620 (N_18620,N_18462,N_18481);
xor U18621 (N_18621,N_18271,N_18445);
xnor U18622 (N_18622,N_18282,N_18275);
and U18623 (N_18623,N_18432,N_18286);
or U18624 (N_18624,N_18397,N_18372);
nand U18625 (N_18625,N_18353,N_18419);
or U18626 (N_18626,N_18345,N_18377);
xnor U18627 (N_18627,N_18440,N_18360);
xnor U18628 (N_18628,N_18260,N_18435);
nand U18629 (N_18629,N_18490,N_18437);
and U18630 (N_18630,N_18420,N_18443);
nand U18631 (N_18631,N_18263,N_18483);
xor U18632 (N_18632,N_18428,N_18276);
nand U18633 (N_18633,N_18276,N_18259);
and U18634 (N_18634,N_18362,N_18407);
nand U18635 (N_18635,N_18444,N_18384);
nand U18636 (N_18636,N_18391,N_18423);
and U18637 (N_18637,N_18264,N_18498);
or U18638 (N_18638,N_18424,N_18494);
and U18639 (N_18639,N_18278,N_18437);
nand U18640 (N_18640,N_18470,N_18384);
nor U18641 (N_18641,N_18431,N_18317);
xor U18642 (N_18642,N_18467,N_18361);
or U18643 (N_18643,N_18259,N_18274);
or U18644 (N_18644,N_18361,N_18497);
nor U18645 (N_18645,N_18348,N_18312);
or U18646 (N_18646,N_18357,N_18459);
nand U18647 (N_18647,N_18409,N_18306);
nor U18648 (N_18648,N_18253,N_18426);
nor U18649 (N_18649,N_18489,N_18452);
and U18650 (N_18650,N_18428,N_18479);
xnor U18651 (N_18651,N_18405,N_18451);
xnor U18652 (N_18652,N_18479,N_18350);
xor U18653 (N_18653,N_18408,N_18485);
and U18654 (N_18654,N_18351,N_18265);
nand U18655 (N_18655,N_18374,N_18414);
xnor U18656 (N_18656,N_18314,N_18475);
and U18657 (N_18657,N_18414,N_18321);
nand U18658 (N_18658,N_18267,N_18452);
xor U18659 (N_18659,N_18437,N_18487);
xor U18660 (N_18660,N_18488,N_18324);
or U18661 (N_18661,N_18383,N_18487);
nand U18662 (N_18662,N_18300,N_18469);
or U18663 (N_18663,N_18329,N_18467);
and U18664 (N_18664,N_18444,N_18264);
or U18665 (N_18665,N_18479,N_18302);
and U18666 (N_18666,N_18323,N_18499);
nand U18667 (N_18667,N_18433,N_18269);
or U18668 (N_18668,N_18327,N_18326);
and U18669 (N_18669,N_18438,N_18348);
nor U18670 (N_18670,N_18412,N_18423);
xor U18671 (N_18671,N_18356,N_18492);
xor U18672 (N_18672,N_18371,N_18288);
xor U18673 (N_18673,N_18482,N_18456);
nor U18674 (N_18674,N_18283,N_18499);
nand U18675 (N_18675,N_18441,N_18454);
nand U18676 (N_18676,N_18448,N_18353);
and U18677 (N_18677,N_18345,N_18259);
or U18678 (N_18678,N_18297,N_18375);
xnor U18679 (N_18679,N_18493,N_18276);
xnor U18680 (N_18680,N_18355,N_18390);
and U18681 (N_18681,N_18395,N_18418);
xor U18682 (N_18682,N_18365,N_18321);
xnor U18683 (N_18683,N_18258,N_18330);
xor U18684 (N_18684,N_18365,N_18302);
xnor U18685 (N_18685,N_18328,N_18387);
nor U18686 (N_18686,N_18471,N_18401);
and U18687 (N_18687,N_18344,N_18309);
or U18688 (N_18688,N_18470,N_18267);
or U18689 (N_18689,N_18407,N_18253);
or U18690 (N_18690,N_18333,N_18487);
or U18691 (N_18691,N_18368,N_18444);
xor U18692 (N_18692,N_18425,N_18270);
xor U18693 (N_18693,N_18371,N_18344);
xnor U18694 (N_18694,N_18379,N_18410);
xnor U18695 (N_18695,N_18314,N_18445);
and U18696 (N_18696,N_18365,N_18382);
and U18697 (N_18697,N_18294,N_18250);
or U18698 (N_18698,N_18341,N_18299);
xor U18699 (N_18699,N_18391,N_18394);
nand U18700 (N_18700,N_18496,N_18260);
xnor U18701 (N_18701,N_18397,N_18421);
xnor U18702 (N_18702,N_18450,N_18261);
nor U18703 (N_18703,N_18257,N_18288);
or U18704 (N_18704,N_18485,N_18422);
xnor U18705 (N_18705,N_18426,N_18484);
nor U18706 (N_18706,N_18385,N_18486);
xor U18707 (N_18707,N_18450,N_18373);
nor U18708 (N_18708,N_18339,N_18328);
nor U18709 (N_18709,N_18330,N_18316);
and U18710 (N_18710,N_18258,N_18355);
and U18711 (N_18711,N_18469,N_18393);
and U18712 (N_18712,N_18450,N_18455);
nand U18713 (N_18713,N_18278,N_18380);
or U18714 (N_18714,N_18459,N_18278);
or U18715 (N_18715,N_18358,N_18284);
nand U18716 (N_18716,N_18258,N_18349);
nand U18717 (N_18717,N_18265,N_18305);
and U18718 (N_18718,N_18309,N_18311);
nor U18719 (N_18719,N_18251,N_18378);
or U18720 (N_18720,N_18261,N_18325);
or U18721 (N_18721,N_18338,N_18272);
or U18722 (N_18722,N_18299,N_18309);
or U18723 (N_18723,N_18419,N_18497);
and U18724 (N_18724,N_18314,N_18264);
nand U18725 (N_18725,N_18496,N_18392);
and U18726 (N_18726,N_18337,N_18345);
nand U18727 (N_18727,N_18477,N_18256);
nor U18728 (N_18728,N_18401,N_18275);
or U18729 (N_18729,N_18321,N_18474);
or U18730 (N_18730,N_18288,N_18256);
nor U18731 (N_18731,N_18341,N_18431);
nand U18732 (N_18732,N_18331,N_18282);
nor U18733 (N_18733,N_18378,N_18278);
or U18734 (N_18734,N_18416,N_18403);
nand U18735 (N_18735,N_18465,N_18265);
nor U18736 (N_18736,N_18312,N_18441);
xnor U18737 (N_18737,N_18344,N_18393);
nor U18738 (N_18738,N_18394,N_18279);
or U18739 (N_18739,N_18331,N_18361);
xor U18740 (N_18740,N_18433,N_18410);
nor U18741 (N_18741,N_18492,N_18348);
nand U18742 (N_18742,N_18297,N_18270);
xor U18743 (N_18743,N_18426,N_18414);
nand U18744 (N_18744,N_18499,N_18440);
nor U18745 (N_18745,N_18366,N_18313);
xnor U18746 (N_18746,N_18474,N_18455);
and U18747 (N_18747,N_18333,N_18417);
nor U18748 (N_18748,N_18407,N_18455);
or U18749 (N_18749,N_18473,N_18418);
nor U18750 (N_18750,N_18583,N_18541);
xor U18751 (N_18751,N_18510,N_18511);
and U18752 (N_18752,N_18749,N_18545);
or U18753 (N_18753,N_18527,N_18721);
nand U18754 (N_18754,N_18692,N_18648);
or U18755 (N_18755,N_18723,N_18626);
or U18756 (N_18756,N_18575,N_18645);
and U18757 (N_18757,N_18611,N_18730);
nand U18758 (N_18758,N_18675,N_18620);
and U18759 (N_18759,N_18742,N_18514);
nand U18760 (N_18760,N_18549,N_18586);
or U18761 (N_18761,N_18561,N_18665);
and U18762 (N_18762,N_18668,N_18650);
or U18763 (N_18763,N_18555,N_18604);
nor U18764 (N_18764,N_18515,N_18580);
nand U18765 (N_18765,N_18588,N_18568);
and U18766 (N_18766,N_18571,N_18567);
and U18767 (N_18767,N_18554,N_18577);
nand U18768 (N_18768,N_18590,N_18520);
nor U18769 (N_18769,N_18512,N_18735);
and U18770 (N_18770,N_18748,N_18632);
or U18771 (N_18771,N_18625,N_18621);
xnor U18772 (N_18772,N_18582,N_18695);
xnor U18773 (N_18773,N_18722,N_18731);
xnor U18774 (N_18774,N_18635,N_18663);
or U18775 (N_18775,N_18506,N_18534);
or U18776 (N_18776,N_18562,N_18595);
nand U18777 (N_18777,N_18629,N_18741);
nand U18778 (N_18778,N_18740,N_18610);
or U18779 (N_18779,N_18680,N_18696);
and U18780 (N_18780,N_18553,N_18652);
nand U18781 (N_18781,N_18678,N_18523);
nand U18782 (N_18782,N_18596,N_18634);
xnor U18783 (N_18783,N_18603,N_18594);
nand U18784 (N_18784,N_18747,N_18616);
nor U18785 (N_18785,N_18538,N_18533);
nand U18786 (N_18786,N_18711,N_18720);
and U18787 (N_18787,N_18623,N_18737);
xnor U18788 (N_18788,N_18618,N_18684);
nor U18789 (N_18789,N_18671,N_18544);
and U18790 (N_18790,N_18592,N_18513);
nand U18791 (N_18791,N_18507,N_18660);
nand U18792 (N_18792,N_18615,N_18704);
nand U18793 (N_18793,N_18669,N_18727);
or U18794 (N_18794,N_18529,N_18563);
xnor U18795 (N_18795,N_18526,N_18681);
nor U18796 (N_18796,N_18716,N_18698);
nand U18797 (N_18797,N_18589,N_18724);
nor U18798 (N_18798,N_18560,N_18569);
and U18799 (N_18799,N_18733,N_18504);
nand U18800 (N_18800,N_18519,N_18656);
nor U18801 (N_18801,N_18536,N_18729);
nand U18802 (N_18802,N_18518,N_18736);
xnor U18803 (N_18803,N_18734,N_18712);
xor U18804 (N_18804,N_18543,N_18651);
xnor U18805 (N_18805,N_18664,N_18581);
xor U18806 (N_18806,N_18714,N_18593);
and U18807 (N_18807,N_18641,N_18535);
nor U18808 (N_18808,N_18732,N_18591);
and U18809 (N_18809,N_18584,N_18574);
or U18810 (N_18810,N_18700,N_18649);
nor U18811 (N_18811,N_18636,N_18717);
and U18812 (N_18812,N_18646,N_18706);
or U18813 (N_18813,N_18579,N_18532);
xor U18814 (N_18814,N_18710,N_18633);
and U18815 (N_18815,N_18674,N_18631);
or U18816 (N_18816,N_18559,N_18661);
nor U18817 (N_18817,N_18540,N_18556);
xnor U18818 (N_18818,N_18707,N_18701);
and U18819 (N_18819,N_18564,N_18743);
and U18820 (N_18820,N_18531,N_18642);
nor U18821 (N_18821,N_18677,N_18600);
xnor U18822 (N_18822,N_18546,N_18522);
or U18823 (N_18823,N_18597,N_18726);
and U18824 (N_18824,N_18558,N_18551);
nor U18825 (N_18825,N_18718,N_18672);
and U18826 (N_18826,N_18682,N_18637);
xnor U18827 (N_18827,N_18570,N_18690);
or U18828 (N_18828,N_18622,N_18548);
nand U18829 (N_18829,N_18628,N_18517);
and U18830 (N_18830,N_18697,N_18667);
or U18831 (N_18831,N_18508,N_18601);
nand U18832 (N_18832,N_18509,N_18599);
nand U18833 (N_18833,N_18657,N_18606);
nor U18834 (N_18834,N_18576,N_18537);
nand U18835 (N_18835,N_18638,N_18566);
or U18836 (N_18836,N_18687,N_18686);
xnor U18837 (N_18837,N_18525,N_18713);
nand U18838 (N_18838,N_18608,N_18542);
or U18839 (N_18839,N_18524,N_18676);
and U18840 (N_18840,N_18573,N_18502);
or U18841 (N_18841,N_18503,N_18719);
nor U18842 (N_18842,N_18501,N_18688);
xnor U18843 (N_18843,N_18739,N_18539);
nand U18844 (N_18844,N_18557,N_18613);
and U18845 (N_18845,N_18644,N_18528);
xor U18846 (N_18846,N_18679,N_18619);
or U18847 (N_18847,N_18715,N_18630);
xor U18848 (N_18848,N_18516,N_18612);
or U18849 (N_18849,N_18673,N_18550);
and U18850 (N_18850,N_18659,N_18640);
nand U18851 (N_18851,N_18666,N_18702);
and U18852 (N_18852,N_18614,N_18605);
and U18853 (N_18853,N_18552,N_18653);
nor U18854 (N_18854,N_18689,N_18662);
nor U18855 (N_18855,N_18699,N_18685);
and U18856 (N_18856,N_18598,N_18703);
or U18857 (N_18857,N_18607,N_18578);
or U18858 (N_18858,N_18744,N_18643);
nand U18859 (N_18859,N_18530,N_18500);
and U18860 (N_18860,N_18521,N_18617);
xor U18861 (N_18861,N_18705,N_18738);
or U18862 (N_18862,N_18639,N_18654);
or U18863 (N_18863,N_18647,N_18572);
and U18864 (N_18864,N_18655,N_18683);
nand U18865 (N_18865,N_18602,N_18728);
and U18866 (N_18866,N_18547,N_18694);
nor U18867 (N_18867,N_18691,N_18587);
xor U18868 (N_18868,N_18624,N_18565);
and U18869 (N_18869,N_18746,N_18693);
or U18870 (N_18870,N_18709,N_18708);
and U18871 (N_18871,N_18658,N_18505);
xnor U18872 (N_18872,N_18585,N_18745);
xor U18873 (N_18873,N_18725,N_18609);
nand U18874 (N_18874,N_18670,N_18627);
xnor U18875 (N_18875,N_18606,N_18520);
or U18876 (N_18876,N_18734,N_18583);
xor U18877 (N_18877,N_18673,N_18660);
nand U18878 (N_18878,N_18587,N_18748);
nand U18879 (N_18879,N_18672,N_18710);
or U18880 (N_18880,N_18575,N_18559);
or U18881 (N_18881,N_18503,N_18591);
xnor U18882 (N_18882,N_18674,N_18569);
nand U18883 (N_18883,N_18535,N_18613);
and U18884 (N_18884,N_18657,N_18647);
and U18885 (N_18885,N_18590,N_18730);
nor U18886 (N_18886,N_18709,N_18724);
nand U18887 (N_18887,N_18558,N_18500);
nor U18888 (N_18888,N_18746,N_18708);
xnor U18889 (N_18889,N_18688,N_18733);
xnor U18890 (N_18890,N_18735,N_18720);
nand U18891 (N_18891,N_18532,N_18502);
and U18892 (N_18892,N_18579,N_18593);
xnor U18893 (N_18893,N_18661,N_18639);
or U18894 (N_18894,N_18640,N_18639);
and U18895 (N_18895,N_18501,N_18723);
and U18896 (N_18896,N_18743,N_18574);
nand U18897 (N_18897,N_18537,N_18583);
and U18898 (N_18898,N_18693,N_18608);
or U18899 (N_18899,N_18590,N_18648);
nor U18900 (N_18900,N_18659,N_18690);
or U18901 (N_18901,N_18512,N_18623);
xnor U18902 (N_18902,N_18558,N_18709);
and U18903 (N_18903,N_18626,N_18622);
nand U18904 (N_18904,N_18549,N_18654);
nand U18905 (N_18905,N_18637,N_18573);
nand U18906 (N_18906,N_18622,N_18697);
xnor U18907 (N_18907,N_18638,N_18654);
nor U18908 (N_18908,N_18573,N_18748);
nor U18909 (N_18909,N_18637,N_18749);
and U18910 (N_18910,N_18724,N_18516);
nor U18911 (N_18911,N_18677,N_18521);
or U18912 (N_18912,N_18745,N_18556);
nor U18913 (N_18913,N_18581,N_18740);
nand U18914 (N_18914,N_18616,N_18523);
nand U18915 (N_18915,N_18731,N_18568);
and U18916 (N_18916,N_18635,N_18514);
xor U18917 (N_18917,N_18570,N_18667);
or U18918 (N_18918,N_18646,N_18662);
nand U18919 (N_18919,N_18515,N_18641);
nand U18920 (N_18920,N_18582,N_18663);
and U18921 (N_18921,N_18573,N_18575);
xor U18922 (N_18922,N_18689,N_18567);
xor U18923 (N_18923,N_18669,N_18668);
and U18924 (N_18924,N_18508,N_18628);
xor U18925 (N_18925,N_18566,N_18506);
and U18926 (N_18926,N_18686,N_18564);
nand U18927 (N_18927,N_18620,N_18537);
nand U18928 (N_18928,N_18676,N_18532);
nand U18929 (N_18929,N_18739,N_18612);
xnor U18930 (N_18930,N_18728,N_18633);
xnor U18931 (N_18931,N_18698,N_18731);
and U18932 (N_18932,N_18745,N_18661);
nand U18933 (N_18933,N_18668,N_18728);
nand U18934 (N_18934,N_18541,N_18595);
or U18935 (N_18935,N_18675,N_18555);
and U18936 (N_18936,N_18624,N_18563);
nand U18937 (N_18937,N_18509,N_18715);
and U18938 (N_18938,N_18540,N_18741);
xor U18939 (N_18939,N_18639,N_18605);
nor U18940 (N_18940,N_18554,N_18592);
nand U18941 (N_18941,N_18735,N_18601);
and U18942 (N_18942,N_18513,N_18621);
or U18943 (N_18943,N_18577,N_18509);
or U18944 (N_18944,N_18736,N_18728);
or U18945 (N_18945,N_18663,N_18638);
nor U18946 (N_18946,N_18571,N_18613);
nand U18947 (N_18947,N_18557,N_18636);
or U18948 (N_18948,N_18691,N_18595);
or U18949 (N_18949,N_18522,N_18636);
or U18950 (N_18950,N_18625,N_18545);
xor U18951 (N_18951,N_18689,N_18686);
nor U18952 (N_18952,N_18585,N_18712);
nor U18953 (N_18953,N_18629,N_18694);
or U18954 (N_18954,N_18561,N_18714);
xor U18955 (N_18955,N_18514,N_18715);
nand U18956 (N_18956,N_18614,N_18747);
nand U18957 (N_18957,N_18562,N_18554);
and U18958 (N_18958,N_18535,N_18520);
xnor U18959 (N_18959,N_18533,N_18613);
nor U18960 (N_18960,N_18688,N_18661);
nand U18961 (N_18961,N_18739,N_18508);
and U18962 (N_18962,N_18677,N_18643);
xor U18963 (N_18963,N_18561,N_18577);
nor U18964 (N_18964,N_18613,N_18516);
nand U18965 (N_18965,N_18689,N_18658);
xnor U18966 (N_18966,N_18616,N_18604);
nand U18967 (N_18967,N_18539,N_18546);
nor U18968 (N_18968,N_18697,N_18602);
or U18969 (N_18969,N_18665,N_18634);
xnor U18970 (N_18970,N_18650,N_18705);
xor U18971 (N_18971,N_18697,N_18677);
or U18972 (N_18972,N_18599,N_18618);
xor U18973 (N_18973,N_18716,N_18645);
nand U18974 (N_18974,N_18650,N_18530);
or U18975 (N_18975,N_18727,N_18716);
and U18976 (N_18976,N_18671,N_18619);
xor U18977 (N_18977,N_18590,N_18530);
or U18978 (N_18978,N_18607,N_18690);
and U18979 (N_18979,N_18639,N_18568);
or U18980 (N_18980,N_18611,N_18674);
xnor U18981 (N_18981,N_18584,N_18705);
and U18982 (N_18982,N_18634,N_18637);
nor U18983 (N_18983,N_18688,N_18740);
and U18984 (N_18984,N_18699,N_18553);
and U18985 (N_18985,N_18625,N_18529);
or U18986 (N_18986,N_18665,N_18647);
and U18987 (N_18987,N_18540,N_18612);
and U18988 (N_18988,N_18684,N_18626);
nor U18989 (N_18989,N_18725,N_18590);
xnor U18990 (N_18990,N_18505,N_18727);
and U18991 (N_18991,N_18529,N_18522);
nand U18992 (N_18992,N_18603,N_18540);
xnor U18993 (N_18993,N_18744,N_18687);
and U18994 (N_18994,N_18676,N_18653);
or U18995 (N_18995,N_18635,N_18685);
nor U18996 (N_18996,N_18644,N_18625);
and U18997 (N_18997,N_18736,N_18606);
xor U18998 (N_18998,N_18523,N_18629);
or U18999 (N_18999,N_18701,N_18723);
xnor U19000 (N_19000,N_18883,N_18810);
and U19001 (N_19001,N_18971,N_18953);
nand U19002 (N_19002,N_18757,N_18928);
or U19003 (N_19003,N_18903,N_18947);
and U19004 (N_19004,N_18997,N_18799);
or U19005 (N_19005,N_18802,N_18864);
and U19006 (N_19006,N_18789,N_18801);
xnor U19007 (N_19007,N_18887,N_18846);
xor U19008 (N_19008,N_18870,N_18929);
nand U19009 (N_19009,N_18845,N_18817);
or U19010 (N_19010,N_18826,N_18995);
nor U19011 (N_19011,N_18835,N_18889);
or U19012 (N_19012,N_18772,N_18793);
xor U19013 (N_19013,N_18879,N_18967);
nor U19014 (N_19014,N_18920,N_18898);
nor U19015 (N_19015,N_18976,N_18983);
xnor U19016 (N_19016,N_18834,N_18798);
xnor U19017 (N_19017,N_18923,N_18950);
nor U19018 (N_19018,N_18999,N_18972);
or U19019 (N_19019,N_18814,N_18838);
and U19020 (N_19020,N_18832,N_18763);
nor U19021 (N_19021,N_18932,N_18811);
xnor U19022 (N_19022,N_18969,N_18818);
nor U19023 (N_19023,N_18994,N_18877);
nor U19024 (N_19024,N_18911,N_18904);
or U19025 (N_19025,N_18998,N_18958);
nand U19026 (N_19026,N_18952,N_18823);
or U19027 (N_19027,N_18852,N_18984);
and U19028 (N_19028,N_18987,N_18899);
xor U19029 (N_19029,N_18865,N_18780);
xnor U19030 (N_19030,N_18821,N_18931);
xnor U19031 (N_19031,N_18943,N_18848);
nor U19032 (N_19032,N_18766,N_18769);
xnor U19033 (N_19033,N_18996,N_18888);
nand U19034 (N_19034,N_18840,N_18890);
nor U19035 (N_19035,N_18939,N_18886);
or U19036 (N_19036,N_18918,N_18804);
nor U19037 (N_19037,N_18849,N_18800);
nor U19038 (N_19038,N_18940,N_18963);
or U19039 (N_19039,N_18831,N_18820);
nand U19040 (N_19040,N_18839,N_18938);
nand U19041 (N_19041,N_18988,N_18842);
nor U19042 (N_19042,N_18768,N_18841);
xor U19043 (N_19043,N_18776,N_18822);
nand U19044 (N_19044,N_18854,N_18782);
nand U19045 (N_19045,N_18990,N_18765);
nand U19046 (N_19046,N_18751,N_18773);
xnor U19047 (N_19047,N_18993,N_18827);
xnor U19048 (N_19048,N_18921,N_18863);
and U19049 (N_19049,N_18790,N_18975);
nor U19050 (N_19050,N_18753,N_18891);
nor U19051 (N_19051,N_18926,N_18964);
xor U19052 (N_19052,N_18901,N_18942);
and U19053 (N_19053,N_18833,N_18853);
nand U19054 (N_19054,N_18896,N_18760);
or U19055 (N_19055,N_18869,N_18795);
or U19056 (N_19056,N_18770,N_18927);
or U19057 (N_19057,N_18992,N_18837);
or U19058 (N_19058,N_18978,N_18847);
and U19059 (N_19059,N_18933,N_18968);
nand U19060 (N_19060,N_18755,N_18881);
or U19061 (N_19061,N_18915,N_18961);
xor U19062 (N_19062,N_18989,N_18862);
xor U19063 (N_19063,N_18778,N_18917);
nor U19064 (N_19064,N_18924,N_18761);
xor U19065 (N_19065,N_18794,N_18966);
or U19066 (N_19066,N_18944,N_18791);
and U19067 (N_19067,N_18949,N_18985);
nor U19068 (N_19068,N_18764,N_18872);
xnor U19069 (N_19069,N_18959,N_18752);
or U19070 (N_19070,N_18851,N_18874);
or U19071 (N_19071,N_18829,N_18965);
or U19072 (N_19072,N_18797,N_18981);
nor U19073 (N_19073,N_18905,N_18819);
or U19074 (N_19074,N_18914,N_18775);
xnor U19075 (N_19075,N_18805,N_18785);
nand U19076 (N_19076,N_18876,N_18912);
xnor U19077 (N_19077,N_18957,N_18930);
and U19078 (N_19078,N_18784,N_18759);
or U19079 (N_19079,N_18808,N_18825);
xnor U19080 (N_19080,N_18894,N_18777);
xor U19081 (N_19081,N_18910,N_18960);
or U19082 (N_19082,N_18945,N_18856);
xnor U19083 (N_19083,N_18936,N_18908);
and U19084 (N_19084,N_18884,N_18878);
xnor U19085 (N_19085,N_18935,N_18902);
nor U19086 (N_19086,N_18892,N_18774);
and U19087 (N_19087,N_18974,N_18844);
xor U19088 (N_19088,N_18803,N_18781);
xor U19089 (N_19089,N_18893,N_18962);
nand U19090 (N_19090,N_18900,N_18867);
nor U19091 (N_19091,N_18855,N_18948);
xnor U19092 (N_19092,N_18828,N_18812);
nor U19093 (N_19093,N_18946,N_18758);
nor U19094 (N_19094,N_18913,N_18934);
nand U19095 (N_19095,N_18792,N_18980);
and U19096 (N_19096,N_18859,N_18941);
or U19097 (N_19097,N_18991,N_18880);
and U19098 (N_19098,N_18875,N_18788);
and U19099 (N_19099,N_18809,N_18925);
or U19100 (N_19100,N_18882,N_18807);
nor U19101 (N_19101,N_18750,N_18857);
or U19102 (N_19102,N_18895,N_18850);
nand U19103 (N_19103,N_18871,N_18906);
or U19104 (N_19104,N_18771,N_18786);
xnor U19105 (N_19105,N_18813,N_18815);
or U19106 (N_19106,N_18922,N_18973);
nor U19107 (N_19107,N_18954,N_18982);
and U19108 (N_19108,N_18783,N_18956);
nand U19109 (N_19109,N_18885,N_18909);
or U19110 (N_19110,N_18860,N_18779);
xor U19111 (N_19111,N_18897,N_18868);
and U19112 (N_19112,N_18843,N_18977);
and U19113 (N_19113,N_18907,N_18787);
and U19114 (N_19114,N_18951,N_18873);
nand U19115 (N_19115,N_18767,N_18866);
nand U19116 (N_19116,N_18979,N_18916);
nor U19117 (N_19117,N_18970,N_18937);
or U19118 (N_19118,N_18816,N_18861);
nand U19119 (N_19119,N_18955,N_18754);
xor U19120 (N_19120,N_18986,N_18919);
or U19121 (N_19121,N_18830,N_18806);
nand U19122 (N_19122,N_18858,N_18836);
or U19123 (N_19123,N_18756,N_18824);
nor U19124 (N_19124,N_18762,N_18796);
and U19125 (N_19125,N_18929,N_18960);
nor U19126 (N_19126,N_18960,N_18875);
or U19127 (N_19127,N_18970,N_18843);
and U19128 (N_19128,N_18957,N_18880);
xnor U19129 (N_19129,N_18913,N_18953);
xor U19130 (N_19130,N_18951,N_18967);
nand U19131 (N_19131,N_18879,N_18759);
nand U19132 (N_19132,N_18911,N_18881);
or U19133 (N_19133,N_18834,N_18870);
xnor U19134 (N_19134,N_18845,N_18789);
xnor U19135 (N_19135,N_18883,N_18808);
or U19136 (N_19136,N_18889,N_18866);
and U19137 (N_19137,N_18999,N_18931);
or U19138 (N_19138,N_18860,N_18820);
nor U19139 (N_19139,N_18846,N_18787);
and U19140 (N_19140,N_18972,N_18787);
and U19141 (N_19141,N_18792,N_18788);
or U19142 (N_19142,N_18924,N_18838);
xor U19143 (N_19143,N_18977,N_18751);
and U19144 (N_19144,N_18897,N_18976);
or U19145 (N_19145,N_18838,N_18808);
and U19146 (N_19146,N_18821,N_18809);
and U19147 (N_19147,N_18753,N_18883);
or U19148 (N_19148,N_18780,N_18766);
or U19149 (N_19149,N_18892,N_18924);
nand U19150 (N_19150,N_18986,N_18964);
nor U19151 (N_19151,N_18753,N_18942);
nor U19152 (N_19152,N_18993,N_18825);
or U19153 (N_19153,N_18978,N_18852);
nor U19154 (N_19154,N_18858,N_18781);
nand U19155 (N_19155,N_18785,N_18883);
or U19156 (N_19156,N_18756,N_18985);
nand U19157 (N_19157,N_18779,N_18831);
or U19158 (N_19158,N_18917,N_18755);
or U19159 (N_19159,N_18914,N_18968);
and U19160 (N_19160,N_18828,N_18974);
nor U19161 (N_19161,N_18935,N_18774);
nor U19162 (N_19162,N_18811,N_18854);
or U19163 (N_19163,N_18758,N_18854);
and U19164 (N_19164,N_18848,N_18809);
nand U19165 (N_19165,N_18938,N_18900);
nor U19166 (N_19166,N_18828,N_18770);
nor U19167 (N_19167,N_18920,N_18973);
nor U19168 (N_19168,N_18972,N_18934);
xnor U19169 (N_19169,N_18872,N_18769);
nor U19170 (N_19170,N_18953,N_18851);
nor U19171 (N_19171,N_18936,N_18780);
or U19172 (N_19172,N_18865,N_18933);
xor U19173 (N_19173,N_18844,N_18874);
nand U19174 (N_19174,N_18915,N_18767);
nor U19175 (N_19175,N_18871,N_18883);
xnor U19176 (N_19176,N_18857,N_18920);
nor U19177 (N_19177,N_18860,N_18923);
or U19178 (N_19178,N_18826,N_18863);
and U19179 (N_19179,N_18934,N_18908);
nand U19180 (N_19180,N_18865,N_18775);
nand U19181 (N_19181,N_18839,N_18969);
xnor U19182 (N_19182,N_18766,N_18835);
and U19183 (N_19183,N_18991,N_18940);
nand U19184 (N_19184,N_18755,N_18920);
or U19185 (N_19185,N_18960,N_18897);
nor U19186 (N_19186,N_18823,N_18888);
and U19187 (N_19187,N_18768,N_18884);
nor U19188 (N_19188,N_18945,N_18952);
nand U19189 (N_19189,N_18989,N_18804);
nor U19190 (N_19190,N_18967,N_18837);
or U19191 (N_19191,N_18995,N_18921);
nand U19192 (N_19192,N_18832,N_18757);
or U19193 (N_19193,N_18818,N_18848);
nor U19194 (N_19194,N_18971,N_18788);
nor U19195 (N_19195,N_18911,N_18897);
nor U19196 (N_19196,N_18910,N_18974);
nor U19197 (N_19197,N_18837,N_18949);
nand U19198 (N_19198,N_18993,N_18883);
xnor U19199 (N_19199,N_18816,N_18932);
xor U19200 (N_19200,N_18884,N_18962);
or U19201 (N_19201,N_18939,N_18771);
or U19202 (N_19202,N_18758,N_18989);
xor U19203 (N_19203,N_18922,N_18945);
nor U19204 (N_19204,N_18769,N_18858);
or U19205 (N_19205,N_18881,N_18772);
or U19206 (N_19206,N_18811,N_18758);
nand U19207 (N_19207,N_18929,N_18764);
or U19208 (N_19208,N_18963,N_18978);
xor U19209 (N_19209,N_18953,N_18918);
and U19210 (N_19210,N_18966,N_18965);
nand U19211 (N_19211,N_18924,N_18952);
xor U19212 (N_19212,N_18971,N_18765);
or U19213 (N_19213,N_18849,N_18835);
nor U19214 (N_19214,N_18933,N_18973);
nor U19215 (N_19215,N_18898,N_18916);
and U19216 (N_19216,N_18786,N_18893);
xnor U19217 (N_19217,N_18874,N_18993);
or U19218 (N_19218,N_18908,N_18983);
nand U19219 (N_19219,N_18806,N_18948);
xnor U19220 (N_19220,N_18964,N_18827);
or U19221 (N_19221,N_18942,N_18807);
nand U19222 (N_19222,N_18982,N_18770);
nand U19223 (N_19223,N_18977,N_18877);
and U19224 (N_19224,N_18988,N_18954);
xnor U19225 (N_19225,N_18947,N_18803);
nor U19226 (N_19226,N_18823,N_18926);
or U19227 (N_19227,N_18956,N_18820);
xnor U19228 (N_19228,N_18987,N_18773);
xor U19229 (N_19229,N_18912,N_18880);
xor U19230 (N_19230,N_18911,N_18808);
nand U19231 (N_19231,N_18851,N_18830);
nor U19232 (N_19232,N_18958,N_18876);
or U19233 (N_19233,N_18763,N_18897);
xor U19234 (N_19234,N_18897,N_18861);
nor U19235 (N_19235,N_18903,N_18783);
nor U19236 (N_19236,N_18936,N_18769);
and U19237 (N_19237,N_18878,N_18860);
nor U19238 (N_19238,N_18772,N_18788);
nand U19239 (N_19239,N_18932,N_18795);
nand U19240 (N_19240,N_18930,N_18995);
or U19241 (N_19241,N_18800,N_18898);
and U19242 (N_19242,N_18996,N_18928);
nand U19243 (N_19243,N_18954,N_18899);
or U19244 (N_19244,N_18946,N_18831);
nand U19245 (N_19245,N_18958,N_18783);
xor U19246 (N_19246,N_18866,N_18968);
xor U19247 (N_19247,N_18973,N_18838);
or U19248 (N_19248,N_18989,N_18974);
and U19249 (N_19249,N_18984,N_18961);
and U19250 (N_19250,N_19058,N_19223);
or U19251 (N_19251,N_19104,N_19222);
nand U19252 (N_19252,N_19081,N_19126);
nand U19253 (N_19253,N_19216,N_19097);
nor U19254 (N_19254,N_19240,N_19162);
or U19255 (N_19255,N_19008,N_19110);
xor U19256 (N_19256,N_19027,N_19115);
or U19257 (N_19257,N_19070,N_19158);
nor U19258 (N_19258,N_19225,N_19049);
or U19259 (N_19259,N_19221,N_19028);
and U19260 (N_19260,N_19085,N_19201);
nor U19261 (N_19261,N_19154,N_19103);
nand U19262 (N_19262,N_19005,N_19146);
xnor U19263 (N_19263,N_19203,N_19247);
and U19264 (N_19264,N_19161,N_19117);
nand U19265 (N_19265,N_19093,N_19025);
and U19266 (N_19266,N_19013,N_19129);
or U19267 (N_19267,N_19205,N_19003);
nor U19268 (N_19268,N_19077,N_19113);
xor U19269 (N_19269,N_19140,N_19194);
nand U19270 (N_19270,N_19053,N_19060);
and U19271 (N_19271,N_19121,N_19030);
nor U19272 (N_19272,N_19153,N_19232);
or U19273 (N_19273,N_19213,N_19196);
or U19274 (N_19274,N_19209,N_19190);
and U19275 (N_19275,N_19174,N_19242);
nor U19276 (N_19276,N_19214,N_19165);
and U19277 (N_19277,N_19130,N_19208);
or U19278 (N_19278,N_19197,N_19160);
xor U19279 (N_19279,N_19017,N_19220);
or U19280 (N_19280,N_19148,N_19163);
xnor U19281 (N_19281,N_19012,N_19187);
nand U19282 (N_19282,N_19231,N_19050);
nor U19283 (N_19283,N_19075,N_19212);
and U19284 (N_19284,N_19227,N_19082);
nor U19285 (N_19285,N_19037,N_19135);
nor U19286 (N_19286,N_19167,N_19061);
nor U19287 (N_19287,N_19238,N_19177);
nor U19288 (N_19288,N_19079,N_19229);
nand U19289 (N_19289,N_19006,N_19001);
nand U19290 (N_19290,N_19226,N_19087);
nor U19291 (N_19291,N_19096,N_19189);
xor U19292 (N_19292,N_19084,N_19233);
nand U19293 (N_19293,N_19074,N_19172);
or U19294 (N_19294,N_19132,N_19092);
xnor U19295 (N_19295,N_19032,N_19236);
xnor U19296 (N_19296,N_19109,N_19199);
nand U19297 (N_19297,N_19106,N_19241);
xor U19298 (N_19298,N_19243,N_19180);
and U19299 (N_19299,N_19059,N_19054);
nand U19300 (N_19300,N_19175,N_19184);
or U19301 (N_19301,N_19064,N_19206);
xor U19302 (N_19302,N_19089,N_19157);
nand U19303 (N_19303,N_19105,N_19086);
nand U19304 (N_19304,N_19088,N_19218);
nor U19305 (N_19305,N_19038,N_19234);
nand U19306 (N_19306,N_19024,N_19185);
and U19307 (N_19307,N_19246,N_19048);
nand U19308 (N_19308,N_19090,N_19239);
or U19309 (N_19309,N_19098,N_19188);
nand U19310 (N_19310,N_19034,N_19202);
xnor U19311 (N_19311,N_19021,N_19237);
or U19312 (N_19312,N_19128,N_19230);
or U19313 (N_19313,N_19124,N_19036);
xnor U19314 (N_19314,N_19009,N_19022);
nand U19315 (N_19315,N_19011,N_19156);
xor U19316 (N_19316,N_19219,N_19072);
or U19317 (N_19317,N_19091,N_19111);
or U19318 (N_19318,N_19136,N_19108);
xor U19319 (N_19319,N_19083,N_19047);
nor U19320 (N_19320,N_19080,N_19004);
nand U19321 (N_19321,N_19198,N_19204);
xnor U19322 (N_19322,N_19186,N_19051);
and U19323 (N_19323,N_19137,N_19014);
nand U19324 (N_19324,N_19062,N_19195);
and U19325 (N_19325,N_19041,N_19057);
and U19326 (N_19326,N_19122,N_19141);
xnor U19327 (N_19327,N_19248,N_19245);
nor U19328 (N_19328,N_19018,N_19071);
or U19329 (N_19329,N_19023,N_19033);
nor U19330 (N_19330,N_19235,N_19120);
nand U19331 (N_19331,N_19191,N_19138);
xor U19332 (N_19332,N_19010,N_19101);
xor U19333 (N_19333,N_19144,N_19176);
xnor U19334 (N_19334,N_19002,N_19015);
nor U19335 (N_19335,N_19200,N_19042);
xor U19336 (N_19336,N_19149,N_19169);
and U19337 (N_19337,N_19249,N_19078);
nor U19338 (N_19338,N_19094,N_19244);
nand U19339 (N_19339,N_19118,N_19007);
nor U19340 (N_19340,N_19112,N_19065);
or U19341 (N_19341,N_19147,N_19166);
or U19342 (N_19342,N_19178,N_19073);
or U19343 (N_19343,N_19170,N_19139);
nand U19344 (N_19344,N_19134,N_19045);
or U19345 (N_19345,N_19133,N_19182);
nand U19346 (N_19346,N_19211,N_19164);
and U19347 (N_19347,N_19044,N_19020);
or U19348 (N_19348,N_19179,N_19107);
and U19349 (N_19349,N_19100,N_19046);
nor U19350 (N_19350,N_19102,N_19040);
nand U19351 (N_19351,N_19039,N_19035);
xnor U19352 (N_19352,N_19055,N_19114);
or U19353 (N_19353,N_19183,N_19043);
or U19354 (N_19354,N_19207,N_19069);
nand U19355 (N_19355,N_19068,N_19142);
or U19356 (N_19356,N_19143,N_19152);
and U19357 (N_19357,N_19215,N_19159);
xnor U19358 (N_19358,N_19063,N_19168);
nor U19359 (N_19359,N_19145,N_19125);
or U19360 (N_19360,N_19095,N_19016);
or U19361 (N_19361,N_19076,N_19193);
or U19362 (N_19362,N_19066,N_19067);
nor U19363 (N_19363,N_19019,N_19029);
and U19364 (N_19364,N_19099,N_19127);
xnor U19365 (N_19365,N_19131,N_19123);
and U19366 (N_19366,N_19155,N_19056);
nand U19367 (N_19367,N_19052,N_19119);
nand U19368 (N_19368,N_19217,N_19228);
or U19369 (N_19369,N_19000,N_19151);
and U19370 (N_19370,N_19192,N_19224);
and U19371 (N_19371,N_19150,N_19173);
or U19372 (N_19372,N_19026,N_19031);
nor U19373 (N_19373,N_19116,N_19181);
xnor U19374 (N_19374,N_19210,N_19171);
and U19375 (N_19375,N_19076,N_19238);
nand U19376 (N_19376,N_19029,N_19147);
and U19377 (N_19377,N_19226,N_19222);
xor U19378 (N_19378,N_19098,N_19059);
xor U19379 (N_19379,N_19028,N_19225);
nand U19380 (N_19380,N_19121,N_19110);
nor U19381 (N_19381,N_19231,N_19208);
xnor U19382 (N_19382,N_19188,N_19230);
nand U19383 (N_19383,N_19203,N_19210);
nor U19384 (N_19384,N_19113,N_19021);
xnor U19385 (N_19385,N_19194,N_19088);
or U19386 (N_19386,N_19047,N_19219);
nand U19387 (N_19387,N_19031,N_19221);
nor U19388 (N_19388,N_19156,N_19178);
and U19389 (N_19389,N_19003,N_19203);
nor U19390 (N_19390,N_19231,N_19207);
nor U19391 (N_19391,N_19181,N_19029);
and U19392 (N_19392,N_19217,N_19214);
xnor U19393 (N_19393,N_19086,N_19075);
nand U19394 (N_19394,N_19115,N_19243);
nand U19395 (N_19395,N_19179,N_19022);
xnor U19396 (N_19396,N_19003,N_19099);
and U19397 (N_19397,N_19051,N_19016);
and U19398 (N_19398,N_19037,N_19063);
or U19399 (N_19399,N_19041,N_19211);
nor U19400 (N_19400,N_19029,N_19219);
or U19401 (N_19401,N_19164,N_19210);
nor U19402 (N_19402,N_19084,N_19185);
nor U19403 (N_19403,N_19102,N_19041);
xor U19404 (N_19404,N_19103,N_19153);
and U19405 (N_19405,N_19243,N_19098);
nand U19406 (N_19406,N_19073,N_19198);
nand U19407 (N_19407,N_19164,N_19110);
nor U19408 (N_19408,N_19133,N_19059);
nand U19409 (N_19409,N_19069,N_19055);
xnor U19410 (N_19410,N_19175,N_19137);
nand U19411 (N_19411,N_19128,N_19047);
and U19412 (N_19412,N_19059,N_19142);
xnor U19413 (N_19413,N_19068,N_19221);
nand U19414 (N_19414,N_19050,N_19181);
xnor U19415 (N_19415,N_19021,N_19078);
or U19416 (N_19416,N_19082,N_19045);
or U19417 (N_19417,N_19233,N_19079);
or U19418 (N_19418,N_19249,N_19114);
nand U19419 (N_19419,N_19047,N_19151);
nor U19420 (N_19420,N_19145,N_19036);
and U19421 (N_19421,N_19108,N_19081);
nor U19422 (N_19422,N_19188,N_19089);
nand U19423 (N_19423,N_19238,N_19022);
nor U19424 (N_19424,N_19089,N_19224);
or U19425 (N_19425,N_19057,N_19195);
and U19426 (N_19426,N_19043,N_19224);
or U19427 (N_19427,N_19011,N_19031);
xnor U19428 (N_19428,N_19147,N_19009);
nand U19429 (N_19429,N_19027,N_19087);
or U19430 (N_19430,N_19231,N_19085);
nor U19431 (N_19431,N_19205,N_19204);
nand U19432 (N_19432,N_19150,N_19078);
nor U19433 (N_19433,N_19014,N_19152);
and U19434 (N_19434,N_19124,N_19029);
or U19435 (N_19435,N_19034,N_19077);
and U19436 (N_19436,N_19246,N_19003);
nor U19437 (N_19437,N_19084,N_19222);
nand U19438 (N_19438,N_19105,N_19195);
and U19439 (N_19439,N_19217,N_19081);
and U19440 (N_19440,N_19005,N_19049);
nor U19441 (N_19441,N_19187,N_19017);
or U19442 (N_19442,N_19114,N_19196);
and U19443 (N_19443,N_19048,N_19025);
and U19444 (N_19444,N_19073,N_19227);
xor U19445 (N_19445,N_19066,N_19035);
nor U19446 (N_19446,N_19234,N_19114);
nor U19447 (N_19447,N_19086,N_19151);
xnor U19448 (N_19448,N_19013,N_19004);
or U19449 (N_19449,N_19191,N_19004);
nand U19450 (N_19450,N_19027,N_19143);
or U19451 (N_19451,N_19129,N_19206);
xnor U19452 (N_19452,N_19113,N_19133);
nand U19453 (N_19453,N_19100,N_19234);
and U19454 (N_19454,N_19122,N_19239);
nor U19455 (N_19455,N_19063,N_19198);
nand U19456 (N_19456,N_19085,N_19167);
xor U19457 (N_19457,N_19213,N_19199);
nand U19458 (N_19458,N_19026,N_19123);
nor U19459 (N_19459,N_19017,N_19057);
nor U19460 (N_19460,N_19027,N_19101);
nand U19461 (N_19461,N_19152,N_19246);
xor U19462 (N_19462,N_19073,N_19098);
and U19463 (N_19463,N_19221,N_19240);
nor U19464 (N_19464,N_19033,N_19096);
xnor U19465 (N_19465,N_19148,N_19130);
nor U19466 (N_19466,N_19068,N_19025);
xor U19467 (N_19467,N_19046,N_19198);
or U19468 (N_19468,N_19111,N_19212);
nor U19469 (N_19469,N_19055,N_19200);
and U19470 (N_19470,N_19217,N_19182);
or U19471 (N_19471,N_19049,N_19022);
nor U19472 (N_19472,N_19140,N_19052);
or U19473 (N_19473,N_19130,N_19053);
and U19474 (N_19474,N_19245,N_19034);
or U19475 (N_19475,N_19142,N_19185);
or U19476 (N_19476,N_19123,N_19069);
nand U19477 (N_19477,N_19092,N_19000);
nor U19478 (N_19478,N_19121,N_19247);
and U19479 (N_19479,N_19185,N_19226);
and U19480 (N_19480,N_19131,N_19145);
nor U19481 (N_19481,N_19134,N_19070);
or U19482 (N_19482,N_19187,N_19106);
nand U19483 (N_19483,N_19188,N_19209);
or U19484 (N_19484,N_19140,N_19026);
xor U19485 (N_19485,N_19186,N_19199);
nor U19486 (N_19486,N_19097,N_19122);
nand U19487 (N_19487,N_19184,N_19150);
or U19488 (N_19488,N_19120,N_19089);
nand U19489 (N_19489,N_19192,N_19183);
or U19490 (N_19490,N_19197,N_19186);
nand U19491 (N_19491,N_19086,N_19117);
xnor U19492 (N_19492,N_19203,N_19082);
nor U19493 (N_19493,N_19131,N_19167);
or U19494 (N_19494,N_19134,N_19087);
nand U19495 (N_19495,N_19081,N_19033);
xor U19496 (N_19496,N_19136,N_19017);
nor U19497 (N_19497,N_19101,N_19153);
and U19498 (N_19498,N_19160,N_19135);
xnor U19499 (N_19499,N_19162,N_19017);
and U19500 (N_19500,N_19419,N_19277);
nor U19501 (N_19501,N_19487,N_19427);
or U19502 (N_19502,N_19283,N_19269);
xnor U19503 (N_19503,N_19418,N_19420);
nand U19504 (N_19504,N_19356,N_19262);
and U19505 (N_19505,N_19297,N_19441);
xnor U19506 (N_19506,N_19494,N_19351);
and U19507 (N_19507,N_19453,N_19349);
and U19508 (N_19508,N_19443,N_19445);
xnor U19509 (N_19509,N_19478,N_19455);
xor U19510 (N_19510,N_19329,N_19369);
and U19511 (N_19511,N_19339,N_19331);
nor U19512 (N_19512,N_19258,N_19392);
xor U19513 (N_19513,N_19447,N_19401);
xnor U19514 (N_19514,N_19257,N_19300);
nand U19515 (N_19515,N_19379,N_19433);
xor U19516 (N_19516,N_19407,N_19492);
or U19517 (N_19517,N_19322,N_19346);
nand U19518 (N_19518,N_19358,N_19426);
nand U19519 (N_19519,N_19363,N_19411);
and U19520 (N_19520,N_19293,N_19345);
nor U19521 (N_19521,N_19467,N_19298);
nand U19522 (N_19522,N_19348,N_19472);
and U19523 (N_19523,N_19442,N_19308);
nand U19524 (N_19524,N_19384,N_19481);
xnor U19525 (N_19525,N_19250,N_19422);
nand U19526 (N_19526,N_19326,N_19370);
or U19527 (N_19527,N_19458,N_19273);
nor U19528 (N_19528,N_19254,N_19367);
nor U19529 (N_19529,N_19333,N_19284);
or U19530 (N_19530,N_19385,N_19383);
or U19531 (N_19531,N_19495,N_19354);
xnor U19532 (N_19532,N_19275,N_19311);
and U19533 (N_19533,N_19347,N_19464);
xnor U19534 (N_19534,N_19402,N_19394);
or U19535 (N_19535,N_19395,N_19372);
nand U19536 (N_19536,N_19412,N_19266);
or U19537 (N_19537,N_19431,N_19473);
nand U19538 (N_19538,N_19287,N_19475);
xor U19539 (N_19539,N_19360,N_19474);
and U19540 (N_19540,N_19320,N_19336);
xor U19541 (N_19541,N_19373,N_19424);
or U19542 (N_19542,N_19327,N_19406);
and U19543 (N_19543,N_19353,N_19325);
nand U19544 (N_19544,N_19398,N_19310);
or U19545 (N_19545,N_19355,N_19261);
nand U19546 (N_19546,N_19324,N_19342);
xor U19547 (N_19547,N_19461,N_19334);
xnor U19548 (N_19548,N_19299,N_19312);
xnor U19549 (N_19549,N_19439,N_19432);
xor U19550 (N_19550,N_19465,N_19399);
xor U19551 (N_19551,N_19486,N_19425);
nand U19552 (N_19552,N_19255,N_19305);
and U19553 (N_19553,N_19286,N_19251);
nand U19554 (N_19554,N_19476,N_19393);
or U19555 (N_19555,N_19404,N_19276);
nand U19556 (N_19556,N_19289,N_19382);
and U19557 (N_19557,N_19389,N_19253);
and U19558 (N_19558,N_19361,N_19391);
nand U19559 (N_19559,N_19375,N_19341);
and U19560 (N_19560,N_19381,N_19498);
and U19561 (N_19561,N_19491,N_19352);
and U19562 (N_19562,N_19471,N_19405);
xor U19563 (N_19563,N_19479,N_19428);
and U19564 (N_19564,N_19314,N_19301);
and U19565 (N_19565,N_19417,N_19376);
nand U19566 (N_19566,N_19462,N_19499);
nor U19567 (N_19567,N_19414,N_19282);
or U19568 (N_19568,N_19400,N_19350);
nand U19569 (N_19569,N_19252,N_19386);
nor U19570 (N_19570,N_19469,N_19271);
nand U19571 (N_19571,N_19264,N_19430);
nor U19572 (N_19572,N_19456,N_19323);
xor U19573 (N_19573,N_19449,N_19270);
xor U19574 (N_19574,N_19313,N_19489);
xnor U19575 (N_19575,N_19497,N_19484);
and U19576 (N_19576,N_19330,N_19446);
or U19577 (N_19577,N_19396,N_19332);
nor U19578 (N_19578,N_19291,N_19377);
nor U19579 (N_19579,N_19496,N_19304);
or U19580 (N_19580,N_19267,N_19328);
or U19581 (N_19581,N_19468,N_19294);
nand U19582 (N_19582,N_19268,N_19437);
and U19583 (N_19583,N_19480,N_19357);
and U19584 (N_19584,N_19344,N_19317);
nand U19585 (N_19585,N_19337,N_19338);
nor U19586 (N_19586,N_19315,N_19485);
nor U19587 (N_19587,N_19260,N_19272);
or U19588 (N_19588,N_19470,N_19285);
xnor U19589 (N_19589,N_19340,N_19416);
nand U19590 (N_19590,N_19335,N_19454);
or U19591 (N_19591,N_19397,N_19316);
nor U19592 (N_19592,N_19448,N_19483);
nor U19593 (N_19593,N_19278,N_19388);
xnor U19594 (N_19594,N_19477,N_19256);
or U19595 (N_19595,N_19374,N_19364);
or U19596 (N_19596,N_19365,N_19434);
and U19597 (N_19597,N_19290,N_19288);
nor U19598 (N_19598,N_19265,N_19410);
nand U19599 (N_19599,N_19380,N_19281);
xor U19600 (N_19600,N_19415,N_19295);
nand U19601 (N_19601,N_19429,N_19413);
nand U19602 (N_19602,N_19321,N_19451);
nor U19603 (N_19603,N_19343,N_19490);
or U19604 (N_19604,N_19309,N_19459);
xnor U19605 (N_19605,N_19368,N_19318);
nand U19606 (N_19606,N_19452,N_19307);
or U19607 (N_19607,N_19440,N_19296);
nand U19608 (N_19608,N_19435,N_19493);
and U19609 (N_19609,N_19444,N_19423);
nand U19610 (N_19610,N_19306,N_19450);
nor U19611 (N_19611,N_19403,N_19378);
nor U19612 (N_19612,N_19390,N_19460);
and U19613 (N_19613,N_19302,N_19482);
xnor U19614 (N_19614,N_19259,N_19466);
or U19615 (N_19615,N_19438,N_19359);
and U19616 (N_19616,N_19362,N_19457);
or U19617 (N_19617,N_19436,N_19366);
or U19618 (N_19618,N_19463,N_19279);
nand U19619 (N_19619,N_19371,N_19387);
xor U19620 (N_19620,N_19292,N_19274);
and U19621 (N_19621,N_19303,N_19319);
or U19622 (N_19622,N_19280,N_19409);
nand U19623 (N_19623,N_19263,N_19488);
nor U19624 (N_19624,N_19408,N_19421);
nor U19625 (N_19625,N_19366,N_19386);
xnor U19626 (N_19626,N_19463,N_19286);
xnor U19627 (N_19627,N_19431,N_19262);
nand U19628 (N_19628,N_19476,N_19477);
nor U19629 (N_19629,N_19262,N_19355);
and U19630 (N_19630,N_19380,N_19369);
and U19631 (N_19631,N_19348,N_19351);
nor U19632 (N_19632,N_19438,N_19323);
nor U19633 (N_19633,N_19484,N_19466);
xor U19634 (N_19634,N_19262,N_19403);
nor U19635 (N_19635,N_19307,N_19379);
xnor U19636 (N_19636,N_19381,N_19399);
nor U19637 (N_19637,N_19357,N_19379);
or U19638 (N_19638,N_19286,N_19305);
or U19639 (N_19639,N_19273,N_19452);
or U19640 (N_19640,N_19485,N_19368);
xor U19641 (N_19641,N_19416,N_19261);
nor U19642 (N_19642,N_19379,N_19359);
or U19643 (N_19643,N_19360,N_19477);
and U19644 (N_19644,N_19358,N_19449);
nor U19645 (N_19645,N_19315,N_19368);
nor U19646 (N_19646,N_19479,N_19444);
and U19647 (N_19647,N_19366,N_19486);
xnor U19648 (N_19648,N_19466,N_19335);
xnor U19649 (N_19649,N_19331,N_19467);
nor U19650 (N_19650,N_19398,N_19253);
nand U19651 (N_19651,N_19455,N_19322);
nand U19652 (N_19652,N_19374,N_19450);
xor U19653 (N_19653,N_19345,N_19407);
or U19654 (N_19654,N_19261,N_19337);
xor U19655 (N_19655,N_19295,N_19321);
xor U19656 (N_19656,N_19427,N_19286);
or U19657 (N_19657,N_19376,N_19374);
nand U19658 (N_19658,N_19487,N_19300);
and U19659 (N_19659,N_19326,N_19256);
or U19660 (N_19660,N_19499,N_19293);
nand U19661 (N_19661,N_19279,N_19482);
or U19662 (N_19662,N_19430,N_19445);
and U19663 (N_19663,N_19400,N_19326);
xor U19664 (N_19664,N_19417,N_19402);
or U19665 (N_19665,N_19395,N_19493);
xnor U19666 (N_19666,N_19490,N_19339);
nor U19667 (N_19667,N_19302,N_19344);
nor U19668 (N_19668,N_19316,N_19429);
nor U19669 (N_19669,N_19433,N_19317);
nand U19670 (N_19670,N_19321,N_19469);
nand U19671 (N_19671,N_19388,N_19449);
nand U19672 (N_19672,N_19480,N_19391);
xnor U19673 (N_19673,N_19357,N_19395);
nand U19674 (N_19674,N_19373,N_19435);
nor U19675 (N_19675,N_19311,N_19254);
xor U19676 (N_19676,N_19474,N_19257);
or U19677 (N_19677,N_19388,N_19324);
nand U19678 (N_19678,N_19394,N_19484);
xnor U19679 (N_19679,N_19353,N_19404);
or U19680 (N_19680,N_19255,N_19491);
and U19681 (N_19681,N_19389,N_19415);
and U19682 (N_19682,N_19441,N_19478);
or U19683 (N_19683,N_19352,N_19451);
or U19684 (N_19684,N_19290,N_19452);
nand U19685 (N_19685,N_19499,N_19389);
and U19686 (N_19686,N_19381,N_19313);
nand U19687 (N_19687,N_19490,N_19280);
and U19688 (N_19688,N_19300,N_19252);
nor U19689 (N_19689,N_19407,N_19312);
and U19690 (N_19690,N_19453,N_19284);
nor U19691 (N_19691,N_19293,N_19381);
xor U19692 (N_19692,N_19258,N_19496);
and U19693 (N_19693,N_19273,N_19455);
and U19694 (N_19694,N_19345,N_19408);
or U19695 (N_19695,N_19297,N_19490);
and U19696 (N_19696,N_19386,N_19274);
nor U19697 (N_19697,N_19385,N_19323);
xnor U19698 (N_19698,N_19361,N_19312);
xor U19699 (N_19699,N_19482,N_19280);
and U19700 (N_19700,N_19451,N_19442);
xor U19701 (N_19701,N_19282,N_19438);
nand U19702 (N_19702,N_19345,N_19288);
nor U19703 (N_19703,N_19422,N_19303);
nor U19704 (N_19704,N_19491,N_19290);
and U19705 (N_19705,N_19425,N_19386);
or U19706 (N_19706,N_19486,N_19350);
and U19707 (N_19707,N_19328,N_19452);
xor U19708 (N_19708,N_19464,N_19300);
nand U19709 (N_19709,N_19448,N_19387);
xor U19710 (N_19710,N_19412,N_19293);
nand U19711 (N_19711,N_19371,N_19469);
and U19712 (N_19712,N_19478,N_19317);
and U19713 (N_19713,N_19357,N_19261);
nand U19714 (N_19714,N_19470,N_19397);
nor U19715 (N_19715,N_19436,N_19324);
nand U19716 (N_19716,N_19397,N_19369);
nor U19717 (N_19717,N_19464,N_19487);
nor U19718 (N_19718,N_19267,N_19470);
and U19719 (N_19719,N_19272,N_19440);
or U19720 (N_19720,N_19401,N_19288);
nand U19721 (N_19721,N_19436,N_19421);
or U19722 (N_19722,N_19494,N_19261);
nor U19723 (N_19723,N_19420,N_19304);
or U19724 (N_19724,N_19487,N_19407);
nor U19725 (N_19725,N_19438,N_19440);
nand U19726 (N_19726,N_19439,N_19326);
and U19727 (N_19727,N_19335,N_19413);
xnor U19728 (N_19728,N_19370,N_19285);
nand U19729 (N_19729,N_19368,N_19363);
xnor U19730 (N_19730,N_19452,N_19283);
nor U19731 (N_19731,N_19321,N_19423);
or U19732 (N_19732,N_19307,N_19456);
xor U19733 (N_19733,N_19380,N_19461);
and U19734 (N_19734,N_19288,N_19429);
or U19735 (N_19735,N_19388,N_19459);
xor U19736 (N_19736,N_19257,N_19421);
or U19737 (N_19737,N_19376,N_19386);
nor U19738 (N_19738,N_19253,N_19355);
xor U19739 (N_19739,N_19322,N_19268);
nand U19740 (N_19740,N_19295,N_19392);
nor U19741 (N_19741,N_19366,N_19297);
xnor U19742 (N_19742,N_19336,N_19287);
nor U19743 (N_19743,N_19406,N_19268);
and U19744 (N_19744,N_19387,N_19454);
nand U19745 (N_19745,N_19379,N_19358);
and U19746 (N_19746,N_19486,N_19477);
and U19747 (N_19747,N_19459,N_19460);
and U19748 (N_19748,N_19435,N_19269);
and U19749 (N_19749,N_19357,N_19322);
and U19750 (N_19750,N_19512,N_19743);
and U19751 (N_19751,N_19585,N_19688);
or U19752 (N_19752,N_19611,N_19605);
xor U19753 (N_19753,N_19593,N_19599);
nand U19754 (N_19754,N_19625,N_19730);
xor U19755 (N_19755,N_19542,N_19639);
nand U19756 (N_19756,N_19624,N_19604);
or U19757 (N_19757,N_19650,N_19598);
or U19758 (N_19758,N_19551,N_19581);
nand U19759 (N_19759,N_19547,N_19591);
or U19760 (N_19760,N_19642,N_19669);
or U19761 (N_19761,N_19531,N_19519);
xnor U19762 (N_19762,N_19686,N_19541);
and U19763 (N_19763,N_19655,N_19528);
nor U19764 (N_19764,N_19731,N_19539);
nand U19765 (N_19765,N_19631,N_19594);
and U19766 (N_19766,N_19566,N_19746);
and U19767 (N_19767,N_19646,N_19663);
nand U19768 (N_19768,N_19725,N_19678);
nor U19769 (N_19769,N_19535,N_19703);
nor U19770 (N_19770,N_19580,N_19682);
xor U19771 (N_19771,N_19706,N_19608);
xor U19772 (N_19772,N_19576,N_19516);
or U19773 (N_19773,N_19732,N_19737);
or U19774 (N_19774,N_19671,N_19662);
nand U19775 (N_19775,N_19696,N_19677);
nand U19776 (N_19776,N_19514,N_19565);
xnor U19777 (N_19777,N_19652,N_19592);
or U19778 (N_19778,N_19596,N_19569);
nand U19779 (N_19779,N_19672,N_19716);
nand U19780 (N_19780,N_19616,N_19530);
and U19781 (N_19781,N_19659,N_19717);
xor U19782 (N_19782,N_19618,N_19545);
or U19783 (N_19783,N_19649,N_19713);
nor U19784 (N_19784,N_19544,N_19513);
nand U19785 (N_19785,N_19620,N_19546);
nor U19786 (N_19786,N_19634,N_19734);
nor U19787 (N_19787,N_19562,N_19638);
and U19788 (N_19788,N_19644,N_19505);
xor U19789 (N_19789,N_19708,N_19681);
nand U19790 (N_19790,N_19572,N_19670);
or U19791 (N_19791,N_19548,N_19709);
nand U19792 (N_19792,N_19532,N_19691);
or U19793 (N_19793,N_19595,N_19658);
nor U19794 (N_19794,N_19651,N_19582);
nor U19795 (N_19795,N_19578,N_19502);
nor U19796 (N_19796,N_19629,N_19515);
xor U19797 (N_19797,N_19715,N_19522);
or U19798 (N_19798,N_19571,N_19590);
xor U19799 (N_19799,N_19632,N_19720);
nand U19800 (N_19800,N_19729,N_19584);
nor U19801 (N_19801,N_19518,N_19735);
nand U19802 (N_19802,N_19517,N_19614);
nor U19803 (N_19803,N_19603,N_19683);
xor U19804 (N_19804,N_19647,N_19510);
xnor U19805 (N_19805,N_19674,N_19742);
or U19806 (N_19806,N_19586,N_19733);
nor U19807 (N_19807,N_19553,N_19657);
or U19808 (N_19808,N_19719,N_19701);
xnor U19809 (N_19809,N_19570,N_19643);
and U19810 (N_19810,N_19702,N_19692);
nor U19811 (N_19811,N_19741,N_19635);
nand U19812 (N_19812,N_19567,N_19689);
or U19813 (N_19813,N_19648,N_19601);
nand U19814 (N_19814,N_19557,N_19690);
nor U19815 (N_19815,N_19602,N_19685);
xor U19816 (N_19816,N_19588,N_19537);
nor U19817 (N_19817,N_19687,N_19525);
xor U19818 (N_19818,N_19527,N_19558);
xor U19819 (N_19819,N_19587,N_19640);
nor U19820 (N_19820,N_19694,N_19543);
xnor U19821 (N_19821,N_19641,N_19676);
and U19822 (N_19822,N_19549,N_19724);
nand U19823 (N_19823,N_19526,N_19607);
nand U19824 (N_19824,N_19529,N_19501);
xnor U19825 (N_19825,N_19653,N_19597);
nand U19826 (N_19826,N_19728,N_19710);
nand U19827 (N_19827,N_19705,N_19711);
or U19828 (N_19828,N_19656,N_19666);
or U19829 (N_19829,N_19538,N_19628);
xor U19830 (N_19830,N_19577,N_19712);
or U19831 (N_19831,N_19612,N_19606);
nand U19832 (N_19832,N_19660,N_19748);
nor U19833 (N_19833,N_19574,N_19745);
and U19834 (N_19834,N_19697,N_19508);
or U19835 (N_19835,N_19668,N_19739);
nor U19836 (N_19836,N_19667,N_19619);
and U19837 (N_19837,N_19665,N_19573);
or U19838 (N_19838,N_19698,N_19673);
nand U19839 (N_19839,N_19700,N_19507);
or U19840 (N_19840,N_19533,N_19699);
nor U19841 (N_19841,N_19523,N_19500);
xnor U19842 (N_19842,N_19654,N_19622);
nor U19843 (N_19843,N_19600,N_19684);
nor U19844 (N_19844,N_19693,N_19534);
or U19845 (N_19845,N_19661,N_19559);
nor U19846 (N_19846,N_19749,N_19550);
or U19847 (N_19847,N_19718,N_19536);
nand U19848 (N_19848,N_19621,N_19560);
and U19849 (N_19849,N_19579,N_19563);
nand U19850 (N_19850,N_19723,N_19617);
or U19851 (N_19851,N_19583,N_19675);
nor U19852 (N_19852,N_19626,N_19540);
and U19853 (N_19853,N_19589,N_19524);
and U19854 (N_19854,N_19636,N_19554);
nand U19855 (N_19855,N_19727,N_19568);
or U19856 (N_19856,N_19645,N_19726);
xnor U19857 (N_19857,N_19736,N_19503);
nor U19858 (N_19858,N_19609,N_19637);
nor U19859 (N_19859,N_19610,N_19627);
or U19860 (N_19860,N_19561,N_19679);
nand U19861 (N_19861,N_19504,N_19521);
xnor U19862 (N_19862,N_19707,N_19722);
nand U19863 (N_19863,N_19613,N_19564);
nand U19864 (N_19864,N_19511,N_19714);
nor U19865 (N_19865,N_19738,N_19633);
or U19866 (N_19866,N_19630,N_19721);
or U19867 (N_19867,N_19520,N_19695);
nand U19868 (N_19868,N_19680,N_19704);
nor U19869 (N_19869,N_19552,N_19744);
xnor U19870 (N_19870,N_19615,N_19575);
and U19871 (N_19871,N_19623,N_19740);
and U19872 (N_19872,N_19664,N_19509);
and U19873 (N_19873,N_19747,N_19506);
xor U19874 (N_19874,N_19556,N_19555);
or U19875 (N_19875,N_19592,N_19572);
or U19876 (N_19876,N_19689,N_19571);
and U19877 (N_19877,N_19501,N_19583);
xor U19878 (N_19878,N_19532,N_19597);
or U19879 (N_19879,N_19532,N_19533);
xor U19880 (N_19880,N_19501,N_19532);
nor U19881 (N_19881,N_19628,N_19661);
or U19882 (N_19882,N_19563,N_19646);
and U19883 (N_19883,N_19691,N_19720);
nand U19884 (N_19884,N_19678,N_19669);
nand U19885 (N_19885,N_19576,N_19640);
and U19886 (N_19886,N_19669,N_19668);
or U19887 (N_19887,N_19747,N_19566);
or U19888 (N_19888,N_19547,N_19747);
nand U19889 (N_19889,N_19533,N_19688);
or U19890 (N_19890,N_19560,N_19667);
xnor U19891 (N_19891,N_19621,N_19721);
or U19892 (N_19892,N_19685,N_19645);
and U19893 (N_19893,N_19578,N_19518);
nand U19894 (N_19894,N_19690,N_19617);
or U19895 (N_19895,N_19671,N_19716);
and U19896 (N_19896,N_19548,N_19547);
nor U19897 (N_19897,N_19520,N_19542);
nand U19898 (N_19898,N_19600,N_19572);
or U19899 (N_19899,N_19530,N_19665);
xor U19900 (N_19900,N_19734,N_19623);
nand U19901 (N_19901,N_19592,N_19621);
or U19902 (N_19902,N_19633,N_19509);
nor U19903 (N_19903,N_19622,N_19707);
nor U19904 (N_19904,N_19611,N_19720);
and U19905 (N_19905,N_19652,N_19686);
and U19906 (N_19906,N_19527,N_19530);
nand U19907 (N_19907,N_19673,N_19743);
nand U19908 (N_19908,N_19681,N_19616);
or U19909 (N_19909,N_19616,N_19663);
nor U19910 (N_19910,N_19534,N_19639);
nor U19911 (N_19911,N_19505,N_19587);
and U19912 (N_19912,N_19521,N_19560);
xnor U19913 (N_19913,N_19554,N_19584);
and U19914 (N_19914,N_19740,N_19693);
nand U19915 (N_19915,N_19626,N_19741);
xnor U19916 (N_19916,N_19548,N_19602);
xnor U19917 (N_19917,N_19711,N_19637);
or U19918 (N_19918,N_19601,N_19618);
nand U19919 (N_19919,N_19742,N_19735);
and U19920 (N_19920,N_19568,N_19547);
or U19921 (N_19921,N_19660,N_19540);
nor U19922 (N_19922,N_19600,N_19744);
nor U19923 (N_19923,N_19588,N_19600);
nand U19924 (N_19924,N_19657,N_19741);
and U19925 (N_19925,N_19544,N_19668);
or U19926 (N_19926,N_19626,N_19724);
or U19927 (N_19927,N_19623,N_19554);
and U19928 (N_19928,N_19640,N_19558);
and U19929 (N_19929,N_19512,N_19732);
and U19930 (N_19930,N_19610,N_19643);
nor U19931 (N_19931,N_19598,N_19570);
or U19932 (N_19932,N_19664,N_19508);
xor U19933 (N_19933,N_19707,N_19601);
and U19934 (N_19934,N_19591,N_19636);
nor U19935 (N_19935,N_19563,N_19640);
nor U19936 (N_19936,N_19674,N_19663);
and U19937 (N_19937,N_19587,N_19701);
and U19938 (N_19938,N_19555,N_19740);
nand U19939 (N_19939,N_19594,N_19721);
or U19940 (N_19940,N_19530,N_19622);
and U19941 (N_19941,N_19606,N_19625);
or U19942 (N_19942,N_19727,N_19710);
and U19943 (N_19943,N_19520,N_19597);
or U19944 (N_19944,N_19687,N_19650);
nand U19945 (N_19945,N_19680,N_19547);
nor U19946 (N_19946,N_19579,N_19520);
nor U19947 (N_19947,N_19566,N_19730);
and U19948 (N_19948,N_19505,N_19597);
and U19949 (N_19949,N_19623,N_19749);
nor U19950 (N_19950,N_19715,N_19536);
xor U19951 (N_19951,N_19588,N_19702);
and U19952 (N_19952,N_19631,N_19672);
and U19953 (N_19953,N_19570,N_19641);
nand U19954 (N_19954,N_19723,N_19725);
xnor U19955 (N_19955,N_19735,N_19575);
nor U19956 (N_19956,N_19633,N_19634);
nor U19957 (N_19957,N_19697,N_19736);
and U19958 (N_19958,N_19677,N_19546);
and U19959 (N_19959,N_19506,N_19552);
nand U19960 (N_19960,N_19563,N_19730);
and U19961 (N_19961,N_19625,N_19743);
or U19962 (N_19962,N_19515,N_19683);
and U19963 (N_19963,N_19537,N_19659);
nor U19964 (N_19964,N_19516,N_19649);
and U19965 (N_19965,N_19547,N_19732);
nor U19966 (N_19966,N_19619,N_19569);
xor U19967 (N_19967,N_19648,N_19570);
or U19968 (N_19968,N_19515,N_19649);
nand U19969 (N_19969,N_19716,N_19509);
nor U19970 (N_19970,N_19632,N_19657);
nor U19971 (N_19971,N_19631,N_19698);
or U19972 (N_19972,N_19683,N_19647);
nor U19973 (N_19973,N_19648,N_19611);
xnor U19974 (N_19974,N_19713,N_19703);
or U19975 (N_19975,N_19691,N_19638);
or U19976 (N_19976,N_19618,N_19547);
and U19977 (N_19977,N_19620,N_19556);
or U19978 (N_19978,N_19738,N_19666);
and U19979 (N_19979,N_19742,N_19704);
or U19980 (N_19980,N_19540,N_19702);
nand U19981 (N_19981,N_19681,N_19727);
xnor U19982 (N_19982,N_19550,N_19515);
or U19983 (N_19983,N_19723,N_19634);
nand U19984 (N_19984,N_19702,N_19566);
or U19985 (N_19985,N_19629,N_19643);
nand U19986 (N_19986,N_19554,N_19544);
xor U19987 (N_19987,N_19564,N_19668);
or U19988 (N_19988,N_19571,N_19714);
nor U19989 (N_19989,N_19640,N_19588);
nand U19990 (N_19990,N_19582,N_19592);
and U19991 (N_19991,N_19583,N_19643);
xor U19992 (N_19992,N_19555,N_19560);
xor U19993 (N_19993,N_19667,N_19708);
xor U19994 (N_19994,N_19545,N_19582);
nand U19995 (N_19995,N_19673,N_19658);
xor U19996 (N_19996,N_19705,N_19608);
or U19997 (N_19997,N_19730,N_19571);
or U19998 (N_19998,N_19655,N_19588);
nor U19999 (N_19999,N_19574,N_19657);
or U20000 (N_20000,N_19795,N_19968);
nor U20001 (N_20001,N_19991,N_19847);
xor U20002 (N_20002,N_19850,N_19871);
or U20003 (N_20003,N_19934,N_19937);
xor U20004 (N_20004,N_19780,N_19884);
and U20005 (N_20005,N_19929,N_19851);
nand U20006 (N_20006,N_19965,N_19918);
nand U20007 (N_20007,N_19858,N_19814);
nor U20008 (N_20008,N_19774,N_19901);
nand U20009 (N_20009,N_19981,N_19865);
nor U20010 (N_20010,N_19803,N_19950);
and U20011 (N_20011,N_19882,N_19764);
xor U20012 (N_20012,N_19872,N_19878);
nand U20013 (N_20013,N_19952,N_19769);
and U20014 (N_20014,N_19927,N_19943);
nand U20015 (N_20015,N_19870,N_19778);
and U20016 (N_20016,N_19921,N_19958);
and U20017 (N_20017,N_19854,N_19794);
nand U20018 (N_20018,N_19941,N_19869);
and U20019 (N_20019,N_19938,N_19829);
or U20020 (N_20020,N_19860,N_19856);
nor U20021 (N_20021,N_19779,N_19907);
nand U20022 (N_20022,N_19786,N_19959);
nand U20023 (N_20023,N_19857,N_19784);
nor U20024 (N_20024,N_19966,N_19839);
and U20025 (N_20025,N_19842,N_19964);
nand U20026 (N_20026,N_19834,N_19888);
and U20027 (N_20027,N_19848,N_19935);
or U20028 (N_20028,N_19910,N_19924);
nor U20029 (N_20029,N_19824,N_19886);
and U20030 (N_20030,N_19763,N_19751);
xor U20031 (N_20031,N_19999,N_19852);
or U20032 (N_20032,N_19862,N_19951);
xnor U20033 (N_20033,N_19996,N_19953);
or U20034 (N_20034,N_19987,N_19917);
and U20035 (N_20035,N_19796,N_19787);
nand U20036 (N_20036,N_19873,N_19883);
nand U20037 (N_20037,N_19876,N_19930);
nor U20038 (N_20038,N_19802,N_19904);
or U20039 (N_20039,N_19790,N_19838);
nor U20040 (N_20040,N_19864,N_19980);
nand U20041 (N_20041,N_19759,N_19819);
nand U20042 (N_20042,N_19977,N_19785);
and U20043 (N_20043,N_19788,N_19885);
and U20044 (N_20044,N_19755,N_19978);
nand U20045 (N_20045,N_19781,N_19775);
nor U20046 (N_20046,N_19811,N_19773);
xnor U20047 (N_20047,N_19813,N_19815);
xnor U20048 (N_20048,N_19890,N_19900);
or U20049 (N_20049,N_19758,N_19843);
or U20050 (N_20050,N_19822,N_19954);
and U20051 (N_20051,N_19939,N_19949);
nor U20052 (N_20052,N_19932,N_19754);
or U20053 (N_20053,N_19853,N_19906);
nand U20054 (N_20054,N_19891,N_19836);
xnor U20055 (N_20055,N_19875,N_19762);
nor U20056 (N_20056,N_19892,N_19925);
or U20057 (N_20057,N_19989,N_19783);
and U20058 (N_20058,N_19806,N_19776);
nand U20059 (N_20059,N_19970,N_19793);
xnor U20060 (N_20060,N_19902,N_19753);
nand U20061 (N_20061,N_19947,N_19936);
nand U20062 (N_20062,N_19957,N_19805);
nor U20063 (N_20063,N_19913,N_19919);
and U20064 (N_20064,N_19782,N_19797);
xor U20065 (N_20065,N_19899,N_19933);
nor U20066 (N_20066,N_19940,N_19923);
nor U20067 (N_20067,N_19757,N_19993);
or U20068 (N_20068,N_19750,N_19897);
nor U20069 (N_20069,N_19967,N_19920);
xnor U20070 (N_20070,N_19789,N_19816);
nand U20071 (N_20071,N_19976,N_19800);
xor U20072 (N_20072,N_19861,N_19817);
nand U20073 (N_20073,N_19828,N_19889);
xor U20074 (N_20074,N_19955,N_19825);
and U20075 (N_20075,N_19770,N_19974);
and U20076 (N_20076,N_19863,N_19879);
xor U20077 (N_20077,N_19922,N_19804);
nor U20078 (N_20078,N_19792,N_19948);
and U20079 (N_20079,N_19835,N_19926);
or U20080 (N_20080,N_19761,N_19820);
xor U20081 (N_20081,N_19983,N_19812);
or U20082 (N_20082,N_19903,N_19752);
xnor U20083 (N_20083,N_19821,N_19969);
nand U20084 (N_20084,N_19975,N_19931);
nand U20085 (N_20085,N_19830,N_19945);
xor U20086 (N_20086,N_19960,N_19840);
nand U20087 (N_20087,N_19928,N_19859);
nand U20088 (N_20088,N_19961,N_19818);
and U20089 (N_20089,N_19881,N_19801);
nand U20090 (N_20090,N_19971,N_19767);
xnor U20091 (N_20091,N_19867,N_19877);
nand U20092 (N_20092,N_19988,N_19837);
nand U20093 (N_20093,N_19810,N_19849);
nand U20094 (N_20094,N_19893,N_19942);
or U20095 (N_20095,N_19963,N_19998);
and U20096 (N_20096,N_19972,N_19791);
or U20097 (N_20097,N_19798,N_19855);
nor U20098 (N_20098,N_19909,N_19896);
or U20099 (N_20099,N_19777,N_19990);
and U20100 (N_20100,N_19915,N_19911);
and U20101 (N_20101,N_19880,N_19973);
xor U20102 (N_20102,N_19841,N_19823);
and U20103 (N_20103,N_19760,N_19765);
nor U20104 (N_20104,N_19912,N_19831);
nand U20105 (N_20105,N_19808,N_19895);
nand U20106 (N_20106,N_19956,N_19944);
nor U20107 (N_20107,N_19826,N_19799);
and U20108 (N_20108,N_19986,N_19898);
nor U20109 (N_20109,N_19908,N_19833);
nor U20110 (N_20110,N_19756,N_19844);
and U20111 (N_20111,N_19962,N_19868);
and U20112 (N_20112,N_19771,N_19887);
or U20113 (N_20113,N_19866,N_19772);
or U20114 (N_20114,N_19846,N_19916);
and U20115 (N_20115,N_19874,N_19894);
xnor U20116 (N_20116,N_19994,N_19807);
nor U20117 (N_20117,N_19827,N_19905);
or U20118 (N_20118,N_19992,N_19997);
xnor U20119 (N_20119,N_19995,N_19768);
nor U20120 (N_20120,N_19979,N_19809);
xnor U20121 (N_20121,N_19946,N_19914);
or U20122 (N_20122,N_19845,N_19985);
or U20123 (N_20123,N_19984,N_19766);
nor U20124 (N_20124,N_19832,N_19982);
nand U20125 (N_20125,N_19966,N_19908);
nand U20126 (N_20126,N_19824,N_19948);
nor U20127 (N_20127,N_19801,N_19942);
and U20128 (N_20128,N_19956,N_19923);
xnor U20129 (N_20129,N_19754,N_19832);
nand U20130 (N_20130,N_19800,N_19911);
and U20131 (N_20131,N_19843,N_19868);
and U20132 (N_20132,N_19879,N_19982);
or U20133 (N_20133,N_19784,N_19954);
and U20134 (N_20134,N_19765,N_19999);
and U20135 (N_20135,N_19868,N_19856);
or U20136 (N_20136,N_19952,N_19751);
and U20137 (N_20137,N_19852,N_19768);
and U20138 (N_20138,N_19910,N_19900);
nor U20139 (N_20139,N_19773,N_19857);
nor U20140 (N_20140,N_19821,N_19865);
and U20141 (N_20141,N_19898,N_19932);
nor U20142 (N_20142,N_19968,N_19798);
nor U20143 (N_20143,N_19761,N_19856);
nand U20144 (N_20144,N_19752,N_19841);
or U20145 (N_20145,N_19899,N_19859);
or U20146 (N_20146,N_19940,N_19996);
nor U20147 (N_20147,N_19827,N_19891);
xnor U20148 (N_20148,N_19762,N_19974);
and U20149 (N_20149,N_19796,N_19869);
and U20150 (N_20150,N_19990,N_19779);
nand U20151 (N_20151,N_19994,N_19980);
and U20152 (N_20152,N_19878,N_19864);
nor U20153 (N_20153,N_19824,N_19977);
and U20154 (N_20154,N_19785,N_19891);
and U20155 (N_20155,N_19851,N_19762);
nor U20156 (N_20156,N_19949,N_19824);
xor U20157 (N_20157,N_19821,N_19819);
xnor U20158 (N_20158,N_19975,N_19836);
xnor U20159 (N_20159,N_19832,N_19813);
nor U20160 (N_20160,N_19846,N_19771);
nor U20161 (N_20161,N_19880,N_19791);
nor U20162 (N_20162,N_19789,N_19987);
nor U20163 (N_20163,N_19891,N_19954);
or U20164 (N_20164,N_19860,N_19779);
nand U20165 (N_20165,N_19950,N_19913);
and U20166 (N_20166,N_19811,N_19790);
and U20167 (N_20167,N_19882,N_19817);
nor U20168 (N_20168,N_19961,N_19779);
and U20169 (N_20169,N_19970,N_19760);
xor U20170 (N_20170,N_19866,N_19824);
xnor U20171 (N_20171,N_19894,N_19770);
nor U20172 (N_20172,N_19810,N_19951);
and U20173 (N_20173,N_19809,N_19780);
or U20174 (N_20174,N_19774,N_19991);
and U20175 (N_20175,N_19809,N_19835);
nand U20176 (N_20176,N_19837,N_19917);
xnor U20177 (N_20177,N_19978,N_19885);
and U20178 (N_20178,N_19774,N_19982);
or U20179 (N_20179,N_19931,N_19819);
nor U20180 (N_20180,N_19926,N_19965);
xor U20181 (N_20181,N_19776,N_19787);
nand U20182 (N_20182,N_19947,N_19945);
nand U20183 (N_20183,N_19834,N_19906);
nand U20184 (N_20184,N_19920,N_19936);
xnor U20185 (N_20185,N_19894,N_19814);
nor U20186 (N_20186,N_19980,N_19937);
or U20187 (N_20187,N_19854,N_19819);
nor U20188 (N_20188,N_19979,N_19753);
and U20189 (N_20189,N_19754,N_19864);
nor U20190 (N_20190,N_19886,N_19941);
nand U20191 (N_20191,N_19844,N_19853);
nor U20192 (N_20192,N_19757,N_19955);
xnor U20193 (N_20193,N_19930,N_19775);
or U20194 (N_20194,N_19937,N_19933);
xor U20195 (N_20195,N_19928,N_19923);
nor U20196 (N_20196,N_19883,N_19886);
or U20197 (N_20197,N_19858,N_19767);
xnor U20198 (N_20198,N_19882,N_19916);
or U20199 (N_20199,N_19930,N_19767);
xor U20200 (N_20200,N_19983,N_19897);
and U20201 (N_20201,N_19781,N_19907);
and U20202 (N_20202,N_19869,N_19750);
nand U20203 (N_20203,N_19905,N_19863);
nor U20204 (N_20204,N_19830,N_19958);
or U20205 (N_20205,N_19905,N_19853);
and U20206 (N_20206,N_19922,N_19963);
nor U20207 (N_20207,N_19813,N_19760);
and U20208 (N_20208,N_19863,N_19797);
xnor U20209 (N_20209,N_19750,N_19999);
and U20210 (N_20210,N_19936,N_19768);
nand U20211 (N_20211,N_19772,N_19913);
xor U20212 (N_20212,N_19799,N_19805);
nor U20213 (N_20213,N_19767,N_19875);
and U20214 (N_20214,N_19980,N_19779);
nor U20215 (N_20215,N_19925,N_19966);
and U20216 (N_20216,N_19814,N_19972);
nand U20217 (N_20217,N_19980,N_19925);
nor U20218 (N_20218,N_19871,N_19848);
and U20219 (N_20219,N_19986,N_19951);
xor U20220 (N_20220,N_19982,N_19964);
or U20221 (N_20221,N_19857,N_19974);
and U20222 (N_20222,N_19894,N_19841);
nor U20223 (N_20223,N_19994,N_19785);
or U20224 (N_20224,N_19900,N_19985);
nor U20225 (N_20225,N_19752,N_19892);
nor U20226 (N_20226,N_19994,N_19938);
nand U20227 (N_20227,N_19760,N_19855);
or U20228 (N_20228,N_19847,N_19976);
nand U20229 (N_20229,N_19919,N_19812);
and U20230 (N_20230,N_19979,N_19915);
nor U20231 (N_20231,N_19835,N_19909);
and U20232 (N_20232,N_19981,N_19817);
and U20233 (N_20233,N_19958,N_19882);
and U20234 (N_20234,N_19879,N_19953);
xnor U20235 (N_20235,N_19778,N_19946);
xor U20236 (N_20236,N_19778,N_19918);
and U20237 (N_20237,N_19979,N_19910);
nand U20238 (N_20238,N_19906,N_19941);
or U20239 (N_20239,N_19773,N_19756);
nor U20240 (N_20240,N_19867,N_19889);
xnor U20241 (N_20241,N_19912,N_19780);
and U20242 (N_20242,N_19771,N_19948);
nand U20243 (N_20243,N_19874,N_19953);
nor U20244 (N_20244,N_19846,N_19987);
xnor U20245 (N_20245,N_19969,N_19893);
nand U20246 (N_20246,N_19853,N_19967);
xor U20247 (N_20247,N_19816,N_19828);
nand U20248 (N_20248,N_19791,N_19902);
nand U20249 (N_20249,N_19863,N_19942);
and U20250 (N_20250,N_20127,N_20165);
nor U20251 (N_20251,N_20122,N_20123);
nor U20252 (N_20252,N_20095,N_20135);
nand U20253 (N_20253,N_20089,N_20164);
nand U20254 (N_20254,N_20137,N_20209);
nor U20255 (N_20255,N_20020,N_20147);
or U20256 (N_20256,N_20110,N_20138);
and U20257 (N_20257,N_20094,N_20004);
or U20258 (N_20258,N_20150,N_20016);
nand U20259 (N_20259,N_20036,N_20051);
nor U20260 (N_20260,N_20074,N_20023);
xnor U20261 (N_20261,N_20242,N_20172);
and U20262 (N_20262,N_20182,N_20133);
nor U20263 (N_20263,N_20039,N_20047);
and U20264 (N_20264,N_20218,N_20140);
nand U20265 (N_20265,N_20007,N_20021);
nand U20266 (N_20266,N_20104,N_20158);
or U20267 (N_20267,N_20118,N_20102);
and U20268 (N_20268,N_20083,N_20119);
and U20269 (N_20269,N_20238,N_20049);
or U20270 (N_20270,N_20205,N_20189);
xor U20271 (N_20271,N_20130,N_20243);
nor U20272 (N_20272,N_20009,N_20213);
or U20273 (N_20273,N_20234,N_20220);
nand U20274 (N_20274,N_20066,N_20202);
and U20275 (N_20275,N_20204,N_20241);
nor U20276 (N_20276,N_20156,N_20141);
nand U20277 (N_20277,N_20224,N_20173);
or U20278 (N_20278,N_20225,N_20237);
or U20279 (N_20279,N_20113,N_20120);
or U20280 (N_20280,N_20149,N_20197);
nor U20281 (N_20281,N_20201,N_20244);
xor U20282 (N_20282,N_20131,N_20179);
or U20283 (N_20283,N_20005,N_20162);
xnor U20284 (N_20284,N_20246,N_20111);
xnor U20285 (N_20285,N_20192,N_20067);
nor U20286 (N_20286,N_20105,N_20228);
nor U20287 (N_20287,N_20041,N_20203);
xnor U20288 (N_20288,N_20035,N_20029);
nand U20289 (N_20289,N_20177,N_20084);
nand U20290 (N_20290,N_20198,N_20152);
nand U20291 (N_20291,N_20062,N_20043);
and U20292 (N_20292,N_20145,N_20044);
nor U20293 (N_20293,N_20154,N_20157);
and U20294 (N_20294,N_20163,N_20134);
nand U20295 (N_20295,N_20030,N_20055);
or U20296 (N_20296,N_20183,N_20239);
nand U20297 (N_20297,N_20178,N_20229);
nor U20298 (N_20298,N_20143,N_20139);
xor U20299 (N_20299,N_20175,N_20245);
and U20300 (N_20300,N_20000,N_20033);
nand U20301 (N_20301,N_20099,N_20249);
and U20302 (N_20302,N_20223,N_20012);
or U20303 (N_20303,N_20187,N_20010);
nor U20304 (N_20304,N_20231,N_20057);
nand U20305 (N_20305,N_20210,N_20003);
and U20306 (N_20306,N_20235,N_20046);
nor U20307 (N_20307,N_20216,N_20226);
nor U20308 (N_20308,N_20195,N_20121);
and U20309 (N_20309,N_20194,N_20028);
nor U20310 (N_20310,N_20093,N_20193);
and U20311 (N_20311,N_20077,N_20159);
nor U20312 (N_20312,N_20236,N_20085);
and U20313 (N_20313,N_20176,N_20115);
xor U20314 (N_20314,N_20160,N_20103);
nor U20315 (N_20315,N_20180,N_20106);
or U20316 (N_20316,N_20082,N_20060);
or U20317 (N_20317,N_20166,N_20206);
nor U20318 (N_20318,N_20017,N_20240);
nand U20319 (N_20319,N_20171,N_20070);
nor U20320 (N_20320,N_20190,N_20098);
nand U20321 (N_20321,N_20058,N_20230);
and U20322 (N_20322,N_20136,N_20001);
and U20323 (N_20323,N_20169,N_20031);
and U20324 (N_20324,N_20091,N_20038);
nand U20325 (N_20325,N_20073,N_20013);
xnor U20326 (N_20326,N_20097,N_20087);
and U20327 (N_20327,N_20219,N_20072);
nand U20328 (N_20328,N_20018,N_20132);
or U20329 (N_20329,N_20185,N_20126);
or U20330 (N_20330,N_20034,N_20068);
nand U20331 (N_20331,N_20222,N_20037);
nor U20332 (N_20332,N_20191,N_20148);
nor U20333 (N_20333,N_20188,N_20100);
nand U20334 (N_20334,N_20088,N_20170);
xnor U20335 (N_20335,N_20011,N_20196);
or U20336 (N_20336,N_20101,N_20125);
or U20337 (N_20337,N_20096,N_20221);
or U20338 (N_20338,N_20151,N_20080);
or U20339 (N_20339,N_20129,N_20076);
and U20340 (N_20340,N_20014,N_20040);
nor U20341 (N_20341,N_20059,N_20167);
nand U20342 (N_20342,N_20006,N_20247);
nor U20343 (N_20343,N_20065,N_20075);
or U20344 (N_20344,N_20215,N_20050);
xor U20345 (N_20345,N_20045,N_20061);
nor U20346 (N_20346,N_20153,N_20109);
and U20347 (N_20347,N_20002,N_20124);
nor U20348 (N_20348,N_20181,N_20108);
and U20349 (N_20349,N_20056,N_20008);
nand U20350 (N_20350,N_20015,N_20026);
nand U20351 (N_20351,N_20032,N_20211);
or U20352 (N_20352,N_20248,N_20144);
xnor U20353 (N_20353,N_20117,N_20107);
nor U20354 (N_20354,N_20042,N_20071);
and U20355 (N_20355,N_20214,N_20022);
and U20356 (N_20356,N_20128,N_20079);
nand U20357 (N_20357,N_20161,N_20052);
nor U20358 (N_20358,N_20233,N_20217);
nand U20359 (N_20359,N_20232,N_20208);
or U20360 (N_20360,N_20048,N_20025);
nor U20361 (N_20361,N_20212,N_20054);
or U20362 (N_20362,N_20200,N_20227);
or U20363 (N_20363,N_20146,N_20168);
xnor U20364 (N_20364,N_20199,N_20090);
nor U20365 (N_20365,N_20027,N_20092);
nor U20366 (N_20366,N_20207,N_20069);
nor U20367 (N_20367,N_20114,N_20186);
xnor U20368 (N_20368,N_20053,N_20155);
xor U20369 (N_20369,N_20174,N_20064);
and U20370 (N_20370,N_20112,N_20086);
nand U20371 (N_20371,N_20024,N_20116);
nor U20372 (N_20372,N_20081,N_20019);
nor U20373 (N_20373,N_20063,N_20142);
nor U20374 (N_20374,N_20184,N_20078);
nor U20375 (N_20375,N_20031,N_20177);
and U20376 (N_20376,N_20191,N_20233);
nand U20377 (N_20377,N_20000,N_20248);
nor U20378 (N_20378,N_20148,N_20156);
or U20379 (N_20379,N_20206,N_20248);
or U20380 (N_20380,N_20096,N_20007);
and U20381 (N_20381,N_20014,N_20179);
and U20382 (N_20382,N_20053,N_20022);
nand U20383 (N_20383,N_20014,N_20005);
and U20384 (N_20384,N_20077,N_20080);
and U20385 (N_20385,N_20036,N_20076);
and U20386 (N_20386,N_20197,N_20024);
and U20387 (N_20387,N_20060,N_20162);
or U20388 (N_20388,N_20061,N_20101);
or U20389 (N_20389,N_20085,N_20098);
nor U20390 (N_20390,N_20032,N_20087);
or U20391 (N_20391,N_20037,N_20210);
and U20392 (N_20392,N_20127,N_20052);
and U20393 (N_20393,N_20211,N_20125);
nand U20394 (N_20394,N_20115,N_20242);
and U20395 (N_20395,N_20096,N_20158);
nand U20396 (N_20396,N_20218,N_20225);
nor U20397 (N_20397,N_20150,N_20069);
xnor U20398 (N_20398,N_20094,N_20228);
or U20399 (N_20399,N_20190,N_20093);
nand U20400 (N_20400,N_20131,N_20142);
or U20401 (N_20401,N_20163,N_20001);
or U20402 (N_20402,N_20126,N_20094);
nor U20403 (N_20403,N_20007,N_20138);
xnor U20404 (N_20404,N_20002,N_20228);
or U20405 (N_20405,N_20032,N_20097);
nand U20406 (N_20406,N_20049,N_20118);
or U20407 (N_20407,N_20067,N_20003);
and U20408 (N_20408,N_20015,N_20127);
nor U20409 (N_20409,N_20144,N_20011);
or U20410 (N_20410,N_20222,N_20041);
and U20411 (N_20411,N_20190,N_20007);
nor U20412 (N_20412,N_20243,N_20027);
nand U20413 (N_20413,N_20047,N_20202);
xnor U20414 (N_20414,N_20019,N_20104);
or U20415 (N_20415,N_20249,N_20183);
or U20416 (N_20416,N_20011,N_20185);
and U20417 (N_20417,N_20091,N_20243);
nand U20418 (N_20418,N_20025,N_20205);
or U20419 (N_20419,N_20091,N_20151);
and U20420 (N_20420,N_20198,N_20051);
or U20421 (N_20421,N_20058,N_20241);
nand U20422 (N_20422,N_20059,N_20156);
nor U20423 (N_20423,N_20079,N_20049);
or U20424 (N_20424,N_20146,N_20121);
and U20425 (N_20425,N_20053,N_20198);
nand U20426 (N_20426,N_20108,N_20223);
xor U20427 (N_20427,N_20052,N_20185);
and U20428 (N_20428,N_20186,N_20054);
or U20429 (N_20429,N_20120,N_20171);
and U20430 (N_20430,N_20120,N_20130);
xnor U20431 (N_20431,N_20147,N_20177);
and U20432 (N_20432,N_20249,N_20234);
xor U20433 (N_20433,N_20025,N_20120);
and U20434 (N_20434,N_20186,N_20217);
and U20435 (N_20435,N_20093,N_20050);
nor U20436 (N_20436,N_20134,N_20084);
or U20437 (N_20437,N_20062,N_20077);
nand U20438 (N_20438,N_20191,N_20171);
xnor U20439 (N_20439,N_20131,N_20046);
nor U20440 (N_20440,N_20065,N_20217);
or U20441 (N_20441,N_20128,N_20077);
nand U20442 (N_20442,N_20158,N_20134);
xor U20443 (N_20443,N_20178,N_20099);
or U20444 (N_20444,N_20184,N_20072);
nor U20445 (N_20445,N_20071,N_20058);
or U20446 (N_20446,N_20029,N_20026);
and U20447 (N_20447,N_20015,N_20164);
and U20448 (N_20448,N_20013,N_20048);
nor U20449 (N_20449,N_20132,N_20104);
nor U20450 (N_20450,N_20239,N_20090);
or U20451 (N_20451,N_20216,N_20224);
and U20452 (N_20452,N_20143,N_20171);
or U20453 (N_20453,N_20248,N_20109);
nor U20454 (N_20454,N_20194,N_20071);
nor U20455 (N_20455,N_20241,N_20111);
nor U20456 (N_20456,N_20182,N_20107);
nand U20457 (N_20457,N_20147,N_20189);
nand U20458 (N_20458,N_20204,N_20023);
nor U20459 (N_20459,N_20124,N_20134);
nand U20460 (N_20460,N_20076,N_20064);
and U20461 (N_20461,N_20078,N_20197);
nor U20462 (N_20462,N_20167,N_20029);
nand U20463 (N_20463,N_20240,N_20237);
nand U20464 (N_20464,N_20017,N_20230);
nor U20465 (N_20465,N_20138,N_20071);
or U20466 (N_20466,N_20148,N_20237);
or U20467 (N_20467,N_20018,N_20078);
and U20468 (N_20468,N_20099,N_20198);
nor U20469 (N_20469,N_20150,N_20127);
and U20470 (N_20470,N_20248,N_20183);
xor U20471 (N_20471,N_20108,N_20073);
and U20472 (N_20472,N_20049,N_20235);
and U20473 (N_20473,N_20006,N_20045);
and U20474 (N_20474,N_20016,N_20053);
or U20475 (N_20475,N_20100,N_20189);
and U20476 (N_20476,N_20045,N_20170);
and U20477 (N_20477,N_20247,N_20091);
xnor U20478 (N_20478,N_20122,N_20070);
and U20479 (N_20479,N_20249,N_20150);
or U20480 (N_20480,N_20122,N_20017);
or U20481 (N_20481,N_20223,N_20126);
nand U20482 (N_20482,N_20129,N_20060);
or U20483 (N_20483,N_20167,N_20181);
or U20484 (N_20484,N_20147,N_20039);
and U20485 (N_20485,N_20047,N_20101);
nor U20486 (N_20486,N_20173,N_20176);
nand U20487 (N_20487,N_20015,N_20194);
xnor U20488 (N_20488,N_20211,N_20006);
or U20489 (N_20489,N_20236,N_20002);
xor U20490 (N_20490,N_20017,N_20004);
or U20491 (N_20491,N_20176,N_20033);
xnor U20492 (N_20492,N_20056,N_20134);
or U20493 (N_20493,N_20043,N_20229);
nor U20494 (N_20494,N_20188,N_20022);
xor U20495 (N_20495,N_20214,N_20164);
xnor U20496 (N_20496,N_20166,N_20094);
or U20497 (N_20497,N_20222,N_20209);
or U20498 (N_20498,N_20140,N_20040);
xor U20499 (N_20499,N_20051,N_20100);
and U20500 (N_20500,N_20414,N_20253);
or U20501 (N_20501,N_20379,N_20297);
nand U20502 (N_20502,N_20452,N_20351);
or U20503 (N_20503,N_20401,N_20305);
nand U20504 (N_20504,N_20399,N_20377);
or U20505 (N_20505,N_20482,N_20266);
or U20506 (N_20506,N_20328,N_20353);
or U20507 (N_20507,N_20393,N_20289);
nand U20508 (N_20508,N_20259,N_20494);
nor U20509 (N_20509,N_20417,N_20485);
and U20510 (N_20510,N_20406,N_20416);
xor U20511 (N_20511,N_20283,N_20250);
and U20512 (N_20512,N_20394,N_20324);
or U20513 (N_20513,N_20313,N_20465);
nand U20514 (N_20514,N_20350,N_20486);
or U20515 (N_20515,N_20273,N_20407);
xnor U20516 (N_20516,N_20489,N_20308);
nor U20517 (N_20517,N_20337,N_20371);
nand U20518 (N_20518,N_20488,N_20293);
nor U20519 (N_20519,N_20443,N_20309);
and U20520 (N_20520,N_20338,N_20478);
or U20521 (N_20521,N_20476,N_20357);
nor U20522 (N_20522,N_20360,N_20453);
nand U20523 (N_20523,N_20397,N_20498);
nor U20524 (N_20524,N_20497,N_20472);
or U20525 (N_20525,N_20369,N_20320);
nand U20526 (N_20526,N_20356,N_20451);
or U20527 (N_20527,N_20358,N_20280);
nor U20528 (N_20528,N_20348,N_20368);
and U20529 (N_20529,N_20372,N_20285);
nor U20530 (N_20530,N_20256,N_20400);
xor U20531 (N_20531,N_20439,N_20435);
nor U20532 (N_20532,N_20267,N_20387);
and U20533 (N_20533,N_20463,N_20466);
or U20534 (N_20534,N_20340,N_20271);
nand U20535 (N_20535,N_20449,N_20262);
or U20536 (N_20536,N_20496,N_20291);
or U20537 (N_20537,N_20345,N_20475);
nor U20538 (N_20538,N_20403,N_20269);
xor U20539 (N_20539,N_20433,N_20464);
nand U20540 (N_20540,N_20410,N_20275);
and U20541 (N_20541,N_20299,N_20479);
nand U20542 (N_20542,N_20391,N_20318);
xnor U20543 (N_20543,N_20359,N_20390);
or U20544 (N_20544,N_20481,N_20252);
nand U20545 (N_20545,N_20336,N_20376);
nand U20546 (N_20546,N_20321,N_20314);
nor U20547 (N_20547,N_20362,N_20278);
or U20548 (N_20548,N_20460,N_20491);
nand U20549 (N_20549,N_20347,N_20396);
nor U20550 (N_20550,N_20366,N_20296);
and U20551 (N_20551,N_20263,N_20438);
or U20552 (N_20552,N_20402,N_20290);
xor U20553 (N_20553,N_20343,N_20431);
xnor U20554 (N_20554,N_20454,N_20427);
nand U20555 (N_20555,N_20447,N_20474);
xnor U20556 (N_20556,N_20361,N_20257);
xor U20557 (N_20557,N_20395,N_20346);
and U20558 (N_20558,N_20493,N_20270);
xnor U20559 (N_20559,N_20388,N_20317);
nand U20560 (N_20560,N_20286,N_20277);
nor U20561 (N_20561,N_20331,N_20327);
nor U20562 (N_20562,N_20419,N_20384);
or U20563 (N_20563,N_20445,N_20484);
and U20564 (N_20564,N_20440,N_20332);
and U20565 (N_20565,N_20492,N_20382);
xor U20566 (N_20566,N_20292,N_20375);
or U20567 (N_20567,N_20272,N_20373);
nand U20568 (N_20568,N_20398,N_20349);
or U20569 (N_20569,N_20300,N_20261);
or U20570 (N_20570,N_20279,N_20436);
and U20571 (N_20571,N_20430,N_20378);
nand U20572 (N_20572,N_20483,N_20381);
and U20573 (N_20573,N_20455,N_20499);
xor U20574 (N_20574,N_20477,N_20469);
nor U20575 (N_20575,N_20344,N_20404);
and U20576 (N_20576,N_20423,N_20330);
and U20577 (N_20577,N_20386,N_20354);
and U20578 (N_20578,N_20473,N_20298);
xor U20579 (N_20579,N_20258,N_20458);
or U20580 (N_20580,N_20255,N_20428);
and U20581 (N_20581,N_20325,N_20312);
or U20582 (N_20582,N_20306,N_20471);
nand U20583 (N_20583,N_20364,N_20322);
or U20584 (N_20584,N_20374,N_20462);
or U20585 (N_20585,N_20304,N_20412);
nand U20586 (N_20586,N_20422,N_20487);
xnor U20587 (N_20587,N_20281,N_20326);
nand U20588 (N_20588,N_20315,N_20495);
xnor U20589 (N_20589,N_20264,N_20444);
or U20590 (N_20590,N_20333,N_20265);
or U20591 (N_20591,N_20480,N_20461);
nand U20592 (N_20592,N_20418,N_20284);
nand U20593 (N_20593,N_20307,N_20339);
nand U20594 (N_20594,N_20335,N_20434);
and U20595 (N_20595,N_20301,N_20303);
or U20596 (N_20596,N_20254,N_20490);
xnor U20597 (N_20597,N_20367,N_20457);
nand U20598 (N_20598,N_20355,N_20385);
and U20599 (N_20599,N_20310,N_20302);
nand U20600 (N_20600,N_20425,N_20442);
xnor U20601 (N_20601,N_20380,N_20329);
and U20602 (N_20602,N_20450,N_20413);
or U20603 (N_20603,N_20365,N_20415);
nor U20604 (N_20604,N_20311,N_20295);
or U20605 (N_20605,N_20342,N_20323);
and U20606 (N_20606,N_20287,N_20459);
and U20607 (N_20607,N_20467,N_20432);
and U20608 (N_20608,N_20352,N_20429);
or U20609 (N_20609,N_20334,N_20319);
xor U20610 (N_20610,N_20421,N_20408);
or U20611 (N_20611,N_20363,N_20260);
nor U20612 (N_20612,N_20316,N_20441);
nand U20613 (N_20613,N_20370,N_20409);
or U20614 (N_20614,N_20437,N_20446);
and U20615 (N_20615,N_20282,N_20389);
or U20616 (N_20616,N_20456,N_20411);
and U20617 (N_20617,N_20274,N_20341);
or U20618 (N_20618,N_20294,N_20420);
xnor U20619 (N_20619,N_20251,N_20468);
or U20620 (N_20620,N_20426,N_20288);
nor U20621 (N_20621,N_20276,N_20268);
and U20622 (N_20622,N_20383,N_20405);
or U20623 (N_20623,N_20424,N_20392);
or U20624 (N_20624,N_20470,N_20448);
and U20625 (N_20625,N_20315,N_20486);
or U20626 (N_20626,N_20314,N_20323);
and U20627 (N_20627,N_20380,N_20424);
xor U20628 (N_20628,N_20358,N_20461);
nor U20629 (N_20629,N_20398,N_20360);
nor U20630 (N_20630,N_20256,N_20432);
and U20631 (N_20631,N_20459,N_20367);
or U20632 (N_20632,N_20424,N_20479);
nand U20633 (N_20633,N_20313,N_20319);
xnor U20634 (N_20634,N_20265,N_20341);
or U20635 (N_20635,N_20276,N_20394);
and U20636 (N_20636,N_20286,N_20389);
nor U20637 (N_20637,N_20493,N_20257);
nor U20638 (N_20638,N_20395,N_20344);
nor U20639 (N_20639,N_20359,N_20271);
xor U20640 (N_20640,N_20429,N_20266);
nor U20641 (N_20641,N_20407,N_20363);
nand U20642 (N_20642,N_20261,N_20349);
xor U20643 (N_20643,N_20354,N_20481);
and U20644 (N_20644,N_20458,N_20469);
nor U20645 (N_20645,N_20250,N_20450);
or U20646 (N_20646,N_20311,N_20413);
nor U20647 (N_20647,N_20478,N_20420);
and U20648 (N_20648,N_20400,N_20322);
and U20649 (N_20649,N_20313,N_20475);
and U20650 (N_20650,N_20301,N_20299);
or U20651 (N_20651,N_20414,N_20484);
nor U20652 (N_20652,N_20348,N_20333);
nor U20653 (N_20653,N_20288,N_20364);
or U20654 (N_20654,N_20482,N_20489);
nor U20655 (N_20655,N_20317,N_20423);
nand U20656 (N_20656,N_20352,N_20329);
and U20657 (N_20657,N_20349,N_20339);
or U20658 (N_20658,N_20264,N_20402);
xnor U20659 (N_20659,N_20410,N_20336);
nand U20660 (N_20660,N_20460,N_20345);
or U20661 (N_20661,N_20280,N_20279);
xnor U20662 (N_20662,N_20367,N_20379);
or U20663 (N_20663,N_20290,N_20498);
and U20664 (N_20664,N_20466,N_20478);
or U20665 (N_20665,N_20445,N_20449);
xor U20666 (N_20666,N_20441,N_20284);
and U20667 (N_20667,N_20457,N_20278);
nand U20668 (N_20668,N_20360,N_20419);
nand U20669 (N_20669,N_20255,N_20426);
or U20670 (N_20670,N_20263,N_20399);
and U20671 (N_20671,N_20323,N_20403);
nand U20672 (N_20672,N_20343,N_20329);
nor U20673 (N_20673,N_20313,N_20328);
nand U20674 (N_20674,N_20379,N_20271);
or U20675 (N_20675,N_20482,N_20488);
nor U20676 (N_20676,N_20283,N_20269);
and U20677 (N_20677,N_20469,N_20472);
nand U20678 (N_20678,N_20417,N_20418);
or U20679 (N_20679,N_20317,N_20471);
nand U20680 (N_20680,N_20341,N_20262);
xnor U20681 (N_20681,N_20435,N_20266);
nand U20682 (N_20682,N_20253,N_20426);
xor U20683 (N_20683,N_20494,N_20321);
xnor U20684 (N_20684,N_20461,N_20366);
and U20685 (N_20685,N_20297,N_20489);
or U20686 (N_20686,N_20351,N_20454);
and U20687 (N_20687,N_20303,N_20269);
nand U20688 (N_20688,N_20366,N_20398);
nor U20689 (N_20689,N_20332,N_20323);
and U20690 (N_20690,N_20347,N_20300);
nand U20691 (N_20691,N_20274,N_20320);
nand U20692 (N_20692,N_20457,N_20482);
and U20693 (N_20693,N_20358,N_20481);
and U20694 (N_20694,N_20274,N_20411);
nor U20695 (N_20695,N_20355,N_20406);
and U20696 (N_20696,N_20418,N_20256);
and U20697 (N_20697,N_20363,N_20298);
or U20698 (N_20698,N_20382,N_20482);
nand U20699 (N_20699,N_20347,N_20271);
xnor U20700 (N_20700,N_20373,N_20470);
nand U20701 (N_20701,N_20364,N_20269);
and U20702 (N_20702,N_20404,N_20476);
nand U20703 (N_20703,N_20389,N_20422);
or U20704 (N_20704,N_20333,N_20328);
or U20705 (N_20705,N_20451,N_20355);
xor U20706 (N_20706,N_20356,N_20384);
or U20707 (N_20707,N_20484,N_20271);
xnor U20708 (N_20708,N_20430,N_20345);
nor U20709 (N_20709,N_20403,N_20418);
xnor U20710 (N_20710,N_20495,N_20310);
xnor U20711 (N_20711,N_20371,N_20342);
and U20712 (N_20712,N_20268,N_20496);
nor U20713 (N_20713,N_20290,N_20284);
nand U20714 (N_20714,N_20470,N_20440);
nand U20715 (N_20715,N_20485,N_20286);
or U20716 (N_20716,N_20258,N_20290);
nand U20717 (N_20717,N_20488,N_20434);
or U20718 (N_20718,N_20346,N_20341);
xor U20719 (N_20719,N_20370,N_20397);
nand U20720 (N_20720,N_20271,N_20324);
or U20721 (N_20721,N_20307,N_20369);
or U20722 (N_20722,N_20431,N_20465);
nand U20723 (N_20723,N_20359,N_20306);
nand U20724 (N_20724,N_20299,N_20358);
nor U20725 (N_20725,N_20361,N_20433);
nor U20726 (N_20726,N_20396,N_20344);
or U20727 (N_20727,N_20263,N_20307);
or U20728 (N_20728,N_20497,N_20386);
nand U20729 (N_20729,N_20396,N_20473);
or U20730 (N_20730,N_20412,N_20465);
nor U20731 (N_20731,N_20447,N_20337);
nand U20732 (N_20732,N_20287,N_20393);
nor U20733 (N_20733,N_20489,N_20370);
or U20734 (N_20734,N_20490,N_20297);
or U20735 (N_20735,N_20336,N_20384);
and U20736 (N_20736,N_20326,N_20440);
xnor U20737 (N_20737,N_20289,N_20383);
nand U20738 (N_20738,N_20422,N_20464);
xnor U20739 (N_20739,N_20454,N_20388);
or U20740 (N_20740,N_20340,N_20345);
or U20741 (N_20741,N_20353,N_20261);
or U20742 (N_20742,N_20328,N_20454);
or U20743 (N_20743,N_20280,N_20415);
and U20744 (N_20744,N_20420,N_20434);
or U20745 (N_20745,N_20450,N_20448);
xnor U20746 (N_20746,N_20384,N_20405);
or U20747 (N_20747,N_20255,N_20252);
xnor U20748 (N_20748,N_20442,N_20303);
or U20749 (N_20749,N_20408,N_20324);
or U20750 (N_20750,N_20729,N_20645);
nand U20751 (N_20751,N_20646,N_20541);
nand U20752 (N_20752,N_20746,N_20523);
nor U20753 (N_20753,N_20555,N_20640);
nand U20754 (N_20754,N_20508,N_20522);
and U20755 (N_20755,N_20588,N_20744);
and U20756 (N_20756,N_20677,N_20520);
and U20757 (N_20757,N_20561,N_20727);
nand U20758 (N_20758,N_20509,N_20650);
xnor U20759 (N_20759,N_20535,N_20660);
or U20760 (N_20760,N_20601,N_20696);
xor U20761 (N_20761,N_20745,N_20639);
or U20762 (N_20762,N_20705,N_20649);
xor U20763 (N_20763,N_20662,N_20558);
or U20764 (N_20764,N_20512,N_20593);
xor U20765 (N_20765,N_20518,N_20557);
nor U20766 (N_20766,N_20681,N_20618);
and U20767 (N_20767,N_20570,N_20576);
xnor U20768 (N_20768,N_20595,N_20679);
and U20769 (N_20769,N_20655,N_20678);
xor U20770 (N_20770,N_20687,N_20702);
or U20771 (N_20771,N_20513,N_20693);
xor U20772 (N_20772,N_20537,N_20721);
nor U20773 (N_20773,N_20565,N_20502);
or U20774 (N_20774,N_20673,N_20562);
nand U20775 (N_20775,N_20553,N_20619);
and U20776 (N_20776,N_20574,N_20590);
nand U20777 (N_20777,N_20586,N_20686);
and U20778 (N_20778,N_20572,N_20566);
nand U20779 (N_20779,N_20547,N_20549);
nand U20780 (N_20780,N_20628,N_20675);
nor U20781 (N_20781,N_20610,N_20609);
nor U20782 (N_20782,N_20706,N_20667);
xor U20783 (N_20783,N_20669,N_20592);
nor U20784 (N_20784,N_20584,N_20680);
or U20785 (N_20785,N_20642,N_20691);
and U20786 (N_20786,N_20538,N_20585);
xnor U20787 (N_20787,N_20536,N_20560);
or U20788 (N_20788,N_20500,N_20615);
nor U20789 (N_20789,N_20632,N_20551);
or U20790 (N_20790,N_20652,N_20703);
or U20791 (N_20791,N_20730,N_20511);
or U20792 (N_20792,N_20713,N_20731);
nand U20793 (N_20793,N_20550,N_20738);
xnor U20794 (N_20794,N_20622,N_20682);
nor U20795 (N_20795,N_20736,N_20666);
nand U20796 (N_20796,N_20689,N_20578);
nor U20797 (N_20797,N_20748,N_20626);
xor U20798 (N_20798,N_20505,N_20657);
nand U20799 (N_20799,N_20659,N_20621);
xor U20800 (N_20800,N_20644,N_20651);
or U20801 (N_20801,N_20563,N_20577);
or U20802 (N_20802,N_20514,N_20737);
and U20803 (N_20803,N_20741,N_20698);
or U20804 (N_20804,N_20725,N_20631);
and U20805 (N_20805,N_20583,N_20743);
nor U20806 (N_20806,N_20569,N_20596);
nand U20807 (N_20807,N_20732,N_20587);
xnor U20808 (N_20808,N_20692,N_20740);
or U20809 (N_20809,N_20603,N_20726);
and U20810 (N_20810,N_20665,N_20571);
or U20811 (N_20811,N_20539,N_20575);
nand U20812 (N_20812,N_20717,N_20684);
nor U20813 (N_20813,N_20529,N_20749);
or U20814 (N_20814,N_20720,N_20735);
nand U20815 (N_20815,N_20739,N_20641);
xor U20816 (N_20816,N_20625,N_20567);
and U20817 (N_20817,N_20733,N_20519);
nand U20818 (N_20818,N_20531,N_20715);
and U20819 (N_20819,N_20580,N_20579);
or U20820 (N_20820,N_20525,N_20707);
nor U20821 (N_20821,N_20616,N_20637);
or U20822 (N_20822,N_20668,N_20724);
xnor U20823 (N_20823,N_20542,N_20709);
xor U20824 (N_20824,N_20672,N_20697);
nor U20825 (N_20825,N_20663,N_20545);
and U20826 (N_20826,N_20544,N_20582);
nor U20827 (N_20827,N_20712,N_20515);
nor U20828 (N_20828,N_20643,N_20552);
xnor U20829 (N_20829,N_20629,N_20636);
or U20830 (N_20830,N_20510,N_20647);
nand U20831 (N_20831,N_20704,N_20676);
xor U20832 (N_20832,N_20611,N_20633);
or U20833 (N_20833,N_20589,N_20613);
nor U20834 (N_20834,N_20530,N_20701);
nand U20835 (N_20835,N_20614,N_20653);
nor U20836 (N_20836,N_20671,N_20699);
xnor U20837 (N_20837,N_20658,N_20564);
nor U20838 (N_20838,N_20714,N_20620);
nor U20839 (N_20839,N_20548,N_20591);
xor U20840 (N_20840,N_20528,N_20521);
and U20841 (N_20841,N_20627,N_20608);
xnor U20842 (N_20842,N_20599,N_20594);
nor U20843 (N_20843,N_20656,N_20661);
and U20844 (N_20844,N_20638,N_20607);
nand U20845 (N_20845,N_20598,N_20718);
xor U20846 (N_20846,N_20606,N_20524);
or U20847 (N_20847,N_20554,N_20747);
nor U20848 (N_20848,N_20602,N_20600);
nand U20849 (N_20849,N_20734,N_20534);
nor U20850 (N_20850,N_20501,N_20504);
and U20851 (N_20851,N_20722,N_20617);
and U20852 (N_20852,N_20664,N_20742);
xor U20853 (N_20853,N_20695,N_20581);
nor U20854 (N_20854,N_20708,N_20543);
nand U20855 (N_20855,N_20605,N_20711);
or U20856 (N_20856,N_20694,N_20573);
and U20857 (N_20857,N_20700,N_20532);
nor U20858 (N_20858,N_20630,N_20604);
nand U20859 (N_20859,N_20503,N_20623);
nor U20860 (N_20860,N_20688,N_20728);
and U20861 (N_20861,N_20710,N_20506);
xnor U20862 (N_20862,N_20533,N_20719);
or U20863 (N_20863,N_20723,N_20674);
xor U20864 (N_20864,N_20683,N_20527);
nand U20865 (N_20865,N_20635,N_20516);
nand U20866 (N_20866,N_20654,N_20540);
or U20867 (N_20867,N_20670,N_20526);
and U20868 (N_20868,N_20634,N_20507);
nand U20869 (N_20869,N_20690,N_20559);
xor U20870 (N_20870,N_20546,N_20568);
nand U20871 (N_20871,N_20685,N_20517);
or U20872 (N_20872,N_20716,N_20624);
nand U20873 (N_20873,N_20648,N_20612);
xnor U20874 (N_20874,N_20597,N_20556);
nor U20875 (N_20875,N_20577,N_20682);
or U20876 (N_20876,N_20533,N_20606);
and U20877 (N_20877,N_20692,N_20643);
or U20878 (N_20878,N_20729,N_20716);
or U20879 (N_20879,N_20571,N_20663);
or U20880 (N_20880,N_20627,N_20702);
xor U20881 (N_20881,N_20719,N_20740);
xor U20882 (N_20882,N_20550,N_20669);
xor U20883 (N_20883,N_20584,N_20736);
xnor U20884 (N_20884,N_20712,N_20723);
xnor U20885 (N_20885,N_20565,N_20677);
nor U20886 (N_20886,N_20671,N_20577);
nor U20887 (N_20887,N_20561,N_20547);
nand U20888 (N_20888,N_20635,N_20747);
xor U20889 (N_20889,N_20540,N_20690);
xor U20890 (N_20890,N_20650,N_20597);
nand U20891 (N_20891,N_20647,N_20748);
nand U20892 (N_20892,N_20747,N_20719);
xor U20893 (N_20893,N_20527,N_20641);
nand U20894 (N_20894,N_20506,N_20657);
and U20895 (N_20895,N_20527,N_20535);
nor U20896 (N_20896,N_20507,N_20671);
and U20897 (N_20897,N_20655,N_20642);
nor U20898 (N_20898,N_20511,N_20552);
or U20899 (N_20899,N_20658,N_20705);
nand U20900 (N_20900,N_20503,N_20704);
xor U20901 (N_20901,N_20526,N_20549);
nor U20902 (N_20902,N_20660,N_20586);
xor U20903 (N_20903,N_20520,N_20624);
or U20904 (N_20904,N_20526,N_20619);
and U20905 (N_20905,N_20539,N_20596);
or U20906 (N_20906,N_20728,N_20523);
xor U20907 (N_20907,N_20645,N_20650);
nor U20908 (N_20908,N_20724,N_20636);
or U20909 (N_20909,N_20673,N_20502);
or U20910 (N_20910,N_20635,N_20697);
and U20911 (N_20911,N_20642,N_20606);
or U20912 (N_20912,N_20539,N_20549);
nand U20913 (N_20913,N_20652,N_20551);
and U20914 (N_20914,N_20663,N_20568);
xnor U20915 (N_20915,N_20708,N_20715);
and U20916 (N_20916,N_20684,N_20723);
and U20917 (N_20917,N_20536,N_20605);
or U20918 (N_20918,N_20738,N_20602);
nand U20919 (N_20919,N_20617,N_20630);
nor U20920 (N_20920,N_20611,N_20681);
nand U20921 (N_20921,N_20731,N_20639);
nor U20922 (N_20922,N_20677,N_20735);
nor U20923 (N_20923,N_20581,N_20729);
nor U20924 (N_20924,N_20678,N_20689);
xor U20925 (N_20925,N_20696,N_20525);
nor U20926 (N_20926,N_20628,N_20701);
nor U20927 (N_20927,N_20617,N_20700);
nand U20928 (N_20928,N_20699,N_20643);
or U20929 (N_20929,N_20633,N_20741);
or U20930 (N_20930,N_20569,N_20544);
and U20931 (N_20931,N_20699,N_20573);
or U20932 (N_20932,N_20569,N_20532);
and U20933 (N_20933,N_20697,N_20575);
nand U20934 (N_20934,N_20602,N_20638);
or U20935 (N_20935,N_20539,N_20668);
and U20936 (N_20936,N_20562,N_20532);
nor U20937 (N_20937,N_20608,N_20711);
xor U20938 (N_20938,N_20638,N_20576);
and U20939 (N_20939,N_20545,N_20681);
or U20940 (N_20940,N_20678,N_20545);
and U20941 (N_20941,N_20652,N_20576);
xor U20942 (N_20942,N_20706,N_20669);
xor U20943 (N_20943,N_20522,N_20666);
nor U20944 (N_20944,N_20556,N_20702);
or U20945 (N_20945,N_20527,N_20558);
nand U20946 (N_20946,N_20514,N_20532);
and U20947 (N_20947,N_20546,N_20673);
or U20948 (N_20948,N_20634,N_20601);
nor U20949 (N_20949,N_20572,N_20654);
xor U20950 (N_20950,N_20575,N_20739);
nand U20951 (N_20951,N_20530,N_20629);
and U20952 (N_20952,N_20650,N_20665);
nor U20953 (N_20953,N_20739,N_20632);
nand U20954 (N_20954,N_20558,N_20724);
or U20955 (N_20955,N_20504,N_20682);
or U20956 (N_20956,N_20609,N_20680);
or U20957 (N_20957,N_20569,N_20604);
xor U20958 (N_20958,N_20644,N_20706);
or U20959 (N_20959,N_20686,N_20631);
nand U20960 (N_20960,N_20522,N_20518);
or U20961 (N_20961,N_20590,N_20569);
nand U20962 (N_20962,N_20504,N_20647);
and U20963 (N_20963,N_20747,N_20609);
nand U20964 (N_20964,N_20502,N_20642);
nor U20965 (N_20965,N_20718,N_20624);
or U20966 (N_20966,N_20556,N_20731);
nor U20967 (N_20967,N_20681,N_20540);
nor U20968 (N_20968,N_20601,N_20683);
xnor U20969 (N_20969,N_20532,N_20537);
or U20970 (N_20970,N_20677,N_20607);
and U20971 (N_20971,N_20658,N_20604);
nand U20972 (N_20972,N_20552,N_20693);
nand U20973 (N_20973,N_20569,N_20572);
and U20974 (N_20974,N_20735,N_20732);
nand U20975 (N_20975,N_20737,N_20599);
nand U20976 (N_20976,N_20634,N_20715);
or U20977 (N_20977,N_20549,N_20583);
or U20978 (N_20978,N_20574,N_20643);
nand U20979 (N_20979,N_20672,N_20572);
nand U20980 (N_20980,N_20639,N_20718);
nor U20981 (N_20981,N_20722,N_20534);
or U20982 (N_20982,N_20664,N_20637);
and U20983 (N_20983,N_20660,N_20635);
nor U20984 (N_20984,N_20531,N_20690);
nand U20985 (N_20985,N_20611,N_20695);
or U20986 (N_20986,N_20580,N_20677);
and U20987 (N_20987,N_20649,N_20719);
or U20988 (N_20988,N_20584,N_20586);
xnor U20989 (N_20989,N_20574,N_20637);
xnor U20990 (N_20990,N_20736,N_20631);
xnor U20991 (N_20991,N_20547,N_20564);
and U20992 (N_20992,N_20598,N_20530);
or U20993 (N_20993,N_20622,N_20608);
and U20994 (N_20994,N_20672,N_20557);
or U20995 (N_20995,N_20674,N_20598);
nand U20996 (N_20996,N_20632,N_20741);
nand U20997 (N_20997,N_20667,N_20555);
xnor U20998 (N_20998,N_20680,N_20704);
xor U20999 (N_20999,N_20631,N_20622);
xor U21000 (N_21000,N_20844,N_20871);
or U21001 (N_21001,N_20779,N_20921);
nand U21002 (N_21002,N_20822,N_20919);
nand U21003 (N_21003,N_20854,N_20966);
and U21004 (N_21004,N_20958,N_20814);
nand U21005 (N_21005,N_20894,N_20913);
xor U21006 (N_21006,N_20990,N_20988);
nor U21007 (N_21007,N_20781,N_20905);
nor U21008 (N_21008,N_20794,N_20908);
nand U21009 (N_21009,N_20791,N_20785);
xnor U21010 (N_21010,N_20956,N_20878);
or U21011 (N_21011,N_20750,N_20889);
nor U21012 (N_21012,N_20825,N_20768);
or U21013 (N_21013,N_20997,N_20827);
nor U21014 (N_21014,N_20954,N_20796);
xnor U21015 (N_21015,N_20893,N_20992);
nand U21016 (N_21016,N_20898,N_20982);
nor U21017 (N_21017,N_20974,N_20979);
nand U21018 (N_21018,N_20873,N_20863);
and U21019 (N_21019,N_20955,N_20776);
nor U21020 (N_21020,N_20927,N_20883);
or U21021 (N_21021,N_20876,N_20900);
nor U21022 (N_21022,N_20906,N_20769);
xor U21023 (N_21023,N_20763,N_20853);
nor U21024 (N_21024,N_20952,N_20849);
nand U21025 (N_21025,N_20887,N_20820);
nand U21026 (N_21026,N_20939,N_20999);
and U21027 (N_21027,N_20882,N_20777);
and U21028 (N_21028,N_20759,N_20874);
nor U21029 (N_21029,N_20751,N_20856);
nand U21030 (N_21030,N_20766,N_20957);
nor U21031 (N_21031,N_20783,N_20864);
or U21032 (N_21032,N_20753,N_20931);
or U21033 (N_21033,N_20869,N_20852);
nor U21034 (N_21034,N_20802,N_20773);
xor U21035 (N_21035,N_20870,N_20860);
or U21036 (N_21036,N_20929,N_20885);
nor U21037 (N_21037,N_20760,N_20810);
nand U21038 (N_21038,N_20943,N_20805);
and U21039 (N_21039,N_20800,N_20808);
nand U21040 (N_21040,N_20786,N_20924);
nor U21041 (N_21041,N_20841,N_20976);
or U21042 (N_21042,N_20964,N_20946);
and U21043 (N_21043,N_20961,N_20950);
nand U21044 (N_21044,N_20821,N_20945);
nor U21045 (N_21045,N_20948,N_20770);
xor U21046 (N_21046,N_20847,N_20754);
nor U21047 (N_21047,N_20914,N_20771);
nand U21048 (N_21048,N_20923,N_20891);
or U21049 (N_21049,N_20840,N_20940);
or U21050 (N_21050,N_20843,N_20888);
nand U21051 (N_21051,N_20793,N_20767);
and U21052 (N_21052,N_20823,N_20970);
xor U21053 (N_21053,N_20787,N_20971);
nand U21054 (N_21054,N_20816,N_20835);
xor U21055 (N_21055,N_20792,N_20831);
or U21056 (N_21056,N_20764,N_20757);
and U21057 (N_21057,N_20934,N_20829);
or U21058 (N_21058,N_20755,N_20765);
nand U21059 (N_21059,N_20915,N_20903);
xnor U21060 (N_21060,N_20809,N_20951);
xnor U21061 (N_21061,N_20758,N_20987);
nor U21062 (N_21062,N_20911,N_20818);
nor U21063 (N_21063,N_20833,N_20995);
nand U21064 (N_21064,N_20965,N_20817);
nor U21065 (N_21065,N_20895,N_20813);
and U21066 (N_21066,N_20925,N_20868);
nor U21067 (N_21067,N_20930,N_20944);
nand U21068 (N_21068,N_20967,N_20941);
nand U21069 (N_21069,N_20973,N_20837);
nand U21070 (N_21070,N_20932,N_20910);
and U21071 (N_21071,N_20865,N_20761);
xor U21072 (N_21072,N_20993,N_20811);
nand U21073 (N_21073,N_20782,N_20828);
nand U21074 (N_21074,N_20928,N_20953);
nor U21075 (N_21075,N_20806,N_20866);
or U21076 (N_21076,N_20949,N_20846);
xor U21077 (N_21077,N_20807,N_20851);
xnor U21078 (N_21078,N_20922,N_20935);
nand U21079 (N_21079,N_20875,N_20798);
or U21080 (N_21080,N_20980,N_20937);
or U21081 (N_21081,N_20855,N_20861);
nor U21082 (N_21082,N_20969,N_20886);
nand U21083 (N_21083,N_20872,N_20819);
nand U21084 (N_21084,N_20983,N_20963);
nor U21085 (N_21085,N_20890,N_20830);
nor U21086 (N_21086,N_20978,N_20884);
and U21087 (N_21087,N_20904,N_20772);
or U21088 (N_21088,N_20892,N_20838);
xnor U21089 (N_21089,N_20877,N_20784);
or U21090 (N_21090,N_20762,N_20752);
nor U21091 (N_21091,N_20909,N_20857);
nand U21092 (N_21092,N_20879,N_20901);
or U21093 (N_21093,N_20858,N_20880);
nand U21094 (N_21094,N_20826,N_20920);
nor U21095 (N_21095,N_20832,N_20850);
nand U21096 (N_21096,N_20795,N_20789);
and U21097 (N_21097,N_20801,N_20859);
or U21098 (N_21098,N_20975,N_20839);
nand U21099 (N_21099,N_20862,N_20899);
nor U21100 (N_21100,N_20836,N_20998);
nor U21101 (N_21101,N_20962,N_20834);
or U21102 (N_21102,N_20881,N_20942);
nor U21103 (N_21103,N_20989,N_20756);
and U21104 (N_21104,N_20824,N_20918);
or U21105 (N_21105,N_20947,N_20896);
or U21106 (N_21106,N_20959,N_20994);
nor U21107 (N_21107,N_20778,N_20972);
nand U21108 (N_21108,N_20985,N_20788);
and U21109 (N_21109,N_20775,N_20799);
xor U21110 (N_21110,N_20803,N_20977);
xnor U21111 (N_21111,N_20842,N_20933);
nand U21112 (N_21112,N_20902,N_20968);
xor U21113 (N_21113,N_20960,N_20867);
xor U21114 (N_21114,N_20938,N_20981);
nor U21115 (N_21115,N_20774,N_20815);
xnor U21116 (N_21116,N_20926,N_20986);
or U21117 (N_21117,N_20790,N_20804);
nand U21118 (N_21118,N_20780,N_20897);
or U21119 (N_21119,N_20916,N_20912);
or U21120 (N_21120,N_20996,N_20845);
or U21121 (N_21121,N_20907,N_20797);
or U21122 (N_21122,N_20991,N_20917);
xnor U21123 (N_21123,N_20936,N_20812);
nor U21124 (N_21124,N_20848,N_20984);
xnor U21125 (N_21125,N_20880,N_20925);
or U21126 (N_21126,N_20833,N_20940);
nor U21127 (N_21127,N_20895,N_20830);
nand U21128 (N_21128,N_20850,N_20871);
or U21129 (N_21129,N_20837,N_20986);
xor U21130 (N_21130,N_20785,N_20835);
nor U21131 (N_21131,N_20981,N_20958);
nand U21132 (N_21132,N_20885,N_20994);
xnor U21133 (N_21133,N_20755,N_20868);
nor U21134 (N_21134,N_20874,N_20853);
xnor U21135 (N_21135,N_20800,N_20851);
or U21136 (N_21136,N_20812,N_20944);
xor U21137 (N_21137,N_20756,N_20991);
nor U21138 (N_21138,N_20832,N_20823);
nor U21139 (N_21139,N_20848,N_20868);
nand U21140 (N_21140,N_20941,N_20874);
xor U21141 (N_21141,N_20954,N_20961);
and U21142 (N_21142,N_20991,N_20961);
or U21143 (N_21143,N_20879,N_20945);
nor U21144 (N_21144,N_20845,N_20878);
nand U21145 (N_21145,N_20840,N_20760);
or U21146 (N_21146,N_20826,N_20872);
or U21147 (N_21147,N_20899,N_20996);
nor U21148 (N_21148,N_20909,N_20840);
nor U21149 (N_21149,N_20917,N_20861);
nand U21150 (N_21150,N_20885,N_20789);
or U21151 (N_21151,N_20898,N_20883);
or U21152 (N_21152,N_20892,N_20958);
and U21153 (N_21153,N_20932,N_20751);
and U21154 (N_21154,N_20998,N_20775);
and U21155 (N_21155,N_20925,N_20930);
xor U21156 (N_21156,N_20796,N_20998);
xor U21157 (N_21157,N_20842,N_20920);
or U21158 (N_21158,N_20816,N_20920);
xnor U21159 (N_21159,N_20891,N_20831);
or U21160 (N_21160,N_20817,N_20806);
and U21161 (N_21161,N_20803,N_20889);
and U21162 (N_21162,N_20852,N_20966);
and U21163 (N_21163,N_20795,N_20953);
and U21164 (N_21164,N_20887,N_20909);
or U21165 (N_21165,N_20924,N_20998);
and U21166 (N_21166,N_20899,N_20890);
nor U21167 (N_21167,N_20947,N_20909);
nor U21168 (N_21168,N_20896,N_20753);
nand U21169 (N_21169,N_20938,N_20997);
nor U21170 (N_21170,N_20802,N_20806);
xnor U21171 (N_21171,N_20840,N_20774);
nor U21172 (N_21172,N_20768,N_20939);
xnor U21173 (N_21173,N_20790,N_20839);
nand U21174 (N_21174,N_20784,N_20933);
nor U21175 (N_21175,N_20936,N_20980);
xnor U21176 (N_21176,N_20910,N_20964);
and U21177 (N_21177,N_20895,N_20838);
and U21178 (N_21178,N_20932,N_20979);
nand U21179 (N_21179,N_20798,N_20825);
nor U21180 (N_21180,N_20907,N_20950);
or U21181 (N_21181,N_20874,N_20978);
xor U21182 (N_21182,N_20936,N_20848);
or U21183 (N_21183,N_20840,N_20843);
nor U21184 (N_21184,N_20958,N_20974);
and U21185 (N_21185,N_20900,N_20808);
and U21186 (N_21186,N_20882,N_20789);
nand U21187 (N_21187,N_20806,N_20974);
nand U21188 (N_21188,N_20932,N_20870);
and U21189 (N_21189,N_20898,N_20787);
xor U21190 (N_21190,N_20887,N_20914);
nand U21191 (N_21191,N_20750,N_20764);
and U21192 (N_21192,N_20784,N_20770);
nand U21193 (N_21193,N_20955,N_20917);
nor U21194 (N_21194,N_20890,N_20934);
or U21195 (N_21195,N_20760,N_20964);
nand U21196 (N_21196,N_20832,N_20881);
xor U21197 (N_21197,N_20806,N_20907);
nor U21198 (N_21198,N_20925,N_20768);
nand U21199 (N_21199,N_20773,N_20954);
and U21200 (N_21200,N_20900,N_20971);
nand U21201 (N_21201,N_20943,N_20890);
nand U21202 (N_21202,N_20829,N_20806);
nand U21203 (N_21203,N_20794,N_20938);
xor U21204 (N_21204,N_20805,N_20753);
and U21205 (N_21205,N_20760,N_20945);
nor U21206 (N_21206,N_20938,N_20907);
nand U21207 (N_21207,N_20883,N_20762);
or U21208 (N_21208,N_20920,N_20953);
nor U21209 (N_21209,N_20765,N_20855);
and U21210 (N_21210,N_20842,N_20841);
and U21211 (N_21211,N_20943,N_20796);
or U21212 (N_21212,N_20852,N_20801);
nand U21213 (N_21213,N_20892,N_20751);
nand U21214 (N_21214,N_20788,N_20862);
nand U21215 (N_21215,N_20808,N_20813);
xor U21216 (N_21216,N_20864,N_20844);
and U21217 (N_21217,N_20760,N_20997);
xnor U21218 (N_21218,N_20840,N_20789);
or U21219 (N_21219,N_20995,N_20983);
xor U21220 (N_21220,N_20985,N_20947);
nor U21221 (N_21221,N_20924,N_20796);
nor U21222 (N_21222,N_20985,N_20997);
and U21223 (N_21223,N_20959,N_20773);
xor U21224 (N_21224,N_20841,N_20924);
nor U21225 (N_21225,N_20873,N_20823);
nor U21226 (N_21226,N_20752,N_20939);
nand U21227 (N_21227,N_20759,N_20800);
nor U21228 (N_21228,N_20940,N_20908);
and U21229 (N_21229,N_20986,N_20778);
nand U21230 (N_21230,N_20885,N_20839);
nor U21231 (N_21231,N_20800,N_20994);
or U21232 (N_21232,N_20846,N_20869);
nand U21233 (N_21233,N_20944,N_20955);
and U21234 (N_21234,N_20986,N_20992);
and U21235 (N_21235,N_20782,N_20917);
and U21236 (N_21236,N_20826,N_20908);
and U21237 (N_21237,N_20786,N_20868);
xor U21238 (N_21238,N_20923,N_20797);
nand U21239 (N_21239,N_20965,N_20834);
xnor U21240 (N_21240,N_20833,N_20984);
or U21241 (N_21241,N_20990,N_20783);
or U21242 (N_21242,N_20774,N_20918);
nor U21243 (N_21243,N_20953,N_20865);
and U21244 (N_21244,N_20997,N_20852);
nor U21245 (N_21245,N_20925,N_20923);
xor U21246 (N_21246,N_20899,N_20896);
and U21247 (N_21247,N_20854,N_20955);
nand U21248 (N_21248,N_20897,N_20825);
xor U21249 (N_21249,N_20984,N_20821);
nand U21250 (N_21250,N_21207,N_21112);
or U21251 (N_21251,N_21167,N_21211);
xnor U21252 (N_21252,N_21005,N_21230);
nand U21253 (N_21253,N_21198,N_21091);
nand U21254 (N_21254,N_21032,N_21035);
and U21255 (N_21255,N_21240,N_21241);
nor U21256 (N_21256,N_21131,N_21093);
and U21257 (N_21257,N_21094,N_21084);
nor U21258 (N_21258,N_21036,N_21164);
or U21259 (N_21259,N_21182,N_21158);
xor U21260 (N_21260,N_21090,N_21049);
or U21261 (N_21261,N_21234,N_21119);
nor U21262 (N_21262,N_21033,N_21030);
or U21263 (N_21263,N_21161,N_21008);
and U21264 (N_21264,N_21229,N_21059);
nand U21265 (N_21265,N_21097,N_21022);
xnor U21266 (N_21266,N_21102,N_21144);
xor U21267 (N_21267,N_21141,N_21219);
nand U21268 (N_21268,N_21203,N_21130);
or U21269 (N_21269,N_21075,N_21154);
and U21270 (N_21270,N_21007,N_21125);
nor U21271 (N_21271,N_21113,N_21047);
xor U21272 (N_21272,N_21108,N_21222);
xnor U21273 (N_21273,N_21180,N_21175);
xor U21274 (N_21274,N_21089,N_21146);
nand U21275 (N_21275,N_21124,N_21190);
or U21276 (N_21276,N_21208,N_21233);
or U21277 (N_21277,N_21103,N_21074);
nor U21278 (N_21278,N_21128,N_21186);
or U21279 (N_21279,N_21053,N_21083);
or U21280 (N_21280,N_21012,N_21137);
nand U21281 (N_21281,N_21179,N_21026);
nor U21282 (N_21282,N_21189,N_21244);
or U21283 (N_21283,N_21236,N_21187);
and U21284 (N_21284,N_21243,N_21088);
nor U21285 (N_21285,N_21153,N_21016);
or U21286 (N_21286,N_21065,N_21212);
nor U21287 (N_21287,N_21028,N_21239);
nor U21288 (N_21288,N_21126,N_21087);
nand U21289 (N_21289,N_21117,N_21116);
nor U21290 (N_21290,N_21148,N_21226);
nand U21291 (N_21291,N_21122,N_21041);
or U21292 (N_21292,N_21004,N_21155);
or U21293 (N_21293,N_21058,N_21051);
xor U21294 (N_21294,N_21159,N_21216);
nor U21295 (N_21295,N_21095,N_21199);
nand U21296 (N_21296,N_21101,N_21066);
or U21297 (N_21297,N_21168,N_21061);
or U21298 (N_21298,N_21152,N_21062);
or U21299 (N_21299,N_21224,N_21021);
xor U21300 (N_21300,N_21118,N_21092);
and U21301 (N_21301,N_21225,N_21071);
nand U21302 (N_21302,N_21185,N_21178);
or U21303 (N_21303,N_21166,N_21121);
nor U21304 (N_21304,N_21143,N_21115);
or U21305 (N_21305,N_21214,N_21248);
nand U21306 (N_21306,N_21184,N_21160);
or U21307 (N_21307,N_21165,N_21170);
nand U21308 (N_21308,N_21015,N_21191);
or U21309 (N_21309,N_21150,N_21157);
or U21310 (N_21310,N_21140,N_21106);
and U21311 (N_21311,N_21023,N_21055);
or U21312 (N_21312,N_21238,N_21162);
nand U21313 (N_21313,N_21034,N_21227);
xor U21314 (N_21314,N_21018,N_21046);
and U21315 (N_21315,N_21001,N_21109);
nor U21316 (N_21316,N_21174,N_21242);
xnor U21317 (N_21317,N_21194,N_21070);
xnor U21318 (N_21318,N_21151,N_21200);
xnor U21319 (N_21319,N_21085,N_21134);
or U21320 (N_21320,N_21006,N_21147);
and U21321 (N_21321,N_21024,N_21223);
nand U21322 (N_21322,N_21042,N_21107);
xnor U21323 (N_21323,N_21082,N_21086);
nor U21324 (N_21324,N_21218,N_21120);
nand U21325 (N_21325,N_21081,N_21247);
or U21326 (N_21326,N_21073,N_21017);
or U21327 (N_21327,N_21000,N_21176);
nand U21328 (N_21328,N_21009,N_21209);
or U21329 (N_21329,N_21213,N_21079);
xnor U21330 (N_21330,N_21098,N_21099);
nor U21331 (N_21331,N_21056,N_21245);
or U21332 (N_21332,N_21169,N_21052);
nor U21333 (N_21333,N_21249,N_21206);
and U21334 (N_21334,N_21096,N_21123);
nor U21335 (N_21335,N_21132,N_21172);
nand U21336 (N_21336,N_21135,N_21156);
and U21337 (N_21337,N_21020,N_21193);
nand U21338 (N_21338,N_21142,N_21205);
nor U21339 (N_21339,N_21011,N_21063);
nor U21340 (N_21340,N_21068,N_21013);
nand U21341 (N_21341,N_21138,N_21003);
nand U21342 (N_21342,N_21067,N_21171);
and U21343 (N_21343,N_21105,N_21215);
nor U21344 (N_21344,N_21204,N_21183);
and U21345 (N_21345,N_21010,N_21043);
or U21346 (N_21346,N_21111,N_21181);
nor U21347 (N_21347,N_21202,N_21235);
nor U21348 (N_21348,N_21192,N_21031);
nor U21349 (N_21349,N_21054,N_21195);
nand U21350 (N_21350,N_21237,N_21136);
nand U21351 (N_21351,N_21228,N_21027);
nand U21352 (N_21352,N_21173,N_21076);
nor U21353 (N_21353,N_21045,N_21014);
and U21354 (N_21354,N_21040,N_21114);
or U21355 (N_21355,N_21078,N_21069);
xor U21356 (N_21356,N_21246,N_21197);
xor U21357 (N_21357,N_21231,N_21057);
or U21358 (N_21358,N_21196,N_21100);
xnor U21359 (N_21359,N_21232,N_21129);
and U21360 (N_21360,N_21037,N_21110);
nand U21361 (N_21361,N_21133,N_21077);
and U21362 (N_21362,N_21050,N_21201);
and U21363 (N_21363,N_21025,N_21210);
and U21364 (N_21364,N_21044,N_21019);
and U21365 (N_21365,N_21039,N_21177);
xnor U21366 (N_21366,N_21217,N_21002);
nor U21367 (N_21367,N_21072,N_21127);
nor U21368 (N_21368,N_21188,N_21029);
and U21369 (N_21369,N_21145,N_21064);
nor U21370 (N_21370,N_21221,N_21220);
and U21371 (N_21371,N_21149,N_21038);
nand U21372 (N_21372,N_21048,N_21060);
xnor U21373 (N_21373,N_21139,N_21163);
nor U21374 (N_21374,N_21080,N_21104);
xor U21375 (N_21375,N_21161,N_21005);
nor U21376 (N_21376,N_21099,N_21146);
nor U21377 (N_21377,N_21054,N_21013);
xor U21378 (N_21378,N_21033,N_21096);
xnor U21379 (N_21379,N_21107,N_21013);
xnor U21380 (N_21380,N_21119,N_21049);
or U21381 (N_21381,N_21209,N_21197);
and U21382 (N_21382,N_21183,N_21201);
xnor U21383 (N_21383,N_21192,N_21191);
and U21384 (N_21384,N_21162,N_21090);
nor U21385 (N_21385,N_21195,N_21052);
and U21386 (N_21386,N_21208,N_21029);
or U21387 (N_21387,N_21199,N_21059);
nand U21388 (N_21388,N_21081,N_21193);
nor U21389 (N_21389,N_21135,N_21073);
xor U21390 (N_21390,N_21060,N_21243);
and U21391 (N_21391,N_21102,N_21085);
xor U21392 (N_21392,N_21061,N_21053);
or U21393 (N_21393,N_21119,N_21070);
and U21394 (N_21394,N_21072,N_21065);
nor U21395 (N_21395,N_21140,N_21021);
xor U21396 (N_21396,N_21127,N_21115);
nand U21397 (N_21397,N_21019,N_21243);
nand U21398 (N_21398,N_21089,N_21064);
xnor U21399 (N_21399,N_21140,N_21138);
nor U21400 (N_21400,N_21067,N_21005);
xnor U21401 (N_21401,N_21229,N_21103);
nor U21402 (N_21402,N_21131,N_21163);
nor U21403 (N_21403,N_21195,N_21017);
nand U21404 (N_21404,N_21112,N_21135);
nor U21405 (N_21405,N_21029,N_21138);
or U21406 (N_21406,N_21066,N_21086);
and U21407 (N_21407,N_21190,N_21180);
and U21408 (N_21408,N_21078,N_21244);
and U21409 (N_21409,N_21198,N_21189);
nand U21410 (N_21410,N_21076,N_21247);
and U21411 (N_21411,N_21051,N_21130);
or U21412 (N_21412,N_21104,N_21135);
or U21413 (N_21413,N_21221,N_21119);
nor U21414 (N_21414,N_21065,N_21135);
nand U21415 (N_21415,N_21003,N_21139);
nand U21416 (N_21416,N_21168,N_21219);
nor U21417 (N_21417,N_21027,N_21141);
xnor U21418 (N_21418,N_21040,N_21081);
nor U21419 (N_21419,N_21154,N_21006);
or U21420 (N_21420,N_21038,N_21008);
xnor U21421 (N_21421,N_21038,N_21097);
or U21422 (N_21422,N_21195,N_21012);
nand U21423 (N_21423,N_21173,N_21110);
xnor U21424 (N_21424,N_21017,N_21157);
nand U21425 (N_21425,N_21238,N_21042);
or U21426 (N_21426,N_21226,N_21072);
nor U21427 (N_21427,N_21146,N_21091);
xnor U21428 (N_21428,N_21175,N_21188);
or U21429 (N_21429,N_21086,N_21148);
nor U21430 (N_21430,N_21239,N_21070);
xor U21431 (N_21431,N_21219,N_21043);
and U21432 (N_21432,N_21120,N_21008);
nor U21433 (N_21433,N_21043,N_21012);
xor U21434 (N_21434,N_21069,N_21055);
nor U21435 (N_21435,N_21139,N_21065);
and U21436 (N_21436,N_21191,N_21195);
and U21437 (N_21437,N_21207,N_21177);
nand U21438 (N_21438,N_21097,N_21169);
nor U21439 (N_21439,N_21172,N_21146);
nand U21440 (N_21440,N_21028,N_21196);
nor U21441 (N_21441,N_21014,N_21007);
nor U21442 (N_21442,N_21179,N_21098);
and U21443 (N_21443,N_21214,N_21126);
xor U21444 (N_21444,N_21031,N_21167);
nand U21445 (N_21445,N_21009,N_21026);
and U21446 (N_21446,N_21020,N_21101);
nand U21447 (N_21447,N_21242,N_21155);
xor U21448 (N_21448,N_21028,N_21174);
and U21449 (N_21449,N_21107,N_21175);
or U21450 (N_21450,N_21190,N_21123);
or U21451 (N_21451,N_21107,N_21002);
or U21452 (N_21452,N_21142,N_21047);
and U21453 (N_21453,N_21077,N_21165);
or U21454 (N_21454,N_21193,N_21088);
nor U21455 (N_21455,N_21169,N_21215);
and U21456 (N_21456,N_21249,N_21031);
and U21457 (N_21457,N_21246,N_21241);
or U21458 (N_21458,N_21056,N_21237);
or U21459 (N_21459,N_21196,N_21077);
xor U21460 (N_21460,N_21138,N_21230);
xnor U21461 (N_21461,N_21132,N_21221);
xnor U21462 (N_21462,N_21230,N_21218);
xnor U21463 (N_21463,N_21034,N_21137);
or U21464 (N_21464,N_21105,N_21061);
xnor U21465 (N_21465,N_21125,N_21155);
and U21466 (N_21466,N_21036,N_21048);
nor U21467 (N_21467,N_21136,N_21123);
nor U21468 (N_21468,N_21034,N_21219);
xor U21469 (N_21469,N_21227,N_21129);
or U21470 (N_21470,N_21070,N_21153);
or U21471 (N_21471,N_21077,N_21117);
nor U21472 (N_21472,N_21090,N_21008);
nor U21473 (N_21473,N_21148,N_21038);
or U21474 (N_21474,N_21112,N_21239);
nor U21475 (N_21475,N_21217,N_21123);
or U21476 (N_21476,N_21186,N_21244);
nand U21477 (N_21477,N_21158,N_21080);
nand U21478 (N_21478,N_21077,N_21235);
and U21479 (N_21479,N_21097,N_21194);
nor U21480 (N_21480,N_21040,N_21206);
nor U21481 (N_21481,N_21151,N_21082);
and U21482 (N_21482,N_21056,N_21130);
or U21483 (N_21483,N_21220,N_21023);
nor U21484 (N_21484,N_21224,N_21071);
or U21485 (N_21485,N_21183,N_21052);
xor U21486 (N_21486,N_21073,N_21190);
nor U21487 (N_21487,N_21162,N_21050);
xnor U21488 (N_21488,N_21193,N_21024);
nor U21489 (N_21489,N_21210,N_21211);
or U21490 (N_21490,N_21052,N_21119);
nand U21491 (N_21491,N_21009,N_21182);
xor U21492 (N_21492,N_21064,N_21207);
xor U21493 (N_21493,N_21083,N_21009);
xor U21494 (N_21494,N_21125,N_21096);
nor U21495 (N_21495,N_21101,N_21184);
nor U21496 (N_21496,N_21119,N_21016);
nor U21497 (N_21497,N_21172,N_21044);
nand U21498 (N_21498,N_21131,N_21011);
and U21499 (N_21499,N_21048,N_21038);
nand U21500 (N_21500,N_21389,N_21416);
xor U21501 (N_21501,N_21273,N_21424);
and U21502 (N_21502,N_21284,N_21276);
nor U21503 (N_21503,N_21368,N_21342);
nor U21504 (N_21504,N_21443,N_21381);
and U21505 (N_21505,N_21252,N_21287);
xnor U21506 (N_21506,N_21331,N_21433);
nor U21507 (N_21507,N_21417,N_21472);
xor U21508 (N_21508,N_21267,N_21322);
nand U21509 (N_21509,N_21492,N_21372);
xor U21510 (N_21510,N_21312,N_21283);
or U21511 (N_21511,N_21373,N_21401);
xor U21512 (N_21512,N_21423,N_21396);
nand U21513 (N_21513,N_21409,N_21386);
nand U21514 (N_21514,N_21347,N_21338);
xnor U21515 (N_21515,N_21364,N_21297);
or U21516 (N_21516,N_21366,N_21350);
xor U21517 (N_21517,N_21304,N_21448);
and U21518 (N_21518,N_21463,N_21337);
nor U21519 (N_21519,N_21392,N_21482);
nand U21520 (N_21520,N_21407,N_21324);
xor U21521 (N_21521,N_21285,N_21481);
or U21522 (N_21522,N_21260,N_21346);
or U21523 (N_21523,N_21288,N_21329);
and U21524 (N_21524,N_21311,N_21266);
nand U21525 (N_21525,N_21484,N_21320);
and U21526 (N_21526,N_21441,N_21485);
nor U21527 (N_21527,N_21442,N_21315);
nand U21528 (N_21528,N_21460,N_21480);
nor U21529 (N_21529,N_21325,N_21253);
nor U21530 (N_21530,N_21499,N_21357);
xnor U21531 (N_21531,N_21387,N_21299);
nand U21532 (N_21532,N_21292,N_21457);
nor U21533 (N_21533,N_21279,N_21272);
nor U21534 (N_21534,N_21493,N_21393);
xor U21535 (N_21535,N_21256,N_21374);
nor U21536 (N_21536,N_21413,N_21455);
nand U21537 (N_21537,N_21269,N_21388);
and U21538 (N_21538,N_21470,N_21486);
or U21539 (N_21539,N_21262,N_21384);
and U21540 (N_21540,N_21349,N_21420);
nand U21541 (N_21541,N_21425,N_21362);
and U21542 (N_21542,N_21345,N_21308);
xor U21543 (N_21543,N_21278,N_21497);
nor U21544 (N_21544,N_21261,N_21487);
nand U21545 (N_21545,N_21316,N_21453);
nor U21546 (N_21546,N_21437,N_21495);
nand U21547 (N_21547,N_21264,N_21302);
and U21548 (N_21548,N_21479,N_21319);
nand U21549 (N_21549,N_21268,N_21490);
and U21550 (N_21550,N_21491,N_21395);
xnor U21551 (N_21551,N_21469,N_21456);
nand U21552 (N_21552,N_21418,N_21277);
or U21553 (N_21553,N_21436,N_21390);
or U21554 (N_21554,N_21294,N_21430);
xnor U21555 (N_21555,N_21280,N_21363);
nor U21556 (N_21556,N_21310,N_21477);
nand U21557 (N_21557,N_21449,N_21377);
or U21558 (N_21558,N_21429,N_21348);
or U21559 (N_21559,N_21394,N_21274);
or U21560 (N_21560,N_21414,N_21265);
and U21561 (N_21561,N_21452,N_21307);
nand U21562 (N_21562,N_21333,N_21353);
and U21563 (N_21563,N_21400,N_21286);
xor U21564 (N_21564,N_21376,N_21275);
xor U21565 (N_21565,N_21451,N_21444);
nand U21566 (N_21566,N_21257,N_21271);
or U21567 (N_21567,N_21295,N_21270);
nand U21568 (N_21568,N_21422,N_21440);
nand U21569 (N_21569,N_21411,N_21447);
nor U21570 (N_21570,N_21334,N_21321);
and U21571 (N_21571,N_21313,N_21309);
and U21572 (N_21572,N_21306,N_21323);
nand U21573 (N_21573,N_21359,N_21370);
nor U21574 (N_21574,N_21300,N_21379);
or U21575 (N_21575,N_21317,N_21415);
nor U21576 (N_21576,N_21406,N_21468);
or U21577 (N_21577,N_21314,N_21459);
nor U21578 (N_21578,N_21466,N_21410);
nor U21579 (N_21579,N_21475,N_21450);
or U21580 (N_21580,N_21467,N_21296);
nor U21581 (N_21581,N_21385,N_21361);
and U21582 (N_21582,N_21305,N_21426);
or U21583 (N_21583,N_21496,N_21258);
or U21584 (N_21584,N_21371,N_21369);
and U21585 (N_21585,N_21488,N_21378);
xor U21586 (N_21586,N_21340,N_21489);
or U21587 (N_21587,N_21335,N_21397);
or U21588 (N_21588,N_21291,N_21365);
or U21589 (N_21589,N_21408,N_21399);
and U21590 (N_21590,N_21380,N_21458);
or U21591 (N_21591,N_21259,N_21398);
xnor U21592 (N_21592,N_21327,N_21328);
nor U21593 (N_21593,N_21356,N_21427);
or U21594 (N_21594,N_21464,N_21344);
or U21595 (N_21595,N_21498,N_21251);
and U21596 (N_21596,N_21465,N_21355);
and U21597 (N_21597,N_21339,N_21494);
and U21598 (N_21598,N_21434,N_21330);
or U21599 (N_21599,N_21383,N_21461);
nand U21600 (N_21600,N_21419,N_21412);
nand U21601 (N_21601,N_21336,N_21382);
nand U21602 (N_21602,N_21352,N_21405);
xor U21603 (N_21603,N_21250,N_21298);
xor U21604 (N_21604,N_21332,N_21293);
nor U21605 (N_21605,N_21282,N_21476);
or U21606 (N_21606,N_21303,N_21255);
and U21607 (N_21607,N_21326,N_21290);
nor U21608 (N_21608,N_21471,N_21289);
and U21609 (N_21609,N_21351,N_21254);
xor U21610 (N_21610,N_21478,N_21341);
nand U21611 (N_21611,N_21281,N_21428);
nor U21612 (N_21612,N_21438,N_21462);
and U21613 (N_21613,N_21318,N_21403);
xor U21614 (N_21614,N_21421,N_21431);
xor U21615 (N_21615,N_21360,N_21435);
xor U21616 (N_21616,N_21263,N_21375);
and U21617 (N_21617,N_21454,N_21483);
nand U21618 (N_21618,N_21404,N_21354);
nand U21619 (N_21619,N_21445,N_21391);
nor U21620 (N_21620,N_21432,N_21474);
and U21621 (N_21621,N_21358,N_21446);
xor U21622 (N_21622,N_21402,N_21367);
xor U21623 (N_21623,N_21301,N_21343);
nand U21624 (N_21624,N_21439,N_21473);
xnor U21625 (N_21625,N_21393,N_21274);
nand U21626 (N_21626,N_21446,N_21381);
and U21627 (N_21627,N_21425,N_21316);
nand U21628 (N_21628,N_21419,N_21446);
xor U21629 (N_21629,N_21497,N_21365);
nand U21630 (N_21630,N_21377,N_21443);
xnor U21631 (N_21631,N_21469,N_21387);
xnor U21632 (N_21632,N_21370,N_21462);
or U21633 (N_21633,N_21274,N_21280);
nand U21634 (N_21634,N_21383,N_21422);
and U21635 (N_21635,N_21318,N_21408);
nand U21636 (N_21636,N_21257,N_21337);
nand U21637 (N_21637,N_21391,N_21494);
nor U21638 (N_21638,N_21413,N_21492);
xnor U21639 (N_21639,N_21325,N_21447);
and U21640 (N_21640,N_21313,N_21338);
nor U21641 (N_21641,N_21436,N_21295);
nand U21642 (N_21642,N_21304,N_21257);
nor U21643 (N_21643,N_21346,N_21429);
xnor U21644 (N_21644,N_21447,N_21306);
and U21645 (N_21645,N_21307,N_21394);
xor U21646 (N_21646,N_21313,N_21262);
nand U21647 (N_21647,N_21277,N_21349);
or U21648 (N_21648,N_21405,N_21367);
and U21649 (N_21649,N_21408,N_21322);
nand U21650 (N_21650,N_21337,N_21449);
and U21651 (N_21651,N_21311,N_21290);
nor U21652 (N_21652,N_21342,N_21325);
nand U21653 (N_21653,N_21461,N_21413);
xor U21654 (N_21654,N_21308,N_21301);
nand U21655 (N_21655,N_21270,N_21387);
and U21656 (N_21656,N_21366,N_21298);
xor U21657 (N_21657,N_21376,N_21314);
nand U21658 (N_21658,N_21477,N_21441);
nor U21659 (N_21659,N_21418,N_21396);
and U21660 (N_21660,N_21378,N_21286);
and U21661 (N_21661,N_21470,N_21256);
or U21662 (N_21662,N_21470,N_21434);
xor U21663 (N_21663,N_21393,N_21325);
xor U21664 (N_21664,N_21269,N_21403);
xnor U21665 (N_21665,N_21428,N_21352);
or U21666 (N_21666,N_21413,N_21498);
xnor U21667 (N_21667,N_21253,N_21390);
or U21668 (N_21668,N_21399,N_21280);
or U21669 (N_21669,N_21329,N_21365);
xor U21670 (N_21670,N_21447,N_21261);
nand U21671 (N_21671,N_21431,N_21291);
nor U21672 (N_21672,N_21394,N_21301);
xnor U21673 (N_21673,N_21449,N_21386);
or U21674 (N_21674,N_21357,N_21474);
xnor U21675 (N_21675,N_21460,N_21415);
nand U21676 (N_21676,N_21401,N_21413);
nor U21677 (N_21677,N_21447,N_21320);
nand U21678 (N_21678,N_21387,N_21352);
and U21679 (N_21679,N_21364,N_21317);
nor U21680 (N_21680,N_21373,N_21488);
nor U21681 (N_21681,N_21293,N_21390);
nor U21682 (N_21682,N_21383,N_21282);
xnor U21683 (N_21683,N_21453,N_21250);
and U21684 (N_21684,N_21387,N_21394);
and U21685 (N_21685,N_21260,N_21311);
nor U21686 (N_21686,N_21286,N_21331);
nand U21687 (N_21687,N_21277,N_21495);
nand U21688 (N_21688,N_21377,N_21339);
nand U21689 (N_21689,N_21484,N_21367);
and U21690 (N_21690,N_21459,N_21443);
or U21691 (N_21691,N_21266,N_21297);
nand U21692 (N_21692,N_21472,N_21477);
xor U21693 (N_21693,N_21275,N_21286);
nor U21694 (N_21694,N_21490,N_21250);
nand U21695 (N_21695,N_21362,N_21499);
nand U21696 (N_21696,N_21307,N_21354);
nor U21697 (N_21697,N_21495,N_21349);
xor U21698 (N_21698,N_21482,N_21371);
xor U21699 (N_21699,N_21409,N_21499);
xnor U21700 (N_21700,N_21340,N_21254);
nand U21701 (N_21701,N_21356,N_21300);
nor U21702 (N_21702,N_21265,N_21397);
or U21703 (N_21703,N_21345,N_21359);
nand U21704 (N_21704,N_21426,N_21419);
and U21705 (N_21705,N_21415,N_21301);
xnor U21706 (N_21706,N_21482,N_21346);
and U21707 (N_21707,N_21474,N_21312);
xor U21708 (N_21708,N_21425,N_21255);
or U21709 (N_21709,N_21349,N_21280);
xor U21710 (N_21710,N_21404,N_21342);
nand U21711 (N_21711,N_21378,N_21386);
nand U21712 (N_21712,N_21482,N_21362);
nor U21713 (N_21713,N_21266,N_21336);
or U21714 (N_21714,N_21255,N_21458);
or U21715 (N_21715,N_21400,N_21458);
and U21716 (N_21716,N_21478,N_21287);
or U21717 (N_21717,N_21416,N_21277);
nand U21718 (N_21718,N_21403,N_21441);
nand U21719 (N_21719,N_21396,N_21288);
and U21720 (N_21720,N_21479,N_21315);
and U21721 (N_21721,N_21327,N_21388);
nand U21722 (N_21722,N_21416,N_21438);
nor U21723 (N_21723,N_21274,N_21251);
and U21724 (N_21724,N_21455,N_21323);
or U21725 (N_21725,N_21312,N_21451);
xor U21726 (N_21726,N_21343,N_21467);
and U21727 (N_21727,N_21463,N_21498);
nand U21728 (N_21728,N_21275,N_21281);
xor U21729 (N_21729,N_21311,N_21469);
or U21730 (N_21730,N_21450,N_21314);
nor U21731 (N_21731,N_21296,N_21379);
nand U21732 (N_21732,N_21392,N_21371);
nand U21733 (N_21733,N_21456,N_21262);
and U21734 (N_21734,N_21425,N_21392);
xnor U21735 (N_21735,N_21252,N_21335);
and U21736 (N_21736,N_21260,N_21436);
nand U21737 (N_21737,N_21386,N_21447);
nand U21738 (N_21738,N_21415,N_21440);
nand U21739 (N_21739,N_21359,N_21324);
or U21740 (N_21740,N_21416,N_21376);
or U21741 (N_21741,N_21454,N_21317);
nand U21742 (N_21742,N_21389,N_21335);
or U21743 (N_21743,N_21362,N_21290);
or U21744 (N_21744,N_21364,N_21406);
or U21745 (N_21745,N_21459,N_21352);
or U21746 (N_21746,N_21495,N_21496);
or U21747 (N_21747,N_21435,N_21375);
nor U21748 (N_21748,N_21263,N_21498);
nor U21749 (N_21749,N_21274,N_21415);
xor U21750 (N_21750,N_21582,N_21526);
or U21751 (N_21751,N_21665,N_21550);
or U21752 (N_21752,N_21622,N_21643);
xnor U21753 (N_21753,N_21569,N_21630);
nor U21754 (N_21754,N_21577,N_21590);
nor U21755 (N_21755,N_21508,N_21707);
and U21756 (N_21756,N_21558,N_21517);
or U21757 (N_21757,N_21518,N_21657);
nor U21758 (N_21758,N_21604,N_21602);
or U21759 (N_21759,N_21715,N_21731);
or U21760 (N_21760,N_21624,N_21658);
or U21761 (N_21761,N_21685,N_21503);
xnor U21762 (N_21762,N_21573,N_21677);
xor U21763 (N_21763,N_21509,N_21721);
nand U21764 (N_21764,N_21530,N_21554);
xnor U21765 (N_21765,N_21571,N_21623);
nand U21766 (N_21766,N_21686,N_21559);
and U21767 (N_21767,N_21626,N_21621);
and U21768 (N_21768,N_21676,N_21709);
nand U21769 (N_21769,N_21639,N_21565);
nor U21770 (N_21770,N_21638,N_21738);
and U21771 (N_21771,N_21633,N_21730);
nand U21772 (N_21772,N_21743,N_21524);
nor U21773 (N_21773,N_21544,N_21516);
nand U21774 (N_21774,N_21732,N_21549);
and U21775 (N_21775,N_21736,N_21652);
nand U21776 (N_21776,N_21596,N_21695);
nor U21777 (N_21777,N_21661,N_21586);
and U21778 (N_21778,N_21741,N_21555);
nand U21779 (N_21779,N_21522,N_21728);
xnor U21780 (N_21780,N_21607,N_21581);
and U21781 (N_21781,N_21616,N_21647);
xnor U21782 (N_21782,N_21557,N_21696);
xnor U21783 (N_21783,N_21748,N_21585);
xnor U21784 (N_21784,N_21689,N_21690);
xor U21785 (N_21785,N_21574,N_21556);
nand U21786 (N_21786,N_21603,N_21575);
nor U21787 (N_21787,N_21663,N_21649);
nand U21788 (N_21788,N_21561,N_21727);
xnor U21789 (N_21789,N_21683,N_21505);
nand U21790 (N_21790,N_21668,N_21708);
and U21791 (N_21791,N_21651,N_21700);
xor U21792 (N_21792,N_21594,N_21535);
xor U21793 (N_21793,N_21742,N_21546);
and U21794 (N_21794,N_21548,N_21547);
or U21795 (N_21795,N_21667,N_21655);
nand U21796 (N_21796,N_21591,N_21684);
nor U21797 (N_21797,N_21629,N_21606);
and U21798 (N_21798,N_21560,N_21619);
xor U21799 (N_21799,N_21527,N_21501);
nand U21800 (N_21800,N_21678,N_21679);
or U21801 (N_21801,N_21553,N_21609);
or U21802 (N_21802,N_21567,N_21618);
xnor U21803 (N_21803,N_21739,N_21510);
nor U21804 (N_21804,N_21611,N_21566);
or U21805 (N_21805,N_21534,N_21533);
or U21806 (N_21806,N_21694,N_21515);
and U21807 (N_21807,N_21514,N_21726);
xor U21808 (N_21808,N_21697,N_21541);
and U21809 (N_21809,N_21744,N_21532);
or U21810 (N_21810,N_21674,N_21712);
nor U21811 (N_21811,N_21713,N_21507);
xor U21812 (N_21812,N_21531,N_21664);
nor U21813 (N_21813,N_21592,N_21576);
xnor U21814 (N_21814,N_21710,N_21543);
nand U21815 (N_21815,N_21737,N_21552);
nand U21816 (N_21816,N_21698,N_21653);
and U21817 (N_21817,N_21660,N_21579);
nand U21818 (N_21818,N_21650,N_21570);
nor U21819 (N_21819,N_21646,N_21719);
nor U21820 (N_21820,N_21687,N_21589);
nor U21821 (N_21821,N_21529,N_21747);
and U21822 (N_21822,N_21680,N_21714);
nor U21823 (N_21823,N_21613,N_21513);
and U21824 (N_21824,N_21627,N_21625);
nor U21825 (N_21825,N_21733,N_21724);
xnor U21826 (N_21826,N_21703,N_21662);
nor U21827 (N_21827,N_21669,N_21525);
nor U21828 (N_21828,N_21631,N_21745);
or U21829 (N_21829,N_21608,N_21578);
nor U21830 (N_21830,N_21614,N_21654);
nor U21831 (N_21831,N_21598,N_21628);
or U21832 (N_21832,N_21634,N_21644);
and U21833 (N_21833,N_21682,N_21722);
xnor U21834 (N_21834,N_21540,N_21641);
nand U21835 (N_21835,N_21520,N_21672);
nand U21836 (N_21836,N_21615,N_21718);
or U21837 (N_21837,N_21562,N_21610);
or U21838 (N_21838,N_21681,N_21725);
xor U21839 (N_21839,N_21572,N_21519);
and U21840 (N_21840,N_21723,N_21666);
xor U21841 (N_21841,N_21563,N_21706);
nor U21842 (N_21842,N_21605,N_21512);
nand U21843 (N_21843,N_21595,N_21701);
xor U21844 (N_21844,N_21692,N_21538);
and U21845 (N_21845,N_21564,N_21716);
nor U21846 (N_21846,N_21539,N_21587);
nor U21847 (N_21847,N_21659,N_21601);
nand U21848 (N_21848,N_21599,N_21537);
nor U21849 (N_21849,N_21506,N_21521);
nor U21850 (N_21850,N_21632,N_21500);
nand U21851 (N_21851,N_21584,N_21691);
and U21852 (N_21852,N_21511,N_21597);
or U21853 (N_21853,N_21536,N_21648);
nand U21854 (N_21854,N_21528,N_21729);
or U21855 (N_21855,N_21673,N_21612);
and U21856 (N_21856,N_21568,N_21749);
and U21857 (N_21857,N_21656,N_21688);
nand U21858 (N_21858,N_21502,N_21617);
and U21859 (N_21859,N_21675,N_21545);
or U21860 (N_21860,N_21551,N_21671);
nand U21861 (N_21861,N_21735,N_21593);
and U21862 (N_21862,N_21635,N_21637);
xnor U21863 (N_21863,N_21734,N_21740);
or U21864 (N_21864,N_21702,N_21542);
xor U21865 (N_21865,N_21720,N_21704);
nand U21866 (N_21866,N_21620,N_21645);
and U21867 (N_21867,N_21523,N_21580);
or U21868 (N_21868,N_21693,N_21636);
xor U21869 (N_21869,N_21583,N_21504);
or U21870 (N_21870,N_21588,N_21705);
or U21871 (N_21871,N_21711,N_21670);
nor U21872 (N_21872,N_21746,N_21640);
or U21873 (N_21873,N_21642,N_21717);
nor U21874 (N_21874,N_21699,N_21600);
xor U21875 (N_21875,N_21529,N_21543);
and U21876 (N_21876,N_21701,N_21703);
and U21877 (N_21877,N_21658,N_21715);
nand U21878 (N_21878,N_21603,N_21667);
nand U21879 (N_21879,N_21664,N_21547);
or U21880 (N_21880,N_21536,N_21727);
xnor U21881 (N_21881,N_21604,N_21529);
xor U21882 (N_21882,N_21708,N_21570);
nor U21883 (N_21883,N_21619,N_21702);
xnor U21884 (N_21884,N_21595,N_21586);
nand U21885 (N_21885,N_21516,N_21526);
or U21886 (N_21886,N_21678,N_21649);
and U21887 (N_21887,N_21705,N_21623);
nand U21888 (N_21888,N_21600,N_21506);
xor U21889 (N_21889,N_21729,N_21658);
or U21890 (N_21890,N_21588,N_21601);
and U21891 (N_21891,N_21713,N_21601);
and U21892 (N_21892,N_21738,N_21634);
nand U21893 (N_21893,N_21714,N_21664);
and U21894 (N_21894,N_21717,N_21707);
xnor U21895 (N_21895,N_21718,N_21719);
or U21896 (N_21896,N_21714,N_21724);
nand U21897 (N_21897,N_21558,N_21736);
nand U21898 (N_21898,N_21617,N_21606);
or U21899 (N_21899,N_21737,N_21617);
nor U21900 (N_21900,N_21539,N_21566);
xnor U21901 (N_21901,N_21723,N_21556);
and U21902 (N_21902,N_21701,N_21737);
or U21903 (N_21903,N_21576,N_21728);
xor U21904 (N_21904,N_21523,N_21611);
nor U21905 (N_21905,N_21531,N_21652);
xor U21906 (N_21906,N_21513,N_21669);
nor U21907 (N_21907,N_21603,N_21528);
or U21908 (N_21908,N_21697,N_21654);
nor U21909 (N_21909,N_21568,N_21740);
nor U21910 (N_21910,N_21502,N_21711);
or U21911 (N_21911,N_21553,N_21709);
or U21912 (N_21912,N_21546,N_21618);
or U21913 (N_21913,N_21723,N_21726);
or U21914 (N_21914,N_21564,N_21536);
nor U21915 (N_21915,N_21613,N_21620);
and U21916 (N_21916,N_21628,N_21637);
or U21917 (N_21917,N_21534,N_21515);
xor U21918 (N_21918,N_21730,N_21651);
and U21919 (N_21919,N_21651,N_21568);
xnor U21920 (N_21920,N_21500,N_21620);
or U21921 (N_21921,N_21604,N_21570);
nor U21922 (N_21922,N_21598,N_21736);
or U21923 (N_21923,N_21566,N_21556);
xor U21924 (N_21924,N_21547,N_21737);
and U21925 (N_21925,N_21638,N_21678);
or U21926 (N_21926,N_21665,N_21588);
and U21927 (N_21927,N_21560,N_21575);
nand U21928 (N_21928,N_21672,N_21512);
xor U21929 (N_21929,N_21566,N_21529);
or U21930 (N_21930,N_21617,N_21697);
and U21931 (N_21931,N_21557,N_21510);
or U21932 (N_21932,N_21518,N_21547);
and U21933 (N_21933,N_21723,N_21631);
or U21934 (N_21934,N_21729,N_21686);
or U21935 (N_21935,N_21722,N_21621);
or U21936 (N_21936,N_21727,N_21518);
or U21937 (N_21937,N_21544,N_21748);
and U21938 (N_21938,N_21710,N_21741);
nand U21939 (N_21939,N_21739,N_21714);
xnor U21940 (N_21940,N_21597,N_21608);
nor U21941 (N_21941,N_21514,N_21741);
or U21942 (N_21942,N_21650,N_21683);
nor U21943 (N_21943,N_21599,N_21558);
and U21944 (N_21944,N_21567,N_21736);
or U21945 (N_21945,N_21634,N_21720);
xor U21946 (N_21946,N_21745,N_21723);
nor U21947 (N_21947,N_21517,N_21625);
xnor U21948 (N_21948,N_21521,N_21593);
or U21949 (N_21949,N_21695,N_21564);
nand U21950 (N_21950,N_21732,N_21593);
nor U21951 (N_21951,N_21686,N_21591);
nand U21952 (N_21952,N_21656,N_21615);
nand U21953 (N_21953,N_21707,N_21626);
and U21954 (N_21954,N_21614,N_21744);
nand U21955 (N_21955,N_21527,N_21609);
or U21956 (N_21956,N_21701,N_21522);
nor U21957 (N_21957,N_21508,N_21546);
and U21958 (N_21958,N_21667,N_21616);
or U21959 (N_21959,N_21707,N_21534);
xor U21960 (N_21960,N_21607,N_21578);
and U21961 (N_21961,N_21710,N_21522);
or U21962 (N_21962,N_21532,N_21646);
and U21963 (N_21963,N_21592,N_21654);
or U21964 (N_21964,N_21621,N_21607);
or U21965 (N_21965,N_21554,N_21723);
and U21966 (N_21966,N_21641,N_21737);
and U21967 (N_21967,N_21571,N_21566);
nand U21968 (N_21968,N_21609,N_21572);
xnor U21969 (N_21969,N_21691,N_21616);
nor U21970 (N_21970,N_21559,N_21503);
nor U21971 (N_21971,N_21693,N_21611);
nand U21972 (N_21972,N_21716,N_21607);
xnor U21973 (N_21973,N_21672,N_21749);
or U21974 (N_21974,N_21509,N_21661);
or U21975 (N_21975,N_21666,N_21566);
or U21976 (N_21976,N_21702,N_21535);
xnor U21977 (N_21977,N_21640,N_21590);
xor U21978 (N_21978,N_21578,N_21691);
xor U21979 (N_21979,N_21659,N_21650);
nor U21980 (N_21980,N_21731,N_21526);
xnor U21981 (N_21981,N_21516,N_21508);
xor U21982 (N_21982,N_21567,N_21645);
nor U21983 (N_21983,N_21748,N_21504);
and U21984 (N_21984,N_21683,N_21739);
nand U21985 (N_21985,N_21638,N_21719);
nor U21986 (N_21986,N_21696,N_21659);
nor U21987 (N_21987,N_21589,N_21742);
nor U21988 (N_21988,N_21525,N_21582);
nand U21989 (N_21989,N_21513,N_21530);
or U21990 (N_21990,N_21696,N_21502);
nand U21991 (N_21991,N_21530,N_21633);
xor U21992 (N_21992,N_21554,N_21727);
or U21993 (N_21993,N_21633,N_21744);
or U21994 (N_21994,N_21555,N_21719);
or U21995 (N_21995,N_21573,N_21609);
nor U21996 (N_21996,N_21535,N_21618);
nor U21997 (N_21997,N_21631,N_21689);
xor U21998 (N_21998,N_21640,N_21696);
or U21999 (N_21999,N_21533,N_21681);
nor U22000 (N_22000,N_21753,N_21994);
xnor U22001 (N_22001,N_21970,N_21864);
nor U22002 (N_22002,N_21826,N_21978);
or U22003 (N_22003,N_21906,N_21751);
xor U22004 (N_22004,N_21819,N_21984);
nor U22005 (N_22005,N_21892,N_21769);
xnor U22006 (N_22006,N_21818,N_21794);
xnor U22007 (N_22007,N_21985,N_21814);
and U22008 (N_22008,N_21950,N_21971);
and U22009 (N_22009,N_21874,N_21815);
nand U22010 (N_22010,N_21807,N_21983);
nand U22011 (N_22011,N_21841,N_21792);
nor U22012 (N_22012,N_21924,N_21925);
nand U22013 (N_22013,N_21945,N_21827);
nor U22014 (N_22014,N_21776,N_21943);
nor U22015 (N_22015,N_21833,N_21907);
xor U22016 (N_22016,N_21887,N_21796);
xor U22017 (N_22017,N_21884,N_21804);
or U22018 (N_22018,N_21850,N_21997);
nor U22019 (N_22019,N_21918,N_21834);
or U22020 (N_22020,N_21910,N_21810);
or U22021 (N_22021,N_21991,N_21846);
nor U22022 (N_22022,N_21988,N_21771);
xnor U22023 (N_22023,N_21889,N_21823);
nor U22024 (N_22024,N_21876,N_21858);
nor U22025 (N_22025,N_21806,N_21830);
and U22026 (N_22026,N_21932,N_21953);
and U22027 (N_22027,N_21966,N_21999);
and U22028 (N_22028,N_21960,N_21765);
and U22029 (N_22029,N_21852,N_21759);
nor U22030 (N_22030,N_21904,N_21940);
and U22031 (N_22031,N_21779,N_21878);
nor U22032 (N_22032,N_21798,N_21962);
or U22033 (N_22033,N_21908,N_21927);
or U22034 (N_22034,N_21800,N_21861);
and U22035 (N_22035,N_21770,N_21898);
xor U22036 (N_22036,N_21871,N_21831);
or U22037 (N_22037,N_21903,N_21885);
or U22038 (N_22038,N_21787,N_21987);
and U22039 (N_22039,N_21965,N_21901);
nand U22040 (N_22040,N_21845,N_21890);
nand U22041 (N_22041,N_21762,N_21956);
xnor U22042 (N_22042,N_21964,N_21990);
or U22043 (N_22043,N_21767,N_21877);
nor U22044 (N_22044,N_21754,N_21784);
and U22045 (N_22045,N_21774,N_21848);
nor U22046 (N_22046,N_21844,N_21855);
and U22047 (N_22047,N_21959,N_21857);
and U22048 (N_22048,N_21905,N_21808);
xor U22049 (N_22049,N_21875,N_21803);
nor U22050 (N_22050,N_21811,N_21790);
or U22051 (N_22051,N_21763,N_21926);
nand U22052 (N_22052,N_21842,N_21923);
and U22053 (N_22053,N_21851,N_21872);
nor U22054 (N_22054,N_21981,N_21828);
or U22055 (N_22055,N_21891,N_21952);
or U22056 (N_22056,N_21799,N_21882);
nor U22057 (N_22057,N_21934,N_21752);
nand U22058 (N_22058,N_21993,N_21791);
xor U22059 (N_22059,N_21941,N_21995);
nand U22060 (N_22060,N_21757,N_21942);
nor U22061 (N_22061,N_21822,N_21775);
nand U22062 (N_22062,N_21977,N_21946);
xnor U22063 (N_22063,N_21756,N_21836);
nand U22064 (N_22064,N_21860,N_21854);
nor U22065 (N_22065,N_21761,N_21972);
nand U22066 (N_22066,N_21782,N_21802);
or U22067 (N_22067,N_21768,N_21989);
and U22068 (N_22068,N_21938,N_21772);
and U22069 (N_22069,N_21829,N_21979);
or U22070 (N_22070,N_21982,N_21902);
nand U22071 (N_22071,N_21840,N_21849);
xnor U22072 (N_22072,N_21781,N_21880);
nand U22073 (N_22073,N_21760,N_21866);
xor U22074 (N_22074,N_21996,N_21967);
and U22075 (N_22075,N_21859,N_21974);
nand U22076 (N_22076,N_21937,N_21879);
nand U22077 (N_22077,N_21935,N_21912);
or U22078 (N_22078,N_21816,N_21986);
and U22079 (N_22079,N_21973,N_21963);
or U22080 (N_22080,N_21976,N_21881);
or U22081 (N_22081,N_21773,N_21980);
nor U22082 (N_22082,N_21958,N_21856);
nand U22083 (N_22083,N_21894,N_21969);
nand U22084 (N_22084,N_21788,N_21916);
xor U22085 (N_22085,N_21883,N_21886);
or U22086 (N_22086,N_21862,N_21843);
xor U22087 (N_22087,N_21931,N_21949);
nor U22088 (N_22088,N_21913,N_21939);
nand U22089 (N_22089,N_21783,N_21920);
or U22090 (N_22090,N_21915,N_21832);
nand U22091 (N_22091,N_21780,N_21928);
or U22092 (N_22092,N_21839,N_21786);
nand U22093 (N_22093,N_21936,N_21897);
nand U22094 (N_22094,N_21896,N_21930);
or U22095 (N_22095,N_21888,N_21873);
nor U22096 (N_22096,N_21863,N_21865);
and U22097 (N_22097,N_21755,N_21955);
and U22098 (N_22098,N_21801,N_21911);
nand U22099 (N_22099,N_21870,N_21805);
xor U22100 (N_22100,N_21948,N_21922);
xor U22101 (N_22101,N_21793,N_21868);
xnor U22102 (N_22102,N_21933,N_21758);
or U22103 (N_22103,N_21951,N_21824);
xnor U22104 (N_22104,N_21813,N_21992);
nand U22105 (N_22105,N_21789,N_21820);
nand U22106 (N_22106,N_21847,N_21817);
and U22107 (N_22107,N_21968,N_21821);
nand U22108 (N_22108,N_21869,N_21809);
and U22109 (N_22109,N_21853,N_21917);
nand U22110 (N_22110,N_21921,N_21895);
nor U22111 (N_22111,N_21838,N_21812);
nand U22112 (N_22112,N_21909,N_21835);
or U22113 (N_22113,N_21914,N_21778);
or U22114 (N_22114,N_21929,N_21998);
and U22115 (N_22115,N_21961,N_21750);
or U22116 (N_22116,N_21766,N_21919);
and U22117 (N_22117,N_21777,N_21944);
nor U22118 (N_22118,N_21764,N_21795);
nand U22119 (N_22119,N_21947,N_21900);
nor U22120 (N_22120,N_21954,N_21899);
or U22121 (N_22121,N_21893,N_21785);
nor U22122 (N_22122,N_21975,N_21867);
or U22123 (N_22123,N_21825,N_21957);
and U22124 (N_22124,N_21797,N_21837);
nand U22125 (N_22125,N_21951,N_21825);
nand U22126 (N_22126,N_21799,N_21922);
or U22127 (N_22127,N_21768,N_21936);
xnor U22128 (N_22128,N_21822,N_21847);
nand U22129 (N_22129,N_21944,N_21953);
nor U22130 (N_22130,N_21835,N_21896);
nor U22131 (N_22131,N_21914,N_21993);
and U22132 (N_22132,N_21831,N_21956);
and U22133 (N_22133,N_21901,N_21902);
nor U22134 (N_22134,N_21823,N_21772);
xor U22135 (N_22135,N_21917,N_21868);
and U22136 (N_22136,N_21852,N_21849);
nand U22137 (N_22137,N_21962,N_21961);
and U22138 (N_22138,N_21821,N_21850);
nand U22139 (N_22139,N_21884,N_21913);
xnor U22140 (N_22140,N_21993,N_21943);
nor U22141 (N_22141,N_21969,N_21814);
or U22142 (N_22142,N_21984,N_21809);
nor U22143 (N_22143,N_21931,N_21796);
xnor U22144 (N_22144,N_21768,N_21962);
nor U22145 (N_22145,N_21769,N_21924);
and U22146 (N_22146,N_21980,N_21896);
nand U22147 (N_22147,N_21763,N_21773);
nor U22148 (N_22148,N_21837,N_21937);
nand U22149 (N_22149,N_21817,N_21923);
nor U22150 (N_22150,N_21852,N_21877);
nor U22151 (N_22151,N_21812,N_21942);
nand U22152 (N_22152,N_21852,N_21782);
or U22153 (N_22153,N_21807,N_21770);
or U22154 (N_22154,N_21829,N_21981);
and U22155 (N_22155,N_21806,N_21819);
or U22156 (N_22156,N_21803,N_21923);
nor U22157 (N_22157,N_21837,N_21909);
xnor U22158 (N_22158,N_21963,N_21930);
and U22159 (N_22159,N_21923,N_21909);
nor U22160 (N_22160,N_21810,N_21846);
xnor U22161 (N_22161,N_21864,N_21767);
or U22162 (N_22162,N_21934,N_21759);
nor U22163 (N_22163,N_21881,N_21765);
and U22164 (N_22164,N_21887,N_21790);
nand U22165 (N_22165,N_21823,N_21793);
nor U22166 (N_22166,N_21859,N_21899);
nor U22167 (N_22167,N_21987,N_21960);
or U22168 (N_22168,N_21791,N_21957);
nor U22169 (N_22169,N_21815,N_21882);
xor U22170 (N_22170,N_21859,N_21892);
nand U22171 (N_22171,N_21764,N_21768);
and U22172 (N_22172,N_21881,N_21960);
nand U22173 (N_22173,N_21896,N_21829);
nand U22174 (N_22174,N_21766,N_21995);
and U22175 (N_22175,N_21939,N_21753);
nand U22176 (N_22176,N_21918,N_21866);
xor U22177 (N_22177,N_21783,N_21806);
and U22178 (N_22178,N_21833,N_21760);
nand U22179 (N_22179,N_21985,N_21881);
or U22180 (N_22180,N_21952,N_21823);
nand U22181 (N_22181,N_21894,N_21785);
nor U22182 (N_22182,N_21787,N_21889);
nand U22183 (N_22183,N_21934,N_21939);
xor U22184 (N_22184,N_21969,N_21755);
and U22185 (N_22185,N_21860,N_21939);
nand U22186 (N_22186,N_21888,N_21810);
or U22187 (N_22187,N_21903,N_21764);
or U22188 (N_22188,N_21963,N_21920);
nand U22189 (N_22189,N_21996,N_21769);
xnor U22190 (N_22190,N_21960,N_21797);
nand U22191 (N_22191,N_21944,N_21874);
xnor U22192 (N_22192,N_21851,N_21910);
xnor U22193 (N_22193,N_21885,N_21816);
and U22194 (N_22194,N_21969,N_21882);
nor U22195 (N_22195,N_21916,N_21836);
or U22196 (N_22196,N_21827,N_21968);
nor U22197 (N_22197,N_21964,N_21831);
and U22198 (N_22198,N_21997,N_21978);
xnor U22199 (N_22199,N_21795,N_21796);
or U22200 (N_22200,N_21796,N_21779);
nor U22201 (N_22201,N_21775,N_21929);
nand U22202 (N_22202,N_21834,N_21926);
or U22203 (N_22203,N_21783,N_21926);
or U22204 (N_22204,N_21792,N_21778);
or U22205 (N_22205,N_21954,N_21941);
xnor U22206 (N_22206,N_21765,N_21895);
or U22207 (N_22207,N_21828,N_21999);
nand U22208 (N_22208,N_21975,N_21959);
nor U22209 (N_22209,N_21941,N_21857);
nor U22210 (N_22210,N_21873,N_21790);
xor U22211 (N_22211,N_21786,N_21756);
or U22212 (N_22212,N_21754,N_21839);
or U22213 (N_22213,N_21920,N_21915);
or U22214 (N_22214,N_21831,N_21800);
nor U22215 (N_22215,N_21818,N_21965);
nor U22216 (N_22216,N_21995,N_21900);
nand U22217 (N_22217,N_21756,N_21804);
nor U22218 (N_22218,N_21932,N_21859);
nor U22219 (N_22219,N_21775,N_21840);
or U22220 (N_22220,N_21891,N_21777);
and U22221 (N_22221,N_21842,N_21858);
or U22222 (N_22222,N_21898,N_21993);
nand U22223 (N_22223,N_21908,N_21904);
or U22224 (N_22224,N_21804,N_21831);
nand U22225 (N_22225,N_21910,N_21955);
nor U22226 (N_22226,N_21893,N_21882);
xor U22227 (N_22227,N_21833,N_21920);
nor U22228 (N_22228,N_21780,N_21965);
xnor U22229 (N_22229,N_21806,N_21861);
xnor U22230 (N_22230,N_21869,N_21940);
nor U22231 (N_22231,N_21868,N_21920);
and U22232 (N_22232,N_21771,N_21870);
and U22233 (N_22233,N_21818,N_21846);
and U22234 (N_22234,N_21981,N_21897);
nand U22235 (N_22235,N_21883,N_21920);
nand U22236 (N_22236,N_21785,N_21950);
and U22237 (N_22237,N_21805,N_21947);
and U22238 (N_22238,N_21826,N_21958);
or U22239 (N_22239,N_21919,N_21753);
nor U22240 (N_22240,N_21888,N_21762);
or U22241 (N_22241,N_21902,N_21843);
nor U22242 (N_22242,N_21878,N_21809);
nand U22243 (N_22243,N_21834,N_21837);
and U22244 (N_22244,N_21908,N_21967);
nor U22245 (N_22245,N_21823,N_21850);
or U22246 (N_22246,N_21813,N_21778);
nor U22247 (N_22247,N_21895,N_21902);
and U22248 (N_22248,N_21921,N_21922);
nand U22249 (N_22249,N_21869,N_21849);
nor U22250 (N_22250,N_22165,N_22128);
xor U22251 (N_22251,N_22050,N_22046);
nand U22252 (N_22252,N_22166,N_22077);
nand U22253 (N_22253,N_22090,N_22002);
nand U22254 (N_22254,N_22204,N_22173);
xnor U22255 (N_22255,N_22034,N_22213);
or U22256 (N_22256,N_22247,N_22125);
or U22257 (N_22257,N_22172,N_22178);
xor U22258 (N_22258,N_22001,N_22197);
xnor U22259 (N_22259,N_22071,N_22214);
nand U22260 (N_22260,N_22237,N_22124);
or U22261 (N_22261,N_22037,N_22176);
and U22262 (N_22262,N_22228,N_22210);
and U22263 (N_22263,N_22069,N_22087);
or U22264 (N_22264,N_22147,N_22007);
xor U22265 (N_22265,N_22132,N_22015);
xnor U22266 (N_22266,N_22004,N_22045);
nor U22267 (N_22267,N_22133,N_22168);
nand U22268 (N_22268,N_22026,N_22032);
and U22269 (N_22269,N_22221,N_22096);
nor U22270 (N_22270,N_22070,N_22160);
xnor U22271 (N_22271,N_22218,N_22126);
or U22272 (N_22272,N_22021,N_22079);
and U22273 (N_22273,N_22056,N_22158);
and U22274 (N_22274,N_22140,N_22177);
and U22275 (N_22275,N_22123,N_22036);
nor U22276 (N_22276,N_22058,N_22208);
nor U22277 (N_22277,N_22103,N_22149);
nand U22278 (N_22278,N_22047,N_22244);
xor U22279 (N_22279,N_22187,N_22235);
nor U22280 (N_22280,N_22006,N_22199);
xnor U22281 (N_22281,N_22141,N_22193);
nor U22282 (N_22282,N_22150,N_22089);
and U22283 (N_22283,N_22086,N_22175);
nand U22284 (N_22284,N_22152,N_22039);
nand U22285 (N_22285,N_22061,N_22144);
nor U22286 (N_22286,N_22008,N_22170);
nand U22287 (N_22287,N_22113,N_22022);
and U22288 (N_22288,N_22234,N_22183);
or U22289 (N_22289,N_22188,N_22027);
nor U22290 (N_22290,N_22114,N_22020);
nand U22291 (N_22291,N_22182,N_22143);
or U22292 (N_22292,N_22005,N_22179);
nand U22293 (N_22293,N_22053,N_22206);
and U22294 (N_22294,N_22035,N_22076);
nor U22295 (N_22295,N_22084,N_22192);
nor U22296 (N_22296,N_22003,N_22196);
or U22297 (N_22297,N_22085,N_22131);
and U22298 (N_22298,N_22013,N_22105);
and U22299 (N_22299,N_22029,N_22216);
xor U22300 (N_22300,N_22109,N_22043);
and U22301 (N_22301,N_22014,N_22238);
and U22302 (N_22302,N_22195,N_22054);
xnor U22303 (N_22303,N_22138,N_22059);
xor U22304 (N_22304,N_22151,N_22052);
and U22305 (N_22305,N_22055,N_22010);
or U22306 (N_22306,N_22211,N_22023);
nand U22307 (N_22307,N_22135,N_22049);
nor U22308 (N_22308,N_22137,N_22242);
nor U22309 (N_22309,N_22107,N_22142);
nand U22310 (N_22310,N_22012,N_22134);
and U22311 (N_22311,N_22217,N_22119);
or U22312 (N_22312,N_22220,N_22062);
and U22313 (N_22313,N_22091,N_22122);
nor U22314 (N_22314,N_22060,N_22117);
and U22315 (N_22315,N_22102,N_22030);
or U22316 (N_22316,N_22148,N_22240);
and U22317 (N_22317,N_22121,N_22145);
and U22318 (N_22318,N_22153,N_22190);
and U22319 (N_22319,N_22154,N_22174);
nor U22320 (N_22320,N_22223,N_22156);
xor U22321 (N_22321,N_22248,N_22180);
xnor U22322 (N_22322,N_22212,N_22232);
or U22323 (N_22323,N_22019,N_22202);
and U22324 (N_22324,N_22215,N_22073);
nor U22325 (N_22325,N_22163,N_22233);
nand U22326 (N_22326,N_22207,N_22246);
nor U22327 (N_22327,N_22028,N_22129);
xor U22328 (N_22328,N_22249,N_22189);
xor U22329 (N_22329,N_22000,N_22038);
or U22330 (N_22330,N_22093,N_22205);
nor U22331 (N_22331,N_22241,N_22078);
and U22332 (N_22332,N_22094,N_22009);
nor U22333 (N_22333,N_22081,N_22057);
xor U22334 (N_22334,N_22031,N_22225);
and U22335 (N_22335,N_22167,N_22245);
or U22336 (N_22336,N_22067,N_22229);
xor U22337 (N_22337,N_22191,N_22044);
nand U22338 (N_22338,N_22181,N_22161);
and U22339 (N_22339,N_22231,N_22186);
xor U22340 (N_22340,N_22018,N_22164);
or U22341 (N_22341,N_22100,N_22112);
xnor U22342 (N_22342,N_22230,N_22184);
nor U22343 (N_22343,N_22101,N_22104);
xor U22344 (N_22344,N_22146,N_22169);
nand U22345 (N_22345,N_22194,N_22130);
and U22346 (N_22346,N_22155,N_22108);
nand U22347 (N_22347,N_22092,N_22025);
nand U22348 (N_22348,N_22064,N_22222);
and U22349 (N_22349,N_22097,N_22095);
nor U22350 (N_22350,N_22157,N_22236);
xor U22351 (N_22351,N_22051,N_22041);
and U22352 (N_22352,N_22042,N_22082);
nor U22353 (N_22353,N_22016,N_22219);
and U22354 (N_22354,N_22098,N_22068);
nand U22355 (N_22355,N_22224,N_22162);
or U22356 (N_22356,N_22110,N_22198);
and U22357 (N_22357,N_22106,N_22239);
and U22358 (N_22358,N_22011,N_22111);
xor U22359 (N_22359,N_22118,N_22171);
or U22360 (N_22360,N_22033,N_22116);
xnor U22361 (N_22361,N_22209,N_22024);
and U22362 (N_22362,N_22120,N_22066);
or U22363 (N_22363,N_22099,N_22226);
or U22364 (N_22364,N_22185,N_22203);
or U22365 (N_22365,N_22083,N_22201);
nor U22366 (N_22366,N_22200,N_22074);
xor U22367 (N_22367,N_22063,N_22139);
nor U22368 (N_22368,N_22075,N_22115);
nor U22369 (N_22369,N_22243,N_22136);
nor U22370 (N_22370,N_22088,N_22159);
nand U22371 (N_22371,N_22127,N_22072);
nand U22372 (N_22372,N_22048,N_22227);
and U22373 (N_22373,N_22017,N_22080);
and U22374 (N_22374,N_22040,N_22065);
xor U22375 (N_22375,N_22235,N_22177);
xor U22376 (N_22376,N_22019,N_22137);
nor U22377 (N_22377,N_22236,N_22131);
or U22378 (N_22378,N_22183,N_22117);
nand U22379 (N_22379,N_22013,N_22149);
nand U22380 (N_22380,N_22168,N_22131);
nor U22381 (N_22381,N_22022,N_22228);
nand U22382 (N_22382,N_22227,N_22058);
nor U22383 (N_22383,N_22217,N_22027);
xor U22384 (N_22384,N_22060,N_22088);
and U22385 (N_22385,N_22066,N_22215);
xnor U22386 (N_22386,N_22078,N_22149);
nand U22387 (N_22387,N_22126,N_22022);
and U22388 (N_22388,N_22089,N_22245);
xnor U22389 (N_22389,N_22112,N_22013);
or U22390 (N_22390,N_22126,N_22149);
nand U22391 (N_22391,N_22222,N_22129);
or U22392 (N_22392,N_22046,N_22120);
nand U22393 (N_22393,N_22218,N_22095);
or U22394 (N_22394,N_22099,N_22122);
nor U22395 (N_22395,N_22156,N_22108);
nand U22396 (N_22396,N_22048,N_22234);
and U22397 (N_22397,N_22242,N_22099);
nor U22398 (N_22398,N_22085,N_22061);
nand U22399 (N_22399,N_22132,N_22222);
nor U22400 (N_22400,N_22180,N_22095);
nand U22401 (N_22401,N_22082,N_22039);
nor U22402 (N_22402,N_22143,N_22081);
nor U22403 (N_22403,N_22057,N_22217);
nor U22404 (N_22404,N_22188,N_22170);
nor U22405 (N_22405,N_22191,N_22181);
nand U22406 (N_22406,N_22016,N_22201);
nand U22407 (N_22407,N_22059,N_22224);
or U22408 (N_22408,N_22147,N_22081);
xor U22409 (N_22409,N_22214,N_22166);
or U22410 (N_22410,N_22031,N_22238);
xor U22411 (N_22411,N_22071,N_22215);
or U22412 (N_22412,N_22092,N_22103);
xor U22413 (N_22413,N_22118,N_22109);
nor U22414 (N_22414,N_22059,N_22060);
or U22415 (N_22415,N_22231,N_22090);
and U22416 (N_22416,N_22151,N_22000);
nor U22417 (N_22417,N_22103,N_22001);
and U22418 (N_22418,N_22181,N_22109);
nor U22419 (N_22419,N_22216,N_22021);
xor U22420 (N_22420,N_22193,N_22052);
nand U22421 (N_22421,N_22205,N_22098);
and U22422 (N_22422,N_22199,N_22148);
xnor U22423 (N_22423,N_22165,N_22066);
and U22424 (N_22424,N_22055,N_22016);
or U22425 (N_22425,N_22075,N_22029);
nor U22426 (N_22426,N_22198,N_22191);
nand U22427 (N_22427,N_22173,N_22238);
or U22428 (N_22428,N_22017,N_22203);
nand U22429 (N_22429,N_22199,N_22054);
and U22430 (N_22430,N_22225,N_22132);
or U22431 (N_22431,N_22063,N_22126);
nand U22432 (N_22432,N_22231,N_22059);
xor U22433 (N_22433,N_22216,N_22160);
nand U22434 (N_22434,N_22175,N_22069);
and U22435 (N_22435,N_22159,N_22093);
or U22436 (N_22436,N_22099,N_22165);
or U22437 (N_22437,N_22232,N_22038);
or U22438 (N_22438,N_22012,N_22064);
and U22439 (N_22439,N_22034,N_22249);
xor U22440 (N_22440,N_22033,N_22074);
nor U22441 (N_22441,N_22239,N_22249);
nor U22442 (N_22442,N_22208,N_22017);
or U22443 (N_22443,N_22213,N_22218);
nand U22444 (N_22444,N_22003,N_22115);
and U22445 (N_22445,N_22248,N_22088);
nor U22446 (N_22446,N_22151,N_22248);
nand U22447 (N_22447,N_22080,N_22141);
nand U22448 (N_22448,N_22083,N_22184);
xor U22449 (N_22449,N_22192,N_22191);
xnor U22450 (N_22450,N_22128,N_22177);
and U22451 (N_22451,N_22185,N_22209);
or U22452 (N_22452,N_22078,N_22171);
or U22453 (N_22453,N_22003,N_22136);
nor U22454 (N_22454,N_22046,N_22091);
and U22455 (N_22455,N_22086,N_22246);
nor U22456 (N_22456,N_22247,N_22072);
xnor U22457 (N_22457,N_22190,N_22110);
nand U22458 (N_22458,N_22156,N_22226);
and U22459 (N_22459,N_22146,N_22109);
and U22460 (N_22460,N_22196,N_22117);
and U22461 (N_22461,N_22209,N_22025);
or U22462 (N_22462,N_22196,N_22037);
nand U22463 (N_22463,N_22067,N_22112);
or U22464 (N_22464,N_22048,N_22166);
xnor U22465 (N_22465,N_22115,N_22100);
nand U22466 (N_22466,N_22195,N_22105);
xor U22467 (N_22467,N_22173,N_22116);
and U22468 (N_22468,N_22115,N_22059);
nand U22469 (N_22469,N_22228,N_22061);
and U22470 (N_22470,N_22154,N_22104);
and U22471 (N_22471,N_22005,N_22128);
or U22472 (N_22472,N_22237,N_22014);
and U22473 (N_22473,N_22119,N_22122);
xnor U22474 (N_22474,N_22021,N_22209);
or U22475 (N_22475,N_22149,N_22009);
nand U22476 (N_22476,N_22025,N_22189);
nor U22477 (N_22477,N_22192,N_22046);
nor U22478 (N_22478,N_22080,N_22162);
or U22479 (N_22479,N_22192,N_22028);
or U22480 (N_22480,N_22039,N_22000);
or U22481 (N_22481,N_22135,N_22183);
and U22482 (N_22482,N_22043,N_22080);
nand U22483 (N_22483,N_22109,N_22040);
nand U22484 (N_22484,N_22070,N_22219);
and U22485 (N_22485,N_22203,N_22057);
or U22486 (N_22486,N_22066,N_22108);
and U22487 (N_22487,N_22073,N_22170);
xor U22488 (N_22488,N_22178,N_22113);
nor U22489 (N_22489,N_22047,N_22208);
and U22490 (N_22490,N_22151,N_22032);
nor U22491 (N_22491,N_22172,N_22061);
nor U22492 (N_22492,N_22149,N_22020);
nand U22493 (N_22493,N_22033,N_22169);
or U22494 (N_22494,N_22208,N_22140);
xor U22495 (N_22495,N_22134,N_22032);
or U22496 (N_22496,N_22177,N_22025);
and U22497 (N_22497,N_22069,N_22181);
or U22498 (N_22498,N_22224,N_22211);
or U22499 (N_22499,N_22107,N_22241);
nand U22500 (N_22500,N_22464,N_22311);
nor U22501 (N_22501,N_22498,N_22415);
xor U22502 (N_22502,N_22257,N_22483);
and U22503 (N_22503,N_22380,N_22383);
nand U22504 (N_22504,N_22492,N_22486);
nand U22505 (N_22505,N_22470,N_22473);
and U22506 (N_22506,N_22284,N_22456);
and U22507 (N_22507,N_22396,N_22419);
xnor U22508 (N_22508,N_22333,N_22294);
xor U22509 (N_22509,N_22378,N_22427);
xnor U22510 (N_22510,N_22295,N_22409);
nor U22511 (N_22511,N_22421,N_22286);
and U22512 (N_22512,N_22264,N_22366);
nor U22513 (N_22513,N_22389,N_22491);
nand U22514 (N_22514,N_22263,N_22426);
or U22515 (N_22515,N_22318,N_22394);
and U22516 (N_22516,N_22350,N_22434);
nand U22517 (N_22517,N_22292,N_22254);
or U22518 (N_22518,N_22462,N_22250);
or U22519 (N_22519,N_22407,N_22327);
nor U22520 (N_22520,N_22324,N_22251);
and U22521 (N_22521,N_22382,N_22276);
or U22522 (N_22522,N_22340,N_22277);
nand U22523 (N_22523,N_22479,N_22290);
and U22524 (N_22524,N_22354,N_22410);
nor U22525 (N_22525,N_22321,N_22372);
nor U22526 (N_22526,N_22283,N_22417);
nand U22527 (N_22527,N_22377,N_22465);
nor U22528 (N_22528,N_22402,N_22336);
nor U22529 (N_22529,N_22332,N_22412);
nor U22530 (N_22530,N_22365,N_22315);
and U22531 (N_22531,N_22397,N_22379);
nand U22532 (N_22532,N_22270,N_22446);
xor U22533 (N_22533,N_22369,N_22356);
nor U22534 (N_22534,N_22476,N_22307);
and U22535 (N_22535,N_22301,N_22346);
nor U22536 (N_22536,N_22450,N_22393);
and U22537 (N_22537,N_22285,N_22256);
xnor U22538 (N_22538,N_22337,N_22425);
nor U22539 (N_22539,N_22291,N_22288);
nand U22540 (N_22540,N_22414,N_22430);
nor U22541 (N_22541,N_22310,N_22422);
xnor U22542 (N_22542,N_22439,N_22384);
or U22543 (N_22543,N_22323,N_22469);
xor U22544 (N_22544,N_22253,N_22472);
nor U22545 (N_22545,N_22347,N_22268);
nand U22546 (N_22546,N_22388,N_22448);
or U22547 (N_22547,N_22305,N_22437);
nor U22548 (N_22548,N_22304,N_22339);
xnor U22549 (N_22549,N_22341,N_22271);
and U22550 (N_22550,N_22278,N_22406);
and U22551 (N_22551,N_22424,N_22490);
and U22552 (N_22552,N_22420,N_22474);
and U22553 (N_22553,N_22322,N_22466);
or U22554 (N_22554,N_22451,N_22403);
nand U22555 (N_22555,N_22289,N_22381);
or U22556 (N_22556,N_22261,N_22463);
and U22557 (N_22557,N_22260,N_22471);
and U22558 (N_22558,N_22404,N_22262);
nand U22559 (N_22559,N_22494,N_22440);
nand U22560 (N_22560,N_22478,N_22413);
nor U22561 (N_22561,N_22441,N_22280);
and U22562 (N_22562,N_22468,N_22461);
and U22563 (N_22563,N_22438,N_22416);
and U22564 (N_22564,N_22258,N_22338);
nand U22565 (N_22565,N_22480,N_22391);
nand U22566 (N_22566,N_22309,N_22267);
and U22567 (N_22567,N_22429,N_22458);
xor U22568 (N_22568,N_22488,N_22320);
and U22569 (N_22569,N_22395,N_22489);
nor U22570 (N_22570,N_22445,N_22319);
and U22571 (N_22571,N_22411,N_22298);
and U22572 (N_22572,N_22436,N_22455);
xnor U22573 (N_22573,N_22457,N_22392);
nand U22574 (N_22574,N_22433,N_22368);
and U22575 (N_22575,N_22360,N_22447);
and U22576 (N_22576,N_22475,N_22477);
xnor U22577 (N_22577,N_22266,N_22355);
nor U22578 (N_22578,N_22385,N_22370);
nand U22579 (N_22579,N_22373,N_22444);
nand U22580 (N_22580,N_22431,N_22459);
xor U22581 (N_22581,N_22316,N_22330);
nand U22582 (N_22582,N_22317,N_22481);
xor U22583 (N_22583,N_22374,N_22497);
nor U22584 (N_22584,N_22428,N_22273);
and U22585 (N_22585,N_22496,N_22442);
and U22586 (N_22586,N_22252,N_22255);
xor U22587 (N_22587,N_22265,N_22493);
xnor U22588 (N_22588,N_22281,N_22453);
and U22589 (N_22589,N_22303,N_22400);
and U22590 (N_22590,N_22335,N_22334);
or U22591 (N_22591,N_22423,N_22387);
nor U22592 (N_22592,N_22358,N_22325);
or U22593 (N_22593,N_22357,N_22367);
or U22594 (N_22594,N_22484,N_22326);
or U22595 (N_22595,N_22432,N_22499);
xnor U22596 (N_22596,N_22308,N_22454);
or U22597 (N_22597,N_22482,N_22351);
or U22598 (N_22598,N_22259,N_22269);
nand U22599 (N_22599,N_22343,N_22296);
and U22600 (N_22600,N_22306,N_22460);
nor U22601 (N_22601,N_22279,N_22353);
xnor U22602 (N_22602,N_22274,N_22328);
or U22603 (N_22603,N_22362,N_22345);
xor U22604 (N_22604,N_22299,N_22361);
xnor U22605 (N_22605,N_22399,N_22408);
nand U22606 (N_22606,N_22375,N_22435);
nand U22607 (N_22607,N_22297,N_22287);
or U22608 (N_22608,N_22352,N_22452);
xor U22609 (N_22609,N_22376,N_22331);
nor U22610 (N_22610,N_22342,N_22398);
or U22611 (N_22611,N_22418,N_22293);
xor U22612 (N_22612,N_22344,N_22302);
nand U22613 (N_22613,N_22467,N_22371);
xnor U22614 (N_22614,N_22390,N_22487);
xor U22615 (N_22615,N_22312,N_22329);
nand U22616 (N_22616,N_22313,N_22386);
or U22617 (N_22617,N_22405,N_22349);
and U22618 (N_22618,N_22359,N_22348);
nand U22619 (N_22619,N_22401,N_22272);
or U22620 (N_22620,N_22282,N_22363);
and U22621 (N_22621,N_22443,N_22495);
or U22622 (N_22622,N_22485,N_22275);
xor U22623 (N_22623,N_22449,N_22314);
xnor U22624 (N_22624,N_22300,N_22364);
nand U22625 (N_22625,N_22479,N_22252);
or U22626 (N_22626,N_22316,N_22389);
or U22627 (N_22627,N_22365,N_22473);
or U22628 (N_22628,N_22395,N_22280);
nand U22629 (N_22629,N_22273,N_22434);
nand U22630 (N_22630,N_22449,N_22320);
and U22631 (N_22631,N_22304,N_22257);
xor U22632 (N_22632,N_22329,N_22310);
nand U22633 (N_22633,N_22357,N_22499);
nand U22634 (N_22634,N_22454,N_22424);
nand U22635 (N_22635,N_22311,N_22286);
nor U22636 (N_22636,N_22325,N_22338);
nor U22637 (N_22637,N_22328,N_22288);
xnor U22638 (N_22638,N_22353,N_22298);
nand U22639 (N_22639,N_22339,N_22429);
or U22640 (N_22640,N_22299,N_22442);
or U22641 (N_22641,N_22280,N_22366);
xor U22642 (N_22642,N_22459,N_22283);
or U22643 (N_22643,N_22497,N_22494);
and U22644 (N_22644,N_22495,N_22407);
nand U22645 (N_22645,N_22488,N_22386);
nand U22646 (N_22646,N_22324,N_22340);
nand U22647 (N_22647,N_22491,N_22437);
nor U22648 (N_22648,N_22304,N_22355);
nor U22649 (N_22649,N_22423,N_22309);
nand U22650 (N_22650,N_22470,N_22286);
xor U22651 (N_22651,N_22272,N_22330);
and U22652 (N_22652,N_22442,N_22294);
or U22653 (N_22653,N_22456,N_22423);
nand U22654 (N_22654,N_22259,N_22283);
nor U22655 (N_22655,N_22397,N_22424);
xnor U22656 (N_22656,N_22348,N_22350);
xnor U22657 (N_22657,N_22486,N_22484);
and U22658 (N_22658,N_22375,N_22351);
and U22659 (N_22659,N_22413,N_22353);
nand U22660 (N_22660,N_22283,N_22479);
or U22661 (N_22661,N_22391,N_22389);
xnor U22662 (N_22662,N_22266,N_22402);
nor U22663 (N_22663,N_22407,N_22256);
nor U22664 (N_22664,N_22337,N_22261);
nand U22665 (N_22665,N_22286,N_22312);
or U22666 (N_22666,N_22327,N_22457);
nor U22667 (N_22667,N_22294,N_22295);
nand U22668 (N_22668,N_22424,N_22301);
xor U22669 (N_22669,N_22460,N_22473);
and U22670 (N_22670,N_22292,N_22256);
or U22671 (N_22671,N_22480,N_22448);
or U22672 (N_22672,N_22291,N_22274);
or U22673 (N_22673,N_22284,N_22325);
nor U22674 (N_22674,N_22326,N_22330);
nor U22675 (N_22675,N_22282,N_22354);
and U22676 (N_22676,N_22445,N_22252);
nor U22677 (N_22677,N_22452,N_22267);
xnor U22678 (N_22678,N_22273,N_22304);
nor U22679 (N_22679,N_22331,N_22318);
and U22680 (N_22680,N_22437,N_22271);
nand U22681 (N_22681,N_22382,N_22278);
or U22682 (N_22682,N_22390,N_22456);
and U22683 (N_22683,N_22252,N_22274);
nor U22684 (N_22684,N_22427,N_22312);
nor U22685 (N_22685,N_22487,N_22396);
nor U22686 (N_22686,N_22446,N_22253);
and U22687 (N_22687,N_22443,N_22324);
nand U22688 (N_22688,N_22403,N_22429);
and U22689 (N_22689,N_22409,N_22487);
nand U22690 (N_22690,N_22449,N_22294);
or U22691 (N_22691,N_22283,N_22420);
nor U22692 (N_22692,N_22312,N_22412);
or U22693 (N_22693,N_22259,N_22289);
and U22694 (N_22694,N_22262,N_22382);
and U22695 (N_22695,N_22463,N_22387);
and U22696 (N_22696,N_22459,N_22406);
nor U22697 (N_22697,N_22279,N_22296);
and U22698 (N_22698,N_22313,N_22472);
or U22699 (N_22699,N_22283,N_22425);
xnor U22700 (N_22700,N_22269,N_22258);
nor U22701 (N_22701,N_22332,N_22449);
nor U22702 (N_22702,N_22344,N_22428);
nand U22703 (N_22703,N_22309,N_22269);
nor U22704 (N_22704,N_22445,N_22387);
and U22705 (N_22705,N_22480,N_22460);
nor U22706 (N_22706,N_22420,N_22432);
or U22707 (N_22707,N_22258,N_22476);
nor U22708 (N_22708,N_22452,N_22481);
xor U22709 (N_22709,N_22268,N_22285);
or U22710 (N_22710,N_22327,N_22370);
and U22711 (N_22711,N_22458,N_22342);
nor U22712 (N_22712,N_22306,N_22261);
xnor U22713 (N_22713,N_22460,N_22355);
xor U22714 (N_22714,N_22467,N_22350);
nor U22715 (N_22715,N_22303,N_22410);
and U22716 (N_22716,N_22299,N_22310);
and U22717 (N_22717,N_22261,N_22250);
xor U22718 (N_22718,N_22339,N_22435);
nand U22719 (N_22719,N_22428,N_22380);
or U22720 (N_22720,N_22451,N_22398);
or U22721 (N_22721,N_22361,N_22327);
and U22722 (N_22722,N_22426,N_22399);
xor U22723 (N_22723,N_22441,N_22271);
or U22724 (N_22724,N_22397,N_22422);
and U22725 (N_22725,N_22311,N_22321);
nand U22726 (N_22726,N_22457,N_22499);
nand U22727 (N_22727,N_22422,N_22452);
and U22728 (N_22728,N_22291,N_22323);
nand U22729 (N_22729,N_22381,N_22329);
xnor U22730 (N_22730,N_22294,N_22370);
nor U22731 (N_22731,N_22438,N_22403);
nand U22732 (N_22732,N_22397,N_22314);
nor U22733 (N_22733,N_22278,N_22316);
and U22734 (N_22734,N_22292,N_22318);
or U22735 (N_22735,N_22353,N_22489);
and U22736 (N_22736,N_22272,N_22373);
and U22737 (N_22737,N_22489,N_22392);
xnor U22738 (N_22738,N_22330,N_22453);
or U22739 (N_22739,N_22493,N_22302);
xor U22740 (N_22740,N_22317,N_22364);
nand U22741 (N_22741,N_22386,N_22304);
or U22742 (N_22742,N_22379,N_22257);
nor U22743 (N_22743,N_22488,N_22455);
and U22744 (N_22744,N_22486,N_22395);
and U22745 (N_22745,N_22403,N_22326);
xor U22746 (N_22746,N_22295,N_22423);
or U22747 (N_22747,N_22441,N_22305);
or U22748 (N_22748,N_22410,N_22391);
or U22749 (N_22749,N_22364,N_22427);
or U22750 (N_22750,N_22548,N_22589);
nor U22751 (N_22751,N_22526,N_22665);
nand U22752 (N_22752,N_22585,N_22714);
or U22753 (N_22753,N_22541,N_22501);
xor U22754 (N_22754,N_22690,N_22532);
xor U22755 (N_22755,N_22545,N_22582);
nor U22756 (N_22756,N_22617,N_22540);
nor U22757 (N_22757,N_22591,N_22558);
and U22758 (N_22758,N_22517,N_22745);
nand U22759 (N_22759,N_22514,N_22522);
nor U22760 (N_22760,N_22503,N_22542);
or U22761 (N_22761,N_22638,N_22587);
nor U22762 (N_22762,N_22721,N_22635);
nand U22763 (N_22763,N_22523,N_22544);
or U22764 (N_22764,N_22709,N_22741);
nor U22765 (N_22765,N_22736,N_22533);
nand U22766 (N_22766,N_22670,N_22686);
or U22767 (N_22767,N_22537,N_22563);
nand U22768 (N_22768,N_22551,N_22715);
nand U22769 (N_22769,N_22718,N_22625);
nor U22770 (N_22770,N_22534,N_22643);
xor U22771 (N_22771,N_22560,N_22681);
nor U22772 (N_22772,N_22703,N_22680);
xor U22773 (N_22773,N_22621,N_22504);
nor U22774 (N_22774,N_22570,N_22575);
or U22775 (N_22775,N_22691,N_22521);
and U22776 (N_22776,N_22595,N_22692);
nand U22777 (N_22777,N_22720,N_22586);
or U22778 (N_22778,N_22528,N_22612);
nand U22779 (N_22779,N_22655,N_22530);
nor U22780 (N_22780,N_22505,N_22525);
and U22781 (N_22781,N_22644,N_22737);
and U22782 (N_22782,N_22529,N_22576);
or U22783 (N_22783,N_22704,N_22669);
xor U22784 (N_22784,N_22664,N_22674);
nor U22785 (N_22785,N_22510,N_22749);
nor U22786 (N_22786,N_22557,N_22642);
xnor U22787 (N_22787,N_22512,N_22663);
xnor U22788 (N_22788,N_22717,N_22668);
nor U22789 (N_22789,N_22746,N_22539);
nand U22790 (N_22790,N_22619,N_22614);
nand U22791 (N_22791,N_22622,N_22699);
xnor U22792 (N_22792,N_22659,N_22683);
or U22793 (N_22793,N_22700,N_22698);
nor U22794 (N_22794,N_22590,N_22584);
nor U22795 (N_22795,N_22553,N_22506);
or U22796 (N_22796,N_22599,N_22613);
and U22797 (N_22797,N_22682,N_22733);
nor U22798 (N_22798,N_22743,N_22742);
or U22799 (N_22799,N_22675,N_22687);
xor U22800 (N_22800,N_22711,N_22645);
and U22801 (N_22801,N_22724,N_22607);
xnor U22802 (N_22802,N_22623,N_22535);
nor U22803 (N_22803,N_22660,N_22511);
or U22804 (N_22804,N_22549,N_22654);
nor U22805 (N_22805,N_22605,N_22732);
nor U22806 (N_22806,N_22729,N_22565);
or U22807 (N_22807,N_22731,N_22578);
nor U22808 (N_22808,N_22601,N_22610);
xnor U22809 (N_22809,N_22726,N_22564);
nand U22810 (N_22810,N_22673,N_22705);
nor U22811 (N_22811,N_22609,N_22689);
nor U22812 (N_22812,N_22627,N_22616);
or U22813 (N_22813,N_22649,N_22624);
or U22814 (N_22814,N_22571,N_22566);
xor U22815 (N_22815,N_22581,N_22628);
or U22816 (N_22816,N_22502,N_22516);
or U22817 (N_22817,N_22580,N_22620);
and U22818 (N_22818,N_22588,N_22611);
and U22819 (N_22819,N_22600,N_22583);
nand U22820 (N_22820,N_22694,N_22688);
nor U22821 (N_22821,N_22547,N_22573);
or U22822 (N_22822,N_22738,N_22730);
or U22823 (N_22823,N_22739,N_22536);
and U22824 (N_22824,N_22646,N_22671);
nand U22825 (N_22825,N_22555,N_22693);
nand U22826 (N_22826,N_22615,N_22662);
or U22827 (N_22827,N_22719,N_22507);
or U22828 (N_22828,N_22546,N_22631);
and U22829 (N_22829,N_22722,N_22626);
and U22830 (N_22830,N_22712,N_22740);
or U22831 (N_22831,N_22716,N_22597);
nand U22832 (N_22832,N_22658,N_22672);
xor U22833 (N_22833,N_22592,N_22697);
nand U22834 (N_22834,N_22708,N_22574);
and U22835 (N_22835,N_22667,N_22596);
nand U22836 (N_22836,N_22608,N_22543);
nand U22837 (N_22837,N_22676,N_22677);
nor U22838 (N_22838,N_22579,N_22515);
and U22839 (N_22839,N_22706,N_22652);
nand U22840 (N_22840,N_22509,N_22524);
and U22841 (N_22841,N_22651,N_22657);
nand U22842 (N_22842,N_22701,N_22648);
nand U22843 (N_22843,N_22513,N_22508);
nor U22844 (N_22844,N_22598,N_22561);
and U22845 (N_22845,N_22527,N_22647);
nor U22846 (N_22846,N_22710,N_22538);
nor U22847 (N_22847,N_22639,N_22684);
or U22848 (N_22848,N_22725,N_22678);
or U22849 (N_22849,N_22637,N_22666);
and U22850 (N_22850,N_22661,N_22653);
and U22851 (N_22851,N_22630,N_22735);
nor U22852 (N_22852,N_22695,N_22707);
or U22853 (N_22853,N_22696,N_22594);
or U22854 (N_22854,N_22572,N_22618);
or U22855 (N_22855,N_22569,N_22632);
nor U22856 (N_22856,N_22556,N_22679);
xnor U22857 (N_22857,N_22641,N_22685);
or U22858 (N_22858,N_22640,N_22747);
nand U22859 (N_22859,N_22734,N_22603);
nand U22860 (N_22860,N_22723,N_22744);
nand U22861 (N_22861,N_22500,N_22604);
xnor U22862 (N_22862,N_22713,N_22702);
nor U22863 (N_22863,N_22577,N_22519);
nand U22864 (N_22864,N_22633,N_22636);
nor U22865 (N_22865,N_22520,N_22602);
nor U22866 (N_22866,N_22562,N_22629);
and U22867 (N_22867,N_22727,N_22748);
xor U22868 (N_22868,N_22518,N_22550);
xnor U22869 (N_22869,N_22656,N_22650);
and U22870 (N_22870,N_22634,N_22728);
or U22871 (N_22871,N_22593,N_22552);
xor U22872 (N_22872,N_22554,N_22567);
xor U22873 (N_22873,N_22559,N_22606);
xor U22874 (N_22874,N_22568,N_22531);
nor U22875 (N_22875,N_22635,N_22592);
nor U22876 (N_22876,N_22650,N_22606);
or U22877 (N_22877,N_22570,N_22669);
xor U22878 (N_22878,N_22665,N_22683);
nor U22879 (N_22879,N_22501,N_22696);
and U22880 (N_22880,N_22594,N_22531);
nand U22881 (N_22881,N_22546,N_22677);
nor U22882 (N_22882,N_22630,N_22595);
xor U22883 (N_22883,N_22639,N_22624);
nor U22884 (N_22884,N_22577,N_22624);
or U22885 (N_22885,N_22544,N_22728);
nand U22886 (N_22886,N_22589,N_22530);
and U22887 (N_22887,N_22631,N_22727);
nor U22888 (N_22888,N_22594,N_22557);
and U22889 (N_22889,N_22678,N_22720);
xnor U22890 (N_22890,N_22568,N_22718);
nor U22891 (N_22891,N_22717,N_22657);
xnor U22892 (N_22892,N_22512,N_22598);
or U22893 (N_22893,N_22721,N_22672);
nor U22894 (N_22894,N_22633,N_22605);
or U22895 (N_22895,N_22684,N_22628);
xnor U22896 (N_22896,N_22595,N_22681);
nor U22897 (N_22897,N_22506,N_22708);
nor U22898 (N_22898,N_22500,N_22596);
nor U22899 (N_22899,N_22576,N_22648);
nand U22900 (N_22900,N_22563,N_22724);
xnor U22901 (N_22901,N_22657,N_22556);
nand U22902 (N_22902,N_22715,N_22677);
xor U22903 (N_22903,N_22734,N_22557);
and U22904 (N_22904,N_22686,N_22558);
or U22905 (N_22905,N_22697,N_22516);
and U22906 (N_22906,N_22551,N_22695);
nand U22907 (N_22907,N_22584,N_22621);
xor U22908 (N_22908,N_22707,N_22545);
nand U22909 (N_22909,N_22596,N_22709);
xnor U22910 (N_22910,N_22594,N_22554);
or U22911 (N_22911,N_22509,N_22599);
nand U22912 (N_22912,N_22648,N_22732);
or U22913 (N_22913,N_22687,N_22734);
xnor U22914 (N_22914,N_22540,N_22532);
nand U22915 (N_22915,N_22531,N_22723);
nor U22916 (N_22916,N_22506,N_22586);
nand U22917 (N_22917,N_22640,N_22517);
nor U22918 (N_22918,N_22690,N_22630);
and U22919 (N_22919,N_22686,N_22625);
or U22920 (N_22920,N_22609,N_22650);
or U22921 (N_22921,N_22739,N_22590);
nor U22922 (N_22922,N_22698,N_22599);
nand U22923 (N_22923,N_22598,N_22623);
nand U22924 (N_22924,N_22500,N_22728);
xor U22925 (N_22925,N_22666,N_22653);
or U22926 (N_22926,N_22671,N_22526);
nor U22927 (N_22927,N_22584,N_22518);
nor U22928 (N_22928,N_22746,N_22675);
nand U22929 (N_22929,N_22600,N_22642);
or U22930 (N_22930,N_22633,N_22738);
nor U22931 (N_22931,N_22573,N_22530);
nor U22932 (N_22932,N_22524,N_22717);
xnor U22933 (N_22933,N_22516,N_22614);
and U22934 (N_22934,N_22744,N_22514);
nor U22935 (N_22935,N_22659,N_22532);
nor U22936 (N_22936,N_22720,N_22572);
and U22937 (N_22937,N_22604,N_22677);
nor U22938 (N_22938,N_22681,N_22533);
nand U22939 (N_22939,N_22616,N_22626);
nor U22940 (N_22940,N_22503,N_22553);
and U22941 (N_22941,N_22664,N_22500);
nand U22942 (N_22942,N_22683,N_22523);
nor U22943 (N_22943,N_22721,N_22613);
and U22944 (N_22944,N_22735,N_22552);
xor U22945 (N_22945,N_22556,N_22609);
or U22946 (N_22946,N_22665,N_22658);
xor U22947 (N_22947,N_22527,N_22542);
or U22948 (N_22948,N_22539,N_22717);
xnor U22949 (N_22949,N_22709,N_22723);
nand U22950 (N_22950,N_22739,N_22664);
nand U22951 (N_22951,N_22543,N_22717);
nand U22952 (N_22952,N_22595,N_22521);
xor U22953 (N_22953,N_22569,N_22555);
and U22954 (N_22954,N_22679,N_22637);
nand U22955 (N_22955,N_22655,N_22732);
nor U22956 (N_22956,N_22547,N_22512);
nor U22957 (N_22957,N_22560,N_22702);
and U22958 (N_22958,N_22697,N_22713);
nor U22959 (N_22959,N_22666,N_22722);
nand U22960 (N_22960,N_22522,N_22671);
and U22961 (N_22961,N_22722,N_22674);
or U22962 (N_22962,N_22587,N_22572);
or U22963 (N_22963,N_22619,N_22558);
and U22964 (N_22964,N_22725,N_22528);
xnor U22965 (N_22965,N_22664,N_22671);
nor U22966 (N_22966,N_22669,N_22516);
or U22967 (N_22967,N_22615,N_22638);
nor U22968 (N_22968,N_22663,N_22647);
and U22969 (N_22969,N_22719,N_22675);
or U22970 (N_22970,N_22710,N_22687);
nor U22971 (N_22971,N_22723,N_22638);
xnor U22972 (N_22972,N_22555,N_22559);
xor U22973 (N_22973,N_22666,N_22711);
nand U22974 (N_22974,N_22557,N_22695);
or U22975 (N_22975,N_22517,N_22582);
nor U22976 (N_22976,N_22552,N_22632);
or U22977 (N_22977,N_22549,N_22536);
xnor U22978 (N_22978,N_22706,N_22565);
xor U22979 (N_22979,N_22730,N_22629);
nor U22980 (N_22980,N_22553,N_22739);
xor U22981 (N_22981,N_22567,N_22696);
xnor U22982 (N_22982,N_22600,N_22746);
nor U22983 (N_22983,N_22715,N_22659);
and U22984 (N_22984,N_22704,N_22593);
nand U22985 (N_22985,N_22704,N_22711);
and U22986 (N_22986,N_22599,N_22722);
or U22987 (N_22987,N_22709,N_22584);
xor U22988 (N_22988,N_22706,N_22661);
nand U22989 (N_22989,N_22699,N_22696);
and U22990 (N_22990,N_22748,N_22523);
nor U22991 (N_22991,N_22543,N_22722);
and U22992 (N_22992,N_22626,N_22681);
nand U22993 (N_22993,N_22582,N_22569);
nand U22994 (N_22994,N_22604,N_22705);
nand U22995 (N_22995,N_22598,N_22681);
or U22996 (N_22996,N_22647,N_22683);
or U22997 (N_22997,N_22664,N_22647);
and U22998 (N_22998,N_22677,N_22577);
nand U22999 (N_22999,N_22529,N_22747);
xnor U23000 (N_23000,N_22912,N_22783);
and U23001 (N_23001,N_22774,N_22815);
nand U23002 (N_23002,N_22973,N_22988);
nor U23003 (N_23003,N_22817,N_22952);
or U23004 (N_23004,N_22916,N_22757);
or U23005 (N_23005,N_22970,N_22854);
xnor U23006 (N_23006,N_22870,N_22798);
nor U23007 (N_23007,N_22879,N_22908);
and U23008 (N_23008,N_22990,N_22834);
and U23009 (N_23009,N_22826,N_22764);
or U23010 (N_23010,N_22956,N_22806);
or U23011 (N_23011,N_22779,N_22794);
nand U23012 (N_23012,N_22957,N_22963);
and U23013 (N_23013,N_22781,N_22902);
nand U23014 (N_23014,N_22769,N_22895);
and U23015 (N_23015,N_22775,N_22814);
or U23016 (N_23016,N_22993,N_22937);
and U23017 (N_23017,N_22832,N_22796);
nand U23018 (N_23018,N_22965,N_22843);
nand U23019 (N_23019,N_22761,N_22995);
xnor U23020 (N_23020,N_22984,N_22864);
or U23021 (N_23021,N_22992,N_22987);
or U23022 (N_23022,N_22837,N_22959);
nand U23023 (N_23023,N_22808,N_22771);
and U23024 (N_23024,N_22760,N_22768);
nor U23025 (N_23025,N_22894,N_22942);
and U23026 (N_23026,N_22891,N_22818);
nand U23027 (N_23027,N_22800,N_22866);
or U23028 (N_23028,N_22919,N_22979);
nor U23029 (N_23029,N_22903,N_22960);
nand U23030 (N_23030,N_22869,N_22876);
nor U23031 (N_23031,N_22861,N_22999);
xor U23032 (N_23032,N_22889,N_22933);
or U23033 (N_23033,N_22994,N_22822);
or U23034 (N_23034,N_22780,N_22838);
nand U23035 (N_23035,N_22953,N_22897);
or U23036 (N_23036,N_22788,N_22976);
nor U23037 (N_23037,N_22947,N_22921);
nor U23038 (N_23038,N_22874,N_22886);
and U23039 (N_23039,N_22823,N_22765);
and U23040 (N_23040,N_22844,N_22930);
nand U23041 (N_23041,N_22940,N_22962);
or U23042 (N_23042,N_22905,N_22888);
nand U23043 (N_23043,N_22782,N_22941);
xor U23044 (N_23044,N_22972,N_22885);
xnor U23045 (N_23045,N_22918,N_22829);
nor U23046 (N_23046,N_22898,N_22816);
or U23047 (N_23047,N_22899,N_22954);
or U23048 (N_23048,N_22911,N_22753);
nand U23049 (N_23049,N_22758,N_22901);
nand U23050 (N_23050,N_22880,N_22910);
and U23051 (N_23051,N_22878,N_22938);
xor U23052 (N_23052,N_22945,N_22849);
or U23053 (N_23053,N_22896,N_22801);
nand U23054 (N_23054,N_22795,N_22991);
nor U23055 (N_23055,N_22985,N_22777);
or U23056 (N_23056,N_22871,N_22858);
and U23057 (N_23057,N_22872,N_22950);
nand U23058 (N_23058,N_22873,N_22920);
nor U23059 (N_23059,N_22755,N_22913);
and U23060 (N_23060,N_22907,N_22852);
and U23061 (N_23061,N_22939,N_22935);
xor U23062 (N_23062,N_22958,N_22917);
nand U23063 (N_23063,N_22846,N_22867);
nor U23064 (N_23064,N_22751,N_22949);
nand U23065 (N_23065,N_22791,N_22830);
or U23066 (N_23066,N_22857,N_22778);
nand U23067 (N_23067,N_22936,N_22975);
xnor U23068 (N_23068,N_22803,N_22763);
xnor U23069 (N_23069,N_22804,N_22859);
or U23070 (N_23070,N_22797,N_22847);
nor U23071 (N_23071,N_22883,N_22759);
and U23072 (N_23072,N_22853,N_22807);
xnor U23073 (N_23073,N_22827,N_22835);
nor U23074 (N_23074,N_22934,N_22932);
xnor U23075 (N_23075,N_22851,N_22772);
xor U23076 (N_23076,N_22825,N_22974);
and U23077 (N_23077,N_22929,N_22997);
nand U23078 (N_23078,N_22892,N_22948);
and U23079 (N_23079,N_22931,N_22865);
and U23080 (N_23080,N_22922,N_22978);
nor U23081 (N_23081,N_22875,N_22924);
nor U23082 (N_23082,N_22983,N_22811);
or U23083 (N_23083,N_22840,N_22980);
and U23084 (N_23084,N_22792,N_22845);
nor U23085 (N_23085,N_22951,N_22848);
nor U23086 (N_23086,N_22785,N_22833);
nor U23087 (N_23087,N_22812,N_22943);
or U23088 (N_23088,N_22836,N_22955);
nor U23089 (N_23089,N_22828,N_22906);
xor U23090 (N_23090,N_22961,N_22813);
or U23091 (N_23091,N_22809,N_22754);
nand U23092 (N_23092,N_22868,N_22773);
xor U23093 (N_23093,N_22799,N_22762);
nand U23094 (N_23094,N_22900,N_22810);
or U23095 (N_23095,N_22914,N_22882);
and U23096 (N_23096,N_22776,N_22789);
or U23097 (N_23097,N_22786,N_22770);
and U23098 (N_23098,N_22971,N_22821);
or U23099 (N_23099,N_22968,N_22881);
xnor U23100 (N_23100,N_22909,N_22752);
or U23101 (N_23101,N_22904,N_22927);
nor U23102 (N_23102,N_22856,N_22944);
xnor U23103 (N_23103,N_22824,N_22925);
xor U23104 (N_23104,N_22767,N_22977);
nand U23105 (N_23105,N_22862,N_22989);
nor U23106 (N_23106,N_22887,N_22998);
or U23107 (N_23107,N_22819,N_22831);
and U23108 (N_23108,N_22784,N_22750);
nand U23109 (N_23109,N_22928,N_22839);
or U23110 (N_23110,N_22884,N_22802);
and U23111 (N_23111,N_22842,N_22969);
nand U23112 (N_23112,N_22850,N_22793);
or U23113 (N_23113,N_22926,N_22946);
and U23114 (N_23114,N_22805,N_22996);
and U23115 (N_23115,N_22841,N_22820);
or U23116 (N_23116,N_22982,N_22766);
nor U23117 (N_23117,N_22893,N_22890);
nand U23118 (N_23118,N_22966,N_22915);
nand U23119 (N_23119,N_22967,N_22964);
xor U23120 (N_23120,N_22855,N_22981);
nand U23121 (N_23121,N_22923,N_22877);
nor U23122 (N_23122,N_22986,N_22863);
nor U23123 (N_23123,N_22790,N_22756);
nand U23124 (N_23124,N_22787,N_22860);
and U23125 (N_23125,N_22896,N_22904);
and U23126 (N_23126,N_22976,N_22809);
nor U23127 (N_23127,N_22753,N_22850);
and U23128 (N_23128,N_22830,N_22767);
nor U23129 (N_23129,N_22940,N_22990);
xnor U23130 (N_23130,N_22960,N_22832);
or U23131 (N_23131,N_22942,N_22976);
nor U23132 (N_23132,N_22943,N_22893);
and U23133 (N_23133,N_22963,N_22775);
nand U23134 (N_23134,N_22964,N_22937);
xnor U23135 (N_23135,N_22755,N_22813);
nor U23136 (N_23136,N_22920,N_22802);
nor U23137 (N_23137,N_22874,N_22974);
xnor U23138 (N_23138,N_22769,N_22998);
xnor U23139 (N_23139,N_22796,N_22806);
xor U23140 (N_23140,N_22982,N_22983);
or U23141 (N_23141,N_22827,N_22954);
and U23142 (N_23142,N_22802,N_22753);
nor U23143 (N_23143,N_22786,N_22941);
or U23144 (N_23144,N_22805,N_22773);
xor U23145 (N_23145,N_22813,N_22789);
nor U23146 (N_23146,N_22954,N_22907);
nand U23147 (N_23147,N_22869,N_22922);
nand U23148 (N_23148,N_22909,N_22929);
or U23149 (N_23149,N_22874,N_22779);
xor U23150 (N_23150,N_22916,N_22771);
or U23151 (N_23151,N_22901,N_22821);
nor U23152 (N_23152,N_22802,N_22767);
nand U23153 (N_23153,N_22869,N_22830);
nand U23154 (N_23154,N_22752,N_22860);
xnor U23155 (N_23155,N_22888,N_22825);
or U23156 (N_23156,N_22853,N_22822);
nand U23157 (N_23157,N_22961,N_22947);
nand U23158 (N_23158,N_22964,N_22791);
or U23159 (N_23159,N_22916,N_22908);
xnor U23160 (N_23160,N_22967,N_22948);
nand U23161 (N_23161,N_22858,N_22823);
xnor U23162 (N_23162,N_22952,N_22758);
xor U23163 (N_23163,N_22900,N_22915);
or U23164 (N_23164,N_22933,N_22770);
nor U23165 (N_23165,N_22859,N_22960);
nor U23166 (N_23166,N_22868,N_22899);
nand U23167 (N_23167,N_22833,N_22797);
xor U23168 (N_23168,N_22915,N_22950);
and U23169 (N_23169,N_22902,N_22889);
xnor U23170 (N_23170,N_22769,N_22922);
or U23171 (N_23171,N_22918,N_22864);
nand U23172 (N_23172,N_22844,N_22856);
xor U23173 (N_23173,N_22984,N_22853);
or U23174 (N_23174,N_22926,N_22850);
nor U23175 (N_23175,N_22970,N_22753);
nor U23176 (N_23176,N_22944,N_22838);
nand U23177 (N_23177,N_22808,N_22767);
nor U23178 (N_23178,N_22766,N_22845);
xnor U23179 (N_23179,N_22923,N_22996);
and U23180 (N_23180,N_22804,N_22962);
xor U23181 (N_23181,N_22847,N_22779);
xnor U23182 (N_23182,N_22908,N_22823);
nand U23183 (N_23183,N_22910,N_22938);
nor U23184 (N_23184,N_22942,N_22830);
xor U23185 (N_23185,N_22767,N_22878);
nor U23186 (N_23186,N_22913,N_22812);
nor U23187 (N_23187,N_22824,N_22806);
or U23188 (N_23188,N_22806,N_22817);
or U23189 (N_23189,N_22822,N_22806);
xnor U23190 (N_23190,N_22775,N_22912);
nand U23191 (N_23191,N_22792,N_22892);
and U23192 (N_23192,N_22969,N_22924);
or U23193 (N_23193,N_22752,N_22871);
nand U23194 (N_23194,N_22893,N_22871);
and U23195 (N_23195,N_22856,N_22955);
and U23196 (N_23196,N_22982,N_22756);
or U23197 (N_23197,N_22958,N_22893);
and U23198 (N_23198,N_22754,N_22832);
nand U23199 (N_23199,N_22910,N_22889);
nand U23200 (N_23200,N_22869,N_22935);
or U23201 (N_23201,N_22984,N_22991);
nor U23202 (N_23202,N_22839,N_22788);
nand U23203 (N_23203,N_22829,N_22834);
and U23204 (N_23204,N_22956,N_22824);
nor U23205 (N_23205,N_22907,N_22980);
and U23206 (N_23206,N_22871,N_22784);
nor U23207 (N_23207,N_22872,N_22801);
or U23208 (N_23208,N_22781,N_22750);
xnor U23209 (N_23209,N_22810,N_22987);
and U23210 (N_23210,N_22813,N_22994);
nand U23211 (N_23211,N_22756,N_22875);
and U23212 (N_23212,N_22765,N_22891);
xor U23213 (N_23213,N_22750,N_22842);
and U23214 (N_23214,N_22950,N_22910);
nand U23215 (N_23215,N_22965,N_22767);
or U23216 (N_23216,N_22771,N_22944);
and U23217 (N_23217,N_22809,N_22759);
xnor U23218 (N_23218,N_22920,N_22862);
nor U23219 (N_23219,N_22802,N_22766);
or U23220 (N_23220,N_22858,N_22801);
nand U23221 (N_23221,N_22772,N_22779);
xor U23222 (N_23222,N_22896,N_22892);
xnor U23223 (N_23223,N_22990,N_22781);
xnor U23224 (N_23224,N_22967,N_22957);
nor U23225 (N_23225,N_22909,N_22824);
and U23226 (N_23226,N_22924,N_22980);
nand U23227 (N_23227,N_22795,N_22755);
nand U23228 (N_23228,N_22888,N_22981);
or U23229 (N_23229,N_22797,N_22933);
or U23230 (N_23230,N_22924,N_22818);
nor U23231 (N_23231,N_22875,N_22953);
nand U23232 (N_23232,N_22792,N_22854);
xor U23233 (N_23233,N_22853,N_22933);
or U23234 (N_23234,N_22760,N_22894);
nor U23235 (N_23235,N_22995,N_22937);
or U23236 (N_23236,N_22769,N_22938);
and U23237 (N_23237,N_22924,N_22837);
nand U23238 (N_23238,N_22840,N_22774);
or U23239 (N_23239,N_22998,N_22916);
xnor U23240 (N_23240,N_22979,N_22833);
and U23241 (N_23241,N_22857,N_22773);
nand U23242 (N_23242,N_22899,N_22830);
xor U23243 (N_23243,N_22775,N_22794);
xor U23244 (N_23244,N_22828,N_22915);
nor U23245 (N_23245,N_22788,N_22766);
and U23246 (N_23246,N_22864,N_22806);
nand U23247 (N_23247,N_22750,N_22922);
or U23248 (N_23248,N_22965,N_22892);
nor U23249 (N_23249,N_22770,N_22963);
or U23250 (N_23250,N_23183,N_23010);
or U23251 (N_23251,N_23068,N_23117);
nand U23252 (N_23252,N_23075,N_23085);
nor U23253 (N_23253,N_23009,N_23052);
or U23254 (N_23254,N_23189,N_23166);
nor U23255 (N_23255,N_23160,N_23057);
or U23256 (N_23256,N_23081,N_23011);
and U23257 (N_23257,N_23237,N_23236);
nor U23258 (N_23258,N_23029,N_23061);
or U23259 (N_23259,N_23123,N_23245);
xnor U23260 (N_23260,N_23216,N_23227);
nor U23261 (N_23261,N_23148,N_23008);
xnor U23262 (N_23262,N_23139,N_23230);
xnor U23263 (N_23263,N_23226,N_23122);
nor U23264 (N_23264,N_23003,N_23133);
or U23265 (N_23265,N_23149,N_23062);
nor U23266 (N_23266,N_23113,N_23004);
xor U23267 (N_23267,N_23209,N_23036);
and U23268 (N_23268,N_23221,N_23198);
nand U23269 (N_23269,N_23048,N_23238);
and U23270 (N_23270,N_23042,N_23231);
xor U23271 (N_23271,N_23172,N_23080);
nor U23272 (N_23272,N_23083,N_23091);
or U23273 (N_23273,N_23088,N_23024);
nand U23274 (N_23274,N_23144,N_23035);
nand U23275 (N_23275,N_23059,N_23072);
or U23276 (N_23276,N_23194,N_23214);
or U23277 (N_23277,N_23007,N_23246);
or U23278 (N_23278,N_23224,N_23050);
nand U23279 (N_23279,N_23067,N_23154);
nor U23280 (N_23280,N_23200,N_23031);
nand U23281 (N_23281,N_23065,N_23126);
xor U23282 (N_23282,N_23199,N_23235);
or U23283 (N_23283,N_23056,N_23193);
nor U23284 (N_23284,N_23162,N_23016);
and U23285 (N_23285,N_23114,N_23188);
and U23286 (N_23286,N_23186,N_23131);
nor U23287 (N_23287,N_23096,N_23181);
xnor U23288 (N_23288,N_23101,N_23248);
nor U23289 (N_23289,N_23156,N_23129);
and U23290 (N_23290,N_23225,N_23190);
xor U23291 (N_23291,N_23157,N_23093);
or U23292 (N_23292,N_23141,N_23058);
and U23293 (N_23293,N_23137,N_23147);
and U23294 (N_23294,N_23218,N_23026);
or U23295 (N_23295,N_23241,N_23146);
and U23296 (N_23296,N_23159,N_23006);
or U23297 (N_23297,N_23046,N_23111);
or U23298 (N_23298,N_23039,N_23185);
and U23299 (N_23299,N_23210,N_23105);
xnor U23300 (N_23300,N_23098,N_23204);
xor U23301 (N_23301,N_23213,N_23140);
or U23302 (N_23302,N_23234,N_23182);
nor U23303 (N_23303,N_23138,N_23176);
nand U23304 (N_23304,N_23041,N_23047);
xnor U23305 (N_23305,N_23195,N_23247);
nor U23306 (N_23306,N_23028,N_23175);
nor U23307 (N_23307,N_23171,N_23021);
and U23308 (N_23308,N_23196,N_23032);
nand U23309 (N_23309,N_23066,N_23106);
or U23310 (N_23310,N_23002,N_23121);
or U23311 (N_23311,N_23120,N_23040);
or U23312 (N_23312,N_23125,N_23242);
and U23313 (N_23313,N_23124,N_23037);
or U23314 (N_23314,N_23135,N_23102);
and U23315 (N_23315,N_23012,N_23243);
nor U23316 (N_23316,N_23233,N_23043);
xnor U23317 (N_23317,N_23060,N_23071);
nor U23318 (N_23318,N_23019,N_23220);
and U23319 (N_23319,N_23084,N_23000);
nor U23320 (N_23320,N_23086,N_23119);
or U23321 (N_23321,N_23173,N_23107);
nand U23322 (N_23322,N_23184,N_23094);
nand U23323 (N_23323,N_23078,N_23150);
or U23324 (N_23324,N_23134,N_23142);
nor U23325 (N_23325,N_23178,N_23153);
and U23326 (N_23326,N_23112,N_23151);
and U23327 (N_23327,N_23223,N_23201);
nand U23328 (N_23328,N_23211,N_23217);
xor U23329 (N_23329,N_23179,N_23023);
xor U23330 (N_23330,N_23158,N_23079);
xor U23331 (N_23331,N_23064,N_23099);
xnor U23332 (N_23332,N_23239,N_23167);
nand U23333 (N_23333,N_23013,N_23015);
and U23334 (N_23334,N_23128,N_23203);
or U23335 (N_23335,N_23053,N_23110);
and U23336 (N_23336,N_23087,N_23130);
nand U23337 (N_23337,N_23116,N_23180);
xnor U23338 (N_23338,N_23027,N_23169);
nand U23339 (N_23339,N_23069,N_23082);
and U23340 (N_23340,N_23145,N_23033);
xnor U23341 (N_23341,N_23097,N_23100);
and U23342 (N_23342,N_23034,N_23155);
nand U23343 (N_23343,N_23055,N_23073);
xnor U23344 (N_23344,N_23104,N_23118);
and U23345 (N_23345,N_23174,N_23161);
and U23346 (N_23346,N_23170,N_23074);
nand U23347 (N_23347,N_23207,N_23014);
nor U23348 (N_23348,N_23208,N_23232);
nor U23349 (N_23349,N_23168,N_23109);
xnor U23350 (N_23350,N_23077,N_23020);
and U23351 (N_23351,N_23018,N_23001);
and U23352 (N_23352,N_23244,N_23132);
xnor U23353 (N_23353,N_23022,N_23044);
xor U23354 (N_23354,N_23038,N_23219);
nand U23355 (N_23355,N_23212,N_23249);
and U23356 (N_23356,N_23005,N_23076);
and U23357 (N_23357,N_23192,N_23187);
nand U23358 (N_23358,N_23215,N_23228);
xnor U23359 (N_23359,N_23229,N_23070);
nand U23360 (N_23360,N_23063,N_23089);
or U23361 (N_23361,N_23051,N_23205);
or U23362 (N_23362,N_23152,N_23202);
nand U23363 (N_23363,N_23115,N_23095);
and U23364 (N_23364,N_23049,N_23103);
nand U23365 (N_23365,N_23143,N_23206);
nor U23366 (N_23366,N_23164,N_23045);
nor U23367 (N_23367,N_23127,N_23191);
xor U23368 (N_23368,N_23092,N_23197);
nor U23369 (N_23369,N_23163,N_23017);
xnor U23370 (N_23370,N_23090,N_23222);
and U23371 (N_23371,N_23025,N_23054);
or U23372 (N_23372,N_23030,N_23240);
xor U23373 (N_23373,N_23136,N_23177);
and U23374 (N_23374,N_23108,N_23165);
nor U23375 (N_23375,N_23000,N_23242);
nor U23376 (N_23376,N_23206,N_23068);
or U23377 (N_23377,N_23233,N_23223);
xor U23378 (N_23378,N_23112,N_23023);
and U23379 (N_23379,N_23056,N_23214);
and U23380 (N_23380,N_23026,N_23163);
xor U23381 (N_23381,N_23045,N_23037);
nand U23382 (N_23382,N_23165,N_23081);
and U23383 (N_23383,N_23012,N_23062);
and U23384 (N_23384,N_23205,N_23070);
nor U23385 (N_23385,N_23117,N_23243);
or U23386 (N_23386,N_23081,N_23180);
or U23387 (N_23387,N_23183,N_23116);
xor U23388 (N_23388,N_23130,N_23082);
xor U23389 (N_23389,N_23239,N_23204);
or U23390 (N_23390,N_23201,N_23057);
nand U23391 (N_23391,N_23082,N_23196);
or U23392 (N_23392,N_23061,N_23247);
or U23393 (N_23393,N_23211,N_23231);
and U23394 (N_23394,N_23092,N_23072);
and U23395 (N_23395,N_23206,N_23036);
nand U23396 (N_23396,N_23207,N_23050);
or U23397 (N_23397,N_23037,N_23089);
or U23398 (N_23398,N_23135,N_23022);
nor U23399 (N_23399,N_23043,N_23141);
and U23400 (N_23400,N_23087,N_23145);
nand U23401 (N_23401,N_23131,N_23190);
xnor U23402 (N_23402,N_23084,N_23072);
nor U23403 (N_23403,N_23084,N_23156);
nor U23404 (N_23404,N_23005,N_23218);
or U23405 (N_23405,N_23201,N_23002);
nand U23406 (N_23406,N_23139,N_23222);
nand U23407 (N_23407,N_23043,N_23199);
xnor U23408 (N_23408,N_23171,N_23139);
xnor U23409 (N_23409,N_23214,N_23070);
nor U23410 (N_23410,N_23053,N_23203);
or U23411 (N_23411,N_23119,N_23200);
or U23412 (N_23412,N_23122,N_23224);
xnor U23413 (N_23413,N_23098,N_23150);
nor U23414 (N_23414,N_23050,N_23241);
nor U23415 (N_23415,N_23227,N_23131);
nand U23416 (N_23416,N_23184,N_23041);
xor U23417 (N_23417,N_23202,N_23080);
and U23418 (N_23418,N_23209,N_23145);
or U23419 (N_23419,N_23032,N_23246);
and U23420 (N_23420,N_23181,N_23142);
xor U23421 (N_23421,N_23124,N_23159);
xnor U23422 (N_23422,N_23204,N_23026);
or U23423 (N_23423,N_23023,N_23217);
nand U23424 (N_23424,N_23080,N_23012);
or U23425 (N_23425,N_23072,N_23125);
or U23426 (N_23426,N_23044,N_23127);
xor U23427 (N_23427,N_23088,N_23111);
xnor U23428 (N_23428,N_23069,N_23213);
xor U23429 (N_23429,N_23021,N_23095);
or U23430 (N_23430,N_23051,N_23025);
or U23431 (N_23431,N_23007,N_23076);
or U23432 (N_23432,N_23085,N_23141);
or U23433 (N_23433,N_23068,N_23233);
or U23434 (N_23434,N_23059,N_23092);
xnor U23435 (N_23435,N_23104,N_23205);
nor U23436 (N_23436,N_23045,N_23114);
xnor U23437 (N_23437,N_23092,N_23116);
nor U23438 (N_23438,N_23215,N_23041);
xor U23439 (N_23439,N_23134,N_23031);
and U23440 (N_23440,N_23180,N_23220);
nor U23441 (N_23441,N_23210,N_23151);
nand U23442 (N_23442,N_23172,N_23132);
and U23443 (N_23443,N_23221,N_23173);
nand U23444 (N_23444,N_23207,N_23064);
and U23445 (N_23445,N_23217,N_23075);
nor U23446 (N_23446,N_23118,N_23205);
or U23447 (N_23447,N_23176,N_23128);
xor U23448 (N_23448,N_23085,N_23059);
xor U23449 (N_23449,N_23062,N_23006);
nand U23450 (N_23450,N_23245,N_23051);
nor U23451 (N_23451,N_23119,N_23163);
and U23452 (N_23452,N_23180,N_23233);
xnor U23453 (N_23453,N_23190,N_23054);
and U23454 (N_23454,N_23097,N_23177);
xor U23455 (N_23455,N_23074,N_23025);
nand U23456 (N_23456,N_23116,N_23173);
nor U23457 (N_23457,N_23236,N_23140);
xnor U23458 (N_23458,N_23065,N_23102);
and U23459 (N_23459,N_23038,N_23064);
nand U23460 (N_23460,N_23191,N_23059);
nor U23461 (N_23461,N_23148,N_23209);
and U23462 (N_23462,N_23003,N_23040);
nor U23463 (N_23463,N_23016,N_23051);
nor U23464 (N_23464,N_23068,N_23003);
or U23465 (N_23465,N_23000,N_23024);
nor U23466 (N_23466,N_23215,N_23235);
nand U23467 (N_23467,N_23169,N_23138);
and U23468 (N_23468,N_23074,N_23210);
or U23469 (N_23469,N_23185,N_23155);
xor U23470 (N_23470,N_23136,N_23211);
or U23471 (N_23471,N_23248,N_23199);
xor U23472 (N_23472,N_23161,N_23193);
nor U23473 (N_23473,N_23113,N_23166);
nand U23474 (N_23474,N_23064,N_23139);
nand U23475 (N_23475,N_23015,N_23080);
xor U23476 (N_23476,N_23135,N_23162);
nand U23477 (N_23477,N_23103,N_23063);
and U23478 (N_23478,N_23120,N_23205);
nand U23479 (N_23479,N_23043,N_23082);
nand U23480 (N_23480,N_23011,N_23189);
and U23481 (N_23481,N_23160,N_23102);
or U23482 (N_23482,N_23196,N_23057);
or U23483 (N_23483,N_23242,N_23067);
or U23484 (N_23484,N_23094,N_23229);
or U23485 (N_23485,N_23118,N_23213);
nor U23486 (N_23486,N_23057,N_23063);
nand U23487 (N_23487,N_23111,N_23165);
and U23488 (N_23488,N_23095,N_23038);
xnor U23489 (N_23489,N_23232,N_23198);
or U23490 (N_23490,N_23204,N_23087);
nand U23491 (N_23491,N_23089,N_23194);
and U23492 (N_23492,N_23026,N_23093);
xor U23493 (N_23493,N_23112,N_23058);
nand U23494 (N_23494,N_23189,N_23156);
xnor U23495 (N_23495,N_23171,N_23178);
xnor U23496 (N_23496,N_23178,N_23114);
or U23497 (N_23497,N_23107,N_23065);
nor U23498 (N_23498,N_23164,N_23138);
xnor U23499 (N_23499,N_23060,N_23056);
and U23500 (N_23500,N_23250,N_23397);
nor U23501 (N_23501,N_23329,N_23252);
nand U23502 (N_23502,N_23491,N_23301);
and U23503 (N_23503,N_23404,N_23422);
nand U23504 (N_23504,N_23416,N_23409);
xor U23505 (N_23505,N_23369,N_23350);
nand U23506 (N_23506,N_23298,N_23407);
or U23507 (N_23507,N_23282,N_23293);
or U23508 (N_23508,N_23291,N_23492);
nor U23509 (N_23509,N_23382,N_23365);
or U23510 (N_23510,N_23493,N_23489);
xnor U23511 (N_23511,N_23454,N_23332);
nor U23512 (N_23512,N_23356,N_23432);
nor U23513 (N_23513,N_23488,N_23473);
or U23514 (N_23514,N_23261,N_23352);
nor U23515 (N_23515,N_23391,N_23343);
nand U23516 (N_23516,N_23364,N_23286);
or U23517 (N_23517,N_23274,N_23482);
and U23518 (N_23518,N_23460,N_23277);
or U23519 (N_23519,N_23424,N_23484);
and U23520 (N_23520,N_23344,N_23314);
and U23521 (N_23521,N_23318,N_23411);
or U23522 (N_23522,N_23387,N_23323);
nand U23523 (N_23523,N_23372,N_23430);
nand U23524 (N_23524,N_23358,N_23464);
and U23525 (N_23525,N_23302,N_23283);
nor U23526 (N_23526,N_23434,N_23326);
nor U23527 (N_23527,N_23384,N_23266);
or U23528 (N_23528,N_23295,N_23325);
and U23529 (N_23529,N_23459,N_23486);
and U23530 (N_23530,N_23285,N_23334);
nor U23531 (N_23531,N_23386,N_23374);
xor U23532 (N_23532,N_23353,N_23475);
or U23533 (N_23533,N_23457,N_23273);
and U23534 (N_23534,N_23275,N_23453);
and U23535 (N_23535,N_23461,N_23467);
nor U23536 (N_23536,N_23466,N_23462);
or U23537 (N_23537,N_23417,N_23414);
xor U23538 (N_23538,N_23481,N_23324);
or U23539 (N_23539,N_23485,N_23476);
nor U23540 (N_23540,N_23494,N_23395);
xor U23541 (N_23541,N_23435,N_23477);
nor U23542 (N_23542,N_23465,N_23284);
xnor U23543 (N_23543,N_23471,N_23310);
or U23544 (N_23544,N_23499,N_23342);
or U23545 (N_23545,N_23394,N_23357);
and U23546 (N_23546,N_23483,N_23319);
xnor U23547 (N_23547,N_23498,N_23479);
or U23548 (N_23548,N_23495,N_23315);
nor U23549 (N_23549,N_23260,N_23415);
or U23550 (N_23550,N_23402,N_23289);
xor U23551 (N_23551,N_23253,N_23333);
and U23552 (N_23552,N_23428,N_23442);
nand U23553 (N_23553,N_23383,N_23292);
nand U23554 (N_23554,N_23309,N_23406);
nor U23555 (N_23555,N_23472,N_23456);
xnor U23556 (N_23556,N_23346,N_23355);
nand U23557 (N_23557,N_23392,N_23449);
nor U23558 (N_23558,N_23276,N_23373);
xor U23559 (N_23559,N_23308,N_23251);
nor U23560 (N_23560,N_23311,N_23267);
or U23561 (N_23561,N_23371,N_23367);
xor U23562 (N_23562,N_23307,N_23487);
or U23563 (N_23563,N_23412,N_23450);
xnor U23564 (N_23564,N_23349,N_23431);
or U23565 (N_23565,N_23306,N_23321);
nor U23566 (N_23566,N_23296,N_23354);
xor U23567 (N_23567,N_23294,N_23375);
nor U23568 (N_23568,N_23288,N_23256);
nor U23569 (N_23569,N_23388,N_23497);
nand U23570 (N_23570,N_23351,N_23341);
nand U23571 (N_23571,N_23259,N_23418);
xnor U23572 (N_23572,N_23257,N_23303);
nand U23573 (N_23573,N_23389,N_23437);
or U23574 (N_23574,N_23444,N_23413);
nor U23575 (N_23575,N_23421,N_23265);
and U23576 (N_23576,N_23470,N_23451);
and U23577 (N_23577,N_23279,N_23328);
and U23578 (N_23578,N_23452,N_23370);
nand U23579 (N_23579,N_23270,N_23340);
xor U23580 (N_23580,N_23366,N_23455);
nor U23581 (N_23581,N_23377,N_23446);
nor U23582 (N_23582,N_23320,N_23438);
nor U23583 (N_23583,N_23447,N_23338);
and U23584 (N_23584,N_23269,N_23255);
nor U23585 (N_23585,N_23268,N_23474);
and U23586 (N_23586,N_23339,N_23316);
xor U23587 (N_23587,N_23300,N_23496);
nand U23588 (N_23588,N_23401,N_23399);
or U23589 (N_23589,N_23322,N_23336);
or U23590 (N_23590,N_23290,N_23448);
nor U23591 (N_23591,N_23490,N_23425);
and U23592 (N_23592,N_23480,N_23385);
or U23593 (N_23593,N_23436,N_23376);
and U23594 (N_23594,N_23304,N_23441);
xnor U23595 (N_23595,N_23419,N_23433);
and U23596 (N_23596,N_23458,N_23272);
and U23597 (N_23597,N_23312,N_23263);
xor U23598 (N_23598,N_23400,N_23330);
and U23599 (N_23599,N_23405,N_23396);
or U23600 (N_23600,N_23297,N_23403);
and U23601 (N_23601,N_23381,N_23271);
nand U23602 (N_23602,N_23426,N_23468);
or U23603 (N_23603,N_23313,N_23258);
nand U23604 (N_23604,N_23360,N_23347);
nand U23605 (N_23605,N_23439,N_23345);
and U23606 (N_23606,N_23254,N_23363);
and U23607 (N_23607,N_23393,N_23378);
xor U23608 (N_23608,N_23429,N_23335);
or U23609 (N_23609,N_23359,N_23287);
and U23610 (N_23610,N_23445,N_23410);
xor U23611 (N_23611,N_23362,N_23262);
nand U23612 (N_23612,N_23443,N_23427);
or U23613 (N_23613,N_23299,N_23281);
and U23614 (N_23614,N_23423,N_23390);
nand U23615 (N_23615,N_23348,N_23469);
and U23616 (N_23616,N_23280,N_23398);
or U23617 (N_23617,N_23380,N_23305);
and U23618 (N_23618,N_23264,N_23379);
nor U23619 (N_23619,N_23368,N_23278);
xor U23620 (N_23620,N_23408,N_23463);
xor U23621 (N_23621,N_23317,N_23420);
or U23622 (N_23622,N_23331,N_23327);
or U23623 (N_23623,N_23478,N_23440);
and U23624 (N_23624,N_23337,N_23361);
xnor U23625 (N_23625,N_23456,N_23283);
and U23626 (N_23626,N_23375,N_23367);
and U23627 (N_23627,N_23302,N_23251);
or U23628 (N_23628,N_23409,N_23404);
nor U23629 (N_23629,N_23274,N_23298);
xor U23630 (N_23630,N_23444,N_23346);
or U23631 (N_23631,N_23492,N_23441);
xnor U23632 (N_23632,N_23335,N_23399);
or U23633 (N_23633,N_23404,N_23285);
and U23634 (N_23634,N_23412,N_23319);
and U23635 (N_23635,N_23289,N_23310);
nand U23636 (N_23636,N_23330,N_23278);
and U23637 (N_23637,N_23490,N_23443);
nor U23638 (N_23638,N_23358,N_23422);
and U23639 (N_23639,N_23414,N_23408);
xnor U23640 (N_23640,N_23339,N_23483);
or U23641 (N_23641,N_23436,N_23257);
xor U23642 (N_23642,N_23291,N_23478);
nor U23643 (N_23643,N_23327,N_23367);
nor U23644 (N_23644,N_23458,N_23318);
nand U23645 (N_23645,N_23445,N_23286);
or U23646 (N_23646,N_23494,N_23497);
nand U23647 (N_23647,N_23342,N_23283);
xor U23648 (N_23648,N_23253,N_23434);
and U23649 (N_23649,N_23260,N_23424);
and U23650 (N_23650,N_23456,N_23261);
and U23651 (N_23651,N_23366,N_23305);
xor U23652 (N_23652,N_23251,N_23282);
and U23653 (N_23653,N_23422,N_23406);
and U23654 (N_23654,N_23468,N_23267);
or U23655 (N_23655,N_23448,N_23298);
xnor U23656 (N_23656,N_23498,N_23268);
xnor U23657 (N_23657,N_23294,N_23413);
or U23658 (N_23658,N_23353,N_23450);
or U23659 (N_23659,N_23346,N_23446);
xnor U23660 (N_23660,N_23251,N_23389);
nand U23661 (N_23661,N_23357,N_23416);
xnor U23662 (N_23662,N_23478,N_23427);
xnor U23663 (N_23663,N_23256,N_23299);
nor U23664 (N_23664,N_23378,N_23463);
nor U23665 (N_23665,N_23332,N_23496);
and U23666 (N_23666,N_23261,N_23413);
nor U23667 (N_23667,N_23287,N_23495);
nor U23668 (N_23668,N_23483,N_23445);
xnor U23669 (N_23669,N_23386,N_23396);
xnor U23670 (N_23670,N_23276,N_23479);
or U23671 (N_23671,N_23445,N_23296);
xnor U23672 (N_23672,N_23260,N_23329);
xnor U23673 (N_23673,N_23322,N_23379);
or U23674 (N_23674,N_23471,N_23343);
nand U23675 (N_23675,N_23444,N_23382);
nor U23676 (N_23676,N_23368,N_23250);
xor U23677 (N_23677,N_23430,N_23421);
xnor U23678 (N_23678,N_23345,N_23495);
nand U23679 (N_23679,N_23273,N_23477);
nor U23680 (N_23680,N_23426,N_23347);
nor U23681 (N_23681,N_23457,N_23492);
xnor U23682 (N_23682,N_23372,N_23330);
and U23683 (N_23683,N_23408,N_23354);
or U23684 (N_23684,N_23398,N_23456);
nand U23685 (N_23685,N_23376,N_23480);
xnor U23686 (N_23686,N_23270,N_23309);
or U23687 (N_23687,N_23467,N_23317);
nand U23688 (N_23688,N_23458,N_23345);
nand U23689 (N_23689,N_23282,N_23346);
nor U23690 (N_23690,N_23432,N_23399);
or U23691 (N_23691,N_23307,N_23349);
xnor U23692 (N_23692,N_23492,N_23287);
and U23693 (N_23693,N_23282,N_23382);
or U23694 (N_23694,N_23335,N_23292);
nor U23695 (N_23695,N_23286,N_23401);
xor U23696 (N_23696,N_23461,N_23254);
and U23697 (N_23697,N_23487,N_23252);
nand U23698 (N_23698,N_23486,N_23334);
or U23699 (N_23699,N_23466,N_23491);
and U23700 (N_23700,N_23417,N_23287);
or U23701 (N_23701,N_23288,N_23343);
nor U23702 (N_23702,N_23374,N_23337);
nor U23703 (N_23703,N_23302,N_23370);
xor U23704 (N_23704,N_23444,N_23361);
xor U23705 (N_23705,N_23285,N_23401);
nor U23706 (N_23706,N_23349,N_23277);
nor U23707 (N_23707,N_23273,N_23495);
xor U23708 (N_23708,N_23400,N_23267);
or U23709 (N_23709,N_23486,N_23419);
and U23710 (N_23710,N_23390,N_23394);
nand U23711 (N_23711,N_23439,N_23258);
xor U23712 (N_23712,N_23335,N_23419);
and U23713 (N_23713,N_23379,N_23313);
nor U23714 (N_23714,N_23264,N_23419);
nor U23715 (N_23715,N_23356,N_23353);
xnor U23716 (N_23716,N_23463,N_23288);
nor U23717 (N_23717,N_23489,N_23443);
xor U23718 (N_23718,N_23321,N_23463);
or U23719 (N_23719,N_23481,N_23295);
nor U23720 (N_23720,N_23337,N_23412);
or U23721 (N_23721,N_23301,N_23498);
or U23722 (N_23722,N_23329,N_23287);
and U23723 (N_23723,N_23429,N_23373);
nor U23724 (N_23724,N_23315,N_23251);
nor U23725 (N_23725,N_23436,N_23433);
nor U23726 (N_23726,N_23480,N_23329);
nand U23727 (N_23727,N_23373,N_23489);
nor U23728 (N_23728,N_23464,N_23396);
nor U23729 (N_23729,N_23492,N_23394);
nand U23730 (N_23730,N_23452,N_23358);
or U23731 (N_23731,N_23403,N_23494);
and U23732 (N_23732,N_23316,N_23370);
xnor U23733 (N_23733,N_23403,N_23324);
xor U23734 (N_23734,N_23368,N_23395);
or U23735 (N_23735,N_23331,N_23397);
or U23736 (N_23736,N_23385,N_23331);
and U23737 (N_23737,N_23396,N_23275);
nor U23738 (N_23738,N_23356,N_23404);
xor U23739 (N_23739,N_23347,N_23405);
nor U23740 (N_23740,N_23324,N_23406);
or U23741 (N_23741,N_23341,N_23435);
nand U23742 (N_23742,N_23325,N_23344);
or U23743 (N_23743,N_23420,N_23412);
nor U23744 (N_23744,N_23262,N_23268);
or U23745 (N_23745,N_23274,N_23414);
nor U23746 (N_23746,N_23468,N_23463);
or U23747 (N_23747,N_23463,N_23467);
and U23748 (N_23748,N_23306,N_23477);
and U23749 (N_23749,N_23330,N_23485);
and U23750 (N_23750,N_23637,N_23543);
xor U23751 (N_23751,N_23672,N_23713);
xor U23752 (N_23752,N_23620,N_23722);
and U23753 (N_23753,N_23639,N_23731);
xor U23754 (N_23754,N_23697,N_23734);
and U23755 (N_23755,N_23729,N_23636);
nand U23756 (N_23756,N_23524,N_23580);
and U23757 (N_23757,N_23599,N_23522);
xor U23758 (N_23758,N_23727,N_23571);
and U23759 (N_23759,N_23631,N_23605);
nand U23760 (N_23760,N_23583,N_23572);
nor U23761 (N_23761,N_23525,N_23558);
xnor U23762 (N_23762,N_23628,N_23655);
xor U23763 (N_23763,N_23533,N_23516);
xor U23764 (N_23764,N_23500,N_23621);
nor U23765 (N_23765,N_23632,N_23553);
and U23766 (N_23766,N_23712,N_23579);
or U23767 (N_23767,N_23741,N_23619);
xnor U23768 (N_23768,N_23596,N_23681);
nand U23769 (N_23769,N_23577,N_23548);
nor U23770 (N_23770,N_23567,N_23640);
xor U23771 (N_23771,N_23728,N_23616);
nor U23772 (N_23772,N_23534,N_23531);
nor U23773 (N_23773,N_23562,N_23663);
or U23774 (N_23774,N_23529,N_23746);
nand U23775 (N_23775,N_23647,N_23740);
xor U23776 (N_23776,N_23506,N_23603);
xnor U23777 (N_23777,N_23608,N_23673);
nand U23778 (N_23778,N_23724,N_23634);
and U23779 (N_23779,N_23625,N_23638);
and U23780 (N_23780,N_23610,N_23536);
nor U23781 (N_23781,N_23660,N_23704);
nand U23782 (N_23782,N_23554,N_23749);
and U23783 (N_23783,N_23699,N_23748);
xnor U23784 (N_23784,N_23508,N_23617);
nor U23785 (N_23785,N_23578,N_23645);
and U23786 (N_23786,N_23544,N_23698);
xnor U23787 (N_23787,N_23745,N_23664);
and U23788 (N_23788,N_23670,N_23703);
nand U23789 (N_23789,N_23515,N_23503);
or U23790 (N_23790,N_23582,N_23726);
and U23791 (N_23791,N_23505,N_23595);
nor U23792 (N_23792,N_23733,N_23611);
nor U23793 (N_23793,N_23566,N_23549);
nor U23794 (N_23794,N_23584,N_23623);
xor U23795 (N_23795,N_23714,N_23707);
and U23796 (N_23796,N_23570,N_23642);
nor U23797 (N_23797,N_23666,N_23658);
or U23798 (N_23798,N_23569,N_23512);
and U23799 (N_23799,N_23565,N_23545);
or U23800 (N_23800,N_23564,N_23648);
nand U23801 (N_23801,N_23626,N_23618);
xnor U23802 (N_23802,N_23541,N_23652);
or U23803 (N_23803,N_23735,N_23687);
nor U23804 (N_23804,N_23592,N_23744);
xnor U23805 (N_23805,N_23743,N_23560);
and U23806 (N_23806,N_23513,N_23688);
nor U23807 (N_23807,N_23527,N_23723);
and U23808 (N_23808,N_23604,N_23725);
and U23809 (N_23809,N_23598,N_23700);
nor U23810 (N_23810,N_23683,N_23693);
or U23811 (N_23811,N_23504,N_23574);
xor U23812 (N_23812,N_23588,N_23606);
xor U23813 (N_23813,N_23706,N_23718);
or U23814 (N_23814,N_23613,N_23667);
or U23815 (N_23815,N_23650,N_23563);
nand U23816 (N_23816,N_23550,N_23542);
xnor U23817 (N_23817,N_23641,N_23518);
and U23818 (N_23818,N_23736,N_23556);
nor U23819 (N_23819,N_23682,N_23539);
nor U23820 (N_23820,N_23523,N_23708);
and U23821 (N_23821,N_23679,N_23609);
nor U23822 (N_23822,N_23691,N_23695);
xor U23823 (N_23823,N_23649,N_23624);
nand U23824 (N_23824,N_23643,N_23555);
and U23825 (N_23825,N_23719,N_23677);
nand U23826 (N_23826,N_23546,N_23528);
nand U23827 (N_23827,N_23559,N_23520);
and U23828 (N_23828,N_23674,N_23540);
xor U23829 (N_23829,N_23573,N_23747);
nand U23830 (N_23830,N_23737,N_23690);
and U23831 (N_23831,N_23709,N_23684);
nand U23832 (N_23832,N_23615,N_23517);
nor U23833 (N_23833,N_23702,N_23717);
and U23834 (N_23834,N_23600,N_23591);
and U23835 (N_23835,N_23501,N_23644);
and U23836 (N_23836,N_23535,N_23685);
nor U23837 (N_23837,N_23659,N_23680);
nand U23838 (N_23838,N_23594,N_23711);
nor U23839 (N_23839,N_23590,N_23689);
xor U23840 (N_23840,N_23742,N_23509);
xnor U23841 (N_23841,N_23581,N_23557);
nor U23842 (N_23842,N_23614,N_23710);
or U23843 (N_23843,N_23510,N_23507);
and U23844 (N_23844,N_23519,N_23701);
or U23845 (N_23845,N_23538,N_23576);
nor U23846 (N_23846,N_23502,N_23597);
and U23847 (N_23847,N_23694,N_23732);
xnor U23848 (N_23848,N_23716,N_23568);
xnor U23849 (N_23849,N_23657,N_23721);
nor U23850 (N_23850,N_23738,N_23547);
xor U23851 (N_23851,N_23671,N_23715);
and U23852 (N_23852,N_23653,N_23654);
nand U23853 (N_23853,N_23665,N_23651);
xnor U23854 (N_23854,N_23602,N_23589);
nor U23855 (N_23855,N_23633,N_23530);
and U23856 (N_23856,N_23669,N_23696);
xor U23857 (N_23857,N_23635,N_23686);
nor U23858 (N_23858,N_23739,N_23593);
nand U23859 (N_23859,N_23678,N_23551);
xor U23860 (N_23860,N_23612,N_23526);
or U23861 (N_23861,N_23629,N_23552);
and U23862 (N_23862,N_23675,N_23662);
nand U23863 (N_23863,N_23627,N_23622);
xor U23864 (N_23864,N_23607,N_23587);
or U23865 (N_23865,N_23561,N_23521);
xnor U23866 (N_23866,N_23514,N_23532);
xor U23867 (N_23867,N_23537,N_23575);
or U23868 (N_23868,N_23705,N_23676);
and U23869 (N_23869,N_23730,N_23720);
and U23870 (N_23870,N_23586,N_23601);
or U23871 (N_23871,N_23692,N_23668);
xor U23872 (N_23872,N_23646,N_23585);
nor U23873 (N_23873,N_23661,N_23511);
or U23874 (N_23874,N_23630,N_23656);
nor U23875 (N_23875,N_23686,N_23707);
and U23876 (N_23876,N_23569,N_23728);
or U23877 (N_23877,N_23574,N_23661);
or U23878 (N_23878,N_23678,N_23546);
and U23879 (N_23879,N_23628,N_23718);
nand U23880 (N_23880,N_23565,N_23566);
nor U23881 (N_23881,N_23537,N_23620);
nor U23882 (N_23882,N_23624,N_23667);
and U23883 (N_23883,N_23654,N_23658);
and U23884 (N_23884,N_23624,N_23572);
nand U23885 (N_23885,N_23539,N_23663);
or U23886 (N_23886,N_23616,N_23566);
nor U23887 (N_23887,N_23695,N_23676);
and U23888 (N_23888,N_23530,N_23702);
xor U23889 (N_23889,N_23719,N_23720);
or U23890 (N_23890,N_23555,N_23616);
nand U23891 (N_23891,N_23587,N_23647);
nor U23892 (N_23892,N_23672,N_23571);
and U23893 (N_23893,N_23638,N_23582);
and U23894 (N_23894,N_23572,N_23577);
nor U23895 (N_23895,N_23597,N_23690);
or U23896 (N_23896,N_23608,N_23678);
xnor U23897 (N_23897,N_23689,N_23544);
and U23898 (N_23898,N_23700,N_23607);
or U23899 (N_23899,N_23601,N_23725);
and U23900 (N_23900,N_23739,N_23743);
and U23901 (N_23901,N_23693,N_23568);
nand U23902 (N_23902,N_23533,N_23717);
nor U23903 (N_23903,N_23679,N_23678);
nand U23904 (N_23904,N_23554,N_23718);
and U23905 (N_23905,N_23707,N_23639);
nand U23906 (N_23906,N_23628,N_23644);
and U23907 (N_23907,N_23667,N_23539);
and U23908 (N_23908,N_23662,N_23573);
nand U23909 (N_23909,N_23539,N_23578);
and U23910 (N_23910,N_23625,N_23688);
nor U23911 (N_23911,N_23717,N_23671);
nor U23912 (N_23912,N_23683,N_23557);
or U23913 (N_23913,N_23702,N_23505);
nor U23914 (N_23914,N_23724,N_23514);
and U23915 (N_23915,N_23602,N_23641);
xor U23916 (N_23916,N_23692,N_23624);
nor U23917 (N_23917,N_23697,N_23523);
xor U23918 (N_23918,N_23682,N_23513);
or U23919 (N_23919,N_23658,N_23512);
xnor U23920 (N_23920,N_23625,N_23722);
and U23921 (N_23921,N_23623,N_23664);
nor U23922 (N_23922,N_23728,N_23618);
and U23923 (N_23923,N_23739,N_23577);
and U23924 (N_23924,N_23643,N_23733);
nor U23925 (N_23925,N_23618,N_23622);
or U23926 (N_23926,N_23503,N_23579);
or U23927 (N_23927,N_23540,N_23689);
or U23928 (N_23928,N_23730,N_23616);
nand U23929 (N_23929,N_23721,N_23673);
nand U23930 (N_23930,N_23513,N_23500);
and U23931 (N_23931,N_23509,N_23582);
nor U23932 (N_23932,N_23608,N_23662);
or U23933 (N_23933,N_23529,N_23644);
xor U23934 (N_23934,N_23514,N_23590);
and U23935 (N_23935,N_23739,N_23682);
and U23936 (N_23936,N_23717,N_23744);
xnor U23937 (N_23937,N_23594,N_23608);
xor U23938 (N_23938,N_23715,N_23738);
xor U23939 (N_23939,N_23555,N_23638);
nand U23940 (N_23940,N_23646,N_23580);
and U23941 (N_23941,N_23644,N_23557);
nor U23942 (N_23942,N_23627,N_23560);
or U23943 (N_23943,N_23599,N_23660);
nor U23944 (N_23944,N_23534,N_23624);
nor U23945 (N_23945,N_23589,N_23591);
nand U23946 (N_23946,N_23564,N_23552);
and U23947 (N_23947,N_23613,N_23623);
and U23948 (N_23948,N_23525,N_23621);
and U23949 (N_23949,N_23723,N_23672);
nor U23950 (N_23950,N_23637,N_23545);
nor U23951 (N_23951,N_23566,N_23612);
xor U23952 (N_23952,N_23631,N_23539);
nor U23953 (N_23953,N_23608,N_23574);
or U23954 (N_23954,N_23547,N_23556);
nand U23955 (N_23955,N_23672,N_23648);
xor U23956 (N_23956,N_23665,N_23518);
nand U23957 (N_23957,N_23599,N_23668);
nand U23958 (N_23958,N_23626,N_23741);
xnor U23959 (N_23959,N_23611,N_23567);
or U23960 (N_23960,N_23651,N_23673);
or U23961 (N_23961,N_23681,N_23568);
nand U23962 (N_23962,N_23684,N_23707);
nand U23963 (N_23963,N_23558,N_23700);
and U23964 (N_23964,N_23638,N_23669);
nor U23965 (N_23965,N_23737,N_23623);
nor U23966 (N_23966,N_23638,N_23567);
and U23967 (N_23967,N_23582,N_23581);
nand U23968 (N_23968,N_23596,N_23730);
nand U23969 (N_23969,N_23708,N_23692);
nand U23970 (N_23970,N_23619,N_23736);
nor U23971 (N_23971,N_23564,N_23677);
nor U23972 (N_23972,N_23532,N_23531);
nor U23973 (N_23973,N_23561,N_23746);
xnor U23974 (N_23974,N_23607,N_23500);
nand U23975 (N_23975,N_23531,N_23566);
nand U23976 (N_23976,N_23659,N_23510);
and U23977 (N_23977,N_23688,N_23666);
nor U23978 (N_23978,N_23616,N_23561);
and U23979 (N_23979,N_23543,N_23618);
nand U23980 (N_23980,N_23560,N_23576);
xnor U23981 (N_23981,N_23522,N_23535);
and U23982 (N_23982,N_23604,N_23715);
xor U23983 (N_23983,N_23668,N_23611);
or U23984 (N_23984,N_23725,N_23632);
or U23985 (N_23985,N_23570,N_23682);
xnor U23986 (N_23986,N_23639,N_23596);
xor U23987 (N_23987,N_23681,N_23720);
nor U23988 (N_23988,N_23749,N_23517);
xor U23989 (N_23989,N_23668,N_23682);
xnor U23990 (N_23990,N_23578,N_23739);
and U23991 (N_23991,N_23577,N_23723);
nor U23992 (N_23992,N_23638,N_23563);
and U23993 (N_23993,N_23715,N_23628);
and U23994 (N_23994,N_23517,N_23661);
or U23995 (N_23995,N_23648,N_23724);
nand U23996 (N_23996,N_23571,N_23656);
xnor U23997 (N_23997,N_23633,N_23595);
nor U23998 (N_23998,N_23603,N_23589);
nor U23999 (N_23999,N_23687,N_23710);
or U24000 (N_24000,N_23902,N_23921);
or U24001 (N_24001,N_23847,N_23994);
nand U24002 (N_24002,N_23796,N_23785);
or U24003 (N_24003,N_23923,N_23954);
nor U24004 (N_24004,N_23838,N_23788);
nand U24005 (N_24005,N_23776,N_23861);
nor U24006 (N_24006,N_23967,N_23859);
nand U24007 (N_24007,N_23901,N_23894);
or U24008 (N_24008,N_23879,N_23778);
nor U24009 (N_24009,N_23871,N_23928);
and U24010 (N_24010,N_23961,N_23878);
nand U24011 (N_24011,N_23781,N_23854);
nand U24012 (N_24012,N_23951,N_23987);
or U24013 (N_24013,N_23813,N_23754);
and U24014 (N_24014,N_23822,N_23899);
nand U24015 (N_24015,N_23929,N_23832);
and U24016 (N_24016,N_23874,N_23770);
nor U24017 (N_24017,N_23803,N_23927);
nor U24018 (N_24018,N_23942,N_23938);
xnor U24019 (N_24019,N_23905,N_23933);
nor U24020 (N_24020,N_23876,N_23889);
or U24021 (N_24021,N_23913,N_23774);
or U24022 (N_24022,N_23896,N_23880);
xnor U24023 (N_24023,N_23970,N_23763);
and U24024 (N_24024,N_23910,N_23771);
nor U24025 (N_24025,N_23953,N_23988);
xnor U24026 (N_24026,N_23858,N_23891);
or U24027 (N_24027,N_23780,N_23996);
nand U24028 (N_24028,N_23978,N_23823);
nand U24029 (N_24029,N_23924,N_23941);
and U24030 (N_24030,N_23869,N_23958);
nor U24031 (N_24031,N_23909,N_23947);
xnor U24032 (N_24032,N_23831,N_23758);
or U24033 (N_24033,N_23751,N_23786);
nand U24034 (N_24034,N_23868,N_23794);
xnor U24035 (N_24035,N_23989,N_23912);
xnor U24036 (N_24036,N_23969,N_23790);
or U24037 (N_24037,N_23965,N_23801);
nor U24038 (N_24038,N_23990,N_23952);
and U24039 (N_24039,N_23852,N_23973);
and U24040 (N_24040,N_23853,N_23864);
nand U24041 (N_24041,N_23837,N_23768);
nand U24042 (N_24042,N_23904,N_23963);
xor U24043 (N_24043,N_23971,N_23860);
and U24044 (N_24044,N_23883,N_23885);
and U24045 (N_24045,N_23760,N_23810);
xnor U24046 (N_24046,N_23907,N_23811);
nand U24047 (N_24047,N_23759,N_23882);
nand U24048 (N_24048,N_23946,N_23979);
and U24049 (N_24049,N_23931,N_23993);
and U24050 (N_24050,N_23908,N_23920);
and U24051 (N_24051,N_23805,N_23750);
nand U24052 (N_24052,N_23962,N_23886);
nand U24053 (N_24053,N_23799,N_23765);
and U24054 (N_24054,N_23764,N_23911);
nor U24055 (N_24055,N_23890,N_23866);
xor U24056 (N_24056,N_23752,N_23782);
nor U24057 (N_24057,N_23888,N_23976);
nor U24058 (N_24058,N_23812,N_23795);
or U24059 (N_24059,N_23769,N_23793);
nand U24060 (N_24060,N_23857,N_23809);
and U24061 (N_24061,N_23991,N_23862);
or U24062 (N_24062,N_23992,N_23835);
nor U24063 (N_24063,N_23825,N_23802);
nand U24064 (N_24064,N_23834,N_23893);
nor U24065 (N_24065,N_23843,N_23791);
nand U24066 (N_24066,N_23981,N_23915);
and U24067 (N_24067,N_23856,N_23959);
or U24068 (N_24068,N_23818,N_23887);
nor U24069 (N_24069,N_23950,N_23877);
xnor U24070 (N_24070,N_23944,N_23895);
and U24071 (N_24071,N_23982,N_23819);
nand U24072 (N_24072,N_23966,N_23919);
nor U24073 (N_24073,N_23997,N_23974);
nand U24074 (N_24074,N_23755,N_23836);
or U24075 (N_24075,N_23984,N_23867);
nor U24076 (N_24076,N_23936,N_23817);
xor U24077 (N_24077,N_23772,N_23829);
or U24078 (N_24078,N_23828,N_23872);
or U24079 (N_24079,N_23766,N_23998);
and U24080 (N_24080,N_23848,N_23850);
or U24081 (N_24081,N_23851,N_23964);
xnor U24082 (N_24082,N_23881,N_23922);
nor U24083 (N_24083,N_23884,N_23995);
nand U24084 (N_24084,N_23784,N_23841);
or U24085 (N_24085,N_23846,N_23949);
or U24086 (N_24086,N_23849,N_23808);
nand U24087 (N_24087,N_23925,N_23903);
nand U24088 (N_24088,N_23972,N_23789);
and U24089 (N_24089,N_23945,N_23756);
nor U24090 (N_24090,N_23757,N_23892);
or U24091 (N_24091,N_23804,N_23968);
nand U24092 (N_24092,N_23821,N_23792);
nand U24093 (N_24093,N_23798,N_23870);
or U24094 (N_24094,N_23948,N_23839);
or U24095 (N_24095,N_23827,N_23762);
xnor U24096 (N_24096,N_23773,N_23845);
and U24097 (N_24097,N_23906,N_23975);
nor U24098 (N_24098,N_23999,N_23783);
nand U24099 (N_24099,N_23943,N_23873);
or U24100 (N_24100,N_23806,N_23957);
nand U24101 (N_24101,N_23955,N_23918);
nand U24102 (N_24102,N_23977,N_23914);
nor U24103 (N_24103,N_23986,N_23797);
nand U24104 (N_24104,N_23844,N_23863);
or U24105 (N_24105,N_23800,N_23807);
xnor U24106 (N_24106,N_23917,N_23815);
or U24107 (N_24107,N_23767,N_23830);
or U24108 (N_24108,N_23814,N_23932);
and U24109 (N_24109,N_23934,N_23935);
nand U24110 (N_24110,N_23816,N_23840);
or U24111 (N_24111,N_23960,N_23956);
nand U24112 (N_24112,N_23939,N_23940);
xnor U24113 (N_24113,N_23898,N_23930);
nand U24114 (N_24114,N_23753,N_23842);
and U24115 (N_24115,N_23826,N_23824);
nand U24116 (N_24116,N_23900,N_23865);
nor U24117 (N_24117,N_23937,N_23875);
and U24118 (N_24118,N_23916,N_23897);
or U24119 (N_24119,N_23761,N_23926);
xnor U24120 (N_24120,N_23787,N_23775);
xnor U24121 (N_24121,N_23983,N_23833);
xnor U24122 (N_24122,N_23820,N_23980);
xnor U24123 (N_24123,N_23777,N_23855);
and U24124 (N_24124,N_23985,N_23779);
and U24125 (N_24125,N_23987,N_23907);
xnor U24126 (N_24126,N_23912,N_23901);
nand U24127 (N_24127,N_23928,N_23772);
nand U24128 (N_24128,N_23949,N_23884);
xnor U24129 (N_24129,N_23824,N_23841);
or U24130 (N_24130,N_23855,N_23868);
nand U24131 (N_24131,N_23792,N_23830);
nor U24132 (N_24132,N_23865,N_23834);
nor U24133 (N_24133,N_23968,N_23898);
nand U24134 (N_24134,N_23915,N_23900);
or U24135 (N_24135,N_23871,N_23985);
xor U24136 (N_24136,N_23956,N_23951);
nor U24137 (N_24137,N_23789,N_23946);
nor U24138 (N_24138,N_23995,N_23898);
nor U24139 (N_24139,N_23901,N_23763);
or U24140 (N_24140,N_23752,N_23813);
or U24141 (N_24141,N_23934,N_23966);
xnor U24142 (N_24142,N_23873,N_23894);
or U24143 (N_24143,N_23927,N_23977);
xor U24144 (N_24144,N_23912,N_23945);
xor U24145 (N_24145,N_23898,N_23771);
or U24146 (N_24146,N_23914,N_23927);
nand U24147 (N_24147,N_23811,N_23806);
nor U24148 (N_24148,N_23848,N_23759);
and U24149 (N_24149,N_23863,N_23890);
nor U24150 (N_24150,N_23753,N_23913);
xnor U24151 (N_24151,N_23883,N_23926);
or U24152 (N_24152,N_23999,N_23899);
and U24153 (N_24153,N_23992,N_23917);
or U24154 (N_24154,N_23881,N_23923);
nor U24155 (N_24155,N_23927,N_23930);
and U24156 (N_24156,N_23909,N_23853);
or U24157 (N_24157,N_23753,N_23755);
or U24158 (N_24158,N_23930,N_23806);
or U24159 (N_24159,N_23776,N_23879);
nor U24160 (N_24160,N_23794,N_23791);
or U24161 (N_24161,N_23862,N_23785);
nand U24162 (N_24162,N_23964,N_23882);
nand U24163 (N_24163,N_23920,N_23837);
nand U24164 (N_24164,N_23990,N_23856);
and U24165 (N_24165,N_23756,N_23837);
nand U24166 (N_24166,N_23783,N_23835);
nand U24167 (N_24167,N_23798,N_23834);
nand U24168 (N_24168,N_23859,N_23771);
xnor U24169 (N_24169,N_23816,N_23815);
or U24170 (N_24170,N_23889,N_23893);
nor U24171 (N_24171,N_23811,N_23840);
nor U24172 (N_24172,N_23791,N_23789);
and U24173 (N_24173,N_23977,N_23946);
or U24174 (N_24174,N_23766,N_23848);
and U24175 (N_24175,N_23884,N_23750);
or U24176 (N_24176,N_23975,N_23822);
xor U24177 (N_24177,N_23878,N_23791);
nand U24178 (N_24178,N_23840,N_23799);
or U24179 (N_24179,N_23855,N_23841);
nand U24180 (N_24180,N_23903,N_23819);
nand U24181 (N_24181,N_23902,N_23976);
nand U24182 (N_24182,N_23867,N_23864);
nand U24183 (N_24183,N_23792,N_23890);
xor U24184 (N_24184,N_23968,N_23849);
or U24185 (N_24185,N_23988,N_23848);
and U24186 (N_24186,N_23860,N_23778);
nor U24187 (N_24187,N_23811,N_23942);
and U24188 (N_24188,N_23935,N_23820);
nor U24189 (N_24189,N_23999,N_23889);
nor U24190 (N_24190,N_23882,N_23975);
or U24191 (N_24191,N_23790,N_23979);
and U24192 (N_24192,N_23876,N_23964);
or U24193 (N_24193,N_23887,N_23899);
nand U24194 (N_24194,N_23934,N_23930);
xor U24195 (N_24195,N_23795,N_23978);
xnor U24196 (N_24196,N_23913,N_23755);
or U24197 (N_24197,N_23777,N_23895);
or U24198 (N_24198,N_23805,N_23869);
nor U24199 (N_24199,N_23934,N_23764);
nand U24200 (N_24200,N_23880,N_23953);
xor U24201 (N_24201,N_23854,N_23938);
xnor U24202 (N_24202,N_23922,N_23783);
xor U24203 (N_24203,N_23824,N_23946);
and U24204 (N_24204,N_23986,N_23868);
xnor U24205 (N_24205,N_23765,N_23943);
or U24206 (N_24206,N_23762,N_23958);
nor U24207 (N_24207,N_23804,N_23758);
nand U24208 (N_24208,N_23846,N_23843);
nor U24209 (N_24209,N_23828,N_23896);
nand U24210 (N_24210,N_23991,N_23853);
nor U24211 (N_24211,N_23900,N_23768);
nor U24212 (N_24212,N_23923,N_23755);
nand U24213 (N_24213,N_23955,N_23876);
xnor U24214 (N_24214,N_23765,N_23830);
or U24215 (N_24215,N_23967,N_23908);
nor U24216 (N_24216,N_23971,N_23789);
and U24217 (N_24217,N_23945,N_23758);
or U24218 (N_24218,N_23835,N_23773);
nor U24219 (N_24219,N_23780,N_23853);
or U24220 (N_24220,N_23800,N_23832);
and U24221 (N_24221,N_23773,N_23979);
nand U24222 (N_24222,N_23765,N_23994);
or U24223 (N_24223,N_23947,N_23970);
nor U24224 (N_24224,N_23891,N_23821);
nor U24225 (N_24225,N_23815,N_23949);
and U24226 (N_24226,N_23917,N_23761);
nand U24227 (N_24227,N_23908,N_23882);
nand U24228 (N_24228,N_23871,N_23971);
xor U24229 (N_24229,N_23796,N_23854);
nor U24230 (N_24230,N_23877,N_23901);
and U24231 (N_24231,N_23816,N_23952);
nand U24232 (N_24232,N_23798,N_23904);
nor U24233 (N_24233,N_23870,N_23954);
nand U24234 (N_24234,N_23879,N_23790);
nor U24235 (N_24235,N_23780,N_23794);
nand U24236 (N_24236,N_23806,N_23950);
and U24237 (N_24237,N_23786,N_23998);
or U24238 (N_24238,N_23923,N_23995);
nor U24239 (N_24239,N_23828,N_23941);
nor U24240 (N_24240,N_23871,N_23972);
nand U24241 (N_24241,N_23791,N_23826);
nor U24242 (N_24242,N_23957,N_23918);
xor U24243 (N_24243,N_23866,N_23919);
and U24244 (N_24244,N_23925,N_23877);
xor U24245 (N_24245,N_23843,N_23982);
and U24246 (N_24246,N_23815,N_23925);
or U24247 (N_24247,N_23818,N_23945);
or U24248 (N_24248,N_23905,N_23974);
xnor U24249 (N_24249,N_23999,N_23907);
or U24250 (N_24250,N_24248,N_24247);
or U24251 (N_24251,N_24232,N_24174);
nor U24252 (N_24252,N_24024,N_24236);
nor U24253 (N_24253,N_24159,N_24198);
nand U24254 (N_24254,N_24243,N_24003);
nand U24255 (N_24255,N_24212,N_24222);
nand U24256 (N_24256,N_24218,N_24092);
nand U24257 (N_24257,N_24191,N_24093);
nand U24258 (N_24258,N_24165,N_24001);
nor U24259 (N_24259,N_24000,N_24123);
nand U24260 (N_24260,N_24061,N_24105);
xor U24261 (N_24261,N_24082,N_24115);
nor U24262 (N_24262,N_24068,N_24245);
nand U24263 (N_24263,N_24089,N_24186);
nand U24264 (N_24264,N_24055,N_24112);
nor U24265 (N_24265,N_24106,N_24064);
nand U24266 (N_24266,N_24086,N_24228);
or U24267 (N_24267,N_24080,N_24065);
nand U24268 (N_24268,N_24150,N_24196);
and U24269 (N_24269,N_24201,N_24234);
xor U24270 (N_24270,N_24079,N_24244);
nor U24271 (N_24271,N_24163,N_24107);
and U24272 (N_24272,N_24227,N_24205);
nor U24273 (N_24273,N_24019,N_24135);
or U24274 (N_24274,N_24169,N_24182);
nor U24275 (N_24275,N_24179,N_24039);
and U24276 (N_24276,N_24155,N_24184);
xnor U24277 (N_24277,N_24108,N_24011);
xor U24278 (N_24278,N_24237,N_24113);
nand U24279 (N_24279,N_24208,N_24072);
nand U24280 (N_24280,N_24056,N_24129);
nor U24281 (N_24281,N_24131,N_24091);
nand U24282 (N_24282,N_24118,N_24062);
and U24283 (N_24283,N_24020,N_24181);
and U24284 (N_24284,N_24120,N_24054);
nand U24285 (N_24285,N_24008,N_24073);
and U24286 (N_24286,N_24199,N_24197);
xor U24287 (N_24287,N_24033,N_24002);
nor U24288 (N_24288,N_24211,N_24180);
or U24289 (N_24289,N_24136,N_24214);
or U24290 (N_24290,N_24134,N_24032);
and U24291 (N_24291,N_24206,N_24226);
nor U24292 (N_24292,N_24176,N_24058);
and U24293 (N_24293,N_24042,N_24238);
nand U24294 (N_24294,N_24172,N_24235);
and U24295 (N_24295,N_24048,N_24220);
or U24296 (N_24296,N_24027,N_24192);
nand U24297 (N_24297,N_24034,N_24233);
nor U24298 (N_24298,N_24170,N_24195);
xnor U24299 (N_24299,N_24037,N_24030);
xor U24300 (N_24300,N_24066,N_24126);
or U24301 (N_24301,N_24230,N_24242);
and U24302 (N_24302,N_24188,N_24146);
or U24303 (N_24303,N_24140,N_24095);
or U24304 (N_24304,N_24138,N_24088);
xor U24305 (N_24305,N_24046,N_24043);
or U24306 (N_24306,N_24096,N_24216);
and U24307 (N_24307,N_24189,N_24026);
nand U24308 (N_24308,N_24153,N_24207);
xor U24309 (N_24309,N_24083,N_24156);
nand U24310 (N_24310,N_24204,N_24125);
nor U24311 (N_24311,N_24006,N_24109);
nand U24312 (N_24312,N_24117,N_24012);
and U24313 (N_24313,N_24071,N_24124);
or U24314 (N_24314,N_24009,N_24110);
nor U24315 (N_24315,N_24147,N_24098);
nor U24316 (N_24316,N_24087,N_24029);
or U24317 (N_24317,N_24041,N_24161);
nand U24318 (N_24318,N_24215,N_24239);
nand U24319 (N_24319,N_24219,N_24246);
nor U24320 (N_24320,N_24075,N_24040);
nand U24321 (N_24321,N_24101,N_24178);
or U24322 (N_24322,N_24194,N_24004);
nand U24323 (N_24323,N_24139,N_24240);
and U24324 (N_24324,N_24154,N_24097);
nor U24325 (N_24325,N_24221,N_24052);
xnor U24326 (N_24326,N_24187,N_24078);
nor U24327 (N_24327,N_24016,N_24103);
nor U24328 (N_24328,N_24070,N_24177);
and U24329 (N_24329,N_24144,N_24128);
xor U24330 (N_24330,N_24085,N_24158);
and U24331 (N_24331,N_24059,N_24143);
or U24332 (N_24332,N_24133,N_24148);
and U24333 (N_24333,N_24152,N_24047);
xnor U24334 (N_24334,N_24121,N_24209);
xnor U24335 (N_24335,N_24044,N_24217);
or U24336 (N_24336,N_24005,N_24094);
nand U24337 (N_24337,N_24132,N_24022);
and U24338 (N_24338,N_24060,N_24183);
or U24339 (N_24339,N_24090,N_24137);
and U24340 (N_24340,N_24167,N_24210);
and U24341 (N_24341,N_24151,N_24031);
nand U24342 (N_24342,N_24007,N_24229);
nor U24343 (N_24343,N_24076,N_24074);
or U24344 (N_24344,N_24099,N_24223);
and U24345 (N_24345,N_24077,N_24200);
xor U24346 (N_24346,N_24035,N_24014);
and U24347 (N_24347,N_24053,N_24203);
or U24348 (N_24348,N_24225,N_24119);
xnor U24349 (N_24349,N_24231,N_24185);
nand U24350 (N_24350,N_24067,N_24104);
or U24351 (N_24351,N_24051,N_24175);
xnor U24352 (N_24352,N_24036,N_24122);
and U24353 (N_24353,N_24018,N_24213);
nor U24354 (N_24354,N_24157,N_24013);
nand U24355 (N_24355,N_24130,N_24193);
xor U24356 (N_24356,N_24141,N_24164);
or U24357 (N_24357,N_24049,N_24168);
xnor U24358 (N_24358,N_24241,N_24084);
nor U24359 (N_24359,N_24162,N_24111);
or U24360 (N_24360,N_24149,N_24114);
or U24361 (N_24361,N_24045,N_24160);
or U24362 (N_24362,N_24063,N_24166);
nor U24363 (N_24363,N_24069,N_24017);
or U24364 (N_24364,N_24010,N_24224);
nor U24365 (N_24365,N_24102,N_24038);
nor U24366 (N_24366,N_24100,N_24173);
nor U24367 (N_24367,N_24023,N_24249);
xnor U24368 (N_24368,N_24025,N_24116);
nor U24369 (N_24369,N_24021,N_24171);
and U24370 (N_24370,N_24202,N_24142);
nand U24371 (N_24371,N_24057,N_24190);
nand U24372 (N_24372,N_24127,N_24081);
nor U24373 (N_24373,N_24050,N_24028);
and U24374 (N_24374,N_24015,N_24145);
nand U24375 (N_24375,N_24109,N_24005);
or U24376 (N_24376,N_24148,N_24182);
and U24377 (N_24377,N_24239,N_24101);
and U24378 (N_24378,N_24228,N_24182);
and U24379 (N_24379,N_24061,N_24239);
nor U24380 (N_24380,N_24199,N_24159);
and U24381 (N_24381,N_24239,N_24136);
and U24382 (N_24382,N_24088,N_24054);
nor U24383 (N_24383,N_24192,N_24194);
and U24384 (N_24384,N_24215,N_24011);
and U24385 (N_24385,N_24134,N_24191);
xor U24386 (N_24386,N_24080,N_24091);
xnor U24387 (N_24387,N_24096,N_24107);
and U24388 (N_24388,N_24026,N_24235);
nor U24389 (N_24389,N_24060,N_24146);
xor U24390 (N_24390,N_24133,N_24023);
nor U24391 (N_24391,N_24011,N_24142);
or U24392 (N_24392,N_24191,N_24128);
nor U24393 (N_24393,N_24010,N_24059);
or U24394 (N_24394,N_24185,N_24089);
and U24395 (N_24395,N_24221,N_24100);
and U24396 (N_24396,N_24132,N_24050);
nand U24397 (N_24397,N_24228,N_24125);
xor U24398 (N_24398,N_24177,N_24238);
nand U24399 (N_24399,N_24179,N_24180);
xor U24400 (N_24400,N_24220,N_24231);
xor U24401 (N_24401,N_24082,N_24012);
nand U24402 (N_24402,N_24030,N_24185);
and U24403 (N_24403,N_24024,N_24154);
and U24404 (N_24404,N_24172,N_24072);
and U24405 (N_24405,N_24166,N_24234);
and U24406 (N_24406,N_24026,N_24149);
and U24407 (N_24407,N_24199,N_24144);
nor U24408 (N_24408,N_24170,N_24175);
and U24409 (N_24409,N_24223,N_24071);
nor U24410 (N_24410,N_24168,N_24234);
nor U24411 (N_24411,N_24074,N_24136);
or U24412 (N_24412,N_24232,N_24224);
and U24413 (N_24413,N_24240,N_24159);
or U24414 (N_24414,N_24078,N_24035);
and U24415 (N_24415,N_24194,N_24071);
or U24416 (N_24416,N_24053,N_24111);
nor U24417 (N_24417,N_24152,N_24241);
xnor U24418 (N_24418,N_24057,N_24161);
nand U24419 (N_24419,N_24131,N_24080);
xor U24420 (N_24420,N_24015,N_24129);
xnor U24421 (N_24421,N_24164,N_24068);
xor U24422 (N_24422,N_24109,N_24197);
or U24423 (N_24423,N_24018,N_24205);
nor U24424 (N_24424,N_24119,N_24057);
nand U24425 (N_24425,N_24073,N_24138);
or U24426 (N_24426,N_24041,N_24132);
nor U24427 (N_24427,N_24161,N_24018);
nor U24428 (N_24428,N_24173,N_24144);
and U24429 (N_24429,N_24148,N_24008);
xnor U24430 (N_24430,N_24224,N_24013);
nand U24431 (N_24431,N_24049,N_24201);
or U24432 (N_24432,N_24153,N_24236);
nor U24433 (N_24433,N_24059,N_24156);
nor U24434 (N_24434,N_24065,N_24066);
nand U24435 (N_24435,N_24233,N_24073);
and U24436 (N_24436,N_24035,N_24191);
xor U24437 (N_24437,N_24237,N_24104);
and U24438 (N_24438,N_24139,N_24038);
nand U24439 (N_24439,N_24232,N_24150);
nand U24440 (N_24440,N_24211,N_24095);
and U24441 (N_24441,N_24187,N_24088);
nor U24442 (N_24442,N_24186,N_24225);
or U24443 (N_24443,N_24079,N_24150);
nand U24444 (N_24444,N_24145,N_24159);
nor U24445 (N_24445,N_24154,N_24031);
and U24446 (N_24446,N_24154,N_24242);
nor U24447 (N_24447,N_24240,N_24017);
xnor U24448 (N_24448,N_24232,N_24145);
xnor U24449 (N_24449,N_24077,N_24084);
or U24450 (N_24450,N_24184,N_24182);
and U24451 (N_24451,N_24086,N_24114);
nor U24452 (N_24452,N_24088,N_24020);
nand U24453 (N_24453,N_24009,N_24236);
xnor U24454 (N_24454,N_24210,N_24091);
and U24455 (N_24455,N_24147,N_24163);
xnor U24456 (N_24456,N_24214,N_24040);
nor U24457 (N_24457,N_24042,N_24137);
or U24458 (N_24458,N_24243,N_24074);
xnor U24459 (N_24459,N_24070,N_24011);
xor U24460 (N_24460,N_24003,N_24057);
xor U24461 (N_24461,N_24086,N_24169);
nor U24462 (N_24462,N_24188,N_24139);
and U24463 (N_24463,N_24212,N_24083);
xor U24464 (N_24464,N_24224,N_24186);
xor U24465 (N_24465,N_24244,N_24041);
nor U24466 (N_24466,N_24138,N_24182);
nand U24467 (N_24467,N_24016,N_24035);
nor U24468 (N_24468,N_24192,N_24123);
and U24469 (N_24469,N_24017,N_24248);
or U24470 (N_24470,N_24189,N_24156);
xnor U24471 (N_24471,N_24165,N_24104);
xor U24472 (N_24472,N_24020,N_24005);
nor U24473 (N_24473,N_24176,N_24191);
or U24474 (N_24474,N_24040,N_24037);
nand U24475 (N_24475,N_24069,N_24176);
or U24476 (N_24476,N_24087,N_24108);
or U24477 (N_24477,N_24116,N_24188);
nor U24478 (N_24478,N_24125,N_24156);
or U24479 (N_24479,N_24067,N_24041);
nand U24480 (N_24480,N_24048,N_24214);
nand U24481 (N_24481,N_24231,N_24127);
and U24482 (N_24482,N_24231,N_24014);
nand U24483 (N_24483,N_24035,N_24154);
nor U24484 (N_24484,N_24174,N_24079);
and U24485 (N_24485,N_24005,N_24043);
and U24486 (N_24486,N_24055,N_24177);
nand U24487 (N_24487,N_24182,N_24192);
xor U24488 (N_24488,N_24018,N_24077);
xnor U24489 (N_24489,N_24100,N_24045);
or U24490 (N_24490,N_24105,N_24025);
and U24491 (N_24491,N_24030,N_24015);
or U24492 (N_24492,N_24050,N_24048);
nor U24493 (N_24493,N_24046,N_24198);
nand U24494 (N_24494,N_24017,N_24081);
nor U24495 (N_24495,N_24084,N_24130);
nor U24496 (N_24496,N_24247,N_24153);
and U24497 (N_24497,N_24234,N_24220);
xnor U24498 (N_24498,N_24227,N_24151);
or U24499 (N_24499,N_24056,N_24248);
nor U24500 (N_24500,N_24326,N_24356);
and U24501 (N_24501,N_24488,N_24306);
nor U24502 (N_24502,N_24355,N_24255);
nor U24503 (N_24503,N_24386,N_24440);
nand U24504 (N_24504,N_24343,N_24481);
xnor U24505 (N_24505,N_24412,N_24480);
or U24506 (N_24506,N_24435,N_24381);
nor U24507 (N_24507,N_24459,N_24484);
and U24508 (N_24508,N_24325,N_24417);
xor U24509 (N_24509,N_24348,N_24449);
nand U24510 (N_24510,N_24323,N_24316);
xor U24511 (N_24511,N_24422,N_24437);
and U24512 (N_24512,N_24457,N_24486);
nor U24513 (N_24513,N_24401,N_24446);
or U24514 (N_24514,N_24405,N_24317);
xnor U24515 (N_24515,N_24463,N_24290);
and U24516 (N_24516,N_24278,N_24336);
or U24517 (N_24517,N_24396,N_24363);
nor U24518 (N_24518,N_24431,N_24297);
nor U24519 (N_24519,N_24420,N_24456);
xor U24520 (N_24520,N_24337,N_24478);
xor U24521 (N_24521,N_24320,N_24364);
nor U24522 (N_24522,N_24257,N_24303);
nor U24523 (N_24523,N_24309,N_24485);
nor U24524 (N_24524,N_24347,N_24376);
xnor U24525 (N_24525,N_24362,N_24461);
xor U24526 (N_24526,N_24310,N_24366);
xor U24527 (N_24527,N_24274,N_24395);
nand U24528 (N_24528,N_24380,N_24379);
nor U24529 (N_24529,N_24474,N_24400);
nand U24530 (N_24530,N_24349,N_24258);
or U24531 (N_24531,N_24436,N_24443);
nand U24532 (N_24532,N_24373,N_24361);
nand U24533 (N_24533,N_24406,N_24399);
and U24534 (N_24534,N_24460,N_24477);
nor U24535 (N_24535,N_24334,N_24368);
nor U24536 (N_24536,N_24266,N_24332);
and U24537 (N_24537,N_24352,N_24359);
or U24538 (N_24538,N_24479,N_24445);
nand U24539 (N_24539,N_24353,N_24264);
xnor U24540 (N_24540,N_24282,N_24433);
or U24541 (N_24541,N_24263,N_24495);
nand U24542 (N_24542,N_24447,N_24298);
xnor U24543 (N_24543,N_24410,N_24487);
and U24544 (N_24544,N_24341,N_24421);
nor U24545 (N_24545,N_24434,N_24415);
nand U24546 (N_24546,N_24441,N_24358);
or U24547 (N_24547,N_24398,N_24491);
and U24548 (N_24548,N_24393,N_24322);
or U24549 (N_24549,N_24284,N_24419);
or U24550 (N_24550,N_24252,N_24388);
nand U24551 (N_24551,N_24344,N_24319);
nand U24552 (N_24552,N_24345,N_24453);
nand U24553 (N_24553,N_24360,N_24372);
or U24554 (N_24554,N_24288,N_24413);
xor U24555 (N_24555,N_24296,N_24267);
nand U24556 (N_24556,N_24275,N_24408);
or U24557 (N_24557,N_24466,N_24301);
nand U24558 (N_24558,N_24467,N_24383);
and U24559 (N_24559,N_24307,N_24472);
nand U24560 (N_24560,N_24494,N_24462);
and U24561 (N_24561,N_24283,N_24351);
and U24562 (N_24562,N_24450,N_24304);
nor U24563 (N_24563,N_24286,N_24251);
and U24564 (N_24564,N_24276,N_24370);
xor U24565 (N_24565,N_24483,N_24254);
nand U24566 (N_24566,N_24311,N_24490);
nor U24567 (N_24567,N_24272,N_24496);
xor U24568 (N_24568,N_24369,N_24279);
xnor U24569 (N_24569,N_24354,N_24497);
or U24570 (N_24570,N_24375,N_24492);
xnor U24571 (N_24571,N_24365,N_24295);
nor U24572 (N_24572,N_24302,N_24292);
and U24573 (N_24573,N_24385,N_24259);
xor U24574 (N_24574,N_24493,N_24262);
or U24575 (N_24575,N_24414,N_24423);
xor U24576 (N_24576,N_24430,N_24285);
nor U24577 (N_24577,N_24260,N_24394);
nand U24578 (N_24578,N_24464,N_24338);
and U24579 (N_24579,N_24328,N_24287);
xor U24580 (N_24580,N_24291,N_24397);
nand U24581 (N_24581,N_24499,N_24498);
or U24582 (N_24582,N_24468,N_24470);
nand U24583 (N_24583,N_24293,N_24416);
or U24584 (N_24584,N_24432,N_24411);
xor U24585 (N_24585,N_24313,N_24407);
nand U24586 (N_24586,N_24321,N_24329);
nor U24587 (N_24587,N_24357,N_24439);
xor U24588 (N_24588,N_24340,N_24438);
or U24589 (N_24589,N_24327,N_24444);
nand U24590 (N_24590,N_24427,N_24346);
nor U24591 (N_24591,N_24305,N_24335);
nand U24592 (N_24592,N_24403,N_24271);
or U24593 (N_24593,N_24425,N_24330);
nand U24594 (N_24594,N_24473,N_24308);
or U24595 (N_24595,N_24424,N_24418);
nand U24596 (N_24596,N_24268,N_24280);
or U24597 (N_24597,N_24350,N_24384);
xor U24598 (N_24598,N_24442,N_24489);
nand U24599 (N_24599,N_24402,N_24390);
nor U24600 (N_24600,N_24318,N_24333);
or U24601 (N_24601,N_24451,N_24458);
nor U24602 (N_24602,N_24324,N_24331);
or U24603 (N_24603,N_24250,N_24367);
nor U24604 (N_24604,N_24371,N_24312);
xnor U24605 (N_24605,N_24315,N_24314);
and U24606 (N_24606,N_24476,N_24392);
and U24607 (N_24607,N_24339,N_24265);
and U24608 (N_24608,N_24382,N_24387);
and U24609 (N_24609,N_24269,N_24299);
or U24610 (N_24610,N_24391,N_24452);
nor U24611 (N_24611,N_24389,N_24253);
or U24612 (N_24612,N_24273,N_24374);
nand U24613 (N_24613,N_24454,N_24455);
nor U24614 (N_24614,N_24469,N_24482);
or U24615 (N_24615,N_24289,N_24429);
nand U24616 (N_24616,N_24378,N_24404);
nand U24617 (N_24617,N_24294,N_24281);
nor U24618 (N_24618,N_24342,N_24465);
nand U24619 (N_24619,N_24277,N_24448);
nand U24620 (N_24620,N_24270,N_24428);
xor U24621 (N_24621,N_24377,N_24300);
xnor U24622 (N_24622,N_24471,N_24256);
nand U24623 (N_24623,N_24261,N_24409);
or U24624 (N_24624,N_24426,N_24475);
and U24625 (N_24625,N_24306,N_24301);
or U24626 (N_24626,N_24471,N_24384);
or U24627 (N_24627,N_24329,N_24400);
and U24628 (N_24628,N_24453,N_24441);
nor U24629 (N_24629,N_24259,N_24368);
nor U24630 (N_24630,N_24269,N_24356);
and U24631 (N_24631,N_24406,N_24384);
or U24632 (N_24632,N_24320,N_24335);
nand U24633 (N_24633,N_24493,N_24328);
and U24634 (N_24634,N_24251,N_24442);
xnor U24635 (N_24635,N_24284,N_24267);
xnor U24636 (N_24636,N_24450,N_24387);
xor U24637 (N_24637,N_24444,N_24322);
or U24638 (N_24638,N_24351,N_24486);
or U24639 (N_24639,N_24353,N_24352);
or U24640 (N_24640,N_24299,N_24289);
and U24641 (N_24641,N_24279,N_24309);
xnor U24642 (N_24642,N_24280,N_24352);
and U24643 (N_24643,N_24281,N_24493);
nand U24644 (N_24644,N_24342,N_24482);
and U24645 (N_24645,N_24359,N_24252);
and U24646 (N_24646,N_24365,N_24480);
nand U24647 (N_24647,N_24487,N_24450);
xor U24648 (N_24648,N_24394,N_24289);
nand U24649 (N_24649,N_24427,N_24358);
or U24650 (N_24650,N_24345,N_24436);
nor U24651 (N_24651,N_24306,N_24426);
nor U24652 (N_24652,N_24273,N_24479);
xnor U24653 (N_24653,N_24458,N_24462);
and U24654 (N_24654,N_24270,N_24310);
nand U24655 (N_24655,N_24396,N_24452);
xor U24656 (N_24656,N_24443,N_24434);
and U24657 (N_24657,N_24251,N_24297);
nor U24658 (N_24658,N_24306,N_24257);
or U24659 (N_24659,N_24373,N_24250);
xor U24660 (N_24660,N_24311,N_24283);
nor U24661 (N_24661,N_24277,N_24488);
nor U24662 (N_24662,N_24254,N_24314);
xor U24663 (N_24663,N_24435,N_24420);
or U24664 (N_24664,N_24406,N_24389);
and U24665 (N_24665,N_24384,N_24382);
nor U24666 (N_24666,N_24276,N_24315);
or U24667 (N_24667,N_24498,N_24395);
nand U24668 (N_24668,N_24431,N_24430);
xnor U24669 (N_24669,N_24453,N_24405);
nand U24670 (N_24670,N_24312,N_24285);
xnor U24671 (N_24671,N_24295,N_24423);
xor U24672 (N_24672,N_24454,N_24400);
xor U24673 (N_24673,N_24384,N_24392);
nor U24674 (N_24674,N_24446,N_24351);
or U24675 (N_24675,N_24474,N_24260);
nand U24676 (N_24676,N_24489,N_24311);
and U24677 (N_24677,N_24382,N_24266);
xnor U24678 (N_24678,N_24375,N_24261);
nor U24679 (N_24679,N_24425,N_24383);
or U24680 (N_24680,N_24251,N_24407);
nor U24681 (N_24681,N_24492,N_24359);
nor U24682 (N_24682,N_24390,N_24287);
nor U24683 (N_24683,N_24338,N_24333);
and U24684 (N_24684,N_24445,N_24376);
xnor U24685 (N_24685,N_24401,N_24445);
nand U24686 (N_24686,N_24454,N_24287);
xor U24687 (N_24687,N_24496,N_24395);
or U24688 (N_24688,N_24257,N_24358);
xor U24689 (N_24689,N_24296,N_24359);
or U24690 (N_24690,N_24312,N_24313);
or U24691 (N_24691,N_24489,N_24470);
xor U24692 (N_24692,N_24400,N_24331);
nand U24693 (N_24693,N_24352,N_24372);
and U24694 (N_24694,N_24431,N_24370);
nor U24695 (N_24695,N_24498,N_24260);
and U24696 (N_24696,N_24266,N_24341);
and U24697 (N_24697,N_24474,N_24351);
xnor U24698 (N_24698,N_24434,N_24370);
or U24699 (N_24699,N_24425,N_24453);
and U24700 (N_24700,N_24325,N_24342);
xnor U24701 (N_24701,N_24499,N_24448);
nand U24702 (N_24702,N_24343,N_24312);
nor U24703 (N_24703,N_24343,N_24369);
or U24704 (N_24704,N_24349,N_24408);
nand U24705 (N_24705,N_24289,N_24449);
or U24706 (N_24706,N_24468,N_24260);
nand U24707 (N_24707,N_24461,N_24274);
or U24708 (N_24708,N_24368,N_24486);
xnor U24709 (N_24709,N_24480,N_24377);
nand U24710 (N_24710,N_24420,N_24309);
xnor U24711 (N_24711,N_24409,N_24392);
xnor U24712 (N_24712,N_24326,N_24370);
or U24713 (N_24713,N_24480,N_24473);
or U24714 (N_24714,N_24376,N_24267);
nand U24715 (N_24715,N_24355,N_24413);
nand U24716 (N_24716,N_24392,N_24429);
nand U24717 (N_24717,N_24404,N_24372);
nor U24718 (N_24718,N_24406,N_24449);
and U24719 (N_24719,N_24455,N_24344);
or U24720 (N_24720,N_24451,N_24479);
and U24721 (N_24721,N_24452,N_24309);
nand U24722 (N_24722,N_24441,N_24381);
nor U24723 (N_24723,N_24262,N_24496);
nand U24724 (N_24724,N_24365,N_24418);
and U24725 (N_24725,N_24300,N_24316);
or U24726 (N_24726,N_24382,N_24464);
xnor U24727 (N_24727,N_24405,N_24286);
nor U24728 (N_24728,N_24454,N_24263);
and U24729 (N_24729,N_24472,N_24372);
nor U24730 (N_24730,N_24499,N_24474);
xor U24731 (N_24731,N_24451,N_24497);
or U24732 (N_24732,N_24255,N_24437);
and U24733 (N_24733,N_24426,N_24388);
nor U24734 (N_24734,N_24394,N_24301);
nor U24735 (N_24735,N_24368,N_24272);
nand U24736 (N_24736,N_24431,N_24339);
xnor U24737 (N_24737,N_24287,N_24312);
nor U24738 (N_24738,N_24404,N_24325);
nor U24739 (N_24739,N_24346,N_24330);
or U24740 (N_24740,N_24446,N_24470);
or U24741 (N_24741,N_24392,N_24438);
or U24742 (N_24742,N_24414,N_24301);
and U24743 (N_24743,N_24413,N_24292);
nor U24744 (N_24744,N_24474,N_24297);
and U24745 (N_24745,N_24326,N_24271);
nand U24746 (N_24746,N_24329,N_24308);
nand U24747 (N_24747,N_24315,N_24338);
or U24748 (N_24748,N_24264,N_24385);
nor U24749 (N_24749,N_24464,N_24274);
or U24750 (N_24750,N_24501,N_24599);
or U24751 (N_24751,N_24631,N_24544);
xor U24752 (N_24752,N_24612,N_24585);
nor U24753 (N_24753,N_24548,N_24524);
or U24754 (N_24754,N_24639,N_24511);
nor U24755 (N_24755,N_24626,N_24689);
nor U24756 (N_24756,N_24651,N_24623);
and U24757 (N_24757,N_24742,N_24546);
and U24758 (N_24758,N_24620,N_24654);
xnor U24759 (N_24759,N_24641,N_24520);
xnor U24760 (N_24760,N_24568,N_24660);
nor U24761 (N_24761,N_24642,N_24703);
nand U24762 (N_24762,N_24658,N_24622);
nor U24763 (N_24763,N_24556,N_24722);
and U24764 (N_24764,N_24694,N_24743);
xnor U24765 (N_24765,N_24578,N_24704);
nor U24766 (N_24766,N_24664,N_24738);
xnor U24767 (N_24767,N_24611,N_24618);
xnor U24768 (N_24768,N_24507,N_24676);
nand U24769 (N_24769,N_24557,N_24636);
nor U24770 (N_24770,N_24593,N_24597);
and U24771 (N_24771,N_24627,N_24613);
nor U24772 (N_24772,N_24691,N_24734);
xor U24773 (N_24773,N_24523,N_24635);
or U24774 (N_24774,N_24619,N_24659);
nand U24775 (N_24775,N_24579,N_24615);
or U24776 (N_24776,N_24736,N_24560);
nand U24777 (N_24777,N_24514,N_24528);
xor U24778 (N_24778,N_24649,N_24540);
xnor U24779 (N_24779,N_24569,N_24707);
nand U24780 (N_24780,N_24705,N_24666);
or U24781 (N_24781,N_24632,N_24522);
and U24782 (N_24782,N_24679,N_24698);
or U24783 (N_24783,N_24706,N_24504);
xnor U24784 (N_24784,N_24720,N_24576);
nand U24785 (N_24785,N_24749,N_24564);
nor U24786 (N_24786,N_24602,N_24638);
xnor U24787 (N_24787,N_24739,N_24737);
and U24788 (N_24788,N_24532,N_24603);
and U24789 (N_24789,N_24616,N_24625);
nand U24790 (N_24790,N_24633,N_24509);
or U24791 (N_24791,N_24656,N_24589);
nand U24792 (N_24792,N_24673,N_24601);
and U24793 (N_24793,N_24541,N_24617);
xnor U24794 (N_24794,N_24688,N_24590);
and U24795 (N_24795,N_24567,N_24515);
xor U24796 (N_24796,N_24566,N_24655);
and U24797 (N_24797,N_24693,N_24628);
nor U24798 (N_24798,N_24549,N_24561);
xnor U24799 (N_24799,N_24735,N_24592);
and U24800 (N_24800,N_24558,N_24591);
and U24801 (N_24801,N_24637,N_24526);
nor U24802 (N_24802,N_24701,N_24500);
xor U24803 (N_24803,N_24510,N_24685);
and U24804 (N_24804,N_24624,N_24634);
xnor U24805 (N_24805,N_24729,N_24723);
nand U24806 (N_24806,N_24724,N_24586);
nand U24807 (N_24807,N_24594,N_24537);
nor U24808 (N_24808,N_24669,N_24554);
and U24809 (N_24809,N_24745,N_24667);
and U24810 (N_24810,N_24527,N_24551);
nand U24811 (N_24811,N_24552,N_24605);
xor U24812 (N_24812,N_24539,N_24695);
nor U24813 (N_24813,N_24748,N_24502);
nor U24814 (N_24814,N_24702,N_24555);
xor U24815 (N_24815,N_24683,N_24580);
nand U24816 (N_24816,N_24512,N_24595);
nor U24817 (N_24817,N_24686,N_24696);
nor U24818 (N_24818,N_24503,N_24645);
nor U24819 (N_24819,N_24550,N_24740);
xor U24820 (N_24820,N_24531,N_24516);
or U24821 (N_24821,N_24690,N_24728);
nor U24822 (N_24822,N_24674,N_24600);
nand U24823 (N_24823,N_24741,N_24682);
and U24824 (N_24824,N_24699,N_24726);
xor U24825 (N_24825,N_24610,N_24731);
or U24826 (N_24826,N_24542,N_24647);
or U24827 (N_24827,N_24521,N_24572);
nor U24828 (N_24828,N_24574,N_24614);
nand U24829 (N_24829,N_24543,N_24577);
and U24830 (N_24830,N_24680,N_24534);
nor U24831 (N_24831,N_24662,N_24732);
or U24832 (N_24832,N_24675,N_24583);
nor U24833 (N_24833,N_24506,N_24747);
nand U24834 (N_24834,N_24584,N_24665);
and U24835 (N_24835,N_24529,N_24671);
and U24836 (N_24836,N_24663,N_24668);
nor U24837 (N_24837,N_24536,N_24709);
xnor U24838 (N_24838,N_24629,N_24657);
or U24839 (N_24839,N_24652,N_24681);
or U24840 (N_24840,N_24746,N_24713);
nor U24841 (N_24841,N_24717,N_24714);
nor U24842 (N_24842,N_24607,N_24609);
or U24843 (N_24843,N_24643,N_24547);
xor U24844 (N_24844,N_24710,N_24582);
nor U24845 (N_24845,N_24648,N_24533);
nor U24846 (N_24846,N_24684,N_24604);
nand U24847 (N_24847,N_24565,N_24587);
nor U24848 (N_24848,N_24640,N_24596);
nand U24849 (N_24849,N_24545,N_24508);
nor U24850 (N_24850,N_24559,N_24733);
nor U24851 (N_24851,N_24575,N_24530);
xnor U24852 (N_24852,N_24563,N_24708);
nor U24853 (N_24853,N_24700,N_24571);
xnor U24854 (N_24854,N_24715,N_24744);
nand U24855 (N_24855,N_24513,N_24678);
nor U24856 (N_24856,N_24677,N_24598);
or U24857 (N_24857,N_24653,N_24581);
nor U24858 (N_24858,N_24608,N_24650);
nor U24859 (N_24859,N_24730,N_24517);
xor U24860 (N_24860,N_24719,N_24692);
xor U24861 (N_24861,N_24712,N_24725);
or U24862 (N_24862,N_24711,N_24630);
xor U24863 (N_24863,N_24525,N_24687);
or U24864 (N_24864,N_24727,N_24646);
or U24865 (N_24865,N_24505,N_24672);
nor U24866 (N_24866,N_24644,N_24716);
and U24867 (N_24867,N_24519,N_24718);
nand U24868 (N_24868,N_24573,N_24606);
or U24869 (N_24869,N_24661,N_24538);
xnor U24870 (N_24870,N_24535,N_24670);
or U24871 (N_24871,N_24518,N_24721);
and U24872 (N_24872,N_24697,N_24621);
or U24873 (N_24873,N_24588,N_24553);
nor U24874 (N_24874,N_24570,N_24562);
xnor U24875 (N_24875,N_24550,N_24708);
nand U24876 (N_24876,N_24566,N_24583);
xor U24877 (N_24877,N_24547,N_24543);
nand U24878 (N_24878,N_24602,N_24581);
or U24879 (N_24879,N_24584,N_24540);
and U24880 (N_24880,N_24545,N_24568);
xnor U24881 (N_24881,N_24633,N_24642);
nand U24882 (N_24882,N_24576,N_24534);
xnor U24883 (N_24883,N_24706,N_24664);
or U24884 (N_24884,N_24697,N_24583);
nand U24885 (N_24885,N_24617,N_24546);
or U24886 (N_24886,N_24706,N_24705);
or U24887 (N_24887,N_24744,N_24725);
or U24888 (N_24888,N_24696,N_24735);
and U24889 (N_24889,N_24676,N_24645);
nand U24890 (N_24890,N_24698,N_24532);
xor U24891 (N_24891,N_24522,N_24615);
nand U24892 (N_24892,N_24693,N_24722);
or U24893 (N_24893,N_24708,N_24636);
and U24894 (N_24894,N_24534,N_24639);
or U24895 (N_24895,N_24572,N_24678);
or U24896 (N_24896,N_24528,N_24614);
and U24897 (N_24897,N_24664,N_24696);
and U24898 (N_24898,N_24703,N_24568);
and U24899 (N_24899,N_24739,N_24724);
nand U24900 (N_24900,N_24740,N_24681);
xnor U24901 (N_24901,N_24547,N_24575);
xor U24902 (N_24902,N_24728,N_24669);
and U24903 (N_24903,N_24548,N_24670);
and U24904 (N_24904,N_24577,N_24580);
and U24905 (N_24905,N_24695,N_24645);
and U24906 (N_24906,N_24528,N_24741);
nand U24907 (N_24907,N_24644,N_24674);
and U24908 (N_24908,N_24560,N_24745);
nand U24909 (N_24909,N_24641,N_24720);
nand U24910 (N_24910,N_24682,N_24565);
nand U24911 (N_24911,N_24661,N_24737);
or U24912 (N_24912,N_24541,N_24597);
or U24913 (N_24913,N_24664,N_24555);
nand U24914 (N_24914,N_24545,N_24517);
and U24915 (N_24915,N_24744,N_24612);
xor U24916 (N_24916,N_24544,N_24601);
nand U24917 (N_24917,N_24592,N_24571);
and U24918 (N_24918,N_24535,N_24603);
and U24919 (N_24919,N_24644,N_24638);
and U24920 (N_24920,N_24651,N_24715);
nor U24921 (N_24921,N_24571,N_24643);
xnor U24922 (N_24922,N_24587,N_24638);
nor U24923 (N_24923,N_24710,N_24722);
nand U24924 (N_24924,N_24613,N_24538);
xnor U24925 (N_24925,N_24664,N_24532);
or U24926 (N_24926,N_24741,N_24627);
nand U24927 (N_24927,N_24594,N_24614);
nor U24928 (N_24928,N_24731,N_24583);
nand U24929 (N_24929,N_24542,N_24657);
nor U24930 (N_24930,N_24557,N_24672);
nand U24931 (N_24931,N_24686,N_24660);
and U24932 (N_24932,N_24663,N_24713);
or U24933 (N_24933,N_24624,N_24548);
nor U24934 (N_24934,N_24572,N_24611);
nor U24935 (N_24935,N_24626,N_24511);
and U24936 (N_24936,N_24695,N_24627);
or U24937 (N_24937,N_24677,N_24674);
nand U24938 (N_24938,N_24630,N_24733);
or U24939 (N_24939,N_24525,N_24574);
or U24940 (N_24940,N_24510,N_24578);
and U24941 (N_24941,N_24542,N_24551);
or U24942 (N_24942,N_24694,N_24612);
xnor U24943 (N_24943,N_24624,N_24578);
or U24944 (N_24944,N_24689,N_24715);
and U24945 (N_24945,N_24716,N_24715);
xnor U24946 (N_24946,N_24628,N_24687);
or U24947 (N_24947,N_24701,N_24569);
nor U24948 (N_24948,N_24576,N_24626);
xnor U24949 (N_24949,N_24608,N_24569);
and U24950 (N_24950,N_24662,N_24617);
nor U24951 (N_24951,N_24657,N_24618);
and U24952 (N_24952,N_24671,N_24735);
xnor U24953 (N_24953,N_24559,N_24714);
and U24954 (N_24954,N_24518,N_24526);
xor U24955 (N_24955,N_24542,N_24525);
nand U24956 (N_24956,N_24727,N_24578);
xor U24957 (N_24957,N_24601,N_24540);
or U24958 (N_24958,N_24594,N_24696);
nor U24959 (N_24959,N_24665,N_24617);
nor U24960 (N_24960,N_24648,N_24610);
nand U24961 (N_24961,N_24629,N_24679);
nand U24962 (N_24962,N_24608,N_24564);
xnor U24963 (N_24963,N_24716,N_24534);
nor U24964 (N_24964,N_24655,N_24545);
xnor U24965 (N_24965,N_24584,N_24535);
nor U24966 (N_24966,N_24665,N_24625);
and U24967 (N_24967,N_24732,N_24537);
nand U24968 (N_24968,N_24583,N_24539);
xor U24969 (N_24969,N_24584,N_24611);
or U24970 (N_24970,N_24633,N_24537);
or U24971 (N_24971,N_24518,N_24604);
nand U24972 (N_24972,N_24624,N_24661);
xor U24973 (N_24973,N_24604,N_24637);
nand U24974 (N_24974,N_24600,N_24529);
nand U24975 (N_24975,N_24562,N_24653);
and U24976 (N_24976,N_24616,N_24542);
nand U24977 (N_24977,N_24746,N_24717);
nand U24978 (N_24978,N_24616,N_24640);
nor U24979 (N_24979,N_24534,N_24603);
and U24980 (N_24980,N_24609,N_24697);
xor U24981 (N_24981,N_24600,N_24629);
and U24982 (N_24982,N_24715,N_24693);
xor U24983 (N_24983,N_24717,N_24749);
xnor U24984 (N_24984,N_24515,N_24660);
nor U24985 (N_24985,N_24529,N_24608);
nand U24986 (N_24986,N_24712,N_24599);
or U24987 (N_24987,N_24667,N_24561);
and U24988 (N_24988,N_24640,N_24511);
or U24989 (N_24989,N_24514,N_24734);
nor U24990 (N_24990,N_24561,N_24648);
xnor U24991 (N_24991,N_24599,N_24571);
xor U24992 (N_24992,N_24644,N_24503);
or U24993 (N_24993,N_24547,N_24594);
or U24994 (N_24994,N_24527,N_24562);
and U24995 (N_24995,N_24603,N_24712);
nand U24996 (N_24996,N_24530,N_24599);
and U24997 (N_24997,N_24739,N_24633);
xor U24998 (N_24998,N_24656,N_24586);
xor U24999 (N_24999,N_24546,N_24638);
or UO_0 (O_0,N_24909,N_24852);
nand UO_1 (O_1,N_24990,N_24775);
nand UO_2 (O_2,N_24883,N_24930);
and UO_3 (O_3,N_24803,N_24842);
or UO_4 (O_4,N_24816,N_24908);
nor UO_5 (O_5,N_24906,N_24953);
nor UO_6 (O_6,N_24937,N_24806);
nor UO_7 (O_7,N_24823,N_24768);
nand UO_8 (O_8,N_24794,N_24925);
nor UO_9 (O_9,N_24993,N_24856);
nand UO_10 (O_10,N_24877,N_24973);
or UO_11 (O_11,N_24870,N_24858);
nand UO_12 (O_12,N_24840,N_24972);
nor UO_13 (O_13,N_24761,N_24766);
or UO_14 (O_14,N_24989,N_24923);
nand UO_15 (O_15,N_24977,N_24765);
nor UO_16 (O_16,N_24907,N_24792);
xnor UO_17 (O_17,N_24891,N_24848);
nor UO_18 (O_18,N_24785,N_24833);
xnor UO_19 (O_19,N_24886,N_24996);
or UO_20 (O_20,N_24876,N_24922);
and UO_21 (O_21,N_24959,N_24924);
nand UO_22 (O_22,N_24936,N_24821);
nor UO_23 (O_23,N_24798,N_24797);
nor UO_24 (O_24,N_24865,N_24914);
or UO_25 (O_25,N_24897,N_24793);
or UO_26 (O_26,N_24763,N_24957);
nand UO_27 (O_27,N_24931,N_24903);
or UO_28 (O_28,N_24934,N_24967);
xnor UO_29 (O_29,N_24758,N_24902);
nand UO_30 (O_30,N_24815,N_24759);
or UO_31 (O_31,N_24955,N_24942);
or UO_32 (O_32,N_24752,N_24772);
or UO_33 (O_33,N_24963,N_24829);
nor UO_34 (O_34,N_24928,N_24974);
and UO_35 (O_35,N_24978,N_24893);
xnor UO_36 (O_36,N_24911,N_24968);
nor UO_37 (O_37,N_24777,N_24818);
nor UO_38 (O_38,N_24874,N_24976);
xor UO_39 (O_39,N_24795,N_24921);
nor UO_40 (O_40,N_24807,N_24884);
or UO_41 (O_41,N_24912,N_24875);
and UO_42 (O_42,N_24846,N_24756);
xnor UO_43 (O_43,N_24979,N_24796);
nor UO_44 (O_44,N_24952,N_24787);
nand UO_45 (O_45,N_24982,N_24764);
xor UO_46 (O_46,N_24769,N_24905);
nor UO_47 (O_47,N_24830,N_24898);
xor UO_48 (O_48,N_24809,N_24853);
and UO_49 (O_49,N_24994,N_24887);
nand UO_50 (O_50,N_24948,N_24827);
and UO_51 (O_51,N_24760,N_24981);
xnor UO_52 (O_52,N_24814,N_24826);
xor UO_53 (O_53,N_24944,N_24938);
xor UO_54 (O_54,N_24780,N_24799);
or UO_55 (O_55,N_24885,N_24986);
and UO_56 (O_56,N_24790,N_24964);
and UO_57 (O_57,N_24867,N_24854);
xor UO_58 (O_58,N_24834,N_24776);
nor UO_59 (O_59,N_24956,N_24782);
or UO_60 (O_60,N_24770,N_24961);
nand UO_61 (O_61,N_24863,N_24890);
nor UO_62 (O_62,N_24926,N_24836);
xnor UO_63 (O_63,N_24917,N_24941);
or UO_64 (O_64,N_24958,N_24839);
and UO_65 (O_65,N_24800,N_24945);
or UO_66 (O_66,N_24753,N_24998);
or UO_67 (O_67,N_24828,N_24755);
and UO_68 (O_68,N_24789,N_24757);
nor UO_69 (O_69,N_24824,N_24879);
and UO_70 (O_70,N_24889,N_24985);
nor UO_71 (O_71,N_24849,N_24966);
nor UO_72 (O_72,N_24820,N_24983);
nand UO_73 (O_73,N_24949,N_24951);
and UO_74 (O_74,N_24892,N_24847);
and UO_75 (O_75,N_24791,N_24954);
nand UO_76 (O_76,N_24817,N_24947);
nor UO_77 (O_77,N_24916,N_24751);
xnor UO_78 (O_78,N_24771,N_24943);
xor UO_79 (O_79,N_24881,N_24940);
nor UO_80 (O_80,N_24811,N_24813);
nor UO_81 (O_81,N_24910,N_24971);
and UO_82 (O_82,N_24841,N_24988);
or UO_83 (O_83,N_24918,N_24786);
nor UO_84 (O_84,N_24975,N_24869);
or UO_85 (O_85,N_24984,N_24901);
nor UO_86 (O_86,N_24950,N_24946);
xor UO_87 (O_87,N_24774,N_24778);
or UO_88 (O_88,N_24805,N_24992);
and UO_89 (O_89,N_24788,N_24812);
and UO_90 (O_90,N_24845,N_24880);
xnor UO_91 (O_91,N_24933,N_24873);
xor UO_92 (O_92,N_24860,N_24932);
or UO_93 (O_93,N_24851,N_24804);
nand UO_94 (O_94,N_24832,N_24750);
nor UO_95 (O_95,N_24837,N_24825);
xor UO_96 (O_96,N_24965,N_24808);
nand UO_97 (O_97,N_24991,N_24915);
or UO_98 (O_98,N_24822,N_24920);
or UO_99 (O_99,N_24871,N_24838);
nand UO_100 (O_100,N_24857,N_24831);
nand UO_101 (O_101,N_24802,N_24779);
nor UO_102 (O_102,N_24882,N_24844);
nor UO_103 (O_103,N_24850,N_24754);
or UO_104 (O_104,N_24919,N_24960);
nor UO_105 (O_105,N_24894,N_24962);
nand UO_106 (O_106,N_24801,N_24861);
xor UO_107 (O_107,N_24866,N_24868);
or UO_108 (O_108,N_24997,N_24872);
nand UO_109 (O_109,N_24896,N_24935);
nor UO_110 (O_110,N_24899,N_24970);
nand UO_111 (O_111,N_24781,N_24995);
or UO_112 (O_112,N_24862,N_24987);
or UO_113 (O_113,N_24864,N_24810);
or UO_114 (O_114,N_24843,N_24767);
nand UO_115 (O_115,N_24888,N_24939);
or UO_116 (O_116,N_24900,N_24904);
and UO_117 (O_117,N_24784,N_24980);
xor UO_118 (O_118,N_24855,N_24969);
nand UO_119 (O_119,N_24859,N_24927);
nand UO_120 (O_120,N_24895,N_24783);
nand UO_121 (O_121,N_24819,N_24929);
or UO_122 (O_122,N_24762,N_24835);
and UO_123 (O_123,N_24878,N_24999);
or UO_124 (O_124,N_24913,N_24773);
nand UO_125 (O_125,N_24907,N_24775);
xnor UO_126 (O_126,N_24914,N_24883);
and UO_127 (O_127,N_24851,N_24944);
or UO_128 (O_128,N_24975,N_24817);
and UO_129 (O_129,N_24997,N_24857);
or UO_130 (O_130,N_24978,N_24957);
nand UO_131 (O_131,N_24963,N_24918);
or UO_132 (O_132,N_24864,N_24768);
xor UO_133 (O_133,N_24967,N_24985);
xnor UO_134 (O_134,N_24813,N_24893);
nor UO_135 (O_135,N_24808,N_24943);
xnor UO_136 (O_136,N_24882,N_24764);
and UO_137 (O_137,N_24821,N_24822);
or UO_138 (O_138,N_24919,N_24797);
nand UO_139 (O_139,N_24936,N_24961);
nor UO_140 (O_140,N_24864,N_24829);
nand UO_141 (O_141,N_24861,N_24879);
nand UO_142 (O_142,N_24885,N_24909);
nor UO_143 (O_143,N_24995,N_24950);
and UO_144 (O_144,N_24828,N_24901);
nor UO_145 (O_145,N_24868,N_24862);
and UO_146 (O_146,N_24988,N_24930);
or UO_147 (O_147,N_24765,N_24857);
nor UO_148 (O_148,N_24796,N_24829);
nor UO_149 (O_149,N_24911,N_24801);
nand UO_150 (O_150,N_24983,N_24971);
nand UO_151 (O_151,N_24947,N_24940);
nor UO_152 (O_152,N_24917,N_24783);
or UO_153 (O_153,N_24860,N_24895);
nor UO_154 (O_154,N_24839,N_24777);
and UO_155 (O_155,N_24992,N_24756);
nor UO_156 (O_156,N_24774,N_24751);
or UO_157 (O_157,N_24910,N_24859);
or UO_158 (O_158,N_24901,N_24996);
and UO_159 (O_159,N_24966,N_24867);
and UO_160 (O_160,N_24783,N_24801);
and UO_161 (O_161,N_24901,N_24951);
or UO_162 (O_162,N_24954,N_24961);
nand UO_163 (O_163,N_24956,N_24786);
nand UO_164 (O_164,N_24936,N_24843);
xnor UO_165 (O_165,N_24769,N_24806);
and UO_166 (O_166,N_24964,N_24999);
nor UO_167 (O_167,N_24933,N_24915);
nor UO_168 (O_168,N_24897,N_24802);
nand UO_169 (O_169,N_24895,N_24816);
nand UO_170 (O_170,N_24760,N_24853);
or UO_171 (O_171,N_24858,N_24953);
nand UO_172 (O_172,N_24919,N_24907);
nor UO_173 (O_173,N_24848,N_24835);
nor UO_174 (O_174,N_24756,N_24859);
nand UO_175 (O_175,N_24924,N_24964);
or UO_176 (O_176,N_24950,N_24784);
xnor UO_177 (O_177,N_24810,N_24964);
or UO_178 (O_178,N_24979,N_24995);
and UO_179 (O_179,N_24792,N_24928);
xnor UO_180 (O_180,N_24870,N_24781);
and UO_181 (O_181,N_24980,N_24842);
nand UO_182 (O_182,N_24754,N_24887);
xor UO_183 (O_183,N_24811,N_24750);
nand UO_184 (O_184,N_24967,N_24773);
nand UO_185 (O_185,N_24914,N_24784);
nand UO_186 (O_186,N_24970,N_24965);
nor UO_187 (O_187,N_24832,N_24802);
or UO_188 (O_188,N_24794,N_24924);
and UO_189 (O_189,N_24793,N_24762);
and UO_190 (O_190,N_24818,N_24984);
nand UO_191 (O_191,N_24779,N_24769);
or UO_192 (O_192,N_24885,N_24830);
xnor UO_193 (O_193,N_24801,N_24767);
nand UO_194 (O_194,N_24993,N_24757);
xnor UO_195 (O_195,N_24930,N_24757);
nor UO_196 (O_196,N_24917,N_24884);
or UO_197 (O_197,N_24860,N_24845);
nand UO_198 (O_198,N_24971,N_24750);
xnor UO_199 (O_199,N_24822,N_24803);
nand UO_200 (O_200,N_24837,N_24751);
nor UO_201 (O_201,N_24793,N_24922);
nand UO_202 (O_202,N_24822,N_24869);
nand UO_203 (O_203,N_24846,N_24820);
nand UO_204 (O_204,N_24988,N_24845);
nor UO_205 (O_205,N_24908,N_24821);
xor UO_206 (O_206,N_24901,N_24912);
nor UO_207 (O_207,N_24948,N_24872);
nand UO_208 (O_208,N_24896,N_24850);
or UO_209 (O_209,N_24850,N_24967);
xor UO_210 (O_210,N_24826,N_24994);
nand UO_211 (O_211,N_24779,N_24985);
nor UO_212 (O_212,N_24809,N_24925);
or UO_213 (O_213,N_24978,N_24987);
or UO_214 (O_214,N_24822,N_24788);
and UO_215 (O_215,N_24803,N_24841);
xnor UO_216 (O_216,N_24779,N_24971);
nand UO_217 (O_217,N_24952,N_24954);
nand UO_218 (O_218,N_24815,N_24891);
and UO_219 (O_219,N_24844,N_24911);
or UO_220 (O_220,N_24824,N_24853);
nand UO_221 (O_221,N_24839,N_24754);
nor UO_222 (O_222,N_24780,N_24863);
or UO_223 (O_223,N_24879,N_24848);
xnor UO_224 (O_224,N_24949,N_24907);
xnor UO_225 (O_225,N_24791,N_24751);
or UO_226 (O_226,N_24790,N_24810);
and UO_227 (O_227,N_24803,N_24895);
nand UO_228 (O_228,N_24922,N_24900);
nand UO_229 (O_229,N_24956,N_24909);
or UO_230 (O_230,N_24791,N_24899);
xor UO_231 (O_231,N_24821,N_24914);
nand UO_232 (O_232,N_24827,N_24972);
nand UO_233 (O_233,N_24959,N_24840);
and UO_234 (O_234,N_24769,N_24921);
or UO_235 (O_235,N_24877,N_24774);
nor UO_236 (O_236,N_24897,N_24920);
nand UO_237 (O_237,N_24882,N_24973);
nand UO_238 (O_238,N_24967,N_24953);
or UO_239 (O_239,N_24933,N_24828);
and UO_240 (O_240,N_24806,N_24869);
or UO_241 (O_241,N_24810,N_24819);
or UO_242 (O_242,N_24880,N_24946);
nor UO_243 (O_243,N_24769,N_24823);
or UO_244 (O_244,N_24829,N_24975);
nand UO_245 (O_245,N_24845,N_24805);
or UO_246 (O_246,N_24851,N_24792);
nand UO_247 (O_247,N_24911,N_24781);
or UO_248 (O_248,N_24961,N_24766);
or UO_249 (O_249,N_24904,N_24866);
xnor UO_250 (O_250,N_24960,N_24892);
nand UO_251 (O_251,N_24870,N_24962);
xor UO_252 (O_252,N_24991,N_24949);
xor UO_253 (O_253,N_24971,N_24772);
and UO_254 (O_254,N_24872,N_24868);
or UO_255 (O_255,N_24797,N_24997);
xor UO_256 (O_256,N_24818,N_24779);
and UO_257 (O_257,N_24853,N_24783);
nor UO_258 (O_258,N_24913,N_24834);
nand UO_259 (O_259,N_24788,N_24995);
nor UO_260 (O_260,N_24923,N_24941);
nand UO_261 (O_261,N_24900,N_24770);
nor UO_262 (O_262,N_24773,N_24836);
xor UO_263 (O_263,N_24856,N_24938);
nand UO_264 (O_264,N_24859,N_24831);
and UO_265 (O_265,N_24898,N_24955);
and UO_266 (O_266,N_24810,N_24956);
nand UO_267 (O_267,N_24921,N_24925);
and UO_268 (O_268,N_24827,N_24762);
nand UO_269 (O_269,N_24859,N_24897);
nor UO_270 (O_270,N_24938,N_24995);
nand UO_271 (O_271,N_24920,N_24974);
nand UO_272 (O_272,N_24856,N_24800);
nand UO_273 (O_273,N_24788,N_24918);
and UO_274 (O_274,N_24948,N_24814);
nor UO_275 (O_275,N_24763,N_24976);
and UO_276 (O_276,N_24993,N_24816);
nand UO_277 (O_277,N_24797,N_24781);
nor UO_278 (O_278,N_24782,N_24948);
and UO_279 (O_279,N_24951,N_24927);
xor UO_280 (O_280,N_24980,N_24808);
nand UO_281 (O_281,N_24873,N_24897);
nand UO_282 (O_282,N_24973,N_24878);
and UO_283 (O_283,N_24884,N_24810);
xnor UO_284 (O_284,N_24986,N_24859);
and UO_285 (O_285,N_24921,N_24859);
or UO_286 (O_286,N_24892,N_24780);
xor UO_287 (O_287,N_24992,N_24815);
xnor UO_288 (O_288,N_24817,N_24884);
or UO_289 (O_289,N_24762,N_24881);
nand UO_290 (O_290,N_24796,N_24800);
or UO_291 (O_291,N_24966,N_24831);
and UO_292 (O_292,N_24875,N_24812);
and UO_293 (O_293,N_24970,N_24856);
nor UO_294 (O_294,N_24829,N_24890);
nand UO_295 (O_295,N_24756,N_24986);
nand UO_296 (O_296,N_24950,N_24817);
nor UO_297 (O_297,N_24989,N_24814);
and UO_298 (O_298,N_24891,N_24752);
or UO_299 (O_299,N_24956,N_24930);
nor UO_300 (O_300,N_24978,N_24804);
or UO_301 (O_301,N_24752,N_24948);
or UO_302 (O_302,N_24844,N_24867);
nor UO_303 (O_303,N_24938,N_24796);
or UO_304 (O_304,N_24753,N_24941);
and UO_305 (O_305,N_24972,N_24825);
nand UO_306 (O_306,N_24858,N_24826);
and UO_307 (O_307,N_24810,N_24758);
or UO_308 (O_308,N_24802,N_24986);
nor UO_309 (O_309,N_24957,N_24789);
and UO_310 (O_310,N_24797,N_24869);
and UO_311 (O_311,N_24853,N_24849);
xor UO_312 (O_312,N_24843,N_24835);
nor UO_313 (O_313,N_24884,N_24819);
nand UO_314 (O_314,N_24891,N_24913);
or UO_315 (O_315,N_24909,N_24906);
nand UO_316 (O_316,N_24961,N_24933);
nand UO_317 (O_317,N_24908,N_24799);
nand UO_318 (O_318,N_24771,N_24991);
xor UO_319 (O_319,N_24899,N_24784);
or UO_320 (O_320,N_24798,N_24776);
xnor UO_321 (O_321,N_24940,N_24866);
xor UO_322 (O_322,N_24922,N_24906);
xnor UO_323 (O_323,N_24866,N_24859);
nand UO_324 (O_324,N_24863,N_24809);
or UO_325 (O_325,N_24854,N_24913);
nand UO_326 (O_326,N_24932,N_24783);
nor UO_327 (O_327,N_24877,N_24809);
nor UO_328 (O_328,N_24894,N_24840);
nor UO_329 (O_329,N_24827,N_24942);
nor UO_330 (O_330,N_24753,N_24942);
and UO_331 (O_331,N_24939,N_24836);
or UO_332 (O_332,N_24895,N_24962);
xnor UO_333 (O_333,N_24865,N_24791);
or UO_334 (O_334,N_24758,N_24780);
xor UO_335 (O_335,N_24780,N_24795);
nand UO_336 (O_336,N_24820,N_24799);
and UO_337 (O_337,N_24991,N_24777);
and UO_338 (O_338,N_24853,N_24895);
nand UO_339 (O_339,N_24991,N_24934);
and UO_340 (O_340,N_24830,N_24791);
nor UO_341 (O_341,N_24803,N_24903);
or UO_342 (O_342,N_24885,N_24875);
xnor UO_343 (O_343,N_24817,N_24899);
and UO_344 (O_344,N_24898,N_24899);
nand UO_345 (O_345,N_24966,N_24995);
nand UO_346 (O_346,N_24838,N_24994);
xnor UO_347 (O_347,N_24835,N_24859);
or UO_348 (O_348,N_24850,N_24959);
and UO_349 (O_349,N_24884,N_24755);
nand UO_350 (O_350,N_24970,N_24884);
nand UO_351 (O_351,N_24750,N_24915);
and UO_352 (O_352,N_24948,N_24771);
nor UO_353 (O_353,N_24836,N_24815);
and UO_354 (O_354,N_24915,N_24864);
and UO_355 (O_355,N_24807,N_24888);
nand UO_356 (O_356,N_24931,N_24754);
and UO_357 (O_357,N_24818,N_24919);
nor UO_358 (O_358,N_24896,N_24773);
nor UO_359 (O_359,N_24808,N_24995);
and UO_360 (O_360,N_24877,N_24791);
xnor UO_361 (O_361,N_24873,N_24753);
nor UO_362 (O_362,N_24879,N_24996);
nor UO_363 (O_363,N_24945,N_24975);
and UO_364 (O_364,N_24889,N_24961);
xor UO_365 (O_365,N_24908,N_24847);
or UO_366 (O_366,N_24899,N_24929);
and UO_367 (O_367,N_24965,N_24908);
or UO_368 (O_368,N_24912,N_24841);
or UO_369 (O_369,N_24957,N_24952);
or UO_370 (O_370,N_24905,N_24945);
nand UO_371 (O_371,N_24800,N_24980);
nor UO_372 (O_372,N_24877,N_24944);
nor UO_373 (O_373,N_24844,N_24790);
xnor UO_374 (O_374,N_24787,N_24808);
nand UO_375 (O_375,N_24947,N_24928);
xor UO_376 (O_376,N_24806,N_24890);
or UO_377 (O_377,N_24946,N_24822);
nor UO_378 (O_378,N_24751,N_24804);
xor UO_379 (O_379,N_24847,N_24792);
or UO_380 (O_380,N_24857,N_24853);
and UO_381 (O_381,N_24980,N_24879);
nor UO_382 (O_382,N_24876,N_24775);
and UO_383 (O_383,N_24794,N_24932);
nor UO_384 (O_384,N_24802,N_24865);
and UO_385 (O_385,N_24772,N_24905);
xor UO_386 (O_386,N_24909,N_24984);
xor UO_387 (O_387,N_24754,N_24779);
nand UO_388 (O_388,N_24981,N_24953);
nor UO_389 (O_389,N_24963,N_24877);
nand UO_390 (O_390,N_24895,N_24753);
and UO_391 (O_391,N_24988,N_24946);
xor UO_392 (O_392,N_24946,N_24920);
xnor UO_393 (O_393,N_24812,N_24888);
nor UO_394 (O_394,N_24870,N_24755);
or UO_395 (O_395,N_24781,N_24813);
and UO_396 (O_396,N_24882,N_24872);
nand UO_397 (O_397,N_24863,N_24879);
and UO_398 (O_398,N_24821,N_24875);
xor UO_399 (O_399,N_24839,N_24914);
nor UO_400 (O_400,N_24985,N_24914);
xnor UO_401 (O_401,N_24768,N_24775);
xor UO_402 (O_402,N_24810,N_24874);
and UO_403 (O_403,N_24770,N_24929);
or UO_404 (O_404,N_24841,N_24889);
and UO_405 (O_405,N_24996,N_24760);
nand UO_406 (O_406,N_24886,N_24919);
and UO_407 (O_407,N_24833,N_24967);
and UO_408 (O_408,N_24852,N_24832);
nor UO_409 (O_409,N_24782,N_24765);
nand UO_410 (O_410,N_24841,N_24799);
or UO_411 (O_411,N_24984,N_24980);
xor UO_412 (O_412,N_24767,N_24770);
or UO_413 (O_413,N_24955,N_24944);
xnor UO_414 (O_414,N_24751,N_24937);
nor UO_415 (O_415,N_24867,N_24919);
and UO_416 (O_416,N_24868,N_24897);
and UO_417 (O_417,N_24952,N_24878);
and UO_418 (O_418,N_24919,N_24821);
xor UO_419 (O_419,N_24895,N_24989);
xor UO_420 (O_420,N_24975,N_24889);
nand UO_421 (O_421,N_24810,N_24897);
and UO_422 (O_422,N_24754,N_24897);
nor UO_423 (O_423,N_24780,N_24815);
or UO_424 (O_424,N_24985,N_24986);
nor UO_425 (O_425,N_24908,N_24870);
nor UO_426 (O_426,N_24860,N_24978);
and UO_427 (O_427,N_24921,N_24835);
nand UO_428 (O_428,N_24900,N_24942);
or UO_429 (O_429,N_24930,N_24802);
or UO_430 (O_430,N_24888,N_24752);
or UO_431 (O_431,N_24824,N_24959);
xor UO_432 (O_432,N_24969,N_24753);
xnor UO_433 (O_433,N_24930,N_24780);
or UO_434 (O_434,N_24857,N_24981);
xor UO_435 (O_435,N_24973,N_24755);
and UO_436 (O_436,N_24999,N_24983);
or UO_437 (O_437,N_24842,N_24905);
nand UO_438 (O_438,N_24888,N_24922);
xnor UO_439 (O_439,N_24907,N_24904);
or UO_440 (O_440,N_24795,N_24995);
or UO_441 (O_441,N_24974,N_24993);
or UO_442 (O_442,N_24829,N_24922);
or UO_443 (O_443,N_24792,N_24768);
and UO_444 (O_444,N_24779,N_24755);
or UO_445 (O_445,N_24980,N_24878);
and UO_446 (O_446,N_24805,N_24768);
nor UO_447 (O_447,N_24963,N_24989);
nand UO_448 (O_448,N_24916,N_24769);
and UO_449 (O_449,N_24821,N_24931);
and UO_450 (O_450,N_24881,N_24849);
and UO_451 (O_451,N_24964,N_24836);
nor UO_452 (O_452,N_24862,N_24973);
nor UO_453 (O_453,N_24875,N_24891);
nand UO_454 (O_454,N_24878,N_24961);
xnor UO_455 (O_455,N_24961,N_24847);
nor UO_456 (O_456,N_24893,N_24833);
nor UO_457 (O_457,N_24935,N_24794);
nor UO_458 (O_458,N_24997,N_24800);
or UO_459 (O_459,N_24817,N_24786);
or UO_460 (O_460,N_24995,N_24903);
nand UO_461 (O_461,N_24805,N_24972);
and UO_462 (O_462,N_24817,N_24895);
xnor UO_463 (O_463,N_24993,N_24872);
and UO_464 (O_464,N_24774,N_24938);
and UO_465 (O_465,N_24853,N_24911);
nor UO_466 (O_466,N_24927,N_24888);
or UO_467 (O_467,N_24779,N_24813);
nor UO_468 (O_468,N_24847,N_24987);
or UO_469 (O_469,N_24866,N_24949);
xnor UO_470 (O_470,N_24771,N_24760);
nor UO_471 (O_471,N_24929,N_24807);
nand UO_472 (O_472,N_24999,N_24754);
or UO_473 (O_473,N_24945,N_24994);
or UO_474 (O_474,N_24812,N_24903);
nand UO_475 (O_475,N_24759,N_24903);
and UO_476 (O_476,N_24866,N_24915);
or UO_477 (O_477,N_24988,N_24783);
or UO_478 (O_478,N_24960,N_24762);
nor UO_479 (O_479,N_24990,N_24860);
nor UO_480 (O_480,N_24818,N_24931);
or UO_481 (O_481,N_24964,N_24993);
and UO_482 (O_482,N_24888,N_24765);
or UO_483 (O_483,N_24885,N_24801);
or UO_484 (O_484,N_24963,N_24968);
nor UO_485 (O_485,N_24793,N_24938);
nor UO_486 (O_486,N_24860,N_24910);
nor UO_487 (O_487,N_24805,N_24790);
xnor UO_488 (O_488,N_24865,N_24936);
nand UO_489 (O_489,N_24803,N_24871);
xor UO_490 (O_490,N_24854,N_24835);
nand UO_491 (O_491,N_24805,N_24978);
xnor UO_492 (O_492,N_24957,N_24984);
nand UO_493 (O_493,N_24956,N_24839);
nor UO_494 (O_494,N_24996,N_24874);
nor UO_495 (O_495,N_24863,N_24786);
or UO_496 (O_496,N_24902,N_24910);
nand UO_497 (O_497,N_24904,N_24805);
nor UO_498 (O_498,N_24764,N_24933);
and UO_499 (O_499,N_24944,N_24770);
nand UO_500 (O_500,N_24884,N_24994);
nand UO_501 (O_501,N_24893,N_24943);
nand UO_502 (O_502,N_24845,N_24862);
nand UO_503 (O_503,N_24862,N_24863);
xor UO_504 (O_504,N_24905,N_24866);
xnor UO_505 (O_505,N_24863,N_24967);
and UO_506 (O_506,N_24808,N_24810);
and UO_507 (O_507,N_24786,N_24841);
nand UO_508 (O_508,N_24876,N_24943);
nor UO_509 (O_509,N_24844,N_24980);
and UO_510 (O_510,N_24851,N_24898);
and UO_511 (O_511,N_24827,N_24806);
nor UO_512 (O_512,N_24930,N_24895);
xnor UO_513 (O_513,N_24893,N_24840);
nor UO_514 (O_514,N_24811,N_24927);
nor UO_515 (O_515,N_24949,N_24829);
xor UO_516 (O_516,N_24878,N_24880);
and UO_517 (O_517,N_24912,N_24863);
or UO_518 (O_518,N_24981,N_24766);
nor UO_519 (O_519,N_24906,N_24847);
nand UO_520 (O_520,N_24776,N_24901);
nand UO_521 (O_521,N_24982,N_24984);
or UO_522 (O_522,N_24930,N_24755);
and UO_523 (O_523,N_24809,N_24787);
nand UO_524 (O_524,N_24948,N_24997);
nand UO_525 (O_525,N_24797,N_24907);
nor UO_526 (O_526,N_24920,N_24808);
nand UO_527 (O_527,N_24852,N_24768);
nand UO_528 (O_528,N_24807,N_24906);
nor UO_529 (O_529,N_24992,N_24996);
or UO_530 (O_530,N_24832,N_24881);
xnor UO_531 (O_531,N_24909,N_24875);
nor UO_532 (O_532,N_24800,N_24809);
nor UO_533 (O_533,N_24855,N_24963);
xnor UO_534 (O_534,N_24884,N_24993);
xnor UO_535 (O_535,N_24966,N_24895);
and UO_536 (O_536,N_24869,N_24796);
nand UO_537 (O_537,N_24778,N_24913);
nor UO_538 (O_538,N_24859,N_24992);
xnor UO_539 (O_539,N_24891,N_24755);
and UO_540 (O_540,N_24779,N_24883);
xnor UO_541 (O_541,N_24988,N_24976);
nor UO_542 (O_542,N_24856,N_24751);
nor UO_543 (O_543,N_24759,N_24898);
xor UO_544 (O_544,N_24979,N_24936);
or UO_545 (O_545,N_24779,N_24944);
or UO_546 (O_546,N_24758,N_24886);
xor UO_547 (O_547,N_24793,N_24967);
or UO_548 (O_548,N_24959,N_24765);
nor UO_549 (O_549,N_24972,N_24962);
or UO_550 (O_550,N_24835,N_24960);
xor UO_551 (O_551,N_24887,N_24966);
and UO_552 (O_552,N_24902,N_24841);
nand UO_553 (O_553,N_24964,N_24755);
xor UO_554 (O_554,N_24796,N_24753);
nand UO_555 (O_555,N_24890,N_24975);
or UO_556 (O_556,N_24784,N_24971);
and UO_557 (O_557,N_24917,N_24955);
xor UO_558 (O_558,N_24829,N_24762);
or UO_559 (O_559,N_24969,N_24772);
nor UO_560 (O_560,N_24751,N_24886);
nor UO_561 (O_561,N_24980,N_24991);
nand UO_562 (O_562,N_24993,N_24914);
xor UO_563 (O_563,N_24893,N_24779);
nor UO_564 (O_564,N_24934,N_24928);
and UO_565 (O_565,N_24774,N_24984);
xnor UO_566 (O_566,N_24772,N_24849);
nand UO_567 (O_567,N_24755,N_24960);
and UO_568 (O_568,N_24766,N_24930);
nand UO_569 (O_569,N_24789,N_24883);
and UO_570 (O_570,N_24812,N_24997);
xnor UO_571 (O_571,N_24854,N_24992);
xnor UO_572 (O_572,N_24787,N_24870);
nand UO_573 (O_573,N_24957,N_24753);
or UO_574 (O_574,N_24953,N_24942);
and UO_575 (O_575,N_24928,N_24797);
and UO_576 (O_576,N_24817,N_24858);
nor UO_577 (O_577,N_24942,N_24878);
xor UO_578 (O_578,N_24868,N_24941);
nor UO_579 (O_579,N_24936,N_24911);
xor UO_580 (O_580,N_24954,N_24825);
nand UO_581 (O_581,N_24829,N_24797);
xnor UO_582 (O_582,N_24905,N_24965);
xnor UO_583 (O_583,N_24896,N_24895);
or UO_584 (O_584,N_24986,N_24770);
nand UO_585 (O_585,N_24970,N_24984);
nor UO_586 (O_586,N_24885,N_24997);
xnor UO_587 (O_587,N_24900,N_24810);
and UO_588 (O_588,N_24965,N_24946);
or UO_589 (O_589,N_24953,N_24925);
and UO_590 (O_590,N_24950,N_24965);
nand UO_591 (O_591,N_24998,N_24843);
and UO_592 (O_592,N_24927,N_24842);
and UO_593 (O_593,N_24935,N_24760);
xor UO_594 (O_594,N_24944,N_24812);
nor UO_595 (O_595,N_24932,N_24752);
nand UO_596 (O_596,N_24859,N_24874);
xor UO_597 (O_597,N_24961,N_24885);
or UO_598 (O_598,N_24978,N_24903);
nand UO_599 (O_599,N_24841,N_24999);
nor UO_600 (O_600,N_24887,N_24927);
and UO_601 (O_601,N_24972,N_24798);
nor UO_602 (O_602,N_24968,N_24832);
nor UO_603 (O_603,N_24964,N_24829);
or UO_604 (O_604,N_24823,N_24945);
nor UO_605 (O_605,N_24833,N_24966);
xor UO_606 (O_606,N_24909,N_24901);
nand UO_607 (O_607,N_24868,N_24777);
and UO_608 (O_608,N_24883,N_24962);
nand UO_609 (O_609,N_24892,N_24810);
xnor UO_610 (O_610,N_24896,N_24758);
xnor UO_611 (O_611,N_24781,N_24902);
xnor UO_612 (O_612,N_24911,N_24814);
nand UO_613 (O_613,N_24769,N_24774);
nor UO_614 (O_614,N_24834,N_24887);
nor UO_615 (O_615,N_24773,N_24972);
and UO_616 (O_616,N_24839,N_24937);
nor UO_617 (O_617,N_24865,N_24926);
nor UO_618 (O_618,N_24762,N_24797);
nand UO_619 (O_619,N_24921,N_24860);
and UO_620 (O_620,N_24756,N_24865);
xnor UO_621 (O_621,N_24981,N_24940);
nor UO_622 (O_622,N_24931,N_24820);
nor UO_623 (O_623,N_24913,N_24770);
and UO_624 (O_624,N_24990,N_24781);
and UO_625 (O_625,N_24849,N_24949);
and UO_626 (O_626,N_24800,N_24928);
and UO_627 (O_627,N_24777,N_24877);
nand UO_628 (O_628,N_24807,N_24935);
and UO_629 (O_629,N_24783,N_24984);
and UO_630 (O_630,N_24774,N_24793);
or UO_631 (O_631,N_24864,N_24982);
nand UO_632 (O_632,N_24761,N_24903);
xor UO_633 (O_633,N_24930,N_24986);
and UO_634 (O_634,N_24902,N_24860);
nand UO_635 (O_635,N_24986,N_24928);
and UO_636 (O_636,N_24981,N_24989);
xnor UO_637 (O_637,N_24856,N_24815);
nor UO_638 (O_638,N_24817,N_24783);
nor UO_639 (O_639,N_24767,N_24958);
xnor UO_640 (O_640,N_24788,N_24777);
nand UO_641 (O_641,N_24912,N_24897);
nand UO_642 (O_642,N_24974,N_24969);
xnor UO_643 (O_643,N_24820,N_24908);
and UO_644 (O_644,N_24906,N_24758);
or UO_645 (O_645,N_24882,N_24754);
and UO_646 (O_646,N_24954,N_24948);
nor UO_647 (O_647,N_24758,N_24894);
nor UO_648 (O_648,N_24792,N_24776);
or UO_649 (O_649,N_24756,N_24934);
xor UO_650 (O_650,N_24790,N_24891);
xor UO_651 (O_651,N_24812,N_24893);
or UO_652 (O_652,N_24975,N_24850);
nand UO_653 (O_653,N_24769,N_24950);
and UO_654 (O_654,N_24944,N_24891);
xor UO_655 (O_655,N_24941,N_24938);
nand UO_656 (O_656,N_24794,N_24791);
and UO_657 (O_657,N_24961,N_24892);
and UO_658 (O_658,N_24806,N_24836);
or UO_659 (O_659,N_24880,N_24910);
or UO_660 (O_660,N_24800,N_24822);
nand UO_661 (O_661,N_24895,N_24820);
and UO_662 (O_662,N_24924,N_24960);
and UO_663 (O_663,N_24790,N_24905);
xnor UO_664 (O_664,N_24961,N_24752);
and UO_665 (O_665,N_24913,N_24769);
xor UO_666 (O_666,N_24878,N_24771);
or UO_667 (O_667,N_24756,N_24835);
xor UO_668 (O_668,N_24911,N_24785);
and UO_669 (O_669,N_24844,N_24913);
nor UO_670 (O_670,N_24953,N_24962);
nand UO_671 (O_671,N_24934,N_24987);
nand UO_672 (O_672,N_24934,N_24867);
or UO_673 (O_673,N_24889,N_24984);
and UO_674 (O_674,N_24859,N_24822);
nand UO_675 (O_675,N_24815,N_24938);
xor UO_676 (O_676,N_24777,N_24884);
nor UO_677 (O_677,N_24916,N_24806);
nor UO_678 (O_678,N_24827,N_24904);
nand UO_679 (O_679,N_24808,N_24875);
xnor UO_680 (O_680,N_24881,N_24948);
or UO_681 (O_681,N_24860,N_24907);
xnor UO_682 (O_682,N_24750,N_24880);
nor UO_683 (O_683,N_24968,N_24754);
nor UO_684 (O_684,N_24991,N_24977);
nand UO_685 (O_685,N_24797,N_24902);
nand UO_686 (O_686,N_24935,N_24879);
nor UO_687 (O_687,N_24840,N_24872);
nand UO_688 (O_688,N_24962,N_24771);
xnor UO_689 (O_689,N_24809,N_24902);
and UO_690 (O_690,N_24785,N_24838);
or UO_691 (O_691,N_24817,N_24940);
nor UO_692 (O_692,N_24759,N_24940);
and UO_693 (O_693,N_24988,N_24821);
nor UO_694 (O_694,N_24883,N_24938);
xor UO_695 (O_695,N_24752,N_24846);
and UO_696 (O_696,N_24789,N_24755);
xor UO_697 (O_697,N_24999,N_24854);
nor UO_698 (O_698,N_24994,N_24970);
nand UO_699 (O_699,N_24979,N_24784);
nand UO_700 (O_700,N_24896,N_24787);
or UO_701 (O_701,N_24935,N_24764);
and UO_702 (O_702,N_24761,N_24835);
xnor UO_703 (O_703,N_24846,N_24777);
and UO_704 (O_704,N_24947,N_24919);
or UO_705 (O_705,N_24763,N_24879);
nand UO_706 (O_706,N_24841,N_24837);
or UO_707 (O_707,N_24923,N_24771);
nor UO_708 (O_708,N_24865,N_24835);
nand UO_709 (O_709,N_24898,N_24986);
nand UO_710 (O_710,N_24955,N_24997);
nor UO_711 (O_711,N_24901,N_24960);
and UO_712 (O_712,N_24961,N_24989);
nand UO_713 (O_713,N_24888,N_24894);
xnor UO_714 (O_714,N_24920,N_24880);
nor UO_715 (O_715,N_24898,N_24758);
or UO_716 (O_716,N_24897,N_24914);
nor UO_717 (O_717,N_24969,N_24803);
or UO_718 (O_718,N_24939,N_24906);
and UO_719 (O_719,N_24840,N_24996);
nor UO_720 (O_720,N_24883,N_24910);
nand UO_721 (O_721,N_24907,N_24755);
xor UO_722 (O_722,N_24865,N_24905);
xor UO_723 (O_723,N_24923,N_24890);
or UO_724 (O_724,N_24857,N_24988);
or UO_725 (O_725,N_24839,N_24981);
or UO_726 (O_726,N_24791,N_24938);
or UO_727 (O_727,N_24937,N_24962);
xor UO_728 (O_728,N_24794,N_24907);
and UO_729 (O_729,N_24892,N_24799);
nor UO_730 (O_730,N_24939,N_24999);
nand UO_731 (O_731,N_24852,N_24779);
nand UO_732 (O_732,N_24797,N_24890);
nor UO_733 (O_733,N_24910,N_24908);
xnor UO_734 (O_734,N_24969,N_24921);
and UO_735 (O_735,N_24964,N_24838);
or UO_736 (O_736,N_24991,N_24930);
nor UO_737 (O_737,N_24893,N_24948);
nor UO_738 (O_738,N_24887,N_24971);
nand UO_739 (O_739,N_24891,N_24878);
and UO_740 (O_740,N_24888,N_24780);
and UO_741 (O_741,N_24933,N_24972);
nand UO_742 (O_742,N_24896,N_24937);
and UO_743 (O_743,N_24846,N_24960);
xnor UO_744 (O_744,N_24833,N_24769);
and UO_745 (O_745,N_24769,N_24997);
or UO_746 (O_746,N_24764,N_24973);
nand UO_747 (O_747,N_24979,N_24752);
nor UO_748 (O_748,N_24790,N_24757);
and UO_749 (O_749,N_24954,N_24829);
nor UO_750 (O_750,N_24773,N_24992);
and UO_751 (O_751,N_24985,N_24857);
nand UO_752 (O_752,N_24900,N_24790);
or UO_753 (O_753,N_24888,N_24903);
or UO_754 (O_754,N_24877,N_24827);
or UO_755 (O_755,N_24902,N_24899);
nand UO_756 (O_756,N_24806,N_24960);
xor UO_757 (O_757,N_24959,N_24930);
and UO_758 (O_758,N_24822,N_24973);
nand UO_759 (O_759,N_24815,N_24880);
nand UO_760 (O_760,N_24756,N_24955);
or UO_761 (O_761,N_24756,N_24967);
nor UO_762 (O_762,N_24991,N_24826);
nor UO_763 (O_763,N_24799,N_24945);
and UO_764 (O_764,N_24901,N_24759);
and UO_765 (O_765,N_24752,N_24916);
nand UO_766 (O_766,N_24789,N_24872);
nor UO_767 (O_767,N_24896,N_24927);
nor UO_768 (O_768,N_24937,N_24923);
nor UO_769 (O_769,N_24872,N_24812);
or UO_770 (O_770,N_24821,N_24923);
nor UO_771 (O_771,N_24757,N_24799);
or UO_772 (O_772,N_24874,N_24809);
nand UO_773 (O_773,N_24777,N_24754);
nor UO_774 (O_774,N_24920,N_24957);
nand UO_775 (O_775,N_24893,N_24929);
nor UO_776 (O_776,N_24808,N_24962);
or UO_777 (O_777,N_24942,N_24855);
or UO_778 (O_778,N_24899,N_24948);
xor UO_779 (O_779,N_24922,N_24770);
nor UO_780 (O_780,N_24751,N_24826);
nor UO_781 (O_781,N_24988,N_24775);
or UO_782 (O_782,N_24967,N_24993);
nand UO_783 (O_783,N_24963,N_24967);
or UO_784 (O_784,N_24804,N_24881);
and UO_785 (O_785,N_24797,N_24911);
and UO_786 (O_786,N_24851,N_24809);
xnor UO_787 (O_787,N_24953,N_24851);
or UO_788 (O_788,N_24928,N_24958);
nor UO_789 (O_789,N_24952,N_24859);
or UO_790 (O_790,N_24859,N_24949);
nor UO_791 (O_791,N_24859,N_24871);
nor UO_792 (O_792,N_24837,N_24927);
nor UO_793 (O_793,N_24894,N_24965);
nand UO_794 (O_794,N_24787,N_24751);
xor UO_795 (O_795,N_24798,N_24778);
and UO_796 (O_796,N_24958,N_24819);
nand UO_797 (O_797,N_24864,N_24792);
and UO_798 (O_798,N_24763,N_24872);
nand UO_799 (O_799,N_24939,N_24973);
nor UO_800 (O_800,N_24875,N_24782);
or UO_801 (O_801,N_24877,N_24958);
nor UO_802 (O_802,N_24913,N_24756);
xnor UO_803 (O_803,N_24821,N_24845);
or UO_804 (O_804,N_24849,N_24816);
nor UO_805 (O_805,N_24800,N_24773);
nor UO_806 (O_806,N_24796,N_24836);
nor UO_807 (O_807,N_24944,N_24959);
and UO_808 (O_808,N_24822,N_24752);
nor UO_809 (O_809,N_24999,N_24906);
or UO_810 (O_810,N_24902,N_24960);
nor UO_811 (O_811,N_24813,N_24948);
and UO_812 (O_812,N_24828,N_24909);
or UO_813 (O_813,N_24988,N_24768);
and UO_814 (O_814,N_24902,N_24940);
nor UO_815 (O_815,N_24837,N_24768);
and UO_816 (O_816,N_24938,N_24818);
xor UO_817 (O_817,N_24813,N_24816);
xnor UO_818 (O_818,N_24754,N_24985);
nand UO_819 (O_819,N_24847,N_24944);
and UO_820 (O_820,N_24910,N_24885);
and UO_821 (O_821,N_24943,N_24760);
nand UO_822 (O_822,N_24976,N_24824);
or UO_823 (O_823,N_24791,N_24903);
and UO_824 (O_824,N_24786,N_24770);
and UO_825 (O_825,N_24976,N_24765);
and UO_826 (O_826,N_24879,N_24777);
nor UO_827 (O_827,N_24753,N_24890);
and UO_828 (O_828,N_24782,N_24794);
nor UO_829 (O_829,N_24906,N_24759);
or UO_830 (O_830,N_24754,N_24874);
nor UO_831 (O_831,N_24750,N_24857);
nor UO_832 (O_832,N_24908,N_24999);
xnor UO_833 (O_833,N_24974,N_24909);
and UO_834 (O_834,N_24875,N_24921);
nor UO_835 (O_835,N_24895,N_24754);
or UO_836 (O_836,N_24754,N_24990);
xnor UO_837 (O_837,N_24807,N_24976);
or UO_838 (O_838,N_24895,N_24784);
or UO_839 (O_839,N_24804,N_24997);
and UO_840 (O_840,N_24861,N_24886);
and UO_841 (O_841,N_24755,N_24839);
or UO_842 (O_842,N_24948,N_24949);
nor UO_843 (O_843,N_24768,N_24962);
nor UO_844 (O_844,N_24923,N_24815);
or UO_845 (O_845,N_24846,N_24817);
nor UO_846 (O_846,N_24983,N_24887);
and UO_847 (O_847,N_24900,N_24872);
or UO_848 (O_848,N_24987,N_24886);
nand UO_849 (O_849,N_24966,N_24782);
and UO_850 (O_850,N_24814,N_24865);
and UO_851 (O_851,N_24990,N_24961);
nor UO_852 (O_852,N_24941,N_24764);
nand UO_853 (O_853,N_24973,N_24853);
nor UO_854 (O_854,N_24929,N_24793);
nor UO_855 (O_855,N_24964,N_24817);
or UO_856 (O_856,N_24819,N_24893);
nor UO_857 (O_857,N_24948,N_24897);
and UO_858 (O_858,N_24952,N_24863);
and UO_859 (O_859,N_24964,N_24797);
nor UO_860 (O_860,N_24924,N_24803);
nor UO_861 (O_861,N_24823,N_24855);
and UO_862 (O_862,N_24822,N_24807);
and UO_863 (O_863,N_24859,N_24772);
or UO_864 (O_864,N_24794,N_24920);
xor UO_865 (O_865,N_24951,N_24820);
xnor UO_866 (O_866,N_24868,N_24821);
xor UO_867 (O_867,N_24817,N_24757);
nand UO_868 (O_868,N_24947,N_24876);
or UO_869 (O_869,N_24764,N_24917);
xor UO_870 (O_870,N_24771,N_24754);
nand UO_871 (O_871,N_24989,N_24831);
xor UO_872 (O_872,N_24756,N_24887);
xor UO_873 (O_873,N_24846,N_24809);
xor UO_874 (O_874,N_24908,N_24974);
nor UO_875 (O_875,N_24858,N_24992);
nor UO_876 (O_876,N_24778,N_24970);
and UO_877 (O_877,N_24875,N_24836);
or UO_878 (O_878,N_24788,N_24923);
or UO_879 (O_879,N_24762,N_24807);
nor UO_880 (O_880,N_24833,N_24923);
nand UO_881 (O_881,N_24836,N_24750);
nor UO_882 (O_882,N_24960,N_24950);
xnor UO_883 (O_883,N_24803,N_24812);
xor UO_884 (O_884,N_24771,N_24997);
or UO_885 (O_885,N_24902,N_24956);
or UO_886 (O_886,N_24900,N_24884);
and UO_887 (O_887,N_24991,N_24840);
and UO_888 (O_888,N_24844,N_24879);
xor UO_889 (O_889,N_24931,N_24846);
nor UO_890 (O_890,N_24810,N_24910);
or UO_891 (O_891,N_24912,N_24756);
and UO_892 (O_892,N_24848,N_24863);
and UO_893 (O_893,N_24814,N_24752);
nor UO_894 (O_894,N_24829,N_24765);
nand UO_895 (O_895,N_24865,N_24774);
nor UO_896 (O_896,N_24920,N_24860);
xnor UO_897 (O_897,N_24760,N_24997);
xor UO_898 (O_898,N_24960,N_24832);
xnor UO_899 (O_899,N_24792,N_24982);
or UO_900 (O_900,N_24919,N_24767);
or UO_901 (O_901,N_24834,N_24984);
or UO_902 (O_902,N_24993,N_24943);
nor UO_903 (O_903,N_24937,N_24809);
and UO_904 (O_904,N_24884,N_24885);
nor UO_905 (O_905,N_24892,N_24957);
or UO_906 (O_906,N_24952,N_24816);
and UO_907 (O_907,N_24990,N_24891);
xnor UO_908 (O_908,N_24785,N_24938);
or UO_909 (O_909,N_24779,N_24789);
xnor UO_910 (O_910,N_24862,N_24775);
xnor UO_911 (O_911,N_24768,N_24879);
xor UO_912 (O_912,N_24893,N_24829);
nand UO_913 (O_913,N_24881,N_24772);
nor UO_914 (O_914,N_24841,N_24990);
xnor UO_915 (O_915,N_24936,N_24799);
nor UO_916 (O_916,N_24845,N_24901);
or UO_917 (O_917,N_24763,N_24965);
or UO_918 (O_918,N_24804,N_24750);
and UO_919 (O_919,N_24929,N_24782);
xor UO_920 (O_920,N_24859,N_24783);
nor UO_921 (O_921,N_24964,N_24807);
and UO_922 (O_922,N_24940,N_24825);
and UO_923 (O_923,N_24981,N_24844);
and UO_924 (O_924,N_24917,N_24939);
nand UO_925 (O_925,N_24979,N_24908);
nor UO_926 (O_926,N_24838,N_24790);
or UO_927 (O_927,N_24770,N_24794);
nor UO_928 (O_928,N_24867,N_24935);
and UO_929 (O_929,N_24778,N_24941);
or UO_930 (O_930,N_24764,N_24983);
nand UO_931 (O_931,N_24841,N_24808);
nor UO_932 (O_932,N_24870,N_24832);
or UO_933 (O_933,N_24882,N_24989);
nor UO_934 (O_934,N_24912,N_24950);
or UO_935 (O_935,N_24858,N_24788);
nor UO_936 (O_936,N_24787,N_24933);
nor UO_937 (O_937,N_24771,N_24842);
nand UO_938 (O_938,N_24826,N_24945);
nand UO_939 (O_939,N_24976,N_24953);
nand UO_940 (O_940,N_24840,N_24988);
xnor UO_941 (O_941,N_24937,N_24964);
xor UO_942 (O_942,N_24974,N_24922);
and UO_943 (O_943,N_24863,N_24983);
xor UO_944 (O_944,N_24767,N_24968);
nor UO_945 (O_945,N_24879,N_24892);
xor UO_946 (O_946,N_24975,N_24967);
nor UO_947 (O_947,N_24814,N_24824);
nand UO_948 (O_948,N_24994,N_24793);
xnor UO_949 (O_949,N_24864,N_24755);
xor UO_950 (O_950,N_24934,N_24965);
nand UO_951 (O_951,N_24948,N_24818);
nor UO_952 (O_952,N_24771,N_24899);
and UO_953 (O_953,N_24942,N_24947);
xnor UO_954 (O_954,N_24899,N_24828);
nor UO_955 (O_955,N_24928,N_24848);
and UO_956 (O_956,N_24876,N_24960);
nand UO_957 (O_957,N_24784,N_24827);
nor UO_958 (O_958,N_24852,N_24879);
or UO_959 (O_959,N_24798,N_24887);
nor UO_960 (O_960,N_24878,N_24839);
nor UO_961 (O_961,N_24988,N_24779);
and UO_962 (O_962,N_24835,N_24982);
xnor UO_963 (O_963,N_24824,N_24857);
nor UO_964 (O_964,N_24819,N_24987);
nand UO_965 (O_965,N_24757,N_24756);
or UO_966 (O_966,N_24778,N_24883);
and UO_967 (O_967,N_24961,N_24893);
nor UO_968 (O_968,N_24911,N_24945);
or UO_969 (O_969,N_24787,N_24805);
or UO_970 (O_970,N_24918,N_24992);
nor UO_971 (O_971,N_24925,N_24812);
xor UO_972 (O_972,N_24865,N_24750);
xor UO_973 (O_973,N_24822,N_24899);
nor UO_974 (O_974,N_24778,N_24833);
or UO_975 (O_975,N_24893,N_24769);
and UO_976 (O_976,N_24755,N_24904);
nand UO_977 (O_977,N_24924,N_24797);
and UO_978 (O_978,N_24870,N_24817);
xor UO_979 (O_979,N_24982,N_24955);
or UO_980 (O_980,N_24977,N_24954);
nand UO_981 (O_981,N_24880,N_24998);
nand UO_982 (O_982,N_24799,N_24913);
nand UO_983 (O_983,N_24857,N_24948);
or UO_984 (O_984,N_24858,N_24819);
or UO_985 (O_985,N_24992,N_24863);
nand UO_986 (O_986,N_24754,N_24827);
or UO_987 (O_987,N_24900,N_24804);
nand UO_988 (O_988,N_24869,N_24872);
nor UO_989 (O_989,N_24849,N_24751);
nor UO_990 (O_990,N_24841,N_24956);
xnor UO_991 (O_991,N_24751,N_24768);
and UO_992 (O_992,N_24944,N_24875);
xnor UO_993 (O_993,N_24806,N_24811);
xor UO_994 (O_994,N_24793,N_24754);
and UO_995 (O_995,N_24930,N_24750);
nor UO_996 (O_996,N_24925,N_24820);
nand UO_997 (O_997,N_24972,N_24771);
nand UO_998 (O_998,N_24853,N_24832);
nand UO_999 (O_999,N_24912,N_24846);
nor UO_1000 (O_1000,N_24864,N_24961);
and UO_1001 (O_1001,N_24920,N_24886);
or UO_1002 (O_1002,N_24855,N_24758);
or UO_1003 (O_1003,N_24945,N_24930);
nand UO_1004 (O_1004,N_24777,N_24764);
xor UO_1005 (O_1005,N_24805,N_24783);
xnor UO_1006 (O_1006,N_24835,N_24819);
xor UO_1007 (O_1007,N_24908,N_24789);
or UO_1008 (O_1008,N_24798,N_24851);
and UO_1009 (O_1009,N_24890,N_24956);
and UO_1010 (O_1010,N_24821,N_24757);
and UO_1011 (O_1011,N_24771,N_24765);
xnor UO_1012 (O_1012,N_24807,N_24934);
nand UO_1013 (O_1013,N_24844,N_24945);
xor UO_1014 (O_1014,N_24815,N_24777);
xnor UO_1015 (O_1015,N_24946,N_24910);
and UO_1016 (O_1016,N_24873,N_24799);
and UO_1017 (O_1017,N_24859,N_24808);
or UO_1018 (O_1018,N_24973,N_24871);
nor UO_1019 (O_1019,N_24862,N_24974);
nor UO_1020 (O_1020,N_24800,N_24982);
and UO_1021 (O_1021,N_24970,N_24843);
nor UO_1022 (O_1022,N_24759,N_24960);
or UO_1023 (O_1023,N_24786,N_24844);
or UO_1024 (O_1024,N_24909,N_24960);
and UO_1025 (O_1025,N_24885,N_24846);
and UO_1026 (O_1026,N_24789,N_24771);
nor UO_1027 (O_1027,N_24910,N_24760);
and UO_1028 (O_1028,N_24826,N_24885);
and UO_1029 (O_1029,N_24824,N_24855);
xor UO_1030 (O_1030,N_24824,N_24790);
nand UO_1031 (O_1031,N_24836,N_24922);
nor UO_1032 (O_1032,N_24909,N_24765);
and UO_1033 (O_1033,N_24845,N_24974);
nor UO_1034 (O_1034,N_24948,N_24985);
and UO_1035 (O_1035,N_24905,N_24869);
and UO_1036 (O_1036,N_24795,N_24758);
nand UO_1037 (O_1037,N_24784,N_24947);
or UO_1038 (O_1038,N_24944,N_24777);
nor UO_1039 (O_1039,N_24885,N_24954);
and UO_1040 (O_1040,N_24908,N_24829);
nand UO_1041 (O_1041,N_24789,N_24995);
and UO_1042 (O_1042,N_24876,N_24909);
xor UO_1043 (O_1043,N_24788,N_24813);
and UO_1044 (O_1044,N_24750,N_24776);
and UO_1045 (O_1045,N_24920,N_24899);
nand UO_1046 (O_1046,N_24823,N_24806);
and UO_1047 (O_1047,N_24837,N_24932);
nand UO_1048 (O_1048,N_24852,N_24815);
and UO_1049 (O_1049,N_24998,N_24826);
nand UO_1050 (O_1050,N_24787,N_24922);
or UO_1051 (O_1051,N_24886,N_24782);
nand UO_1052 (O_1052,N_24994,N_24819);
and UO_1053 (O_1053,N_24867,N_24932);
nand UO_1054 (O_1054,N_24817,N_24995);
nand UO_1055 (O_1055,N_24979,N_24850);
and UO_1056 (O_1056,N_24874,N_24751);
xnor UO_1057 (O_1057,N_24895,N_24968);
and UO_1058 (O_1058,N_24826,N_24808);
nor UO_1059 (O_1059,N_24770,N_24838);
xor UO_1060 (O_1060,N_24854,N_24906);
nand UO_1061 (O_1061,N_24814,N_24941);
or UO_1062 (O_1062,N_24757,N_24978);
or UO_1063 (O_1063,N_24937,N_24934);
or UO_1064 (O_1064,N_24803,N_24827);
nor UO_1065 (O_1065,N_24924,N_24784);
nor UO_1066 (O_1066,N_24765,N_24889);
xnor UO_1067 (O_1067,N_24774,N_24960);
nor UO_1068 (O_1068,N_24804,N_24877);
xor UO_1069 (O_1069,N_24990,N_24883);
or UO_1070 (O_1070,N_24843,N_24846);
xnor UO_1071 (O_1071,N_24994,N_24922);
nor UO_1072 (O_1072,N_24800,N_24799);
xor UO_1073 (O_1073,N_24827,N_24901);
and UO_1074 (O_1074,N_24754,N_24934);
nor UO_1075 (O_1075,N_24762,N_24872);
nand UO_1076 (O_1076,N_24956,N_24914);
or UO_1077 (O_1077,N_24959,N_24934);
nand UO_1078 (O_1078,N_24827,N_24937);
nand UO_1079 (O_1079,N_24764,N_24924);
and UO_1080 (O_1080,N_24795,N_24752);
xnor UO_1081 (O_1081,N_24906,N_24901);
nand UO_1082 (O_1082,N_24826,N_24975);
nand UO_1083 (O_1083,N_24799,N_24831);
xnor UO_1084 (O_1084,N_24995,N_24831);
and UO_1085 (O_1085,N_24815,N_24995);
xor UO_1086 (O_1086,N_24752,N_24755);
nor UO_1087 (O_1087,N_24768,N_24763);
and UO_1088 (O_1088,N_24770,N_24869);
nand UO_1089 (O_1089,N_24837,N_24988);
or UO_1090 (O_1090,N_24911,N_24850);
nand UO_1091 (O_1091,N_24781,N_24844);
nor UO_1092 (O_1092,N_24942,N_24935);
nand UO_1093 (O_1093,N_24824,N_24961);
or UO_1094 (O_1094,N_24983,N_24981);
nand UO_1095 (O_1095,N_24823,N_24763);
nor UO_1096 (O_1096,N_24936,N_24750);
nor UO_1097 (O_1097,N_24811,N_24770);
and UO_1098 (O_1098,N_24986,N_24854);
or UO_1099 (O_1099,N_24983,N_24991);
nor UO_1100 (O_1100,N_24827,N_24875);
or UO_1101 (O_1101,N_24798,N_24919);
nand UO_1102 (O_1102,N_24961,N_24757);
and UO_1103 (O_1103,N_24986,N_24921);
nand UO_1104 (O_1104,N_24775,N_24916);
or UO_1105 (O_1105,N_24939,N_24912);
nand UO_1106 (O_1106,N_24933,N_24955);
and UO_1107 (O_1107,N_24826,N_24817);
xnor UO_1108 (O_1108,N_24788,N_24861);
nor UO_1109 (O_1109,N_24856,N_24897);
xnor UO_1110 (O_1110,N_24939,N_24848);
xnor UO_1111 (O_1111,N_24886,N_24780);
nand UO_1112 (O_1112,N_24799,N_24840);
or UO_1113 (O_1113,N_24877,N_24949);
nand UO_1114 (O_1114,N_24960,N_24792);
nor UO_1115 (O_1115,N_24757,N_24884);
nor UO_1116 (O_1116,N_24953,N_24982);
nand UO_1117 (O_1117,N_24929,N_24814);
nand UO_1118 (O_1118,N_24959,N_24955);
nor UO_1119 (O_1119,N_24830,N_24949);
nand UO_1120 (O_1120,N_24853,N_24886);
xor UO_1121 (O_1121,N_24814,N_24765);
nand UO_1122 (O_1122,N_24788,N_24882);
nor UO_1123 (O_1123,N_24825,N_24996);
xnor UO_1124 (O_1124,N_24770,N_24954);
and UO_1125 (O_1125,N_24750,N_24903);
xnor UO_1126 (O_1126,N_24773,N_24885);
and UO_1127 (O_1127,N_24999,N_24853);
or UO_1128 (O_1128,N_24750,N_24798);
nor UO_1129 (O_1129,N_24981,N_24799);
or UO_1130 (O_1130,N_24849,N_24759);
nor UO_1131 (O_1131,N_24764,N_24895);
nand UO_1132 (O_1132,N_24772,N_24860);
and UO_1133 (O_1133,N_24770,N_24885);
nand UO_1134 (O_1134,N_24928,N_24868);
xor UO_1135 (O_1135,N_24833,N_24791);
and UO_1136 (O_1136,N_24825,N_24948);
or UO_1137 (O_1137,N_24979,N_24966);
or UO_1138 (O_1138,N_24980,N_24966);
or UO_1139 (O_1139,N_24927,N_24861);
and UO_1140 (O_1140,N_24840,N_24822);
and UO_1141 (O_1141,N_24841,N_24966);
and UO_1142 (O_1142,N_24826,N_24949);
nand UO_1143 (O_1143,N_24813,N_24823);
nand UO_1144 (O_1144,N_24767,N_24810);
nor UO_1145 (O_1145,N_24875,N_24761);
nor UO_1146 (O_1146,N_24962,N_24983);
or UO_1147 (O_1147,N_24893,N_24764);
xnor UO_1148 (O_1148,N_24787,N_24916);
xnor UO_1149 (O_1149,N_24988,N_24750);
nand UO_1150 (O_1150,N_24868,N_24826);
nor UO_1151 (O_1151,N_24981,N_24759);
xor UO_1152 (O_1152,N_24795,N_24956);
or UO_1153 (O_1153,N_24911,N_24892);
and UO_1154 (O_1154,N_24790,N_24756);
nor UO_1155 (O_1155,N_24912,N_24864);
nand UO_1156 (O_1156,N_24819,N_24753);
or UO_1157 (O_1157,N_24983,N_24989);
nand UO_1158 (O_1158,N_24971,N_24877);
nand UO_1159 (O_1159,N_24999,N_24845);
nor UO_1160 (O_1160,N_24913,N_24874);
nor UO_1161 (O_1161,N_24793,N_24902);
or UO_1162 (O_1162,N_24966,N_24874);
nand UO_1163 (O_1163,N_24994,N_24905);
xor UO_1164 (O_1164,N_24849,N_24937);
and UO_1165 (O_1165,N_24985,N_24992);
or UO_1166 (O_1166,N_24801,N_24773);
or UO_1167 (O_1167,N_24884,N_24995);
or UO_1168 (O_1168,N_24864,N_24969);
nand UO_1169 (O_1169,N_24762,N_24893);
nand UO_1170 (O_1170,N_24916,N_24834);
or UO_1171 (O_1171,N_24802,N_24818);
and UO_1172 (O_1172,N_24883,N_24995);
xor UO_1173 (O_1173,N_24914,N_24763);
nor UO_1174 (O_1174,N_24802,N_24938);
or UO_1175 (O_1175,N_24857,N_24907);
and UO_1176 (O_1176,N_24871,N_24798);
nand UO_1177 (O_1177,N_24983,N_24776);
or UO_1178 (O_1178,N_24942,N_24907);
xnor UO_1179 (O_1179,N_24833,N_24912);
nor UO_1180 (O_1180,N_24943,N_24768);
or UO_1181 (O_1181,N_24942,N_24761);
nor UO_1182 (O_1182,N_24780,N_24940);
nand UO_1183 (O_1183,N_24777,N_24942);
nor UO_1184 (O_1184,N_24918,N_24975);
nand UO_1185 (O_1185,N_24804,N_24890);
xor UO_1186 (O_1186,N_24788,N_24773);
nand UO_1187 (O_1187,N_24764,N_24925);
nand UO_1188 (O_1188,N_24760,N_24780);
nand UO_1189 (O_1189,N_24818,N_24905);
xor UO_1190 (O_1190,N_24906,N_24920);
nor UO_1191 (O_1191,N_24929,N_24833);
and UO_1192 (O_1192,N_24952,N_24805);
xor UO_1193 (O_1193,N_24886,N_24795);
nor UO_1194 (O_1194,N_24912,N_24761);
or UO_1195 (O_1195,N_24992,N_24796);
or UO_1196 (O_1196,N_24819,N_24812);
xnor UO_1197 (O_1197,N_24780,N_24890);
nor UO_1198 (O_1198,N_24832,N_24911);
and UO_1199 (O_1199,N_24800,N_24999);
nand UO_1200 (O_1200,N_24888,N_24933);
nand UO_1201 (O_1201,N_24765,N_24781);
and UO_1202 (O_1202,N_24818,N_24769);
nand UO_1203 (O_1203,N_24893,N_24789);
nand UO_1204 (O_1204,N_24836,N_24762);
nand UO_1205 (O_1205,N_24926,N_24777);
and UO_1206 (O_1206,N_24864,N_24906);
nor UO_1207 (O_1207,N_24823,N_24936);
nand UO_1208 (O_1208,N_24794,N_24942);
xor UO_1209 (O_1209,N_24817,N_24871);
and UO_1210 (O_1210,N_24803,N_24879);
and UO_1211 (O_1211,N_24856,N_24775);
xor UO_1212 (O_1212,N_24819,N_24798);
or UO_1213 (O_1213,N_24973,N_24772);
or UO_1214 (O_1214,N_24799,N_24935);
nand UO_1215 (O_1215,N_24918,N_24986);
nand UO_1216 (O_1216,N_24842,N_24807);
or UO_1217 (O_1217,N_24993,N_24874);
nand UO_1218 (O_1218,N_24820,N_24970);
and UO_1219 (O_1219,N_24913,N_24919);
and UO_1220 (O_1220,N_24957,N_24985);
nor UO_1221 (O_1221,N_24772,N_24872);
nand UO_1222 (O_1222,N_24784,N_24778);
nor UO_1223 (O_1223,N_24824,N_24858);
nor UO_1224 (O_1224,N_24929,N_24891);
or UO_1225 (O_1225,N_24999,N_24792);
nand UO_1226 (O_1226,N_24890,N_24838);
or UO_1227 (O_1227,N_24773,N_24961);
nor UO_1228 (O_1228,N_24883,N_24759);
or UO_1229 (O_1229,N_24892,N_24927);
nor UO_1230 (O_1230,N_24910,N_24781);
and UO_1231 (O_1231,N_24981,N_24915);
nand UO_1232 (O_1232,N_24902,N_24864);
xor UO_1233 (O_1233,N_24949,N_24954);
xor UO_1234 (O_1234,N_24820,N_24937);
xnor UO_1235 (O_1235,N_24889,N_24930);
nor UO_1236 (O_1236,N_24936,N_24813);
or UO_1237 (O_1237,N_24804,N_24790);
nor UO_1238 (O_1238,N_24910,N_24773);
or UO_1239 (O_1239,N_24835,N_24889);
nand UO_1240 (O_1240,N_24868,N_24870);
and UO_1241 (O_1241,N_24793,N_24965);
nor UO_1242 (O_1242,N_24895,N_24981);
and UO_1243 (O_1243,N_24816,N_24894);
nand UO_1244 (O_1244,N_24990,N_24930);
nand UO_1245 (O_1245,N_24886,N_24851);
nand UO_1246 (O_1246,N_24820,N_24907);
and UO_1247 (O_1247,N_24913,N_24976);
nor UO_1248 (O_1248,N_24919,N_24979);
xor UO_1249 (O_1249,N_24828,N_24811);
or UO_1250 (O_1250,N_24851,N_24880);
and UO_1251 (O_1251,N_24988,N_24782);
or UO_1252 (O_1252,N_24759,N_24768);
nand UO_1253 (O_1253,N_24771,N_24954);
nor UO_1254 (O_1254,N_24907,N_24987);
nor UO_1255 (O_1255,N_24790,N_24836);
nor UO_1256 (O_1256,N_24994,N_24966);
nor UO_1257 (O_1257,N_24923,N_24807);
nor UO_1258 (O_1258,N_24863,N_24833);
and UO_1259 (O_1259,N_24969,N_24886);
or UO_1260 (O_1260,N_24892,N_24918);
or UO_1261 (O_1261,N_24946,N_24957);
xnor UO_1262 (O_1262,N_24777,N_24795);
or UO_1263 (O_1263,N_24825,N_24965);
nand UO_1264 (O_1264,N_24839,N_24855);
nor UO_1265 (O_1265,N_24805,N_24997);
xnor UO_1266 (O_1266,N_24978,N_24902);
nand UO_1267 (O_1267,N_24928,N_24851);
nor UO_1268 (O_1268,N_24980,N_24792);
xor UO_1269 (O_1269,N_24760,N_24955);
nand UO_1270 (O_1270,N_24837,N_24964);
nor UO_1271 (O_1271,N_24755,N_24810);
or UO_1272 (O_1272,N_24887,N_24875);
or UO_1273 (O_1273,N_24887,N_24934);
nor UO_1274 (O_1274,N_24969,N_24882);
nand UO_1275 (O_1275,N_24930,N_24823);
nor UO_1276 (O_1276,N_24843,N_24775);
nand UO_1277 (O_1277,N_24872,N_24988);
nand UO_1278 (O_1278,N_24780,N_24896);
nand UO_1279 (O_1279,N_24993,N_24763);
and UO_1280 (O_1280,N_24819,N_24913);
or UO_1281 (O_1281,N_24839,N_24840);
nand UO_1282 (O_1282,N_24829,N_24932);
nand UO_1283 (O_1283,N_24755,N_24771);
nor UO_1284 (O_1284,N_24978,N_24999);
xor UO_1285 (O_1285,N_24991,N_24860);
nor UO_1286 (O_1286,N_24997,N_24932);
and UO_1287 (O_1287,N_24995,N_24864);
xor UO_1288 (O_1288,N_24952,N_24887);
or UO_1289 (O_1289,N_24766,N_24790);
nor UO_1290 (O_1290,N_24775,N_24898);
and UO_1291 (O_1291,N_24953,N_24803);
and UO_1292 (O_1292,N_24795,N_24905);
or UO_1293 (O_1293,N_24993,N_24916);
and UO_1294 (O_1294,N_24755,N_24993);
xnor UO_1295 (O_1295,N_24806,N_24915);
xnor UO_1296 (O_1296,N_24752,N_24853);
nor UO_1297 (O_1297,N_24769,N_24919);
and UO_1298 (O_1298,N_24753,N_24912);
xor UO_1299 (O_1299,N_24795,N_24898);
nor UO_1300 (O_1300,N_24764,N_24923);
xnor UO_1301 (O_1301,N_24890,N_24849);
and UO_1302 (O_1302,N_24950,N_24816);
nor UO_1303 (O_1303,N_24977,N_24850);
or UO_1304 (O_1304,N_24969,N_24972);
nand UO_1305 (O_1305,N_24796,N_24803);
xnor UO_1306 (O_1306,N_24999,N_24911);
nand UO_1307 (O_1307,N_24813,N_24875);
and UO_1308 (O_1308,N_24967,N_24811);
nand UO_1309 (O_1309,N_24952,N_24794);
nor UO_1310 (O_1310,N_24859,N_24939);
or UO_1311 (O_1311,N_24997,N_24935);
or UO_1312 (O_1312,N_24900,N_24789);
nand UO_1313 (O_1313,N_24939,N_24815);
nand UO_1314 (O_1314,N_24804,N_24776);
or UO_1315 (O_1315,N_24844,N_24789);
xnor UO_1316 (O_1316,N_24958,N_24787);
nand UO_1317 (O_1317,N_24765,N_24932);
nand UO_1318 (O_1318,N_24927,N_24847);
nand UO_1319 (O_1319,N_24761,N_24856);
xor UO_1320 (O_1320,N_24986,N_24751);
xor UO_1321 (O_1321,N_24799,N_24857);
or UO_1322 (O_1322,N_24823,N_24918);
nand UO_1323 (O_1323,N_24803,N_24951);
and UO_1324 (O_1324,N_24971,N_24988);
or UO_1325 (O_1325,N_24780,N_24970);
nand UO_1326 (O_1326,N_24992,N_24903);
nand UO_1327 (O_1327,N_24757,N_24855);
nand UO_1328 (O_1328,N_24941,N_24782);
xnor UO_1329 (O_1329,N_24823,N_24992);
nor UO_1330 (O_1330,N_24913,N_24788);
nor UO_1331 (O_1331,N_24776,N_24934);
xnor UO_1332 (O_1332,N_24897,N_24958);
xor UO_1333 (O_1333,N_24885,N_24943);
nor UO_1334 (O_1334,N_24903,N_24945);
nand UO_1335 (O_1335,N_24783,N_24762);
nor UO_1336 (O_1336,N_24869,N_24750);
or UO_1337 (O_1337,N_24824,N_24850);
nor UO_1338 (O_1338,N_24757,N_24973);
nor UO_1339 (O_1339,N_24776,N_24953);
or UO_1340 (O_1340,N_24958,N_24873);
nor UO_1341 (O_1341,N_24865,N_24995);
xnor UO_1342 (O_1342,N_24787,N_24759);
xor UO_1343 (O_1343,N_24766,N_24998);
or UO_1344 (O_1344,N_24986,N_24887);
nand UO_1345 (O_1345,N_24982,N_24947);
and UO_1346 (O_1346,N_24775,N_24771);
xnor UO_1347 (O_1347,N_24849,N_24801);
nor UO_1348 (O_1348,N_24818,N_24890);
and UO_1349 (O_1349,N_24913,N_24820);
or UO_1350 (O_1350,N_24894,N_24988);
xor UO_1351 (O_1351,N_24802,N_24814);
and UO_1352 (O_1352,N_24875,N_24931);
nand UO_1353 (O_1353,N_24771,N_24797);
nor UO_1354 (O_1354,N_24996,N_24821);
and UO_1355 (O_1355,N_24986,N_24936);
nand UO_1356 (O_1356,N_24876,N_24980);
nand UO_1357 (O_1357,N_24914,N_24860);
and UO_1358 (O_1358,N_24910,N_24856);
and UO_1359 (O_1359,N_24815,N_24907);
nand UO_1360 (O_1360,N_24831,N_24945);
nand UO_1361 (O_1361,N_24785,N_24928);
nor UO_1362 (O_1362,N_24906,N_24870);
nor UO_1363 (O_1363,N_24931,N_24943);
nand UO_1364 (O_1364,N_24957,N_24924);
nor UO_1365 (O_1365,N_24820,N_24864);
nand UO_1366 (O_1366,N_24769,N_24762);
and UO_1367 (O_1367,N_24782,N_24949);
nand UO_1368 (O_1368,N_24872,N_24933);
nand UO_1369 (O_1369,N_24871,N_24952);
or UO_1370 (O_1370,N_24901,N_24795);
nor UO_1371 (O_1371,N_24887,N_24751);
nor UO_1372 (O_1372,N_24861,N_24903);
nor UO_1373 (O_1373,N_24921,N_24942);
or UO_1374 (O_1374,N_24751,N_24976);
nand UO_1375 (O_1375,N_24928,N_24768);
or UO_1376 (O_1376,N_24794,N_24996);
nand UO_1377 (O_1377,N_24941,N_24848);
or UO_1378 (O_1378,N_24803,N_24766);
and UO_1379 (O_1379,N_24901,N_24924);
nand UO_1380 (O_1380,N_24860,N_24824);
xor UO_1381 (O_1381,N_24917,N_24854);
or UO_1382 (O_1382,N_24824,N_24951);
and UO_1383 (O_1383,N_24967,N_24825);
nor UO_1384 (O_1384,N_24760,N_24937);
and UO_1385 (O_1385,N_24754,N_24982);
nand UO_1386 (O_1386,N_24991,N_24776);
nand UO_1387 (O_1387,N_24813,N_24994);
nand UO_1388 (O_1388,N_24851,N_24797);
nand UO_1389 (O_1389,N_24924,N_24938);
and UO_1390 (O_1390,N_24854,N_24846);
and UO_1391 (O_1391,N_24833,N_24881);
nand UO_1392 (O_1392,N_24907,N_24778);
or UO_1393 (O_1393,N_24900,N_24833);
nor UO_1394 (O_1394,N_24899,N_24979);
nand UO_1395 (O_1395,N_24836,N_24948);
nand UO_1396 (O_1396,N_24972,N_24986);
and UO_1397 (O_1397,N_24951,N_24925);
nand UO_1398 (O_1398,N_24890,N_24946);
and UO_1399 (O_1399,N_24974,N_24842);
nor UO_1400 (O_1400,N_24955,N_24953);
nand UO_1401 (O_1401,N_24796,N_24947);
nor UO_1402 (O_1402,N_24842,N_24788);
nand UO_1403 (O_1403,N_24786,N_24987);
or UO_1404 (O_1404,N_24995,N_24767);
nand UO_1405 (O_1405,N_24837,N_24764);
and UO_1406 (O_1406,N_24822,N_24786);
xnor UO_1407 (O_1407,N_24976,N_24919);
nand UO_1408 (O_1408,N_24834,N_24969);
xnor UO_1409 (O_1409,N_24903,N_24954);
nand UO_1410 (O_1410,N_24861,N_24852);
nand UO_1411 (O_1411,N_24921,N_24815);
xor UO_1412 (O_1412,N_24873,N_24831);
nor UO_1413 (O_1413,N_24802,N_24956);
nand UO_1414 (O_1414,N_24938,N_24904);
xnor UO_1415 (O_1415,N_24804,N_24996);
xor UO_1416 (O_1416,N_24842,N_24810);
nand UO_1417 (O_1417,N_24943,N_24921);
nor UO_1418 (O_1418,N_24926,N_24875);
and UO_1419 (O_1419,N_24844,N_24992);
or UO_1420 (O_1420,N_24882,N_24795);
xnor UO_1421 (O_1421,N_24830,N_24798);
xnor UO_1422 (O_1422,N_24845,N_24810);
xor UO_1423 (O_1423,N_24815,N_24803);
or UO_1424 (O_1424,N_24815,N_24974);
nand UO_1425 (O_1425,N_24926,N_24759);
xor UO_1426 (O_1426,N_24981,N_24868);
xor UO_1427 (O_1427,N_24952,N_24779);
or UO_1428 (O_1428,N_24839,N_24963);
or UO_1429 (O_1429,N_24950,N_24757);
and UO_1430 (O_1430,N_24879,N_24942);
and UO_1431 (O_1431,N_24755,N_24989);
nor UO_1432 (O_1432,N_24776,N_24928);
nand UO_1433 (O_1433,N_24910,N_24851);
xnor UO_1434 (O_1434,N_24941,N_24787);
xnor UO_1435 (O_1435,N_24804,N_24879);
xnor UO_1436 (O_1436,N_24968,N_24867);
xor UO_1437 (O_1437,N_24901,N_24865);
and UO_1438 (O_1438,N_24952,N_24925);
and UO_1439 (O_1439,N_24791,N_24785);
and UO_1440 (O_1440,N_24897,N_24828);
or UO_1441 (O_1441,N_24942,N_24896);
nand UO_1442 (O_1442,N_24968,N_24964);
nor UO_1443 (O_1443,N_24843,N_24851);
or UO_1444 (O_1444,N_24767,N_24864);
nand UO_1445 (O_1445,N_24838,N_24828);
nor UO_1446 (O_1446,N_24802,N_24890);
nor UO_1447 (O_1447,N_24911,N_24869);
nand UO_1448 (O_1448,N_24894,N_24892);
and UO_1449 (O_1449,N_24849,N_24891);
nor UO_1450 (O_1450,N_24917,N_24763);
and UO_1451 (O_1451,N_24766,N_24825);
and UO_1452 (O_1452,N_24999,N_24816);
and UO_1453 (O_1453,N_24780,N_24768);
or UO_1454 (O_1454,N_24846,N_24824);
or UO_1455 (O_1455,N_24986,N_24755);
nor UO_1456 (O_1456,N_24963,N_24941);
xnor UO_1457 (O_1457,N_24821,N_24965);
or UO_1458 (O_1458,N_24988,N_24871);
and UO_1459 (O_1459,N_24773,N_24769);
nor UO_1460 (O_1460,N_24989,N_24984);
nand UO_1461 (O_1461,N_24788,N_24879);
or UO_1462 (O_1462,N_24984,N_24956);
or UO_1463 (O_1463,N_24914,N_24769);
and UO_1464 (O_1464,N_24943,N_24769);
nor UO_1465 (O_1465,N_24868,N_24779);
or UO_1466 (O_1466,N_24919,N_24833);
or UO_1467 (O_1467,N_24881,N_24781);
or UO_1468 (O_1468,N_24842,N_24906);
xor UO_1469 (O_1469,N_24763,N_24839);
nor UO_1470 (O_1470,N_24962,N_24939);
nand UO_1471 (O_1471,N_24973,N_24807);
nand UO_1472 (O_1472,N_24871,N_24950);
and UO_1473 (O_1473,N_24760,N_24810);
xor UO_1474 (O_1474,N_24801,N_24925);
xor UO_1475 (O_1475,N_24761,N_24962);
nand UO_1476 (O_1476,N_24826,N_24898);
nor UO_1477 (O_1477,N_24783,N_24827);
xnor UO_1478 (O_1478,N_24832,N_24872);
or UO_1479 (O_1479,N_24875,N_24865);
nor UO_1480 (O_1480,N_24751,N_24842);
and UO_1481 (O_1481,N_24952,N_24899);
and UO_1482 (O_1482,N_24992,N_24982);
nor UO_1483 (O_1483,N_24986,N_24862);
and UO_1484 (O_1484,N_24969,N_24819);
nand UO_1485 (O_1485,N_24896,N_24864);
xor UO_1486 (O_1486,N_24886,N_24899);
and UO_1487 (O_1487,N_24879,N_24793);
or UO_1488 (O_1488,N_24829,N_24870);
xor UO_1489 (O_1489,N_24915,N_24921);
or UO_1490 (O_1490,N_24828,N_24809);
nand UO_1491 (O_1491,N_24854,N_24997);
nand UO_1492 (O_1492,N_24863,N_24898);
and UO_1493 (O_1493,N_24786,N_24916);
nand UO_1494 (O_1494,N_24816,N_24910);
xnor UO_1495 (O_1495,N_24942,N_24904);
xor UO_1496 (O_1496,N_24755,N_24908);
and UO_1497 (O_1497,N_24991,N_24935);
or UO_1498 (O_1498,N_24939,N_24882);
nand UO_1499 (O_1499,N_24864,N_24849);
and UO_1500 (O_1500,N_24807,N_24879);
nand UO_1501 (O_1501,N_24825,N_24997);
xor UO_1502 (O_1502,N_24802,N_24935);
or UO_1503 (O_1503,N_24779,N_24824);
xor UO_1504 (O_1504,N_24781,N_24974);
xnor UO_1505 (O_1505,N_24922,N_24923);
or UO_1506 (O_1506,N_24848,N_24865);
nor UO_1507 (O_1507,N_24799,N_24995);
or UO_1508 (O_1508,N_24979,N_24934);
nand UO_1509 (O_1509,N_24981,N_24969);
nand UO_1510 (O_1510,N_24818,N_24992);
and UO_1511 (O_1511,N_24923,N_24816);
nand UO_1512 (O_1512,N_24815,N_24972);
nor UO_1513 (O_1513,N_24854,N_24840);
nand UO_1514 (O_1514,N_24801,N_24944);
and UO_1515 (O_1515,N_24945,N_24943);
and UO_1516 (O_1516,N_24808,N_24822);
or UO_1517 (O_1517,N_24778,N_24921);
and UO_1518 (O_1518,N_24989,N_24864);
or UO_1519 (O_1519,N_24832,N_24752);
or UO_1520 (O_1520,N_24806,N_24982);
nand UO_1521 (O_1521,N_24940,N_24919);
nand UO_1522 (O_1522,N_24925,N_24816);
and UO_1523 (O_1523,N_24825,N_24772);
or UO_1524 (O_1524,N_24831,N_24771);
nand UO_1525 (O_1525,N_24816,N_24871);
and UO_1526 (O_1526,N_24793,N_24909);
nor UO_1527 (O_1527,N_24983,N_24875);
xnor UO_1528 (O_1528,N_24964,N_24802);
or UO_1529 (O_1529,N_24969,N_24962);
xnor UO_1530 (O_1530,N_24774,N_24845);
or UO_1531 (O_1531,N_24953,N_24948);
or UO_1532 (O_1532,N_24930,N_24934);
xnor UO_1533 (O_1533,N_24899,N_24940);
xnor UO_1534 (O_1534,N_24949,N_24850);
nor UO_1535 (O_1535,N_24784,N_24934);
or UO_1536 (O_1536,N_24917,N_24798);
or UO_1537 (O_1537,N_24783,N_24818);
xnor UO_1538 (O_1538,N_24947,N_24808);
nand UO_1539 (O_1539,N_24977,N_24892);
or UO_1540 (O_1540,N_24754,N_24758);
and UO_1541 (O_1541,N_24764,N_24779);
xnor UO_1542 (O_1542,N_24840,N_24888);
nor UO_1543 (O_1543,N_24914,N_24754);
xor UO_1544 (O_1544,N_24871,N_24858);
or UO_1545 (O_1545,N_24765,N_24788);
nand UO_1546 (O_1546,N_24775,N_24857);
xor UO_1547 (O_1547,N_24884,N_24772);
nand UO_1548 (O_1548,N_24917,N_24755);
nand UO_1549 (O_1549,N_24864,N_24894);
or UO_1550 (O_1550,N_24904,N_24959);
nor UO_1551 (O_1551,N_24850,N_24939);
and UO_1552 (O_1552,N_24816,N_24814);
nor UO_1553 (O_1553,N_24926,N_24755);
nor UO_1554 (O_1554,N_24894,N_24782);
nor UO_1555 (O_1555,N_24981,N_24931);
nand UO_1556 (O_1556,N_24798,N_24949);
nand UO_1557 (O_1557,N_24893,N_24905);
xor UO_1558 (O_1558,N_24848,N_24810);
nand UO_1559 (O_1559,N_24917,N_24914);
xor UO_1560 (O_1560,N_24926,N_24851);
nand UO_1561 (O_1561,N_24889,N_24901);
nand UO_1562 (O_1562,N_24786,N_24979);
and UO_1563 (O_1563,N_24783,N_24833);
nor UO_1564 (O_1564,N_24815,N_24845);
xnor UO_1565 (O_1565,N_24967,N_24955);
xnor UO_1566 (O_1566,N_24768,N_24907);
and UO_1567 (O_1567,N_24869,N_24925);
nor UO_1568 (O_1568,N_24904,N_24914);
xnor UO_1569 (O_1569,N_24778,N_24910);
or UO_1570 (O_1570,N_24867,N_24862);
or UO_1571 (O_1571,N_24766,N_24884);
and UO_1572 (O_1572,N_24752,N_24906);
nor UO_1573 (O_1573,N_24829,N_24764);
nor UO_1574 (O_1574,N_24816,N_24926);
nor UO_1575 (O_1575,N_24896,N_24956);
nor UO_1576 (O_1576,N_24768,N_24859);
nor UO_1577 (O_1577,N_24996,N_24791);
xor UO_1578 (O_1578,N_24771,N_24919);
and UO_1579 (O_1579,N_24963,N_24853);
or UO_1580 (O_1580,N_24954,N_24907);
nand UO_1581 (O_1581,N_24979,N_24959);
nor UO_1582 (O_1582,N_24892,N_24828);
nand UO_1583 (O_1583,N_24778,N_24860);
nand UO_1584 (O_1584,N_24969,N_24955);
nor UO_1585 (O_1585,N_24850,N_24801);
or UO_1586 (O_1586,N_24941,N_24872);
nand UO_1587 (O_1587,N_24867,N_24995);
and UO_1588 (O_1588,N_24757,N_24785);
or UO_1589 (O_1589,N_24768,N_24999);
nand UO_1590 (O_1590,N_24822,N_24941);
and UO_1591 (O_1591,N_24892,N_24785);
nor UO_1592 (O_1592,N_24863,N_24995);
nand UO_1593 (O_1593,N_24904,N_24975);
and UO_1594 (O_1594,N_24917,N_24926);
and UO_1595 (O_1595,N_24770,N_24849);
or UO_1596 (O_1596,N_24808,N_24793);
xnor UO_1597 (O_1597,N_24833,N_24763);
and UO_1598 (O_1598,N_24935,N_24998);
nor UO_1599 (O_1599,N_24951,N_24802);
nor UO_1600 (O_1600,N_24827,N_24880);
and UO_1601 (O_1601,N_24811,N_24977);
or UO_1602 (O_1602,N_24832,N_24817);
nor UO_1603 (O_1603,N_24781,N_24785);
and UO_1604 (O_1604,N_24986,N_24805);
and UO_1605 (O_1605,N_24761,N_24932);
and UO_1606 (O_1606,N_24785,N_24952);
or UO_1607 (O_1607,N_24756,N_24905);
nor UO_1608 (O_1608,N_24931,N_24993);
or UO_1609 (O_1609,N_24960,N_24986);
nor UO_1610 (O_1610,N_24877,N_24807);
or UO_1611 (O_1611,N_24889,N_24866);
nand UO_1612 (O_1612,N_24966,N_24754);
and UO_1613 (O_1613,N_24918,N_24951);
xnor UO_1614 (O_1614,N_24924,N_24967);
xor UO_1615 (O_1615,N_24982,N_24750);
and UO_1616 (O_1616,N_24949,N_24852);
nor UO_1617 (O_1617,N_24937,N_24759);
nor UO_1618 (O_1618,N_24907,N_24935);
nand UO_1619 (O_1619,N_24876,N_24820);
nand UO_1620 (O_1620,N_24908,N_24963);
xnor UO_1621 (O_1621,N_24870,N_24876);
and UO_1622 (O_1622,N_24822,N_24867);
and UO_1623 (O_1623,N_24975,N_24814);
or UO_1624 (O_1624,N_24959,N_24913);
nor UO_1625 (O_1625,N_24968,N_24996);
nand UO_1626 (O_1626,N_24826,N_24973);
xnor UO_1627 (O_1627,N_24957,N_24808);
nor UO_1628 (O_1628,N_24778,N_24944);
nor UO_1629 (O_1629,N_24987,N_24885);
or UO_1630 (O_1630,N_24953,N_24809);
nand UO_1631 (O_1631,N_24916,N_24919);
xnor UO_1632 (O_1632,N_24890,N_24793);
nor UO_1633 (O_1633,N_24759,N_24881);
nand UO_1634 (O_1634,N_24766,N_24972);
nand UO_1635 (O_1635,N_24750,N_24968);
nor UO_1636 (O_1636,N_24964,N_24846);
nand UO_1637 (O_1637,N_24876,N_24807);
nand UO_1638 (O_1638,N_24850,N_24952);
nand UO_1639 (O_1639,N_24817,N_24894);
or UO_1640 (O_1640,N_24988,N_24777);
and UO_1641 (O_1641,N_24925,N_24931);
nor UO_1642 (O_1642,N_24948,N_24910);
xnor UO_1643 (O_1643,N_24932,N_24986);
nor UO_1644 (O_1644,N_24757,N_24755);
nor UO_1645 (O_1645,N_24778,N_24836);
or UO_1646 (O_1646,N_24887,N_24901);
nand UO_1647 (O_1647,N_24857,N_24984);
nor UO_1648 (O_1648,N_24845,N_24998);
or UO_1649 (O_1649,N_24999,N_24997);
xor UO_1650 (O_1650,N_24933,N_24831);
or UO_1651 (O_1651,N_24755,N_24956);
and UO_1652 (O_1652,N_24829,N_24971);
xnor UO_1653 (O_1653,N_24782,N_24967);
nand UO_1654 (O_1654,N_24797,N_24969);
xnor UO_1655 (O_1655,N_24837,N_24844);
and UO_1656 (O_1656,N_24973,N_24863);
and UO_1657 (O_1657,N_24875,N_24980);
and UO_1658 (O_1658,N_24999,N_24884);
xor UO_1659 (O_1659,N_24999,N_24780);
and UO_1660 (O_1660,N_24793,N_24917);
or UO_1661 (O_1661,N_24816,N_24935);
or UO_1662 (O_1662,N_24990,N_24792);
xor UO_1663 (O_1663,N_24911,N_24916);
nand UO_1664 (O_1664,N_24951,N_24913);
and UO_1665 (O_1665,N_24991,N_24800);
nand UO_1666 (O_1666,N_24782,N_24834);
or UO_1667 (O_1667,N_24821,N_24928);
and UO_1668 (O_1668,N_24932,N_24797);
nand UO_1669 (O_1669,N_24966,N_24821);
nand UO_1670 (O_1670,N_24757,N_24776);
nand UO_1671 (O_1671,N_24866,N_24804);
nand UO_1672 (O_1672,N_24810,N_24855);
and UO_1673 (O_1673,N_24822,N_24959);
xnor UO_1674 (O_1674,N_24819,N_24911);
nand UO_1675 (O_1675,N_24780,N_24878);
nor UO_1676 (O_1676,N_24995,N_24958);
and UO_1677 (O_1677,N_24812,N_24859);
nand UO_1678 (O_1678,N_24972,N_24897);
or UO_1679 (O_1679,N_24894,N_24885);
nor UO_1680 (O_1680,N_24769,N_24973);
or UO_1681 (O_1681,N_24846,N_24774);
nor UO_1682 (O_1682,N_24836,N_24759);
and UO_1683 (O_1683,N_24849,N_24804);
and UO_1684 (O_1684,N_24844,N_24922);
nor UO_1685 (O_1685,N_24865,N_24762);
xor UO_1686 (O_1686,N_24825,N_24908);
nand UO_1687 (O_1687,N_24893,N_24886);
or UO_1688 (O_1688,N_24814,N_24922);
nor UO_1689 (O_1689,N_24996,N_24943);
nor UO_1690 (O_1690,N_24763,N_24783);
nor UO_1691 (O_1691,N_24857,N_24979);
or UO_1692 (O_1692,N_24887,N_24808);
and UO_1693 (O_1693,N_24975,N_24896);
xnor UO_1694 (O_1694,N_24772,N_24945);
and UO_1695 (O_1695,N_24922,N_24898);
nor UO_1696 (O_1696,N_24990,N_24987);
nand UO_1697 (O_1697,N_24764,N_24993);
xor UO_1698 (O_1698,N_24857,N_24793);
nor UO_1699 (O_1699,N_24864,N_24987);
nand UO_1700 (O_1700,N_24982,N_24988);
and UO_1701 (O_1701,N_24953,N_24999);
xnor UO_1702 (O_1702,N_24932,N_24845);
nand UO_1703 (O_1703,N_24798,N_24980);
and UO_1704 (O_1704,N_24975,N_24947);
xor UO_1705 (O_1705,N_24988,N_24808);
nor UO_1706 (O_1706,N_24789,N_24988);
xnor UO_1707 (O_1707,N_24935,N_24755);
and UO_1708 (O_1708,N_24856,N_24971);
and UO_1709 (O_1709,N_24885,N_24808);
nand UO_1710 (O_1710,N_24974,N_24892);
nor UO_1711 (O_1711,N_24825,N_24883);
nor UO_1712 (O_1712,N_24861,N_24935);
xnor UO_1713 (O_1713,N_24752,N_24790);
or UO_1714 (O_1714,N_24879,N_24820);
and UO_1715 (O_1715,N_24840,N_24927);
nand UO_1716 (O_1716,N_24829,N_24832);
xnor UO_1717 (O_1717,N_24773,N_24765);
nand UO_1718 (O_1718,N_24933,N_24832);
or UO_1719 (O_1719,N_24942,N_24933);
and UO_1720 (O_1720,N_24993,N_24849);
xnor UO_1721 (O_1721,N_24788,N_24871);
nand UO_1722 (O_1722,N_24872,N_24810);
xnor UO_1723 (O_1723,N_24803,N_24848);
or UO_1724 (O_1724,N_24841,N_24984);
nand UO_1725 (O_1725,N_24793,N_24765);
xor UO_1726 (O_1726,N_24771,N_24791);
nor UO_1727 (O_1727,N_24791,N_24812);
nand UO_1728 (O_1728,N_24940,N_24777);
or UO_1729 (O_1729,N_24889,N_24968);
nand UO_1730 (O_1730,N_24940,N_24790);
nor UO_1731 (O_1731,N_24880,N_24896);
nor UO_1732 (O_1732,N_24776,N_24784);
and UO_1733 (O_1733,N_24767,N_24753);
or UO_1734 (O_1734,N_24834,N_24847);
or UO_1735 (O_1735,N_24776,N_24841);
nor UO_1736 (O_1736,N_24941,N_24943);
or UO_1737 (O_1737,N_24902,N_24832);
nand UO_1738 (O_1738,N_24878,N_24986);
or UO_1739 (O_1739,N_24821,N_24765);
or UO_1740 (O_1740,N_24912,N_24985);
nor UO_1741 (O_1741,N_24805,N_24814);
nand UO_1742 (O_1742,N_24807,N_24902);
and UO_1743 (O_1743,N_24891,N_24900);
xnor UO_1744 (O_1744,N_24822,N_24915);
nor UO_1745 (O_1745,N_24980,N_24845);
nand UO_1746 (O_1746,N_24979,N_24898);
nand UO_1747 (O_1747,N_24911,N_24957);
or UO_1748 (O_1748,N_24882,N_24871);
and UO_1749 (O_1749,N_24796,N_24776);
or UO_1750 (O_1750,N_24793,N_24810);
nor UO_1751 (O_1751,N_24905,N_24991);
nand UO_1752 (O_1752,N_24918,N_24828);
nand UO_1753 (O_1753,N_24792,N_24797);
nor UO_1754 (O_1754,N_24802,N_24838);
and UO_1755 (O_1755,N_24900,N_24767);
xnor UO_1756 (O_1756,N_24969,N_24874);
xor UO_1757 (O_1757,N_24981,N_24847);
xor UO_1758 (O_1758,N_24849,N_24928);
xor UO_1759 (O_1759,N_24875,N_24838);
xor UO_1760 (O_1760,N_24960,N_24896);
nor UO_1761 (O_1761,N_24917,N_24850);
or UO_1762 (O_1762,N_24968,N_24992);
or UO_1763 (O_1763,N_24877,N_24799);
nor UO_1764 (O_1764,N_24832,N_24848);
or UO_1765 (O_1765,N_24789,N_24904);
or UO_1766 (O_1766,N_24753,N_24774);
nor UO_1767 (O_1767,N_24769,N_24873);
nand UO_1768 (O_1768,N_24901,N_24982);
or UO_1769 (O_1769,N_24845,N_24808);
nor UO_1770 (O_1770,N_24856,N_24813);
and UO_1771 (O_1771,N_24832,N_24965);
or UO_1772 (O_1772,N_24783,N_24913);
or UO_1773 (O_1773,N_24993,N_24971);
nor UO_1774 (O_1774,N_24890,N_24993);
xor UO_1775 (O_1775,N_24981,N_24794);
nor UO_1776 (O_1776,N_24957,N_24931);
nor UO_1777 (O_1777,N_24970,N_24871);
and UO_1778 (O_1778,N_24999,N_24936);
nor UO_1779 (O_1779,N_24891,N_24844);
and UO_1780 (O_1780,N_24840,N_24941);
and UO_1781 (O_1781,N_24855,N_24865);
nor UO_1782 (O_1782,N_24975,N_24837);
nor UO_1783 (O_1783,N_24840,N_24957);
nor UO_1784 (O_1784,N_24949,N_24856);
and UO_1785 (O_1785,N_24952,N_24921);
and UO_1786 (O_1786,N_24935,N_24875);
nor UO_1787 (O_1787,N_24768,N_24986);
and UO_1788 (O_1788,N_24974,N_24869);
or UO_1789 (O_1789,N_24828,N_24925);
nand UO_1790 (O_1790,N_24865,N_24949);
xnor UO_1791 (O_1791,N_24921,N_24841);
nand UO_1792 (O_1792,N_24930,N_24932);
or UO_1793 (O_1793,N_24951,N_24813);
nand UO_1794 (O_1794,N_24802,N_24845);
and UO_1795 (O_1795,N_24854,N_24839);
xnor UO_1796 (O_1796,N_24883,N_24751);
or UO_1797 (O_1797,N_24832,N_24805);
or UO_1798 (O_1798,N_24856,N_24893);
nor UO_1799 (O_1799,N_24854,N_24811);
or UO_1800 (O_1800,N_24851,N_24878);
nand UO_1801 (O_1801,N_24899,N_24997);
and UO_1802 (O_1802,N_24930,N_24778);
or UO_1803 (O_1803,N_24893,N_24883);
nand UO_1804 (O_1804,N_24830,N_24863);
nor UO_1805 (O_1805,N_24871,N_24961);
or UO_1806 (O_1806,N_24965,N_24850);
or UO_1807 (O_1807,N_24767,N_24806);
nand UO_1808 (O_1808,N_24962,N_24753);
xnor UO_1809 (O_1809,N_24936,N_24977);
or UO_1810 (O_1810,N_24903,N_24897);
or UO_1811 (O_1811,N_24827,N_24980);
or UO_1812 (O_1812,N_24863,N_24823);
nand UO_1813 (O_1813,N_24902,N_24752);
nor UO_1814 (O_1814,N_24983,N_24822);
and UO_1815 (O_1815,N_24966,N_24750);
or UO_1816 (O_1816,N_24850,N_24942);
and UO_1817 (O_1817,N_24933,N_24944);
nor UO_1818 (O_1818,N_24940,N_24846);
or UO_1819 (O_1819,N_24805,N_24879);
nor UO_1820 (O_1820,N_24812,N_24809);
or UO_1821 (O_1821,N_24902,N_24788);
nand UO_1822 (O_1822,N_24991,N_24839);
or UO_1823 (O_1823,N_24862,N_24885);
xor UO_1824 (O_1824,N_24942,N_24876);
nand UO_1825 (O_1825,N_24916,N_24987);
nand UO_1826 (O_1826,N_24805,N_24979);
or UO_1827 (O_1827,N_24940,N_24993);
nand UO_1828 (O_1828,N_24982,N_24966);
nor UO_1829 (O_1829,N_24875,N_24964);
nor UO_1830 (O_1830,N_24816,N_24757);
or UO_1831 (O_1831,N_24956,N_24990);
nand UO_1832 (O_1832,N_24822,N_24990);
nand UO_1833 (O_1833,N_24755,N_24853);
or UO_1834 (O_1834,N_24992,N_24973);
xnor UO_1835 (O_1835,N_24754,N_24807);
or UO_1836 (O_1836,N_24975,N_24963);
or UO_1837 (O_1837,N_24924,N_24786);
or UO_1838 (O_1838,N_24798,N_24773);
or UO_1839 (O_1839,N_24942,N_24772);
xnor UO_1840 (O_1840,N_24877,N_24881);
and UO_1841 (O_1841,N_24914,N_24764);
nor UO_1842 (O_1842,N_24764,N_24845);
or UO_1843 (O_1843,N_24851,N_24876);
nand UO_1844 (O_1844,N_24882,N_24947);
nor UO_1845 (O_1845,N_24869,N_24774);
nor UO_1846 (O_1846,N_24783,N_24778);
or UO_1847 (O_1847,N_24762,N_24866);
and UO_1848 (O_1848,N_24768,N_24992);
nor UO_1849 (O_1849,N_24890,N_24824);
nand UO_1850 (O_1850,N_24992,N_24808);
nor UO_1851 (O_1851,N_24954,N_24816);
nor UO_1852 (O_1852,N_24803,N_24987);
or UO_1853 (O_1853,N_24979,N_24817);
nand UO_1854 (O_1854,N_24992,N_24884);
and UO_1855 (O_1855,N_24801,N_24874);
nand UO_1856 (O_1856,N_24788,N_24835);
or UO_1857 (O_1857,N_24865,N_24753);
nand UO_1858 (O_1858,N_24862,N_24795);
xor UO_1859 (O_1859,N_24752,N_24921);
and UO_1860 (O_1860,N_24957,N_24986);
nand UO_1861 (O_1861,N_24963,N_24930);
or UO_1862 (O_1862,N_24768,N_24797);
nor UO_1863 (O_1863,N_24759,N_24955);
or UO_1864 (O_1864,N_24775,N_24810);
xnor UO_1865 (O_1865,N_24953,N_24939);
nor UO_1866 (O_1866,N_24786,N_24891);
and UO_1867 (O_1867,N_24887,N_24813);
nand UO_1868 (O_1868,N_24790,N_24923);
nand UO_1869 (O_1869,N_24988,N_24979);
and UO_1870 (O_1870,N_24817,N_24914);
nand UO_1871 (O_1871,N_24763,N_24894);
xor UO_1872 (O_1872,N_24756,N_24797);
xnor UO_1873 (O_1873,N_24932,N_24764);
nor UO_1874 (O_1874,N_24795,N_24975);
or UO_1875 (O_1875,N_24820,N_24802);
xor UO_1876 (O_1876,N_24905,N_24924);
xnor UO_1877 (O_1877,N_24778,N_24853);
nor UO_1878 (O_1878,N_24867,N_24857);
or UO_1879 (O_1879,N_24906,N_24809);
nand UO_1880 (O_1880,N_24790,N_24758);
or UO_1881 (O_1881,N_24899,N_24968);
nor UO_1882 (O_1882,N_24895,N_24934);
nor UO_1883 (O_1883,N_24909,N_24898);
and UO_1884 (O_1884,N_24797,N_24941);
nor UO_1885 (O_1885,N_24755,N_24977);
xnor UO_1886 (O_1886,N_24869,N_24960);
and UO_1887 (O_1887,N_24982,N_24876);
nand UO_1888 (O_1888,N_24833,N_24975);
or UO_1889 (O_1889,N_24860,N_24846);
xor UO_1890 (O_1890,N_24752,N_24919);
nor UO_1891 (O_1891,N_24970,N_24851);
and UO_1892 (O_1892,N_24771,N_24960);
nand UO_1893 (O_1893,N_24807,N_24786);
and UO_1894 (O_1894,N_24752,N_24774);
xnor UO_1895 (O_1895,N_24790,N_24871);
xnor UO_1896 (O_1896,N_24924,N_24802);
nand UO_1897 (O_1897,N_24914,N_24796);
xor UO_1898 (O_1898,N_24859,N_24892);
xor UO_1899 (O_1899,N_24855,N_24884);
xor UO_1900 (O_1900,N_24891,N_24969);
and UO_1901 (O_1901,N_24874,N_24900);
xor UO_1902 (O_1902,N_24863,N_24750);
or UO_1903 (O_1903,N_24779,N_24873);
nand UO_1904 (O_1904,N_24750,N_24792);
or UO_1905 (O_1905,N_24877,N_24784);
and UO_1906 (O_1906,N_24807,N_24917);
and UO_1907 (O_1907,N_24758,N_24899);
and UO_1908 (O_1908,N_24906,N_24988);
nor UO_1909 (O_1909,N_24903,N_24982);
nor UO_1910 (O_1910,N_24787,N_24975);
nand UO_1911 (O_1911,N_24783,N_24941);
or UO_1912 (O_1912,N_24888,N_24834);
nand UO_1913 (O_1913,N_24872,N_24839);
or UO_1914 (O_1914,N_24989,N_24938);
xor UO_1915 (O_1915,N_24968,N_24822);
nor UO_1916 (O_1916,N_24825,N_24789);
xnor UO_1917 (O_1917,N_24888,N_24867);
xor UO_1918 (O_1918,N_24935,N_24789);
or UO_1919 (O_1919,N_24959,N_24804);
xnor UO_1920 (O_1920,N_24946,N_24810);
xor UO_1921 (O_1921,N_24921,N_24801);
and UO_1922 (O_1922,N_24948,N_24986);
nor UO_1923 (O_1923,N_24779,N_24895);
xnor UO_1924 (O_1924,N_24835,N_24925);
nand UO_1925 (O_1925,N_24863,N_24914);
xor UO_1926 (O_1926,N_24977,N_24799);
or UO_1927 (O_1927,N_24864,N_24774);
xnor UO_1928 (O_1928,N_24957,N_24848);
nand UO_1929 (O_1929,N_24750,N_24882);
and UO_1930 (O_1930,N_24990,N_24895);
xnor UO_1931 (O_1931,N_24809,N_24842);
nor UO_1932 (O_1932,N_24927,N_24917);
nor UO_1933 (O_1933,N_24907,N_24995);
or UO_1934 (O_1934,N_24941,N_24960);
xnor UO_1935 (O_1935,N_24922,N_24915);
nand UO_1936 (O_1936,N_24852,N_24765);
nor UO_1937 (O_1937,N_24778,N_24844);
nor UO_1938 (O_1938,N_24865,N_24898);
or UO_1939 (O_1939,N_24823,N_24987);
nor UO_1940 (O_1940,N_24962,N_24803);
xor UO_1941 (O_1941,N_24937,N_24814);
nand UO_1942 (O_1942,N_24896,N_24944);
xnor UO_1943 (O_1943,N_24792,N_24766);
or UO_1944 (O_1944,N_24964,N_24904);
nand UO_1945 (O_1945,N_24946,N_24911);
or UO_1946 (O_1946,N_24818,N_24966);
xor UO_1947 (O_1947,N_24917,N_24861);
nor UO_1948 (O_1948,N_24934,N_24919);
nand UO_1949 (O_1949,N_24900,N_24964);
xor UO_1950 (O_1950,N_24882,N_24863);
or UO_1951 (O_1951,N_24918,N_24765);
nand UO_1952 (O_1952,N_24990,N_24915);
xnor UO_1953 (O_1953,N_24763,N_24955);
nor UO_1954 (O_1954,N_24993,N_24786);
nand UO_1955 (O_1955,N_24912,N_24879);
or UO_1956 (O_1956,N_24808,N_24752);
and UO_1957 (O_1957,N_24786,N_24792);
and UO_1958 (O_1958,N_24821,N_24987);
nor UO_1959 (O_1959,N_24909,N_24902);
and UO_1960 (O_1960,N_24955,N_24849);
and UO_1961 (O_1961,N_24781,N_24883);
xnor UO_1962 (O_1962,N_24827,N_24801);
nor UO_1963 (O_1963,N_24831,N_24938);
nor UO_1964 (O_1964,N_24873,N_24760);
or UO_1965 (O_1965,N_24982,N_24857);
and UO_1966 (O_1966,N_24814,N_24839);
nand UO_1967 (O_1967,N_24904,N_24819);
nand UO_1968 (O_1968,N_24955,N_24771);
nand UO_1969 (O_1969,N_24856,N_24960);
nor UO_1970 (O_1970,N_24942,N_24768);
or UO_1971 (O_1971,N_24895,N_24871);
nand UO_1972 (O_1972,N_24853,N_24942);
xor UO_1973 (O_1973,N_24876,N_24806);
and UO_1974 (O_1974,N_24980,N_24941);
or UO_1975 (O_1975,N_24819,N_24968);
xor UO_1976 (O_1976,N_24814,N_24773);
or UO_1977 (O_1977,N_24816,N_24802);
and UO_1978 (O_1978,N_24755,N_24872);
xnor UO_1979 (O_1979,N_24958,N_24918);
and UO_1980 (O_1980,N_24909,N_24920);
xor UO_1981 (O_1981,N_24924,N_24953);
nand UO_1982 (O_1982,N_24820,N_24945);
nand UO_1983 (O_1983,N_24762,N_24986);
nor UO_1984 (O_1984,N_24913,N_24868);
nand UO_1985 (O_1985,N_24870,N_24902);
nand UO_1986 (O_1986,N_24806,N_24918);
xor UO_1987 (O_1987,N_24963,N_24772);
nor UO_1988 (O_1988,N_24967,N_24767);
xor UO_1989 (O_1989,N_24968,N_24898);
or UO_1990 (O_1990,N_24906,N_24926);
and UO_1991 (O_1991,N_24757,N_24968);
and UO_1992 (O_1992,N_24854,N_24772);
or UO_1993 (O_1993,N_24883,N_24996);
nor UO_1994 (O_1994,N_24963,N_24958);
or UO_1995 (O_1995,N_24834,N_24901);
nor UO_1996 (O_1996,N_24992,N_24824);
nand UO_1997 (O_1997,N_24847,N_24996);
and UO_1998 (O_1998,N_24913,N_24864);
xnor UO_1999 (O_1999,N_24806,N_24939);
xor UO_2000 (O_2000,N_24926,N_24751);
nor UO_2001 (O_2001,N_24891,N_24827);
or UO_2002 (O_2002,N_24978,N_24758);
or UO_2003 (O_2003,N_24962,N_24935);
nand UO_2004 (O_2004,N_24904,N_24887);
nor UO_2005 (O_2005,N_24924,N_24820);
and UO_2006 (O_2006,N_24777,N_24947);
or UO_2007 (O_2007,N_24803,N_24885);
and UO_2008 (O_2008,N_24840,N_24895);
or UO_2009 (O_2009,N_24991,N_24961);
or UO_2010 (O_2010,N_24849,N_24952);
nand UO_2011 (O_2011,N_24840,N_24804);
or UO_2012 (O_2012,N_24932,N_24865);
or UO_2013 (O_2013,N_24988,N_24991);
nand UO_2014 (O_2014,N_24831,N_24920);
nor UO_2015 (O_2015,N_24898,N_24954);
xnor UO_2016 (O_2016,N_24871,N_24776);
nand UO_2017 (O_2017,N_24817,N_24889);
nor UO_2018 (O_2018,N_24839,N_24944);
nand UO_2019 (O_2019,N_24911,N_24967);
xnor UO_2020 (O_2020,N_24963,N_24959);
xnor UO_2021 (O_2021,N_24887,N_24786);
or UO_2022 (O_2022,N_24835,N_24844);
and UO_2023 (O_2023,N_24897,N_24922);
or UO_2024 (O_2024,N_24989,N_24982);
and UO_2025 (O_2025,N_24990,N_24853);
and UO_2026 (O_2026,N_24835,N_24999);
and UO_2027 (O_2027,N_24911,N_24971);
and UO_2028 (O_2028,N_24777,N_24994);
nand UO_2029 (O_2029,N_24994,N_24770);
or UO_2030 (O_2030,N_24854,N_24943);
nor UO_2031 (O_2031,N_24989,N_24985);
or UO_2032 (O_2032,N_24896,N_24902);
nand UO_2033 (O_2033,N_24917,N_24825);
nor UO_2034 (O_2034,N_24843,N_24906);
xnor UO_2035 (O_2035,N_24882,N_24952);
nand UO_2036 (O_2036,N_24808,N_24916);
xnor UO_2037 (O_2037,N_24926,N_24820);
xnor UO_2038 (O_2038,N_24924,N_24771);
nor UO_2039 (O_2039,N_24766,N_24807);
and UO_2040 (O_2040,N_24885,N_24890);
and UO_2041 (O_2041,N_24802,N_24973);
or UO_2042 (O_2042,N_24963,N_24906);
or UO_2043 (O_2043,N_24870,N_24767);
or UO_2044 (O_2044,N_24764,N_24766);
nor UO_2045 (O_2045,N_24764,N_24888);
nor UO_2046 (O_2046,N_24991,N_24969);
xnor UO_2047 (O_2047,N_24992,N_24776);
nor UO_2048 (O_2048,N_24923,N_24930);
and UO_2049 (O_2049,N_24969,N_24900);
or UO_2050 (O_2050,N_24939,N_24952);
or UO_2051 (O_2051,N_24972,N_24869);
nand UO_2052 (O_2052,N_24960,N_24767);
or UO_2053 (O_2053,N_24796,N_24873);
or UO_2054 (O_2054,N_24753,N_24821);
or UO_2055 (O_2055,N_24920,N_24778);
or UO_2056 (O_2056,N_24991,N_24846);
xnor UO_2057 (O_2057,N_24938,N_24853);
nand UO_2058 (O_2058,N_24777,N_24883);
nor UO_2059 (O_2059,N_24905,N_24927);
nand UO_2060 (O_2060,N_24997,N_24995);
and UO_2061 (O_2061,N_24998,N_24996);
nor UO_2062 (O_2062,N_24963,N_24888);
nand UO_2063 (O_2063,N_24837,N_24990);
nand UO_2064 (O_2064,N_24848,N_24821);
nand UO_2065 (O_2065,N_24938,N_24751);
and UO_2066 (O_2066,N_24847,N_24843);
xnor UO_2067 (O_2067,N_24876,N_24868);
nor UO_2068 (O_2068,N_24792,N_24807);
nand UO_2069 (O_2069,N_24789,N_24949);
xnor UO_2070 (O_2070,N_24999,N_24922);
and UO_2071 (O_2071,N_24925,N_24752);
xnor UO_2072 (O_2072,N_24757,N_24925);
nand UO_2073 (O_2073,N_24967,N_24797);
and UO_2074 (O_2074,N_24873,N_24768);
nand UO_2075 (O_2075,N_24946,N_24876);
nand UO_2076 (O_2076,N_24759,N_24976);
nor UO_2077 (O_2077,N_24847,N_24880);
xor UO_2078 (O_2078,N_24875,N_24914);
xor UO_2079 (O_2079,N_24983,N_24996);
xor UO_2080 (O_2080,N_24789,N_24782);
nor UO_2081 (O_2081,N_24987,N_24947);
nor UO_2082 (O_2082,N_24970,N_24801);
nand UO_2083 (O_2083,N_24788,N_24930);
or UO_2084 (O_2084,N_24937,N_24750);
xor UO_2085 (O_2085,N_24841,N_24813);
xnor UO_2086 (O_2086,N_24811,N_24946);
nor UO_2087 (O_2087,N_24792,N_24857);
or UO_2088 (O_2088,N_24832,N_24843);
nor UO_2089 (O_2089,N_24770,N_24984);
nand UO_2090 (O_2090,N_24848,N_24924);
nand UO_2091 (O_2091,N_24844,N_24842);
and UO_2092 (O_2092,N_24926,N_24754);
nand UO_2093 (O_2093,N_24979,N_24964);
nor UO_2094 (O_2094,N_24959,N_24810);
xnor UO_2095 (O_2095,N_24870,N_24773);
or UO_2096 (O_2096,N_24966,N_24789);
xor UO_2097 (O_2097,N_24967,N_24889);
or UO_2098 (O_2098,N_24982,N_24875);
or UO_2099 (O_2099,N_24983,N_24842);
and UO_2100 (O_2100,N_24773,N_24933);
and UO_2101 (O_2101,N_24907,N_24984);
and UO_2102 (O_2102,N_24999,N_24839);
nand UO_2103 (O_2103,N_24838,N_24764);
or UO_2104 (O_2104,N_24775,N_24874);
nor UO_2105 (O_2105,N_24828,N_24819);
nand UO_2106 (O_2106,N_24912,N_24813);
and UO_2107 (O_2107,N_24880,N_24939);
xnor UO_2108 (O_2108,N_24776,N_24916);
and UO_2109 (O_2109,N_24843,N_24819);
xnor UO_2110 (O_2110,N_24923,N_24813);
and UO_2111 (O_2111,N_24996,N_24759);
xnor UO_2112 (O_2112,N_24900,N_24889);
or UO_2113 (O_2113,N_24864,N_24943);
nor UO_2114 (O_2114,N_24853,N_24987);
nand UO_2115 (O_2115,N_24981,N_24992);
and UO_2116 (O_2116,N_24915,N_24785);
and UO_2117 (O_2117,N_24937,N_24777);
and UO_2118 (O_2118,N_24814,N_24879);
nand UO_2119 (O_2119,N_24988,N_24940);
or UO_2120 (O_2120,N_24751,N_24802);
nor UO_2121 (O_2121,N_24835,N_24922);
nand UO_2122 (O_2122,N_24877,N_24873);
or UO_2123 (O_2123,N_24821,N_24964);
nor UO_2124 (O_2124,N_24870,N_24905);
nor UO_2125 (O_2125,N_24873,N_24961);
xnor UO_2126 (O_2126,N_24926,N_24981);
or UO_2127 (O_2127,N_24985,N_24830);
and UO_2128 (O_2128,N_24853,N_24828);
xnor UO_2129 (O_2129,N_24932,N_24943);
and UO_2130 (O_2130,N_24788,N_24870);
or UO_2131 (O_2131,N_24869,N_24839);
or UO_2132 (O_2132,N_24957,N_24997);
nand UO_2133 (O_2133,N_24764,N_24964);
nor UO_2134 (O_2134,N_24849,N_24977);
and UO_2135 (O_2135,N_24989,N_24860);
nand UO_2136 (O_2136,N_24990,N_24910);
or UO_2137 (O_2137,N_24912,N_24925);
or UO_2138 (O_2138,N_24827,N_24834);
and UO_2139 (O_2139,N_24773,N_24949);
or UO_2140 (O_2140,N_24884,N_24924);
or UO_2141 (O_2141,N_24778,N_24796);
nor UO_2142 (O_2142,N_24754,N_24979);
nor UO_2143 (O_2143,N_24782,N_24799);
xnor UO_2144 (O_2144,N_24771,N_24852);
nor UO_2145 (O_2145,N_24940,N_24776);
and UO_2146 (O_2146,N_24753,N_24785);
xor UO_2147 (O_2147,N_24938,N_24854);
or UO_2148 (O_2148,N_24838,N_24798);
or UO_2149 (O_2149,N_24865,N_24917);
and UO_2150 (O_2150,N_24812,N_24971);
xnor UO_2151 (O_2151,N_24932,N_24924);
or UO_2152 (O_2152,N_24952,N_24770);
nor UO_2153 (O_2153,N_24757,N_24801);
xnor UO_2154 (O_2154,N_24767,N_24811);
and UO_2155 (O_2155,N_24958,N_24862);
and UO_2156 (O_2156,N_24948,N_24817);
xor UO_2157 (O_2157,N_24822,N_24889);
nand UO_2158 (O_2158,N_24788,N_24950);
xnor UO_2159 (O_2159,N_24805,N_24915);
or UO_2160 (O_2160,N_24857,N_24845);
or UO_2161 (O_2161,N_24767,N_24856);
and UO_2162 (O_2162,N_24841,N_24774);
and UO_2163 (O_2163,N_24818,N_24847);
xor UO_2164 (O_2164,N_24973,N_24972);
or UO_2165 (O_2165,N_24882,N_24859);
xnor UO_2166 (O_2166,N_24795,N_24785);
or UO_2167 (O_2167,N_24753,N_24869);
xnor UO_2168 (O_2168,N_24845,N_24817);
nand UO_2169 (O_2169,N_24972,N_24756);
nand UO_2170 (O_2170,N_24856,N_24802);
xor UO_2171 (O_2171,N_24859,N_24853);
nor UO_2172 (O_2172,N_24873,N_24800);
and UO_2173 (O_2173,N_24981,N_24922);
or UO_2174 (O_2174,N_24863,N_24875);
nor UO_2175 (O_2175,N_24928,N_24906);
or UO_2176 (O_2176,N_24816,N_24836);
and UO_2177 (O_2177,N_24797,N_24878);
nor UO_2178 (O_2178,N_24896,N_24907);
and UO_2179 (O_2179,N_24864,N_24840);
or UO_2180 (O_2180,N_24931,N_24954);
or UO_2181 (O_2181,N_24802,N_24766);
or UO_2182 (O_2182,N_24880,N_24825);
and UO_2183 (O_2183,N_24981,N_24886);
nand UO_2184 (O_2184,N_24776,N_24782);
and UO_2185 (O_2185,N_24974,N_24775);
and UO_2186 (O_2186,N_24857,N_24766);
and UO_2187 (O_2187,N_24761,N_24911);
and UO_2188 (O_2188,N_24967,N_24875);
xnor UO_2189 (O_2189,N_24804,N_24764);
or UO_2190 (O_2190,N_24756,N_24769);
or UO_2191 (O_2191,N_24850,N_24954);
nand UO_2192 (O_2192,N_24926,N_24802);
nand UO_2193 (O_2193,N_24845,N_24831);
and UO_2194 (O_2194,N_24778,N_24916);
nor UO_2195 (O_2195,N_24950,N_24847);
or UO_2196 (O_2196,N_24946,N_24866);
xor UO_2197 (O_2197,N_24965,N_24956);
and UO_2198 (O_2198,N_24979,N_24783);
or UO_2199 (O_2199,N_24762,N_24877);
or UO_2200 (O_2200,N_24979,N_24973);
nand UO_2201 (O_2201,N_24852,N_24881);
and UO_2202 (O_2202,N_24808,N_24755);
xor UO_2203 (O_2203,N_24885,N_24838);
and UO_2204 (O_2204,N_24752,N_24753);
or UO_2205 (O_2205,N_24887,N_24825);
or UO_2206 (O_2206,N_24958,N_24778);
nor UO_2207 (O_2207,N_24766,N_24994);
and UO_2208 (O_2208,N_24808,N_24919);
nor UO_2209 (O_2209,N_24775,N_24993);
xor UO_2210 (O_2210,N_24851,N_24935);
nand UO_2211 (O_2211,N_24934,N_24854);
or UO_2212 (O_2212,N_24930,N_24774);
xnor UO_2213 (O_2213,N_24969,N_24812);
or UO_2214 (O_2214,N_24954,N_24998);
xor UO_2215 (O_2215,N_24811,N_24969);
nand UO_2216 (O_2216,N_24906,N_24863);
and UO_2217 (O_2217,N_24932,N_24916);
and UO_2218 (O_2218,N_24884,N_24770);
xor UO_2219 (O_2219,N_24964,N_24983);
or UO_2220 (O_2220,N_24937,N_24882);
xnor UO_2221 (O_2221,N_24844,N_24916);
and UO_2222 (O_2222,N_24868,N_24900);
nor UO_2223 (O_2223,N_24793,N_24776);
xor UO_2224 (O_2224,N_24900,N_24966);
nand UO_2225 (O_2225,N_24860,N_24909);
nand UO_2226 (O_2226,N_24817,N_24952);
nor UO_2227 (O_2227,N_24969,N_24774);
nand UO_2228 (O_2228,N_24947,N_24886);
or UO_2229 (O_2229,N_24841,N_24955);
and UO_2230 (O_2230,N_24923,N_24939);
xor UO_2231 (O_2231,N_24918,N_24939);
nand UO_2232 (O_2232,N_24868,N_24962);
nor UO_2233 (O_2233,N_24918,N_24964);
nand UO_2234 (O_2234,N_24962,N_24802);
or UO_2235 (O_2235,N_24972,N_24843);
or UO_2236 (O_2236,N_24758,N_24824);
nand UO_2237 (O_2237,N_24944,N_24920);
nand UO_2238 (O_2238,N_24835,N_24881);
and UO_2239 (O_2239,N_24782,N_24818);
xnor UO_2240 (O_2240,N_24966,N_24934);
and UO_2241 (O_2241,N_24851,N_24958);
or UO_2242 (O_2242,N_24932,N_24803);
xor UO_2243 (O_2243,N_24938,N_24827);
xnor UO_2244 (O_2244,N_24891,N_24758);
nor UO_2245 (O_2245,N_24840,N_24961);
nor UO_2246 (O_2246,N_24912,N_24887);
xnor UO_2247 (O_2247,N_24867,N_24763);
nor UO_2248 (O_2248,N_24886,N_24774);
nor UO_2249 (O_2249,N_24900,N_24800);
nor UO_2250 (O_2250,N_24786,N_24758);
nand UO_2251 (O_2251,N_24840,N_24832);
nand UO_2252 (O_2252,N_24967,N_24935);
xnor UO_2253 (O_2253,N_24949,N_24751);
or UO_2254 (O_2254,N_24838,N_24903);
nand UO_2255 (O_2255,N_24901,N_24928);
nor UO_2256 (O_2256,N_24854,N_24754);
xor UO_2257 (O_2257,N_24999,N_24969);
and UO_2258 (O_2258,N_24755,N_24751);
nor UO_2259 (O_2259,N_24880,N_24871);
and UO_2260 (O_2260,N_24963,N_24950);
xnor UO_2261 (O_2261,N_24993,N_24811);
nand UO_2262 (O_2262,N_24834,N_24818);
and UO_2263 (O_2263,N_24934,N_24896);
xnor UO_2264 (O_2264,N_24809,N_24786);
xor UO_2265 (O_2265,N_24911,N_24859);
xor UO_2266 (O_2266,N_24844,N_24950);
or UO_2267 (O_2267,N_24805,N_24844);
nand UO_2268 (O_2268,N_24795,N_24896);
or UO_2269 (O_2269,N_24891,N_24894);
xor UO_2270 (O_2270,N_24826,N_24976);
or UO_2271 (O_2271,N_24770,N_24882);
and UO_2272 (O_2272,N_24959,N_24800);
xnor UO_2273 (O_2273,N_24829,N_24817);
nand UO_2274 (O_2274,N_24839,N_24879);
nand UO_2275 (O_2275,N_24763,N_24979);
and UO_2276 (O_2276,N_24970,N_24959);
or UO_2277 (O_2277,N_24853,N_24982);
nand UO_2278 (O_2278,N_24888,N_24951);
xor UO_2279 (O_2279,N_24903,N_24763);
or UO_2280 (O_2280,N_24939,N_24804);
nand UO_2281 (O_2281,N_24899,N_24916);
and UO_2282 (O_2282,N_24787,N_24986);
nor UO_2283 (O_2283,N_24764,N_24949);
nor UO_2284 (O_2284,N_24797,N_24922);
nor UO_2285 (O_2285,N_24868,N_24975);
xor UO_2286 (O_2286,N_24971,N_24847);
and UO_2287 (O_2287,N_24839,N_24753);
nor UO_2288 (O_2288,N_24984,N_24886);
and UO_2289 (O_2289,N_24930,N_24756);
nand UO_2290 (O_2290,N_24938,N_24953);
or UO_2291 (O_2291,N_24892,N_24953);
nand UO_2292 (O_2292,N_24856,N_24987);
or UO_2293 (O_2293,N_24901,N_24791);
and UO_2294 (O_2294,N_24829,N_24996);
nand UO_2295 (O_2295,N_24762,N_24969);
xnor UO_2296 (O_2296,N_24793,N_24999);
or UO_2297 (O_2297,N_24880,N_24832);
or UO_2298 (O_2298,N_24867,N_24972);
nor UO_2299 (O_2299,N_24821,N_24912);
nand UO_2300 (O_2300,N_24982,N_24946);
nand UO_2301 (O_2301,N_24791,N_24955);
or UO_2302 (O_2302,N_24885,N_24942);
nor UO_2303 (O_2303,N_24969,N_24920);
and UO_2304 (O_2304,N_24903,N_24907);
nor UO_2305 (O_2305,N_24966,N_24775);
nor UO_2306 (O_2306,N_24777,N_24850);
nor UO_2307 (O_2307,N_24839,N_24851);
nand UO_2308 (O_2308,N_24832,N_24808);
or UO_2309 (O_2309,N_24954,N_24758);
and UO_2310 (O_2310,N_24899,N_24802);
and UO_2311 (O_2311,N_24925,N_24914);
or UO_2312 (O_2312,N_24928,N_24853);
nand UO_2313 (O_2313,N_24898,N_24921);
and UO_2314 (O_2314,N_24952,N_24979);
and UO_2315 (O_2315,N_24843,N_24811);
nor UO_2316 (O_2316,N_24890,N_24906);
xor UO_2317 (O_2317,N_24774,N_24758);
xnor UO_2318 (O_2318,N_24859,N_24975);
and UO_2319 (O_2319,N_24806,N_24874);
xor UO_2320 (O_2320,N_24833,N_24931);
and UO_2321 (O_2321,N_24906,N_24907);
nor UO_2322 (O_2322,N_24976,N_24921);
nor UO_2323 (O_2323,N_24839,N_24949);
or UO_2324 (O_2324,N_24994,N_24974);
xor UO_2325 (O_2325,N_24888,N_24932);
or UO_2326 (O_2326,N_24985,N_24979);
xor UO_2327 (O_2327,N_24852,N_24989);
or UO_2328 (O_2328,N_24893,N_24818);
or UO_2329 (O_2329,N_24953,N_24782);
nand UO_2330 (O_2330,N_24920,N_24839);
and UO_2331 (O_2331,N_24988,N_24908);
and UO_2332 (O_2332,N_24898,N_24884);
nand UO_2333 (O_2333,N_24906,N_24777);
and UO_2334 (O_2334,N_24830,N_24934);
or UO_2335 (O_2335,N_24795,N_24969);
xnor UO_2336 (O_2336,N_24991,N_24867);
or UO_2337 (O_2337,N_24856,N_24786);
nor UO_2338 (O_2338,N_24774,N_24888);
nor UO_2339 (O_2339,N_24990,N_24870);
and UO_2340 (O_2340,N_24900,N_24816);
nand UO_2341 (O_2341,N_24755,N_24901);
nand UO_2342 (O_2342,N_24780,N_24834);
and UO_2343 (O_2343,N_24848,N_24816);
nand UO_2344 (O_2344,N_24908,N_24919);
nor UO_2345 (O_2345,N_24980,N_24850);
xnor UO_2346 (O_2346,N_24857,N_24778);
xnor UO_2347 (O_2347,N_24894,N_24819);
xnor UO_2348 (O_2348,N_24871,N_24884);
and UO_2349 (O_2349,N_24753,N_24906);
nand UO_2350 (O_2350,N_24941,N_24755);
nor UO_2351 (O_2351,N_24971,N_24855);
xor UO_2352 (O_2352,N_24835,N_24823);
or UO_2353 (O_2353,N_24929,N_24851);
nand UO_2354 (O_2354,N_24777,N_24964);
or UO_2355 (O_2355,N_24992,N_24932);
nor UO_2356 (O_2356,N_24840,N_24793);
or UO_2357 (O_2357,N_24963,N_24762);
and UO_2358 (O_2358,N_24968,N_24913);
nand UO_2359 (O_2359,N_24964,N_24891);
xnor UO_2360 (O_2360,N_24917,N_24785);
xor UO_2361 (O_2361,N_24823,N_24834);
nor UO_2362 (O_2362,N_24865,N_24918);
xor UO_2363 (O_2363,N_24876,N_24959);
or UO_2364 (O_2364,N_24969,N_24996);
nor UO_2365 (O_2365,N_24779,N_24904);
nor UO_2366 (O_2366,N_24758,N_24779);
xor UO_2367 (O_2367,N_24853,N_24865);
nor UO_2368 (O_2368,N_24917,N_24866);
nand UO_2369 (O_2369,N_24820,N_24885);
nand UO_2370 (O_2370,N_24980,N_24772);
nor UO_2371 (O_2371,N_24894,N_24797);
and UO_2372 (O_2372,N_24801,N_24852);
and UO_2373 (O_2373,N_24990,N_24960);
nor UO_2374 (O_2374,N_24793,N_24916);
and UO_2375 (O_2375,N_24899,N_24825);
and UO_2376 (O_2376,N_24766,N_24905);
nand UO_2377 (O_2377,N_24794,N_24983);
and UO_2378 (O_2378,N_24962,N_24814);
nor UO_2379 (O_2379,N_24850,N_24773);
xor UO_2380 (O_2380,N_24916,N_24839);
nor UO_2381 (O_2381,N_24801,N_24971);
xnor UO_2382 (O_2382,N_24781,N_24847);
xor UO_2383 (O_2383,N_24765,N_24764);
and UO_2384 (O_2384,N_24978,N_24823);
xnor UO_2385 (O_2385,N_24764,N_24919);
and UO_2386 (O_2386,N_24785,N_24923);
and UO_2387 (O_2387,N_24941,N_24843);
nand UO_2388 (O_2388,N_24889,N_24815);
nand UO_2389 (O_2389,N_24879,N_24984);
nand UO_2390 (O_2390,N_24970,N_24993);
and UO_2391 (O_2391,N_24967,N_24998);
xor UO_2392 (O_2392,N_24865,N_24763);
nor UO_2393 (O_2393,N_24781,N_24783);
nand UO_2394 (O_2394,N_24873,N_24834);
nand UO_2395 (O_2395,N_24756,N_24954);
nor UO_2396 (O_2396,N_24798,N_24897);
and UO_2397 (O_2397,N_24855,N_24857);
nand UO_2398 (O_2398,N_24969,N_24861);
nor UO_2399 (O_2399,N_24857,N_24884);
and UO_2400 (O_2400,N_24983,N_24782);
nor UO_2401 (O_2401,N_24909,N_24943);
nand UO_2402 (O_2402,N_24806,N_24761);
nand UO_2403 (O_2403,N_24955,N_24974);
or UO_2404 (O_2404,N_24932,N_24779);
xnor UO_2405 (O_2405,N_24916,N_24949);
or UO_2406 (O_2406,N_24877,N_24759);
nor UO_2407 (O_2407,N_24788,N_24889);
xnor UO_2408 (O_2408,N_24846,N_24926);
or UO_2409 (O_2409,N_24787,N_24754);
nand UO_2410 (O_2410,N_24847,N_24949);
nand UO_2411 (O_2411,N_24859,N_24815);
and UO_2412 (O_2412,N_24823,N_24951);
xnor UO_2413 (O_2413,N_24853,N_24852);
nand UO_2414 (O_2414,N_24798,N_24883);
or UO_2415 (O_2415,N_24926,N_24987);
nand UO_2416 (O_2416,N_24782,N_24851);
xor UO_2417 (O_2417,N_24934,N_24851);
xnor UO_2418 (O_2418,N_24809,N_24821);
xor UO_2419 (O_2419,N_24760,N_24916);
xnor UO_2420 (O_2420,N_24797,N_24988);
xnor UO_2421 (O_2421,N_24759,N_24989);
nor UO_2422 (O_2422,N_24871,N_24820);
or UO_2423 (O_2423,N_24892,N_24972);
and UO_2424 (O_2424,N_24965,N_24888);
nor UO_2425 (O_2425,N_24883,N_24840);
nor UO_2426 (O_2426,N_24987,N_24796);
nor UO_2427 (O_2427,N_24917,N_24833);
nor UO_2428 (O_2428,N_24837,N_24895);
and UO_2429 (O_2429,N_24772,N_24985);
nor UO_2430 (O_2430,N_24826,N_24777);
nor UO_2431 (O_2431,N_24994,N_24875);
or UO_2432 (O_2432,N_24781,N_24864);
and UO_2433 (O_2433,N_24959,N_24808);
or UO_2434 (O_2434,N_24850,N_24858);
nand UO_2435 (O_2435,N_24770,N_24806);
nand UO_2436 (O_2436,N_24922,N_24852);
xor UO_2437 (O_2437,N_24788,N_24993);
nor UO_2438 (O_2438,N_24952,N_24776);
nor UO_2439 (O_2439,N_24830,N_24957);
or UO_2440 (O_2440,N_24800,N_24828);
and UO_2441 (O_2441,N_24959,N_24859);
nand UO_2442 (O_2442,N_24953,N_24904);
xnor UO_2443 (O_2443,N_24760,N_24932);
or UO_2444 (O_2444,N_24987,N_24952);
xor UO_2445 (O_2445,N_24753,N_24970);
nand UO_2446 (O_2446,N_24783,N_24972);
and UO_2447 (O_2447,N_24940,N_24944);
and UO_2448 (O_2448,N_24764,N_24977);
and UO_2449 (O_2449,N_24993,N_24855);
or UO_2450 (O_2450,N_24878,N_24956);
nor UO_2451 (O_2451,N_24787,N_24752);
xor UO_2452 (O_2452,N_24966,N_24768);
or UO_2453 (O_2453,N_24855,N_24849);
nor UO_2454 (O_2454,N_24801,N_24862);
or UO_2455 (O_2455,N_24883,N_24782);
or UO_2456 (O_2456,N_24977,N_24972);
and UO_2457 (O_2457,N_24948,N_24854);
nor UO_2458 (O_2458,N_24793,N_24791);
or UO_2459 (O_2459,N_24793,N_24836);
nor UO_2460 (O_2460,N_24751,N_24884);
and UO_2461 (O_2461,N_24951,N_24905);
or UO_2462 (O_2462,N_24832,N_24882);
xnor UO_2463 (O_2463,N_24966,N_24919);
nand UO_2464 (O_2464,N_24814,N_24925);
xnor UO_2465 (O_2465,N_24920,N_24875);
nand UO_2466 (O_2466,N_24908,N_24856);
or UO_2467 (O_2467,N_24794,N_24778);
xor UO_2468 (O_2468,N_24890,N_24755);
and UO_2469 (O_2469,N_24978,N_24833);
nor UO_2470 (O_2470,N_24848,N_24913);
nor UO_2471 (O_2471,N_24806,N_24809);
xor UO_2472 (O_2472,N_24805,N_24939);
and UO_2473 (O_2473,N_24926,N_24801);
xor UO_2474 (O_2474,N_24885,N_24796);
and UO_2475 (O_2475,N_24758,N_24869);
nor UO_2476 (O_2476,N_24955,N_24903);
xnor UO_2477 (O_2477,N_24897,N_24779);
and UO_2478 (O_2478,N_24761,N_24830);
or UO_2479 (O_2479,N_24935,N_24973);
xor UO_2480 (O_2480,N_24941,N_24834);
nor UO_2481 (O_2481,N_24871,N_24991);
nand UO_2482 (O_2482,N_24940,N_24815);
or UO_2483 (O_2483,N_24951,N_24938);
nand UO_2484 (O_2484,N_24784,N_24896);
xor UO_2485 (O_2485,N_24885,N_24916);
or UO_2486 (O_2486,N_24942,N_24912);
and UO_2487 (O_2487,N_24908,N_24773);
nor UO_2488 (O_2488,N_24917,N_24852);
xor UO_2489 (O_2489,N_24994,N_24957);
or UO_2490 (O_2490,N_24813,N_24988);
and UO_2491 (O_2491,N_24951,N_24912);
xor UO_2492 (O_2492,N_24950,N_24994);
or UO_2493 (O_2493,N_24967,N_24776);
or UO_2494 (O_2494,N_24983,N_24883);
nand UO_2495 (O_2495,N_24836,N_24807);
xor UO_2496 (O_2496,N_24980,N_24762);
xor UO_2497 (O_2497,N_24955,N_24902);
nor UO_2498 (O_2498,N_24959,N_24870);
nand UO_2499 (O_2499,N_24866,N_24913);
nor UO_2500 (O_2500,N_24848,N_24889);
nand UO_2501 (O_2501,N_24892,N_24826);
nor UO_2502 (O_2502,N_24934,N_24790);
or UO_2503 (O_2503,N_24767,N_24976);
or UO_2504 (O_2504,N_24916,N_24847);
nand UO_2505 (O_2505,N_24965,N_24869);
and UO_2506 (O_2506,N_24972,N_24881);
nor UO_2507 (O_2507,N_24863,N_24923);
xnor UO_2508 (O_2508,N_24757,N_24869);
xnor UO_2509 (O_2509,N_24869,N_24769);
nand UO_2510 (O_2510,N_24782,N_24919);
and UO_2511 (O_2511,N_24754,N_24819);
nand UO_2512 (O_2512,N_24958,N_24886);
and UO_2513 (O_2513,N_24899,N_24985);
nand UO_2514 (O_2514,N_24926,N_24772);
or UO_2515 (O_2515,N_24903,N_24802);
nand UO_2516 (O_2516,N_24848,N_24951);
nor UO_2517 (O_2517,N_24876,N_24964);
and UO_2518 (O_2518,N_24946,N_24833);
and UO_2519 (O_2519,N_24917,N_24877);
nor UO_2520 (O_2520,N_24775,N_24981);
and UO_2521 (O_2521,N_24956,N_24847);
nor UO_2522 (O_2522,N_24976,N_24989);
xnor UO_2523 (O_2523,N_24944,N_24771);
xnor UO_2524 (O_2524,N_24945,N_24759);
or UO_2525 (O_2525,N_24795,N_24871);
xnor UO_2526 (O_2526,N_24921,N_24750);
nand UO_2527 (O_2527,N_24766,N_24896);
and UO_2528 (O_2528,N_24761,N_24804);
nand UO_2529 (O_2529,N_24860,N_24885);
nor UO_2530 (O_2530,N_24970,N_24852);
nor UO_2531 (O_2531,N_24890,N_24860);
nor UO_2532 (O_2532,N_24858,N_24865);
and UO_2533 (O_2533,N_24952,N_24978);
xor UO_2534 (O_2534,N_24973,N_24919);
xor UO_2535 (O_2535,N_24991,N_24954);
nor UO_2536 (O_2536,N_24804,N_24795);
nand UO_2537 (O_2537,N_24838,N_24822);
or UO_2538 (O_2538,N_24818,N_24889);
nor UO_2539 (O_2539,N_24857,N_24784);
xor UO_2540 (O_2540,N_24963,N_24913);
or UO_2541 (O_2541,N_24876,N_24798);
or UO_2542 (O_2542,N_24814,N_24762);
nor UO_2543 (O_2543,N_24940,N_24808);
xnor UO_2544 (O_2544,N_24878,N_24806);
or UO_2545 (O_2545,N_24905,N_24784);
nand UO_2546 (O_2546,N_24795,N_24848);
xnor UO_2547 (O_2547,N_24896,N_24852);
xnor UO_2548 (O_2548,N_24806,N_24949);
nor UO_2549 (O_2549,N_24867,N_24778);
and UO_2550 (O_2550,N_24971,N_24979);
nor UO_2551 (O_2551,N_24804,N_24823);
and UO_2552 (O_2552,N_24773,N_24840);
and UO_2553 (O_2553,N_24785,N_24930);
xor UO_2554 (O_2554,N_24838,N_24939);
xnor UO_2555 (O_2555,N_24869,N_24881);
nand UO_2556 (O_2556,N_24928,N_24811);
nand UO_2557 (O_2557,N_24808,N_24879);
or UO_2558 (O_2558,N_24794,N_24872);
nor UO_2559 (O_2559,N_24899,N_24881);
or UO_2560 (O_2560,N_24891,N_24954);
xor UO_2561 (O_2561,N_24993,N_24781);
and UO_2562 (O_2562,N_24768,N_24960);
and UO_2563 (O_2563,N_24930,N_24926);
and UO_2564 (O_2564,N_24839,N_24900);
and UO_2565 (O_2565,N_24807,N_24911);
nor UO_2566 (O_2566,N_24982,N_24939);
nor UO_2567 (O_2567,N_24850,N_24940);
or UO_2568 (O_2568,N_24949,N_24939);
or UO_2569 (O_2569,N_24907,N_24802);
or UO_2570 (O_2570,N_24857,N_24777);
or UO_2571 (O_2571,N_24987,N_24793);
and UO_2572 (O_2572,N_24790,N_24833);
nor UO_2573 (O_2573,N_24847,N_24970);
nor UO_2574 (O_2574,N_24910,N_24967);
nand UO_2575 (O_2575,N_24896,N_24933);
nor UO_2576 (O_2576,N_24968,N_24967);
xnor UO_2577 (O_2577,N_24847,N_24941);
or UO_2578 (O_2578,N_24753,N_24794);
nand UO_2579 (O_2579,N_24989,N_24844);
and UO_2580 (O_2580,N_24863,N_24884);
xnor UO_2581 (O_2581,N_24776,N_24907);
nand UO_2582 (O_2582,N_24795,N_24928);
and UO_2583 (O_2583,N_24971,N_24816);
xnor UO_2584 (O_2584,N_24884,N_24914);
or UO_2585 (O_2585,N_24783,N_24967);
xor UO_2586 (O_2586,N_24952,N_24808);
or UO_2587 (O_2587,N_24962,N_24954);
nor UO_2588 (O_2588,N_24838,N_24752);
xnor UO_2589 (O_2589,N_24779,N_24766);
nor UO_2590 (O_2590,N_24824,N_24921);
or UO_2591 (O_2591,N_24813,N_24940);
nand UO_2592 (O_2592,N_24856,N_24963);
nor UO_2593 (O_2593,N_24856,N_24920);
or UO_2594 (O_2594,N_24772,N_24892);
nand UO_2595 (O_2595,N_24773,N_24983);
nand UO_2596 (O_2596,N_24914,N_24840);
or UO_2597 (O_2597,N_24990,N_24788);
or UO_2598 (O_2598,N_24825,N_24836);
xnor UO_2599 (O_2599,N_24759,N_24846);
xnor UO_2600 (O_2600,N_24867,N_24837);
nand UO_2601 (O_2601,N_24910,N_24817);
or UO_2602 (O_2602,N_24981,N_24947);
or UO_2603 (O_2603,N_24951,N_24757);
and UO_2604 (O_2604,N_24796,N_24821);
or UO_2605 (O_2605,N_24976,N_24881);
nand UO_2606 (O_2606,N_24826,N_24950);
or UO_2607 (O_2607,N_24792,N_24979);
nor UO_2608 (O_2608,N_24756,N_24900);
or UO_2609 (O_2609,N_24866,N_24851);
xor UO_2610 (O_2610,N_24791,N_24971);
nand UO_2611 (O_2611,N_24928,N_24984);
nand UO_2612 (O_2612,N_24896,N_24873);
and UO_2613 (O_2613,N_24906,N_24979);
xnor UO_2614 (O_2614,N_24762,N_24763);
nor UO_2615 (O_2615,N_24872,N_24807);
xor UO_2616 (O_2616,N_24842,N_24963);
and UO_2617 (O_2617,N_24755,N_24954);
and UO_2618 (O_2618,N_24955,N_24965);
nor UO_2619 (O_2619,N_24820,N_24862);
or UO_2620 (O_2620,N_24864,N_24816);
or UO_2621 (O_2621,N_24832,N_24766);
or UO_2622 (O_2622,N_24801,N_24975);
xnor UO_2623 (O_2623,N_24953,N_24841);
nor UO_2624 (O_2624,N_24795,N_24863);
or UO_2625 (O_2625,N_24769,N_24802);
xnor UO_2626 (O_2626,N_24914,N_24939);
nand UO_2627 (O_2627,N_24814,N_24837);
xor UO_2628 (O_2628,N_24824,N_24933);
nor UO_2629 (O_2629,N_24918,N_24770);
xor UO_2630 (O_2630,N_24804,N_24896);
and UO_2631 (O_2631,N_24881,N_24969);
or UO_2632 (O_2632,N_24926,N_24938);
or UO_2633 (O_2633,N_24854,N_24919);
xnor UO_2634 (O_2634,N_24934,N_24980);
nand UO_2635 (O_2635,N_24760,N_24761);
nand UO_2636 (O_2636,N_24833,N_24771);
xnor UO_2637 (O_2637,N_24963,N_24907);
or UO_2638 (O_2638,N_24947,N_24980);
and UO_2639 (O_2639,N_24963,N_24872);
nand UO_2640 (O_2640,N_24876,N_24873);
and UO_2641 (O_2641,N_24759,N_24938);
nand UO_2642 (O_2642,N_24792,N_24947);
and UO_2643 (O_2643,N_24897,N_24945);
and UO_2644 (O_2644,N_24774,N_24926);
nor UO_2645 (O_2645,N_24803,N_24916);
nor UO_2646 (O_2646,N_24915,N_24885);
and UO_2647 (O_2647,N_24886,N_24998);
nor UO_2648 (O_2648,N_24860,N_24759);
and UO_2649 (O_2649,N_24921,N_24994);
nand UO_2650 (O_2650,N_24996,N_24766);
xor UO_2651 (O_2651,N_24825,N_24756);
xor UO_2652 (O_2652,N_24989,N_24888);
xnor UO_2653 (O_2653,N_24787,N_24862);
nand UO_2654 (O_2654,N_24819,N_24845);
or UO_2655 (O_2655,N_24882,N_24962);
nor UO_2656 (O_2656,N_24796,N_24818);
or UO_2657 (O_2657,N_24885,N_24861);
nand UO_2658 (O_2658,N_24785,N_24977);
and UO_2659 (O_2659,N_24823,N_24790);
nor UO_2660 (O_2660,N_24866,N_24771);
xnor UO_2661 (O_2661,N_24970,N_24988);
xnor UO_2662 (O_2662,N_24900,N_24886);
nand UO_2663 (O_2663,N_24969,N_24956);
or UO_2664 (O_2664,N_24995,N_24999);
nor UO_2665 (O_2665,N_24835,N_24964);
xnor UO_2666 (O_2666,N_24909,N_24955);
nand UO_2667 (O_2667,N_24781,N_24876);
and UO_2668 (O_2668,N_24926,N_24916);
or UO_2669 (O_2669,N_24870,N_24823);
xnor UO_2670 (O_2670,N_24973,N_24895);
or UO_2671 (O_2671,N_24804,N_24882);
nor UO_2672 (O_2672,N_24871,N_24801);
xor UO_2673 (O_2673,N_24766,N_24818);
xnor UO_2674 (O_2674,N_24901,N_24873);
nand UO_2675 (O_2675,N_24979,N_24779);
nand UO_2676 (O_2676,N_24791,N_24878);
nor UO_2677 (O_2677,N_24921,N_24853);
xor UO_2678 (O_2678,N_24932,N_24770);
xnor UO_2679 (O_2679,N_24882,N_24858);
xor UO_2680 (O_2680,N_24828,N_24795);
nor UO_2681 (O_2681,N_24947,N_24823);
nor UO_2682 (O_2682,N_24903,N_24754);
xnor UO_2683 (O_2683,N_24851,N_24949);
or UO_2684 (O_2684,N_24917,N_24831);
or UO_2685 (O_2685,N_24858,N_24909);
and UO_2686 (O_2686,N_24781,N_24790);
nor UO_2687 (O_2687,N_24843,N_24786);
xnor UO_2688 (O_2688,N_24966,N_24877);
nor UO_2689 (O_2689,N_24817,N_24909);
and UO_2690 (O_2690,N_24922,N_24843);
and UO_2691 (O_2691,N_24865,N_24983);
nor UO_2692 (O_2692,N_24895,N_24856);
or UO_2693 (O_2693,N_24986,N_24857);
nand UO_2694 (O_2694,N_24981,N_24939);
nand UO_2695 (O_2695,N_24894,N_24867);
nand UO_2696 (O_2696,N_24791,N_24839);
xnor UO_2697 (O_2697,N_24797,N_24867);
nor UO_2698 (O_2698,N_24804,N_24841);
nand UO_2699 (O_2699,N_24983,N_24871);
nor UO_2700 (O_2700,N_24909,N_24908);
and UO_2701 (O_2701,N_24948,N_24870);
and UO_2702 (O_2702,N_24781,N_24887);
or UO_2703 (O_2703,N_24895,N_24897);
nor UO_2704 (O_2704,N_24974,N_24947);
or UO_2705 (O_2705,N_24920,N_24910);
nand UO_2706 (O_2706,N_24839,N_24836);
nor UO_2707 (O_2707,N_24829,N_24984);
and UO_2708 (O_2708,N_24828,N_24781);
nand UO_2709 (O_2709,N_24880,N_24786);
nor UO_2710 (O_2710,N_24921,N_24962);
or UO_2711 (O_2711,N_24998,N_24942);
xor UO_2712 (O_2712,N_24752,N_24784);
xor UO_2713 (O_2713,N_24998,N_24979);
nand UO_2714 (O_2714,N_24839,N_24967);
nor UO_2715 (O_2715,N_24886,N_24901);
nand UO_2716 (O_2716,N_24860,N_24954);
xnor UO_2717 (O_2717,N_24878,N_24998);
or UO_2718 (O_2718,N_24766,N_24936);
and UO_2719 (O_2719,N_24811,N_24992);
or UO_2720 (O_2720,N_24921,N_24861);
xnor UO_2721 (O_2721,N_24916,N_24824);
nand UO_2722 (O_2722,N_24830,N_24801);
and UO_2723 (O_2723,N_24855,N_24885);
and UO_2724 (O_2724,N_24813,N_24990);
nand UO_2725 (O_2725,N_24856,N_24994);
nor UO_2726 (O_2726,N_24789,N_24948);
or UO_2727 (O_2727,N_24973,N_24915);
and UO_2728 (O_2728,N_24832,N_24799);
xnor UO_2729 (O_2729,N_24787,N_24874);
nor UO_2730 (O_2730,N_24801,N_24896);
nand UO_2731 (O_2731,N_24997,N_24792);
nor UO_2732 (O_2732,N_24955,N_24931);
nor UO_2733 (O_2733,N_24998,N_24990);
nor UO_2734 (O_2734,N_24805,N_24753);
nor UO_2735 (O_2735,N_24947,N_24896);
nor UO_2736 (O_2736,N_24896,N_24832);
nand UO_2737 (O_2737,N_24786,N_24929);
nand UO_2738 (O_2738,N_24930,N_24961);
or UO_2739 (O_2739,N_24871,N_24808);
xor UO_2740 (O_2740,N_24961,N_24848);
nand UO_2741 (O_2741,N_24879,N_24871);
xnor UO_2742 (O_2742,N_24931,N_24888);
nand UO_2743 (O_2743,N_24789,N_24954);
nor UO_2744 (O_2744,N_24946,N_24869);
xor UO_2745 (O_2745,N_24901,N_24826);
xnor UO_2746 (O_2746,N_24982,N_24765);
or UO_2747 (O_2747,N_24752,N_24946);
xor UO_2748 (O_2748,N_24845,N_24828);
nand UO_2749 (O_2749,N_24825,N_24778);
xor UO_2750 (O_2750,N_24779,N_24770);
xor UO_2751 (O_2751,N_24761,N_24943);
and UO_2752 (O_2752,N_24752,N_24799);
or UO_2753 (O_2753,N_24885,N_24895);
nand UO_2754 (O_2754,N_24805,N_24751);
and UO_2755 (O_2755,N_24990,N_24949);
xor UO_2756 (O_2756,N_24996,N_24818);
nor UO_2757 (O_2757,N_24924,N_24851);
nor UO_2758 (O_2758,N_24817,N_24784);
and UO_2759 (O_2759,N_24982,N_24886);
and UO_2760 (O_2760,N_24942,N_24979);
and UO_2761 (O_2761,N_24845,N_24909);
or UO_2762 (O_2762,N_24758,N_24799);
and UO_2763 (O_2763,N_24947,N_24903);
nand UO_2764 (O_2764,N_24985,N_24775);
xnor UO_2765 (O_2765,N_24769,N_24994);
or UO_2766 (O_2766,N_24937,N_24880);
nor UO_2767 (O_2767,N_24893,N_24806);
nand UO_2768 (O_2768,N_24880,N_24921);
xor UO_2769 (O_2769,N_24882,N_24803);
and UO_2770 (O_2770,N_24818,N_24833);
xnor UO_2771 (O_2771,N_24814,N_24855);
xor UO_2772 (O_2772,N_24780,N_24766);
or UO_2773 (O_2773,N_24860,N_24859);
or UO_2774 (O_2774,N_24878,N_24982);
xnor UO_2775 (O_2775,N_24787,N_24899);
and UO_2776 (O_2776,N_24817,N_24983);
xor UO_2777 (O_2777,N_24952,N_24842);
nand UO_2778 (O_2778,N_24841,N_24904);
or UO_2779 (O_2779,N_24764,N_24931);
and UO_2780 (O_2780,N_24937,N_24900);
nor UO_2781 (O_2781,N_24962,N_24970);
xnor UO_2782 (O_2782,N_24877,N_24768);
xor UO_2783 (O_2783,N_24967,N_24972);
nor UO_2784 (O_2784,N_24805,N_24837);
or UO_2785 (O_2785,N_24905,N_24891);
nor UO_2786 (O_2786,N_24873,N_24778);
and UO_2787 (O_2787,N_24848,N_24988);
or UO_2788 (O_2788,N_24941,N_24870);
nand UO_2789 (O_2789,N_24849,N_24919);
or UO_2790 (O_2790,N_24794,N_24760);
and UO_2791 (O_2791,N_24770,N_24756);
and UO_2792 (O_2792,N_24784,N_24989);
or UO_2793 (O_2793,N_24975,N_24778);
nand UO_2794 (O_2794,N_24980,N_24817);
xor UO_2795 (O_2795,N_24955,N_24877);
or UO_2796 (O_2796,N_24821,N_24778);
nor UO_2797 (O_2797,N_24830,N_24915);
and UO_2798 (O_2798,N_24812,N_24918);
and UO_2799 (O_2799,N_24889,N_24916);
and UO_2800 (O_2800,N_24970,N_24845);
xor UO_2801 (O_2801,N_24972,N_24946);
nand UO_2802 (O_2802,N_24834,N_24866);
and UO_2803 (O_2803,N_24752,N_24957);
and UO_2804 (O_2804,N_24997,N_24876);
and UO_2805 (O_2805,N_24763,N_24918);
nand UO_2806 (O_2806,N_24905,N_24880);
nand UO_2807 (O_2807,N_24810,N_24835);
nor UO_2808 (O_2808,N_24819,N_24806);
xnor UO_2809 (O_2809,N_24901,N_24768);
nand UO_2810 (O_2810,N_24848,N_24974);
nor UO_2811 (O_2811,N_24830,N_24760);
nand UO_2812 (O_2812,N_24894,N_24756);
and UO_2813 (O_2813,N_24759,N_24872);
nand UO_2814 (O_2814,N_24817,N_24978);
and UO_2815 (O_2815,N_24762,N_24988);
and UO_2816 (O_2816,N_24894,N_24847);
nand UO_2817 (O_2817,N_24994,N_24836);
nand UO_2818 (O_2818,N_24945,N_24851);
or UO_2819 (O_2819,N_24957,N_24846);
nor UO_2820 (O_2820,N_24874,N_24921);
nor UO_2821 (O_2821,N_24921,N_24836);
nor UO_2822 (O_2822,N_24822,N_24895);
or UO_2823 (O_2823,N_24925,N_24922);
and UO_2824 (O_2824,N_24800,N_24832);
xnor UO_2825 (O_2825,N_24898,N_24985);
and UO_2826 (O_2826,N_24997,N_24764);
nand UO_2827 (O_2827,N_24987,N_24800);
or UO_2828 (O_2828,N_24980,N_24936);
nor UO_2829 (O_2829,N_24968,N_24799);
and UO_2830 (O_2830,N_24770,N_24769);
nor UO_2831 (O_2831,N_24910,N_24868);
nand UO_2832 (O_2832,N_24883,N_24917);
and UO_2833 (O_2833,N_24982,N_24821);
nand UO_2834 (O_2834,N_24891,N_24851);
or UO_2835 (O_2835,N_24919,N_24823);
and UO_2836 (O_2836,N_24776,N_24993);
xnor UO_2837 (O_2837,N_24958,N_24892);
nor UO_2838 (O_2838,N_24826,N_24882);
xnor UO_2839 (O_2839,N_24836,N_24766);
and UO_2840 (O_2840,N_24771,N_24987);
or UO_2841 (O_2841,N_24945,N_24953);
nor UO_2842 (O_2842,N_24789,N_24915);
or UO_2843 (O_2843,N_24975,N_24794);
xor UO_2844 (O_2844,N_24834,N_24841);
or UO_2845 (O_2845,N_24776,N_24816);
or UO_2846 (O_2846,N_24971,N_24973);
xnor UO_2847 (O_2847,N_24940,N_24796);
and UO_2848 (O_2848,N_24765,N_24910);
nand UO_2849 (O_2849,N_24770,N_24815);
xnor UO_2850 (O_2850,N_24938,N_24758);
and UO_2851 (O_2851,N_24867,N_24947);
nor UO_2852 (O_2852,N_24844,N_24919);
xnor UO_2853 (O_2853,N_24937,N_24925);
xnor UO_2854 (O_2854,N_24969,N_24781);
or UO_2855 (O_2855,N_24880,N_24940);
nand UO_2856 (O_2856,N_24925,N_24823);
or UO_2857 (O_2857,N_24852,N_24945);
xor UO_2858 (O_2858,N_24956,N_24886);
or UO_2859 (O_2859,N_24926,N_24998);
xnor UO_2860 (O_2860,N_24841,N_24819);
and UO_2861 (O_2861,N_24819,N_24889);
nand UO_2862 (O_2862,N_24773,N_24803);
nor UO_2863 (O_2863,N_24938,N_24833);
nand UO_2864 (O_2864,N_24924,N_24824);
nor UO_2865 (O_2865,N_24838,N_24787);
and UO_2866 (O_2866,N_24871,N_24969);
nand UO_2867 (O_2867,N_24837,N_24974);
xnor UO_2868 (O_2868,N_24907,N_24801);
nand UO_2869 (O_2869,N_24997,N_24832);
nor UO_2870 (O_2870,N_24889,N_24870);
and UO_2871 (O_2871,N_24889,N_24949);
nand UO_2872 (O_2872,N_24892,N_24932);
or UO_2873 (O_2873,N_24900,N_24776);
xnor UO_2874 (O_2874,N_24922,N_24892);
or UO_2875 (O_2875,N_24964,N_24957);
nand UO_2876 (O_2876,N_24865,N_24947);
nand UO_2877 (O_2877,N_24902,N_24765);
nor UO_2878 (O_2878,N_24920,N_24866);
xor UO_2879 (O_2879,N_24827,N_24753);
nand UO_2880 (O_2880,N_24961,N_24912);
and UO_2881 (O_2881,N_24992,N_24897);
nand UO_2882 (O_2882,N_24759,N_24789);
and UO_2883 (O_2883,N_24911,N_24752);
or UO_2884 (O_2884,N_24843,N_24857);
or UO_2885 (O_2885,N_24794,N_24915);
nor UO_2886 (O_2886,N_24817,N_24865);
nand UO_2887 (O_2887,N_24897,N_24780);
nor UO_2888 (O_2888,N_24794,N_24852);
or UO_2889 (O_2889,N_24836,N_24931);
nor UO_2890 (O_2890,N_24868,N_24783);
nand UO_2891 (O_2891,N_24860,N_24886);
xnor UO_2892 (O_2892,N_24757,N_24782);
nor UO_2893 (O_2893,N_24804,N_24982);
and UO_2894 (O_2894,N_24892,N_24832);
nand UO_2895 (O_2895,N_24907,N_24901);
and UO_2896 (O_2896,N_24961,N_24774);
xnor UO_2897 (O_2897,N_24817,N_24772);
xnor UO_2898 (O_2898,N_24971,N_24800);
xor UO_2899 (O_2899,N_24761,N_24808);
xnor UO_2900 (O_2900,N_24803,N_24760);
xnor UO_2901 (O_2901,N_24793,N_24777);
and UO_2902 (O_2902,N_24952,N_24758);
xor UO_2903 (O_2903,N_24881,N_24810);
nand UO_2904 (O_2904,N_24988,N_24810);
nor UO_2905 (O_2905,N_24852,N_24919);
xor UO_2906 (O_2906,N_24975,N_24816);
and UO_2907 (O_2907,N_24894,N_24935);
nor UO_2908 (O_2908,N_24948,N_24779);
nor UO_2909 (O_2909,N_24794,N_24773);
nor UO_2910 (O_2910,N_24865,N_24820);
and UO_2911 (O_2911,N_24890,N_24995);
or UO_2912 (O_2912,N_24783,N_24786);
xor UO_2913 (O_2913,N_24866,N_24932);
or UO_2914 (O_2914,N_24803,N_24845);
and UO_2915 (O_2915,N_24863,N_24998);
nor UO_2916 (O_2916,N_24865,N_24874);
and UO_2917 (O_2917,N_24975,N_24948);
nand UO_2918 (O_2918,N_24799,N_24866);
and UO_2919 (O_2919,N_24827,N_24956);
or UO_2920 (O_2920,N_24863,N_24953);
xor UO_2921 (O_2921,N_24920,N_24793);
nand UO_2922 (O_2922,N_24902,N_24985);
nand UO_2923 (O_2923,N_24957,N_24796);
nand UO_2924 (O_2924,N_24881,N_24859);
xor UO_2925 (O_2925,N_24939,N_24897);
and UO_2926 (O_2926,N_24968,N_24872);
or UO_2927 (O_2927,N_24998,N_24840);
xor UO_2928 (O_2928,N_24892,N_24928);
or UO_2929 (O_2929,N_24929,N_24785);
or UO_2930 (O_2930,N_24972,N_24830);
nand UO_2931 (O_2931,N_24808,N_24847);
and UO_2932 (O_2932,N_24853,N_24991);
xnor UO_2933 (O_2933,N_24805,N_24861);
or UO_2934 (O_2934,N_24976,N_24777);
nor UO_2935 (O_2935,N_24946,N_24779);
nand UO_2936 (O_2936,N_24884,N_24830);
and UO_2937 (O_2937,N_24868,N_24793);
nand UO_2938 (O_2938,N_24926,N_24994);
and UO_2939 (O_2939,N_24761,N_24832);
and UO_2940 (O_2940,N_24899,N_24815);
nor UO_2941 (O_2941,N_24794,N_24984);
nand UO_2942 (O_2942,N_24964,N_24902);
nand UO_2943 (O_2943,N_24845,N_24950);
and UO_2944 (O_2944,N_24835,N_24834);
or UO_2945 (O_2945,N_24887,N_24999);
or UO_2946 (O_2946,N_24978,N_24796);
and UO_2947 (O_2947,N_24906,N_24791);
or UO_2948 (O_2948,N_24998,N_24909);
and UO_2949 (O_2949,N_24785,N_24796);
xnor UO_2950 (O_2950,N_24798,N_24788);
nand UO_2951 (O_2951,N_24795,N_24783);
xor UO_2952 (O_2952,N_24957,N_24935);
or UO_2953 (O_2953,N_24991,N_24914);
nand UO_2954 (O_2954,N_24927,N_24906);
and UO_2955 (O_2955,N_24907,N_24883);
or UO_2956 (O_2956,N_24976,N_24981);
and UO_2957 (O_2957,N_24866,N_24793);
xnor UO_2958 (O_2958,N_24928,N_24798);
and UO_2959 (O_2959,N_24973,N_24810);
nor UO_2960 (O_2960,N_24859,N_24842);
xor UO_2961 (O_2961,N_24907,N_24838);
xnor UO_2962 (O_2962,N_24936,N_24900);
or UO_2963 (O_2963,N_24768,N_24954);
or UO_2964 (O_2964,N_24848,N_24890);
nor UO_2965 (O_2965,N_24865,N_24944);
and UO_2966 (O_2966,N_24798,N_24870);
or UO_2967 (O_2967,N_24837,N_24922);
or UO_2968 (O_2968,N_24969,N_24935);
nand UO_2969 (O_2969,N_24800,N_24813);
or UO_2970 (O_2970,N_24827,N_24921);
nand UO_2971 (O_2971,N_24803,N_24997);
nor UO_2972 (O_2972,N_24827,N_24895);
nand UO_2973 (O_2973,N_24901,N_24970);
nand UO_2974 (O_2974,N_24934,N_24925);
xnor UO_2975 (O_2975,N_24811,N_24801);
nor UO_2976 (O_2976,N_24920,N_24877);
or UO_2977 (O_2977,N_24776,N_24865);
and UO_2978 (O_2978,N_24828,N_24872);
or UO_2979 (O_2979,N_24807,N_24820);
nand UO_2980 (O_2980,N_24846,N_24901);
or UO_2981 (O_2981,N_24845,N_24827);
nor UO_2982 (O_2982,N_24901,N_24891);
and UO_2983 (O_2983,N_24899,N_24896);
and UO_2984 (O_2984,N_24836,N_24834);
and UO_2985 (O_2985,N_24784,N_24788);
xnor UO_2986 (O_2986,N_24893,N_24966);
nand UO_2987 (O_2987,N_24750,N_24875);
nand UO_2988 (O_2988,N_24793,N_24797);
nor UO_2989 (O_2989,N_24938,N_24810);
and UO_2990 (O_2990,N_24934,N_24964);
and UO_2991 (O_2991,N_24797,N_24995);
nor UO_2992 (O_2992,N_24896,N_24958);
nor UO_2993 (O_2993,N_24812,N_24935);
or UO_2994 (O_2994,N_24847,N_24810);
nand UO_2995 (O_2995,N_24815,N_24896);
or UO_2996 (O_2996,N_24762,N_24772);
or UO_2997 (O_2997,N_24784,N_24809);
nor UO_2998 (O_2998,N_24833,N_24894);
nand UO_2999 (O_2999,N_24826,N_24919);
endmodule