module basic_500_3000_500_5_levels_5xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
xor U0 (N_0,In_248,In_6);
xnor U1 (N_1,In_22,In_300);
nand U2 (N_2,In_147,In_249);
xnor U3 (N_3,In_168,In_348);
nor U4 (N_4,In_88,In_197);
nand U5 (N_5,In_74,In_241);
or U6 (N_6,In_271,In_400);
nor U7 (N_7,In_252,In_107);
or U8 (N_8,In_481,In_340);
nand U9 (N_9,In_68,In_213);
nor U10 (N_10,In_393,In_386);
xnor U11 (N_11,In_163,In_233);
xnor U12 (N_12,In_414,In_32);
xor U13 (N_13,In_488,In_417);
and U14 (N_14,In_209,In_343);
nand U15 (N_15,In_102,In_442);
or U16 (N_16,In_404,In_322);
or U17 (N_17,In_64,In_367);
nand U18 (N_18,In_302,In_440);
nor U19 (N_19,In_260,In_200);
nor U20 (N_20,In_84,In_114);
nor U21 (N_21,In_287,In_472);
nor U22 (N_22,In_89,In_10);
or U23 (N_23,In_27,In_13);
nand U24 (N_24,In_146,In_336);
nand U25 (N_25,In_191,In_494);
and U26 (N_26,In_223,In_333);
nor U27 (N_27,In_126,In_177);
or U28 (N_28,In_338,In_123);
or U29 (N_29,In_446,In_327);
and U30 (N_30,In_212,In_480);
nand U31 (N_31,In_313,In_101);
or U32 (N_32,In_100,In_144);
and U33 (N_33,In_77,In_479);
xor U34 (N_34,In_225,In_329);
nor U35 (N_35,In_405,In_31);
and U36 (N_36,In_272,In_434);
nand U37 (N_37,In_462,In_162);
or U38 (N_38,In_167,In_58);
nor U39 (N_39,In_80,In_172);
nand U40 (N_40,In_443,In_20);
and U41 (N_41,In_351,In_188);
and U42 (N_42,In_304,In_474);
nand U43 (N_43,In_321,In_16);
nand U44 (N_44,In_421,In_128);
nor U45 (N_45,In_411,In_326);
nand U46 (N_46,In_280,In_360);
and U47 (N_47,In_459,In_425);
and U48 (N_48,In_83,In_237);
nor U49 (N_49,In_268,In_457);
or U50 (N_50,In_218,In_56);
nor U51 (N_51,In_307,In_175);
nand U52 (N_52,In_298,In_432);
xnor U53 (N_53,In_232,In_401);
nand U54 (N_54,In_458,In_49);
and U55 (N_55,In_339,In_52);
nor U56 (N_56,In_255,In_57);
and U57 (N_57,In_246,In_239);
xor U58 (N_58,In_412,In_394);
or U59 (N_59,In_427,In_315);
nand U60 (N_60,In_176,In_62);
and U61 (N_61,In_357,In_452);
nor U62 (N_62,In_413,In_251);
and U63 (N_63,In_433,In_475);
or U64 (N_64,In_464,In_497);
nand U65 (N_65,In_51,In_361);
or U66 (N_66,In_354,In_194);
and U67 (N_67,In_468,In_410);
or U68 (N_68,In_85,In_341);
and U69 (N_69,In_15,In_384);
or U70 (N_70,In_186,In_199);
or U71 (N_71,In_44,In_262);
and U72 (N_72,In_296,In_355);
nor U73 (N_73,In_63,In_403);
nor U74 (N_74,In_283,In_173);
and U75 (N_75,In_495,In_422);
nor U76 (N_76,In_285,In_390);
nand U77 (N_77,In_314,In_149);
or U78 (N_78,In_439,In_39);
or U79 (N_79,In_160,In_184);
nand U80 (N_80,In_30,In_350);
or U81 (N_81,In_129,In_324);
nor U82 (N_82,In_203,In_109);
nand U83 (N_83,In_156,In_273);
or U84 (N_84,In_3,In_353);
nand U85 (N_85,In_483,In_26);
nand U86 (N_86,In_460,In_152);
and U87 (N_87,In_435,In_290);
xnor U88 (N_88,In_36,In_171);
and U89 (N_89,In_112,In_208);
nand U90 (N_90,In_150,In_235);
xnor U91 (N_91,In_37,In_189);
nand U92 (N_92,In_358,In_75);
nor U93 (N_93,In_312,In_447);
and U94 (N_94,In_378,In_8);
nor U95 (N_95,In_202,In_356);
and U96 (N_96,In_477,In_116);
nor U97 (N_97,In_430,In_148);
or U98 (N_98,In_164,In_281);
nand U99 (N_99,In_473,In_375);
and U100 (N_100,In_261,In_206);
or U101 (N_101,In_226,In_115);
nor U102 (N_102,In_242,In_492);
or U103 (N_103,In_106,In_61);
nor U104 (N_104,In_14,In_139);
and U105 (N_105,In_135,In_448);
xor U106 (N_106,In_122,In_381);
nand U107 (N_107,In_337,In_47);
and U108 (N_108,In_486,In_279);
nand U109 (N_109,In_216,In_402);
and U110 (N_110,In_125,In_471);
and U111 (N_111,In_157,In_69);
or U112 (N_112,In_141,In_143);
and U113 (N_113,In_441,In_120);
and U114 (N_114,In_65,In_382);
and U115 (N_115,In_295,In_215);
nand U116 (N_116,In_154,In_470);
nor U117 (N_117,In_220,In_29);
nand U118 (N_118,In_247,In_166);
nor U119 (N_119,In_111,In_396);
and U120 (N_120,In_325,In_124);
nor U121 (N_121,In_119,In_245);
or U122 (N_122,In_418,In_19);
nand U123 (N_123,In_436,In_190);
or U124 (N_124,In_169,In_72);
nand U125 (N_125,In_365,In_376);
and U126 (N_126,In_93,In_210);
xor U127 (N_127,In_294,In_145);
nor U128 (N_128,In_70,In_136);
nor U129 (N_129,In_250,In_416);
xor U130 (N_130,In_289,In_121);
xnor U131 (N_131,In_347,In_159);
xnor U132 (N_132,In_7,In_227);
nand U133 (N_133,In_491,In_383);
nor U134 (N_134,In_11,In_406);
or U135 (N_135,In_269,In_444);
and U136 (N_136,In_317,In_415);
nor U137 (N_137,In_346,In_385);
or U138 (N_138,In_234,In_204);
and U139 (N_139,In_222,In_258);
xor U140 (N_140,In_359,In_224);
and U141 (N_141,In_363,In_437);
nor U142 (N_142,In_463,In_478);
nor U143 (N_143,In_455,In_399);
or U144 (N_144,In_40,In_236);
nor U145 (N_145,In_221,In_257);
or U146 (N_146,In_140,In_345);
nor U147 (N_147,In_398,In_55);
and U148 (N_148,In_332,In_342);
or U149 (N_149,In_370,In_97);
or U150 (N_150,In_466,In_366);
and U151 (N_151,In_277,In_35);
or U152 (N_152,In_498,In_38);
xor U153 (N_153,In_482,In_12);
xnor U154 (N_154,In_161,In_217);
or U155 (N_155,In_110,In_301);
nand U156 (N_156,In_420,In_243);
nand U157 (N_157,In_240,In_132);
and U158 (N_158,In_201,In_305);
and U159 (N_159,In_374,In_87);
xnor U160 (N_160,In_485,In_211);
or U161 (N_161,In_362,In_82);
nand U162 (N_162,In_292,In_253);
and U163 (N_163,In_388,In_306);
and U164 (N_164,In_207,In_45);
xnor U165 (N_165,In_451,In_490);
or U166 (N_166,In_429,In_91);
nor U167 (N_167,In_465,In_1);
nand U168 (N_168,In_407,In_158);
xnor U169 (N_169,In_377,In_219);
or U170 (N_170,In_228,In_489);
and U171 (N_171,In_142,In_5);
or U172 (N_172,In_76,In_183);
nand U173 (N_173,In_259,In_454);
nand U174 (N_174,In_66,In_349);
and U175 (N_175,In_60,In_344);
or U176 (N_176,In_86,In_487);
xnor U177 (N_177,In_395,In_192);
or U178 (N_178,In_270,In_449);
nand U179 (N_179,In_42,In_331);
nor U180 (N_180,In_476,In_73);
nor U181 (N_181,In_310,In_276);
nand U182 (N_182,In_153,In_431);
or U183 (N_183,In_170,In_330);
nand U184 (N_184,In_2,In_92);
or U185 (N_185,In_130,In_379);
and U186 (N_186,In_373,In_34);
and U187 (N_187,In_284,In_81);
nor U188 (N_188,In_364,In_323);
and U189 (N_189,In_67,In_288);
nand U190 (N_190,In_469,In_127);
nor U191 (N_191,In_335,In_181);
and U192 (N_192,In_266,In_320);
nor U193 (N_193,In_182,In_180);
and U194 (N_194,In_275,In_461);
and U195 (N_195,In_371,In_4);
or U196 (N_196,In_178,In_17);
and U197 (N_197,In_291,In_231);
nor U198 (N_198,In_0,In_205);
or U199 (N_199,In_445,In_28);
nand U200 (N_200,In_185,In_264);
and U201 (N_201,In_24,In_419);
or U202 (N_202,In_174,In_18);
and U203 (N_203,In_368,In_450);
nor U204 (N_204,In_21,In_263);
nor U205 (N_205,In_138,In_423);
and U206 (N_206,In_426,In_380);
nor U207 (N_207,In_408,In_155);
and U208 (N_208,In_352,In_267);
nor U209 (N_209,In_195,In_456);
xnor U210 (N_210,In_230,In_95);
nor U211 (N_211,In_94,In_387);
xor U212 (N_212,In_103,In_293);
and U213 (N_213,In_198,In_79);
nor U214 (N_214,In_96,In_274);
nor U215 (N_215,In_229,In_244);
nor U216 (N_216,In_282,In_334);
and U217 (N_217,In_117,In_499);
or U218 (N_218,In_98,In_179);
and U219 (N_219,In_108,In_113);
nor U220 (N_220,In_397,In_286);
nand U221 (N_221,In_134,In_118);
or U222 (N_222,In_328,In_196);
nor U223 (N_223,In_428,In_90);
and U224 (N_224,In_9,In_78);
or U225 (N_225,In_33,In_214);
and U226 (N_226,In_99,In_369);
nand U227 (N_227,In_59,In_25);
xnor U228 (N_228,In_496,In_23);
and U229 (N_229,In_53,In_43);
nand U230 (N_230,In_297,In_467);
and U231 (N_231,In_309,In_318);
nor U232 (N_232,In_303,In_193);
nor U233 (N_233,In_238,In_453);
nor U234 (N_234,In_316,In_104);
and U235 (N_235,In_105,In_256);
xor U236 (N_236,In_187,In_48);
nand U237 (N_237,In_46,In_54);
and U238 (N_238,In_50,In_493);
nand U239 (N_239,In_133,In_151);
nor U240 (N_240,In_311,In_484);
nand U241 (N_241,In_308,In_254);
and U242 (N_242,In_71,In_131);
nand U243 (N_243,In_165,In_278);
nand U244 (N_244,In_391,In_372);
or U245 (N_245,In_265,In_424);
xor U246 (N_246,In_319,In_389);
nand U247 (N_247,In_137,In_409);
xnor U248 (N_248,In_438,In_392);
nor U249 (N_249,In_299,In_41);
and U250 (N_250,In_222,In_93);
and U251 (N_251,In_84,In_215);
nor U252 (N_252,In_77,In_237);
nand U253 (N_253,In_58,In_96);
nor U254 (N_254,In_277,In_57);
nand U255 (N_255,In_23,In_117);
nand U256 (N_256,In_15,In_60);
nand U257 (N_257,In_48,In_353);
or U258 (N_258,In_364,In_2);
nor U259 (N_259,In_167,In_286);
or U260 (N_260,In_415,In_100);
and U261 (N_261,In_297,In_273);
nor U262 (N_262,In_368,In_253);
nand U263 (N_263,In_308,In_474);
and U264 (N_264,In_218,In_97);
or U265 (N_265,In_388,In_450);
nor U266 (N_266,In_9,In_186);
and U267 (N_267,In_110,In_399);
nor U268 (N_268,In_125,In_491);
and U269 (N_269,In_64,In_5);
nor U270 (N_270,In_426,In_293);
xor U271 (N_271,In_468,In_229);
and U272 (N_272,In_203,In_11);
nand U273 (N_273,In_172,In_344);
nand U274 (N_274,In_259,In_400);
nand U275 (N_275,In_497,In_57);
nor U276 (N_276,In_483,In_286);
nor U277 (N_277,In_38,In_430);
and U278 (N_278,In_271,In_346);
and U279 (N_279,In_386,In_334);
or U280 (N_280,In_430,In_456);
xnor U281 (N_281,In_113,In_271);
nand U282 (N_282,In_114,In_168);
and U283 (N_283,In_338,In_119);
and U284 (N_284,In_148,In_422);
or U285 (N_285,In_242,In_261);
xnor U286 (N_286,In_33,In_323);
xor U287 (N_287,In_491,In_149);
nand U288 (N_288,In_244,In_145);
or U289 (N_289,In_447,In_240);
or U290 (N_290,In_299,In_256);
or U291 (N_291,In_153,In_475);
and U292 (N_292,In_99,In_129);
nand U293 (N_293,In_294,In_125);
and U294 (N_294,In_425,In_411);
or U295 (N_295,In_228,In_341);
and U296 (N_296,In_122,In_352);
xnor U297 (N_297,In_74,In_161);
xnor U298 (N_298,In_255,In_385);
or U299 (N_299,In_158,In_43);
or U300 (N_300,In_462,In_61);
xnor U301 (N_301,In_370,In_298);
nand U302 (N_302,In_224,In_407);
nor U303 (N_303,In_334,In_300);
nand U304 (N_304,In_157,In_380);
and U305 (N_305,In_433,In_232);
nor U306 (N_306,In_39,In_364);
nor U307 (N_307,In_477,In_99);
nand U308 (N_308,In_339,In_89);
or U309 (N_309,In_223,In_468);
nor U310 (N_310,In_346,In_184);
nor U311 (N_311,In_200,In_331);
xor U312 (N_312,In_382,In_439);
or U313 (N_313,In_34,In_366);
nand U314 (N_314,In_226,In_19);
and U315 (N_315,In_47,In_53);
or U316 (N_316,In_186,In_59);
nor U317 (N_317,In_313,In_277);
nand U318 (N_318,In_372,In_217);
and U319 (N_319,In_294,In_335);
and U320 (N_320,In_456,In_116);
or U321 (N_321,In_465,In_142);
or U322 (N_322,In_263,In_366);
nand U323 (N_323,In_34,In_6);
or U324 (N_324,In_342,In_291);
or U325 (N_325,In_457,In_58);
or U326 (N_326,In_216,In_206);
or U327 (N_327,In_468,In_368);
nand U328 (N_328,In_202,In_52);
and U329 (N_329,In_210,In_330);
nand U330 (N_330,In_376,In_203);
or U331 (N_331,In_255,In_424);
nand U332 (N_332,In_20,In_470);
or U333 (N_333,In_469,In_344);
xnor U334 (N_334,In_56,In_322);
or U335 (N_335,In_118,In_66);
nor U336 (N_336,In_387,In_225);
nor U337 (N_337,In_44,In_186);
nand U338 (N_338,In_384,In_301);
nor U339 (N_339,In_268,In_446);
xor U340 (N_340,In_395,In_154);
and U341 (N_341,In_440,In_106);
xnor U342 (N_342,In_211,In_319);
nor U343 (N_343,In_5,In_289);
nor U344 (N_344,In_307,In_39);
or U345 (N_345,In_317,In_73);
and U346 (N_346,In_43,In_175);
xnor U347 (N_347,In_428,In_415);
or U348 (N_348,In_312,In_446);
nor U349 (N_349,In_466,In_128);
and U350 (N_350,In_66,In_386);
xnor U351 (N_351,In_19,In_246);
nor U352 (N_352,In_479,In_420);
nor U353 (N_353,In_258,In_265);
nor U354 (N_354,In_180,In_158);
or U355 (N_355,In_74,In_174);
and U356 (N_356,In_81,In_391);
or U357 (N_357,In_67,In_282);
or U358 (N_358,In_178,In_219);
xor U359 (N_359,In_334,In_167);
xor U360 (N_360,In_362,In_157);
and U361 (N_361,In_450,In_62);
nor U362 (N_362,In_446,In_176);
xor U363 (N_363,In_446,In_123);
or U364 (N_364,In_215,In_378);
nor U365 (N_365,In_57,In_168);
or U366 (N_366,In_259,In_240);
nor U367 (N_367,In_189,In_201);
or U368 (N_368,In_180,In_310);
or U369 (N_369,In_459,In_22);
and U370 (N_370,In_337,In_10);
and U371 (N_371,In_161,In_182);
nor U372 (N_372,In_391,In_78);
and U373 (N_373,In_382,In_229);
or U374 (N_374,In_395,In_405);
nor U375 (N_375,In_308,In_202);
or U376 (N_376,In_406,In_317);
xnor U377 (N_377,In_489,In_329);
or U378 (N_378,In_192,In_266);
and U379 (N_379,In_432,In_373);
nand U380 (N_380,In_400,In_108);
nor U381 (N_381,In_172,In_290);
nor U382 (N_382,In_26,In_408);
and U383 (N_383,In_271,In_263);
and U384 (N_384,In_385,In_363);
nand U385 (N_385,In_332,In_310);
nor U386 (N_386,In_480,In_194);
nor U387 (N_387,In_333,In_55);
and U388 (N_388,In_309,In_41);
and U389 (N_389,In_195,In_162);
nand U390 (N_390,In_486,In_7);
nand U391 (N_391,In_276,In_365);
and U392 (N_392,In_479,In_480);
nor U393 (N_393,In_496,In_106);
and U394 (N_394,In_43,In_371);
xnor U395 (N_395,In_299,In_380);
nand U396 (N_396,In_172,In_154);
nor U397 (N_397,In_159,In_195);
nor U398 (N_398,In_332,In_199);
and U399 (N_399,In_232,In_167);
nor U400 (N_400,In_401,In_442);
nand U401 (N_401,In_61,In_6);
or U402 (N_402,In_153,In_137);
and U403 (N_403,In_411,In_222);
nand U404 (N_404,In_339,In_390);
nor U405 (N_405,In_486,In_121);
nand U406 (N_406,In_280,In_103);
and U407 (N_407,In_433,In_434);
or U408 (N_408,In_356,In_390);
and U409 (N_409,In_296,In_297);
or U410 (N_410,In_81,In_249);
or U411 (N_411,In_201,In_464);
nor U412 (N_412,In_317,In_134);
nand U413 (N_413,In_109,In_240);
and U414 (N_414,In_399,In_281);
nand U415 (N_415,In_300,In_349);
nor U416 (N_416,In_334,In_186);
or U417 (N_417,In_21,In_251);
nand U418 (N_418,In_388,In_296);
or U419 (N_419,In_327,In_11);
and U420 (N_420,In_197,In_276);
nor U421 (N_421,In_292,In_472);
nand U422 (N_422,In_225,In_227);
xor U423 (N_423,In_35,In_135);
and U424 (N_424,In_5,In_45);
xnor U425 (N_425,In_196,In_36);
and U426 (N_426,In_328,In_244);
and U427 (N_427,In_432,In_290);
or U428 (N_428,In_138,In_454);
nand U429 (N_429,In_241,In_216);
xor U430 (N_430,In_423,In_246);
or U431 (N_431,In_437,In_59);
and U432 (N_432,In_38,In_148);
nand U433 (N_433,In_418,In_260);
and U434 (N_434,In_217,In_393);
nor U435 (N_435,In_350,In_497);
or U436 (N_436,In_312,In_371);
nor U437 (N_437,In_375,In_496);
and U438 (N_438,In_39,In_55);
nor U439 (N_439,In_174,In_130);
or U440 (N_440,In_388,In_464);
and U441 (N_441,In_134,In_227);
nor U442 (N_442,In_351,In_249);
nor U443 (N_443,In_313,In_251);
nor U444 (N_444,In_118,In_133);
and U445 (N_445,In_111,In_112);
xnor U446 (N_446,In_338,In_458);
nor U447 (N_447,In_428,In_432);
or U448 (N_448,In_291,In_463);
and U449 (N_449,In_484,In_250);
xnor U450 (N_450,In_464,In_297);
or U451 (N_451,In_101,In_438);
nand U452 (N_452,In_330,In_363);
nor U453 (N_453,In_459,In_229);
or U454 (N_454,In_134,In_17);
nor U455 (N_455,In_26,In_52);
nor U456 (N_456,In_206,In_265);
or U457 (N_457,In_180,In_400);
nor U458 (N_458,In_24,In_43);
and U459 (N_459,In_321,In_134);
or U460 (N_460,In_19,In_161);
or U461 (N_461,In_100,In_422);
xnor U462 (N_462,In_82,In_322);
nor U463 (N_463,In_11,In_120);
nand U464 (N_464,In_0,In_405);
xor U465 (N_465,In_83,In_239);
nor U466 (N_466,In_317,In_120);
or U467 (N_467,In_202,In_163);
or U468 (N_468,In_95,In_409);
xnor U469 (N_469,In_170,In_355);
and U470 (N_470,In_27,In_54);
xor U471 (N_471,In_198,In_281);
nor U472 (N_472,In_99,In_117);
nand U473 (N_473,In_464,In_76);
and U474 (N_474,In_488,In_278);
nand U475 (N_475,In_323,In_74);
and U476 (N_476,In_287,In_248);
xor U477 (N_477,In_93,In_297);
and U478 (N_478,In_96,In_136);
xnor U479 (N_479,In_139,In_59);
and U480 (N_480,In_27,In_379);
nor U481 (N_481,In_215,In_334);
xor U482 (N_482,In_336,In_208);
nand U483 (N_483,In_135,In_329);
nand U484 (N_484,In_399,In_153);
nand U485 (N_485,In_264,In_159);
nor U486 (N_486,In_232,In_217);
xor U487 (N_487,In_406,In_175);
nor U488 (N_488,In_473,In_435);
nand U489 (N_489,In_251,In_441);
or U490 (N_490,In_243,In_143);
nand U491 (N_491,In_135,In_161);
and U492 (N_492,In_242,In_233);
nand U493 (N_493,In_288,In_102);
nand U494 (N_494,In_415,In_36);
nor U495 (N_495,In_81,In_208);
or U496 (N_496,In_248,In_422);
nand U497 (N_497,In_42,In_3);
nor U498 (N_498,In_41,In_482);
nand U499 (N_499,In_158,In_214);
and U500 (N_500,In_263,In_411);
and U501 (N_501,In_163,In_286);
nand U502 (N_502,In_414,In_176);
and U503 (N_503,In_120,In_106);
and U504 (N_504,In_146,In_141);
and U505 (N_505,In_300,In_123);
and U506 (N_506,In_344,In_26);
xnor U507 (N_507,In_282,In_111);
nor U508 (N_508,In_161,In_38);
xnor U509 (N_509,In_419,In_174);
nand U510 (N_510,In_449,In_485);
and U511 (N_511,In_406,In_58);
and U512 (N_512,In_201,In_236);
nor U513 (N_513,In_125,In_36);
nand U514 (N_514,In_162,In_343);
nand U515 (N_515,In_40,In_381);
or U516 (N_516,In_207,In_276);
xnor U517 (N_517,In_201,In_192);
or U518 (N_518,In_239,In_274);
or U519 (N_519,In_354,In_344);
or U520 (N_520,In_430,In_245);
nand U521 (N_521,In_114,In_463);
or U522 (N_522,In_170,In_375);
or U523 (N_523,In_93,In_298);
and U524 (N_524,In_4,In_61);
nor U525 (N_525,In_116,In_58);
nor U526 (N_526,In_353,In_213);
or U527 (N_527,In_67,In_187);
nor U528 (N_528,In_205,In_319);
xnor U529 (N_529,In_336,In_280);
nand U530 (N_530,In_310,In_383);
nand U531 (N_531,In_199,In_281);
nand U532 (N_532,In_46,In_322);
nor U533 (N_533,In_438,In_445);
nand U534 (N_534,In_175,In_7);
nor U535 (N_535,In_250,In_257);
xnor U536 (N_536,In_170,In_426);
nor U537 (N_537,In_390,In_54);
or U538 (N_538,In_354,In_176);
nand U539 (N_539,In_58,In_319);
nor U540 (N_540,In_153,In_70);
and U541 (N_541,In_123,In_148);
or U542 (N_542,In_471,In_238);
nand U543 (N_543,In_117,In_476);
nor U544 (N_544,In_472,In_129);
nand U545 (N_545,In_204,In_179);
and U546 (N_546,In_241,In_304);
nand U547 (N_547,In_95,In_110);
and U548 (N_548,In_36,In_390);
nand U549 (N_549,In_91,In_382);
and U550 (N_550,In_0,In_462);
or U551 (N_551,In_348,In_360);
or U552 (N_552,In_367,In_364);
and U553 (N_553,In_284,In_338);
or U554 (N_554,In_267,In_49);
or U555 (N_555,In_146,In_100);
nor U556 (N_556,In_218,In_350);
xor U557 (N_557,In_119,In_81);
nor U558 (N_558,In_226,In_314);
nor U559 (N_559,In_25,In_309);
and U560 (N_560,In_221,In_281);
or U561 (N_561,In_229,In_37);
and U562 (N_562,In_184,In_362);
and U563 (N_563,In_233,In_322);
xor U564 (N_564,In_38,In_323);
nand U565 (N_565,In_52,In_446);
or U566 (N_566,In_461,In_225);
and U567 (N_567,In_43,In_485);
and U568 (N_568,In_254,In_380);
and U569 (N_569,In_178,In_30);
and U570 (N_570,In_221,In_237);
nand U571 (N_571,In_278,In_78);
and U572 (N_572,In_369,In_323);
nor U573 (N_573,In_271,In_335);
or U574 (N_574,In_319,In_381);
and U575 (N_575,In_294,In_366);
or U576 (N_576,In_149,In_269);
nor U577 (N_577,In_63,In_362);
nand U578 (N_578,In_6,In_451);
or U579 (N_579,In_480,In_409);
and U580 (N_580,In_5,In_493);
nand U581 (N_581,In_495,In_147);
nor U582 (N_582,In_317,In_263);
xnor U583 (N_583,In_50,In_359);
and U584 (N_584,In_282,In_81);
nand U585 (N_585,In_268,In_407);
and U586 (N_586,In_240,In_284);
nor U587 (N_587,In_485,In_25);
xor U588 (N_588,In_194,In_404);
nor U589 (N_589,In_293,In_411);
nor U590 (N_590,In_106,In_201);
or U591 (N_591,In_3,In_476);
and U592 (N_592,In_480,In_378);
nor U593 (N_593,In_363,In_2);
nand U594 (N_594,In_211,In_150);
nand U595 (N_595,In_69,In_365);
or U596 (N_596,In_156,In_363);
nor U597 (N_597,In_458,In_259);
xor U598 (N_598,In_424,In_140);
and U599 (N_599,In_365,In_6);
and U600 (N_600,N_342,N_202);
nor U601 (N_601,N_251,N_92);
and U602 (N_602,N_599,N_417);
nand U603 (N_603,N_255,N_381);
or U604 (N_604,N_139,N_332);
nand U605 (N_605,N_545,N_477);
nor U606 (N_606,N_490,N_206);
nor U607 (N_607,N_243,N_248);
and U608 (N_608,N_373,N_108);
and U609 (N_609,N_393,N_355);
or U610 (N_610,N_274,N_386);
and U611 (N_611,N_440,N_569);
nor U612 (N_612,N_285,N_171);
or U613 (N_613,N_264,N_44);
nand U614 (N_614,N_211,N_228);
xnor U615 (N_615,N_90,N_130);
and U616 (N_616,N_563,N_508);
nor U617 (N_617,N_320,N_252);
or U618 (N_618,N_270,N_542);
nand U619 (N_619,N_394,N_395);
nand U620 (N_620,N_256,N_113);
nand U621 (N_621,N_471,N_389);
xor U622 (N_622,N_261,N_297);
nor U623 (N_623,N_445,N_46);
nand U624 (N_624,N_121,N_187);
or U625 (N_625,N_272,N_554);
nand U626 (N_626,N_143,N_539);
and U627 (N_627,N_189,N_109);
or U628 (N_628,N_167,N_402);
nor U629 (N_629,N_472,N_469);
and U630 (N_630,N_336,N_593);
or U631 (N_631,N_6,N_456);
nand U632 (N_632,N_64,N_72);
nand U633 (N_633,N_154,N_492);
and U634 (N_634,N_106,N_334);
and U635 (N_635,N_287,N_78);
and U636 (N_636,N_463,N_147);
and U637 (N_637,N_459,N_458);
nand U638 (N_638,N_565,N_122);
nor U639 (N_639,N_429,N_398);
nand U640 (N_640,N_299,N_521);
nor U641 (N_641,N_451,N_348);
and U642 (N_642,N_260,N_371);
and U643 (N_643,N_250,N_165);
or U644 (N_644,N_128,N_376);
nor U645 (N_645,N_546,N_282);
nand U646 (N_646,N_150,N_367);
and U647 (N_647,N_42,N_192);
nand U648 (N_648,N_68,N_80);
nor U649 (N_649,N_427,N_238);
and U650 (N_650,N_450,N_89);
and U651 (N_651,N_303,N_400);
nor U652 (N_652,N_486,N_49);
nand U653 (N_653,N_170,N_127);
nor U654 (N_654,N_123,N_411);
nand U655 (N_655,N_273,N_333);
and U656 (N_656,N_194,N_421);
nand U657 (N_657,N_489,N_315);
or U658 (N_658,N_4,N_511);
and U659 (N_659,N_153,N_281);
or U660 (N_660,N_319,N_40);
or U661 (N_661,N_77,N_436);
nor U662 (N_662,N_164,N_549);
nor U663 (N_663,N_105,N_91);
xor U664 (N_664,N_364,N_254);
nor U665 (N_665,N_95,N_73);
or U666 (N_666,N_378,N_30);
or U667 (N_667,N_596,N_71);
nor U668 (N_668,N_125,N_218);
nor U669 (N_669,N_535,N_505);
or U670 (N_670,N_326,N_36);
or U671 (N_671,N_488,N_203);
or U672 (N_672,N_96,N_156);
or U673 (N_673,N_135,N_263);
xor U674 (N_674,N_369,N_117);
or U675 (N_675,N_31,N_305);
nor U676 (N_676,N_536,N_406);
nand U677 (N_677,N_45,N_577);
and U678 (N_678,N_144,N_54);
or U679 (N_679,N_559,N_443);
nand U680 (N_680,N_26,N_560);
and U681 (N_681,N_83,N_418);
or U682 (N_682,N_374,N_384);
or U683 (N_683,N_561,N_357);
nor U684 (N_684,N_184,N_541);
and U685 (N_685,N_119,N_358);
xnor U686 (N_686,N_479,N_460);
and U687 (N_687,N_335,N_65);
or U688 (N_688,N_528,N_32);
and U689 (N_689,N_94,N_57);
and U690 (N_690,N_516,N_157);
and U691 (N_691,N_527,N_75);
and U692 (N_692,N_506,N_253);
and U693 (N_693,N_553,N_454);
xor U694 (N_694,N_586,N_377);
nor U695 (N_695,N_216,N_302);
and U696 (N_696,N_1,N_387);
nor U697 (N_697,N_5,N_99);
or U698 (N_698,N_175,N_391);
and U699 (N_699,N_221,N_503);
nor U700 (N_700,N_414,N_268);
or U701 (N_701,N_257,N_465);
xor U702 (N_702,N_115,N_435);
and U703 (N_703,N_455,N_224);
or U704 (N_704,N_292,N_590);
or U705 (N_705,N_431,N_461);
nand U706 (N_706,N_581,N_229);
nor U707 (N_707,N_491,N_310);
and U708 (N_708,N_368,N_370);
or U709 (N_709,N_543,N_12);
xnor U710 (N_710,N_415,N_19);
or U711 (N_711,N_86,N_118);
and U712 (N_712,N_284,N_301);
nand U713 (N_713,N_316,N_317);
nor U714 (N_714,N_512,N_209);
or U715 (N_715,N_448,N_39);
nand U716 (N_716,N_339,N_129);
or U717 (N_717,N_321,N_304);
or U718 (N_718,N_138,N_571);
nand U719 (N_719,N_562,N_37);
nand U720 (N_720,N_379,N_25);
nand U721 (N_721,N_499,N_396);
nand U722 (N_722,N_529,N_227);
and U723 (N_723,N_582,N_483);
xnor U724 (N_724,N_237,N_312);
and U725 (N_725,N_74,N_314);
nand U726 (N_726,N_588,N_169);
or U727 (N_727,N_351,N_515);
and U728 (N_728,N_446,N_331);
or U729 (N_729,N_585,N_425);
and U730 (N_730,N_484,N_423);
nand U731 (N_731,N_311,N_513);
and U732 (N_732,N_204,N_354);
nor U733 (N_733,N_0,N_330);
nand U734 (N_734,N_525,N_519);
or U735 (N_735,N_557,N_61);
nor U736 (N_736,N_361,N_522);
and U737 (N_737,N_579,N_114);
and U738 (N_738,N_85,N_234);
and U739 (N_739,N_344,N_350);
or U740 (N_740,N_592,N_430);
or U741 (N_741,N_172,N_185);
or U742 (N_742,N_176,N_15);
nor U743 (N_743,N_168,N_173);
nand U744 (N_744,N_195,N_244);
nor U745 (N_745,N_28,N_352);
or U746 (N_746,N_152,N_308);
nand U747 (N_747,N_21,N_84);
nand U748 (N_748,N_533,N_27);
or U749 (N_749,N_133,N_322);
nand U750 (N_750,N_294,N_20);
and U751 (N_751,N_145,N_134);
nor U752 (N_752,N_178,N_518);
nor U753 (N_753,N_551,N_56);
nand U754 (N_754,N_382,N_43);
or U755 (N_755,N_366,N_442);
or U756 (N_756,N_517,N_293);
and U757 (N_757,N_7,N_208);
nand U758 (N_758,N_530,N_199);
nor U759 (N_759,N_464,N_179);
and U760 (N_760,N_267,N_69);
nor U761 (N_761,N_29,N_290);
xnor U762 (N_762,N_81,N_365);
or U763 (N_763,N_300,N_307);
nand U764 (N_764,N_52,N_93);
or U765 (N_765,N_385,N_403);
nor U766 (N_766,N_112,N_404);
nor U767 (N_767,N_309,N_452);
nand U768 (N_768,N_475,N_524);
xor U769 (N_769,N_580,N_481);
or U770 (N_770,N_276,N_82);
nor U771 (N_771,N_444,N_555);
nand U772 (N_772,N_23,N_120);
nor U773 (N_773,N_572,N_259);
or U774 (N_774,N_584,N_438);
and U775 (N_775,N_556,N_502);
nor U776 (N_776,N_495,N_102);
nand U777 (N_777,N_498,N_63);
nor U778 (N_778,N_558,N_258);
and U779 (N_779,N_131,N_424);
and U780 (N_780,N_242,N_18);
or U781 (N_781,N_59,N_548);
nand U782 (N_782,N_279,N_283);
nand U783 (N_783,N_507,N_532);
or U784 (N_784,N_589,N_598);
nand U785 (N_785,N_576,N_509);
or U786 (N_786,N_420,N_329);
xnor U787 (N_787,N_34,N_494);
nor U788 (N_788,N_497,N_207);
or U789 (N_789,N_182,N_286);
nor U790 (N_790,N_531,N_70);
xor U791 (N_791,N_269,N_24);
nand U792 (N_792,N_473,N_235);
or U793 (N_793,N_573,N_3);
nand U794 (N_794,N_98,N_186);
or U795 (N_795,N_480,N_514);
nor U796 (N_796,N_289,N_47);
and U797 (N_797,N_587,N_163);
or U798 (N_798,N_233,N_22);
nand U799 (N_799,N_447,N_67);
nand U800 (N_800,N_566,N_466);
and U801 (N_801,N_13,N_280);
nand U802 (N_802,N_564,N_574);
nor U803 (N_803,N_110,N_197);
or U804 (N_804,N_50,N_428);
or U805 (N_805,N_196,N_104);
or U806 (N_806,N_526,N_200);
xor U807 (N_807,N_422,N_328);
or U808 (N_808,N_457,N_213);
or U809 (N_809,N_79,N_485);
nor U810 (N_810,N_180,N_10);
or U811 (N_811,N_338,N_594);
nand U812 (N_812,N_222,N_296);
and U813 (N_813,N_467,N_17);
xor U814 (N_814,N_232,N_340);
and U815 (N_815,N_226,N_583);
nor U816 (N_816,N_439,N_405);
nor U817 (N_817,N_155,N_2);
nor U818 (N_818,N_159,N_388);
nor U819 (N_819,N_552,N_107);
and U820 (N_820,N_38,N_212);
xnor U821 (N_821,N_162,N_160);
xor U822 (N_822,N_158,N_550);
nor U823 (N_823,N_223,N_520);
and U824 (N_824,N_407,N_188);
xnor U825 (N_825,N_575,N_360);
and U826 (N_826,N_409,N_408);
xnor U827 (N_827,N_66,N_327);
or U828 (N_828,N_597,N_537);
nor U829 (N_829,N_240,N_181);
and U830 (N_830,N_399,N_441);
nor U831 (N_831,N_346,N_230);
and U832 (N_832,N_337,N_124);
nor U833 (N_833,N_51,N_141);
nor U834 (N_834,N_220,N_214);
nor U835 (N_835,N_501,N_136);
or U836 (N_836,N_48,N_570);
and U837 (N_837,N_547,N_277);
xnor U838 (N_838,N_397,N_193);
or U839 (N_839,N_380,N_591);
or U840 (N_840,N_433,N_500);
or U841 (N_841,N_298,N_595);
xor U842 (N_842,N_58,N_247);
nor U843 (N_843,N_375,N_60);
nor U844 (N_844,N_217,N_151);
or U845 (N_845,N_271,N_177);
nand U846 (N_846,N_462,N_245);
xnor U847 (N_847,N_246,N_219);
or U848 (N_848,N_190,N_14);
and U849 (N_849,N_205,N_149);
and U850 (N_850,N_11,N_62);
and U851 (N_851,N_359,N_356);
nor U852 (N_852,N_201,N_568);
and U853 (N_853,N_413,N_210);
or U854 (N_854,N_236,N_33);
xor U855 (N_855,N_53,N_410);
nor U856 (N_856,N_324,N_146);
or U857 (N_857,N_278,N_510);
nand U858 (N_858,N_111,N_183);
xor U859 (N_859,N_9,N_87);
nor U860 (N_860,N_241,N_137);
and U861 (N_861,N_496,N_363);
nor U862 (N_862,N_437,N_76);
nand U863 (N_863,N_504,N_493);
or U864 (N_864,N_148,N_372);
nand U865 (N_865,N_215,N_362);
nand U866 (N_866,N_434,N_166);
nor U867 (N_867,N_416,N_453);
and U868 (N_868,N_174,N_140);
or U869 (N_869,N_132,N_347);
nand U870 (N_870,N_392,N_383);
nor U871 (N_871,N_540,N_474);
nand U872 (N_872,N_419,N_318);
or U873 (N_873,N_345,N_103);
nand U874 (N_874,N_126,N_401);
or U875 (N_875,N_313,N_97);
xor U876 (N_876,N_306,N_470);
or U877 (N_877,N_35,N_567);
or U878 (N_878,N_295,N_225);
or U879 (N_879,N_523,N_266);
nand U880 (N_880,N_275,N_476);
and U881 (N_881,N_478,N_142);
and U882 (N_882,N_325,N_100);
xnor U883 (N_883,N_239,N_482);
and U884 (N_884,N_412,N_161);
nor U885 (N_885,N_262,N_291);
nand U886 (N_886,N_534,N_88);
xor U887 (N_887,N_343,N_353);
or U888 (N_888,N_249,N_288);
and U889 (N_889,N_449,N_116);
or U890 (N_890,N_265,N_341);
and U891 (N_891,N_432,N_16);
and U892 (N_892,N_544,N_41);
nor U893 (N_893,N_538,N_55);
or U894 (N_894,N_8,N_578);
nand U895 (N_895,N_349,N_191);
and U896 (N_896,N_101,N_198);
and U897 (N_897,N_323,N_390);
xor U898 (N_898,N_468,N_487);
and U899 (N_899,N_426,N_231);
nand U900 (N_900,N_458,N_82);
nor U901 (N_901,N_508,N_22);
or U902 (N_902,N_180,N_454);
xor U903 (N_903,N_243,N_595);
or U904 (N_904,N_210,N_233);
or U905 (N_905,N_517,N_227);
nor U906 (N_906,N_182,N_354);
or U907 (N_907,N_35,N_328);
nor U908 (N_908,N_567,N_248);
nor U909 (N_909,N_72,N_111);
or U910 (N_910,N_511,N_395);
nand U911 (N_911,N_217,N_379);
nor U912 (N_912,N_587,N_497);
nand U913 (N_913,N_69,N_476);
nand U914 (N_914,N_260,N_335);
and U915 (N_915,N_54,N_12);
nor U916 (N_916,N_591,N_58);
nor U917 (N_917,N_50,N_208);
nor U918 (N_918,N_599,N_510);
nor U919 (N_919,N_118,N_26);
nand U920 (N_920,N_592,N_178);
and U921 (N_921,N_48,N_379);
nand U922 (N_922,N_405,N_153);
nor U923 (N_923,N_537,N_392);
and U924 (N_924,N_298,N_188);
or U925 (N_925,N_248,N_310);
xor U926 (N_926,N_7,N_111);
nand U927 (N_927,N_173,N_140);
nand U928 (N_928,N_458,N_497);
and U929 (N_929,N_145,N_23);
and U930 (N_930,N_258,N_471);
or U931 (N_931,N_74,N_496);
xor U932 (N_932,N_367,N_426);
nor U933 (N_933,N_545,N_136);
xor U934 (N_934,N_88,N_506);
or U935 (N_935,N_457,N_558);
nand U936 (N_936,N_533,N_185);
and U937 (N_937,N_550,N_45);
nand U938 (N_938,N_464,N_194);
and U939 (N_939,N_505,N_393);
and U940 (N_940,N_303,N_9);
nor U941 (N_941,N_598,N_354);
nand U942 (N_942,N_379,N_72);
or U943 (N_943,N_495,N_339);
nand U944 (N_944,N_447,N_584);
nand U945 (N_945,N_518,N_48);
and U946 (N_946,N_327,N_321);
nand U947 (N_947,N_531,N_352);
and U948 (N_948,N_376,N_319);
or U949 (N_949,N_362,N_330);
nand U950 (N_950,N_236,N_133);
nand U951 (N_951,N_163,N_563);
or U952 (N_952,N_375,N_159);
or U953 (N_953,N_92,N_163);
nor U954 (N_954,N_99,N_278);
or U955 (N_955,N_537,N_553);
nand U956 (N_956,N_95,N_311);
nor U957 (N_957,N_381,N_147);
nand U958 (N_958,N_590,N_351);
nand U959 (N_959,N_210,N_49);
nor U960 (N_960,N_254,N_18);
nor U961 (N_961,N_477,N_414);
and U962 (N_962,N_191,N_275);
nand U963 (N_963,N_323,N_147);
and U964 (N_964,N_331,N_258);
nand U965 (N_965,N_178,N_507);
and U966 (N_966,N_470,N_210);
xor U967 (N_967,N_427,N_578);
nor U968 (N_968,N_14,N_407);
nand U969 (N_969,N_525,N_548);
and U970 (N_970,N_330,N_531);
nor U971 (N_971,N_137,N_26);
nor U972 (N_972,N_27,N_344);
nor U973 (N_973,N_221,N_150);
and U974 (N_974,N_429,N_49);
nand U975 (N_975,N_135,N_387);
and U976 (N_976,N_402,N_456);
nor U977 (N_977,N_190,N_154);
and U978 (N_978,N_389,N_447);
nor U979 (N_979,N_512,N_373);
or U980 (N_980,N_267,N_218);
nor U981 (N_981,N_337,N_286);
nor U982 (N_982,N_64,N_457);
nor U983 (N_983,N_169,N_331);
nand U984 (N_984,N_180,N_124);
or U985 (N_985,N_126,N_298);
nor U986 (N_986,N_300,N_374);
nor U987 (N_987,N_399,N_151);
xor U988 (N_988,N_545,N_418);
xnor U989 (N_989,N_354,N_175);
nor U990 (N_990,N_206,N_145);
nand U991 (N_991,N_309,N_114);
nor U992 (N_992,N_13,N_378);
and U993 (N_993,N_399,N_79);
nand U994 (N_994,N_515,N_396);
or U995 (N_995,N_250,N_319);
and U996 (N_996,N_590,N_200);
xnor U997 (N_997,N_452,N_59);
or U998 (N_998,N_584,N_533);
xnor U999 (N_999,N_486,N_115);
and U1000 (N_1000,N_507,N_269);
and U1001 (N_1001,N_510,N_418);
or U1002 (N_1002,N_498,N_507);
and U1003 (N_1003,N_322,N_394);
nand U1004 (N_1004,N_566,N_266);
nand U1005 (N_1005,N_227,N_152);
nor U1006 (N_1006,N_311,N_487);
or U1007 (N_1007,N_406,N_531);
xnor U1008 (N_1008,N_493,N_167);
or U1009 (N_1009,N_188,N_471);
or U1010 (N_1010,N_152,N_179);
nor U1011 (N_1011,N_295,N_426);
or U1012 (N_1012,N_599,N_472);
and U1013 (N_1013,N_573,N_461);
and U1014 (N_1014,N_346,N_427);
nand U1015 (N_1015,N_53,N_474);
nor U1016 (N_1016,N_406,N_186);
and U1017 (N_1017,N_306,N_67);
nor U1018 (N_1018,N_184,N_487);
xnor U1019 (N_1019,N_579,N_153);
nand U1020 (N_1020,N_119,N_537);
nand U1021 (N_1021,N_43,N_62);
nand U1022 (N_1022,N_374,N_463);
or U1023 (N_1023,N_598,N_243);
nand U1024 (N_1024,N_89,N_177);
and U1025 (N_1025,N_438,N_526);
nor U1026 (N_1026,N_174,N_393);
xor U1027 (N_1027,N_27,N_546);
and U1028 (N_1028,N_330,N_165);
nand U1029 (N_1029,N_362,N_237);
and U1030 (N_1030,N_355,N_8);
nand U1031 (N_1031,N_475,N_301);
nor U1032 (N_1032,N_35,N_229);
nor U1033 (N_1033,N_10,N_86);
and U1034 (N_1034,N_210,N_247);
and U1035 (N_1035,N_597,N_491);
and U1036 (N_1036,N_211,N_527);
nor U1037 (N_1037,N_300,N_306);
nor U1038 (N_1038,N_455,N_393);
xor U1039 (N_1039,N_79,N_243);
nand U1040 (N_1040,N_36,N_391);
and U1041 (N_1041,N_336,N_422);
and U1042 (N_1042,N_416,N_81);
nor U1043 (N_1043,N_18,N_275);
nor U1044 (N_1044,N_396,N_572);
nor U1045 (N_1045,N_14,N_362);
nor U1046 (N_1046,N_284,N_73);
or U1047 (N_1047,N_397,N_119);
and U1048 (N_1048,N_225,N_88);
and U1049 (N_1049,N_305,N_569);
nor U1050 (N_1050,N_296,N_82);
xor U1051 (N_1051,N_188,N_119);
and U1052 (N_1052,N_161,N_537);
or U1053 (N_1053,N_77,N_597);
nor U1054 (N_1054,N_509,N_513);
nand U1055 (N_1055,N_329,N_398);
nor U1056 (N_1056,N_498,N_41);
nor U1057 (N_1057,N_490,N_372);
or U1058 (N_1058,N_337,N_43);
xnor U1059 (N_1059,N_70,N_539);
xnor U1060 (N_1060,N_260,N_106);
nand U1061 (N_1061,N_417,N_349);
or U1062 (N_1062,N_342,N_184);
xor U1063 (N_1063,N_197,N_30);
nor U1064 (N_1064,N_99,N_181);
and U1065 (N_1065,N_7,N_31);
nand U1066 (N_1066,N_219,N_426);
or U1067 (N_1067,N_45,N_193);
nand U1068 (N_1068,N_406,N_205);
or U1069 (N_1069,N_562,N_196);
xor U1070 (N_1070,N_407,N_534);
and U1071 (N_1071,N_167,N_246);
nand U1072 (N_1072,N_236,N_26);
or U1073 (N_1073,N_60,N_366);
and U1074 (N_1074,N_355,N_553);
nand U1075 (N_1075,N_67,N_275);
nand U1076 (N_1076,N_202,N_138);
nor U1077 (N_1077,N_70,N_112);
nand U1078 (N_1078,N_91,N_49);
nand U1079 (N_1079,N_329,N_549);
xnor U1080 (N_1080,N_410,N_409);
or U1081 (N_1081,N_317,N_358);
xnor U1082 (N_1082,N_1,N_307);
nor U1083 (N_1083,N_44,N_550);
nand U1084 (N_1084,N_490,N_373);
nor U1085 (N_1085,N_141,N_91);
or U1086 (N_1086,N_374,N_558);
nand U1087 (N_1087,N_337,N_118);
and U1088 (N_1088,N_131,N_47);
xnor U1089 (N_1089,N_555,N_571);
nor U1090 (N_1090,N_399,N_447);
nor U1091 (N_1091,N_280,N_376);
nand U1092 (N_1092,N_58,N_203);
and U1093 (N_1093,N_229,N_134);
xnor U1094 (N_1094,N_587,N_402);
and U1095 (N_1095,N_127,N_34);
or U1096 (N_1096,N_284,N_193);
and U1097 (N_1097,N_160,N_124);
nand U1098 (N_1098,N_494,N_437);
xor U1099 (N_1099,N_11,N_366);
and U1100 (N_1100,N_497,N_55);
and U1101 (N_1101,N_524,N_77);
and U1102 (N_1102,N_575,N_475);
nor U1103 (N_1103,N_337,N_373);
or U1104 (N_1104,N_521,N_350);
and U1105 (N_1105,N_43,N_543);
nor U1106 (N_1106,N_298,N_166);
nand U1107 (N_1107,N_346,N_74);
and U1108 (N_1108,N_216,N_294);
nor U1109 (N_1109,N_141,N_388);
nor U1110 (N_1110,N_209,N_141);
and U1111 (N_1111,N_559,N_407);
and U1112 (N_1112,N_582,N_329);
and U1113 (N_1113,N_274,N_103);
or U1114 (N_1114,N_117,N_147);
nand U1115 (N_1115,N_67,N_177);
and U1116 (N_1116,N_216,N_459);
or U1117 (N_1117,N_174,N_135);
or U1118 (N_1118,N_595,N_218);
and U1119 (N_1119,N_271,N_32);
and U1120 (N_1120,N_388,N_523);
or U1121 (N_1121,N_6,N_142);
and U1122 (N_1122,N_495,N_225);
nor U1123 (N_1123,N_558,N_117);
nand U1124 (N_1124,N_110,N_461);
nor U1125 (N_1125,N_203,N_198);
or U1126 (N_1126,N_596,N_174);
or U1127 (N_1127,N_517,N_300);
and U1128 (N_1128,N_102,N_203);
nand U1129 (N_1129,N_279,N_262);
and U1130 (N_1130,N_474,N_597);
nor U1131 (N_1131,N_219,N_0);
nand U1132 (N_1132,N_86,N_445);
and U1133 (N_1133,N_210,N_461);
nand U1134 (N_1134,N_83,N_380);
nand U1135 (N_1135,N_98,N_373);
or U1136 (N_1136,N_78,N_489);
or U1137 (N_1137,N_472,N_161);
nand U1138 (N_1138,N_173,N_232);
nor U1139 (N_1139,N_515,N_579);
and U1140 (N_1140,N_92,N_181);
nor U1141 (N_1141,N_119,N_381);
or U1142 (N_1142,N_105,N_542);
nor U1143 (N_1143,N_524,N_502);
nand U1144 (N_1144,N_495,N_358);
or U1145 (N_1145,N_48,N_214);
and U1146 (N_1146,N_460,N_418);
and U1147 (N_1147,N_14,N_501);
xnor U1148 (N_1148,N_487,N_431);
or U1149 (N_1149,N_31,N_82);
nand U1150 (N_1150,N_550,N_449);
nand U1151 (N_1151,N_300,N_373);
and U1152 (N_1152,N_397,N_114);
nor U1153 (N_1153,N_526,N_477);
or U1154 (N_1154,N_479,N_223);
nand U1155 (N_1155,N_575,N_524);
nor U1156 (N_1156,N_469,N_47);
and U1157 (N_1157,N_363,N_409);
and U1158 (N_1158,N_424,N_134);
nand U1159 (N_1159,N_488,N_194);
xor U1160 (N_1160,N_585,N_151);
xor U1161 (N_1161,N_304,N_264);
and U1162 (N_1162,N_359,N_582);
or U1163 (N_1163,N_278,N_271);
nor U1164 (N_1164,N_328,N_514);
nand U1165 (N_1165,N_537,N_415);
and U1166 (N_1166,N_453,N_283);
and U1167 (N_1167,N_487,N_131);
and U1168 (N_1168,N_492,N_529);
nand U1169 (N_1169,N_591,N_104);
or U1170 (N_1170,N_212,N_336);
nor U1171 (N_1171,N_12,N_160);
nor U1172 (N_1172,N_492,N_598);
and U1173 (N_1173,N_38,N_270);
or U1174 (N_1174,N_486,N_320);
and U1175 (N_1175,N_369,N_9);
or U1176 (N_1176,N_551,N_554);
and U1177 (N_1177,N_129,N_407);
and U1178 (N_1178,N_297,N_216);
xnor U1179 (N_1179,N_462,N_542);
nand U1180 (N_1180,N_142,N_397);
or U1181 (N_1181,N_357,N_474);
nor U1182 (N_1182,N_541,N_550);
or U1183 (N_1183,N_499,N_123);
and U1184 (N_1184,N_592,N_65);
or U1185 (N_1185,N_284,N_488);
and U1186 (N_1186,N_125,N_224);
nand U1187 (N_1187,N_45,N_404);
or U1188 (N_1188,N_161,N_113);
and U1189 (N_1189,N_435,N_132);
or U1190 (N_1190,N_413,N_184);
nand U1191 (N_1191,N_382,N_69);
or U1192 (N_1192,N_38,N_510);
or U1193 (N_1193,N_530,N_528);
nand U1194 (N_1194,N_465,N_299);
nand U1195 (N_1195,N_239,N_329);
or U1196 (N_1196,N_192,N_567);
nand U1197 (N_1197,N_20,N_110);
and U1198 (N_1198,N_349,N_502);
or U1199 (N_1199,N_274,N_236);
xor U1200 (N_1200,N_767,N_892);
nor U1201 (N_1201,N_654,N_909);
or U1202 (N_1202,N_1129,N_956);
nor U1203 (N_1203,N_801,N_685);
nand U1204 (N_1204,N_998,N_769);
or U1205 (N_1205,N_962,N_1125);
nor U1206 (N_1206,N_938,N_1174);
xnor U1207 (N_1207,N_694,N_754);
nor U1208 (N_1208,N_770,N_882);
nand U1209 (N_1209,N_885,N_838);
nor U1210 (N_1210,N_758,N_789);
or U1211 (N_1211,N_863,N_840);
and U1212 (N_1212,N_939,N_883);
nand U1213 (N_1213,N_1100,N_675);
or U1214 (N_1214,N_1005,N_923);
nand U1215 (N_1215,N_960,N_805);
or U1216 (N_1216,N_827,N_1095);
xnor U1217 (N_1217,N_1172,N_1008);
nor U1218 (N_1218,N_1024,N_1045);
or U1219 (N_1219,N_639,N_611);
or U1220 (N_1220,N_844,N_860);
nor U1221 (N_1221,N_1036,N_1059);
and U1222 (N_1222,N_983,N_705);
and U1223 (N_1223,N_1170,N_944);
nand U1224 (N_1224,N_742,N_776);
or U1225 (N_1225,N_1073,N_899);
and U1226 (N_1226,N_1040,N_1115);
and U1227 (N_1227,N_826,N_622);
nor U1228 (N_1228,N_992,N_1180);
and U1229 (N_1229,N_782,N_804);
nor U1230 (N_1230,N_773,N_709);
xor U1231 (N_1231,N_1034,N_800);
and U1232 (N_1232,N_1199,N_1162);
nand U1233 (N_1233,N_718,N_684);
nor U1234 (N_1234,N_972,N_647);
nand U1235 (N_1235,N_695,N_691);
nor U1236 (N_1236,N_672,N_1065);
and U1237 (N_1237,N_964,N_867);
nor U1238 (N_1238,N_957,N_866);
nor U1239 (N_1239,N_797,N_1193);
or U1240 (N_1240,N_880,N_1013);
nand U1241 (N_1241,N_884,N_1101);
or U1242 (N_1242,N_761,N_1185);
nand U1243 (N_1243,N_603,N_1058);
nor U1244 (N_1244,N_819,N_1016);
nand U1245 (N_1245,N_881,N_706);
xnor U1246 (N_1246,N_728,N_894);
nor U1247 (N_1247,N_913,N_1145);
or U1248 (N_1248,N_976,N_693);
and U1249 (N_1249,N_610,N_1166);
or U1250 (N_1250,N_711,N_793);
or U1251 (N_1251,N_653,N_1075);
and U1252 (N_1252,N_991,N_859);
nor U1253 (N_1253,N_1157,N_868);
nor U1254 (N_1254,N_795,N_919);
xnor U1255 (N_1255,N_1035,N_808);
and U1256 (N_1256,N_936,N_640);
nor U1257 (N_1257,N_621,N_903);
nand U1258 (N_1258,N_974,N_636);
nand U1259 (N_1259,N_616,N_1144);
nand U1260 (N_1260,N_824,N_1022);
and U1261 (N_1261,N_869,N_1176);
and U1262 (N_1262,N_655,N_739);
and U1263 (N_1263,N_674,N_833);
nand U1264 (N_1264,N_916,N_608);
or U1265 (N_1265,N_961,N_949);
xnor U1266 (N_1266,N_900,N_1152);
and U1267 (N_1267,N_1117,N_1028);
and U1268 (N_1268,N_822,N_1140);
xor U1269 (N_1269,N_1088,N_637);
nor U1270 (N_1270,N_785,N_673);
nor U1271 (N_1271,N_721,N_634);
and U1272 (N_1272,N_757,N_988);
and U1273 (N_1273,N_814,N_723);
nor U1274 (N_1274,N_989,N_698);
nand U1275 (N_1275,N_952,N_905);
and U1276 (N_1276,N_835,N_1160);
nand U1277 (N_1277,N_1077,N_1044);
and U1278 (N_1278,N_763,N_1167);
or U1279 (N_1279,N_712,N_690);
nand U1280 (N_1280,N_1063,N_624);
nor U1281 (N_1281,N_813,N_646);
nor U1282 (N_1282,N_652,N_1012);
or U1283 (N_1283,N_715,N_683);
or U1284 (N_1284,N_696,N_745);
or U1285 (N_1285,N_642,N_915);
or U1286 (N_1286,N_807,N_1116);
or U1287 (N_1287,N_1134,N_921);
nor U1288 (N_1288,N_933,N_612);
and U1289 (N_1289,N_837,N_1017);
and U1290 (N_1290,N_1067,N_765);
nor U1291 (N_1291,N_659,N_836);
nand U1292 (N_1292,N_928,N_1025);
nor U1293 (N_1293,N_777,N_663);
xnor U1294 (N_1294,N_978,N_979);
nor U1295 (N_1295,N_1108,N_1099);
nand U1296 (N_1296,N_609,N_902);
and U1297 (N_1297,N_973,N_1014);
and U1298 (N_1298,N_953,N_678);
or U1299 (N_1299,N_970,N_1143);
nor U1300 (N_1300,N_668,N_701);
or U1301 (N_1301,N_604,N_771);
nor U1302 (N_1302,N_656,N_846);
nor U1303 (N_1303,N_716,N_811);
or U1304 (N_1304,N_1197,N_628);
nor U1305 (N_1305,N_1098,N_1078);
and U1306 (N_1306,N_602,N_1027);
and U1307 (N_1307,N_726,N_1018);
and U1308 (N_1308,N_1091,N_1064);
nor U1309 (N_1309,N_889,N_1079);
nor U1310 (N_1310,N_1061,N_852);
and U1311 (N_1311,N_760,N_1010);
and U1312 (N_1312,N_855,N_630);
and U1313 (N_1313,N_743,N_725);
xor U1314 (N_1314,N_911,N_1136);
xnor U1315 (N_1315,N_1090,N_823);
or U1316 (N_1316,N_1119,N_888);
xnor U1317 (N_1317,N_1038,N_831);
nand U1318 (N_1318,N_1131,N_839);
nand U1319 (N_1319,N_687,N_618);
and U1320 (N_1320,N_1050,N_1031);
or U1321 (N_1321,N_748,N_1113);
and U1322 (N_1322,N_1175,N_908);
and U1323 (N_1323,N_922,N_920);
nor U1324 (N_1324,N_768,N_871);
nor U1325 (N_1325,N_699,N_834);
or U1326 (N_1326,N_688,N_649);
nor U1327 (N_1327,N_779,N_1039);
and U1328 (N_1328,N_1198,N_662);
or U1329 (N_1329,N_849,N_932);
xnor U1330 (N_1330,N_906,N_1187);
nand U1331 (N_1331,N_1107,N_682);
and U1332 (N_1332,N_692,N_958);
nand U1333 (N_1333,N_810,N_1135);
and U1334 (N_1334,N_1169,N_1093);
nand U1335 (N_1335,N_1195,N_1142);
nor U1336 (N_1336,N_1094,N_708);
or U1337 (N_1337,N_858,N_1060);
xor U1338 (N_1338,N_806,N_669);
xor U1339 (N_1339,N_778,N_710);
and U1340 (N_1340,N_802,N_650);
nand U1341 (N_1341,N_735,N_862);
nand U1342 (N_1342,N_661,N_635);
nand U1343 (N_1343,N_619,N_766);
nand U1344 (N_1344,N_878,N_1071);
xor U1345 (N_1345,N_910,N_1092);
nor U1346 (N_1346,N_1054,N_781);
or U1347 (N_1347,N_677,N_1041);
and U1348 (N_1348,N_996,N_667);
nand U1349 (N_1349,N_1103,N_1109);
nor U1350 (N_1350,N_798,N_738);
nor U1351 (N_1351,N_843,N_1114);
and U1352 (N_1352,N_1068,N_1019);
nor U1353 (N_1353,N_714,N_1141);
and U1354 (N_1354,N_947,N_1165);
and U1355 (N_1355,N_914,N_1177);
or U1356 (N_1356,N_982,N_887);
nor U1357 (N_1357,N_1189,N_967);
nand U1358 (N_1358,N_857,N_657);
nor U1359 (N_1359,N_741,N_1000);
nand U1360 (N_1360,N_1139,N_803);
nor U1361 (N_1361,N_1179,N_830);
and U1362 (N_1362,N_901,N_1006);
or U1363 (N_1363,N_631,N_1074);
nand U1364 (N_1364,N_997,N_818);
xnor U1365 (N_1365,N_935,N_854);
nor U1366 (N_1366,N_1057,N_736);
or U1367 (N_1367,N_1009,N_815);
or U1368 (N_1368,N_1056,N_876);
nand U1369 (N_1369,N_744,N_1154);
nand U1370 (N_1370,N_1047,N_681);
nand U1371 (N_1371,N_733,N_969);
nand U1372 (N_1372,N_981,N_1032);
and U1373 (N_1373,N_842,N_788);
nand U1374 (N_1374,N_1087,N_792);
xnor U1375 (N_1375,N_633,N_791);
xnor U1376 (N_1376,N_1146,N_1178);
nand U1377 (N_1377,N_945,N_937);
or U1378 (N_1378,N_942,N_845);
nand U1379 (N_1379,N_1021,N_1104);
nor U1380 (N_1380,N_749,N_1046);
and U1381 (N_1381,N_753,N_676);
nor U1382 (N_1382,N_1132,N_848);
and U1383 (N_1383,N_1023,N_1124);
nor U1384 (N_1384,N_898,N_1163);
and U1385 (N_1385,N_877,N_809);
nor U1386 (N_1386,N_1133,N_1155);
nand U1387 (N_1387,N_719,N_1150);
xor U1388 (N_1388,N_1123,N_1004);
nor U1389 (N_1389,N_893,N_703);
xnor U1390 (N_1390,N_751,N_934);
or U1391 (N_1391,N_1171,N_727);
and U1392 (N_1392,N_737,N_1138);
and U1393 (N_1393,N_940,N_1126);
and U1394 (N_1394,N_1184,N_1128);
nand U1395 (N_1395,N_713,N_775);
xor U1396 (N_1396,N_790,N_856);
and U1397 (N_1397,N_643,N_1066);
and U1398 (N_1398,N_984,N_658);
xnor U1399 (N_1399,N_828,N_1149);
and U1400 (N_1400,N_600,N_783);
or U1401 (N_1401,N_886,N_601);
nor U1402 (N_1402,N_774,N_1055);
or U1403 (N_1403,N_787,N_1089);
nor U1404 (N_1404,N_873,N_1049);
or U1405 (N_1405,N_1151,N_671);
and U1406 (N_1406,N_891,N_651);
nand U1407 (N_1407,N_620,N_707);
nand U1408 (N_1408,N_975,N_874);
or U1409 (N_1409,N_924,N_895);
nand U1410 (N_1410,N_613,N_1084);
nor U1411 (N_1411,N_1030,N_762);
nand U1412 (N_1412,N_1080,N_954);
and U1413 (N_1413,N_1148,N_966);
and U1414 (N_1414,N_875,N_1020);
xnor U1415 (N_1415,N_1076,N_980);
nor U1416 (N_1416,N_1147,N_829);
nor U1417 (N_1417,N_985,N_772);
nand U1418 (N_1418,N_1190,N_1026);
nand U1419 (N_1419,N_606,N_1121);
nand U1420 (N_1420,N_977,N_641);
nor U1421 (N_1421,N_955,N_971);
xnor U1422 (N_1422,N_853,N_700);
and U1423 (N_1423,N_1105,N_1081);
nor U1424 (N_1424,N_927,N_1181);
nand U1425 (N_1425,N_821,N_965);
nand U1426 (N_1426,N_680,N_697);
xor U1427 (N_1427,N_948,N_740);
xnor U1428 (N_1428,N_665,N_1096);
nand U1429 (N_1429,N_617,N_1097);
nor U1430 (N_1430,N_926,N_605);
nand U1431 (N_1431,N_930,N_1042);
nor U1432 (N_1432,N_756,N_1069);
nor U1433 (N_1433,N_847,N_1161);
nand U1434 (N_1434,N_1086,N_968);
nand U1435 (N_1435,N_1168,N_764);
nand U1436 (N_1436,N_1072,N_816);
or U1437 (N_1437,N_1082,N_925);
nand U1438 (N_1438,N_931,N_794);
nor U1439 (N_1439,N_625,N_1048);
nor U1440 (N_1440,N_1158,N_1111);
nor U1441 (N_1441,N_912,N_645);
nor U1442 (N_1442,N_1029,N_799);
nand U1443 (N_1443,N_993,N_747);
and U1444 (N_1444,N_626,N_1011);
or U1445 (N_1445,N_720,N_729);
or U1446 (N_1446,N_784,N_1137);
nand U1447 (N_1447,N_1164,N_1130);
and U1448 (N_1448,N_1085,N_679);
nand U1449 (N_1449,N_724,N_896);
nor U1450 (N_1450,N_1153,N_623);
nor U1451 (N_1451,N_832,N_897);
or U1452 (N_1452,N_730,N_786);
or U1453 (N_1453,N_629,N_1102);
nand U1454 (N_1454,N_959,N_1159);
or U1455 (N_1455,N_796,N_750);
nand U1456 (N_1456,N_638,N_1002);
nor U1457 (N_1457,N_689,N_872);
xnor U1458 (N_1458,N_950,N_1183);
or U1459 (N_1459,N_1007,N_1037);
nor U1460 (N_1460,N_780,N_999);
nor U1461 (N_1461,N_755,N_1191);
or U1462 (N_1462,N_1053,N_752);
or U1463 (N_1463,N_904,N_722);
or U1464 (N_1464,N_1051,N_951);
nor U1465 (N_1465,N_734,N_1122);
nand U1466 (N_1466,N_1188,N_917);
or U1467 (N_1467,N_1194,N_1186);
nand U1468 (N_1468,N_1192,N_614);
and U1469 (N_1469,N_946,N_907);
xor U1470 (N_1470,N_1120,N_615);
or U1471 (N_1471,N_850,N_632);
and U1472 (N_1472,N_717,N_1173);
nand U1473 (N_1473,N_1001,N_1118);
and U1474 (N_1474,N_1127,N_759);
nand U1475 (N_1475,N_861,N_1062);
and U1476 (N_1476,N_825,N_704);
and U1477 (N_1477,N_732,N_817);
or U1478 (N_1478,N_890,N_1043);
nand U1479 (N_1479,N_812,N_1015);
or U1480 (N_1480,N_929,N_851);
and U1481 (N_1481,N_879,N_963);
nand U1482 (N_1482,N_731,N_746);
or U1483 (N_1483,N_607,N_627);
nand U1484 (N_1484,N_820,N_870);
and U1485 (N_1485,N_986,N_864);
nand U1486 (N_1486,N_686,N_1052);
or U1487 (N_1487,N_660,N_1033);
or U1488 (N_1488,N_1003,N_648);
and U1489 (N_1489,N_1110,N_1182);
or U1490 (N_1490,N_1083,N_990);
or U1491 (N_1491,N_995,N_994);
xnor U1492 (N_1492,N_987,N_1112);
and U1493 (N_1493,N_865,N_1156);
nor U1494 (N_1494,N_941,N_943);
xor U1495 (N_1495,N_702,N_841);
nand U1496 (N_1496,N_1196,N_664);
and U1497 (N_1497,N_670,N_918);
nand U1498 (N_1498,N_644,N_1070);
nor U1499 (N_1499,N_666,N_1106);
or U1500 (N_1500,N_851,N_817);
or U1501 (N_1501,N_756,N_917);
and U1502 (N_1502,N_875,N_1179);
nand U1503 (N_1503,N_1127,N_1089);
or U1504 (N_1504,N_744,N_1088);
xnor U1505 (N_1505,N_616,N_1159);
or U1506 (N_1506,N_899,N_825);
or U1507 (N_1507,N_1140,N_647);
or U1508 (N_1508,N_652,N_1128);
and U1509 (N_1509,N_654,N_655);
and U1510 (N_1510,N_1063,N_922);
nand U1511 (N_1511,N_991,N_1146);
nor U1512 (N_1512,N_918,N_935);
nand U1513 (N_1513,N_614,N_993);
xnor U1514 (N_1514,N_1090,N_602);
or U1515 (N_1515,N_797,N_671);
nor U1516 (N_1516,N_1144,N_790);
xor U1517 (N_1517,N_1111,N_764);
or U1518 (N_1518,N_1177,N_921);
or U1519 (N_1519,N_1135,N_651);
and U1520 (N_1520,N_1125,N_1016);
nor U1521 (N_1521,N_737,N_854);
nand U1522 (N_1522,N_968,N_1035);
or U1523 (N_1523,N_809,N_1014);
and U1524 (N_1524,N_1134,N_1058);
nor U1525 (N_1525,N_915,N_734);
and U1526 (N_1526,N_904,N_781);
nand U1527 (N_1527,N_684,N_637);
nor U1528 (N_1528,N_691,N_1006);
nor U1529 (N_1529,N_976,N_893);
nor U1530 (N_1530,N_1014,N_684);
nor U1531 (N_1531,N_918,N_743);
nand U1532 (N_1532,N_1037,N_786);
nor U1533 (N_1533,N_925,N_760);
nor U1534 (N_1534,N_779,N_759);
or U1535 (N_1535,N_804,N_723);
nand U1536 (N_1536,N_870,N_612);
nor U1537 (N_1537,N_968,N_811);
and U1538 (N_1538,N_996,N_1067);
and U1539 (N_1539,N_709,N_1119);
and U1540 (N_1540,N_718,N_1080);
or U1541 (N_1541,N_1196,N_808);
nand U1542 (N_1542,N_746,N_848);
nor U1543 (N_1543,N_976,N_862);
nand U1544 (N_1544,N_774,N_743);
nand U1545 (N_1545,N_670,N_628);
nor U1546 (N_1546,N_1136,N_603);
nand U1547 (N_1547,N_738,N_814);
nand U1548 (N_1548,N_1088,N_1017);
xnor U1549 (N_1549,N_990,N_639);
or U1550 (N_1550,N_766,N_1105);
and U1551 (N_1551,N_1190,N_1188);
nor U1552 (N_1552,N_685,N_1112);
nand U1553 (N_1553,N_830,N_601);
xnor U1554 (N_1554,N_818,N_747);
nand U1555 (N_1555,N_925,N_850);
nor U1556 (N_1556,N_1024,N_811);
and U1557 (N_1557,N_988,N_966);
or U1558 (N_1558,N_906,N_611);
nand U1559 (N_1559,N_923,N_648);
nand U1560 (N_1560,N_683,N_671);
xnor U1561 (N_1561,N_919,N_819);
and U1562 (N_1562,N_949,N_917);
nand U1563 (N_1563,N_748,N_877);
and U1564 (N_1564,N_945,N_1093);
and U1565 (N_1565,N_1126,N_1098);
nand U1566 (N_1566,N_1063,N_1131);
or U1567 (N_1567,N_708,N_938);
and U1568 (N_1568,N_751,N_622);
xnor U1569 (N_1569,N_647,N_807);
nor U1570 (N_1570,N_944,N_990);
and U1571 (N_1571,N_994,N_682);
nand U1572 (N_1572,N_719,N_782);
and U1573 (N_1573,N_987,N_920);
nor U1574 (N_1574,N_836,N_744);
xnor U1575 (N_1575,N_702,N_1070);
nand U1576 (N_1576,N_997,N_829);
xnor U1577 (N_1577,N_980,N_1007);
xnor U1578 (N_1578,N_770,N_825);
nand U1579 (N_1579,N_1079,N_1108);
nor U1580 (N_1580,N_916,N_614);
or U1581 (N_1581,N_926,N_921);
nand U1582 (N_1582,N_639,N_894);
nand U1583 (N_1583,N_962,N_908);
nor U1584 (N_1584,N_795,N_792);
or U1585 (N_1585,N_972,N_1083);
or U1586 (N_1586,N_1137,N_683);
and U1587 (N_1587,N_678,N_610);
nor U1588 (N_1588,N_1145,N_740);
xnor U1589 (N_1589,N_797,N_833);
xor U1590 (N_1590,N_1104,N_912);
or U1591 (N_1591,N_726,N_952);
nand U1592 (N_1592,N_1149,N_1041);
nand U1593 (N_1593,N_686,N_985);
nor U1594 (N_1594,N_905,N_651);
or U1595 (N_1595,N_1120,N_908);
or U1596 (N_1596,N_733,N_719);
nand U1597 (N_1597,N_910,N_707);
and U1598 (N_1598,N_851,N_678);
nor U1599 (N_1599,N_1154,N_1032);
nand U1600 (N_1600,N_831,N_1170);
or U1601 (N_1601,N_810,N_780);
or U1602 (N_1602,N_1109,N_657);
and U1603 (N_1603,N_1192,N_1093);
and U1604 (N_1604,N_750,N_659);
nor U1605 (N_1605,N_645,N_715);
or U1606 (N_1606,N_978,N_1148);
xnor U1607 (N_1607,N_925,N_699);
nand U1608 (N_1608,N_718,N_818);
and U1609 (N_1609,N_907,N_722);
nand U1610 (N_1610,N_896,N_692);
or U1611 (N_1611,N_659,N_1178);
or U1612 (N_1612,N_865,N_717);
nor U1613 (N_1613,N_699,N_817);
xor U1614 (N_1614,N_773,N_996);
or U1615 (N_1615,N_705,N_665);
nor U1616 (N_1616,N_1019,N_868);
and U1617 (N_1617,N_1124,N_638);
or U1618 (N_1618,N_988,N_1165);
and U1619 (N_1619,N_1106,N_965);
or U1620 (N_1620,N_923,N_1190);
xnor U1621 (N_1621,N_693,N_890);
nand U1622 (N_1622,N_1015,N_1071);
and U1623 (N_1623,N_917,N_937);
nor U1624 (N_1624,N_862,N_1007);
or U1625 (N_1625,N_796,N_1057);
or U1626 (N_1626,N_720,N_696);
nand U1627 (N_1627,N_807,N_894);
nand U1628 (N_1628,N_600,N_1066);
and U1629 (N_1629,N_739,N_1084);
nand U1630 (N_1630,N_973,N_655);
nand U1631 (N_1631,N_1126,N_982);
or U1632 (N_1632,N_1062,N_1173);
nor U1633 (N_1633,N_1073,N_1093);
and U1634 (N_1634,N_640,N_995);
and U1635 (N_1635,N_713,N_631);
nand U1636 (N_1636,N_996,N_632);
nor U1637 (N_1637,N_1080,N_1179);
nor U1638 (N_1638,N_1098,N_691);
or U1639 (N_1639,N_1026,N_820);
nand U1640 (N_1640,N_832,N_1193);
nor U1641 (N_1641,N_975,N_1094);
nor U1642 (N_1642,N_752,N_838);
and U1643 (N_1643,N_999,N_803);
nor U1644 (N_1644,N_847,N_883);
nor U1645 (N_1645,N_898,N_674);
nand U1646 (N_1646,N_1130,N_674);
nand U1647 (N_1647,N_1009,N_1119);
and U1648 (N_1648,N_852,N_605);
nand U1649 (N_1649,N_692,N_652);
nand U1650 (N_1650,N_1150,N_924);
xor U1651 (N_1651,N_1174,N_993);
nor U1652 (N_1652,N_1143,N_758);
or U1653 (N_1653,N_740,N_733);
nand U1654 (N_1654,N_1066,N_1129);
nand U1655 (N_1655,N_886,N_629);
and U1656 (N_1656,N_838,N_1062);
or U1657 (N_1657,N_1122,N_723);
or U1658 (N_1658,N_1106,N_645);
or U1659 (N_1659,N_732,N_603);
and U1660 (N_1660,N_1046,N_1102);
and U1661 (N_1661,N_1143,N_921);
nor U1662 (N_1662,N_802,N_854);
nand U1663 (N_1663,N_816,N_938);
or U1664 (N_1664,N_603,N_766);
nand U1665 (N_1665,N_706,N_604);
nor U1666 (N_1666,N_678,N_746);
nand U1667 (N_1667,N_914,N_984);
nand U1668 (N_1668,N_1087,N_998);
xor U1669 (N_1669,N_873,N_641);
and U1670 (N_1670,N_916,N_663);
nor U1671 (N_1671,N_1125,N_849);
nor U1672 (N_1672,N_1165,N_1155);
nand U1673 (N_1673,N_1113,N_990);
and U1674 (N_1674,N_943,N_722);
nor U1675 (N_1675,N_804,N_1071);
xor U1676 (N_1676,N_1193,N_1117);
xnor U1677 (N_1677,N_1100,N_643);
and U1678 (N_1678,N_950,N_787);
and U1679 (N_1679,N_844,N_859);
nand U1680 (N_1680,N_668,N_1040);
and U1681 (N_1681,N_1060,N_966);
and U1682 (N_1682,N_853,N_822);
or U1683 (N_1683,N_1148,N_921);
and U1684 (N_1684,N_864,N_905);
nor U1685 (N_1685,N_1087,N_907);
nor U1686 (N_1686,N_838,N_653);
nand U1687 (N_1687,N_884,N_652);
or U1688 (N_1688,N_879,N_730);
nand U1689 (N_1689,N_1195,N_1100);
nor U1690 (N_1690,N_1026,N_727);
nor U1691 (N_1691,N_641,N_1035);
xnor U1692 (N_1692,N_710,N_1031);
or U1693 (N_1693,N_931,N_808);
or U1694 (N_1694,N_766,N_679);
and U1695 (N_1695,N_623,N_1109);
xor U1696 (N_1696,N_898,N_1154);
or U1697 (N_1697,N_1115,N_1014);
nand U1698 (N_1698,N_603,N_1091);
and U1699 (N_1699,N_866,N_916);
or U1700 (N_1700,N_697,N_1002);
nor U1701 (N_1701,N_715,N_1016);
or U1702 (N_1702,N_938,N_704);
nor U1703 (N_1703,N_618,N_875);
nor U1704 (N_1704,N_836,N_1157);
nand U1705 (N_1705,N_754,N_634);
and U1706 (N_1706,N_1107,N_1139);
or U1707 (N_1707,N_940,N_744);
xor U1708 (N_1708,N_1033,N_628);
and U1709 (N_1709,N_762,N_811);
and U1710 (N_1710,N_1012,N_712);
nand U1711 (N_1711,N_612,N_966);
nor U1712 (N_1712,N_807,N_629);
or U1713 (N_1713,N_969,N_1090);
and U1714 (N_1714,N_879,N_757);
nor U1715 (N_1715,N_635,N_869);
nor U1716 (N_1716,N_836,N_1188);
xnor U1717 (N_1717,N_1173,N_1065);
nand U1718 (N_1718,N_790,N_1008);
or U1719 (N_1719,N_843,N_759);
nand U1720 (N_1720,N_697,N_698);
and U1721 (N_1721,N_1098,N_876);
nor U1722 (N_1722,N_637,N_843);
and U1723 (N_1723,N_749,N_823);
or U1724 (N_1724,N_647,N_726);
nor U1725 (N_1725,N_1135,N_955);
and U1726 (N_1726,N_820,N_788);
or U1727 (N_1727,N_863,N_957);
nor U1728 (N_1728,N_1057,N_1040);
and U1729 (N_1729,N_1091,N_1198);
and U1730 (N_1730,N_883,N_792);
nand U1731 (N_1731,N_806,N_832);
or U1732 (N_1732,N_1029,N_915);
nor U1733 (N_1733,N_800,N_1113);
nor U1734 (N_1734,N_1057,N_778);
or U1735 (N_1735,N_1053,N_985);
or U1736 (N_1736,N_984,N_1096);
nand U1737 (N_1737,N_654,N_1110);
nand U1738 (N_1738,N_857,N_702);
nor U1739 (N_1739,N_750,N_742);
nor U1740 (N_1740,N_819,N_823);
and U1741 (N_1741,N_721,N_1097);
nor U1742 (N_1742,N_1190,N_1077);
and U1743 (N_1743,N_888,N_1006);
or U1744 (N_1744,N_875,N_670);
nand U1745 (N_1745,N_829,N_820);
nor U1746 (N_1746,N_1182,N_687);
or U1747 (N_1747,N_716,N_1178);
nor U1748 (N_1748,N_822,N_1065);
xor U1749 (N_1749,N_603,N_634);
or U1750 (N_1750,N_1180,N_889);
or U1751 (N_1751,N_1005,N_1050);
nor U1752 (N_1752,N_700,N_879);
nand U1753 (N_1753,N_1130,N_655);
xor U1754 (N_1754,N_1197,N_971);
xnor U1755 (N_1755,N_766,N_988);
and U1756 (N_1756,N_750,N_727);
or U1757 (N_1757,N_647,N_1100);
nand U1758 (N_1758,N_1180,N_724);
and U1759 (N_1759,N_1194,N_799);
or U1760 (N_1760,N_1126,N_991);
or U1761 (N_1761,N_677,N_842);
xor U1762 (N_1762,N_796,N_1121);
nor U1763 (N_1763,N_745,N_678);
nor U1764 (N_1764,N_877,N_1089);
and U1765 (N_1765,N_908,N_1073);
and U1766 (N_1766,N_713,N_935);
nor U1767 (N_1767,N_707,N_959);
nand U1768 (N_1768,N_680,N_1160);
nand U1769 (N_1769,N_1115,N_1197);
and U1770 (N_1770,N_726,N_1132);
or U1771 (N_1771,N_754,N_840);
nor U1772 (N_1772,N_695,N_716);
nand U1773 (N_1773,N_884,N_1089);
xor U1774 (N_1774,N_742,N_969);
nand U1775 (N_1775,N_885,N_824);
xnor U1776 (N_1776,N_1064,N_1018);
or U1777 (N_1777,N_1144,N_849);
and U1778 (N_1778,N_682,N_761);
and U1779 (N_1779,N_739,N_1174);
nor U1780 (N_1780,N_911,N_1053);
or U1781 (N_1781,N_1069,N_1103);
nand U1782 (N_1782,N_691,N_808);
or U1783 (N_1783,N_861,N_624);
or U1784 (N_1784,N_861,N_908);
and U1785 (N_1785,N_1055,N_685);
and U1786 (N_1786,N_851,N_1006);
nand U1787 (N_1787,N_825,N_815);
or U1788 (N_1788,N_957,N_639);
nor U1789 (N_1789,N_987,N_871);
or U1790 (N_1790,N_700,N_970);
nor U1791 (N_1791,N_741,N_1145);
xnor U1792 (N_1792,N_1054,N_1091);
and U1793 (N_1793,N_672,N_940);
or U1794 (N_1794,N_838,N_680);
nand U1795 (N_1795,N_729,N_1001);
and U1796 (N_1796,N_910,N_1039);
and U1797 (N_1797,N_807,N_1036);
and U1798 (N_1798,N_611,N_1152);
nor U1799 (N_1799,N_936,N_1191);
and U1800 (N_1800,N_1262,N_1782);
and U1801 (N_1801,N_1779,N_1472);
nand U1802 (N_1802,N_1711,N_1726);
nor U1803 (N_1803,N_1468,N_1645);
nand U1804 (N_1804,N_1258,N_1723);
nand U1805 (N_1805,N_1799,N_1390);
nor U1806 (N_1806,N_1225,N_1315);
nor U1807 (N_1807,N_1751,N_1479);
nand U1808 (N_1808,N_1531,N_1559);
nand U1809 (N_1809,N_1244,N_1329);
nor U1810 (N_1810,N_1270,N_1471);
or U1811 (N_1811,N_1647,N_1630);
or U1812 (N_1812,N_1337,N_1210);
or U1813 (N_1813,N_1437,N_1394);
nand U1814 (N_1814,N_1445,N_1469);
and U1815 (N_1815,N_1667,N_1374);
nor U1816 (N_1816,N_1780,N_1538);
nor U1817 (N_1817,N_1633,N_1773);
or U1818 (N_1818,N_1673,N_1528);
and U1819 (N_1819,N_1434,N_1482);
and U1820 (N_1820,N_1429,N_1540);
xor U1821 (N_1821,N_1610,N_1611);
and U1822 (N_1822,N_1478,N_1426);
and U1823 (N_1823,N_1766,N_1509);
or U1824 (N_1824,N_1435,N_1353);
nor U1825 (N_1825,N_1452,N_1288);
nand U1826 (N_1826,N_1397,N_1692);
and U1827 (N_1827,N_1699,N_1688);
and U1828 (N_1828,N_1614,N_1443);
nand U1829 (N_1829,N_1517,N_1295);
nand U1830 (N_1830,N_1696,N_1748);
nand U1831 (N_1831,N_1676,N_1709);
and U1832 (N_1832,N_1551,N_1693);
and U1833 (N_1833,N_1739,N_1318);
and U1834 (N_1834,N_1404,N_1694);
nand U1835 (N_1835,N_1746,N_1798);
nor U1836 (N_1836,N_1489,N_1500);
xnor U1837 (N_1837,N_1408,N_1521);
nand U1838 (N_1838,N_1393,N_1345);
or U1839 (N_1839,N_1402,N_1617);
and U1840 (N_1840,N_1260,N_1439);
nand U1841 (N_1841,N_1259,N_1794);
xnor U1842 (N_1842,N_1275,N_1379);
and U1843 (N_1843,N_1389,N_1367);
and U1844 (N_1844,N_1214,N_1593);
nand U1845 (N_1845,N_1369,N_1573);
and U1846 (N_1846,N_1554,N_1365);
or U1847 (N_1847,N_1226,N_1207);
or U1848 (N_1848,N_1724,N_1741);
and U1849 (N_1849,N_1607,N_1366);
and U1850 (N_1850,N_1771,N_1219);
and U1851 (N_1851,N_1409,N_1406);
and U1852 (N_1852,N_1496,N_1330);
or U1853 (N_1853,N_1555,N_1216);
xnor U1854 (N_1854,N_1255,N_1490);
nand U1855 (N_1855,N_1307,N_1264);
nand U1856 (N_1856,N_1627,N_1632);
nor U1857 (N_1857,N_1356,N_1631);
nand U1858 (N_1858,N_1209,N_1350);
nand U1859 (N_1859,N_1520,N_1564);
nor U1860 (N_1860,N_1513,N_1675);
xnor U1861 (N_1861,N_1338,N_1599);
nand U1862 (N_1862,N_1570,N_1618);
or U1863 (N_1863,N_1299,N_1223);
or U1864 (N_1864,N_1660,N_1227);
and U1865 (N_1865,N_1600,N_1758);
xor U1866 (N_1866,N_1291,N_1728);
nand U1867 (N_1867,N_1240,N_1355);
xor U1868 (N_1868,N_1545,N_1715);
nand U1869 (N_1869,N_1371,N_1273);
nand U1870 (N_1870,N_1677,N_1603);
nand U1871 (N_1871,N_1322,N_1311);
nand U1872 (N_1872,N_1770,N_1348);
or U1873 (N_1873,N_1619,N_1200);
and U1874 (N_1874,N_1313,N_1581);
nor U1875 (N_1875,N_1280,N_1679);
nor U1876 (N_1876,N_1729,N_1312);
nand U1877 (N_1877,N_1380,N_1678);
or U1878 (N_1878,N_1231,N_1297);
and U1879 (N_1879,N_1310,N_1271);
nor U1880 (N_1880,N_1725,N_1671);
and U1881 (N_1881,N_1211,N_1441);
nand U1882 (N_1882,N_1282,N_1720);
nor U1883 (N_1883,N_1563,N_1334);
or U1884 (N_1884,N_1768,N_1341);
nor U1885 (N_1885,N_1762,N_1522);
and U1886 (N_1886,N_1481,N_1668);
nor U1887 (N_1887,N_1612,N_1450);
nand U1888 (N_1888,N_1764,N_1753);
or U1889 (N_1889,N_1533,N_1628);
and U1890 (N_1890,N_1247,N_1689);
and U1891 (N_1891,N_1473,N_1752);
or U1892 (N_1892,N_1651,N_1465);
or U1893 (N_1893,N_1432,N_1743);
and U1894 (N_1894,N_1398,N_1332);
nor U1895 (N_1895,N_1785,N_1646);
and U1896 (N_1896,N_1457,N_1702);
nand U1897 (N_1897,N_1385,N_1681);
nand U1898 (N_1898,N_1582,N_1399);
nand U1899 (N_1899,N_1431,N_1740);
nor U1900 (N_1900,N_1378,N_1727);
xnor U1901 (N_1901,N_1382,N_1384);
nor U1902 (N_1902,N_1598,N_1776);
and U1903 (N_1903,N_1700,N_1623);
or U1904 (N_1904,N_1552,N_1328);
nor U1905 (N_1905,N_1781,N_1407);
xor U1906 (N_1906,N_1640,N_1635);
nor U1907 (N_1907,N_1456,N_1249);
nand U1908 (N_1908,N_1553,N_1228);
nor U1909 (N_1909,N_1707,N_1251);
nand U1910 (N_1910,N_1440,N_1274);
nor U1911 (N_1911,N_1321,N_1281);
nand U1912 (N_1912,N_1622,N_1615);
and U1913 (N_1913,N_1480,N_1324);
xor U1914 (N_1914,N_1524,N_1656);
nand U1915 (N_1915,N_1453,N_1705);
and U1916 (N_1916,N_1601,N_1497);
nand U1917 (N_1917,N_1510,N_1493);
or U1918 (N_1918,N_1745,N_1760);
nor U1919 (N_1919,N_1537,N_1344);
xnor U1920 (N_1920,N_1516,N_1735);
nand U1921 (N_1921,N_1326,N_1518);
nor U1922 (N_1922,N_1508,N_1680);
nand U1923 (N_1923,N_1401,N_1246);
xnor U1924 (N_1924,N_1486,N_1302);
nor U1925 (N_1925,N_1591,N_1738);
nor U1926 (N_1926,N_1423,N_1495);
nor U1927 (N_1927,N_1222,N_1621);
or U1928 (N_1928,N_1579,N_1428);
or U1929 (N_1929,N_1704,N_1477);
xnor U1930 (N_1930,N_1444,N_1596);
nor U1931 (N_1931,N_1761,N_1425);
and U1932 (N_1932,N_1201,N_1525);
and U1933 (N_1933,N_1232,N_1597);
nand U1934 (N_1934,N_1790,N_1286);
or U1935 (N_1935,N_1396,N_1655);
and U1936 (N_1936,N_1784,N_1383);
xor U1937 (N_1937,N_1562,N_1756);
or U1938 (N_1938,N_1224,N_1734);
or U1939 (N_1939,N_1420,N_1484);
xor U1940 (N_1940,N_1265,N_1267);
nand U1941 (N_1941,N_1368,N_1605);
or U1942 (N_1942,N_1463,N_1577);
nor U1943 (N_1943,N_1233,N_1245);
nand U1944 (N_1944,N_1483,N_1400);
or U1945 (N_1945,N_1703,N_1695);
nand U1946 (N_1946,N_1346,N_1590);
nor U1947 (N_1947,N_1215,N_1305);
nand U1948 (N_1948,N_1206,N_1317);
nor U1949 (N_1949,N_1414,N_1664);
xnor U1950 (N_1950,N_1592,N_1774);
xor U1951 (N_1951,N_1716,N_1268);
nand U1952 (N_1952,N_1754,N_1470);
and U1953 (N_1953,N_1543,N_1257);
or U1954 (N_1954,N_1523,N_1212);
or U1955 (N_1955,N_1203,N_1229);
nand U1956 (N_1956,N_1674,N_1519);
xnor U1957 (N_1957,N_1666,N_1360);
nor U1958 (N_1958,N_1301,N_1277);
xnor U1959 (N_1959,N_1625,N_1649);
nand U1960 (N_1960,N_1712,N_1683);
nand U1961 (N_1961,N_1650,N_1672);
nor U1962 (N_1962,N_1218,N_1220);
nand U1963 (N_1963,N_1765,N_1634);
or U1964 (N_1964,N_1648,N_1541);
nand U1965 (N_1965,N_1636,N_1316);
and U1966 (N_1966,N_1609,N_1567);
nor U1967 (N_1967,N_1417,N_1352);
and U1968 (N_1968,N_1658,N_1763);
xnor U1969 (N_1969,N_1349,N_1759);
and U1970 (N_1970,N_1710,N_1418);
and U1971 (N_1971,N_1786,N_1430);
or U1972 (N_1972,N_1661,N_1285);
nor U1973 (N_1973,N_1565,N_1253);
and U1974 (N_1974,N_1487,N_1230);
nand U1975 (N_1975,N_1436,N_1733);
or U1976 (N_1976,N_1419,N_1377);
and U1977 (N_1977,N_1416,N_1732);
nand U1978 (N_1978,N_1340,N_1580);
nor U1979 (N_1979,N_1749,N_1306);
and U1980 (N_1980,N_1514,N_1427);
nor U1981 (N_1981,N_1616,N_1620);
xnor U1982 (N_1982,N_1507,N_1243);
and U1983 (N_1983,N_1354,N_1388);
and U1984 (N_1984,N_1300,N_1363);
xnor U1985 (N_1985,N_1792,N_1641);
and U1986 (N_1986,N_1584,N_1505);
xnor U1987 (N_1987,N_1410,N_1499);
or U1988 (N_1988,N_1325,N_1504);
and U1989 (N_1989,N_1652,N_1204);
and U1990 (N_1990,N_1594,N_1572);
and U1991 (N_1991,N_1358,N_1691);
and U1992 (N_1992,N_1290,N_1789);
nand U1993 (N_1993,N_1604,N_1284);
nand U1994 (N_1994,N_1529,N_1583);
and U1995 (N_1995,N_1461,N_1566);
or U1996 (N_1996,N_1708,N_1239);
xor U1997 (N_1997,N_1298,N_1624);
nand U1998 (N_1998,N_1568,N_1476);
or U1999 (N_1999,N_1278,N_1788);
nand U2000 (N_2000,N_1526,N_1376);
nand U2001 (N_2001,N_1351,N_1539);
or U2002 (N_2002,N_1730,N_1796);
or U2003 (N_2003,N_1775,N_1459);
xor U2004 (N_2004,N_1659,N_1373);
or U2005 (N_2005,N_1670,N_1381);
or U2006 (N_2006,N_1256,N_1455);
xnor U2007 (N_2007,N_1556,N_1475);
nand U2008 (N_2008,N_1248,N_1272);
or U2009 (N_2009,N_1488,N_1767);
nand U2010 (N_2010,N_1532,N_1527);
xnor U2011 (N_2011,N_1663,N_1535);
and U2012 (N_2012,N_1217,N_1602);
or U2013 (N_2013,N_1234,N_1304);
nor U2014 (N_2014,N_1460,N_1783);
and U2015 (N_2015,N_1294,N_1319);
nand U2016 (N_2016,N_1372,N_1357);
or U2017 (N_2017,N_1755,N_1585);
xnor U2018 (N_2018,N_1690,N_1237);
nand U2019 (N_2019,N_1451,N_1442);
and U2020 (N_2020,N_1662,N_1714);
and U2021 (N_2021,N_1778,N_1542);
and U2022 (N_2022,N_1769,N_1731);
nor U2023 (N_2023,N_1558,N_1511);
or U2024 (N_2024,N_1392,N_1467);
and U2025 (N_2025,N_1697,N_1327);
nor U2026 (N_2026,N_1438,N_1424);
or U2027 (N_2027,N_1213,N_1777);
nand U2028 (N_2028,N_1586,N_1506);
and U2029 (N_2029,N_1448,N_1547);
or U2030 (N_2030,N_1464,N_1242);
nor U2031 (N_2031,N_1718,N_1713);
nand U2032 (N_2032,N_1685,N_1362);
nand U2033 (N_2033,N_1787,N_1391);
xnor U2034 (N_2034,N_1613,N_1309);
nor U2035 (N_2035,N_1606,N_1314);
and U2036 (N_2036,N_1576,N_1561);
xnor U2037 (N_2037,N_1386,N_1421);
and U2038 (N_2038,N_1503,N_1269);
nand U2039 (N_2039,N_1462,N_1719);
nand U2040 (N_2040,N_1571,N_1536);
nand U2041 (N_2041,N_1501,N_1331);
xnor U2042 (N_2042,N_1447,N_1706);
or U2043 (N_2043,N_1261,N_1458);
and U2044 (N_2044,N_1335,N_1241);
and U2045 (N_2045,N_1687,N_1422);
nor U2046 (N_2046,N_1221,N_1644);
nor U2047 (N_2047,N_1263,N_1308);
nand U2048 (N_2048,N_1276,N_1474);
and U2049 (N_2049,N_1387,N_1574);
or U2050 (N_2050,N_1544,N_1560);
nand U2051 (N_2051,N_1548,N_1320);
nor U2052 (N_2052,N_1557,N_1657);
and U2053 (N_2053,N_1254,N_1250);
xnor U2054 (N_2054,N_1395,N_1342);
xnor U2055 (N_2055,N_1669,N_1405);
nand U2056 (N_2056,N_1403,N_1293);
nor U2057 (N_2057,N_1236,N_1701);
and U2058 (N_2058,N_1283,N_1772);
nor U2059 (N_2059,N_1653,N_1643);
nor U2060 (N_2060,N_1492,N_1588);
and U2061 (N_2061,N_1266,N_1303);
nor U2062 (N_2062,N_1747,N_1343);
nor U2063 (N_2063,N_1323,N_1608);
and U2064 (N_2064,N_1485,N_1512);
nand U2065 (N_2065,N_1361,N_1546);
nand U2066 (N_2066,N_1642,N_1578);
or U2067 (N_2067,N_1347,N_1534);
nand U2068 (N_2068,N_1684,N_1412);
and U2069 (N_2069,N_1370,N_1289);
nand U2070 (N_2070,N_1411,N_1375);
nand U2071 (N_2071,N_1336,N_1296);
or U2072 (N_2072,N_1717,N_1364);
or U2073 (N_2073,N_1665,N_1515);
or U2074 (N_2074,N_1575,N_1595);
nor U2075 (N_2075,N_1629,N_1433);
nand U2076 (N_2076,N_1279,N_1589);
nand U2077 (N_2077,N_1530,N_1449);
nor U2078 (N_2078,N_1737,N_1498);
nand U2079 (N_2079,N_1626,N_1502);
nand U2080 (N_2080,N_1333,N_1208);
nand U2081 (N_2081,N_1686,N_1292);
and U2082 (N_2082,N_1446,N_1466);
nor U2083 (N_2083,N_1750,N_1736);
and U2084 (N_2084,N_1550,N_1744);
nand U2085 (N_2085,N_1795,N_1494);
or U2086 (N_2086,N_1252,N_1682);
or U2087 (N_2087,N_1793,N_1654);
nand U2088 (N_2088,N_1202,N_1287);
or U2089 (N_2089,N_1454,N_1639);
nor U2090 (N_2090,N_1491,N_1587);
nand U2091 (N_2091,N_1238,N_1569);
or U2092 (N_2092,N_1205,N_1359);
or U2093 (N_2093,N_1742,N_1638);
nor U2094 (N_2094,N_1791,N_1549);
nor U2095 (N_2095,N_1339,N_1797);
nand U2096 (N_2096,N_1415,N_1722);
and U2097 (N_2097,N_1235,N_1637);
and U2098 (N_2098,N_1757,N_1698);
nor U2099 (N_2099,N_1413,N_1721);
nand U2100 (N_2100,N_1739,N_1603);
or U2101 (N_2101,N_1732,N_1762);
nand U2102 (N_2102,N_1654,N_1771);
nor U2103 (N_2103,N_1776,N_1681);
and U2104 (N_2104,N_1685,N_1337);
or U2105 (N_2105,N_1406,N_1414);
xor U2106 (N_2106,N_1508,N_1583);
or U2107 (N_2107,N_1769,N_1552);
nor U2108 (N_2108,N_1265,N_1251);
nand U2109 (N_2109,N_1794,N_1413);
xnor U2110 (N_2110,N_1522,N_1269);
and U2111 (N_2111,N_1725,N_1268);
nor U2112 (N_2112,N_1554,N_1729);
or U2113 (N_2113,N_1240,N_1469);
nor U2114 (N_2114,N_1338,N_1668);
and U2115 (N_2115,N_1731,N_1794);
or U2116 (N_2116,N_1578,N_1212);
xnor U2117 (N_2117,N_1495,N_1330);
xor U2118 (N_2118,N_1439,N_1799);
or U2119 (N_2119,N_1551,N_1606);
nor U2120 (N_2120,N_1259,N_1778);
and U2121 (N_2121,N_1793,N_1401);
or U2122 (N_2122,N_1450,N_1325);
or U2123 (N_2123,N_1452,N_1753);
nor U2124 (N_2124,N_1418,N_1581);
nand U2125 (N_2125,N_1432,N_1277);
nand U2126 (N_2126,N_1299,N_1621);
and U2127 (N_2127,N_1425,N_1276);
or U2128 (N_2128,N_1767,N_1333);
nand U2129 (N_2129,N_1556,N_1778);
nand U2130 (N_2130,N_1737,N_1271);
or U2131 (N_2131,N_1776,N_1602);
or U2132 (N_2132,N_1276,N_1538);
and U2133 (N_2133,N_1670,N_1568);
or U2134 (N_2134,N_1424,N_1550);
or U2135 (N_2135,N_1366,N_1381);
and U2136 (N_2136,N_1295,N_1398);
or U2137 (N_2137,N_1513,N_1534);
or U2138 (N_2138,N_1395,N_1314);
nor U2139 (N_2139,N_1738,N_1519);
and U2140 (N_2140,N_1694,N_1340);
or U2141 (N_2141,N_1443,N_1758);
nand U2142 (N_2142,N_1559,N_1673);
nand U2143 (N_2143,N_1207,N_1739);
nand U2144 (N_2144,N_1739,N_1234);
or U2145 (N_2145,N_1670,N_1236);
nor U2146 (N_2146,N_1732,N_1240);
nor U2147 (N_2147,N_1442,N_1634);
nand U2148 (N_2148,N_1680,N_1223);
and U2149 (N_2149,N_1245,N_1434);
or U2150 (N_2150,N_1550,N_1730);
or U2151 (N_2151,N_1474,N_1410);
nand U2152 (N_2152,N_1236,N_1650);
nand U2153 (N_2153,N_1700,N_1445);
or U2154 (N_2154,N_1726,N_1754);
xor U2155 (N_2155,N_1636,N_1448);
nand U2156 (N_2156,N_1347,N_1276);
and U2157 (N_2157,N_1202,N_1734);
or U2158 (N_2158,N_1630,N_1352);
or U2159 (N_2159,N_1291,N_1710);
nand U2160 (N_2160,N_1363,N_1622);
and U2161 (N_2161,N_1328,N_1293);
or U2162 (N_2162,N_1223,N_1257);
nand U2163 (N_2163,N_1255,N_1538);
nand U2164 (N_2164,N_1300,N_1396);
nand U2165 (N_2165,N_1691,N_1529);
or U2166 (N_2166,N_1232,N_1440);
and U2167 (N_2167,N_1230,N_1338);
and U2168 (N_2168,N_1681,N_1441);
and U2169 (N_2169,N_1347,N_1209);
xor U2170 (N_2170,N_1229,N_1291);
and U2171 (N_2171,N_1332,N_1469);
nand U2172 (N_2172,N_1414,N_1269);
or U2173 (N_2173,N_1666,N_1618);
and U2174 (N_2174,N_1789,N_1678);
nand U2175 (N_2175,N_1470,N_1683);
nor U2176 (N_2176,N_1758,N_1785);
nand U2177 (N_2177,N_1510,N_1465);
and U2178 (N_2178,N_1684,N_1323);
nor U2179 (N_2179,N_1379,N_1579);
nand U2180 (N_2180,N_1617,N_1435);
nand U2181 (N_2181,N_1255,N_1357);
and U2182 (N_2182,N_1273,N_1260);
nand U2183 (N_2183,N_1683,N_1418);
nor U2184 (N_2184,N_1353,N_1365);
nor U2185 (N_2185,N_1474,N_1677);
and U2186 (N_2186,N_1286,N_1725);
and U2187 (N_2187,N_1449,N_1778);
nor U2188 (N_2188,N_1716,N_1771);
nor U2189 (N_2189,N_1795,N_1734);
nor U2190 (N_2190,N_1675,N_1238);
nand U2191 (N_2191,N_1533,N_1208);
and U2192 (N_2192,N_1751,N_1798);
or U2193 (N_2193,N_1664,N_1552);
or U2194 (N_2194,N_1536,N_1542);
or U2195 (N_2195,N_1223,N_1561);
nand U2196 (N_2196,N_1286,N_1264);
or U2197 (N_2197,N_1554,N_1219);
nor U2198 (N_2198,N_1223,N_1716);
and U2199 (N_2199,N_1201,N_1215);
nand U2200 (N_2200,N_1336,N_1450);
or U2201 (N_2201,N_1354,N_1726);
or U2202 (N_2202,N_1513,N_1270);
xor U2203 (N_2203,N_1713,N_1785);
or U2204 (N_2204,N_1394,N_1478);
and U2205 (N_2205,N_1271,N_1407);
and U2206 (N_2206,N_1592,N_1478);
or U2207 (N_2207,N_1729,N_1459);
nor U2208 (N_2208,N_1778,N_1455);
and U2209 (N_2209,N_1233,N_1277);
or U2210 (N_2210,N_1620,N_1295);
xnor U2211 (N_2211,N_1305,N_1738);
or U2212 (N_2212,N_1555,N_1565);
and U2213 (N_2213,N_1280,N_1640);
nand U2214 (N_2214,N_1698,N_1218);
or U2215 (N_2215,N_1772,N_1649);
xnor U2216 (N_2216,N_1644,N_1544);
nand U2217 (N_2217,N_1516,N_1289);
nand U2218 (N_2218,N_1634,N_1632);
or U2219 (N_2219,N_1230,N_1307);
or U2220 (N_2220,N_1749,N_1603);
nor U2221 (N_2221,N_1358,N_1654);
and U2222 (N_2222,N_1662,N_1362);
and U2223 (N_2223,N_1739,N_1615);
nand U2224 (N_2224,N_1223,N_1398);
or U2225 (N_2225,N_1370,N_1754);
or U2226 (N_2226,N_1328,N_1468);
xnor U2227 (N_2227,N_1279,N_1448);
nor U2228 (N_2228,N_1341,N_1271);
nand U2229 (N_2229,N_1459,N_1533);
nor U2230 (N_2230,N_1388,N_1489);
and U2231 (N_2231,N_1774,N_1419);
and U2232 (N_2232,N_1561,N_1756);
nor U2233 (N_2233,N_1271,N_1759);
and U2234 (N_2234,N_1375,N_1204);
nand U2235 (N_2235,N_1385,N_1510);
xnor U2236 (N_2236,N_1756,N_1222);
nor U2237 (N_2237,N_1445,N_1708);
or U2238 (N_2238,N_1674,N_1520);
nor U2239 (N_2239,N_1265,N_1263);
or U2240 (N_2240,N_1705,N_1355);
xnor U2241 (N_2241,N_1545,N_1757);
nand U2242 (N_2242,N_1711,N_1573);
or U2243 (N_2243,N_1300,N_1596);
nand U2244 (N_2244,N_1391,N_1681);
nand U2245 (N_2245,N_1464,N_1745);
xnor U2246 (N_2246,N_1774,N_1349);
xnor U2247 (N_2247,N_1547,N_1556);
nor U2248 (N_2248,N_1261,N_1763);
xnor U2249 (N_2249,N_1696,N_1734);
nor U2250 (N_2250,N_1757,N_1403);
nor U2251 (N_2251,N_1470,N_1235);
or U2252 (N_2252,N_1345,N_1660);
and U2253 (N_2253,N_1252,N_1417);
nor U2254 (N_2254,N_1708,N_1471);
nand U2255 (N_2255,N_1743,N_1653);
nand U2256 (N_2256,N_1356,N_1548);
and U2257 (N_2257,N_1503,N_1459);
nor U2258 (N_2258,N_1356,N_1781);
nor U2259 (N_2259,N_1311,N_1658);
nand U2260 (N_2260,N_1559,N_1588);
or U2261 (N_2261,N_1612,N_1206);
xor U2262 (N_2262,N_1503,N_1754);
nand U2263 (N_2263,N_1411,N_1640);
nor U2264 (N_2264,N_1462,N_1210);
or U2265 (N_2265,N_1796,N_1716);
or U2266 (N_2266,N_1541,N_1790);
nor U2267 (N_2267,N_1307,N_1535);
or U2268 (N_2268,N_1507,N_1339);
nand U2269 (N_2269,N_1249,N_1766);
nor U2270 (N_2270,N_1283,N_1710);
and U2271 (N_2271,N_1477,N_1574);
and U2272 (N_2272,N_1349,N_1534);
nand U2273 (N_2273,N_1239,N_1616);
and U2274 (N_2274,N_1332,N_1301);
nor U2275 (N_2275,N_1455,N_1496);
nor U2276 (N_2276,N_1638,N_1339);
nor U2277 (N_2277,N_1702,N_1418);
xnor U2278 (N_2278,N_1396,N_1200);
nand U2279 (N_2279,N_1674,N_1273);
nand U2280 (N_2280,N_1733,N_1668);
and U2281 (N_2281,N_1634,N_1717);
and U2282 (N_2282,N_1780,N_1404);
or U2283 (N_2283,N_1568,N_1282);
nand U2284 (N_2284,N_1790,N_1770);
nand U2285 (N_2285,N_1715,N_1250);
and U2286 (N_2286,N_1342,N_1285);
or U2287 (N_2287,N_1319,N_1229);
or U2288 (N_2288,N_1592,N_1676);
nand U2289 (N_2289,N_1230,N_1591);
nor U2290 (N_2290,N_1350,N_1677);
or U2291 (N_2291,N_1478,N_1279);
nor U2292 (N_2292,N_1700,N_1489);
and U2293 (N_2293,N_1317,N_1791);
xnor U2294 (N_2294,N_1665,N_1317);
or U2295 (N_2295,N_1714,N_1716);
or U2296 (N_2296,N_1550,N_1394);
nor U2297 (N_2297,N_1424,N_1796);
and U2298 (N_2298,N_1276,N_1242);
nand U2299 (N_2299,N_1226,N_1490);
or U2300 (N_2300,N_1567,N_1301);
and U2301 (N_2301,N_1738,N_1637);
nand U2302 (N_2302,N_1244,N_1401);
nand U2303 (N_2303,N_1309,N_1278);
and U2304 (N_2304,N_1239,N_1518);
nor U2305 (N_2305,N_1246,N_1777);
nand U2306 (N_2306,N_1280,N_1609);
nand U2307 (N_2307,N_1270,N_1279);
nor U2308 (N_2308,N_1393,N_1555);
and U2309 (N_2309,N_1488,N_1284);
nand U2310 (N_2310,N_1785,N_1668);
and U2311 (N_2311,N_1711,N_1232);
and U2312 (N_2312,N_1658,N_1466);
or U2313 (N_2313,N_1280,N_1255);
nand U2314 (N_2314,N_1339,N_1309);
nand U2315 (N_2315,N_1427,N_1385);
nor U2316 (N_2316,N_1206,N_1369);
nand U2317 (N_2317,N_1250,N_1330);
and U2318 (N_2318,N_1616,N_1512);
or U2319 (N_2319,N_1307,N_1581);
and U2320 (N_2320,N_1228,N_1504);
nor U2321 (N_2321,N_1704,N_1367);
nor U2322 (N_2322,N_1715,N_1632);
nor U2323 (N_2323,N_1335,N_1699);
nand U2324 (N_2324,N_1353,N_1461);
nand U2325 (N_2325,N_1771,N_1468);
and U2326 (N_2326,N_1769,N_1702);
xor U2327 (N_2327,N_1202,N_1542);
or U2328 (N_2328,N_1770,N_1387);
nor U2329 (N_2329,N_1664,N_1200);
and U2330 (N_2330,N_1496,N_1762);
nor U2331 (N_2331,N_1752,N_1243);
or U2332 (N_2332,N_1773,N_1369);
nor U2333 (N_2333,N_1360,N_1251);
nor U2334 (N_2334,N_1416,N_1417);
nand U2335 (N_2335,N_1467,N_1502);
and U2336 (N_2336,N_1731,N_1296);
and U2337 (N_2337,N_1433,N_1782);
nor U2338 (N_2338,N_1790,N_1485);
and U2339 (N_2339,N_1620,N_1596);
nand U2340 (N_2340,N_1629,N_1575);
nand U2341 (N_2341,N_1763,N_1390);
nand U2342 (N_2342,N_1329,N_1520);
nand U2343 (N_2343,N_1588,N_1487);
nor U2344 (N_2344,N_1460,N_1668);
or U2345 (N_2345,N_1729,N_1534);
nand U2346 (N_2346,N_1604,N_1471);
nor U2347 (N_2347,N_1451,N_1746);
or U2348 (N_2348,N_1351,N_1340);
nand U2349 (N_2349,N_1753,N_1339);
nor U2350 (N_2350,N_1490,N_1694);
or U2351 (N_2351,N_1311,N_1294);
or U2352 (N_2352,N_1666,N_1239);
nor U2353 (N_2353,N_1346,N_1768);
nor U2354 (N_2354,N_1372,N_1550);
and U2355 (N_2355,N_1636,N_1760);
xor U2356 (N_2356,N_1444,N_1527);
and U2357 (N_2357,N_1733,N_1333);
and U2358 (N_2358,N_1751,N_1541);
xor U2359 (N_2359,N_1419,N_1223);
nor U2360 (N_2360,N_1664,N_1213);
xor U2361 (N_2361,N_1741,N_1311);
nand U2362 (N_2362,N_1602,N_1516);
and U2363 (N_2363,N_1770,N_1729);
and U2364 (N_2364,N_1769,N_1304);
and U2365 (N_2365,N_1550,N_1286);
nor U2366 (N_2366,N_1589,N_1536);
nand U2367 (N_2367,N_1738,N_1249);
xor U2368 (N_2368,N_1336,N_1437);
and U2369 (N_2369,N_1691,N_1798);
or U2370 (N_2370,N_1691,N_1612);
and U2371 (N_2371,N_1355,N_1767);
and U2372 (N_2372,N_1239,N_1210);
or U2373 (N_2373,N_1466,N_1405);
and U2374 (N_2374,N_1598,N_1389);
nand U2375 (N_2375,N_1413,N_1426);
xor U2376 (N_2376,N_1243,N_1590);
and U2377 (N_2377,N_1768,N_1436);
nor U2378 (N_2378,N_1663,N_1615);
nand U2379 (N_2379,N_1206,N_1467);
or U2380 (N_2380,N_1715,N_1563);
and U2381 (N_2381,N_1451,N_1371);
or U2382 (N_2382,N_1602,N_1597);
nand U2383 (N_2383,N_1403,N_1383);
xnor U2384 (N_2384,N_1274,N_1262);
and U2385 (N_2385,N_1574,N_1669);
or U2386 (N_2386,N_1628,N_1785);
and U2387 (N_2387,N_1539,N_1640);
xnor U2388 (N_2388,N_1736,N_1251);
nor U2389 (N_2389,N_1355,N_1526);
nand U2390 (N_2390,N_1760,N_1376);
nand U2391 (N_2391,N_1244,N_1448);
nand U2392 (N_2392,N_1706,N_1552);
nand U2393 (N_2393,N_1520,N_1521);
and U2394 (N_2394,N_1733,N_1244);
xor U2395 (N_2395,N_1630,N_1311);
nand U2396 (N_2396,N_1659,N_1678);
or U2397 (N_2397,N_1343,N_1415);
nor U2398 (N_2398,N_1547,N_1409);
and U2399 (N_2399,N_1608,N_1217);
or U2400 (N_2400,N_2149,N_2074);
xor U2401 (N_2401,N_2263,N_2274);
nor U2402 (N_2402,N_2359,N_1927);
and U2403 (N_2403,N_1851,N_1819);
nand U2404 (N_2404,N_1922,N_2285);
and U2405 (N_2405,N_1946,N_1864);
nand U2406 (N_2406,N_2353,N_2195);
nand U2407 (N_2407,N_1847,N_1941);
nand U2408 (N_2408,N_2165,N_2270);
and U2409 (N_2409,N_2305,N_2054);
nand U2410 (N_2410,N_2355,N_2181);
xnor U2411 (N_2411,N_1848,N_1892);
nor U2412 (N_2412,N_1829,N_2362);
nand U2413 (N_2413,N_1950,N_2255);
nor U2414 (N_2414,N_2217,N_1913);
nor U2415 (N_2415,N_1965,N_2053);
or U2416 (N_2416,N_2135,N_2326);
nand U2417 (N_2417,N_1904,N_1889);
xnor U2418 (N_2418,N_2347,N_1866);
or U2419 (N_2419,N_2016,N_2279);
and U2420 (N_2420,N_1880,N_2090);
xnor U2421 (N_2421,N_2095,N_2057);
and U2422 (N_2422,N_2341,N_2369);
nor U2423 (N_2423,N_1938,N_2246);
nand U2424 (N_2424,N_2184,N_1919);
nor U2425 (N_2425,N_2373,N_1955);
nor U2426 (N_2426,N_2049,N_2204);
nor U2427 (N_2427,N_2121,N_2137);
and U2428 (N_2428,N_1807,N_1850);
nand U2429 (N_2429,N_2360,N_1839);
nor U2430 (N_2430,N_2162,N_2310);
and U2431 (N_2431,N_2019,N_2280);
nor U2432 (N_2432,N_2343,N_2323);
xnor U2433 (N_2433,N_1909,N_2237);
and U2434 (N_2434,N_2157,N_1846);
or U2435 (N_2435,N_1936,N_1893);
and U2436 (N_2436,N_1809,N_1818);
xnor U2437 (N_2437,N_2133,N_1981);
and U2438 (N_2438,N_2115,N_1920);
nand U2439 (N_2439,N_1887,N_2221);
nor U2440 (N_2440,N_2180,N_2236);
nor U2441 (N_2441,N_2116,N_2006);
or U2442 (N_2442,N_2234,N_2030);
and U2443 (N_2443,N_2108,N_1930);
nand U2444 (N_2444,N_2003,N_1836);
nor U2445 (N_2445,N_2245,N_2015);
and U2446 (N_2446,N_1817,N_1979);
nor U2447 (N_2447,N_2174,N_1952);
and U2448 (N_2448,N_1934,N_1823);
nor U2449 (N_2449,N_2242,N_2391);
nand U2450 (N_2450,N_2366,N_2123);
or U2451 (N_2451,N_2315,N_1959);
nor U2452 (N_2452,N_1951,N_1947);
nand U2453 (N_2453,N_2307,N_1885);
or U2454 (N_2454,N_1853,N_2004);
xor U2455 (N_2455,N_1993,N_2260);
and U2456 (N_2456,N_2073,N_2379);
nand U2457 (N_2457,N_1816,N_2088);
nor U2458 (N_2458,N_1967,N_2002);
or U2459 (N_2459,N_2119,N_1970);
nor U2460 (N_2460,N_2316,N_1805);
nand U2461 (N_2461,N_2365,N_2027);
nor U2462 (N_2462,N_2051,N_2215);
or U2463 (N_2463,N_2388,N_2339);
nand U2464 (N_2464,N_1921,N_2302);
nor U2465 (N_2465,N_2346,N_2202);
nand U2466 (N_2466,N_1837,N_1935);
and U2467 (N_2467,N_2257,N_2164);
and U2468 (N_2468,N_2251,N_2120);
xor U2469 (N_2469,N_2161,N_1808);
or U2470 (N_2470,N_1803,N_2044);
or U2471 (N_2471,N_1960,N_2342);
nor U2472 (N_2472,N_1821,N_2062);
nand U2473 (N_2473,N_2334,N_2079);
and U2474 (N_2474,N_1813,N_1881);
and U2475 (N_2475,N_1976,N_2324);
nand U2476 (N_2476,N_2083,N_2213);
or U2477 (N_2477,N_1982,N_1856);
or U2478 (N_2478,N_2264,N_2041);
nor U2479 (N_2479,N_2167,N_1971);
and U2480 (N_2480,N_2332,N_1980);
nor U2481 (N_2481,N_2086,N_1928);
nand U2482 (N_2482,N_2289,N_1958);
or U2483 (N_2483,N_1859,N_1804);
or U2484 (N_2484,N_2265,N_2013);
xnor U2485 (N_2485,N_2144,N_2380);
or U2486 (N_2486,N_1869,N_2278);
nor U2487 (N_2487,N_2361,N_1868);
or U2488 (N_2488,N_2386,N_1814);
or U2489 (N_2489,N_2210,N_1800);
and U2490 (N_2490,N_2169,N_2387);
or U2491 (N_2491,N_1924,N_1992);
nor U2492 (N_2492,N_1974,N_2239);
or U2493 (N_2493,N_1978,N_1811);
nor U2494 (N_2494,N_2099,N_2080);
nand U2495 (N_2495,N_2141,N_2189);
nor U2496 (N_2496,N_2170,N_2131);
nand U2497 (N_2497,N_2291,N_1871);
or U2498 (N_2498,N_2224,N_2211);
xor U2499 (N_2499,N_1945,N_1908);
and U2500 (N_2500,N_2309,N_2018);
and U2501 (N_2501,N_1882,N_1876);
or U2502 (N_2502,N_1875,N_2105);
and U2503 (N_2503,N_1991,N_1990);
and U2504 (N_2504,N_2244,N_1940);
or U2505 (N_2505,N_2089,N_2394);
nand U2506 (N_2506,N_2314,N_2322);
or U2507 (N_2507,N_2273,N_2381);
or U2508 (N_2508,N_2091,N_2025);
nand U2509 (N_2509,N_2101,N_1977);
or U2510 (N_2510,N_2150,N_1884);
nand U2511 (N_2511,N_2243,N_2094);
or U2512 (N_2512,N_2209,N_2038);
and U2513 (N_2513,N_1827,N_2070);
nand U2514 (N_2514,N_2190,N_2392);
or U2515 (N_2515,N_2103,N_2194);
and U2516 (N_2516,N_2299,N_2093);
nor U2517 (N_2517,N_2331,N_1999);
or U2518 (N_2518,N_2247,N_2061);
nor U2519 (N_2519,N_1983,N_2232);
nand U2520 (N_2520,N_2179,N_2153);
or U2521 (N_2521,N_2142,N_1828);
nand U2522 (N_2522,N_2029,N_1943);
or U2523 (N_2523,N_2039,N_1956);
nand U2524 (N_2524,N_2329,N_1831);
and U2525 (N_2525,N_2327,N_2222);
or U2526 (N_2526,N_1933,N_1989);
and U2527 (N_2527,N_2201,N_2178);
nor U2528 (N_2528,N_1898,N_2338);
nor U2529 (N_2529,N_2068,N_1812);
nand U2530 (N_2530,N_1929,N_1902);
and U2531 (N_2531,N_2176,N_2376);
or U2532 (N_2532,N_2272,N_1961);
and U2533 (N_2533,N_1857,N_2253);
nand U2534 (N_2534,N_1824,N_2009);
or U2535 (N_2535,N_2098,N_2218);
nor U2536 (N_2536,N_2235,N_1860);
or U2537 (N_2537,N_2117,N_1877);
and U2538 (N_2538,N_2125,N_2275);
xor U2539 (N_2539,N_2127,N_2320);
or U2540 (N_2540,N_2036,N_2156);
nor U2541 (N_2541,N_2367,N_1833);
and U2542 (N_2542,N_2146,N_1835);
nor U2543 (N_2543,N_2058,N_2357);
xnor U2544 (N_2544,N_2024,N_1916);
and U2545 (N_2545,N_1964,N_2198);
and U2546 (N_2546,N_2321,N_2206);
or U2547 (N_2547,N_2350,N_1858);
xnor U2548 (N_2548,N_1832,N_2268);
xnor U2549 (N_2549,N_2032,N_1843);
nand U2550 (N_2550,N_1942,N_2269);
and U2551 (N_2551,N_1874,N_1997);
and U2552 (N_2552,N_2196,N_2021);
and U2553 (N_2553,N_2152,N_2050);
nor U2554 (N_2554,N_2216,N_2071);
nand U2555 (N_2555,N_1988,N_2191);
nor U2556 (N_2556,N_1912,N_2294);
and U2557 (N_2557,N_2318,N_2284);
or U2558 (N_2558,N_2092,N_1870);
nand U2559 (N_2559,N_1825,N_1998);
nand U2560 (N_2560,N_2220,N_2066);
nor U2561 (N_2561,N_2111,N_2296);
nand U2562 (N_2562,N_2226,N_2182);
nor U2563 (N_2563,N_2124,N_2319);
and U2564 (N_2564,N_2077,N_1901);
nor U2565 (N_2565,N_2122,N_2109);
or U2566 (N_2566,N_2076,N_1822);
xor U2567 (N_2567,N_1899,N_2056);
and U2568 (N_2568,N_2389,N_2290);
xor U2569 (N_2569,N_2328,N_2147);
nand U2570 (N_2570,N_2107,N_2301);
or U2571 (N_2571,N_1830,N_2052);
nor U2572 (N_2572,N_2261,N_2212);
nor U2573 (N_2573,N_2102,N_1954);
nor U2574 (N_2574,N_2340,N_2214);
and U2575 (N_2575,N_2085,N_1939);
or U2576 (N_2576,N_2283,N_2040);
or U2577 (N_2577,N_2368,N_1886);
nand U2578 (N_2578,N_2288,N_2011);
nand U2579 (N_2579,N_1968,N_2172);
nand U2580 (N_2580,N_2370,N_2185);
or U2581 (N_2581,N_1925,N_2267);
nor U2582 (N_2582,N_1944,N_1996);
nand U2583 (N_2583,N_2072,N_2081);
nand U2584 (N_2584,N_2292,N_2129);
nor U2585 (N_2585,N_2037,N_2205);
nor U2586 (N_2586,N_2330,N_2110);
and U2587 (N_2587,N_2100,N_1897);
and U2588 (N_2588,N_1986,N_2384);
and U2589 (N_2589,N_2026,N_2254);
nor U2590 (N_2590,N_2140,N_2000);
nand U2591 (N_2591,N_1973,N_2317);
and U2592 (N_2592,N_2155,N_1948);
nand U2593 (N_2593,N_2145,N_2344);
and U2594 (N_2594,N_2020,N_2397);
or U2595 (N_2595,N_2060,N_1826);
nor U2596 (N_2596,N_2023,N_2175);
nand U2597 (N_2597,N_2252,N_2033);
nor U2598 (N_2598,N_2014,N_1995);
or U2599 (N_2599,N_1895,N_2393);
nand U2600 (N_2600,N_1855,N_1914);
xor U2601 (N_2601,N_2064,N_2250);
and U2602 (N_2602,N_1917,N_2047);
or U2603 (N_2603,N_2306,N_2240);
or U2604 (N_2604,N_2303,N_1863);
and U2605 (N_2605,N_2227,N_2312);
nand U2606 (N_2606,N_2114,N_2112);
and U2607 (N_2607,N_2199,N_1903);
nor U2608 (N_2608,N_2345,N_2304);
and U2609 (N_2609,N_1985,N_1879);
nor U2610 (N_2610,N_2063,N_2363);
and U2611 (N_2611,N_2390,N_2277);
nor U2612 (N_2612,N_2262,N_2385);
or U2613 (N_2613,N_1883,N_2241);
or U2614 (N_2614,N_2351,N_2354);
xnor U2615 (N_2615,N_1878,N_2168);
or U2616 (N_2616,N_1911,N_2139);
nor U2617 (N_2617,N_2042,N_1810);
nor U2618 (N_2618,N_2130,N_2249);
or U2619 (N_2619,N_2067,N_2007);
xor U2620 (N_2620,N_1842,N_2228);
or U2621 (N_2621,N_1834,N_2231);
or U2622 (N_2622,N_2183,N_2046);
nand U2623 (N_2623,N_2356,N_2087);
and U2624 (N_2624,N_2106,N_1918);
and U2625 (N_2625,N_2035,N_2266);
nand U2626 (N_2626,N_2177,N_2300);
nand U2627 (N_2627,N_2143,N_2096);
nor U2628 (N_2628,N_1894,N_2219);
or U2629 (N_2629,N_2311,N_2372);
and U2630 (N_2630,N_2364,N_1854);
nor U2631 (N_2631,N_2282,N_1861);
nand U2632 (N_2632,N_1891,N_1926);
and U2633 (N_2633,N_2259,N_2358);
xor U2634 (N_2634,N_2010,N_2118);
or U2635 (N_2635,N_1910,N_2148);
nor U2636 (N_2636,N_2012,N_2333);
and U2637 (N_2637,N_2078,N_1852);
or U2638 (N_2638,N_1845,N_2097);
and U2639 (N_2639,N_1872,N_2225);
nor U2640 (N_2640,N_2293,N_1867);
or U2641 (N_2641,N_2193,N_2043);
and U2642 (N_2642,N_1994,N_2271);
xor U2643 (N_2643,N_1900,N_2017);
nand U2644 (N_2644,N_2286,N_1838);
or U2645 (N_2645,N_1969,N_2337);
nor U2646 (N_2646,N_2151,N_2138);
and U2647 (N_2647,N_2297,N_1957);
and U2648 (N_2648,N_1931,N_2154);
xor U2649 (N_2649,N_2160,N_2313);
and U2650 (N_2650,N_2163,N_1953);
nor U2651 (N_2651,N_2171,N_2034);
or U2652 (N_2652,N_1820,N_2377);
or U2653 (N_2653,N_1975,N_1849);
nor U2654 (N_2654,N_1806,N_2069);
xor U2655 (N_2655,N_2197,N_2208);
or U2656 (N_2656,N_2159,N_1962);
or U2657 (N_2657,N_1801,N_2001);
nand U2658 (N_2658,N_2383,N_2349);
and U2659 (N_2659,N_1815,N_2203);
and U2660 (N_2660,N_2128,N_2396);
nand U2661 (N_2661,N_2104,N_2045);
and U2662 (N_2662,N_2382,N_1865);
nand U2663 (N_2663,N_2200,N_2113);
nand U2664 (N_2664,N_2336,N_2188);
nor U2665 (N_2665,N_2158,N_2082);
nor U2666 (N_2666,N_2048,N_1972);
xnor U2667 (N_2667,N_1923,N_2031);
or U2668 (N_2668,N_2005,N_2186);
and U2669 (N_2669,N_1890,N_1905);
nor U2670 (N_2670,N_2065,N_2075);
and U2671 (N_2671,N_2371,N_2375);
nor U2672 (N_2672,N_2258,N_2256);
nor U2673 (N_2673,N_1841,N_2238);
nor U2674 (N_2674,N_2192,N_2223);
nand U2675 (N_2675,N_2325,N_2132);
or U2676 (N_2676,N_1896,N_1862);
nor U2677 (N_2677,N_2348,N_1966);
nand U2678 (N_2678,N_2248,N_2276);
and U2679 (N_2679,N_2028,N_1907);
xnor U2680 (N_2680,N_2173,N_1984);
nand U2681 (N_2681,N_2287,N_1873);
nand U2682 (N_2682,N_1906,N_2352);
nor U2683 (N_2683,N_1937,N_1963);
nand U2684 (N_2684,N_2008,N_2298);
nor U2685 (N_2685,N_2229,N_2399);
or U2686 (N_2686,N_2126,N_2295);
or U2687 (N_2687,N_2308,N_2134);
nor U2688 (N_2688,N_2207,N_2022);
nand U2689 (N_2689,N_2136,N_1915);
xor U2690 (N_2690,N_1949,N_2187);
and U2691 (N_2691,N_2335,N_1888);
nor U2692 (N_2692,N_2378,N_2374);
xor U2693 (N_2693,N_1802,N_1987);
and U2694 (N_2694,N_2398,N_2055);
and U2695 (N_2695,N_2084,N_2233);
xnor U2696 (N_2696,N_2281,N_1932);
xor U2697 (N_2697,N_2395,N_2059);
or U2698 (N_2698,N_2230,N_1844);
nor U2699 (N_2699,N_2166,N_1840);
nor U2700 (N_2700,N_2038,N_2046);
xnor U2701 (N_2701,N_1933,N_1854);
and U2702 (N_2702,N_2113,N_2182);
nor U2703 (N_2703,N_1807,N_1953);
nor U2704 (N_2704,N_1857,N_1917);
and U2705 (N_2705,N_1860,N_1940);
and U2706 (N_2706,N_2060,N_2108);
nand U2707 (N_2707,N_2300,N_2389);
or U2708 (N_2708,N_2071,N_2227);
or U2709 (N_2709,N_2025,N_2020);
nand U2710 (N_2710,N_1928,N_2000);
nor U2711 (N_2711,N_2380,N_1924);
and U2712 (N_2712,N_2020,N_1891);
nor U2713 (N_2713,N_2370,N_1906);
and U2714 (N_2714,N_1889,N_2177);
or U2715 (N_2715,N_2208,N_2255);
nand U2716 (N_2716,N_1891,N_1942);
or U2717 (N_2717,N_2159,N_2338);
or U2718 (N_2718,N_2087,N_2184);
nand U2719 (N_2719,N_2088,N_2066);
nand U2720 (N_2720,N_1935,N_2068);
or U2721 (N_2721,N_1947,N_2097);
nand U2722 (N_2722,N_1882,N_2138);
nand U2723 (N_2723,N_2230,N_2206);
nor U2724 (N_2724,N_2101,N_2034);
nand U2725 (N_2725,N_2148,N_2088);
or U2726 (N_2726,N_2395,N_2311);
nand U2727 (N_2727,N_2229,N_1940);
and U2728 (N_2728,N_2355,N_2399);
nor U2729 (N_2729,N_1919,N_2246);
nor U2730 (N_2730,N_1885,N_2394);
and U2731 (N_2731,N_2048,N_2128);
nand U2732 (N_2732,N_2206,N_2264);
or U2733 (N_2733,N_2206,N_2149);
nor U2734 (N_2734,N_2045,N_2298);
or U2735 (N_2735,N_1901,N_2040);
nand U2736 (N_2736,N_2106,N_2267);
nor U2737 (N_2737,N_2244,N_2349);
and U2738 (N_2738,N_2390,N_2248);
nand U2739 (N_2739,N_2176,N_2083);
or U2740 (N_2740,N_1958,N_1998);
nor U2741 (N_2741,N_2193,N_2315);
nand U2742 (N_2742,N_2350,N_1908);
nor U2743 (N_2743,N_2243,N_2154);
nor U2744 (N_2744,N_1884,N_2018);
xor U2745 (N_2745,N_2156,N_2305);
nor U2746 (N_2746,N_1802,N_2148);
and U2747 (N_2747,N_2198,N_1816);
or U2748 (N_2748,N_1945,N_1868);
and U2749 (N_2749,N_1888,N_2193);
nand U2750 (N_2750,N_2024,N_2080);
nand U2751 (N_2751,N_2162,N_2102);
or U2752 (N_2752,N_1890,N_2272);
or U2753 (N_2753,N_1941,N_1977);
xnor U2754 (N_2754,N_2120,N_2194);
nand U2755 (N_2755,N_2260,N_1846);
and U2756 (N_2756,N_1976,N_2084);
and U2757 (N_2757,N_1979,N_1801);
nor U2758 (N_2758,N_2233,N_1961);
or U2759 (N_2759,N_2366,N_2068);
nor U2760 (N_2760,N_2088,N_2374);
or U2761 (N_2761,N_2138,N_2274);
xnor U2762 (N_2762,N_1919,N_2370);
and U2763 (N_2763,N_1901,N_1870);
and U2764 (N_2764,N_2218,N_2255);
nor U2765 (N_2765,N_2242,N_1938);
and U2766 (N_2766,N_1912,N_1978);
nand U2767 (N_2767,N_2186,N_2104);
or U2768 (N_2768,N_2393,N_2318);
nand U2769 (N_2769,N_2369,N_1962);
nor U2770 (N_2770,N_2155,N_2240);
or U2771 (N_2771,N_2158,N_2251);
and U2772 (N_2772,N_1943,N_2223);
nor U2773 (N_2773,N_2076,N_1898);
nand U2774 (N_2774,N_1814,N_2108);
nand U2775 (N_2775,N_2055,N_1906);
and U2776 (N_2776,N_2135,N_2106);
or U2777 (N_2777,N_2061,N_1947);
xor U2778 (N_2778,N_2197,N_2229);
nand U2779 (N_2779,N_1983,N_2325);
and U2780 (N_2780,N_2208,N_2268);
nor U2781 (N_2781,N_2064,N_1929);
and U2782 (N_2782,N_2202,N_2187);
xor U2783 (N_2783,N_2136,N_1995);
nand U2784 (N_2784,N_2352,N_1860);
and U2785 (N_2785,N_2158,N_2337);
and U2786 (N_2786,N_2143,N_2391);
or U2787 (N_2787,N_2386,N_1810);
nand U2788 (N_2788,N_1837,N_1905);
or U2789 (N_2789,N_2350,N_2302);
nand U2790 (N_2790,N_2285,N_2284);
or U2791 (N_2791,N_2320,N_2215);
and U2792 (N_2792,N_2145,N_2105);
xor U2793 (N_2793,N_2193,N_2127);
and U2794 (N_2794,N_2305,N_2100);
and U2795 (N_2795,N_2244,N_2342);
nand U2796 (N_2796,N_2393,N_2124);
nor U2797 (N_2797,N_1896,N_2063);
or U2798 (N_2798,N_1963,N_2224);
and U2799 (N_2799,N_1945,N_1869);
and U2800 (N_2800,N_2229,N_1929);
nand U2801 (N_2801,N_2087,N_2274);
nand U2802 (N_2802,N_1911,N_2388);
nand U2803 (N_2803,N_1959,N_1895);
or U2804 (N_2804,N_1913,N_1835);
nor U2805 (N_2805,N_1992,N_2219);
nand U2806 (N_2806,N_1907,N_1855);
and U2807 (N_2807,N_2210,N_2220);
and U2808 (N_2808,N_1841,N_2389);
nand U2809 (N_2809,N_1957,N_2000);
and U2810 (N_2810,N_1819,N_1990);
nand U2811 (N_2811,N_2100,N_1954);
and U2812 (N_2812,N_2048,N_2007);
and U2813 (N_2813,N_2322,N_2053);
or U2814 (N_2814,N_1962,N_1922);
nand U2815 (N_2815,N_2330,N_2005);
or U2816 (N_2816,N_2115,N_2015);
nor U2817 (N_2817,N_1883,N_2106);
nand U2818 (N_2818,N_1891,N_2088);
xnor U2819 (N_2819,N_1871,N_2270);
nor U2820 (N_2820,N_1857,N_2170);
and U2821 (N_2821,N_2114,N_1836);
and U2822 (N_2822,N_2223,N_2208);
xnor U2823 (N_2823,N_1820,N_1923);
nand U2824 (N_2824,N_2188,N_2354);
nor U2825 (N_2825,N_2273,N_2377);
nand U2826 (N_2826,N_2079,N_1954);
nor U2827 (N_2827,N_2305,N_2293);
nor U2828 (N_2828,N_1977,N_2180);
nand U2829 (N_2829,N_2138,N_2256);
nor U2830 (N_2830,N_2055,N_1983);
nor U2831 (N_2831,N_2155,N_2379);
nor U2832 (N_2832,N_2222,N_1892);
and U2833 (N_2833,N_1959,N_2350);
and U2834 (N_2834,N_1836,N_2054);
and U2835 (N_2835,N_2051,N_2188);
nand U2836 (N_2836,N_1961,N_1898);
or U2837 (N_2837,N_1883,N_2080);
xor U2838 (N_2838,N_1823,N_1872);
or U2839 (N_2839,N_2269,N_2090);
and U2840 (N_2840,N_1921,N_2075);
nand U2841 (N_2841,N_2259,N_1812);
and U2842 (N_2842,N_1929,N_2292);
and U2843 (N_2843,N_2296,N_2306);
or U2844 (N_2844,N_1980,N_2345);
or U2845 (N_2845,N_2172,N_2130);
nor U2846 (N_2846,N_1948,N_2351);
nand U2847 (N_2847,N_2399,N_2257);
nor U2848 (N_2848,N_2350,N_2368);
nor U2849 (N_2849,N_1931,N_1835);
xor U2850 (N_2850,N_1816,N_2365);
or U2851 (N_2851,N_2105,N_2238);
and U2852 (N_2852,N_1896,N_1867);
and U2853 (N_2853,N_2263,N_2381);
xnor U2854 (N_2854,N_2274,N_2090);
nor U2855 (N_2855,N_1823,N_1849);
nor U2856 (N_2856,N_2370,N_1925);
nand U2857 (N_2857,N_2110,N_2268);
nand U2858 (N_2858,N_1886,N_2259);
nand U2859 (N_2859,N_1896,N_2273);
nor U2860 (N_2860,N_1850,N_2095);
nor U2861 (N_2861,N_1823,N_2088);
nor U2862 (N_2862,N_1801,N_2067);
and U2863 (N_2863,N_2268,N_2069);
or U2864 (N_2864,N_2343,N_2061);
or U2865 (N_2865,N_1917,N_1978);
xnor U2866 (N_2866,N_1879,N_1995);
and U2867 (N_2867,N_2002,N_2299);
and U2868 (N_2868,N_2020,N_1927);
and U2869 (N_2869,N_2122,N_2132);
and U2870 (N_2870,N_2338,N_2242);
nor U2871 (N_2871,N_1937,N_1877);
xor U2872 (N_2872,N_2223,N_2064);
and U2873 (N_2873,N_2319,N_2084);
nor U2874 (N_2874,N_2276,N_1919);
xnor U2875 (N_2875,N_2025,N_2039);
or U2876 (N_2876,N_1811,N_1954);
and U2877 (N_2877,N_1984,N_1956);
nand U2878 (N_2878,N_2277,N_2332);
or U2879 (N_2879,N_2147,N_1827);
or U2880 (N_2880,N_2250,N_2318);
or U2881 (N_2881,N_1809,N_2008);
nand U2882 (N_2882,N_2224,N_2005);
nor U2883 (N_2883,N_2262,N_2289);
nor U2884 (N_2884,N_2236,N_2163);
nand U2885 (N_2885,N_2082,N_2185);
or U2886 (N_2886,N_1986,N_2399);
and U2887 (N_2887,N_2009,N_2197);
xor U2888 (N_2888,N_2134,N_2147);
nand U2889 (N_2889,N_2255,N_1878);
nand U2890 (N_2890,N_2287,N_1895);
or U2891 (N_2891,N_2323,N_2181);
nor U2892 (N_2892,N_2078,N_1942);
nand U2893 (N_2893,N_2085,N_2134);
nor U2894 (N_2894,N_2267,N_2169);
nand U2895 (N_2895,N_2073,N_2252);
or U2896 (N_2896,N_2242,N_2020);
xnor U2897 (N_2897,N_1852,N_2087);
and U2898 (N_2898,N_2121,N_1860);
nor U2899 (N_2899,N_2347,N_1823);
or U2900 (N_2900,N_2218,N_1856);
and U2901 (N_2901,N_2042,N_2257);
nand U2902 (N_2902,N_2261,N_1950);
and U2903 (N_2903,N_1948,N_2128);
xnor U2904 (N_2904,N_1987,N_2360);
and U2905 (N_2905,N_2220,N_2035);
and U2906 (N_2906,N_2336,N_2013);
nor U2907 (N_2907,N_2345,N_1879);
and U2908 (N_2908,N_2317,N_2294);
and U2909 (N_2909,N_1872,N_2205);
nand U2910 (N_2910,N_2384,N_2250);
nor U2911 (N_2911,N_2072,N_2231);
nor U2912 (N_2912,N_1983,N_2063);
nor U2913 (N_2913,N_2168,N_2367);
xnor U2914 (N_2914,N_2372,N_1873);
nand U2915 (N_2915,N_2338,N_1950);
or U2916 (N_2916,N_1911,N_2326);
or U2917 (N_2917,N_2150,N_2099);
nand U2918 (N_2918,N_2189,N_1919);
or U2919 (N_2919,N_2013,N_2334);
or U2920 (N_2920,N_1850,N_2325);
and U2921 (N_2921,N_2303,N_1980);
nand U2922 (N_2922,N_2147,N_2108);
xor U2923 (N_2923,N_2085,N_1908);
xnor U2924 (N_2924,N_2183,N_2067);
or U2925 (N_2925,N_2329,N_2106);
or U2926 (N_2926,N_1966,N_2358);
and U2927 (N_2927,N_1932,N_2339);
xor U2928 (N_2928,N_1969,N_2012);
or U2929 (N_2929,N_2313,N_2108);
nand U2930 (N_2930,N_2366,N_1983);
nand U2931 (N_2931,N_1869,N_2318);
or U2932 (N_2932,N_1873,N_2296);
nand U2933 (N_2933,N_1880,N_2071);
nor U2934 (N_2934,N_2162,N_2264);
nand U2935 (N_2935,N_2019,N_2223);
nand U2936 (N_2936,N_2243,N_1943);
nor U2937 (N_2937,N_2270,N_2250);
xnor U2938 (N_2938,N_1902,N_2185);
nor U2939 (N_2939,N_2367,N_1823);
nand U2940 (N_2940,N_2111,N_2384);
or U2941 (N_2941,N_2303,N_2176);
and U2942 (N_2942,N_2193,N_1861);
nor U2943 (N_2943,N_1813,N_2119);
xnor U2944 (N_2944,N_1960,N_2309);
nand U2945 (N_2945,N_2159,N_2021);
nand U2946 (N_2946,N_1842,N_2297);
or U2947 (N_2947,N_2057,N_2302);
nor U2948 (N_2948,N_2090,N_1834);
nand U2949 (N_2949,N_2287,N_2079);
and U2950 (N_2950,N_1860,N_2208);
and U2951 (N_2951,N_2089,N_2275);
and U2952 (N_2952,N_2294,N_2019);
and U2953 (N_2953,N_2159,N_2177);
nand U2954 (N_2954,N_2042,N_1967);
nor U2955 (N_2955,N_1928,N_1920);
nand U2956 (N_2956,N_2168,N_1877);
nor U2957 (N_2957,N_2388,N_2190);
nor U2958 (N_2958,N_1949,N_2098);
nor U2959 (N_2959,N_2394,N_1991);
or U2960 (N_2960,N_2206,N_2236);
and U2961 (N_2961,N_2380,N_2150);
nand U2962 (N_2962,N_1826,N_2070);
nor U2963 (N_2963,N_1842,N_1945);
nand U2964 (N_2964,N_1979,N_2107);
xnor U2965 (N_2965,N_1957,N_2332);
or U2966 (N_2966,N_2062,N_2049);
nor U2967 (N_2967,N_2302,N_1955);
or U2968 (N_2968,N_2284,N_1956);
nor U2969 (N_2969,N_2278,N_2033);
xnor U2970 (N_2970,N_1881,N_2330);
nor U2971 (N_2971,N_2117,N_1916);
or U2972 (N_2972,N_2193,N_1857);
nand U2973 (N_2973,N_1819,N_2208);
and U2974 (N_2974,N_2307,N_1905);
and U2975 (N_2975,N_2346,N_2038);
nand U2976 (N_2976,N_2197,N_1932);
nand U2977 (N_2977,N_2104,N_2072);
nand U2978 (N_2978,N_2393,N_2107);
xnor U2979 (N_2979,N_2246,N_1931);
or U2980 (N_2980,N_2051,N_2019);
xor U2981 (N_2981,N_2224,N_1878);
or U2982 (N_2982,N_1829,N_1915);
and U2983 (N_2983,N_2177,N_2190);
or U2984 (N_2984,N_1867,N_1837);
nand U2985 (N_2985,N_1875,N_2351);
nand U2986 (N_2986,N_1838,N_2388);
nor U2987 (N_2987,N_2265,N_1964);
nor U2988 (N_2988,N_2270,N_2135);
nor U2989 (N_2989,N_1919,N_1997);
nor U2990 (N_2990,N_2312,N_2374);
nand U2991 (N_2991,N_1945,N_2146);
or U2992 (N_2992,N_2027,N_1881);
and U2993 (N_2993,N_1974,N_1817);
nor U2994 (N_2994,N_2086,N_1804);
and U2995 (N_2995,N_2080,N_2073);
xnor U2996 (N_2996,N_2182,N_2033);
nor U2997 (N_2997,N_2258,N_2274);
nor U2998 (N_2998,N_2113,N_2096);
nor U2999 (N_2999,N_2336,N_1929);
nor UO_0 (O_0,N_2998,N_2506);
and UO_1 (O_1,N_2966,N_2935);
and UO_2 (O_2,N_2950,N_2980);
and UO_3 (O_3,N_2789,N_2892);
nand UO_4 (O_4,N_2835,N_2515);
nand UO_5 (O_5,N_2478,N_2837);
nand UO_6 (O_6,N_2903,N_2987);
and UO_7 (O_7,N_2725,N_2617);
and UO_8 (O_8,N_2636,N_2413);
nor UO_9 (O_9,N_2816,N_2425);
or UO_10 (O_10,N_2610,N_2676);
and UO_11 (O_11,N_2955,N_2439);
or UO_12 (O_12,N_2827,N_2778);
and UO_13 (O_13,N_2702,N_2943);
nand UO_14 (O_14,N_2990,N_2929);
or UO_15 (O_15,N_2989,N_2868);
or UO_16 (O_16,N_2641,N_2458);
nor UO_17 (O_17,N_2490,N_2573);
nor UO_18 (O_18,N_2491,N_2708);
nor UO_19 (O_19,N_2700,N_2684);
nand UO_20 (O_20,N_2919,N_2651);
nand UO_21 (O_21,N_2792,N_2685);
and UO_22 (O_22,N_2514,N_2918);
nand UO_23 (O_23,N_2802,N_2488);
nand UO_24 (O_24,N_2462,N_2507);
or UO_25 (O_25,N_2806,N_2587);
xnor UO_26 (O_26,N_2819,N_2597);
or UO_27 (O_27,N_2628,N_2734);
or UO_28 (O_28,N_2770,N_2787);
xor UO_29 (O_29,N_2487,N_2479);
nand UO_30 (O_30,N_2862,N_2761);
or UO_31 (O_31,N_2404,N_2416);
and UO_32 (O_32,N_2591,N_2659);
or UO_33 (O_33,N_2414,N_2695);
nor UO_34 (O_34,N_2775,N_2904);
and UO_35 (O_35,N_2600,N_2483);
and UO_36 (O_36,N_2876,N_2596);
nor UO_37 (O_37,N_2944,N_2457);
and UO_38 (O_38,N_2469,N_2453);
and UO_39 (O_39,N_2531,N_2959);
nor UO_40 (O_40,N_2759,N_2530);
nand UO_41 (O_41,N_2973,N_2732);
nor UO_42 (O_42,N_2454,N_2549);
and UO_43 (O_43,N_2570,N_2670);
nand UO_44 (O_44,N_2664,N_2901);
and UO_45 (O_45,N_2804,N_2814);
and UO_46 (O_46,N_2577,N_2902);
or UO_47 (O_47,N_2466,N_2758);
and UO_48 (O_48,N_2590,N_2602);
or UO_49 (O_49,N_2565,N_2409);
or UO_50 (O_50,N_2848,N_2823);
nand UO_51 (O_51,N_2748,N_2884);
and UO_52 (O_52,N_2535,N_2444);
nor UO_53 (O_53,N_2697,N_2542);
or UO_54 (O_54,N_2709,N_2555);
nand UO_55 (O_55,N_2571,N_2782);
and UO_56 (O_56,N_2502,N_2923);
nand UO_57 (O_57,N_2633,N_2605);
nor UO_58 (O_58,N_2927,N_2908);
nor UO_59 (O_59,N_2871,N_2406);
nand UO_60 (O_60,N_2694,N_2964);
and UO_61 (O_61,N_2441,N_2500);
and UO_62 (O_62,N_2821,N_2863);
or UO_63 (O_63,N_2951,N_2470);
or UO_64 (O_64,N_2681,N_2768);
nor UO_65 (O_65,N_2726,N_2933);
and UO_66 (O_66,N_2949,N_2473);
nand UO_67 (O_67,N_2877,N_2411);
and UO_68 (O_68,N_2632,N_2859);
or UO_69 (O_69,N_2760,N_2757);
nand UO_70 (O_70,N_2885,N_2494);
nand UO_71 (O_71,N_2723,N_2997);
nor UO_72 (O_72,N_2781,N_2522);
or UO_73 (O_73,N_2442,N_2996);
and UO_74 (O_74,N_2679,N_2840);
nor UO_75 (O_75,N_2643,N_2941);
nor UO_76 (O_76,N_2896,N_2578);
or UO_77 (O_77,N_2607,N_2742);
nor UO_78 (O_78,N_2655,N_2661);
or UO_79 (O_79,N_2958,N_2574);
and UO_80 (O_80,N_2735,N_2909);
and UO_81 (O_81,N_2402,N_2471);
and UO_82 (O_82,N_2803,N_2970);
or UO_83 (O_83,N_2558,N_2796);
and UO_84 (O_84,N_2900,N_2513);
or UO_85 (O_85,N_2992,N_2660);
nor UO_86 (O_86,N_2677,N_2603);
nand UO_87 (O_87,N_2833,N_2427);
xor UO_88 (O_88,N_2930,N_2562);
or UO_89 (O_89,N_2707,N_2865);
and UO_90 (O_90,N_2485,N_2747);
nor UO_91 (O_91,N_2773,N_2690);
nor UO_92 (O_92,N_2831,N_2945);
or UO_93 (O_93,N_2873,N_2777);
nor UO_94 (O_94,N_2477,N_2808);
nor UO_95 (O_95,N_2650,N_2851);
or UO_96 (O_96,N_2874,N_2417);
nand UO_97 (O_97,N_2649,N_2640);
or UO_98 (O_98,N_2813,N_2995);
or UO_99 (O_99,N_2853,N_2489);
or UO_100 (O_100,N_2625,N_2893);
nand UO_101 (O_101,N_2436,N_2476);
and UO_102 (O_102,N_2560,N_2461);
and UO_103 (O_103,N_2754,N_2432);
nand UO_104 (O_104,N_2746,N_2745);
or UO_105 (O_105,N_2619,N_2741);
or UO_106 (O_106,N_2701,N_2645);
xnor UO_107 (O_107,N_2484,N_2663);
nand UO_108 (O_108,N_2727,N_2783);
nand UO_109 (O_109,N_2481,N_2836);
or UO_110 (O_110,N_2912,N_2569);
or UO_111 (O_111,N_2637,N_2815);
nand UO_112 (O_112,N_2940,N_2850);
nand UO_113 (O_113,N_2852,N_2431);
nand UO_114 (O_114,N_2673,N_2898);
or UO_115 (O_115,N_2456,N_2843);
nor UO_116 (O_116,N_2631,N_2857);
and UO_117 (O_117,N_2869,N_2811);
or UO_118 (O_118,N_2426,N_2653);
or UO_119 (O_119,N_2960,N_2765);
nand UO_120 (O_120,N_2686,N_2671);
and UO_121 (O_121,N_2864,N_2991);
nand UO_122 (O_122,N_2860,N_2794);
or UO_123 (O_123,N_2688,N_2572);
or UO_124 (O_124,N_2526,N_2675);
or UO_125 (O_125,N_2799,N_2693);
nor UO_126 (O_126,N_2914,N_2744);
nand UO_127 (O_127,N_2638,N_2496);
or UO_128 (O_128,N_2825,N_2972);
nor UO_129 (O_129,N_2762,N_2986);
nor UO_130 (O_130,N_2451,N_2826);
or UO_131 (O_131,N_2769,N_2482);
and UO_132 (O_132,N_2652,N_2517);
or UO_133 (O_133,N_2599,N_2418);
or UO_134 (O_134,N_2962,N_2508);
nor UO_135 (O_135,N_2752,N_2920);
or UO_136 (O_136,N_2849,N_2561);
or UO_137 (O_137,N_2438,N_2576);
xor UO_138 (O_138,N_2475,N_2820);
or UO_139 (O_139,N_2785,N_2447);
and UO_140 (O_140,N_2516,N_2635);
xor UO_141 (O_141,N_2875,N_2527);
and UO_142 (O_142,N_2545,N_2861);
and UO_143 (O_143,N_2780,N_2810);
and UO_144 (O_144,N_2407,N_2548);
or UO_145 (O_145,N_2435,N_2498);
xor UO_146 (O_146,N_2419,N_2867);
nor UO_147 (O_147,N_2907,N_2595);
nor UO_148 (O_148,N_2937,N_2905);
nor UO_149 (O_149,N_2412,N_2683);
and UO_150 (O_150,N_2764,N_2698);
xnor UO_151 (O_151,N_2598,N_2422);
nor UO_152 (O_152,N_2800,N_2467);
xnor UO_153 (O_153,N_2585,N_2609);
xor UO_154 (O_154,N_2566,N_2528);
and UO_155 (O_155,N_2616,N_2968);
and UO_156 (O_156,N_2629,N_2620);
nand UO_157 (O_157,N_2644,N_2739);
nor UO_158 (O_158,N_2805,N_2834);
and UO_159 (O_159,N_2621,N_2463);
nand UO_160 (O_160,N_2556,N_2975);
nor UO_161 (O_161,N_2532,N_2983);
xor UO_162 (O_162,N_2772,N_2845);
nand UO_163 (O_163,N_2984,N_2518);
nor UO_164 (O_164,N_2771,N_2541);
and UO_165 (O_165,N_2446,N_2779);
nand UO_166 (O_166,N_2720,N_2428);
nor UO_167 (O_167,N_2961,N_2567);
nand UO_168 (O_168,N_2776,N_2705);
nand UO_169 (O_169,N_2689,N_2824);
nand UO_170 (O_170,N_2622,N_2988);
nand UO_171 (O_171,N_2812,N_2881);
nor UO_172 (O_172,N_2890,N_2536);
xor UO_173 (O_173,N_2459,N_2588);
or UO_174 (O_174,N_2963,N_2706);
and UO_175 (O_175,N_2829,N_2408);
nand UO_176 (O_176,N_2978,N_2550);
nand UO_177 (O_177,N_2430,N_2818);
or UO_178 (O_178,N_2703,N_2575);
or UO_179 (O_179,N_2928,N_2994);
and UO_180 (O_180,N_2713,N_2552);
nand UO_181 (O_181,N_2795,N_2627);
nor UO_182 (O_182,N_2910,N_2895);
nand UO_183 (O_183,N_2691,N_2942);
xor UO_184 (O_184,N_2533,N_2505);
and UO_185 (O_185,N_2583,N_2630);
nand UO_186 (O_186,N_2433,N_2809);
nand UO_187 (O_187,N_2537,N_2916);
nor UO_188 (O_188,N_2547,N_2969);
xnor UO_189 (O_189,N_2887,N_2455);
or UO_190 (O_190,N_2582,N_2736);
or UO_191 (O_191,N_2728,N_2844);
and UO_192 (O_192,N_2967,N_2906);
nor UO_193 (O_193,N_2985,N_2733);
xor UO_194 (O_194,N_2715,N_2584);
or UO_195 (O_195,N_2618,N_2883);
nand UO_196 (O_196,N_2880,N_2965);
nand UO_197 (O_197,N_2801,N_2750);
and UO_198 (O_198,N_2519,N_2842);
or UO_199 (O_199,N_2790,N_2423);
nor UO_200 (O_200,N_2564,N_2817);
or UO_201 (O_201,N_2434,N_2559);
nor UO_202 (O_202,N_2993,N_2642);
nand UO_203 (O_203,N_2711,N_2882);
nor UO_204 (O_204,N_2678,N_2626);
or UO_205 (O_205,N_2553,N_2510);
or UO_206 (O_206,N_2464,N_2538);
xnor UO_207 (O_207,N_2554,N_2606);
and UO_208 (O_208,N_2639,N_2403);
nor UO_209 (O_209,N_2656,N_2911);
or UO_210 (O_210,N_2551,N_2947);
nand UO_211 (O_211,N_2534,N_2791);
or UO_212 (O_212,N_2957,N_2738);
and UO_213 (O_213,N_2400,N_2615);
nand UO_214 (O_214,N_2717,N_2449);
or UO_215 (O_215,N_2926,N_2604);
xnor UO_216 (O_216,N_2543,N_2841);
nor UO_217 (O_217,N_2523,N_2756);
nand UO_218 (O_218,N_2592,N_2593);
and UO_219 (O_219,N_2828,N_2493);
or UO_220 (O_220,N_2657,N_2539);
or UO_221 (O_221,N_2546,N_2586);
xor UO_222 (O_222,N_2511,N_2714);
nor UO_223 (O_223,N_2886,N_2529);
nand UO_224 (O_224,N_2499,N_2797);
nand UO_225 (O_225,N_2913,N_2401);
or UO_226 (O_226,N_2646,N_2982);
and UO_227 (O_227,N_2594,N_2421);
or UO_228 (O_228,N_2563,N_2872);
or UO_229 (O_229,N_2938,N_2767);
nand UO_230 (O_230,N_2956,N_2870);
and UO_231 (O_231,N_2856,N_2682);
and UO_232 (O_232,N_2953,N_2710);
nor UO_233 (O_233,N_2647,N_2699);
nand UO_234 (O_234,N_2915,N_2472);
or UO_235 (O_235,N_2525,N_2753);
nand UO_236 (O_236,N_2634,N_2474);
nand UO_237 (O_237,N_2974,N_2612);
and UO_238 (O_238,N_2722,N_2879);
nand UO_239 (O_239,N_2492,N_2729);
nand UO_240 (O_240,N_2925,N_2579);
and UO_241 (O_241,N_2838,N_2888);
and UO_242 (O_242,N_2924,N_2503);
or UO_243 (O_243,N_2737,N_2666);
and UO_244 (O_244,N_2763,N_2922);
or UO_245 (O_245,N_2774,N_2410);
nor UO_246 (O_246,N_2465,N_2665);
and UO_247 (O_247,N_2495,N_2999);
or UO_248 (O_248,N_2669,N_2452);
xor UO_249 (O_249,N_2509,N_2524);
or UO_250 (O_250,N_2755,N_2624);
or UO_251 (O_251,N_2846,N_2654);
nand UO_252 (O_252,N_2878,N_2601);
nand UO_253 (O_253,N_2784,N_2497);
nor UO_254 (O_254,N_2889,N_2981);
nor UO_255 (O_255,N_2855,N_2934);
or UO_256 (O_256,N_2420,N_2952);
xor UO_257 (O_257,N_2830,N_2948);
or UO_258 (O_258,N_2674,N_2847);
and UO_259 (O_259,N_2460,N_2501);
nor UO_260 (O_260,N_2445,N_2512);
nor UO_261 (O_261,N_2662,N_2415);
nor UO_262 (O_262,N_2897,N_2839);
and UO_263 (O_263,N_2540,N_2971);
nand UO_264 (O_264,N_2504,N_2623);
nand UO_265 (O_265,N_2719,N_2658);
and UO_266 (O_266,N_2917,N_2440);
and UO_267 (O_267,N_2740,N_2946);
or UO_268 (O_268,N_2749,N_2979);
xor UO_269 (O_269,N_2648,N_2680);
and UO_270 (O_270,N_2832,N_2932);
or UO_271 (O_271,N_2931,N_2443);
and UO_272 (O_272,N_2611,N_2589);
nor UO_273 (O_273,N_2891,N_2712);
nor UO_274 (O_274,N_2480,N_2613);
and UO_275 (O_275,N_2608,N_2894);
nand UO_276 (O_276,N_2486,N_2822);
and UO_277 (O_277,N_2450,N_2696);
xor UO_278 (O_278,N_2793,N_2672);
nand UO_279 (O_279,N_2766,N_2448);
and UO_280 (O_280,N_2521,N_2798);
nor UO_281 (O_281,N_2954,N_2405);
nor UO_282 (O_282,N_2786,N_2568);
nor UO_283 (O_283,N_2544,N_2704);
xor UO_284 (O_284,N_2580,N_2807);
and UO_285 (O_285,N_2718,N_2520);
xor UO_286 (O_286,N_2751,N_2424);
nor UO_287 (O_287,N_2437,N_2788);
or UO_288 (O_288,N_2668,N_2429);
nor UO_289 (O_289,N_2976,N_2921);
nand UO_290 (O_290,N_2716,N_2468);
or UO_291 (O_291,N_2866,N_2667);
and UO_292 (O_292,N_2692,N_2858);
and UO_293 (O_293,N_2557,N_2936);
xnor UO_294 (O_294,N_2730,N_2854);
nand UO_295 (O_295,N_2581,N_2899);
nand UO_296 (O_296,N_2721,N_2743);
nand UO_297 (O_297,N_2724,N_2614);
xnor UO_298 (O_298,N_2731,N_2977);
xnor UO_299 (O_299,N_2687,N_2939);
nor UO_300 (O_300,N_2602,N_2596);
and UO_301 (O_301,N_2668,N_2416);
or UO_302 (O_302,N_2509,N_2501);
and UO_303 (O_303,N_2744,N_2983);
nor UO_304 (O_304,N_2607,N_2674);
nor UO_305 (O_305,N_2885,N_2468);
or UO_306 (O_306,N_2636,N_2619);
nor UO_307 (O_307,N_2630,N_2909);
nor UO_308 (O_308,N_2762,N_2529);
and UO_309 (O_309,N_2657,N_2438);
or UO_310 (O_310,N_2901,N_2725);
and UO_311 (O_311,N_2446,N_2999);
xnor UO_312 (O_312,N_2602,N_2433);
and UO_313 (O_313,N_2737,N_2975);
and UO_314 (O_314,N_2938,N_2576);
nand UO_315 (O_315,N_2609,N_2711);
or UO_316 (O_316,N_2554,N_2706);
nand UO_317 (O_317,N_2838,N_2778);
xor UO_318 (O_318,N_2561,N_2602);
or UO_319 (O_319,N_2670,N_2900);
or UO_320 (O_320,N_2894,N_2998);
nor UO_321 (O_321,N_2919,N_2769);
nand UO_322 (O_322,N_2858,N_2868);
or UO_323 (O_323,N_2801,N_2571);
nor UO_324 (O_324,N_2542,N_2600);
xnor UO_325 (O_325,N_2764,N_2595);
nor UO_326 (O_326,N_2554,N_2544);
and UO_327 (O_327,N_2963,N_2642);
xnor UO_328 (O_328,N_2536,N_2765);
nor UO_329 (O_329,N_2899,N_2435);
and UO_330 (O_330,N_2747,N_2801);
or UO_331 (O_331,N_2988,N_2493);
xnor UO_332 (O_332,N_2797,N_2785);
nand UO_333 (O_333,N_2764,N_2868);
nand UO_334 (O_334,N_2560,N_2591);
or UO_335 (O_335,N_2437,N_2460);
xnor UO_336 (O_336,N_2523,N_2690);
nor UO_337 (O_337,N_2968,N_2447);
xnor UO_338 (O_338,N_2702,N_2874);
or UO_339 (O_339,N_2845,N_2551);
nor UO_340 (O_340,N_2550,N_2458);
or UO_341 (O_341,N_2560,N_2990);
and UO_342 (O_342,N_2457,N_2534);
and UO_343 (O_343,N_2555,N_2602);
nand UO_344 (O_344,N_2687,N_2552);
and UO_345 (O_345,N_2826,N_2613);
nor UO_346 (O_346,N_2423,N_2987);
nor UO_347 (O_347,N_2515,N_2546);
and UO_348 (O_348,N_2482,N_2515);
nand UO_349 (O_349,N_2741,N_2596);
and UO_350 (O_350,N_2760,N_2562);
nor UO_351 (O_351,N_2916,N_2734);
or UO_352 (O_352,N_2627,N_2519);
and UO_353 (O_353,N_2913,N_2816);
or UO_354 (O_354,N_2821,N_2635);
and UO_355 (O_355,N_2741,N_2534);
nor UO_356 (O_356,N_2428,N_2989);
nor UO_357 (O_357,N_2501,N_2494);
or UO_358 (O_358,N_2916,N_2769);
nor UO_359 (O_359,N_2877,N_2980);
or UO_360 (O_360,N_2607,N_2829);
and UO_361 (O_361,N_2763,N_2472);
nand UO_362 (O_362,N_2625,N_2985);
and UO_363 (O_363,N_2786,N_2751);
nand UO_364 (O_364,N_2912,N_2935);
nand UO_365 (O_365,N_2480,N_2490);
or UO_366 (O_366,N_2532,N_2674);
nor UO_367 (O_367,N_2597,N_2583);
or UO_368 (O_368,N_2692,N_2659);
xnor UO_369 (O_369,N_2475,N_2600);
or UO_370 (O_370,N_2468,N_2609);
xnor UO_371 (O_371,N_2890,N_2507);
or UO_372 (O_372,N_2499,N_2798);
xor UO_373 (O_373,N_2758,N_2861);
or UO_374 (O_374,N_2496,N_2462);
nand UO_375 (O_375,N_2533,N_2772);
nor UO_376 (O_376,N_2488,N_2999);
or UO_377 (O_377,N_2923,N_2868);
or UO_378 (O_378,N_2838,N_2723);
and UO_379 (O_379,N_2718,N_2647);
nor UO_380 (O_380,N_2945,N_2713);
and UO_381 (O_381,N_2945,N_2467);
nor UO_382 (O_382,N_2642,N_2578);
nand UO_383 (O_383,N_2593,N_2925);
or UO_384 (O_384,N_2983,N_2401);
nand UO_385 (O_385,N_2914,N_2668);
nand UO_386 (O_386,N_2451,N_2900);
or UO_387 (O_387,N_2460,N_2489);
or UO_388 (O_388,N_2452,N_2668);
or UO_389 (O_389,N_2440,N_2827);
or UO_390 (O_390,N_2474,N_2556);
nor UO_391 (O_391,N_2702,N_2670);
nor UO_392 (O_392,N_2666,N_2777);
nor UO_393 (O_393,N_2748,N_2834);
and UO_394 (O_394,N_2735,N_2730);
nand UO_395 (O_395,N_2426,N_2517);
nor UO_396 (O_396,N_2496,N_2435);
nand UO_397 (O_397,N_2971,N_2976);
nand UO_398 (O_398,N_2494,N_2778);
nor UO_399 (O_399,N_2776,N_2657);
nand UO_400 (O_400,N_2820,N_2549);
and UO_401 (O_401,N_2739,N_2688);
nand UO_402 (O_402,N_2550,N_2575);
nor UO_403 (O_403,N_2519,N_2871);
or UO_404 (O_404,N_2404,N_2562);
and UO_405 (O_405,N_2596,N_2787);
nor UO_406 (O_406,N_2703,N_2955);
nor UO_407 (O_407,N_2557,N_2413);
xor UO_408 (O_408,N_2731,N_2559);
nor UO_409 (O_409,N_2941,N_2851);
or UO_410 (O_410,N_2892,N_2546);
or UO_411 (O_411,N_2554,N_2563);
or UO_412 (O_412,N_2613,N_2511);
and UO_413 (O_413,N_2763,N_2424);
or UO_414 (O_414,N_2435,N_2542);
and UO_415 (O_415,N_2950,N_2840);
nand UO_416 (O_416,N_2883,N_2945);
xnor UO_417 (O_417,N_2568,N_2541);
nand UO_418 (O_418,N_2716,N_2599);
xnor UO_419 (O_419,N_2836,N_2803);
xor UO_420 (O_420,N_2862,N_2815);
nor UO_421 (O_421,N_2806,N_2762);
or UO_422 (O_422,N_2607,N_2544);
nor UO_423 (O_423,N_2991,N_2682);
xor UO_424 (O_424,N_2726,N_2850);
nand UO_425 (O_425,N_2752,N_2839);
nand UO_426 (O_426,N_2711,N_2972);
xnor UO_427 (O_427,N_2723,N_2649);
or UO_428 (O_428,N_2613,N_2667);
nor UO_429 (O_429,N_2612,N_2481);
or UO_430 (O_430,N_2839,N_2435);
nand UO_431 (O_431,N_2917,N_2435);
or UO_432 (O_432,N_2982,N_2539);
or UO_433 (O_433,N_2719,N_2889);
or UO_434 (O_434,N_2594,N_2811);
nor UO_435 (O_435,N_2420,N_2868);
nor UO_436 (O_436,N_2642,N_2529);
nor UO_437 (O_437,N_2447,N_2591);
xnor UO_438 (O_438,N_2908,N_2809);
and UO_439 (O_439,N_2718,N_2427);
xor UO_440 (O_440,N_2716,N_2917);
nand UO_441 (O_441,N_2661,N_2700);
and UO_442 (O_442,N_2987,N_2947);
and UO_443 (O_443,N_2964,N_2697);
nand UO_444 (O_444,N_2689,N_2671);
or UO_445 (O_445,N_2965,N_2836);
or UO_446 (O_446,N_2806,N_2630);
or UO_447 (O_447,N_2911,N_2921);
nand UO_448 (O_448,N_2833,N_2462);
nand UO_449 (O_449,N_2847,N_2999);
or UO_450 (O_450,N_2948,N_2912);
nand UO_451 (O_451,N_2557,N_2929);
or UO_452 (O_452,N_2657,N_2951);
nand UO_453 (O_453,N_2805,N_2868);
or UO_454 (O_454,N_2660,N_2738);
and UO_455 (O_455,N_2717,N_2485);
or UO_456 (O_456,N_2462,N_2941);
nor UO_457 (O_457,N_2798,N_2737);
and UO_458 (O_458,N_2620,N_2723);
nand UO_459 (O_459,N_2924,N_2812);
nor UO_460 (O_460,N_2859,N_2548);
or UO_461 (O_461,N_2865,N_2630);
nand UO_462 (O_462,N_2502,N_2405);
nand UO_463 (O_463,N_2896,N_2412);
xor UO_464 (O_464,N_2814,N_2401);
nand UO_465 (O_465,N_2572,N_2567);
and UO_466 (O_466,N_2762,N_2557);
nand UO_467 (O_467,N_2771,N_2721);
and UO_468 (O_468,N_2414,N_2762);
nand UO_469 (O_469,N_2607,N_2467);
nor UO_470 (O_470,N_2738,N_2665);
nor UO_471 (O_471,N_2721,N_2739);
or UO_472 (O_472,N_2867,N_2443);
nor UO_473 (O_473,N_2741,N_2895);
and UO_474 (O_474,N_2762,N_2663);
nor UO_475 (O_475,N_2529,N_2941);
and UO_476 (O_476,N_2566,N_2526);
and UO_477 (O_477,N_2876,N_2556);
nor UO_478 (O_478,N_2914,N_2946);
nand UO_479 (O_479,N_2588,N_2734);
and UO_480 (O_480,N_2995,N_2414);
or UO_481 (O_481,N_2460,N_2687);
xnor UO_482 (O_482,N_2445,N_2689);
or UO_483 (O_483,N_2652,N_2543);
nor UO_484 (O_484,N_2677,N_2703);
xnor UO_485 (O_485,N_2506,N_2896);
and UO_486 (O_486,N_2644,N_2670);
nand UO_487 (O_487,N_2612,N_2541);
and UO_488 (O_488,N_2676,N_2784);
or UO_489 (O_489,N_2830,N_2856);
nand UO_490 (O_490,N_2999,N_2485);
or UO_491 (O_491,N_2607,N_2478);
or UO_492 (O_492,N_2824,N_2835);
and UO_493 (O_493,N_2830,N_2426);
nand UO_494 (O_494,N_2932,N_2509);
nand UO_495 (O_495,N_2450,N_2876);
or UO_496 (O_496,N_2509,N_2953);
and UO_497 (O_497,N_2741,N_2716);
or UO_498 (O_498,N_2879,N_2891);
nand UO_499 (O_499,N_2484,N_2835);
endmodule