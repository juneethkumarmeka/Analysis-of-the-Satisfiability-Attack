module basic_2000_20000_2500_20_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
and U0 (N_0,In_161,In_671);
and U1 (N_1,In_1127,In_1815);
xor U2 (N_2,In_634,In_1787);
nor U3 (N_3,In_1056,In_1289);
or U4 (N_4,In_1975,In_1008);
or U5 (N_5,In_1088,In_1508);
or U6 (N_6,In_1187,In_29);
nor U7 (N_7,In_1919,In_82);
xnor U8 (N_8,In_1827,In_1599);
nor U9 (N_9,In_22,In_750);
xnor U10 (N_10,In_227,In_1565);
nand U11 (N_11,In_987,In_1171);
or U12 (N_12,In_373,In_1943);
and U13 (N_13,In_225,In_399);
or U14 (N_14,In_997,In_1545);
and U15 (N_15,In_1972,In_1406);
nand U16 (N_16,In_1874,In_617);
and U17 (N_17,In_975,In_1206);
nor U18 (N_18,In_53,In_1712);
and U19 (N_19,In_1090,In_1423);
and U20 (N_20,In_293,In_231);
and U21 (N_21,In_1709,In_569);
xor U22 (N_22,In_1591,In_24);
nand U23 (N_23,In_229,In_802);
nand U24 (N_24,In_482,In_1718);
or U25 (N_25,In_612,In_574);
xnor U26 (N_26,In_343,In_483);
nand U27 (N_27,In_1682,In_1041);
nor U28 (N_28,In_425,In_149);
xor U29 (N_29,In_666,In_1656);
and U30 (N_30,In_9,In_946);
nor U31 (N_31,In_669,In_1906);
and U32 (N_32,In_291,In_1375);
and U33 (N_33,In_1522,In_1634);
or U34 (N_34,In_844,In_675);
nand U35 (N_35,In_89,In_277);
nand U36 (N_36,In_105,In_1715);
xor U37 (N_37,In_285,In_1456);
and U38 (N_38,In_768,In_1266);
and U39 (N_39,In_676,In_1691);
nand U40 (N_40,In_1102,In_523);
nand U41 (N_41,In_1149,In_1885);
or U42 (N_42,In_1109,In_202);
xnor U43 (N_43,In_837,In_1202);
or U44 (N_44,In_1529,In_118);
nor U45 (N_45,In_829,In_1039);
nor U46 (N_46,In_784,In_681);
nor U47 (N_47,In_12,In_723);
nand U48 (N_48,In_969,In_1745);
nand U49 (N_49,In_1214,In_454);
or U50 (N_50,In_387,In_984);
or U51 (N_51,In_487,In_140);
nor U52 (N_52,In_165,In_270);
nand U53 (N_53,In_1777,In_1854);
nor U54 (N_54,In_1161,In_1608);
xnor U55 (N_55,In_1985,In_1458);
and U56 (N_56,In_412,In_155);
nor U57 (N_57,In_1670,In_1875);
xor U58 (N_58,In_1977,In_898);
xor U59 (N_59,In_655,In_958);
nand U60 (N_60,In_1204,In_1926);
xor U61 (N_61,In_1666,In_1821);
xor U62 (N_62,In_1068,In_264);
nand U63 (N_63,In_436,In_1073);
nor U64 (N_64,In_146,In_848);
nand U65 (N_65,In_951,In_154);
xnor U66 (N_66,In_901,In_1841);
xor U67 (N_67,In_1662,In_1574);
nand U68 (N_68,In_55,In_530);
nor U69 (N_69,In_1381,In_1060);
nor U70 (N_70,In_884,In_536);
or U71 (N_71,In_287,In_807);
nand U72 (N_72,In_601,In_1601);
nor U73 (N_73,In_187,In_1525);
nor U74 (N_74,In_1658,In_18);
nand U75 (N_75,In_1462,In_1493);
and U76 (N_76,In_1335,In_101);
or U77 (N_77,In_1640,In_559);
nand U78 (N_78,In_770,In_1627);
nor U79 (N_79,In_1365,In_1108);
nor U80 (N_80,In_532,In_361);
xor U81 (N_81,In_95,In_1105);
or U82 (N_82,In_396,In_581);
and U83 (N_83,In_1195,In_1716);
nor U84 (N_84,In_835,In_185);
nand U85 (N_85,In_1320,In_1075);
or U86 (N_86,In_1879,In_393);
nor U87 (N_87,In_1671,In_1850);
and U88 (N_88,In_1905,In_1891);
xor U89 (N_89,In_663,In_1603);
nor U90 (N_90,In_653,In_467);
nor U91 (N_91,In_236,In_214);
nor U92 (N_92,In_929,In_1776);
and U93 (N_93,In_1596,In_36);
and U94 (N_94,In_1962,In_1723);
xor U95 (N_95,In_145,In_1220);
xnor U96 (N_96,In_628,In_1588);
and U97 (N_97,In_1698,In_917);
and U98 (N_98,In_1693,In_1496);
xnor U99 (N_99,In_221,In_1762);
xnor U100 (N_100,In_607,In_883);
nand U101 (N_101,In_110,In_266);
xnor U102 (N_102,In_709,In_717);
xor U103 (N_103,In_1549,In_534);
nor U104 (N_104,In_1438,In_1274);
xnor U105 (N_105,In_90,In_767);
nand U106 (N_106,In_871,In_1418);
or U107 (N_107,In_1209,In_572);
and U108 (N_108,In_897,In_727);
or U109 (N_109,In_780,In_707);
xnor U110 (N_110,In_1157,In_1865);
and U111 (N_111,In_887,In_970);
xor U112 (N_112,In_1965,In_104);
and U113 (N_113,In_1755,In_326);
and U114 (N_114,In_578,In_45);
and U115 (N_115,In_1048,In_1159);
nand U116 (N_116,In_357,In_732);
or U117 (N_117,In_1675,In_1390);
or U118 (N_118,In_1293,In_1823);
nor U119 (N_119,In_196,In_1194);
nand U120 (N_120,In_510,In_724);
xnor U121 (N_121,In_432,In_228);
xnor U122 (N_122,In_699,In_875);
xor U123 (N_123,In_1654,In_74);
or U124 (N_124,In_1616,In_1870);
nor U125 (N_125,In_1641,In_1559);
nor U126 (N_126,In_347,In_1902);
nand U127 (N_127,In_481,In_128);
and U128 (N_128,In_1425,In_1459);
nor U129 (N_129,In_1292,In_1706);
or U130 (N_130,In_1401,In_8);
xnor U131 (N_131,In_1137,In_1582);
nor U132 (N_132,In_1468,In_862);
xnor U133 (N_133,In_783,In_1339);
xor U134 (N_134,In_1089,In_446);
nor U135 (N_135,In_1746,In_375);
xnor U136 (N_136,In_879,In_1396);
and U137 (N_137,In_1183,In_1642);
and U138 (N_138,In_573,In_1239);
nand U139 (N_139,In_431,In_1415);
xor U140 (N_140,In_1297,In_1753);
nor U141 (N_141,In_988,In_1334);
xor U142 (N_142,In_869,In_596);
xnor U143 (N_143,In_1974,In_469);
or U144 (N_144,In_448,In_1431);
nor U145 (N_145,In_956,In_1853);
nand U146 (N_146,In_1610,In_1125);
xor U147 (N_147,In_1484,In_1688);
and U148 (N_148,In_1534,In_1225);
nor U149 (N_149,In_1483,In_1155);
or U150 (N_150,In_1481,In_1457);
nor U151 (N_151,In_124,In_20);
xor U152 (N_152,In_923,In_504);
or U153 (N_153,In_1578,In_3);
and U154 (N_154,In_1319,In_842);
xnor U155 (N_155,In_400,In_1511);
and U156 (N_156,In_1081,In_1351);
and U157 (N_157,In_1101,In_708);
and U158 (N_158,In_804,In_398);
and U159 (N_159,In_394,In_1208);
nand U160 (N_160,In_260,In_38);
xnor U161 (N_161,In_595,In_1111);
or U162 (N_162,In_1628,In_905);
nand U163 (N_163,In_390,In_1007);
nand U164 (N_164,In_1808,In_1708);
or U165 (N_165,In_1681,In_1734);
or U166 (N_166,In_1349,In_1515);
nor U167 (N_167,In_1021,In_119);
xor U168 (N_168,In_1895,In_881);
nand U169 (N_169,In_1636,In_657);
nand U170 (N_170,In_257,In_664);
or U171 (N_171,In_1011,In_1045);
nor U172 (N_172,In_1028,In_1070);
nor U173 (N_173,In_376,In_1449);
and U174 (N_174,In_1594,In_186);
nand U175 (N_175,In_712,In_1766);
and U176 (N_176,In_1211,In_1846);
and U177 (N_177,In_493,In_735);
and U178 (N_178,In_509,In_518);
or U179 (N_179,In_1480,In_1038);
and U180 (N_180,In_91,In_1908);
nor U181 (N_181,In_283,In_1960);
or U182 (N_182,In_1429,In_543);
nand U183 (N_183,In_942,In_28);
nor U184 (N_184,In_1121,In_1427);
and U185 (N_185,In_160,In_1728);
nor U186 (N_186,In_363,In_834);
nand U187 (N_187,In_1976,In_745);
nand U188 (N_188,In_925,In_1849);
or U189 (N_189,In_379,In_1925);
nand U190 (N_190,In_994,In_1886);
nor U191 (N_191,In_411,In_241);
or U192 (N_192,In_1512,In_1687);
nand U193 (N_193,In_1954,In_716);
xnor U194 (N_194,In_1988,In_1218);
and U195 (N_195,In_1153,In_1702);
or U196 (N_196,In_637,In_1649);
or U197 (N_197,In_301,In_769);
nor U198 (N_198,In_1917,In_1027);
and U199 (N_199,In_129,In_41);
xor U200 (N_200,In_109,In_1852);
xor U201 (N_201,In_1275,In_1347);
and U202 (N_202,In_1667,In_981);
nand U203 (N_203,In_1050,In_544);
and U204 (N_204,In_1122,In_362);
nor U205 (N_205,In_1255,In_1502);
or U206 (N_206,In_1938,In_677);
nor U207 (N_207,In_381,In_405);
nand U208 (N_208,In_344,In_1362);
xor U209 (N_209,In_7,In_1245);
xnor U210 (N_210,In_1686,In_1747);
and U211 (N_211,In_1647,In_451);
nor U212 (N_212,In_1359,In_141);
xor U213 (N_213,In_86,In_1235);
or U214 (N_214,In_1203,In_1848);
nand U215 (N_215,In_113,In_849);
xnor U216 (N_216,In_1788,In_1690);
and U217 (N_217,In_1417,In_395);
nor U218 (N_218,In_1264,In_854);
nor U219 (N_219,In_1424,In_853);
nand U220 (N_220,In_391,In_1949);
xor U221 (N_221,In_670,In_1786);
or U222 (N_222,In_1719,In_58);
and U223 (N_223,In_1998,In_856);
nand U224 (N_224,In_242,In_413);
and U225 (N_225,In_505,In_1022);
nor U226 (N_226,In_1144,In_380);
nor U227 (N_227,In_824,In_1769);
nor U228 (N_228,In_1921,In_56);
and U229 (N_229,In_480,In_384);
and U230 (N_230,In_1129,In_1878);
nor U231 (N_231,In_1439,In_598);
or U232 (N_232,In_526,In_1699);
nor U233 (N_233,In_1343,In_265);
nand U234 (N_234,In_662,In_1311);
nand U235 (N_235,In_1345,In_249);
nand U236 (N_236,In_1552,In_1632);
or U237 (N_237,In_894,In_1781);
nor U238 (N_238,In_588,In_1504);
nor U239 (N_239,In_1200,In_1797);
or U240 (N_240,In_1989,In_1811);
xnor U241 (N_241,In_1802,In_476);
or U242 (N_242,In_694,In_1272);
nor U243 (N_243,In_1013,In_485);
nor U244 (N_244,In_713,In_1579);
xor U245 (N_245,In_1590,In_858);
or U246 (N_246,In_545,In_947);
nor U247 (N_247,In_1333,In_721);
or U248 (N_248,In_441,In_1492);
nor U249 (N_249,In_78,In_765);
xor U250 (N_250,In_537,In_1247);
nand U251 (N_251,In_188,In_1120);
xor U252 (N_252,In_967,In_1765);
nor U253 (N_253,In_439,In_139);
nor U254 (N_254,In_589,In_602);
and U255 (N_255,In_6,In_703);
and U256 (N_256,In_1151,In_54);
xor U257 (N_257,In_323,In_352);
nor U258 (N_258,In_1888,In_1817);
or U259 (N_259,In_126,In_643);
nand U260 (N_260,In_1934,In_410);
or U261 (N_261,In_1475,In_475);
or U262 (N_262,In_1677,In_88);
xor U263 (N_263,In_1744,In_1465);
nor U264 (N_264,In_64,In_909);
or U265 (N_265,In_1800,In_1694);
and U266 (N_266,In_63,In_27);
nor U267 (N_267,In_1500,In_1142);
nand U268 (N_268,In_1497,In_748);
and U269 (N_269,In_1684,In_1665);
nor U270 (N_270,In_564,In_1131);
or U271 (N_271,In_455,In_937);
nor U272 (N_272,In_939,In_191);
and U273 (N_273,In_157,In_255);
xor U274 (N_274,In_1196,In_240);
xor U275 (N_275,In_719,In_198);
and U276 (N_276,In_1831,In_1830);
nand U277 (N_277,In_556,In_121);
nand U278 (N_278,In_1759,In_1657);
nand U279 (N_279,In_616,In_1659);
xor U280 (N_280,In_415,In_1189);
nor U281 (N_281,In_1236,In_302);
xor U282 (N_282,In_1956,In_603);
nand U283 (N_283,In_1792,In_1408);
xnor U284 (N_284,In_1575,In_948);
nor U285 (N_285,In_1778,In_365);
xor U286 (N_286,In_1622,In_1585);
nor U287 (N_287,In_1498,In_739);
or U288 (N_288,In_1625,In_114);
nor U289 (N_289,In_540,In_1298);
nor U290 (N_290,In_1838,In_1863);
nand U291 (N_291,In_785,In_1645);
nand U292 (N_292,In_1093,In_1577);
nor U293 (N_293,In_654,In_576);
xnor U294 (N_294,In_1979,In_740);
and U295 (N_295,In_136,In_1561);
nand U296 (N_296,In_300,In_374);
nor U297 (N_297,In_1257,In_98);
nand U298 (N_298,In_679,In_1652);
and U299 (N_299,In_812,In_685);
xnor U300 (N_300,In_218,In_1543);
or U301 (N_301,In_1807,In_1271);
and U302 (N_302,In_516,In_633);
xnor U303 (N_303,In_1270,In_1637);
nand U304 (N_304,In_1328,In_1533);
and U305 (N_305,In_1971,In_96);
xor U306 (N_306,In_868,In_85);
nor U307 (N_307,In_319,In_1639);
and U308 (N_308,In_219,In_658);
or U309 (N_309,In_430,In_1899);
nor U310 (N_310,In_1689,In_308);
nor U311 (N_311,In_771,In_843);
xnor U312 (N_312,In_850,In_1633);
xnor U313 (N_313,In_652,In_1928);
and U314 (N_314,In_1489,In_1040);
nand U315 (N_315,In_1312,In_1944);
nor U316 (N_316,In_614,In_163);
xor U317 (N_317,In_304,In_1019);
xnor U318 (N_318,In_900,In_1741);
nor U319 (N_319,In_1931,In_1892);
nand U320 (N_320,In_192,In_491);
xnor U321 (N_321,In_312,In_1419);
and U322 (N_322,In_906,In_1826);
xnor U323 (N_323,In_1167,In_1341);
or U324 (N_324,In_1653,In_546);
nor U325 (N_325,In_1606,In_1858);
nor U326 (N_326,In_686,In_507);
xnor U327 (N_327,In_1147,In_1767);
nor U328 (N_328,In_1192,In_207);
nand U329 (N_329,In_120,In_305);
nor U330 (N_330,In_1761,In_1980);
or U331 (N_331,In_1467,In_1047);
and U332 (N_332,In_826,In_1442);
nand U333 (N_333,In_615,In_527);
or U334 (N_334,In_445,In_1933);
nand U335 (N_335,In_907,In_11);
nor U336 (N_336,In_102,In_1619);
xnor U337 (N_337,In_1150,In_1403);
nor U338 (N_338,In_1078,In_857);
xnor U339 (N_339,In_955,In_69);
xor U340 (N_340,In_369,In_865);
nor U341 (N_341,In_1323,In_424);
nor U342 (N_342,In_1384,In_440);
nor U343 (N_343,In_48,In_756);
nand U344 (N_344,In_1607,In_269);
nor U345 (N_345,In_1832,In_180);
and U346 (N_346,In_841,In_1984);
nand U347 (N_347,In_515,In_1941);
and U348 (N_348,In_1923,In_808);
and U349 (N_349,In_1049,In_1057);
nand U350 (N_350,In_1176,In_1791);
xnor U351 (N_351,In_392,In_733);
or U352 (N_352,In_1820,In_806);
nor U353 (N_353,In_281,In_1215);
and U354 (N_354,In_1613,In_1488);
and U355 (N_355,In_1572,In_370);
or U356 (N_356,In_316,In_1182);
and U357 (N_357,In_896,In_926);
and U358 (N_358,In_1082,In_142);
and U359 (N_359,In_1240,In_619);
and U360 (N_360,In_1920,In_10);
and U361 (N_361,In_1179,In_452);
xor U362 (N_362,In_608,In_1112);
or U363 (N_363,In_938,In_1981);
nand U364 (N_364,In_286,In_1281);
nor U365 (N_365,In_1736,In_962);
nor U366 (N_366,In_299,In_1581);
or U367 (N_367,In_1958,In_553);
nand U368 (N_368,In_1764,In_382);
nor U369 (N_369,In_971,In_1360);
and U370 (N_370,In_1420,In_1252);
and U371 (N_371,In_263,In_1623);
nand U372 (N_372,In_1104,In_468);
xnor U373 (N_373,In_704,In_1555);
and U374 (N_374,In_159,In_474);
xor U375 (N_375,In_490,In_1727);
and U376 (N_376,In_1907,In_83);
xor U377 (N_377,In_610,In_99);
or U378 (N_378,In_111,In_416);
nor U379 (N_379,In_60,In_1837);
nand U380 (N_380,In_200,In_645);
and U381 (N_381,In_1638,In_478);
nand U382 (N_382,In_998,In_1097);
nand U383 (N_383,In_1868,In_252);
and U384 (N_384,In_1326,In_1138);
xnor U385 (N_385,In_535,In_746);
nand U386 (N_386,In_1025,In_1517);
and U387 (N_387,In_35,In_903);
nor U388 (N_388,In_1253,In_1435);
nand U389 (N_389,In_580,In_1029);
or U390 (N_390,In_289,In_1969);
nor U391 (N_391,In_93,In_350);
nand U392 (N_392,In_1551,In_1726);
and U393 (N_393,In_1880,In_1617);
xor U394 (N_394,In_1433,In_755);
nor U395 (N_395,In_893,In_33);
or U396 (N_396,In_1205,In_94);
nand U397 (N_397,In_822,In_774);
and U398 (N_398,In_1002,In_1835);
xor U399 (N_399,In_1774,In_1668);
nand U400 (N_400,In_1655,In_1222);
xnor U401 (N_401,In_1422,In_1152);
or U402 (N_402,In_1170,In_1576);
xor U403 (N_403,In_718,In_309);
nand U404 (N_404,In_248,In_220);
and U405 (N_405,In_1066,In_1302);
nor U406 (N_406,In_1069,In_169);
nor U407 (N_407,In_1379,In_39);
and U408 (N_408,In_1986,In_1768);
nand U409 (N_409,In_34,In_1174);
or U410 (N_410,In_720,In_920);
xor U411 (N_411,In_1749,In_1478);
nand U412 (N_412,In_1451,In_1780);
and U413 (N_413,In_13,In_1898);
nand U414 (N_414,In_1141,In_1947);
and U415 (N_415,In_79,In_1190);
nand U416 (N_416,In_1197,In_310);
nand U417 (N_417,In_1454,In_953);
or U418 (N_418,In_1695,In_1304);
nor U419 (N_419,In_689,In_593);
or U420 (N_420,In_371,In_1571);
nor U421 (N_421,In_1404,In_542);
and U422 (N_422,In_423,In_1803);
nor U423 (N_423,In_389,In_1054);
xnor U424 (N_424,In_1893,In_928);
xnor U425 (N_425,In_230,In_1876);
and U426 (N_426,In_174,In_1284);
nor U427 (N_427,In_1946,In_1356);
or U428 (N_428,In_1020,In_1294);
xnor U429 (N_429,In_1630,In_47);
xnor U430 (N_430,In_1096,In_1733);
and U431 (N_431,In_334,In_1828);
nand U432 (N_432,In_43,In_1877);
nor U433 (N_433,In_1894,In_294);
nand U434 (N_434,In_600,In_1859);
xnor U435 (N_435,In_496,In_456);
nor U436 (N_436,In_1995,In_1935);
and U437 (N_437,In_71,In_832);
nand U438 (N_438,In_1554,In_1785);
or U439 (N_439,In_1856,In_566);
xnor U440 (N_440,In_1132,In_1991);
and U441 (N_441,In_1973,In_639);
or U442 (N_442,In_1618,In_125);
xor U443 (N_443,In_705,In_809);
nor U444 (N_444,In_747,In_649);
nand U445 (N_445,In_944,In_1023);
and U446 (N_446,In_453,In_1358);
and U447 (N_447,In_1509,In_1455);
xnor U448 (N_448,In_506,In_427);
nand U449 (N_449,In_1466,In_1626);
and U450 (N_450,In_954,In_1123);
nand U451 (N_451,In_479,In_1321);
xor U452 (N_452,In_729,In_1296);
nor U453 (N_453,In_800,In_223);
nand U454 (N_454,In_514,In_641);
and U455 (N_455,In_1243,In_1524);
xnor U456 (N_456,In_463,In_1177);
nand U457 (N_457,In_648,In_75);
nand U458 (N_458,In_1172,In_656);
or U459 (N_459,In_65,In_1782);
and U460 (N_460,In_62,In_5);
nor U461 (N_461,In_565,In_1737);
nand U462 (N_462,In_1872,In_1268);
and U463 (N_463,In_919,In_1996);
xor U464 (N_464,In_359,In_216);
nand U465 (N_465,In_618,In_122);
or U466 (N_466,In_1446,In_1254);
xnor U467 (N_467,In_674,In_1307);
and U468 (N_468,In_276,In_766);
and U469 (N_469,In_1160,In_199);
or U470 (N_470,In_1077,In_1091);
and U471 (N_471,In_1338,In_1866);
or U472 (N_472,In_1707,In_181);
and U473 (N_473,In_1697,In_1916);
nor U474 (N_474,In_886,In_1535);
nor U475 (N_475,In_358,In_138);
and U476 (N_476,In_1664,In_133);
or U477 (N_477,In_1184,In_1076);
nor U478 (N_478,In_1226,In_1308);
nor U479 (N_479,In_1314,In_682);
and U480 (N_480,In_793,In_959);
or U481 (N_481,In_336,In_1519);
or U482 (N_482,In_345,In_342);
or U483 (N_483,In_1315,In_1487);
nor U484 (N_484,In_1514,In_798);
or U485 (N_485,In_754,In_972);
nand U486 (N_486,In_985,In_1605);
nor U487 (N_487,In_1685,In_1883);
nand U488 (N_488,In_1470,In_1380);
nand U489 (N_489,In_1942,In_1873);
nor U490 (N_490,In_815,In_321);
or U491 (N_491,In_97,In_1553);
nand U492 (N_492,In_1646,In_1374);
or U493 (N_493,In_1373,In_979);
and U494 (N_494,In_1510,In_627);
xor U495 (N_495,In_1825,In_1683);
nand U496 (N_496,In_1904,In_1756);
nand U497 (N_497,In_563,In_642);
or U498 (N_498,In_1644,In_284);
xnor U499 (N_499,In_605,In_204);
nand U500 (N_500,In_148,In_1145);
nor U501 (N_501,In_116,In_52);
xnor U502 (N_502,In_952,In_761);
or U503 (N_503,In_1232,In_1531);
or U504 (N_504,In_976,In_650);
and U505 (N_505,In_1913,In_224);
and U506 (N_506,In_1922,In_466);
nand U507 (N_507,In_1428,In_845);
nor U508 (N_508,In_348,In_484);
nand U509 (N_509,In_1595,In_1700);
nor U510 (N_510,In_684,In_830);
nor U511 (N_511,In_584,In_1348);
nor U512 (N_512,In_1186,In_562);
nor U513 (N_513,In_70,In_778);
or U514 (N_514,In_1386,In_1441);
nand U515 (N_515,In_59,In_1929);
nand U516 (N_516,In_779,In_1754);
and U517 (N_517,In_1523,In_1256);
nor U518 (N_518,In_1717,In_1809);
or U519 (N_519,In_238,In_1609);
and U520 (N_520,In_1635,In_1148);
nand U521 (N_521,In_176,In_1842);
and U522 (N_522,In_1074,In_486);
xor U523 (N_523,In_437,In_1568);
or U524 (N_524,In_715,In_501);
or U525 (N_525,In_1357,In_1889);
nand U526 (N_526,In_1412,In_1355);
nand U527 (N_527,In_983,In_1839);
nor U528 (N_528,In_1250,In_1432);
xnor U529 (N_529,In_1290,In_494);
or U530 (N_530,In_151,In_910);
or U531 (N_531,In_915,In_1461);
xor U532 (N_532,In_421,In_1409);
xnor U533 (N_533,In_753,In_1987);
nor U534 (N_534,In_26,In_706);
xnor U535 (N_535,In_1447,In_1010);
and U536 (N_536,In_46,In_1957);
nor U537 (N_537,In_833,In_882);
and U538 (N_538,In_1165,In_620);
or U539 (N_539,In_1213,In_1673);
nor U540 (N_540,In_517,In_1516);
nor U541 (N_541,In_1146,In_0);
nor U542 (N_542,In_1118,In_1586);
xnor U543 (N_543,In_1789,In_1300);
nand U544 (N_544,In_736,In_173);
xor U545 (N_545,In_930,In_303);
nor U546 (N_546,In_1363,In_1532);
or U547 (N_547,In_1471,In_647);
or U548 (N_548,In_15,In_640);
and U549 (N_549,In_1611,In_582);
nand U550 (N_550,In_190,In_1909);
nand U551 (N_551,In_555,In_1758);
or U552 (N_552,In_1313,In_1847);
nand U553 (N_553,In_1798,In_730);
nor U554 (N_554,In_385,In_1286);
xnor U555 (N_555,In_1421,In_1722);
and U556 (N_556,In_1430,In_714);
and U557 (N_557,In_789,In_1389);
and U558 (N_558,In_57,In_1951);
or U559 (N_559,In_531,In_1237);
or U560 (N_560,In_847,In_1964);
xor U561 (N_561,In_30,In_738);
or U562 (N_562,In_488,In_1169);
or U563 (N_563,In_1721,In_377);
xor U564 (N_564,In_1273,In_1955);
nor U565 (N_565,In_796,In_821);
and U566 (N_566,In_1473,In_888);
or U567 (N_567,In_397,In_213);
nor U568 (N_568,In_1814,In_996);
xnor U569 (N_569,In_541,In_1106);
nor U570 (N_570,In_1259,In_1939);
or U571 (N_571,In_473,In_4);
xnor U572 (N_572,In_777,In_579);
nor U573 (N_573,In_1503,In_673);
xor U574 (N_574,In_859,In_1918);
or U575 (N_575,In_1395,In_693);
and U576 (N_576,In_1799,In_307);
nor U577 (N_577,In_1385,In_794);
and U578 (N_578,In_791,In_1344);
and U579 (N_579,In_683,In_590);
and U580 (N_580,In_1783,In_44);
xnor U581 (N_581,In_813,In_1757);
xor U582 (N_582,In_25,In_1394);
and U583 (N_583,In_889,In_1030);
nor U584 (N_584,In_346,In_823);
or U585 (N_585,In_329,In_1221);
or U586 (N_586,In_106,In_1672);
or U587 (N_587,In_409,In_150);
and U588 (N_588,In_792,In_817);
nand U589 (N_589,In_1738,In_322);
and U590 (N_590,In_776,In_918);
and U591 (N_591,In_1140,In_444);
and U592 (N_592,In_1103,In_1680);
nor U593 (N_593,In_408,In_1017);
or U594 (N_594,In_1134,In_297);
and U595 (N_595,In_168,In_622);
and U596 (N_596,In_1631,In_973);
xnor U597 (N_597,In_1650,In_696);
xnor U598 (N_598,In_1824,In_428);
nor U599 (N_599,In_867,In_722);
xnor U600 (N_600,In_460,In_1064);
nor U601 (N_601,In_103,In_1711);
nor U602 (N_602,In_668,In_960);
xnor U603 (N_603,In_550,In_31);
nand U604 (N_604,In_711,In_651);
and U605 (N_605,In_153,In_1331);
nor U606 (N_606,In_1279,In_1185);
nor U607 (N_607,In_1198,In_1217);
or U608 (N_608,In_1966,In_1032);
xnor U609 (N_609,In_355,In_836);
and U610 (N_610,In_1229,In_1819);
nor U611 (N_611,In_1024,In_672);
nor U612 (N_612,In_1663,In_1570);
and U613 (N_613,In_164,In_356);
xor U614 (N_614,In_575,In_1742);
or U615 (N_615,In_890,In_1887);
nor U616 (N_616,In_678,In_877);
nand U617 (N_617,In_1014,In_1705);
nor U618 (N_618,In_492,In_1772);
or U619 (N_619,In_67,In_876);
nor U620 (N_620,In_1720,In_76);
or U621 (N_621,In_1350,In_968);
nand U622 (N_622,In_37,In_1562);
or U623 (N_623,In_943,In_913);
nand U624 (N_624,In_742,In_1414);
nand U625 (N_625,In_1310,In_1227);
or U626 (N_626,In_1615,In_162);
or U627 (N_627,In_80,In_1952);
or U628 (N_628,In_1937,In_372);
xnor U629 (N_629,In_646,In_349);
and U630 (N_630,In_201,In_1377);
and U631 (N_631,In_1400,In_511);
xor U632 (N_632,In_1915,In_1790);
nand U633 (N_633,In_1536,In_1369);
or U634 (N_634,In_772,In_1262);
or U635 (N_635,In_354,In_1434);
xor U636 (N_636,In_1544,In_1426);
and U637 (N_637,In_1530,In_1862);
nor U638 (N_638,In_1678,In_1114);
xnor U639 (N_639,In_1950,In_1845);
nand U640 (N_640,In_318,In_1527);
and U641 (N_641,In_1464,In_1413);
or U642 (N_642,In_1537,In_1624);
nor U643 (N_643,In_1233,In_577);
xnor U644 (N_644,In_360,In_811);
nand U645 (N_645,In_964,In_1513);
or U646 (N_646,In_512,In_335);
xor U647 (N_647,In_183,In_1936);
nor U648 (N_648,In_1558,In_320);
xor U649 (N_649,In_251,In_1731);
nor U650 (N_650,In_1305,In_1978);
and U651 (N_651,In_127,In_1116);
and U652 (N_652,In_940,In_470);
or U653 (N_653,In_1135,In_1280);
or U654 (N_654,In_1026,In_846);
xnor U655 (N_655,In_2,In_1679);
xnor U656 (N_656,In_591,In_1416);
xnor U657 (N_657,In_922,In_1071);
and U658 (N_658,In_1771,In_982);
or U659 (N_659,In_1042,In_936);
or U660 (N_660,In_625,In_1382);
nor U661 (N_661,In_1822,In_1834);
nand U662 (N_662,In_1486,In_1748);
or U663 (N_663,In_14,In_166);
and U664 (N_664,In_1087,In_549);
or U665 (N_665,In_1330,In_690);
nand U666 (N_666,In_1393,In_551);
nor U667 (N_667,In_1055,In_457);
and U668 (N_668,In_1714,In_1482);
or U669 (N_669,In_737,In_1443);
xnor U670 (N_670,In_1589,In_819);
nor U671 (N_671,In_1156,In_1896);
nand U672 (N_672,In_271,In_855);
nand U673 (N_673,In_1518,In_1676);
and U674 (N_674,In_710,In_611);
nor U675 (N_675,In_760,In_1364);
and U676 (N_676,In_420,In_1246);
and U677 (N_677,In_443,In_801);
and U678 (N_678,In_383,In_1450);
nor U679 (N_679,In_781,In_66);
or U680 (N_680,In_1818,In_144);
or U681 (N_681,In_1361,In_1810);
and U682 (N_682,In_1230,In_560);
nand U683 (N_683,In_980,In_752);
nand U684 (N_684,In_1099,In_1299);
xnor U685 (N_685,In_253,In_665);
nor U686 (N_686,In_1932,In_892);
nand U687 (N_687,In_314,In_1463);
nand U688 (N_688,In_1560,In_695);
or U689 (N_689,In_552,In_1086);
xor U690 (N_690,In_1840,In_503);
xor U691 (N_691,In_1860,In_1813);
and U692 (N_692,In_1477,In_1340);
nand U693 (N_693,In_171,In_233);
xnor U694 (N_694,In_764,In_529);
xor U695 (N_695,In_262,In_1201);
nor U696 (N_696,In_606,In_1547);
and U697 (N_697,In_404,In_571);
xor U698 (N_698,In_254,In_1546);
xnor U699 (N_699,In_609,In_261);
nand U700 (N_700,In_1910,In_1963);
xor U701 (N_701,In_799,In_1005);
and U702 (N_702,In_1336,In_1260);
nor U703 (N_703,In_1216,In_1061);
xnor U704 (N_704,In_353,In_726);
nor U705 (N_705,In_828,In_895);
xnor U706 (N_706,In_1175,In_426);
or U707 (N_707,In_1927,In_1557);
xnor U708 (N_708,In_256,In_325);
and U709 (N_709,In_1354,In_311);
xnor U710 (N_710,In_986,In_137);
xnor U711 (N_711,In_1110,In_1999);
and U712 (N_712,In_586,In_179);
nor U713 (N_713,In_989,In_1538);
nand U714 (N_714,In_366,In_1773);
nor U715 (N_715,In_816,In_290);
and U716 (N_716,In_1324,In_1660);
nand U717 (N_717,In_1126,In_1188);
or U718 (N_718,In_1526,In_680);
xnor U719 (N_719,In_1474,In_629);
nand U720 (N_720,In_1062,In_902);
or U721 (N_721,In_1238,In_222);
xnor U722 (N_722,In_1732,In_749);
nor U723 (N_723,In_1499,In_489);
and U724 (N_724,In_1669,In_561);
and U725 (N_725,In_1540,In_1692);
nor U726 (N_726,In_206,In_1930);
and U727 (N_727,In_1703,In_203);
nor U728 (N_728,In_131,In_1173);
xnor U729 (N_729,In_1805,In_1864);
nor U730 (N_730,In_1648,In_921);
nor U731 (N_731,In_1224,In_741);
nor U732 (N_732,In_1760,In_701);
or U733 (N_733,In_1505,In_414);
xor U734 (N_734,In_1994,In_1882);
and U735 (N_735,In_597,In_557);
or U736 (N_736,In_1861,In_751);
and U737 (N_737,In_1178,In_32);
nand U738 (N_738,In_1012,In_1548);
and U739 (N_739,In_500,In_1643);
and U740 (N_740,In_1583,In_521);
and U741 (N_741,In_1440,In_1378);
and U742 (N_742,In_406,In_613);
nand U743 (N_743,In_1851,In_831);
and U744 (N_744,In_296,In_698);
or U745 (N_745,In_1383,In_433);
nor U746 (N_746,In_61,In_1587);
or U747 (N_747,In_156,In_1436);
nand U748 (N_748,In_1563,In_1083);
nor U749 (N_749,In_1191,In_941);
nor U750 (N_750,In_84,In_340);
or U751 (N_751,In_21,In_1052);
nand U752 (N_752,In_1843,In_1261);
or U753 (N_753,In_1967,In_870);
or U754 (N_754,In_874,In_1444);
and U755 (N_755,In_1193,In_465);
xor U756 (N_756,In_1600,In_1539);
nand U757 (N_757,In_599,In_851);
nor U758 (N_758,In_1033,In_1485);
or U759 (N_759,In_993,In_182);
and U760 (N_760,In_68,In_1479);
and U761 (N_761,In_1735,In_1829);
and U762 (N_762,In_272,In_418);
nand U763 (N_763,In_16,In_247);
nor U764 (N_764,In_1491,In_963);
and U765 (N_765,In_604,In_1065);
xor U766 (N_766,In_1620,In_1521);
or U767 (N_767,In_243,In_932);
or U768 (N_768,In_1107,In_1763);
nand U769 (N_769,In_702,In_966);
nor U770 (N_770,In_554,In_1352);
and U771 (N_771,In_1016,In_1058);
nand U772 (N_772,In_864,In_508);
nor U773 (N_773,In_195,In_1210);
nand U774 (N_774,In_212,In_1696);
nor U775 (N_775,In_1881,In_911);
nor U776 (N_776,In_873,In_1602);
xor U777 (N_777,In_1796,In_934);
nor U778 (N_778,In_1729,In_587);
nor U779 (N_779,In_1469,In_567);
or U780 (N_780,In_497,In_700);
and U781 (N_781,In_1541,In_757);
xnor U782 (N_782,In_306,In_1793);
and U783 (N_783,In_1318,In_471);
nor U784 (N_784,In_1219,In_1051);
xnor U785 (N_785,In_1388,In_891);
nor U786 (N_786,In_1162,In_1372);
or U787 (N_787,In_1006,In_172);
nor U788 (N_788,In_1912,In_1397);
and U789 (N_789,In_525,In_1306);
xnor U790 (N_790,In_1506,In_1228);
nand U791 (N_791,In_332,In_1258);
and U792 (N_792,In_950,In_401);
xor U793 (N_793,In_1871,In_341);
xor U794 (N_794,In_1855,In_1322);
nand U795 (N_795,In_1752,In_1283);
nand U796 (N_796,In_1158,In_351);
nor U797 (N_797,In_1614,In_1405);
or U798 (N_798,In_548,In_1914);
nand U799 (N_799,In_916,In_1704);
nor U800 (N_800,In_403,In_945);
or U801 (N_801,In_852,In_364);
xor U802 (N_802,In_1884,In_1740);
xnor U803 (N_803,In_621,In_1448);
nand U804 (N_804,In_999,In_762);
nand U805 (N_805,In_1143,In_388);
nor U806 (N_806,In_459,In_1795);
or U807 (N_807,In_1399,In_1924);
and U808 (N_808,In_1004,In_1337);
nand U809 (N_809,In_860,In_992);
and U810 (N_810,In_840,In_547);
xor U811 (N_811,In_743,In_1085);
xnor U812 (N_812,In_520,In_1453);
and U813 (N_813,In_193,In_1507);
xnor U814 (N_814,In_1009,In_1003);
and U815 (N_815,In_1542,In_991);
nor U816 (N_816,In_1368,In_333);
and U817 (N_817,In_594,In_795);
nor U818 (N_818,In_1376,In_787);
nor U819 (N_819,In_585,In_17);
or U820 (N_820,In_1410,In_1036);
nor U821 (N_821,In_1325,In_1567);
and U822 (N_822,In_1674,In_1001);
or U823 (N_823,In_1566,In_1730);
nor U824 (N_824,In_667,In_1327);
and U825 (N_825,In_782,In_1168);
nand U826 (N_826,In_1346,In_863);
or U827 (N_827,In_1295,In_1251);
nor U828 (N_828,In_1556,In_1701);
nor U829 (N_829,In_449,In_1015);
nand U830 (N_830,In_592,In_226);
nand U831 (N_831,In_1181,In_1770);
xor U832 (N_832,In_914,In_147);
and U833 (N_833,In_337,In_1833);
and U834 (N_834,In_1550,In_1370);
nor U835 (N_835,In_880,In_538);
nor U836 (N_836,In_1897,In_92);
or U837 (N_837,In_659,In_838);
xnor U838 (N_838,In_1584,In_908);
or U839 (N_839,In_117,In_1180);
xor U840 (N_840,In_167,In_990);
nand U841 (N_841,In_632,In_1495);
nor U842 (N_842,In_189,In_177);
or U843 (N_843,In_644,In_1263);
nor U844 (N_844,In_1139,In_378);
nand U845 (N_845,In_498,In_861);
nand U846 (N_846,In_818,In_744);
xor U847 (N_847,In_539,In_1094);
xnor U848 (N_848,In_234,In_1476);
or U849 (N_849,In_631,In_1604);
and U850 (N_850,In_1098,In_495);
or U851 (N_851,In_623,In_1342);
xnor U852 (N_852,In_1836,In_205);
or U853 (N_853,In_292,In_1391);
nand U854 (N_854,In_935,In_1911);
or U855 (N_855,In_123,In_1816);
or U856 (N_856,In_1046,In_825);
nand U857 (N_857,In_107,In_135);
nand U858 (N_858,In_274,In_635);
nand U859 (N_859,In_73,In_211);
nor U860 (N_860,In_49,In_1043);
and U861 (N_861,In_878,In_1407);
and U862 (N_862,In_1751,In_1593);
and U863 (N_863,In_422,In_1092);
xor U864 (N_864,In_1801,In_1968);
nor U865 (N_865,In_773,In_933);
and U866 (N_866,In_386,In_1940);
nor U867 (N_867,In_583,In_51);
nor U868 (N_868,In_1629,In_1044);
xor U869 (N_869,In_246,In_209);
and U870 (N_870,In_965,In_1724);
xor U871 (N_871,In_1212,In_1367);
nand U872 (N_872,In_1472,In_1316);
xnor U873 (N_873,In_1018,In_931);
xnor U874 (N_874,In_237,In_447);
and U875 (N_875,In_1784,In_108);
nor U876 (N_876,In_1621,In_184);
nor U877 (N_877,In_194,In_924);
nand U878 (N_878,In_464,In_407);
or U879 (N_879,In_660,In_1207);
xnor U880 (N_880,In_1199,In_1857);
and U881 (N_881,In_368,In_278);
or U882 (N_882,In_275,In_1080);
xnor U883 (N_883,In_763,In_77);
nand U884 (N_884,In_1598,In_904);
nand U885 (N_885,In_499,In_1);
and U886 (N_886,In_788,In_429);
nor U887 (N_887,In_1309,In_1775);
xnor U888 (N_888,In_327,In_1961);
nor U889 (N_889,In_1970,In_1990);
nor U890 (N_890,In_1997,In_1779);
nand U891 (N_891,In_417,In_197);
nor U892 (N_892,In_1460,In_1244);
and U893 (N_893,In_558,In_1154);
nand U894 (N_894,In_250,In_687);
and U895 (N_895,In_1329,In_1000);
nand U896 (N_896,In_814,In_178);
or U897 (N_897,In_961,In_1945);
nor U898 (N_898,In_1528,In_298);
nand U899 (N_899,In_1276,In_1794);
xor U900 (N_900,In_524,In_1287);
nand U901 (N_901,In_1901,In_112);
xnor U902 (N_902,In_40,In_1059);
nand U903 (N_903,In_1234,In_502);
nor U904 (N_904,In_1387,In_912);
nand U905 (N_905,In_258,In_279);
nand U906 (N_906,In_624,In_1520);
nand U907 (N_907,In_324,In_450);
nor U908 (N_908,In_1231,In_1804);
nand U909 (N_909,In_775,In_1301);
nand U910 (N_910,In_1445,In_1291);
and U911 (N_911,In_1031,In_72);
and U912 (N_912,In_1166,In_630);
and U913 (N_913,In_885,In_827);
or U914 (N_914,In_132,In_1128);
and U915 (N_915,In_1437,In_1573);
nand U916 (N_916,In_1739,In_1269);
nor U917 (N_917,In_1317,In_215);
nand U918 (N_918,In_245,In_317);
nand U919 (N_919,In_367,In_513);
nor U920 (N_920,In_19,In_1501);
nand U921 (N_921,In_1241,In_280);
and U922 (N_922,In_143,In_528);
and U923 (N_923,In_158,In_1402);
and U924 (N_924,In_688,In_1597);
nor U925 (N_925,In_872,In_1983);
nor U926 (N_926,In_1124,In_438);
nor U927 (N_927,In_1113,In_759);
nand U928 (N_928,In_1136,In_1332);
or U929 (N_929,In_839,In_100);
nor U930 (N_930,In_949,In_1163);
or U931 (N_931,In_731,In_259);
nand U932 (N_932,In_1959,In_1710);
or U933 (N_933,In_786,In_1993);
and U934 (N_934,In_1366,In_50);
xor U935 (N_935,In_115,In_1564);
nor U936 (N_936,In_1072,In_273);
or U937 (N_937,In_1242,In_338);
xnor U938 (N_938,In_313,In_803);
and U939 (N_939,In_1095,In_1267);
or U940 (N_940,In_1713,In_330);
xor U941 (N_941,In_636,In_1119);
nand U942 (N_942,In_995,In_1392);
nand U943 (N_943,In_927,In_1411);
and U944 (N_944,In_1869,In_899);
and U945 (N_945,In_244,In_1288);
xnor U946 (N_946,In_820,In_1900);
nand U947 (N_947,In_435,In_1806);
nor U948 (N_948,In_1651,In_152);
nand U949 (N_949,In_977,In_402);
nand U950 (N_950,In_1248,In_1750);
and U951 (N_951,In_1063,In_282);
and U952 (N_952,In_134,In_1661);
and U953 (N_953,In_1223,In_458);
or U954 (N_954,In_1948,In_1812);
nand U955 (N_955,In_1079,In_692);
nor U956 (N_956,In_797,In_462);
and U957 (N_957,In_1034,In_208);
xnor U958 (N_958,In_1494,In_1084);
xnor U959 (N_959,In_461,In_1115);
or U960 (N_960,In_331,In_758);
nand U961 (N_961,In_1725,In_434);
and U962 (N_962,In_568,In_130);
and U963 (N_963,In_339,In_210);
nand U964 (N_964,In_522,In_175);
nand U965 (N_965,In_239,In_295);
nand U966 (N_966,In_1743,In_1992);
xor U967 (N_967,In_519,In_1282);
or U968 (N_968,In_570,In_697);
nor U969 (N_969,In_81,In_1100);
nor U970 (N_970,In_1035,In_268);
nand U971 (N_971,In_1903,In_232);
nand U972 (N_972,In_328,In_1490);
or U973 (N_973,In_1277,In_725);
nor U974 (N_974,In_442,In_42);
nor U975 (N_975,In_1569,In_1982);
xnor U976 (N_976,In_477,In_1067);
nand U977 (N_977,In_419,In_728);
nor U978 (N_978,In_1053,In_1890);
xor U979 (N_979,In_810,In_1612);
nand U980 (N_980,In_978,In_1164);
or U981 (N_981,In_1953,In_288);
xor U982 (N_982,In_1037,In_638);
or U983 (N_983,In_87,In_315);
and U984 (N_984,In_866,In_1130);
nand U985 (N_985,In_1303,In_1117);
nor U986 (N_986,In_235,In_626);
or U987 (N_987,In_1592,In_661);
or U988 (N_988,In_1371,In_805);
nor U989 (N_989,In_734,In_1867);
or U990 (N_990,In_957,In_1353);
or U991 (N_991,In_1844,In_790);
nor U992 (N_992,In_217,In_691);
nand U993 (N_993,In_472,In_1133);
nand U994 (N_994,In_170,In_1285);
nor U995 (N_995,In_1452,In_23);
or U996 (N_996,In_1265,In_1580);
nor U997 (N_997,In_974,In_1398);
or U998 (N_998,In_1249,In_1278);
xor U999 (N_999,In_267,In_533);
or U1000 (N_1000,N_998,N_905);
nor U1001 (N_1001,N_592,N_896);
nor U1002 (N_1002,N_441,N_555);
nand U1003 (N_1003,N_201,N_384);
and U1004 (N_1004,N_529,N_541);
nand U1005 (N_1005,N_649,N_343);
and U1006 (N_1006,N_62,N_933);
or U1007 (N_1007,N_879,N_178);
and U1008 (N_1008,N_488,N_884);
or U1009 (N_1009,N_18,N_744);
or U1010 (N_1010,N_22,N_74);
and U1011 (N_1011,N_758,N_956);
nor U1012 (N_1012,N_825,N_146);
xor U1013 (N_1013,N_557,N_856);
nand U1014 (N_1014,N_623,N_100);
and U1015 (N_1015,N_280,N_121);
xnor U1016 (N_1016,N_218,N_323);
nor U1017 (N_1017,N_745,N_83);
and U1018 (N_1018,N_590,N_371);
nand U1019 (N_1019,N_571,N_167);
xnor U1020 (N_1020,N_766,N_81);
or U1021 (N_1021,N_250,N_662);
and U1022 (N_1022,N_863,N_138);
or U1023 (N_1023,N_331,N_420);
or U1024 (N_1024,N_411,N_593);
nand U1025 (N_1025,N_834,N_228);
nand U1026 (N_1026,N_47,N_530);
nor U1027 (N_1027,N_97,N_765);
nor U1028 (N_1028,N_542,N_276);
and U1029 (N_1029,N_891,N_365);
xnor U1030 (N_1030,N_775,N_175);
nand U1031 (N_1031,N_715,N_646);
or U1032 (N_1032,N_612,N_814);
nor U1033 (N_1033,N_777,N_379);
nand U1034 (N_1034,N_34,N_33);
nor U1035 (N_1035,N_196,N_174);
xnor U1036 (N_1036,N_561,N_477);
xnor U1037 (N_1037,N_251,N_734);
and U1038 (N_1038,N_215,N_628);
or U1039 (N_1039,N_304,N_566);
and U1040 (N_1040,N_153,N_767);
nand U1041 (N_1041,N_398,N_82);
nor U1042 (N_1042,N_999,N_315);
xnor U1043 (N_1043,N_978,N_110);
xor U1044 (N_1044,N_974,N_476);
xor U1045 (N_1045,N_386,N_728);
nor U1046 (N_1046,N_963,N_988);
and U1047 (N_1047,N_548,N_647);
and U1048 (N_1048,N_327,N_526);
nand U1049 (N_1049,N_602,N_811);
and U1050 (N_1050,N_221,N_869);
or U1051 (N_1051,N_692,N_805);
xnor U1052 (N_1052,N_546,N_847);
and U1053 (N_1053,N_372,N_204);
xnor U1054 (N_1054,N_749,N_6);
and U1055 (N_1055,N_120,N_313);
nor U1056 (N_1056,N_418,N_717);
xnor U1057 (N_1057,N_229,N_536);
and U1058 (N_1058,N_779,N_757);
or U1059 (N_1059,N_684,N_389);
xnor U1060 (N_1060,N_414,N_917);
nor U1061 (N_1061,N_932,N_822);
nor U1062 (N_1062,N_360,N_532);
nand U1063 (N_1063,N_293,N_544);
nand U1064 (N_1064,N_446,N_818);
nor U1065 (N_1065,N_497,N_405);
nor U1066 (N_1066,N_815,N_36);
or U1067 (N_1067,N_867,N_528);
and U1068 (N_1068,N_634,N_622);
xnor U1069 (N_1069,N_984,N_754);
and U1070 (N_1070,N_660,N_244);
xnor U1071 (N_1071,N_392,N_465);
xor U1072 (N_1072,N_579,N_400);
and U1073 (N_1073,N_278,N_443);
nor U1074 (N_1074,N_494,N_816);
xnor U1075 (N_1075,N_898,N_299);
or U1076 (N_1076,N_104,N_720);
and U1077 (N_1077,N_596,N_407);
and U1078 (N_1078,N_58,N_191);
or U1079 (N_1079,N_56,N_923);
xor U1080 (N_1080,N_733,N_194);
or U1081 (N_1081,N_844,N_15);
nand U1082 (N_1082,N_165,N_187);
and U1083 (N_1083,N_514,N_325);
nor U1084 (N_1084,N_243,N_525);
nor U1085 (N_1085,N_145,N_585);
nor U1086 (N_1086,N_394,N_703);
xor U1087 (N_1087,N_283,N_752);
nand U1088 (N_1088,N_179,N_707);
nand U1089 (N_1089,N_479,N_568);
or U1090 (N_1090,N_412,N_272);
nand U1091 (N_1091,N_269,N_506);
or U1092 (N_1092,N_713,N_359);
nand U1093 (N_1093,N_621,N_743);
nand U1094 (N_1094,N_312,N_750);
xor U1095 (N_1095,N_318,N_172);
and U1096 (N_1096,N_252,N_144);
nand U1097 (N_1097,N_42,N_181);
and U1098 (N_1098,N_382,N_116);
or U1099 (N_1099,N_245,N_527);
nor U1100 (N_1100,N_989,N_791);
nor U1101 (N_1101,N_762,N_182);
or U1102 (N_1102,N_613,N_581);
and U1103 (N_1103,N_603,N_729);
and U1104 (N_1104,N_422,N_721);
nor U1105 (N_1105,N_778,N_403);
nor U1106 (N_1106,N_285,N_841);
nand U1107 (N_1107,N_901,N_641);
and U1108 (N_1108,N_375,N_408);
or U1109 (N_1109,N_339,N_358);
nor U1110 (N_1110,N_366,N_550);
nor U1111 (N_1111,N_162,N_404);
and U1112 (N_1112,N_977,N_639);
nor U1113 (N_1113,N_210,N_589);
nand U1114 (N_1114,N_785,N_21);
and U1115 (N_1115,N_888,N_428);
nand U1116 (N_1116,N_421,N_920);
and U1117 (N_1117,N_521,N_483);
nor U1118 (N_1118,N_291,N_85);
or U1119 (N_1119,N_935,N_732);
nand U1120 (N_1120,N_666,N_677);
nor U1121 (N_1121,N_311,N_338);
nor U1122 (N_1122,N_604,N_560);
nand U1123 (N_1123,N_909,N_694);
and U1124 (N_1124,N_595,N_511);
nand U1125 (N_1125,N_334,N_664);
xnor U1126 (N_1126,N_329,N_760);
nor U1127 (N_1127,N_537,N_284);
nand U1128 (N_1128,N_435,N_474);
or U1129 (N_1129,N_918,N_615);
and U1130 (N_1130,N_992,N_580);
nor U1131 (N_1131,N_328,N_129);
and U1132 (N_1132,N_72,N_808);
xor U1133 (N_1133,N_246,N_214);
nand U1134 (N_1134,N_451,N_168);
xnor U1135 (N_1135,N_915,N_256);
xor U1136 (N_1136,N_253,N_468);
nand U1137 (N_1137,N_281,N_876);
nor U1138 (N_1138,N_130,N_960);
xnor U1139 (N_1139,N_13,N_75);
xor U1140 (N_1140,N_57,N_361);
and U1141 (N_1141,N_948,N_682);
or U1142 (N_1142,N_254,N_597);
or U1143 (N_1143,N_79,N_642);
xnor U1144 (N_1144,N_440,N_378);
xnor U1145 (N_1145,N_12,N_286);
xor U1146 (N_1146,N_881,N_473);
or U1147 (N_1147,N_619,N_922);
xor U1148 (N_1148,N_510,N_279);
xor U1149 (N_1149,N_688,N_255);
xor U1150 (N_1150,N_108,N_994);
and U1151 (N_1151,N_906,N_774);
and U1152 (N_1152,N_46,N_836);
nand U1153 (N_1153,N_582,N_309);
or U1154 (N_1154,N_442,N_517);
nand U1155 (N_1155,N_50,N_697);
or U1156 (N_1156,N_310,N_648);
nand U1157 (N_1157,N_868,N_51);
nor U1158 (N_1158,N_349,N_979);
nand U1159 (N_1159,N_410,N_711);
nor U1160 (N_1160,N_300,N_30);
nand U1161 (N_1161,N_678,N_258);
nand U1162 (N_1162,N_340,N_377);
xnor U1163 (N_1163,N_429,N_423);
and U1164 (N_1164,N_89,N_454);
nand U1165 (N_1165,N_24,N_484);
or U1166 (N_1166,N_459,N_681);
nand U1167 (N_1167,N_351,N_601);
and U1168 (N_1168,N_159,N_111);
nor U1169 (N_1169,N_776,N_437);
xnor U1170 (N_1170,N_938,N_887);
and U1171 (N_1171,N_103,N_206);
xnor U1172 (N_1172,N_640,N_14);
or U1173 (N_1173,N_842,N_259);
xor U1174 (N_1174,N_900,N_897);
and U1175 (N_1175,N_190,N_599);
and U1176 (N_1176,N_708,N_335);
nor U1177 (N_1177,N_669,N_516);
nor U1178 (N_1178,N_391,N_320);
xor U1179 (N_1179,N_226,N_96);
nand U1180 (N_1180,N_840,N_80);
xnor U1181 (N_1181,N_128,N_350);
nand U1182 (N_1182,N_23,N_851);
nand U1183 (N_1183,N_983,N_68);
nor U1184 (N_1184,N_629,N_173);
nand U1185 (N_1185,N_157,N_800);
or U1186 (N_1186,N_970,N_444);
nor U1187 (N_1187,N_804,N_60);
nor U1188 (N_1188,N_586,N_142);
xnor U1189 (N_1189,N_94,N_945);
nand U1190 (N_1190,N_263,N_195);
or U1191 (N_1191,N_981,N_10);
and U1192 (N_1192,N_406,N_578);
nor U1193 (N_1193,N_835,N_207);
nor U1194 (N_1194,N_202,N_92);
or U1195 (N_1195,N_342,N_469);
nor U1196 (N_1196,N_726,N_959);
nor U1197 (N_1197,N_990,N_625);
xnor U1198 (N_1198,N_736,N_913);
or U1199 (N_1199,N_176,N_709);
xor U1200 (N_1200,N_376,N_413);
nand U1201 (N_1201,N_559,N_967);
or U1202 (N_1202,N_55,N_569);
xnor U1203 (N_1203,N_702,N_180);
and U1204 (N_1204,N_290,N_951);
nor U1205 (N_1205,N_241,N_806);
nor U1206 (N_1206,N_154,N_871);
nand U1207 (N_1207,N_267,N_0);
nor U1208 (N_1208,N_141,N_993);
and U1209 (N_1209,N_31,N_2);
xor U1210 (N_1210,N_491,N_934);
xor U1211 (N_1211,N_753,N_216);
nor U1212 (N_1212,N_819,N_543);
xnor U1213 (N_1213,N_598,N_558);
nor U1214 (N_1214,N_160,N_158);
or U1215 (N_1215,N_235,N_855);
or U1216 (N_1216,N_499,N_902);
nor U1217 (N_1217,N_953,N_980);
nand U1218 (N_1218,N_430,N_679);
and U1219 (N_1219,N_910,N_606);
xor U1220 (N_1220,N_614,N_921);
and U1221 (N_1221,N_496,N_208);
and U1222 (N_1222,N_368,N_43);
or U1223 (N_1223,N_432,N_883);
nand U1224 (N_1224,N_563,N_770);
or U1225 (N_1225,N_700,N_188);
and U1226 (N_1226,N_231,N_264);
and U1227 (N_1227,N_927,N_831);
and U1228 (N_1228,N_234,N_843);
xnor U1229 (N_1229,N_608,N_357);
nor U1230 (N_1230,N_857,N_540);
nor U1231 (N_1231,N_223,N_904);
or U1232 (N_1232,N_714,N_150);
nor U1233 (N_1233,N_870,N_480);
xor U1234 (N_1234,N_306,N_184);
xnor U1235 (N_1235,N_509,N_508);
nor U1236 (N_1236,N_899,N_824);
or U1237 (N_1237,N_63,N_696);
or U1238 (N_1238,N_725,N_54);
nand U1239 (N_1239,N_88,N_155);
xor U1240 (N_1240,N_746,N_192);
and U1241 (N_1241,N_810,N_633);
nand U1242 (N_1242,N_821,N_973);
nand U1243 (N_1243,N_114,N_59);
nand U1244 (N_1244,N_388,N_799);
or U1245 (N_1245,N_439,N_332);
nor U1246 (N_1246,N_698,N_991);
nor U1247 (N_1247,N_183,N_724);
and U1248 (N_1248,N_803,N_925);
nor U1249 (N_1249,N_886,N_802);
xnor U1250 (N_1250,N_396,N_472);
nor U1251 (N_1251,N_632,N_118);
and U1252 (N_1252,N_106,N_722);
xor U1253 (N_1253,N_519,N_236);
nor U1254 (N_1254,N_737,N_133);
and U1255 (N_1255,N_968,N_270);
and U1256 (N_1256,N_495,N_265);
xor U1257 (N_1257,N_273,N_637);
nand U1258 (N_1258,N_171,N_940);
nand U1259 (N_1259,N_84,N_8);
xor U1260 (N_1260,N_292,N_143);
or U1261 (N_1261,N_149,N_452);
and U1262 (N_1262,N_607,N_237);
nand U1263 (N_1263,N_954,N_591);
and U1264 (N_1264,N_500,N_260);
nand U1265 (N_1265,N_91,N_574);
and U1266 (N_1266,N_820,N_793);
xor U1267 (N_1267,N_796,N_866);
nor U1268 (N_1268,N_217,N_573);
nand U1269 (N_1269,N_7,N_937);
nor U1270 (N_1270,N_277,N_248);
or U1271 (N_1271,N_409,N_319);
nor U1272 (N_1272,N_35,N_780);
xnor U1273 (N_1273,N_735,N_345);
nand U1274 (N_1274,N_661,N_611);
nor U1275 (N_1275,N_424,N_445);
nor U1276 (N_1276,N_807,N_784);
nand U1277 (N_1277,N_303,N_287);
and U1278 (N_1278,N_462,N_798);
nand U1279 (N_1279,N_134,N_322);
nor U1280 (N_1280,N_151,N_39);
nand U1281 (N_1281,N_908,N_211);
nor U1282 (N_1282,N_225,N_756);
or U1283 (N_1283,N_3,N_467);
nor U1284 (N_1284,N_903,N_727);
or U1285 (N_1285,N_513,N_65);
and U1286 (N_1286,N_436,N_498);
and U1287 (N_1287,N_572,N_415);
xor U1288 (N_1288,N_685,N_401);
nand U1289 (N_1289,N_944,N_381);
xnor U1290 (N_1290,N_486,N_169);
nand U1291 (N_1291,N_369,N_25);
nand U1292 (N_1292,N_626,N_553);
nand U1293 (N_1293,N_946,N_124);
xor U1294 (N_1294,N_330,N_665);
or U1295 (N_1295,N_911,N_16);
or U1296 (N_1296,N_296,N_957);
xor U1297 (N_1297,N_222,N_966);
and U1298 (N_1298,N_90,N_1);
nand U1299 (N_1299,N_19,N_773);
nor U1300 (N_1300,N_919,N_164);
nand U1301 (N_1301,N_671,N_152);
nor U1302 (N_1302,N_123,N_177);
nand U1303 (N_1303,N_505,N_958);
nor U1304 (N_1304,N_860,N_249);
nand U1305 (N_1305,N_845,N_538);
nand U1306 (N_1306,N_895,N_431);
nand U1307 (N_1307,N_761,N_268);
xnor U1308 (N_1308,N_38,N_893);
xor U1309 (N_1309,N_242,N_683);
xnor U1310 (N_1310,N_668,N_198);
xor U1311 (N_1311,N_370,N_829);
or U1312 (N_1312,N_140,N_730);
or U1313 (N_1313,N_880,N_274);
nor U1314 (N_1314,N_457,N_333);
or U1315 (N_1315,N_166,N_61);
and U1316 (N_1316,N_336,N_77);
or U1317 (N_1317,N_795,N_565);
nor U1318 (N_1318,N_186,N_507);
nor U1319 (N_1319,N_247,N_645);
and U1320 (N_1320,N_751,N_809);
or U1321 (N_1321,N_849,N_200);
xor U1322 (N_1322,N_240,N_135);
and U1323 (N_1323,N_882,N_986);
and U1324 (N_1324,N_533,N_347);
xor U1325 (N_1325,N_673,N_69);
xnor U1326 (N_1326,N_73,N_651);
or U1327 (N_1327,N_307,N_787);
xor U1328 (N_1328,N_402,N_132);
and U1329 (N_1329,N_971,N_564);
nand U1330 (N_1330,N_433,N_262);
or U1331 (N_1331,N_912,N_41);
xor U1332 (N_1332,N_961,N_219);
nor U1333 (N_1333,N_610,N_878);
xnor U1334 (N_1334,N_119,N_374);
or U1335 (N_1335,N_890,N_20);
and U1336 (N_1336,N_426,N_220);
or U1337 (N_1337,N_363,N_672);
or U1338 (N_1338,N_813,N_636);
or U1339 (N_1339,N_952,N_147);
nand U1340 (N_1340,N_535,N_718);
and U1341 (N_1341,N_926,N_950);
and U1342 (N_1342,N_534,N_383);
nor U1343 (N_1343,N_346,N_570);
or U1344 (N_1344,N_740,N_233);
nand U1345 (N_1345,N_40,N_66);
and U1346 (N_1346,N_837,N_139);
xor U1347 (N_1347,N_355,N_354);
nor U1348 (N_1348,N_101,N_11);
nand U1349 (N_1349,N_487,N_302);
or U1350 (N_1350,N_261,N_489);
and U1351 (N_1351,N_504,N_846);
nand U1352 (N_1352,N_515,N_790);
or U1353 (N_1353,N_972,N_755);
nand U1354 (N_1354,N_481,N_466);
and U1355 (N_1355,N_295,N_832);
and U1356 (N_1356,N_380,N_861);
nor U1357 (N_1357,N_518,N_501);
and U1358 (N_1358,N_742,N_266);
or U1359 (N_1359,N_547,N_224);
or U1360 (N_1360,N_32,N_653);
nand U1361 (N_1361,N_531,N_768);
nand U1362 (N_1362,N_996,N_788);
and U1363 (N_1363,N_131,N_674);
nand U1364 (N_1364,N_781,N_930);
nand U1365 (N_1365,N_448,N_122);
xnor U1366 (N_1366,N_594,N_739);
nor U1367 (N_1367,N_690,N_600);
and U1368 (N_1368,N_390,N_4);
or U1369 (N_1369,N_209,N_556);
xnor U1370 (N_1370,N_667,N_965);
xnor U1371 (N_1371,N_552,N_885);
nand U1372 (N_1372,N_95,N_161);
nor U1373 (N_1373,N_397,N_9);
xor U1374 (N_1374,N_148,N_471);
or U1375 (N_1375,N_759,N_71);
xor U1376 (N_1376,N_828,N_227);
nor U1377 (N_1377,N_635,N_447);
nor U1378 (N_1378,N_456,N_772);
and U1379 (N_1379,N_962,N_826);
and U1380 (N_1380,N_941,N_399);
or U1381 (N_1381,N_156,N_609);
nor U1382 (N_1382,N_102,N_52);
xor U1383 (N_1383,N_271,N_659);
or U1384 (N_1384,N_693,N_213);
nor U1385 (N_1385,N_658,N_282);
xnor U1386 (N_1386,N_109,N_618);
xor U1387 (N_1387,N_584,N_838);
nand U1388 (N_1388,N_324,N_305);
nor U1389 (N_1389,N_907,N_353);
or U1390 (N_1390,N_470,N_852);
nor U1391 (N_1391,N_738,N_64);
and U1392 (N_1392,N_298,N_997);
nand U1393 (N_1393,N_605,N_771);
and U1394 (N_1394,N_337,N_748);
or U1395 (N_1395,N_239,N_126);
nor U1396 (N_1396,N_524,N_823);
nand U1397 (N_1397,N_654,N_475);
and U1398 (N_1398,N_294,N_987);
or U1399 (N_1399,N_434,N_850);
nand U1400 (N_1400,N_719,N_482);
nand U1401 (N_1401,N_689,N_705);
nor U1402 (N_1402,N_947,N_985);
nand U1403 (N_1403,N_655,N_676);
and U1404 (N_1404,N_232,N_630);
or U1405 (N_1405,N_76,N_704);
xnor U1406 (N_1406,N_894,N_549);
xor U1407 (N_1407,N_638,N_943);
and U1408 (N_1408,N_794,N_631);
xor U1409 (N_1409,N_137,N_701);
nor U1410 (N_1410,N_189,N_747);
or U1411 (N_1411,N_301,N_105);
xnor U1412 (N_1412,N_288,N_873);
nand U1413 (N_1413,N_817,N_115);
nand U1414 (N_1414,N_87,N_522);
nand U1415 (N_1415,N_112,N_914);
and U1416 (N_1416,N_93,N_127);
nor U1417 (N_1417,N_341,N_928);
and U1418 (N_1418,N_53,N_620);
nand U1419 (N_1419,N_797,N_710);
nand U1420 (N_1420,N_26,N_872);
or U1421 (N_1421,N_801,N_853);
xor U1422 (N_1422,N_78,N_460);
and U1423 (N_1423,N_769,N_812);
and U1424 (N_1424,N_5,N_859);
or U1425 (N_1425,N_931,N_562);
nor U1426 (N_1426,N_199,N_27);
or U1427 (N_1427,N_539,N_419);
and U1428 (N_1428,N_45,N_575);
nand U1429 (N_1429,N_308,N_364);
or U1430 (N_1430,N_675,N_113);
and U1431 (N_1431,N_789,N_28);
nor U1432 (N_1432,N_699,N_583);
and U1433 (N_1433,N_830,N_975);
nor U1434 (N_1434,N_936,N_716);
xnor U1435 (N_1435,N_877,N_656);
xnor U1436 (N_1436,N_924,N_545);
xor U1437 (N_1437,N_643,N_862);
nand U1438 (N_1438,N_314,N_321);
or U1439 (N_1439,N_949,N_352);
xor U1440 (N_1440,N_731,N_316);
xnor U1441 (N_1441,N_257,N_385);
xnor U1442 (N_1442,N_929,N_848);
xor U1443 (N_1443,N_238,N_670);
xor U1444 (N_1444,N_170,N_512);
or U1445 (N_1445,N_616,N_523);
xor U1446 (N_1446,N_858,N_652);
nand U1447 (N_1447,N_827,N_289);
nor U1448 (N_1448,N_650,N_942);
nand U1449 (N_1449,N_458,N_982);
and U1450 (N_1450,N_67,N_712);
xor U1451 (N_1451,N_764,N_854);
or U1452 (N_1452,N_567,N_98);
and U1453 (N_1453,N_44,N_839);
nor U1454 (N_1454,N_687,N_205);
xnor U1455 (N_1455,N_193,N_461);
nor U1456 (N_1456,N_786,N_464);
nand U1457 (N_1457,N_395,N_502);
nand U1458 (N_1458,N_865,N_478);
or U1459 (N_1459,N_317,N_367);
or U1460 (N_1460,N_617,N_691);
and U1461 (N_1461,N_48,N_577);
nand U1462 (N_1462,N_889,N_763);
nand U1463 (N_1463,N_449,N_520);
nor U1464 (N_1464,N_490,N_356);
xnor U1465 (N_1465,N_723,N_37);
nor U1466 (N_1466,N_969,N_362);
nand U1467 (N_1467,N_17,N_644);
and U1468 (N_1468,N_939,N_453);
xnor U1469 (N_1469,N_663,N_551);
and U1470 (N_1470,N_657,N_86);
nor U1471 (N_1471,N_230,N_163);
nor U1472 (N_1472,N_976,N_493);
nand U1473 (N_1473,N_964,N_455);
nor U1474 (N_1474,N_587,N_29);
nand U1475 (N_1475,N_212,N_916);
nor U1476 (N_1476,N_686,N_326);
xor U1477 (N_1477,N_125,N_427);
xnor U1478 (N_1478,N_792,N_864);
xnor U1479 (N_1479,N_417,N_203);
nor U1480 (N_1480,N_554,N_503);
nand U1481 (N_1481,N_576,N_344);
nand U1482 (N_1482,N_348,N_783);
and U1483 (N_1483,N_680,N_99);
xor U1484 (N_1484,N_393,N_117);
nor U1485 (N_1485,N_387,N_136);
nand U1486 (N_1486,N_874,N_373);
nor U1487 (N_1487,N_463,N_275);
and U1488 (N_1488,N_49,N_624);
nor U1489 (N_1489,N_485,N_197);
or U1490 (N_1490,N_425,N_995);
and U1491 (N_1491,N_695,N_892);
xor U1492 (N_1492,N_627,N_588);
nor U1493 (N_1493,N_450,N_107);
nor U1494 (N_1494,N_185,N_741);
and U1495 (N_1495,N_70,N_297);
nand U1496 (N_1496,N_438,N_955);
or U1497 (N_1497,N_875,N_833);
nor U1498 (N_1498,N_782,N_416);
and U1499 (N_1499,N_706,N_492);
and U1500 (N_1500,N_63,N_686);
nand U1501 (N_1501,N_325,N_981);
and U1502 (N_1502,N_321,N_740);
nor U1503 (N_1503,N_202,N_221);
or U1504 (N_1504,N_536,N_661);
nor U1505 (N_1505,N_958,N_229);
and U1506 (N_1506,N_71,N_737);
or U1507 (N_1507,N_991,N_542);
and U1508 (N_1508,N_281,N_442);
or U1509 (N_1509,N_823,N_483);
or U1510 (N_1510,N_280,N_356);
or U1511 (N_1511,N_130,N_57);
and U1512 (N_1512,N_800,N_553);
xnor U1513 (N_1513,N_904,N_463);
and U1514 (N_1514,N_612,N_109);
or U1515 (N_1515,N_907,N_694);
xnor U1516 (N_1516,N_781,N_692);
or U1517 (N_1517,N_479,N_764);
xnor U1518 (N_1518,N_163,N_158);
and U1519 (N_1519,N_318,N_236);
or U1520 (N_1520,N_763,N_341);
nor U1521 (N_1521,N_49,N_220);
nor U1522 (N_1522,N_276,N_25);
and U1523 (N_1523,N_803,N_970);
or U1524 (N_1524,N_616,N_237);
or U1525 (N_1525,N_53,N_41);
nor U1526 (N_1526,N_765,N_136);
or U1527 (N_1527,N_28,N_871);
xnor U1528 (N_1528,N_496,N_418);
or U1529 (N_1529,N_366,N_558);
and U1530 (N_1530,N_0,N_15);
nor U1531 (N_1531,N_802,N_628);
and U1532 (N_1532,N_751,N_299);
and U1533 (N_1533,N_631,N_985);
and U1534 (N_1534,N_707,N_434);
nand U1535 (N_1535,N_298,N_693);
nand U1536 (N_1536,N_807,N_791);
nor U1537 (N_1537,N_716,N_853);
nand U1538 (N_1538,N_309,N_6);
and U1539 (N_1539,N_536,N_514);
nor U1540 (N_1540,N_143,N_328);
xor U1541 (N_1541,N_519,N_112);
and U1542 (N_1542,N_61,N_489);
or U1543 (N_1543,N_404,N_620);
xor U1544 (N_1544,N_325,N_46);
nand U1545 (N_1545,N_90,N_644);
or U1546 (N_1546,N_400,N_989);
or U1547 (N_1547,N_187,N_723);
nand U1548 (N_1548,N_318,N_577);
xnor U1549 (N_1549,N_283,N_924);
or U1550 (N_1550,N_346,N_402);
xnor U1551 (N_1551,N_255,N_24);
nor U1552 (N_1552,N_14,N_919);
and U1553 (N_1553,N_884,N_397);
or U1554 (N_1554,N_657,N_88);
and U1555 (N_1555,N_844,N_304);
nor U1556 (N_1556,N_887,N_997);
nor U1557 (N_1557,N_702,N_280);
xnor U1558 (N_1558,N_302,N_692);
xnor U1559 (N_1559,N_357,N_363);
xnor U1560 (N_1560,N_55,N_25);
or U1561 (N_1561,N_358,N_828);
and U1562 (N_1562,N_621,N_568);
nor U1563 (N_1563,N_10,N_176);
or U1564 (N_1564,N_906,N_967);
or U1565 (N_1565,N_793,N_463);
and U1566 (N_1566,N_465,N_879);
nor U1567 (N_1567,N_778,N_187);
and U1568 (N_1568,N_508,N_933);
nand U1569 (N_1569,N_657,N_442);
and U1570 (N_1570,N_222,N_608);
or U1571 (N_1571,N_90,N_284);
and U1572 (N_1572,N_761,N_333);
nand U1573 (N_1573,N_248,N_308);
nor U1574 (N_1574,N_536,N_791);
and U1575 (N_1575,N_648,N_404);
or U1576 (N_1576,N_654,N_344);
nor U1577 (N_1577,N_479,N_210);
nor U1578 (N_1578,N_557,N_838);
nor U1579 (N_1579,N_622,N_110);
nand U1580 (N_1580,N_800,N_612);
and U1581 (N_1581,N_319,N_189);
xnor U1582 (N_1582,N_178,N_168);
nand U1583 (N_1583,N_19,N_113);
nor U1584 (N_1584,N_984,N_278);
or U1585 (N_1585,N_950,N_814);
nand U1586 (N_1586,N_422,N_533);
nor U1587 (N_1587,N_650,N_719);
nor U1588 (N_1588,N_558,N_611);
or U1589 (N_1589,N_724,N_477);
nor U1590 (N_1590,N_248,N_226);
and U1591 (N_1591,N_495,N_42);
nor U1592 (N_1592,N_584,N_148);
nor U1593 (N_1593,N_863,N_368);
xnor U1594 (N_1594,N_118,N_856);
nand U1595 (N_1595,N_21,N_197);
xnor U1596 (N_1596,N_825,N_892);
and U1597 (N_1597,N_899,N_948);
nor U1598 (N_1598,N_42,N_823);
and U1599 (N_1599,N_131,N_928);
xor U1600 (N_1600,N_478,N_517);
or U1601 (N_1601,N_328,N_202);
or U1602 (N_1602,N_640,N_58);
nor U1603 (N_1603,N_165,N_769);
nand U1604 (N_1604,N_209,N_575);
nand U1605 (N_1605,N_748,N_562);
nand U1606 (N_1606,N_76,N_709);
or U1607 (N_1607,N_970,N_228);
xnor U1608 (N_1608,N_920,N_800);
and U1609 (N_1609,N_122,N_487);
or U1610 (N_1610,N_120,N_480);
or U1611 (N_1611,N_822,N_35);
nor U1612 (N_1612,N_918,N_834);
or U1613 (N_1613,N_239,N_798);
nor U1614 (N_1614,N_13,N_250);
nand U1615 (N_1615,N_467,N_327);
and U1616 (N_1616,N_722,N_864);
nor U1617 (N_1617,N_88,N_668);
and U1618 (N_1618,N_786,N_291);
nand U1619 (N_1619,N_73,N_333);
and U1620 (N_1620,N_403,N_210);
and U1621 (N_1621,N_537,N_152);
xnor U1622 (N_1622,N_355,N_887);
or U1623 (N_1623,N_386,N_330);
nor U1624 (N_1624,N_895,N_40);
and U1625 (N_1625,N_438,N_186);
xnor U1626 (N_1626,N_803,N_24);
and U1627 (N_1627,N_377,N_97);
or U1628 (N_1628,N_356,N_289);
and U1629 (N_1629,N_161,N_657);
xnor U1630 (N_1630,N_909,N_345);
or U1631 (N_1631,N_695,N_933);
xnor U1632 (N_1632,N_487,N_614);
or U1633 (N_1633,N_775,N_207);
nor U1634 (N_1634,N_295,N_430);
or U1635 (N_1635,N_401,N_74);
nor U1636 (N_1636,N_597,N_355);
or U1637 (N_1637,N_515,N_433);
nand U1638 (N_1638,N_164,N_174);
xor U1639 (N_1639,N_225,N_759);
nand U1640 (N_1640,N_379,N_913);
nor U1641 (N_1641,N_735,N_430);
nor U1642 (N_1642,N_750,N_0);
xor U1643 (N_1643,N_75,N_438);
nand U1644 (N_1644,N_750,N_682);
nand U1645 (N_1645,N_674,N_245);
nor U1646 (N_1646,N_299,N_771);
nor U1647 (N_1647,N_853,N_840);
xnor U1648 (N_1648,N_117,N_984);
and U1649 (N_1649,N_115,N_902);
nor U1650 (N_1650,N_529,N_603);
xnor U1651 (N_1651,N_413,N_20);
or U1652 (N_1652,N_486,N_416);
and U1653 (N_1653,N_96,N_206);
xor U1654 (N_1654,N_515,N_731);
or U1655 (N_1655,N_675,N_300);
xnor U1656 (N_1656,N_440,N_833);
or U1657 (N_1657,N_519,N_782);
nor U1658 (N_1658,N_941,N_432);
xor U1659 (N_1659,N_12,N_891);
nand U1660 (N_1660,N_403,N_388);
nor U1661 (N_1661,N_664,N_852);
xnor U1662 (N_1662,N_764,N_798);
nand U1663 (N_1663,N_497,N_875);
nand U1664 (N_1664,N_199,N_321);
nor U1665 (N_1665,N_581,N_838);
nor U1666 (N_1666,N_959,N_93);
nand U1667 (N_1667,N_926,N_261);
nor U1668 (N_1668,N_71,N_828);
nand U1669 (N_1669,N_758,N_621);
nand U1670 (N_1670,N_237,N_671);
or U1671 (N_1671,N_721,N_955);
xnor U1672 (N_1672,N_53,N_448);
xnor U1673 (N_1673,N_466,N_674);
or U1674 (N_1674,N_370,N_971);
xnor U1675 (N_1675,N_749,N_322);
and U1676 (N_1676,N_936,N_822);
and U1677 (N_1677,N_251,N_230);
nor U1678 (N_1678,N_976,N_622);
xnor U1679 (N_1679,N_67,N_106);
and U1680 (N_1680,N_711,N_412);
nor U1681 (N_1681,N_550,N_675);
xnor U1682 (N_1682,N_26,N_202);
and U1683 (N_1683,N_439,N_378);
and U1684 (N_1684,N_369,N_614);
or U1685 (N_1685,N_76,N_114);
xor U1686 (N_1686,N_739,N_323);
nor U1687 (N_1687,N_552,N_429);
nand U1688 (N_1688,N_911,N_799);
or U1689 (N_1689,N_920,N_496);
or U1690 (N_1690,N_985,N_730);
and U1691 (N_1691,N_706,N_998);
xor U1692 (N_1692,N_419,N_160);
or U1693 (N_1693,N_704,N_508);
xor U1694 (N_1694,N_332,N_653);
and U1695 (N_1695,N_188,N_497);
nand U1696 (N_1696,N_397,N_112);
and U1697 (N_1697,N_725,N_29);
nand U1698 (N_1698,N_703,N_338);
or U1699 (N_1699,N_952,N_575);
or U1700 (N_1700,N_864,N_353);
xnor U1701 (N_1701,N_767,N_373);
nor U1702 (N_1702,N_404,N_997);
or U1703 (N_1703,N_900,N_842);
nor U1704 (N_1704,N_890,N_492);
nor U1705 (N_1705,N_130,N_81);
nor U1706 (N_1706,N_440,N_324);
nor U1707 (N_1707,N_471,N_943);
nor U1708 (N_1708,N_117,N_932);
and U1709 (N_1709,N_905,N_700);
xor U1710 (N_1710,N_164,N_459);
nor U1711 (N_1711,N_570,N_908);
and U1712 (N_1712,N_844,N_605);
nand U1713 (N_1713,N_280,N_447);
nand U1714 (N_1714,N_669,N_12);
or U1715 (N_1715,N_746,N_779);
and U1716 (N_1716,N_63,N_268);
nor U1717 (N_1717,N_710,N_940);
and U1718 (N_1718,N_519,N_579);
nor U1719 (N_1719,N_975,N_494);
nor U1720 (N_1720,N_813,N_320);
and U1721 (N_1721,N_579,N_11);
and U1722 (N_1722,N_691,N_853);
xnor U1723 (N_1723,N_2,N_760);
and U1724 (N_1724,N_161,N_404);
xor U1725 (N_1725,N_783,N_62);
xnor U1726 (N_1726,N_723,N_207);
xor U1727 (N_1727,N_47,N_873);
and U1728 (N_1728,N_761,N_654);
or U1729 (N_1729,N_122,N_641);
and U1730 (N_1730,N_68,N_998);
and U1731 (N_1731,N_597,N_498);
nor U1732 (N_1732,N_212,N_328);
nor U1733 (N_1733,N_284,N_721);
nand U1734 (N_1734,N_174,N_954);
and U1735 (N_1735,N_987,N_284);
nand U1736 (N_1736,N_444,N_317);
xor U1737 (N_1737,N_345,N_131);
or U1738 (N_1738,N_202,N_429);
and U1739 (N_1739,N_683,N_295);
xor U1740 (N_1740,N_476,N_566);
or U1741 (N_1741,N_724,N_23);
nor U1742 (N_1742,N_92,N_430);
or U1743 (N_1743,N_123,N_601);
or U1744 (N_1744,N_412,N_475);
and U1745 (N_1745,N_639,N_771);
and U1746 (N_1746,N_895,N_576);
or U1747 (N_1747,N_965,N_984);
or U1748 (N_1748,N_915,N_386);
nor U1749 (N_1749,N_425,N_493);
and U1750 (N_1750,N_341,N_997);
nor U1751 (N_1751,N_26,N_268);
nand U1752 (N_1752,N_849,N_855);
xnor U1753 (N_1753,N_557,N_44);
nor U1754 (N_1754,N_647,N_622);
or U1755 (N_1755,N_952,N_185);
nor U1756 (N_1756,N_861,N_696);
xor U1757 (N_1757,N_165,N_513);
or U1758 (N_1758,N_917,N_403);
nand U1759 (N_1759,N_530,N_249);
xnor U1760 (N_1760,N_767,N_279);
xor U1761 (N_1761,N_621,N_438);
nor U1762 (N_1762,N_735,N_15);
xor U1763 (N_1763,N_348,N_999);
nand U1764 (N_1764,N_982,N_105);
or U1765 (N_1765,N_195,N_109);
and U1766 (N_1766,N_683,N_486);
nor U1767 (N_1767,N_25,N_151);
and U1768 (N_1768,N_440,N_447);
nand U1769 (N_1769,N_926,N_338);
or U1770 (N_1770,N_615,N_62);
xnor U1771 (N_1771,N_800,N_705);
nor U1772 (N_1772,N_962,N_452);
nand U1773 (N_1773,N_757,N_696);
or U1774 (N_1774,N_922,N_54);
or U1775 (N_1775,N_918,N_617);
xnor U1776 (N_1776,N_421,N_156);
nand U1777 (N_1777,N_310,N_401);
and U1778 (N_1778,N_344,N_533);
or U1779 (N_1779,N_585,N_617);
or U1780 (N_1780,N_387,N_438);
nor U1781 (N_1781,N_318,N_116);
or U1782 (N_1782,N_487,N_23);
and U1783 (N_1783,N_144,N_313);
nand U1784 (N_1784,N_609,N_663);
nor U1785 (N_1785,N_95,N_159);
or U1786 (N_1786,N_116,N_953);
xnor U1787 (N_1787,N_488,N_737);
and U1788 (N_1788,N_494,N_824);
or U1789 (N_1789,N_24,N_893);
and U1790 (N_1790,N_252,N_363);
or U1791 (N_1791,N_546,N_405);
xnor U1792 (N_1792,N_822,N_142);
nand U1793 (N_1793,N_529,N_314);
or U1794 (N_1794,N_810,N_981);
nand U1795 (N_1795,N_900,N_673);
and U1796 (N_1796,N_319,N_304);
and U1797 (N_1797,N_670,N_892);
nand U1798 (N_1798,N_943,N_193);
nor U1799 (N_1799,N_122,N_259);
nand U1800 (N_1800,N_817,N_70);
nand U1801 (N_1801,N_263,N_748);
nand U1802 (N_1802,N_945,N_194);
xnor U1803 (N_1803,N_813,N_187);
nor U1804 (N_1804,N_596,N_182);
and U1805 (N_1805,N_125,N_677);
and U1806 (N_1806,N_646,N_917);
and U1807 (N_1807,N_502,N_334);
or U1808 (N_1808,N_228,N_475);
nand U1809 (N_1809,N_714,N_447);
and U1810 (N_1810,N_476,N_998);
nand U1811 (N_1811,N_930,N_799);
nand U1812 (N_1812,N_233,N_513);
or U1813 (N_1813,N_435,N_268);
or U1814 (N_1814,N_218,N_772);
xnor U1815 (N_1815,N_670,N_833);
or U1816 (N_1816,N_906,N_946);
xnor U1817 (N_1817,N_563,N_521);
or U1818 (N_1818,N_738,N_452);
xnor U1819 (N_1819,N_186,N_671);
nand U1820 (N_1820,N_723,N_118);
xnor U1821 (N_1821,N_541,N_38);
nand U1822 (N_1822,N_608,N_663);
nand U1823 (N_1823,N_888,N_760);
xor U1824 (N_1824,N_899,N_364);
and U1825 (N_1825,N_157,N_223);
and U1826 (N_1826,N_96,N_35);
nand U1827 (N_1827,N_225,N_196);
and U1828 (N_1828,N_321,N_877);
nand U1829 (N_1829,N_359,N_948);
or U1830 (N_1830,N_843,N_338);
xnor U1831 (N_1831,N_312,N_797);
nor U1832 (N_1832,N_296,N_648);
nor U1833 (N_1833,N_138,N_862);
xor U1834 (N_1834,N_953,N_919);
and U1835 (N_1835,N_883,N_60);
or U1836 (N_1836,N_45,N_498);
or U1837 (N_1837,N_453,N_281);
nor U1838 (N_1838,N_269,N_582);
and U1839 (N_1839,N_547,N_972);
and U1840 (N_1840,N_154,N_636);
and U1841 (N_1841,N_64,N_393);
and U1842 (N_1842,N_755,N_531);
xor U1843 (N_1843,N_877,N_743);
and U1844 (N_1844,N_415,N_327);
nor U1845 (N_1845,N_390,N_133);
xnor U1846 (N_1846,N_566,N_965);
nor U1847 (N_1847,N_366,N_85);
nor U1848 (N_1848,N_228,N_443);
nand U1849 (N_1849,N_224,N_727);
or U1850 (N_1850,N_614,N_204);
xnor U1851 (N_1851,N_846,N_850);
or U1852 (N_1852,N_763,N_513);
xnor U1853 (N_1853,N_767,N_186);
xor U1854 (N_1854,N_522,N_260);
nor U1855 (N_1855,N_0,N_142);
nor U1856 (N_1856,N_824,N_613);
and U1857 (N_1857,N_439,N_989);
nor U1858 (N_1858,N_180,N_206);
or U1859 (N_1859,N_597,N_277);
and U1860 (N_1860,N_748,N_908);
and U1861 (N_1861,N_832,N_664);
nor U1862 (N_1862,N_887,N_53);
and U1863 (N_1863,N_688,N_3);
nand U1864 (N_1864,N_983,N_245);
nor U1865 (N_1865,N_833,N_925);
nor U1866 (N_1866,N_966,N_340);
and U1867 (N_1867,N_759,N_553);
nand U1868 (N_1868,N_674,N_400);
nand U1869 (N_1869,N_609,N_922);
xor U1870 (N_1870,N_609,N_153);
or U1871 (N_1871,N_600,N_542);
xnor U1872 (N_1872,N_707,N_529);
nand U1873 (N_1873,N_573,N_641);
or U1874 (N_1874,N_436,N_654);
or U1875 (N_1875,N_564,N_326);
nor U1876 (N_1876,N_983,N_850);
nor U1877 (N_1877,N_860,N_105);
and U1878 (N_1878,N_544,N_536);
nor U1879 (N_1879,N_384,N_974);
nor U1880 (N_1880,N_945,N_40);
and U1881 (N_1881,N_295,N_426);
and U1882 (N_1882,N_759,N_353);
or U1883 (N_1883,N_77,N_259);
nor U1884 (N_1884,N_852,N_98);
xnor U1885 (N_1885,N_847,N_12);
or U1886 (N_1886,N_24,N_692);
or U1887 (N_1887,N_973,N_138);
or U1888 (N_1888,N_946,N_766);
nor U1889 (N_1889,N_124,N_963);
xor U1890 (N_1890,N_837,N_65);
nand U1891 (N_1891,N_504,N_294);
and U1892 (N_1892,N_878,N_343);
nand U1893 (N_1893,N_342,N_145);
nand U1894 (N_1894,N_226,N_863);
or U1895 (N_1895,N_914,N_93);
xor U1896 (N_1896,N_569,N_118);
nand U1897 (N_1897,N_326,N_822);
and U1898 (N_1898,N_79,N_416);
nor U1899 (N_1899,N_966,N_832);
nand U1900 (N_1900,N_452,N_559);
or U1901 (N_1901,N_841,N_964);
nor U1902 (N_1902,N_191,N_465);
nor U1903 (N_1903,N_518,N_367);
xor U1904 (N_1904,N_519,N_938);
xnor U1905 (N_1905,N_459,N_988);
nor U1906 (N_1906,N_379,N_187);
and U1907 (N_1907,N_565,N_212);
xnor U1908 (N_1908,N_551,N_300);
xor U1909 (N_1909,N_64,N_809);
xnor U1910 (N_1910,N_375,N_237);
xnor U1911 (N_1911,N_998,N_460);
and U1912 (N_1912,N_42,N_763);
nor U1913 (N_1913,N_887,N_679);
and U1914 (N_1914,N_769,N_254);
nand U1915 (N_1915,N_297,N_236);
and U1916 (N_1916,N_630,N_7);
or U1917 (N_1917,N_98,N_500);
nand U1918 (N_1918,N_928,N_274);
nand U1919 (N_1919,N_122,N_663);
and U1920 (N_1920,N_266,N_640);
xor U1921 (N_1921,N_183,N_219);
and U1922 (N_1922,N_296,N_810);
nand U1923 (N_1923,N_136,N_428);
and U1924 (N_1924,N_81,N_354);
and U1925 (N_1925,N_752,N_551);
or U1926 (N_1926,N_768,N_626);
and U1927 (N_1927,N_187,N_556);
nor U1928 (N_1928,N_35,N_405);
or U1929 (N_1929,N_663,N_112);
and U1930 (N_1930,N_245,N_621);
or U1931 (N_1931,N_186,N_836);
or U1932 (N_1932,N_833,N_71);
and U1933 (N_1933,N_680,N_91);
xnor U1934 (N_1934,N_221,N_547);
nor U1935 (N_1935,N_347,N_701);
or U1936 (N_1936,N_104,N_230);
or U1937 (N_1937,N_436,N_752);
and U1938 (N_1938,N_624,N_949);
nor U1939 (N_1939,N_118,N_96);
xor U1940 (N_1940,N_443,N_557);
nor U1941 (N_1941,N_177,N_661);
and U1942 (N_1942,N_245,N_948);
nor U1943 (N_1943,N_376,N_998);
nor U1944 (N_1944,N_465,N_358);
nor U1945 (N_1945,N_667,N_357);
and U1946 (N_1946,N_851,N_173);
and U1947 (N_1947,N_253,N_383);
xor U1948 (N_1948,N_429,N_183);
xnor U1949 (N_1949,N_433,N_77);
and U1950 (N_1950,N_371,N_299);
xnor U1951 (N_1951,N_467,N_265);
nor U1952 (N_1952,N_938,N_952);
nor U1953 (N_1953,N_620,N_903);
and U1954 (N_1954,N_386,N_784);
or U1955 (N_1955,N_135,N_897);
and U1956 (N_1956,N_370,N_615);
nor U1957 (N_1957,N_659,N_449);
nand U1958 (N_1958,N_121,N_310);
nor U1959 (N_1959,N_523,N_207);
or U1960 (N_1960,N_730,N_474);
nand U1961 (N_1961,N_929,N_816);
or U1962 (N_1962,N_909,N_365);
xor U1963 (N_1963,N_953,N_431);
xnor U1964 (N_1964,N_955,N_401);
and U1965 (N_1965,N_695,N_369);
xor U1966 (N_1966,N_331,N_773);
xnor U1967 (N_1967,N_715,N_852);
nand U1968 (N_1968,N_582,N_979);
nor U1969 (N_1969,N_928,N_824);
nor U1970 (N_1970,N_96,N_370);
and U1971 (N_1971,N_883,N_81);
xor U1972 (N_1972,N_702,N_655);
nand U1973 (N_1973,N_312,N_987);
xnor U1974 (N_1974,N_6,N_399);
xnor U1975 (N_1975,N_948,N_988);
nand U1976 (N_1976,N_353,N_386);
and U1977 (N_1977,N_154,N_954);
xnor U1978 (N_1978,N_190,N_104);
or U1979 (N_1979,N_801,N_122);
and U1980 (N_1980,N_449,N_237);
or U1981 (N_1981,N_68,N_184);
xnor U1982 (N_1982,N_649,N_457);
or U1983 (N_1983,N_388,N_903);
nand U1984 (N_1984,N_196,N_492);
and U1985 (N_1985,N_263,N_92);
nor U1986 (N_1986,N_978,N_833);
or U1987 (N_1987,N_450,N_382);
or U1988 (N_1988,N_279,N_843);
nand U1989 (N_1989,N_490,N_423);
xnor U1990 (N_1990,N_918,N_342);
or U1991 (N_1991,N_199,N_330);
nand U1992 (N_1992,N_358,N_681);
xor U1993 (N_1993,N_829,N_348);
xor U1994 (N_1994,N_409,N_684);
nand U1995 (N_1995,N_432,N_675);
and U1996 (N_1996,N_497,N_604);
xnor U1997 (N_1997,N_588,N_536);
nor U1998 (N_1998,N_391,N_30);
and U1999 (N_1999,N_910,N_870);
or U2000 (N_2000,N_1946,N_1152);
nand U2001 (N_2001,N_1961,N_1101);
nand U2002 (N_2002,N_1667,N_1330);
and U2003 (N_2003,N_1451,N_1933);
xor U2004 (N_2004,N_1188,N_1621);
nand U2005 (N_2005,N_1637,N_1893);
and U2006 (N_2006,N_1497,N_1529);
or U2007 (N_2007,N_1392,N_1844);
or U2008 (N_2008,N_1161,N_1557);
or U2009 (N_2009,N_1234,N_1346);
xnor U2010 (N_2010,N_1638,N_1652);
nor U2011 (N_2011,N_1579,N_1075);
and U2012 (N_2012,N_1599,N_1746);
and U2013 (N_2013,N_1438,N_1105);
xnor U2014 (N_2014,N_1662,N_1831);
nor U2015 (N_2015,N_1617,N_1390);
xor U2016 (N_2016,N_1805,N_1891);
or U2017 (N_2017,N_1317,N_1928);
nor U2018 (N_2018,N_1711,N_1334);
nand U2019 (N_2019,N_1284,N_1097);
nor U2020 (N_2020,N_1580,N_1439);
and U2021 (N_2021,N_1357,N_1712);
and U2022 (N_2022,N_1403,N_1894);
and U2023 (N_2023,N_1643,N_1151);
and U2024 (N_2024,N_1709,N_1880);
or U2025 (N_2025,N_1061,N_1824);
xnor U2026 (N_2026,N_1764,N_1697);
or U2027 (N_2027,N_1190,N_1794);
nand U2028 (N_2028,N_1807,N_1852);
or U2029 (N_2029,N_1018,N_1810);
and U2030 (N_2030,N_1423,N_1375);
xnor U2031 (N_2031,N_1718,N_1400);
xnor U2032 (N_2032,N_1528,N_1552);
nor U2033 (N_2033,N_1565,N_1885);
xor U2034 (N_2034,N_1297,N_1822);
xnor U2035 (N_2035,N_1465,N_1149);
or U2036 (N_2036,N_1633,N_1780);
nand U2037 (N_2037,N_1993,N_1743);
xnor U2038 (N_2038,N_1548,N_1111);
xnor U2039 (N_2039,N_1737,N_1541);
nor U2040 (N_2040,N_1730,N_1685);
xor U2041 (N_2041,N_1502,N_1514);
or U2042 (N_2042,N_1892,N_1461);
nor U2043 (N_2043,N_1835,N_1607);
and U2044 (N_2044,N_1277,N_1522);
and U2045 (N_2045,N_1694,N_1021);
or U2046 (N_2046,N_1191,N_1542);
nor U2047 (N_2047,N_1750,N_1017);
or U2048 (N_2048,N_1653,N_1814);
or U2049 (N_2049,N_1544,N_1013);
xnor U2050 (N_2050,N_1648,N_1875);
xnor U2051 (N_2051,N_1996,N_1082);
nand U2052 (N_2052,N_1252,N_1449);
nor U2053 (N_2053,N_1328,N_1279);
xor U2054 (N_2054,N_1164,N_1581);
or U2055 (N_2055,N_1184,N_1121);
nor U2056 (N_2056,N_1060,N_1576);
xor U2057 (N_2057,N_1030,N_1942);
and U2058 (N_2058,N_1900,N_1918);
nor U2059 (N_2059,N_1925,N_1872);
or U2060 (N_2060,N_1287,N_1546);
nand U2061 (N_2061,N_1513,N_1717);
nor U2062 (N_2062,N_1235,N_1726);
or U2063 (N_2063,N_1517,N_1310);
and U2064 (N_2064,N_1250,N_1731);
and U2065 (N_2065,N_1887,N_1588);
nor U2066 (N_2066,N_1426,N_1904);
nand U2067 (N_2067,N_1763,N_1558);
nor U2068 (N_2068,N_1257,N_1293);
or U2069 (N_2069,N_1359,N_1367);
xnor U2070 (N_2070,N_1222,N_1406);
xor U2071 (N_2071,N_1864,N_1158);
or U2072 (N_2072,N_1424,N_1670);
nand U2073 (N_2073,N_1698,N_1004);
xor U2074 (N_2074,N_1742,N_1909);
nand U2075 (N_2075,N_1902,N_1353);
nand U2076 (N_2076,N_1285,N_1792);
or U2077 (N_2077,N_1476,N_1006);
nand U2078 (N_2078,N_1421,N_1689);
or U2079 (N_2079,N_1210,N_1138);
nand U2080 (N_2080,N_1821,N_1253);
nor U2081 (N_2081,N_1096,N_1981);
xor U2082 (N_2082,N_1759,N_1059);
xor U2083 (N_2083,N_1244,N_1321);
or U2084 (N_2084,N_1766,N_1224);
or U2085 (N_2085,N_1809,N_1153);
and U2086 (N_2086,N_1614,N_1057);
and U2087 (N_2087,N_1945,N_1562);
and U2088 (N_2088,N_1850,N_1231);
and U2089 (N_2089,N_1309,N_1755);
nand U2090 (N_2090,N_1987,N_1214);
xnor U2091 (N_2091,N_1964,N_1681);
xnor U2092 (N_2092,N_1606,N_1443);
xnor U2093 (N_2093,N_1563,N_1176);
xor U2094 (N_2094,N_1625,N_1770);
or U2095 (N_2095,N_1218,N_1071);
and U2096 (N_2096,N_1765,N_1070);
and U2097 (N_2097,N_1276,N_1661);
and U2098 (N_2098,N_1409,N_1209);
and U2099 (N_2099,N_1237,N_1063);
nand U2100 (N_2100,N_1773,N_1609);
nor U2101 (N_2101,N_1240,N_1073);
xnor U2102 (N_2102,N_1133,N_1586);
nor U2103 (N_2103,N_1725,N_1286);
nor U2104 (N_2104,N_1114,N_1254);
and U2105 (N_2105,N_1380,N_1705);
and U2106 (N_2106,N_1523,N_1693);
or U2107 (N_2107,N_1048,N_1274);
xor U2108 (N_2108,N_1530,N_1171);
nand U2109 (N_2109,N_1640,N_1910);
nand U2110 (N_2110,N_1148,N_1995);
xor U2111 (N_2111,N_1976,N_1147);
nand U2112 (N_2112,N_1116,N_1683);
nand U2113 (N_2113,N_1093,N_1129);
xnor U2114 (N_2114,N_1855,N_1704);
and U2115 (N_2115,N_1427,N_1815);
xor U2116 (N_2116,N_1157,N_1319);
xor U2117 (N_2117,N_1566,N_1054);
xor U2118 (N_2118,N_1354,N_1952);
xnor U2119 (N_2119,N_1913,N_1434);
nand U2120 (N_2120,N_1084,N_1929);
nand U2121 (N_2121,N_1388,N_1947);
nor U2122 (N_2122,N_1592,N_1659);
nand U2123 (N_2123,N_1457,N_1118);
or U2124 (N_2124,N_1641,N_1840);
nor U2125 (N_2125,N_1092,N_1790);
xor U2126 (N_2126,N_1932,N_1487);
and U2127 (N_2127,N_1469,N_1533);
xor U2128 (N_2128,N_1813,N_1361);
xor U2129 (N_2129,N_1965,N_1796);
xor U2130 (N_2130,N_1626,N_1798);
nand U2131 (N_2131,N_1376,N_1168);
or U2132 (N_2132,N_1520,N_1781);
nor U2133 (N_2133,N_1858,N_1401);
nand U2134 (N_2134,N_1554,N_1673);
nand U2135 (N_2135,N_1173,N_1561);
and U2136 (N_2136,N_1671,N_1587);
or U2137 (N_2137,N_1089,N_1037);
nor U2138 (N_2138,N_1348,N_1377);
and U2139 (N_2139,N_1674,N_1682);
xnor U2140 (N_2140,N_1959,N_1786);
nand U2141 (N_2141,N_1972,N_1608);
or U2142 (N_2142,N_1719,N_1771);
xnor U2143 (N_2143,N_1065,N_1124);
nor U2144 (N_2144,N_1255,N_1658);
or U2145 (N_2145,N_1839,N_1833);
xnor U2146 (N_2146,N_1734,N_1564);
and U2147 (N_2147,N_1365,N_1499);
nand U2148 (N_2148,N_1470,N_1373);
nand U2149 (N_2149,N_1249,N_1041);
and U2150 (N_2150,N_1326,N_1405);
or U2151 (N_2151,N_1829,N_1926);
or U2152 (N_2152,N_1701,N_1259);
and U2153 (N_2153,N_1559,N_1495);
or U2154 (N_2154,N_1484,N_1536);
xor U2155 (N_2155,N_1868,N_1318);
xor U2156 (N_2156,N_1733,N_1735);
xnor U2157 (N_2157,N_1068,N_1724);
nand U2158 (N_2158,N_1699,N_1721);
and U2159 (N_2159,N_1355,N_1602);
and U2160 (N_2160,N_1491,N_1990);
and U2161 (N_2161,N_1762,N_1686);
or U2162 (N_2162,N_1370,N_1342);
xnor U2163 (N_2163,N_1791,N_1690);
or U2164 (N_2164,N_1854,N_1534);
nand U2165 (N_2165,N_1509,N_1832);
or U2166 (N_2166,N_1185,N_1146);
nand U2167 (N_2167,N_1782,N_1199);
nand U2168 (N_2168,N_1615,N_1272);
xor U2169 (N_2169,N_1260,N_1710);
or U2170 (N_2170,N_1137,N_1162);
xnor U2171 (N_2171,N_1611,N_1998);
xor U2172 (N_2172,N_1897,N_1539);
or U2173 (N_2173,N_1211,N_1288);
xnor U2174 (N_2174,N_1347,N_1175);
xor U2175 (N_2175,N_1344,N_1033);
nand U2176 (N_2176,N_1371,N_1604);
or U2177 (N_2177,N_1631,N_1408);
nor U2178 (N_2178,N_1908,N_1448);
and U2179 (N_2179,N_1056,N_1582);
and U2180 (N_2180,N_1485,N_1494);
and U2181 (N_2181,N_1714,N_1402);
nor U2182 (N_2182,N_1019,N_1479);
xnor U2183 (N_2183,N_1825,N_1431);
and U2184 (N_2184,N_1795,N_1182);
or U2185 (N_2185,N_1507,N_1198);
nor U2186 (N_2186,N_1715,N_1757);
xnor U2187 (N_2187,N_1226,N_1776);
nand U2188 (N_2188,N_1876,N_1180);
nand U2189 (N_2189,N_1577,N_1512);
xor U2190 (N_2190,N_1200,N_1298);
nor U2191 (N_2191,N_1927,N_1657);
nand U2192 (N_2192,N_1094,N_1843);
nand U2193 (N_2193,N_1302,N_1706);
or U2194 (N_2194,N_1882,N_1139);
and U2195 (N_2195,N_1109,N_1220);
nand U2196 (N_2196,N_1315,N_1119);
nor U2197 (N_2197,N_1797,N_1383);
or U2198 (N_2198,N_1053,N_1740);
xor U2199 (N_2199,N_1258,N_1591);
nand U2200 (N_2200,N_1177,N_1187);
and U2201 (N_2201,N_1201,N_1369);
and U2202 (N_2202,N_1372,N_1213);
xor U2203 (N_2203,N_1335,N_1425);
nor U2204 (N_2204,N_1537,N_1958);
nor U2205 (N_2205,N_1859,N_1675);
and U2206 (N_2206,N_1266,N_1739);
nand U2207 (N_2207,N_1166,N_1189);
and U2208 (N_2208,N_1761,N_1091);
nor U2209 (N_2209,N_1988,N_1837);
nor U2210 (N_2210,N_1051,N_1160);
nand U2211 (N_2211,N_1378,N_1239);
or U2212 (N_2212,N_1610,N_1511);
or U2213 (N_2213,N_1853,N_1108);
nand U2214 (N_2214,N_1951,N_1613);
and U2215 (N_2215,N_1707,N_1280);
nand U2216 (N_2216,N_1247,N_1113);
xnor U2217 (N_2217,N_1263,N_1204);
xor U2218 (N_2218,N_1433,N_1275);
nand U2219 (N_2219,N_1768,N_1440);
nor U2220 (N_2220,N_1174,N_1087);
nand U2221 (N_2221,N_1273,N_1103);
or U2222 (N_2222,N_1603,N_1655);
or U2223 (N_2223,N_1282,N_1314);
nor U2224 (N_2224,N_1464,N_1047);
nand U2225 (N_2225,N_1979,N_1860);
xnor U2226 (N_2226,N_1192,N_1186);
or U2227 (N_2227,N_1281,N_1680);
and U2228 (N_2228,N_1816,N_1881);
and U2229 (N_2229,N_1154,N_1527);
or U2230 (N_2230,N_1635,N_1869);
nand U2231 (N_2231,N_1999,N_1943);
and U2232 (N_2232,N_1769,N_1804);
nand U2233 (N_2233,N_1519,N_1884);
or U2234 (N_2234,N_1538,N_1989);
xnor U2235 (N_2235,N_1008,N_1125);
xnor U2236 (N_2236,N_1473,N_1458);
nand U2237 (N_2237,N_1134,N_1994);
and U2238 (N_2238,N_1379,N_1117);
and U2239 (N_2239,N_1135,N_1622);
and U2240 (N_2240,N_1944,N_1877);
nor U2241 (N_2241,N_1915,N_1624);
xnor U2242 (N_2242,N_1787,N_1551);
nor U2243 (N_2243,N_1264,N_1269);
or U2244 (N_2244,N_1811,N_1352);
xnor U2245 (N_2245,N_1772,N_1744);
nor U2246 (N_2246,N_1144,N_1350);
xnor U2247 (N_2247,N_1395,N_1289);
nand U2248 (N_2248,N_1404,N_1165);
xor U2249 (N_2249,N_1919,N_1336);
xor U2250 (N_2250,N_1687,N_1150);
xor U2251 (N_2251,N_1301,N_1636);
nand U2252 (N_2252,N_1774,N_1903);
xor U2253 (N_2253,N_1356,N_1954);
and U2254 (N_2254,N_1749,N_1058);
nand U2255 (N_2255,N_1906,N_1141);
nor U2256 (N_2256,N_1574,N_1022);
and U2257 (N_2257,N_1142,N_1865);
and U2258 (N_2258,N_1050,N_1038);
xor U2259 (N_2259,N_1616,N_1846);
and U2260 (N_2260,N_1178,N_1741);
or U2261 (N_2261,N_1025,N_1598);
nand U2262 (N_2262,N_1665,N_1651);
nor U2263 (N_2263,N_1463,N_1430);
nor U2264 (N_2264,N_1453,N_1360);
or U2265 (N_2265,N_1696,N_1412);
nor U2266 (N_2266,N_1316,N_1072);
nand U2267 (N_2267,N_1327,N_1767);
xor U2268 (N_2268,N_1332,N_1901);
and U2269 (N_2269,N_1243,N_1306);
xor U2270 (N_2270,N_1027,N_1225);
nor U2271 (N_2271,N_1337,N_1496);
or U2272 (N_2272,N_1397,N_1874);
xnor U2273 (N_2273,N_1802,N_1459);
nor U2274 (N_2274,N_1801,N_1789);
or U2275 (N_2275,N_1248,N_1799);
xor U2276 (N_2276,N_1283,N_1555);
nand U2277 (N_2277,N_1890,N_1632);
and U2278 (N_2278,N_1589,N_1620);
xnor U2279 (N_2279,N_1779,N_1612);
xor U2280 (N_2280,N_1215,N_1110);
and U2281 (N_2281,N_1329,N_1120);
xnor U2282 (N_2282,N_1645,N_1106);
nand U2283 (N_2283,N_1074,N_1886);
and U2284 (N_2284,N_1384,N_1024);
and U2285 (N_2285,N_1196,N_1578);
or U2286 (N_2286,N_1203,N_1510);
xnor U2287 (N_2287,N_1963,N_1806);
or U2288 (N_2288,N_1472,N_1727);
xor U2289 (N_2289,N_1584,N_1679);
nor U2290 (N_2290,N_1723,N_1920);
nor U2291 (N_2291,N_1628,N_1062);
nand U2292 (N_2292,N_1754,N_1341);
and U2293 (N_2293,N_1020,N_1753);
nand U2294 (N_2294,N_1498,N_1011);
and U2295 (N_2295,N_1032,N_1212);
xor U2296 (N_2296,N_1545,N_1251);
nand U2297 (N_2297,N_1575,N_1691);
or U2298 (N_2298,N_1639,N_1623);
and U2299 (N_2299,N_1991,N_1569);
and U2300 (N_2300,N_1703,N_1842);
nand U2301 (N_2301,N_1678,N_1446);
nor U2302 (N_2302,N_1143,N_1123);
xnor U2303 (N_2303,N_1303,N_1834);
xor U2304 (N_2304,N_1418,N_1278);
nand U2305 (N_2305,N_1524,N_1381);
and U2306 (N_2306,N_1728,N_1219);
xor U2307 (N_2307,N_1104,N_1732);
and U2308 (N_2308,N_1629,N_1295);
and U2309 (N_2309,N_1970,N_1444);
nor U2310 (N_2310,N_1800,N_1553);
nand U2311 (N_2311,N_1081,N_1907);
and U2312 (N_2312,N_1879,N_1001);
and U2313 (N_2313,N_1031,N_1899);
nand U2314 (N_2314,N_1873,N_1937);
and U2315 (N_2315,N_1695,N_1107);
nor U2316 (N_2316,N_1593,N_1585);
nand U2317 (N_2317,N_1029,N_1916);
nor U2318 (N_2318,N_1971,N_1163);
and U2319 (N_2319,N_1098,N_1526);
xnor U2320 (N_2320,N_1012,N_1416);
nor U2321 (N_2321,N_1666,N_1304);
nand U2322 (N_2322,N_1751,N_1233);
and U2323 (N_2323,N_1100,N_1036);
xnor U2324 (N_2324,N_1265,N_1745);
or U2325 (N_2325,N_1331,N_1080);
nand U2326 (N_2326,N_1490,N_1847);
nand U2327 (N_2327,N_1155,N_1351);
nor U2328 (N_2328,N_1752,N_1034);
nor U2329 (N_2329,N_1818,N_1362);
nand U2330 (N_2330,N_1169,N_1663);
xor U2331 (N_2331,N_1594,N_1079);
xnor U2332 (N_2332,N_1290,N_1471);
nand U2333 (N_2333,N_1619,N_1760);
xor U2334 (N_2334,N_1992,N_1374);
nand U2335 (N_2335,N_1320,N_1819);
nor U2336 (N_2336,N_1324,N_1066);
nand U2337 (N_2337,N_1827,N_1195);
or U2338 (N_2338,N_1968,N_1040);
nor U2339 (N_2339,N_1338,N_1838);
nor U2340 (N_2340,N_1647,N_1863);
nor U2341 (N_2341,N_1009,N_1938);
nor U2342 (N_2342,N_1812,N_1525);
or U2343 (N_2343,N_1207,N_1261);
xnor U2344 (N_2344,N_1271,N_1478);
nand U2345 (N_2345,N_1078,N_1997);
nor U2346 (N_2346,N_1783,N_1436);
and U2347 (N_2347,N_1128,N_1016);
xor U2348 (N_2348,N_1702,N_1934);
or U2349 (N_2349,N_1560,N_1246);
xnor U2350 (N_2350,N_1966,N_1230);
nand U2351 (N_2351,N_1267,N_1748);
xor U2352 (N_2352,N_1700,N_1911);
and U2353 (N_2353,N_1387,N_1969);
nand U2354 (N_2354,N_1015,N_1851);
xor U2355 (N_2355,N_1339,N_1540);
xor U2356 (N_2356,N_1145,N_1181);
and U2357 (N_2357,N_1922,N_1975);
nor U2358 (N_2358,N_1849,N_1547);
nor U2359 (N_2359,N_1486,N_1956);
nor U2360 (N_2360,N_1193,N_1368);
or U2361 (N_2361,N_1462,N_1262);
nor U2362 (N_2362,N_1597,N_1568);
and U2363 (N_2363,N_1889,N_1898);
nor U2364 (N_2364,N_1441,N_1841);
and U2365 (N_2365,N_1333,N_1052);
xor U2366 (N_2366,N_1500,N_1823);
nor U2367 (N_2367,N_1924,N_1688);
or U2368 (N_2368,N_1127,N_1294);
nand U2369 (N_2369,N_1429,N_1206);
or U2370 (N_2370,N_1986,N_1456);
xor U2371 (N_2371,N_1242,N_1595);
and U2372 (N_2372,N_1729,N_1600);
nand U2373 (N_2373,N_1803,N_1194);
or U2374 (N_2374,N_1112,N_1323);
or U2375 (N_2375,N_1228,N_1758);
nor U2376 (N_2376,N_1217,N_1086);
and U2377 (N_2377,N_1828,N_1618);
and U2378 (N_2378,N_1935,N_1983);
nand U2379 (N_2379,N_1349,N_1516);
nand U2380 (N_2380,N_1345,N_1508);
xor U2381 (N_2381,N_1450,N_1720);
nor U2382 (N_2382,N_1049,N_1090);
or U2383 (N_2383,N_1311,N_1912);
nor U2384 (N_2384,N_1126,N_1982);
nor U2385 (N_2385,N_1002,N_1605);
xor U2386 (N_2386,N_1241,N_1867);
nor U2387 (N_2387,N_1503,N_1571);
nand U2388 (N_2388,N_1026,N_1046);
or U2389 (N_2389,N_1775,N_1895);
and U2390 (N_2390,N_1202,N_1115);
xnor U2391 (N_2391,N_1684,N_1300);
xor U2392 (N_2392,N_1504,N_1023);
nor U2393 (N_2393,N_1039,N_1883);
nor U2394 (N_2394,N_1590,N_1340);
or U2395 (N_2395,N_1393,N_1364);
xnor U2396 (N_2396,N_1205,N_1978);
xor U2397 (N_2397,N_1660,N_1820);
or U2398 (N_2398,N_1437,N_1256);
nand U2399 (N_2399,N_1949,N_1064);
and U2400 (N_2400,N_1567,N_1467);
and U2401 (N_2401,N_1389,N_1322);
nor U2402 (N_2402,N_1291,N_1905);
or U2403 (N_2403,N_1236,N_1848);
or U2404 (N_2404,N_1923,N_1941);
or U2405 (N_2405,N_1197,N_1010);
nand U2406 (N_2406,N_1646,N_1028);
xor U2407 (N_2407,N_1778,N_1043);
or U2408 (N_2408,N_1870,N_1917);
nand U2409 (N_2409,N_1232,N_1325);
xnor U2410 (N_2410,N_1466,N_1055);
or U2411 (N_2411,N_1099,N_1102);
nor U2412 (N_2412,N_1396,N_1422);
nand U2413 (N_2413,N_1268,N_1428);
nand U2414 (N_2414,N_1708,N_1414);
nand U2415 (N_2415,N_1692,N_1131);
nor U2416 (N_2416,N_1948,N_1003);
xnor U2417 (N_2417,N_1627,N_1878);
xnor U2418 (N_2418,N_1420,N_1493);
nand U2419 (N_2419,N_1543,N_1385);
or U2420 (N_2420,N_1394,N_1229);
nor U2421 (N_2421,N_1363,N_1676);
nand U2422 (N_2422,N_1417,N_1386);
or U2423 (N_2423,N_1045,N_1871);
xnor U2424 (N_2424,N_1977,N_1784);
xor U2425 (N_2425,N_1669,N_1296);
xnor U2426 (N_2426,N_1777,N_1305);
and U2427 (N_2427,N_1468,N_1452);
nor U2428 (N_2428,N_1532,N_1140);
xor U2429 (N_2429,N_1179,N_1270);
and U2430 (N_2430,N_1973,N_1088);
and U2431 (N_2431,N_1960,N_1159);
nand U2432 (N_2432,N_1664,N_1245);
or U2433 (N_2433,N_1644,N_1007);
nand U2434 (N_2434,N_1475,N_1014);
xor U2435 (N_2435,N_1411,N_1856);
xnor U2436 (N_2436,N_1649,N_1521);
xnor U2437 (N_2437,N_1005,N_1382);
and U2438 (N_2438,N_1817,N_1531);
or U2439 (N_2439,N_1672,N_1077);
xor U2440 (N_2440,N_1940,N_1857);
or U2441 (N_2441,N_1556,N_1985);
xnor U2442 (N_2442,N_1223,N_1447);
nand U2443 (N_2443,N_1967,N_1419);
or U2444 (N_2444,N_1221,N_1391);
or U2445 (N_2445,N_1454,N_1035);
or U2446 (N_2446,N_1313,N_1515);
nor U2447 (N_2447,N_1489,N_1984);
nand U2448 (N_2448,N_1914,N_1861);
nor U2449 (N_2449,N_1950,N_1980);
and U2450 (N_2450,N_1505,N_1442);
xor U2451 (N_2451,N_1866,N_1067);
nor U2452 (N_2452,N_1845,N_1445);
xor U2453 (N_2453,N_1634,N_1747);
nor U2454 (N_2454,N_1642,N_1930);
nor U2455 (N_2455,N_1896,N_1343);
nor U2456 (N_2456,N_1677,N_1122);
nand U2457 (N_2457,N_1410,N_1482);
or U2458 (N_2458,N_1830,N_1931);
and U2459 (N_2459,N_1518,N_1042);
nor U2460 (N_2460,N_1000,N_1738);
nor U2461 (N_2461,N_1312,N_1481);
and U2462 (N_2462,N_1483,N_1167);
xor U2463 (N_2463,N_1888,N_1474);
and U2464 (N_2464,N_1358,N_1535);
or U2465 (N_2465,N_1955,N_1953);
or U2466 (N_2466,N_1407,N_1366);
and U2467 (N_2467,N_1170,N_1974);
and U2468 (N_2468,N_1501,N_1630);
xor U2469 (N_2469,N_1583,N_1793);
and U2470 (N_2470,N_1808,N_1238);
xor U2471 (N_2471,N_1095,N_1399);
nand U2472 (N_2472,N_1785,N_1208);
nand U2473 (N_2473,N_1716,N_1957);
nor U2474 (N_2474,N_1432,N_1836);
and U2475 (N_2475,N_1435,N_1826);
and U2476 (N_2476,N_1722,N_1083);
nand U2477 (N_2477,N_1398,N_1570);
and U2478 (N_2478,N_1601,N_1460);
nand U2479 (N_2479,N_1921,N_1307);
and U2480 (N_2480,N_1939,N_1455);
or U2481 (N_2481,N_1650,N_1550);
or U2482 (N_2482,N_1573,N_1656);
and U2483 (N_2483,N_1044,N_1132);
xnor U2484 (N_2484,N_1488,N_1172);
nor U2485 (N_2485,N_1477,N_1183);
and U2486 (N_2486,N_1299,N_1572);
and U2487 (N_2487,N_1130,N_1936);
nor U2488 (N_2488,N_1069,N_1506);
nor U2489 (N_2489,N_1756,N_1415);
nand U2490 (N_2490,N_1136,N_1413);
nand U2491 (N_2491,N_1480,N_1713);
or U2492 (N_2492,N_1736,N_1788);
xor U2493 (N_2493,N_1668,N_1492);
nand U2494 (N_2494,N_1216,N_1227);
and U2495 (N_2495,N_1962,N_1308);
xor U2496 (N_2496,N_1156,N_1862);
nand U2497 (N_2497,N_1085,N_1549);
xnor U2498 (N_2498,N_1596,N_1654);
nor U2499 (N_2499,N_1076,N_1292);
or U2500 (N_2500,N_1171,N_1102);
xnor U2501 (N_2501,N_1179,N_1913);
nor U2502 (N_2502,N_1232,N_1799);
nand U2503 (N_2503,N_1732,N_1186);
nor U2504 (N_2504,N_1187,N_1047);
nor U2505 (N_2505,N_1957,N_1928);
or U2506 (N_2506,N_1798,N_1181);
and U2507 (N_2507,N_1031,N_1942);
nor U2508 (N_2508,N_1483,N_1158);
nand U2509 (N_2509,N_1533,N_1509);
and U2510 (N_2510,N_1071,N_1957);
and U2511 (N_2511,N_1261,N_1535);
and U2512 (N_2512,N_1157,N_1875);
xor U2513 (N_2513,N_1028,N_1055);
and U2514 (N_2514,N_1332,N_1846);
or U2515 (N_2515,N_1408,N_1982);
nor U2516 (N_2516,N_1453,N_1877);
and U2517 (N_2517,N_1129,N_1835);
and U2518 (N_2518,N_1294,N_1487);
nor U2519 (N_2519,N_1344,N_1709);
or U2520 (N_2520,N_1537,N_1661);
nor U2521 (N_2521,N_1934,N_1937);
nor U2522 (N_2522,N_1620,N_1760);
nor U2523 (N_2523,N_1215,N_1556);
or U2524 (N_2524,N_1104,N_1105);
or U2525 (N_2525,N_1618,N_1543);
nor U2526 (N_2526,N_1660,N_1807);
nor U2527 (N_2527,N_1589,N_1565);
and U2528 (N_2528,N_1117,N_1054);
nand U2529 (N_2529,N_1942,N_1215);
or U2530 (N_2530,N_1389,N_1978);
xnor U2531 (N_2531,N_1367,N_1943);
or U2532 (N_2532,N_1756,N_1472);
and U2533 (N_2533,N_1569,N_1105);
nor U2534 (N_2534,N_1745,N_1294);
or U2535 (N_2535,N_1184,N_1042);
xor U2536 (N_2536,N_1327,N_1799);
nor U2537 (N_2537,N_1620,N_1258);
nor U2538 (N_2538,N_1592,N_1562);
nor U2539 (N_2539,N_1498,N_1495);
or U2540 (N_2540,N_1203,N_1251);
and U2541 (N_2541,N_1269,N_1891);
xnor U2542 (N_2542,N_1137,N_1045);
nor U2543 (N_2543,N_1434,N_1603);
nor U2544 (N_2544,N_1467,N_1215);
or U2545 (N_2545,N_1849,N_1998);
nand U2546 (N_2546,N_1344,N_1587);
nand U2547 (N_2547,N_1762,N_1452);
or U2548 (N_2548,N_1606,N_1539);
xor U2549 (N_2549,N_1279,N_1587);
nor U2550 (N_2550,N_1670,N_1313);
nor U2551 (N_2551,N_1536,N_1688);
nand U2552 (N_2552,N_1073,N_1126);
xor U2553 (N_2553,N_1273,N_1027);
and U2554 (N_2554,N_1037,N_1791);
or U2555 (N_2555,N_1562,N_1570);
nor U2556 (N_2556,N_1132,N_1674);
and U2557 (N_2557,N_1976,N_1171);
nand U2558 (N_2558,N_1569,N_1711);
nor U2559 (N_2559,N_1210,N_1898);
or U2560 (N_2560,N_1007,N_1301);
nand U2561 (N_2561,N_1288,N_1355);
xnor U2562 (N_2562,N_1982,N_1501);
nand U2563 (N_2563,N_1657,N_1486);
or U2564 (N_2564,N_1605,N_1704);
or U2565 (N_2565,N_1959,N_1606);
nor U2566 (N_2566,N_1577,N_1625);
xnor U2567 (N_2567,N_1133,N_1109);
or U2568 (N_2568,N_1774,N_1513);
or U2569 (N_2569,N_1091,N_1489);
or U2570 (N_2570,N_1226,N_1122);
nand U2571 (N_2571,N_1375,N_1485);
or U2572 (N_2572,N_1682,N_1328);
or U2573 (N_2573,N_1119,N_1412);
nand U2574 (N_2574,N_1544,N_1251);
or U2575 (N_2575,N_1154,N_1476);
or U2576 (N_2576,N_1107,N_1275);
or U2577 (N_2577,N_1735,N_1912);
xor U2578 (N_2578,N_1339,N_1360);
nand U2579 (N_2579,N_1413,N_1399);
nor U2580 (N_2580,N_1307,N_1099);
nor U2581 (N_2581,N_1773,N_1399);
nor U2582 (N_2582,N_1056,N_1474);
or U2583 (N_2583,N_1203,N_1950);
nand U2584 (N_2584,N_1974,N_1999);
or U2585 (N_2585,N_1194,N_1744);
nand U2586 (N_2586,N_1325,N_1475);
and U2587 (N_2587,N_1989,N_1081);
or U2588 (N_2588,N_1243,N_1461);
nor U2589 (N_2589,N_1438,N_1550);
nand U2590 (N_2590,N_1798,N_1674);
xnor U2591 (N_2591,N_1673,N_1413);
nand U2592 (N_2592,N_1185,N_1623);
xor U2593 (N_2593,N_1757,N_1129);
nand U2594 (N_2594,N_1452,N_1330);
nand U2595 (N_2595,N_1025,N_1665);
nand U2596 (N_2596,N_1542,N_1106);
or U2597 (N_2597,N_1545,N_1188);
and U2598 (N_2598,N_1520,N_1763);
and U2599 (N_2599,N_1549,N_1976);
nor U2600 (N_2600,N_1905,N_1618);
and U2601 (N_2601,N_1514,N_1165);
and U2602 (N_2602,N_1305,N_1709);
or U2603 (N_2603,N_1461,N_1015);
nand U2604 (N_2604,N_1450,N_1749);
and U2605 (N_2605,N_1449,N_1142);
and U2606 (N_2606,N_1300,N_1750);
xnor U2607 (N_2607,N_1659,N_1841);
nor U2608 (N_2608,N_1170,N_1777);
xnor U2609 (N_2609,N_1041,N_1819);
or U2610 (N_2610,N_1235,N_1322);
nand U2611 (N_2611,N_1912,N_1360);
xnor U2612 (N_2612,N_1492,N_1931);
xnor U2613 (N_2613,N_1890,N_1788);
nor U2614 (N_2614,N_1703,N_1923);
and U2615 (N_2615,N_1599,N_1734);
and U2616 (N_2616,N_1384,N_1160);
nand U2617 (N_2617,N_1726,N_1203);
nand U2618 (N_2618,N_1958,N_1149);
nor U2619 (N_2619,N_1155,N_1105);
xor U2620 (N_2620,N_1292,N_1083);
and U2621 (N_2621,N_1898,N_1778);
nand U2622 (N_2622,N_1343,N_1419);
xnor U2623 (N_2623,N_1610,N_1897);
and U2624 (N_2624,N_1131,N_1137);
xnor U2625 (N_2625,N_1987,N_1905);
xnor U2626 (N_2626,N_1298,N_1763);
nor U2627 (N_2627,N_1889,N_1848);
or U2628 (N_2628,N_1346,N_1658);
nor U2629 (N_2629,N_1625,N_1696);
or U2630 (N_2630,N_1354,N_1695);
xor U2631 (N_2631,N_1525,N_1003);
xnor U2632 (N_2632,N_1152,N_1031);
or U2633 (N_2633,N_1013,N_1986);
and U2634 (N_2634,N_1705,N_1626);
or U2635 (N_2635,N_1029,N_1574);
xnor U2636 (N_2636,N_1092,N_1208);
nand U2637 (N_2637,N_1868,N_1535);
nand U2638 (N_2638,N_1069,N_1774);
and U2639 (N_2639,N_1115,N_1707);
or U2640 (N_2640,N_1511,N_1018);
xnor U2641 (N_2641,N_1321,N_1295);
xor U2642 (N_2642,N_1175,N_1290);
nand U2643 (N_2643,N_1660,N_1987);
nand U2644 (N_2644,N_1444,N_1673);
and U2645 (N_2645,N_1535,N_1767);
nand U2646 (N_2646,N_1474,N_1539);
xnor U2647 (N_2647,N_1690,N_1039);
or U2648 (N_2648,N_1391,N_1599);
nor U2649 (N_2649,N_1073,N_1928);
nand U2650 (N_2650,N_1109,N_1192);
nor U2651 (N_2651,N_1232,N_1345);
xor U2652 (N_2652,N_1585,N_1952);
nand U2653 (N_2653,N_1665,N_1159);
or U2654 (N_2654,N_1876,N_1940);
nand U2655 (N_2655,N_1620,N_1185);
nand U2656 (N_2656,N_1962,N_1671);
nand U2657 (N_2657,N_1612,N_1969);
xnor U2658 (N_2658,N_1289,N_1130);
nor U2659 (N_2659,N_1989,N_1721);
or U2660 (N_2660,N_1964,N_1666);
xnor U2661 (N_2661,N_1518,N_1096);
and U2662 (N_2662,N_1218,N_1250);
or U2663 (N_2663,N_1964,N_1773);
and U2664 (N_2664,N_1275,N_1894);
xor U2665 (N_2665,N_1793,N_1097);
and U2666 (N_2666,N_1414,N_1295);
nand U2667 (N_2667,N_1502,N_1757);
or U2668 (N_2668,N_1252,N_1624);
nor U2669 (N_2669,N_1696,N_1754);
and U2670 (N_2670,N_1289,N_1468);
nor U2671 (N_2671,N_1265,N_1018);
xor U2672 (N_2672,N_1880,N_1646);
nor U2673 (N_2673,N_1135,N_1345);
and U2674 (N_2674,N_1984,N_1595);
nand U2675 (N_2675,N_1668,N_1376);
nand U2676 (N_2676,N_1499,N_1275);
nand U2677 (N_2677,N_1335,N_1685);
nand U2678 (N_2678,N_1890,N_1673);
xor U2679 (N_2679,N_1139,N_1954);
xnor U2680 (N_2680,N_1113,N_1262);
nand U2681 (N_2681,N_1574,N_1786);
or U2682 (N_2682,N_1808,N_1101);
nand U2683 (N_2683,N_1734,N_1371);
nor U2684 (N_2684,N_1551,N_1142);
and U2685 (N_2685,N_1390,N_1626);
or U2686 (N_2686,N_1528,N_1014);
nand U2687 (N_2687,N_1938,N_1742);
or U2688 (N_2688,N_1267,N_1073);
or U2689 (N_2689,N_1181,N_1879);
xor U2690 (N_2690,N_1632,N_1993);
nor U2691 (N_2691,N_1581,N_1425);
xor U2692 (N_2692,N_1192,N_1108);
nand U2693 (N_2693,N_1456,N_1770);
or U2694 (N_2694,N_1402,N_1883);
nand U2695 (N_2695,N_1829,N_1369);
xnor U2696 (N_2696,N_1333,N_1119);
and U2697 (N_2697,N_1972,N_1929);
nor U2698 (N_2698,N_1397,N_1768);
and U2699 (N_2699,N_1594,N_1571);
and U2700 (N_2700,N_1274,N_1010);
nand U2701 (N_2701,N_1089,N_1433);
or U2702 (N_2702,N_1229,N_1640);
and U2703 (N_2703,N_1074,N_1594);
or U2704 (N_2704,N_1537,N_1446);
xnor U2705 (N_2705,N_1252,N_1758);
or U2706 (N_2706,N_1484,N_1736);
xor U2707 (N_2707,N_1131,N_1080);
nor U2708 (N_2708,N_1411,N_1721);
xor U2709 (N_2709,N_1404,N_1683);
and U2710 (N_2710,N_1072,N_1039);
and U2711 (N_2711,N_1579,N_1883);
and U2712 (N_2712,N_1721,N_1410);
or U2713 (N_2713,N_1695,N_1442);
xor U2714 (N_2714,N_1058,N_1742);
or U2715 (N_2715,N_1666,N_1328);
xnor U2716 (N_2716,N_1752,N_1018);
and U2717 (N_2717,N_1633,N_1158);
nor U2718 (N_2718,N_1277,N_1133);
nor U2719 (N_2719,N_1895,N_1063);
nand U2720 (N_2720,N_1795,N_1541);
or U2721 (N_2721,N_1547,N_1621);
or U2722 (N_2722,N_1164,N_1870);
or U2723 (N_2723,N_1746,N_1558);
and U2724 (N_2724,N_1413,N_1437);
nor U2725 (N_2725,N_1161,N_1097);
nand U2726 (N_2726,N_1832,N_1929);
and U2727 (N_2727,N_1383,N_1284);
or U2728 (N_2728,N_1734,N_1054);
nor U2729 (N_2729,N_1568,N_1671);
xnor U2730 (N_2730,N_1946,N_1373);
or U2731 (N_2731,N_1972,N_1049);
xor U2732 (N_2732,N_1856,N_1070);
or U2733 (N_2733,N_1570,N_1995);
xor U2734 (N_2734,N_1669,N_1171);
or U2735 (N_2735,N_1836,N_1863);
nand U2736 (N_2736,N_1257,N_1396);
nor U2737 (N_2737,N_1523,N_1633);
xor U2738 (N_2738,N_1306,N_1027);
and U2739 (N_2739,N_1152,N_1300);
xnor U2740 (N_2740,N_1932,N_1599);
nor U2741 (N_2741,N_1402,N_1950);
xnor U2742 (N_2742,N_1979,N_1019);
nand U2743 (N_2743,N_1824,N_1145);
or U2744 (N_2744,N_1106,N_1783);
nand U2745 (N_2745,N_1677,N_1000);
nor U2746 (N_2746,N_1582,N_1923);
or U2747 (N_2747,N_1803,N_1834);
or U2748 (N_2748,N_1087,N_1764);
nor U2749 (N_2749,N_1944,N_1598);
or U2750 (N_2750,N_1254,N_1315);
and U2751 (N_2751,N_1827,N_1409);
nand U2752 (N_2752,N_1398,N_1510);
nand U2753 (N_2753,N_1653,N_1402);
xor U2754 (N_2754,N_1627,N_1843);
nor U2755 (N_2755,N_1638,N_1802);
nand U2756 (N_2756,N_1295,N_1537);
nor U2757 (N_2757,N_1309,N_1415);
or U2758 (N_2758,N_1756,N_1433);
nor U2759 (N_2759,N_1588,N_1866);
nand U2760 (N_2760,N_1178,N_1672);
nor U2761 (N_2761,N_1722,N_1902);
nor U2762 (N_2762,N_1234,N_1006);
and U2763 (N_2763,N_1731,N_1816);
and U2764 (N_2764,N_1593,N_1792);
xor U2765 (N_2765,N_1822,N_1779);
or U2766 (N_2766,N_1178,N_1758);
nor U2767 (N_2767,N_1498,N_1765);
or U2768 (N_2768,N_1963,N_1449);
and U2769 (N_2769,N_1418,N_1845);
nor U2770 (N_2770,N_1696,N_1373);
nand U2771 (N_2771,N_1678,N_1688);
nor U2772 (N_2772,N_1360,N_1621);
and U2773 (N_2773,N_1773,N_1636);
nor U2774 (N_2774,N_1879,N_1378);
xnor U2775 (N_2775,N_1514,N_1715);
and U2776 (N_2776,N_1772,N_1784);
or U2777 (N_2777,N_1004,N_1308);
nand U2778 (N_2778,N_1593,N_1669);
xnor U2779 (N_2779,N_1810,N_1028);
nor U2780 (N_2780,N_1924,N_1025);
nor U2781 (N_2781,N_1680,N_1830);
and U2782 (N_2782,N_1581,N_1261);
nand U2783 (N_2783,N_1601,N_1334);
and U2784 (N_2784,N_1723,N_1729);
and U2785 (N_2785,N_1938,N_1503);
or U2786 (N_2786,N_1862,N_1838);
xor U2787 (N_2787,N_1500,N_1470);
xor U2788 (N_2788,N_1619,N_1084);
or U2789 (N_2789,N_1292,N_1501);
and U2790 (N_2790,N_1679,N_1964);
and U2791 (N_2791,N_1495,N_1059);
nor U2792 (N_2792,N_1193,N_1995);
nand U2793 (N_2793,N_1812,N_1458);
and U2794 (N_2794,N_1178,N_1761);
nand U2795 (N_2795,N_1555,N_1659);
and U2796 (N_2796,N_1959,N_1233);
nor U2797 (N_2797,N_1517,N_1589);
and U2798 (N_2798,N_1282,N_1680);
nor U2799 (N_2799,N_1360,N_1324);
nand U2800 (N_2800,N_1186,N_1004);
nand U2801 (N_2801,N_1038,N_1525);
and U2802 (N_2802,N_1280,N_1197);
xnor U2803 (N_2803,N_1027,N_1781);
or U2804 (N_2804,N_1631,N_1697);
and U2805 (N_2805,N_1654,N_1898);
xor U2806 (N_2806,N_1651,N_1462);
xor U2807 (N_2807,N_1919,N_1098);
or U2808 (N_2808,N_1509,N_1594);
and U2809 (N_2809,N_1476,N_1924);
nor U2810 (N_2810,N_1751,N_1005);
or U2811 (N_2811,N_1105,N_1881);
or U2812 (N_2812,N_1681,N_1921);
xor U2813 (N_2813,N_1747,N_1204);
nor U2814 (N_2814,N_1856,N_1919);
nand U2815 (N_2815,N_1436,N_1262);
or U2816 (N_2816,N_1896,N_1677);
nor U2817 (N_2817,N_1549,N_1859);
or U2818 (N_2818,N_1210,N_1277);
xor U2819 (N_2819,N_1891,N_1785);
nand U2820 (N_2820,N_1043,N_1380);
nand U2821 (N_2821,N_1295,N_1875);
xnor U2822 (N_2822,N_1472,N_1212);
nand U2823 (N_2823,N_1776,N_1774);
nor U2824 (N_2824,N_1213,N_1720);
or U2825 (N_2825,N_1860,N_1490);
and U2826 (N_2826,N_1335,N_1859);
nor U2827 (N_2827,N_1955,N_1730);
nor U2828 (N_2828,N_1792,N_1208);
or U2829 (N_2829,N_1732,N_1698);
nor U2830 (N_2830,N_1889,N_1634);
nand U2831 (N_2831,N_1628,N_1882);
or U2832 (N_2832,N_1104,N_1477);
or U2833 (N_2833,N_1532,N_1374);
nor U2834 (N_2834,N_1224,N_1928);
nor U2835 (N_2835,N_1667,N_1364);
or U2836 (N_2836,N_1772,N_1358);
and U2837 (N_2837,N_1217,N_1815);
nor U2838 (N_2838,N_1417,N_1585);
or U2839 (N_2839,N_1702,N_1321);
or U2840 (N_2840,N_1769,N_1507);
nor U2841 (N_2841,N_1600,N_1426);
nor U2842 (N_2842,N_1545,N_1698);
and U2843 (N_2843,N_1136,N_1369);
xor U2844 (N_2844,N_1644,N_1730);
xnor U2845 (N_2845,N_1145,N_1749);
nor U2846 (N_2846,N_1811,N_1343);
and U2847 (N_2847,N_1534,N_1959);
or U2848 (N_2848,N_1910,N_1287);
nor U2849 (N_2849,N_1157,N_1675);
nor U2850 (N_2850,N_1815,N_1441);
nor U2851 (N_2851,N_1478,N_1470);
or U2852 (N_2852,N_1294,N_1122);
nor U2853 (N_2853,N_1791,N_1920);
xor U2854 (N_2854,N_1783,N_1220);
xnor U2855 (N_2855,N_1188,N_1305);
and U2856 (N_2856,N_1440,N_1536);
nor U2857 (N_2857,N_1063,N_1036);
xor U2858 (N_2858,N_1804,N_1489);
nand U2859 (N_2859,N_1419,N_1530);
nand U2860 (N_2860,N_1450,N_1421);
nor U2861 (N_2861,N_1566,N_1988);
or U2862 (N_2862,N_1468,N_1637);
or U2863 (N_2863,N_1682,N_1794);
and U2864 (N_2864,N_1348,N_1222);
nor U2865 (N_2865,N_1976,N_1424);
nor U2866 (N_2866,N_1803,N_1467);
nand U2867 (N_2867,N_1212,N_1329);
or U2868 (N_2868,N_1083,N_1579);
nor U2869 (N_2869,N_1008,N_1240);
nand U2870 (N_2870,N_1360,N_1978);
nor U2871 (N_2871,N_1103,N_1132);
and U2872 (N_2872,N_1312,N_1048);
nand U2873 (N_2873,N_1679,N_1338);
xor U2874 (N_2874,N_1809,N_1752);
and U2875 (N_2875,N_1869,N_1444);
xnor U2876 (N_2876,N_1770,N_1832);
xor U2877 (N_2877,N_1240,N_1348);
or U2878 (N_2878,N_1839,N_1031);
nor U2879 (N_2879,N_1674,N_1083);
nor U2880 (N_2880,N_1004,N_1517);
or U2881 (N_2881,N_1831,N_1319);
or U2882 (N_2882,N_1113,N_1663);
nand U2883 (N_2883,N_1576,N_1625);
nand U2884 (N_2884,N_1098,N_1510);
nor U2885 (N_2885,N_1641,N_1512);
or U2886 (N_2886,N_1303,N_1196);
or U2887 (N_2887,N_1329,N_1318);
and U2888 (N_2888,N_1789,N_1294);
nand U2889 (N_2889,N_1301,N_1396);
nor U2890 (N_2890,N_1117,N_1894);
nand U2891 (N_2891,N_1986,N_1475);
nor U2892 (N_2892,N_1667,N_1391);
xor U2893 (N_2893,N_1251,N_1581);
and U2894 (N_2894,N_1665,N_1850);
nor U2895 (N_2895,N_1719,N_1353);
nor U2896 (N_2896,N_1056,N_1152);
and U2897 (N_2897,N_1631,N_1087);
xor U2898 (N_2898,N_1882,N_1536);
xor U2899 (N_2899,N_1404,N_1790);
or U2900 (N_2900,N_1403,N_1198);
and U2901 (N_2901,N_1151,N_1599);
nand U2902 (N_2902,N_1545,N_1442);
or U2903 (N_2903,N_1661,N_1296);
nand U2904 (N_2904,N_1939,N_1123);
and U2905 (N_2905,N_1187,N_1690);
nand U2906 (N_2906,N_1299,N_1554);
nand U2907 (N_2907,N_1033,N_1518);
and U2908 (N_2908,N_1142,N_1211);
or U2909 (N_2909,N_1034,N_1556);
nand U2910 (N_2910,N_1880,N_1455);
xor U2911 (N_2911,N_1283,N_1896);
nand U2912 (N_2912,N_1525,N_1869);
or U2913 (N_2913,N_1558,N_1410);
nand U2914 (N_2914,N_1523,N_1783);
nand U2915 (N_2915,N_1667,N_1422);
nand U2916 (N_2916,N_1957,N_1760);
or U2917 (N_2917,N_1690,N_1644);
xnor U2918 (N_2918,N_1672,N_1209);
nand U2919 (N_2919,N_1283,N_1922);
nor U2920 (N_2920,N_1065,N_1134);
nand U2921 (N_2921,N_1510,N_1729);
and U2922 (N_2922,N_1816,N_1014);
xnor U2923 (N_2923,N_1809,N_1332);
nor U2924 (N_2924,N_1103,N_1072);
nand U2925 (N_2925,N_1486,N_1175);
or U2926 (N_2926,N_1544,N_1682);
nand U2927 (N_2927,N_1344,N_1597);
xor U2928 (N_2928,N_1257,N_1715);
and U2929 (N_2929,N_1828,N_1645);
nor U2930 (N_2930,N_1491,N_1313);
and U2931 (N_2931,N_1681,N_1601);
nand U2932 (N_2932,N_1074,N_1599);
xnor U2933 (N_2933,N_1487,N_1834);
nand U2934 (N_2934,N_1268,N_1215);
or U2935 (N_2935,N_1765,N_1223);
or U2936 (N_2936,N_1878,N_1272);
and U2937 (N_2937,N_1502,N_1799);
nor U2938 (N_2938,N_1550,N_1463);
nor U2939 (N_2939,N_1826,N_1098);
nand U2940 (N_2940,N_1525,N_1699);
xor U2941 (N_2941,N_1525,N_1903);
xnor U2942 (N_2942,N_1707,N_1734);
and U2943 (N_2943,N_1535,N_1633);
or U2944 (N_2944,N_1022,N_1730);
nand U2945 (N_2945,N_1620,N_1883);
or U2946 (N_2946,N_1503,N_1098);
and U2947 (N_2947,N_1095,N_1758);
nor U2948 (N_2948,N_1839,N_1289);
xor U2949 (N_2949,N_1762,N_1949);
or U2950 (N_2950,N_1608,N_1712);
xnor U2951 (N_2951,N_1224,N_1619);
or U2952 (N_2952,N_1100,N_1970);
and U2953 (N_2953,N_1944,N_1254);
and U2954 (N_2954,N_1361,N_1039);
nor U2955 (N_2955,N_1654,N_1684);
or U2956 (N_2956,N_1208,N_1678);
or U2957 (N_2957,N_1745,N_1537);
nand U2958 (N_2958,N_1253,N_1970);
nor U2959 (N_2959,N_1416,N_1079);
nand U2960 (N_2960,N_1740,N_1424);
nor U2961 (N_2961,N_1862,N_1331);
nor U2962 (N_2962,N_1462,N_1284);
or U2963 (N_2963,N_1280,N_1015);
nor U2964 (N_2964,N_1841,N_1872);
nor U2965 (N_2965,N_1968,N_1850);
or U2966 (N_2966,N_1562,N_1064);
or U2967 (N_2967,N_1012,N_1422);
nand U2968 (N_2968,N_1551,N_1105);
nand U2969 (N_2969,N_1587,N_1024);
or U2970 (N_2970,N_1726,N_1248);
nand U2971 (N_2971,N_1991,N_1485);
nor U2972 (N_2972,N_1724,N_1456);
xnor U2973 (N_2973,N_1952,N_1782);
and U2974 (N_2974,N_1902,N_1216);
or U2975 (N_2975,N_1788,N_1460);
and U2976 (N_2976,N_1497,N_1271);
nand U2977 (N_2977,N_1828,N_1672);
nor U2978 (N_2978,N_1293,N_1804);
xnor U2979 (N_2979,N_1443,N_1415);
or U2980 (N_2980,N_1288,N_1548);
and U2981 (N_2981,N_1643,N_1081);
or U2982 (N_2982,N_1040,N_1864);
xnor U2983 (N_2983,N_1555,N_1075);
or U2984 (N_2984,N_1516,N_1824);
or U2985 (N_2985,N_1644,N_1040);
nor U2986 (N_2986,N_1549,N_1709);
nand U2987 (N_2987,N_1097,N_1466);
xnor U2988 (N_2988,N_1816,N_1190);
nor U2989 (N_2989,N_1397,N_1412);
and U2990 (N_2990,N_1727,N_1313);
xor U2991 (N_2991,N_1049,N_1461);
and U2992 (N_2992,N_1066,N_1280);
and U2993 (N_2993,N_1612,N_1137);
xor U2994 (N_2994,N_1274,N_1574);
nand U2995 (N_2995,N_1481,N_1250);
and U2996 (N_2996,N_1369,N_1834);
nor U2997 (N_2997,N_1426,N_1881);
nand U2998 (N_2998,N_1592,N_1503);
or U2999 (N_2999,N_1894,N_1363);
nor U3000 (N_3000,N_2583,N_2744);
or U3001 (N_3001,N_2747,N_2011);
xnor U3002 (N_3002,N_2914,N_2053);
nand U3003 (N_3003,N_2395,N_2519);
nand U3004 (N_3004,N_2363,N_2778);
or U3005 (N_3005,N_2823,N_2738);
nand U3006 (N_3006,N_2252,N_2824);
nand U3007 (N_3007,N_2806,N_2767);
or U3008 (N_3008,N_2677,N_2568);
xor U3009 (N_3009,N_2024,N_2241);
nor U3010 (N_3010,N_2840,N_2856);
or U3011 (N_3011,N_2885,N_2190);
nand U3012 (N_3012,N_2484,N_2701);
or U3013 (N_3013,N_2996,N_2259);
xnor U3014 (N_3014,N_2348,N_2075);
nor U3015 (N_3015,N_2875,N_2869);
xnor U3016 (N_3016,N_2644,N_2793);
nor U3017 (N_3017,N_2832,N_2740);
and U3018 (N_3018,N_2313,N_2444);
or U3019 (N_3019,N_2043,N_2081);
nor U3020 (N_3020,N_2991,N_2550);
nor U3021 (N_3021,N_2551,N_2238);
xor U3022 (N_3022,N_2896,N_2143);
nor U3023 (N_3023,N_2822,N_2299);
xor U3024 (N_3024,N_2720,N_2347);
nand U3025 (N_3025,N_2023,N_2451);
and U3026 (N_3026,N_2144,N_2138);
xnor U3027 (N_3027,N_2935,N_2052);
nand U3028 (N_3028,N_2650,N_2357);
or U3029 (N_3029,N_2322,N_2157);
nand U3030 (N_3030,N_2697,N_2292);
or U3031 (N_3031,N_2161,N_2243);
and U3032 (N_3032,N_2314,N_2445);
and U3033 (N_3033,N_2850,N_2848);
xnor U3034 (N_3034,N_2761,N_2758);
xor U3035 (N_3035,N_2585,N_2891);
nand U3036 (N_3036,N_2393,N_2189);
and U3037 (N_3037,N_2754,N_2387);
and U3038 (N_3038,N_2984,N_2584);
nand U3039 (N_3039,N_2825,N_2777);
or U3040 (N_3040,N_2063,N_2084);
nand U3041 (N_3041,N_2766,N_2739);
or U3042 (N_3042,N_2477,N_2979);
nor U3043 (N_3043,N_2236,N_2301);
and U3044 (N_3044,N_2741,N_2352);
nor U3045 (N_3045,N_2155,N_2340);
nor U3046 (N_3046,N_2125,N_2006);
nor U3047 (N_3047,N_2337,N_2452);
nand U3048 (N_3048,N_2464,N_2310);
and U3049 (N_3049,N_2315,N_2845);
nor U3050 (N_3050,N_2210,N_2103);
and U3051 (N_3051,N_2226,N_2201);
xor U3052 (N_3052,N_2569,N_2255);
nor U3053 (N_3053,N_2406,N_2779);
nand U3054 (N_3054,N_2405,N_2209);
and U3055 (N_3055,N_2642,N_2366);
and U3056 (N_3056,N_2507,N_2408);
xor U3057 (N_3057,N_2705,N_2272);
nor U3058 (N_3058,N_2102,N_2808);
nor U3059 (N_3059,N_2829,N_2715);
nand U3060 (N_3060,N_2533,N_2244);
and U3061 (N_3061,N_2966,N_2695);
nand U3062 (N_3062,N_2246,N_2265);
nor U3063 (N_3063,N_2199,N_2593);
nand U3064 (N_3064,N_2001,N_2546);
and U3065 (N_3065,N_2294,N_2932);
or U3066 (N_3066,N_2798,N_2578);
nor U3067 (N_3067,N_2819,N_2416);
xnor U3068 (N_3068,N_2906,N_2940);
and U3069 (N_3069,N_2217,N_2909);
xor U3070 (N_3070,N_2517,N_2942);
xnor U3071 (N_3071,N_2400,N_2712);
nor U3072 (N_3072,N_2537,N_2501);
and U3073 (N_3073,N_2689,N_2582);
nor U3074 (N_3074,N_2671,N_2730);
or U3075 (N_3075,N_2344,N_2958);
nand U3076 (N_3076,N_2388,N_2609);
or U3077 (N_3077,N_2723,N_2992);
nor U3078 (N_3078,N_2545,N_2382);
xor U3079 (N_3079,N_2118,N_2888);
and U3080 (N_3080,N_2279,N_2639);
nand U3081 (N_3081,N_2802,N_2604);
nor U3082 (N_3082,N_2918,N_2008);
nor U3083 (N_3083,N_2688,N_2627);
and U3084 (N_3084,N_2605,N_2794);
nand U3085 (N_3085,N_2105,N_2756);
xnor U3086 (N_3086,N_2950,N_2436);
nand U3087 (N_3087,N_2435,N_2101);
nand U3088 (N_3088,N_2775,N_2359);
nand U3089 (N_3089,N_2865,N_2540);
or U3090 (N_3090,N_2805,N_2547);
nor U3091 (N_3091,N_2233,N_2036);
nand U3092 (N_3092,N_2166,N_2629);
nor U3093 (N_3093,N_2580,N_2556);
and U3094 (N_3094,N_2191,N_2197);
and U3095 (N_3095,N_2770,N_2658);
nand U3096 (N_3096,N_2200,N_2768);
nand U3097 (N_3097,N_2474,N_2470);
or U3098 (N_3098,N_2836,N_2413);
xor U3099 (N_3099,N_2354,N_2598);
or U3100 (N_3100,N_2251,N_2543);
nor U3101 (N_3101,N_2085,N_2835);
nor U3102 (N_3102,N_2820,N_2857);
and U3103 (N_3103,N_2208,N_2216);
or U3104 (N_3104,N_2345,N_2659);
xnor U3105 (N_3105,N_2669,N_2681);
or U3106 (N_3106,N_2446,N_2789);
nand U3107 (N_3107,N_2089,N_2266);
nand U3108 (N_3108,N_2367,N_2336);
nor U3109 (N_3109,N_2920,N_2552);
and U3110 (N_3110,N_2643,N_2263);
or U3111 (N_3111,N_2146,N_2019);
xor U3112 (N_3112,N_2130,N_2404);
xnor U3113 (N_3113,N_2311,N_2248);
or U3114 (N_3114,N_2535,N_2432);
or U3115 (N_3115,N_2158,N_2454);
xor U3116 (N_3116,N_2505,N_2046);
and U3117 (N_3117,N_2338,N_2066);
xor U3118 (N_3118,N_2257,N_2792);
and U3119 (N_3119,N_2874,N_2068);
nand U3120 (N_3120,N_2132,N_2734);
or U3121 (N_3121,N_2278,N_2633);
xnor U3122 (N_3122,N_2092,N_2441);
nor U3123 (N_3123,N_2635,N_2087);
and U3124 (N_3124,N_2951,N_2443);
or U3125 (N_3125,N_2884,N_2676);
xnor U3126 (N_3126,N_2440,N_2258);
nor U3127 (N_3127,N_2219,N_2109);
or U3128 (N_3128,N_2119,N_2182);
or U3129 (N_3129,N_2668,N_2973);
nand U3130 (N_3130,N_2468,N_2229);
nand U3131 (N_3131,N_2579,N_2064);
xor U3132 (N_3132,N_2104,N_2523);
and U3133 (N_3133,N_2864,N_2073);
nor U3134 (N_3134,N_2924,N_2800);
nor U3135 (N_3135,N_2780,N_2013);
or U3136 (N_3136,N_2079,N_2462);
nor U3137 (N_3137,N_2370,N_2895);
and U3138 (N_3138,N_2967,N_2287);
or U3139 (N_3139,N_2760,N_2174);
or U3140 (N_3140,N_2649,N_2883);
xnor U3141 (N_3141,N_2458,N_2981);
and U3142 (N_3142,N_2284,N_2675);
or U3143 (N_3143,N_2804,N_2810);
nand U3144 (N_3144,N_2877,N_2486);
nand U3145 (N_3145,N_2274,N_2862);
nor U3146 (N_3146,N_2015,N_2696);
nor U3147 (N_3147,N_2300,N_2149);
or U3148 (N_3148,N_2324,N_2613);
nor U3149 (N_3149,N_2449,N_2686);
and U3150 (N_3150,N_2892,N_2059);
xor U3151 (N_3151,N_2010,N_2323);
nor U3152 (N_3152,N_2047,N_2123);
or U3153 (N_3153,N_2502,N_2070);
nor U3154 (N_3154,N_2306,N_2586);
or U3155 (N_3155,N_2727,N_2271);
or U3156 (N_3156,N_2420,N_2841);
xor U3157 (N_3157,N_2662,N_2719);
xnor U3158 (N_3158,N_2136,N_2687);
nand U3159 (N_3159,N_2709,N_2012);
xor U3160 (N_3160,N_2383,N_2234);
nand U3161 (N_3161,N_2482,N_2751);
xnor U3162 (N_3162,N_2389,N_2009);
nor U3163 (N_3163,N_2964,N_2773);
nor U3164 (N_3164,N_2496,N_2051);
xnor U3165 (N_3165,N_2512,N_2317);
nand U3166 (N_3166,N_2625,N_2384);
xnor U3167 (N_3167,N_2941,N_2492);
xnor U3168 (N_3168,N_2060,N_2706);
and U3169 (N_3169,N_2926,N_2016);
xor U3170 (N_3170,N_2281,N_2142);
or U3171 (N_3171,N_2231,N_2373);
xnor U3172 (N_3172,N_2624,N_2638);
or U3173 (N_3173,N_2227,N_2426);
or U3174 (N_3174,N_2499,N_2156);
and U3175 (N_3175,N_2953,N_2249);
nand U3176 (N_3176,N_2737,N_2150);
xor U3177 (N_3177,N_2530,N_2333);
xnor U3178 (N_3178,N_2980,N_2378);
nand U3179 (N_3179,N_2350,N_2678);
nand U3180 (N_3180,N_2134,N_2776);
nand U3181 (N_3181,N_2375,N_2048);
xor U3182 (N_3182,N_2790,N_2399);
nor U3183 (N_3183,N_2151,N_2276);
xor U3184 (N_3184,N_2831,N_2893);
nand U3185 (N_3185,N_2606,N_2564);
and U3186 (N_3186,N_2974,N_2553);
or U3187 (N_3187,N_2765,N_2392);
and U3188 (N_3188,N_2796,N_2516);
and U3189 (N_3189,N_2423,N_2140);
xnor U3190 (N_3190,N_2970,N_2722);
or U3191 (N_3191,N_2693,N_2448);
or U3192 (N_3192,N_2077,N_2180);
xnor U3193 (N_3193,N_2622,N_2628);
xor U3194 (N_3194,N_2372,N_2901);
xor U3195 (N_3195,N_2503,N_2952);
nand U3196 (N_3196,N_2033,N_2116);
or U3197 (N_3197,N_2341,N_2990);
xnor U3198 (N_3198,N_2721,N_2554);
and U3199 (N_3199,N_2167,N_2514);
xnor U3200 (N_3200,N_2198,N_2963);
xor U3201 (N_3201,N_2853,N_2506);
nor U3202 (N_3202,N_2307,N_2202);
nor U3203 (N_3203,N_2124,N_2031);
and U3204 (N_3204,N_2945,N_2871);
or U3205 (N_3205,N_2025,N_2922);
or U3206 (N_3206,N_2928,N_2529);
or U3207 (N_3207,N_2782,N_2356);
xnor U3208 (N_3208,N_2330,N_2645);
nand U3209 (N_3209,N_2899,N_2817);
nand U3210 (N_3210,N_2193,N_2196);
xnor U3211 (N_3211,N_2524,N_2828);
and U3212 (N_3212,N_2195,N_2478);
nand U3213 (N_3213,N_2746,N_2729);
nand U3214 (N_3214,N_2129,N_2660);
nor U3215 (N_3215,N_2685,N_2342);
xnor U3216 (N_3216,N_2937,N_2612);
xor U3217 (N_3217,N_2139,N_2762);
nand U3218 (N_3218,N_2401,N_2791);
nor U3219 (N_3219,N_2285,N_2457);
xor U3220 (N_3220,N_2250,N_2328);
or U3221 (N_3221,N_2614,N_2528);
nand U3222 (N_3222,N_2018,N_2108);
xor U3223 (N_3223,N_2312,N_2346);
nand U3224 (N_3224,N_2700,N_2954);
nor U3225 (N_3225,N_2785,N_2663);
or U3226 (N_3226,N_2898,N_2931);
nor U3227 (N_3227,N_2293,N_2801);
xnor U3228 (N_3228,N_2597,N_2000);
and U3229 (N_3229,N_2335,N_2807);
xor U3230 (N_3230,N_2083,N_2673);
xor U3231 (N_3231,N_2093,N_2542);
nand U3232 (N_3232,N_2602,N_2419);
xnor U3233 (N_3233,N_2286,N_2131);
xor U3234 (N_3234,N_2106,N_2728);
nand U3235 (N_3235,N_2480,N_2332);
nor U3236 (N_3236,N_2814,N_2757);
and U3237 (N_3237,N_2680,N_2923);
nand U3238 (N_3238,N_2733,N_2071);
and U3239 (N_3239,N_2100,N_2993);
or U3240 (N_3240,N_2570,N_2652);
and U3241 (N_3241,N_2632,N_2647);
xnor U3242 (N_3242,N_2962,N_2165);
nor U3243 (N_3243,N_2913,N_2218);
nor U3244 (N_3244,N_2032,N_2656);
or U3245 (N_3245,N_2122,N_2572);
nor U3246 (N_3246,N_2510,N_2254);
or U3247 (N_3247,N_2107,N_2887);
nor U3248 (N_3248,N_2611,N_2262);
and U3249 (N_3249,N_2170,N_2177);
nor U3250 (N_3250,N_2223,N_2619);
and U3251 (N_3251,N_2058,N_2859);
and U3252 (N_3252,N_2368,N_2925);
nand U3253 (N_3253,N_2753,N_2654);
xnor U3254 (N_3254,N_2969,N_2438);
nand U3255 (N_3255,N_2641,N_2221);
xnor U3256 (N_3256,N_2587,N_2456);
nand U3257 (N_3257,N_2160,N_2475);
or U3258 (N_3258,N_2181,N_2975);
and U3259 (N_3259,N_2225,N_2133);
xor U3260 (N_3260,N_2699,N_2162);
and U3261 (N_3261,N_2826,N_2184);
nor U3262 (N_3262,N_2422,N_2522);
xor U3263 (N_3263,N_2646,N_2799);
or U3264 (N_3264,N_2994,N_2603);
nor U3265 (N_3265,N_2844,N_2186);
and U3266 (N_3266,N_2487,N_2539);
nor U3267 (N_3267,N_2703,N_2041);
or U3268 (N_3268,N_2986,N_2493);
or U3269 (N_3269,N_2168,N_2500);
nand U3270 (N_3270,N_2872,N_2291);
or U3271 (N_3271,N_2921,N_2949);
nor U3272 (N_3272,N_2380,N_2621);
nor U3273 (N_3273,N_2868,N_2490);
nor U3274 (N_3274,N_2434,N_2617);
and U3275 (N_3275,N_2985,N_2711);
nor U3276 (N_3276,N_2188,N_2163);
nand U3277 (N_3277,N_2939,N_2618);
and U3278 (N_3278,N_2704,N_2304);
nand U3279 (N_3279,N_2439,N_2726);
nand U3280 (N_3280,N_2691,N_2082);
nor U3281 (N_3281,N_2636,N_2425);
and U3282 (N_3282,N_2110,N_2904);
and U3283 (N_3283,N_2878,N_2781);
and U3284 (N_3284,N_2096,N_2956);
xnor U3285 (N_3285,N_2067,N_2538);
xnor U3286 (N_3286,N_2890,N_2620);
nand U3287 (N_3287,N_2460,N_2682);
or U3288 (N_3288,N_2215,N_2044);
or U3289 (N_3289,N_2637,N_2424);
nand U3290 (N_3290,N_2090,N_2521);
or U3291 (N_3291,N_2948,N_2289);
and U3292 (N_3292,N_2361,N_2560);
nand U3293 (N_3293,N_2437,N_2900);
nand U3294 (N_3294,N_2398,N_2111);
or U3295 (N_3295,N_2021,N_2837);
nand U3296 (N_3296,N_2852,N_2718);
xor U3297 (N_3297,N_2830,N_2376);
xnor U3298 (N_3298,N_2183,N_2504);
nand U3299 (N_3299,N_2026,N_2206);
nor U3300 (N_3300,N_2957,N_2115);
xnor U3301 (N_3301,N_2567,N_2034);
or U3302 (N_3302,N_2247,N_2412);
or U3303 (N_3303,N_2045,N_2237);
and U3304 (N_3304,N_2783,N_2752);
and U3305 (N_3305,N_2428,N_2938);
and U3306 (N_3306,N_2809,N_2549);
nor U3307 (N_3307,N_2724,N_2288);
and U3308 (N_3308,N_2407,N_2402);
and U3309 (N_3309,N_2472,N_2694);
nand U3310 (N_3310,N_2147,N_2577);
xor U3311 (N_3311,N_2483,N_2999);
nand U3312 (N_3312,N_2745,N_2455);
nor U3313 (N_3313,N_2295,N_2961);
nor U3314 (N_3314,N_2185,N_2467);
or U3315 (N_3315,N_2327,N_2816);
nand U3316 (N_3316,N_2381,N_2880);
xor U3317 (N_3317,N_2450,N_2769);
and U3318 (N_3318,N_2919,N_2318);
nand U3319 (N_3319,N_2471,N_2326);
or U3320 (N_3320,N_2113,N_2651);
nand U3321 (N_3321,N_2847,N_2261);
nand U3322 (N_3322,N_2860,N_2433);
nand U3323 (N_3323,N_2035,N_2911);
xor U3324 (N_3324,N_2520,N_2169);
nor U3325 (N_3325,N_2269,N_2396);
or U3326 (N_3326,N_2098,N_2846);
xnor U3327 (N_3327,N_2273,N_2022);
nand U3328 (N_3328,N_2264,N_2411);
nand U3329 (N_3329,N_2683,N_2665);
nor U3330 (N_3330,N_2204,N_2615);
nor U3331 (N_3331,N_2002,N_2374);
nand U3332 (N_3332,N_2245,N_2971);
and U3333 (N_3333,N_2494,N_2316);
and U3334 (N_3334,N_2735,N_2297);
nand U3335 (N_3335,N_2561,N_2391);
and U3336 (N_3336,N_2091,N_2390);
nor U3337 (N_3337,N_2469,N_2095);
nor U3338 (N_3338,N_2811,N_2054);
xnor U3339 (N_3339,N_2056,N_2972);
or U3340 (N_3340,N_2498,N_2803);
or U3341 (N_3341,N_2086,N_2797);
nand U3342 (N_3342,N_2936,N_2515);
nand U3343 (N_3343,N_2061,N_2566);
nor U3344 (N_3344,N_2959,N_2707);
xor U3345 (N_3345,N_2861,N_2573);
and U3346 (N_3346,N_2187,N_2815);
and U3347 (N_3347,N_2589,N_2159);
nand U3348 (N_3348,N_2518,N_2759);
xor U3349 (N_3349,N_2334,N_2838);
xor U3350 (N_3350,N_2581,N_2296);
nor U3351 (N_3351,N_2369,N_2339);
or U3352 (N_3352,N_2930,N_2447);
and U3353 (N_3353,N_2253,N_2750);
nor U3354 (N_3354,N_2536,N_2988);
xnor U3355 (N_3355,N_2329,N_2145);
and U3356 (N_3356,N_2626,N_2596);
nand U3357 (N_3357,N_2851,N_2321);
xnor U3358 (N_3358,N_2353,N_2302);
and U3359 (N_3359,N_2934,N_2319);
or U3360 (N_3360,N_2179,N_2127);
nand U3361 (N_3361,N_2601,N_2983);
nor U3362 (N_3362,N_2176,N_2866);
or U3363 (N_3363,N_2563,N_2708);
nand U3364 (N_3364,N_2020,N_2473);
or U3365 (N_3365,N_2194,N_2833);
and U3366 (N_3366,N_2591,N_2076);
and U3367 (N_3367,N_2982,N_2927);
nor U3368 (N_3368,N_2213,N_2559);
or U3369 (N_3369,N_2574,N_2164);
or U3370 (N_3370,N_2039,N_2097);
or U3371 (N_3371,N_2842,N_2397);
nor U3372 (N_3372,N_2575,N_2599);
and U3373 (N_3373,N_2476,N_2576);
xor U3374 (N_3374,N_2907,N_2466);
nand U3375 (N_3375,N_2394,N_2485);
or U3376 (N_3376,N_2655,N_2873);
nor U3377 (N_3377,N_2944,N_2929);
nand U3378 (N_3378,N_2128,N_2331);
or U3379 (N_3379,N_2513,N_2879);
xor U3380 (N_3380,N_2371,N_2771);
and U3381 (N_3381,N_2594,N_2672);
nand U3382 (N_3382,N_2784,N_2667);
nor U3383 (N_3383,N_2755,N_2479);
xor U3384 (N_3384,N_2192,N_2038);
xor U3385 (N_3385,N_2690,N_2062);
nand U3386 (N_3386,N_2946,N_2040);
or U3387 (N_3387,N_2894,N_2178);
nor U3388 (N_3388,N_2915,N_2349);
nand U3389 (N_3389,N_2947,N_2812);
and U3390 (N_3390,N_2634,N_2716);
or U3391 (N_3391,N_2481,N_2409);
and U3392 (N_3392,N_2495,N_2117);
or U3393 (N_3393,N_2997,N_2995);
nand U3394 (N_3394,N_2698,N_2239);
or U3395 (N_3395,N_2228,N_2736);
or U3396 (N_3396,N_2453,N_2418);
or U3397 (N_3397,N_2121,N_2674);
and U3398 (N_3398,N_2429,N_2858);
xnor U3399 (N_3399,N_2527,N_2987);
and U3400 (N_3400,N_2014,N_2379);
xnor U3401 (N_3401,N_2653,N_2876);
or U3402 (N_3402,N_2916,N_2277);
nand U3403 (N_3403,N_2787,N_2029);
xor U3404 (N_3404,N_2267,N_2714);
xor U3405 (N_3405,N_2976,N_2558);
nand U3406 (N_3406,N_2153,N_2912);
nand U3407 (N_3407,N_2532,N_2148);
nor U3408 (N_3408,N_2099,N_2640);
and U3409 (N_3409,N_2283,N_2027);
nor U3410 (N_3410,N_2943,N_2415);
nand U3411 (N_3411,N_2965,N_2114);
nand U3412 (N_3412,N_2171,N_2351);
or U3413 (N_3413,N_2005,N_2849);
nor U3414 (N_3414,N_2126,N_2205);
and U3415 (N_3415,N_2212,N_2867);
and U3416 (N_3416,N_2320,N_2902);
xnor U3417 (N_3417,N_2526,N_2275);
xnor U3418 (N_3418,N_2763,N_2430);
xor U3419 (N_3419,N_2616,N_2555);
or U3420 (N_3420,N_2571,N_2431);
nor U3421 (N_3421,N_2224,N_2074);
and U3422 (N_3422,N_2211,N_2303);
and U3423 (N_3423,N_2905,N_2141);
nand U3424 (N_3424,N_2427,N_2525);
nand U3425 (N_3425,N_2630,N_2214);
nand U3426 (N_3426,N_2989,N_2749);
and U3427 (N_3427,N_2855,N_2385);
or U3428 (N_3428,N_2355,N_2960);
or U3429 (N_3429,N_2308,N_2955);
and U3430 (N_3430,N_2137,N_2270);
nand U3431 (N_3431,N_2588,N_2028);
nand U3432 (N_3432,N_2511,N_2508);
nor U3433 (N_3433,N_2631,N_2280);
nand U3434 (N_3434,N_2886,N_2152);
xor U3435 (N_3435,N_2050,N_2112);
nand U3436 (N_3436,N_2078,N_2120);
nor U3437 (N_3437,N_2069,N_2863);
nand U3438 (N_3438,N_2978,N_2818);
or U3439 (N_3439,N_2488,N_2772);
nand U3440 (N_3440,N_2386,N_2461);
or U3441 (N_3441,N_2786,N_2364);
nor U3442 (N_3442,N_2360,N_2094);
or U3443 (N_3443,N_2442,N_2743);
nand U3444 (N_3444,N_2977,N_2203);
xor U3445 (N_3445,N_2702,N_2049);
xor U3446 (N_3446,N_2889,N_2065);
nand U3447 (N_3447,N_2421,N_2154);
xor U3448 (N_3448,N_2713,N_2135);
and U3449 (N_3449,N_2933,N_2595);
nor U3450 (N_3450,N_2897,N_2657);
and U3451 (N_3451,N_2565,N_2623);
nand U3452 (N_3452,N_2534,N_2600);
nand U3453 (N_3453,N_2088,N_2037);
nor U3454 (N_3454,N_2004,N_2666);
nor U3455 (N_3455,N_2207,N_2007);
or U3456 (N_3456,N_2417,N_2232);
and U3457 (N_3457,N_2648,N_2230);
or U3458 (N_3458,N_2240,N_2679);
nand U3459 (N_3459,N_2173,N_2220);
and U3460 (N_3460,N_2732,N_2664);
nand U3461 (N_3461,N_2017,N_2882);
or U3462 (N_3462,N_2541,N_2903);
or U3463 (N_3463,N_2491,N_2821);
or U3464 (N_3464,N_2414,N_2055);
nand U3465 (N_3465,N_2463,N_2030);
nor U3466 (N_3466,N_2410,N_2459);
nor U3467 (N_3467,N_2298,N_2608);
nand U3468 (N_3468,N_2509,N_2057);
nand U3469 (N_3469,N_2692,N_2377);
or U3470 (N_3470,N_2881,N_2268);
xnor U3471 (N_3471,N_2343,N_2764);
nor U3472 (N_3472,N_2607,N_2834);
nand U3473 (N_3473,N_2998,N_2813);
xnor U3474 (N_3474,N_2917,N_2670);
nor U3475 (N_3475,N_2172,N_2003);
or U3476 (N_3476,N_2489,N_2365);
or U3477 (N_3477,N_2731,N_2590);
or U3478 (N_3478,N_2260,N_2774);
and U3479 (N_3479,N_2592,N_2222);
or U3480 (N_3480,N_2309,N_2403);
xor U3481 (N_3481,N_2843,N_2661);
xnor U3482 (N_3482,N_2854,N_2544);
xnor U3483 (N_3483,N_2742,N_2748);
nor U3484 (N_3484,N_2465,N_2242);
xor U3485 (N_3485,N_2325,N_2725);
and U3486 (N_3486,N_2548,N_2531);
xor U3487 (N_3487,N_2710,N_2968);
nand U3488 (N_3488,N_2557,N_2362);
or U3489 (N_3489,N_2175,N_2717);
xor U3490 (N_3490,N_2497,N_2870);
nand U3491 (N_3491,N_2910,N_2042);
xnor U3492 (N_3492,N_2080,N_2562);
or U3493 (N_3493,N_2072,N_2282);
and U3494 (N_3494,N_2235,N_2827);
xnor U3495 (N_3495,N_2305,N_2256);
and U3496 (N_3496,N_2795,N_2290);
and U3497 (N_3497,N_2610,N_2358);
or U3498 (N_3498,N_2908,N_2788);
nand U3499 (N_3499,N_2684,N_2839);
xor U3500 (N_3500,N_2883,N_2850);
and U3501 (N_3501,N_2387,N_2600);
xor U3502 (N_3502,N_2162,N_2784);
nor U3503 (N_3503,N_2843,N_2897);
or U3504 (N_3504,N_2844,N_2628);
nor U3505 (N_3505,N_2485,N_2418);
nor U3506 (N_3506,N_2745,N_2734);
or U3507 (N_3507,N_2014,N_2685);
nor U3508 (N_3508,N_2030,N_2853);
nand U3509 (N_3509,N_2170,N_2805);
nor U3510 (N_3510,N_2715,N_2804);
nor U3511 (N_3511,N_2479,N_2836);
nor U3512 (N_3512,N_2642,N_2774);
nor U3513 (N_3513,N_2123,N_2776);
nand U3514 (N_3514,N_2077,N_2183);
xor U3515 (N_3515,N_2901,N_2957);
and U3516 (N_3516,N_2318,N_2662);
or U3517 (N_3517,N_2657,N_2988);
and U3518 (N_3518,N_2068,N_2131);
nor U3519 (N_3519,N_2391,N_2358);
nor U3520 (N_3520,N_2320,N_2170);
or U3521 (N_3521,N_2568,N_2901);
and U3522 (N_3522,N_2639,N_2189);
xor U3523 (N_3523,N_2650,N_2276);
xnor U3524 (N_3524,N_2231,N_2168);
or U3525 (N_3525,N_2341,N_2456);
and U3526 (N_3526,N_2706,N_2914);
or U3527 (N_3527,N_2100,N_2311);
or U3528 (N_3528,N_2237,N_2256);
nor U3529 (N_3529,N_2731,N_2825);
or U3530 (N_3530,N_2183,N_2876);
or U3531 (N_3531,N_2653,N_2711);
nand U3532 (N_3532,N_2506,N_2563);
or U3533 (N_3533,N_2283,N_2675);
or U3534 (N_3534,N_2652,N_2952);
and U3535 (N_3535,N_2422,N_2837);
and U3536 (N_3536,N_2963,N_2791);
xor U3537 (N_3537,N_2856,N_2670);
xnor U3538 (N_3538,N_2851,N_2861);
xnor U3539 (N_3539,N_2295,N_2512);
and U3540 (N_3540,N_2442,N_2660);
nand U3541 (N_3541,N_2513,N_2833);
and U3542 (N_3542,N_2609,N_2248);
nor U3543 (N_3543,N_2159,N_2809);
nand U3544 (N_3544,N_2840,N_2692);
nand U3545 (N_3545,N_2264,N_2537);
or U3546 (N_3546,N_2141,N_2342);
xnor U3547 (N_3547,N_2027,N_2146);
nor U3548 (N_3548,N_2252,N_2551);
or U3549 (N_3549,N_2567,N_2823);
xnor U3550 (N_3550,N_2786,N_2118);
and U3551 (N_3551,N_2595,N_2683);
nand U3552 (N_3552,N_2533,N_2876);
or U3553 (N_3553,N_2713,N_2107);
and U3554 (N_3554,N_2515,N_2740);
xor U3555 (N_3555,N_2445,N_2008);
nand U3556 (N_3556,N_2048,N_2571);
nor U3557 (N_3557,N_2259,N_2027);
nand U3558 (N_3558,N_2874,N_2822);
and U3559 (N_3559,N_2689,N_2072);
nor U3560 (N_3560,N_2102,N_2215);
nand U3561 (N_3561,N_2021,N_2730);
nor U3562 (N_3562,N_2462,N_2350);
nor U3563 (N_3563,N_2317,N_2019);
nand U3564 (N_3564,N_2466,N_2524);
nor U3565 (N_3565,N_2777,N_2653);
nor U3566 (N_3566,N_2435,N_2003);
xor U3567 (N_3567,N_2765,N_2255);
nand U3568 (N_3568,N_2024,N_2861);
xor U3569 (N_3569,N_2235,N_2003);
or U3570 (N_3570,N_2116,N_2975);
or U3571 (N_3571,N_2954,N_2402);
nand U3572 (N_3572,N_2878,N_2943);
or U3573 (N_3573,N_2600,N_2288);
nand U3574 (N_3574,N_2115,N_2740);
and U3575 (N_3575,N_2257,N_2745);
nand U3576 (N_3576,N_2744,N_2242);
or U3577 (N_3577,N_2461,N_2228);
and U3578 (N_3578,N_2364,N_2993);
nor U3579 (N_3579,N_2651,N_2342);
or U3580 (N_3580,N_2399,N_2279);
xor U3581 (N_3581,N_2539,N_2449);
nor U3582 (N_3582,N_2871,N_2845);
or U3583 (N_3583,N_2912,N_2328);
and U3584 (N_3584,N_2715,N_2419);
nor U3585 (N_3585,N_2668,N_2794);
and U3586 (N_3586,N_2509,N_2197);
nand U3587 (N_3587,N_2577,N_2394);
xor U3588 (N_3588,N_2300,N_2982);
nor U3589 (N_3589,N_2346,N_2322);
or U3590 (N_3590,N_2112,N_2060);
xnor U3591 (N_3591,N_2171,N_2308);
or U3592 (N_3592,N_2681,N_2642);
and U3593 (N_3593,N_2191,N_2417);
nand U3594 (N_3594,N_2726,N_2593);
and U3595 (N_3595,N_2108,N_2840);
nor U3596 (N_3596,N_2063,N_2689);
nor U3597 (N_3597,N_2151,N_2492);
xnor U3598 (N_3598,N_2587,N_2952);
nor U3599 (N_3599,N_2922,N_2155);
nor U3600 (N_3600,N_2192,N_2577);
nand U3601 (N_3601,N_2948,N_2801);
or U3602 (N_3602,N_2013,N_2664);
nand U3603 (N_3603,N_2300,N_2921);
or U3604 (N_3604,N_2098,N_2449);
or U3605 (N_3605,N_2769,N_2820);
nand U3606 (N_3606,N_2542,N_2964);
nor U3607 (N_3607,N_2482,N_2180);
nand U3608 (N_3608,N_2809,N_2377);
nand U3609 (N_3609,N_2824,N_2847);
nand U3610 (N_3610,N_2182,N_2714);
or U3611 (N_3611,N_2112,N_2814);
xor U3612 (N_3612,N_2211,N_2052);
and U3613 (N_3613,N_2766,N_2030);
nand U3614 (N_3614,N_2541,N_2310);
nand U3615 (N_3615,N_2578,N_2351);
nand U3616 (N_3616,N_2858,N_2934);
xnor U3617 (N_3617,N_2479,N_2254);
or U3618 (N_3618,N_2802,N_2979);
nor U3619 (N_3619,N_2643,N_2696);
and U3620 (N_3620,N_2478,N_2759);
xor U3621 (N_3621,N_2046,N_2740);
nand U3622 (N_3622,N_2774,N_2237);
and U3623 (N_3623,N_2832,N_2744);
nand U3624 (N_3624,N_2538,N_2580);
nand U3625 (N_3625,N_2406,N_2165);
xnor U3626 (N_3626,N_2472,N_2862);
nand U3627 (N_3627,N_2024,N_2732);
xor U3628 (N_3628,N_2350,N_2202);
xor U3629 (N_3629,N_2605,N_2645);
and U3630 (N_3630,N_2496,N_2926);
and U3631 (N_3631,N_2061,N_2739);
or U3632 (N_3632,N_2920,N_2500);
and U3633 (N_3633,N_2827,N_2056);
nor U3634 (N_3634,N_2651,N_2480);
nand U3635 (N_3635,N_2310,N_2059);
or U3636 (N_3636,N_2096,N_2894);
nand U3637 (N_3637,N_2654,N_2414);
xor U3638 (N_3638,N_2788,N_2606);
nand U3639 (N_3639,N_2855,N_2382);
or U3640 (N_3640,N_2283,N_2734);
nor U3641 (N_3641,N_2701,N_2985);
or U3642 (N_3642,N_2582,N_2828);
xor U3643 (N_3643,N_2593,N_2004);
xor U3644 (N_3644,N_2898,N_2919);
or U3645 (N_3645,N_2331,N_2253);
and U3646 (N_3646,N_2837,N_2183);
and U3647 (N_3647,N_2887,N_2423);
nor U3648 (N_3648,N_2120,N_2483);
and U3649 (N_3649,N_2626,N_2729);
nor U3650 (N_3650,N_2175,N_2467);
or U3651 (N_3651,N_2476,N_2740);
xnor U3652 (N_3652,N_2319,N_2485);
and U3653 (N_3653,N_2721,N_2273);
nor U3654 (N_3654,N_2169,N_2744);
and U3655 (N_3655,N_2574,N_2646);
nor U3656 (N_3656,N_2148,N_2392);
nor U3657 (N_3657,N_2615,N_2499);
xnor U3658 (N_3658,N_2106,N_2153);
nand U3659 (N_3659,N_2598,N_2935);
nand U3660 (N_3660,N_2427,N_2728);
nor U3661 (N_3661,N_2878,N_2476);
and U3662 (N_3662,N_2619,N_2857);
and U3663 (N_3663,N_2288,N_2848);
and U3664 (N_3664,N_2461,N_2772);
xor U3665 (N_3665,N_2451,N_2800);
xnor U3666 (N_3666,N_2398,N_2868);
or U3667 (N_3667,N_2002,N_2597);
and U3668 (N_3668,N_2302,N_2511);
nor U3669 (N_3669,N_2108,N_2428);
xor U3670 (N_3670,N_2323,N_2781);
and U3671 (N_3671,N_2659,N_2968);
or U3672 (N_3672,N_2155,N_2117);
and U3673 (N_3673,N_2016,N_2059);
nand U3674 (N_3674,N_2308,N_2443);
and U3675 (N_3675,N_2627,N_2896);
nand U3676 (N_3676,N_2453,N_2607);
and U3677 (N_3677,N_2997,N_2701);
or U3678 (N_3678,N_2346,N_2398);
or U3679 (N_3679,N_2676,N_2854);
xnor U3680 (N_3680,N_2537,N_2217);
nand U3681 (N_3681,N_2504,N_2172);
and U3682 (N_3682,N_2614,N_2788);
or U3683 (N_3683,N_2599,N_2988);
xnor U3684 (N_3684,N_2542,N_2859);
or U3685 (N_3685,N_2803,N_2781);
and U3686 (N_3686,N_2864,N_2170);
and U3687 (N_3687,N_2422,N_2723);
xor U3688 (N_3688,N_2626,N_2581);
nand U3689 (N_3689,N_2268,N_2797);
nor U3690 (N_3690,N_2717,N_2185);
xnor U3691 (N_3691,N_2292,N_2604);
or U3692 (N_3692,N_2582,N_2864);
or U3693 (N_3693,N_2512,N_2646);
xnor U3694 (N_3694,N_2506,N_2361);
xor U3695 (N_3695,N_2233,N_2250);
or U3696 (N_3696,N_2017,N_2735);
or U3697 (N_3697,N_2313,N_2212);
nand U3698 (N_3698,N_2348,N_2434);
or U3699 (N_3699,N_2778,N_2219);
xnor U3700 (N_3700,N_2793,N_2790);
and U3701 (N_3701,N_2994,N_2249);
xor U3702 (N_3702,N_2384,N_2247);
or U3703 (N_3703,N_2493,N_2251);
and U3704 (N_3704,N_2735,N_2570);
and U3705 (N_3705,N_2367,N_2625);
or U3706 (N_3706,N_2600,N_2768);
and U3707 (N_3707,N_2711,N_2058);
nand U3708 (N_3708,N_2720,N_2328);
or U3709 (N_3709,N_2355,N_2450);
or U3710 (N_3710,N_2836,N_2311);
xnor U3711 (N_3711,N_2285,N_2652);
or U3712 (N_3712,N_2936,N_2348);
nor U3713 (N_3713,N_2906,N_2909);
nand U3714 (N_3714,N_2505,N_2600);
xor U3715 (N_3715,N_2611,N_2767);
nor U3716 (N_3716,N_2953,N_2394);
nor U3717 (N_3717,N_2055,N_2841);
nor U3718 (N_3718,N_2227,N_2218);
nor U3719 (N_3719,N_2480,N_2726);
or U3720 (N_3720,N_2329,N_2499);
and U3721 (N_3721,N_2936,N_2449);
nand U3722 (N_3722,N_2180,N_2544);
and U3723 (N_3723,N_2647,N_2323);
or U3724 (N_3724,N_2847,N_2254);
and U3725 (N_3725,N_2416,N_2638);
and U3726 (N_3726,N_2836,N_2841);
nor U3727 (N_3727,N_2712,N_2722);
or U3728 (N_3728,N_2305,N_2756);
and U3729 (N_3729,N_2001,N_2776);
and U3730 (N_3730,N_2611,N_2300);
or U3731 (N_3731,N_2025,N_2183);
and U3732 (N_3732,N_2967,N_2503);
and U3733 (N_3733,N_2148,N_2897);
and U3734 (N_3734,N_2400,N_2589);
or U3735 (N_3735,N_2220,N_2745);
and U3736 (N_3736,N_2356,N_2550);
or U3737 (N_3737,N_2328,N_2322);
or U3738 (N_3738,N_2723,N_2951);
nor U3739 (N_3739,N_2295,N_2100);
or U3740 (N_3740,N_2110,N_2144);
or U3741 (N_3741,N_2371,N_2383);
or U3742 (N_3742,N_2444,N_2876);
nor U3743 (N_3743,N_2949,N_2091);
and U3744 (N_3744,N_2498,N_2205);
nand U3745 (N_3745,N_2807,N_2480);
nor U3746 (N_3746,N_2455,N_2092);
nand U3747 (N_3747,N_2122,N_2745);
xnor U3748 (N_3748,N_2343,N_2139);
nand U3749 (N_3749,N_2321,N_2225);
xor U3750 (N_3750,N_2018,N_2151);
and U3751 (N_3751,N_2703,N_2362);
or U3752 (N_3752,N_2714,N_2201);
or U3753 (N_3753,N_2403,N_2203);
xor U3754 (N_3754,N_2704,N_2320);
nand U3755 (N_3755,N_2671,N_2439);
xnor U3756 (N_3756,N_2931,N_2736);
xnor U3757 (N_3757,N_2420,N_2368);
and U3758 (N_3758,N_2601,N_2726);
xnor U3759 (N_3759,N_2764,N_2050);
and U3760 (N_3760,N_2970,N_2048);
nand U3761 (N_3761,N_2151,N_2010);
xnor U3762 (N_3762,N_2625,N_2641);
nand U3763 (N_3763,N_2080,N_2121);
or U3764 (N_3764,N_2392,N_2276);
or U3765 (N_3765,N_2801,N_2510);
nor U3766 (N_3766,N_2468,N_2205);
and U3767 (N_3767,N_2619,N_2480);
xor U3768 (N_3768,N_2981,N_2204);
xor U3769 (N_3769,N_2819,N_2702);
nand U3770 (N_3770,N_2956,N_2998);
and U3771 (N_3771,N_2792,N_2403);
nor U3772 (N_3772,N_2008,N_2600);
or U3773 (N_3773,N_2043,N_2360);
nand U3774 (N_3774,N_2343,N_2260);
or U3775 (N_3775,N_2300,N_2168);
and U3776 (N_3776,N_2595,N_2032);
nor U3777 (N_3777,N_2370,N_2087);
and U3778 (N_3778,N_2563,N_2188);
xnor U3779 (N_3779,N_2671,N_2124);
and U3780 (N_3780,N_2094,N_2052);
and U3781 (N_3781,N_2462,N_2652);
and U3782 (N_3782,N_2637,N_2815);
nand U3783 (N_3783,N_2822,N_2878);
xnor U3784 (N_3784,N_2005,N_2530);
nor U3785 (N_3785,N_2807,N_2199);
nor U3786 (N_3786,N_2222,N_2141);
nor U3787 (N_3787,N_2558,N_2281);
or U3788 (N_3788,N_2215,N_2882);
or U3789 (N_3789,N_2681,N_2311);
nor U3790 (N_3790,N_2916,N_2299);
xor U3791 (N_3791,N_2254,N_2813);
or U3792 (N_3792,N_2755,N_2595);
xor U3793 (N_3793,N_2046,N_2217);
nor U3794 (N_3794,N_2754,N_2325);
xor U3795 (N_3795,N_2185,N_2008);
or U3796 (N_3796,N_2145,N_2506);
nor U3797 (N_3797,N_2378,N_2176);
nor U3798 (N_3798,N_2683,N_2994);
or U3799 (N_3799,N_2512,N_2513);
nor U3800 (N_3800,N_2619,N_2655);
nor U3801 (N_3801,N_2534,N_2936);
nor U3802 (N_3802,N_2764,N_2390);
nor U3803 (N_3803,N_2626,N_2358);
nor U3804 (N_3804,N_2856,N_2321);
nor U3805 (N_3805,N_2030,N_2419);
nand U3806 (N_3806,N_2077,N_2881);
nor U3807 (N_3807,N_2477,N_2485);
nor U3808 (N_3808,N_2428,N_2673);
nor U3809 (N_3809,N_2496,N_2781);
or U3810 (N_3810,N_2833,N_2979);
or U3811 (N_3811,N_2755,N_2654);
xnor U3812 (N_3812,N_2880,N_2404);
nor U3813 (N_3813,N_2065,N_2253);
xor U3814 (N_3814,N_2682,N_2181);
nand U3815 (N_3815,N_2936,N_2049);
and U3816 (N_3816,N_2536,N_2628);
and U3817 (N_3817,N_2582,N_2981);
nor U3818 (N_3818,N_2782,N_2804);
xor U3819 (N_3819,N_2899,N_2538);
and U3820 (N_3820,N_2501,N_2088);
and U3821 (N_3821,N_2428,N_2214);
xnor U3822 (N_3822,N_2218,N_2007);
nor U3823 (N_3823,N_2362,N_2685);
or U3824 (N_3824,N_2375,N_2915);
xor U3825 (N_3825,N_2021,N_2916);
nor U3826 (N_3826,N_2302,N_2264);
and U3827 (N_3827,N_2022,N_2890);
nand U3828 (N_3828,N_2712,N_2214);
and U3829 (N_3829,N_2235,N_2556);
and U3830 (N_3830,N_2903,N_2855);
or U3831 (N_3831,N_2192,N_2176);
nand U3832 (N_3832,N_2897,N_2893);
nand U3833 (N_3833,N_2221,N_2702);
nand U3834 (N_3834,N_2071,N_2529);
or U3835 (N_3835,N_2374,N_2804);
or U3836 (N_3836,N_2508,N_2322);
nor U3837 (N_3837,N_2283,N_2942);
nand U3838 (N_3838,N_2979,N_2261);
xnor U3839 (N_3839,N_2995,N_2394);
nand U3840 (N_3840,N_2783,N_2920);
nor U3841 (N_3841,N_2952,N_2497);
and U3842 (N_3842,N_2176,N_2026);
nand U3843 (N_3843,N_2898,N_2218);
or U3844 (N_3844,N_2174,N_2141);
nand U3845 (N_3845,N_2587,N_2712);
xor U3846 (N_3846,N_2003,N_2707);
or U3847 (N_3847,N_2496,N_2865);
and U3848 (N_3848,N_2236,N_2461);
or U3849 (N_3849,N_2222,N_2637);
or U3850 (N_3850,N_2329,N_2712);
and U3851 (N_3851,N_2021,N_2172);
nand U3852 (N_3852,N_2198,N_2176);
and U3853 (N_3853,N_2203,N_2914);
nor U3854 (N_3854,N_2932,N_2416);
and U3855 (N_3855,N_2436,N_2689);
nor U3856 (N_3856,N_2868,N_2374);
nor U3857 (N_3857,N_2709,N_2153);
or U3858 (N_3858,N_2991,N_2588);
nor U3859 (N_3859,N_2812,N_2486);
nand U3860 (N_3860,N_2787,N_2716);
nor U3861 (N_3861,N_2640,N_2505);
nand U3862 (N_3862,N_2894,N_2713);
and U3863 (N_3863,N_2969,N_2103);
and U3864 (N_3864,N_2354,N_2408);
or U3865 (N_3865,N_2111,N_2726);
nand U3866 (N_3866,N_2362,N_2307);
xor U3867 (N_3867,N_2244,N_2772);
nor U3868 (N_3868,N_2373,N_2212);
nand U3869 (N_3869,N_2410,N_2885);
and U3870 (N_3870,N_2213,N_2355);
nor U3871 (N_3871,N_2366,N_2420);
and U3872 (N_3872,N_2216,N_2292);
and U3873 (N_3873,N_2778,N_2258);
or U3874 (N_3874,N_2010,N_2941);
xor U3875 (N_3875,N_2042,N_2078);
and U3876 (N_3876,N_2314,N_2230);
or U3877 (N_3877,N_2082,N_2331);
nor U3878 (N_3878,N_2157,N_2870);
nor U3879 (N_3879,N_2071,N_2478);
nor U3880 (N_3880,N_2057,N_2217);
nand U3881 (N_3881,N_2030,N_2643);
or U3882 (N_3882,N_2725,N_2504);
xnor U3883 (N_3883,N_2040,N_2615);
or U3884 (N_3884,N_2686,N_2464);
xor U3885 (N_3885,N_2841,N_2081);
nand U3886 (N_3886,N_2781,N_2438);
nand U3887 (N_3887,N_2717,N_2823);
or U3888 (N_3888,N_2768,N_2173);
nor U3889 (N_3889,N_2073,N_2577);
and U3890 (N_3890,N_2223,N_2933);
nor U3891 (N_3891,N_2669,N_2861);
and U3892 (N_3892,N_2392,N_2348);
and U3893 (N_3893,N_2765,N_2496);
and U3894 (N_3894,N_2561,N_2323);
nor U3895 (N_3895,N_2289,N_2086);
nand U3896 (N_3896,N_2722,N_2270);
nand U3897 (N_3897,N_2108,N_2075);
nand U3898 (N_3898,N_2088,N_2173);
or U3899 (N_3899,N_2228,N_2393);
nor U3900 (N_3900,N_2240,N_2188);
or U3901 (N_3901,N_2435,N_2379);
xor U3902 (N_3902,N_2524,N_2334);
nand U3903 (N_3903,N_2465,N_2197);
nand U3904 (N_3904,N_2816,N_2901);
and U3905 (N_3905,N_2692,N_2514);
and U3906 (N_3906,N_2966,N_2492);
and U3907 (N_3907,N_2860,N_2266);
nor U3908 (N_3908,N_2213,N_2260);
xor U3909 (N_3909,N_2873,N_2213);
and U3910 (N_3910,N_2209,N_2863);
nand U3911 (N_3911,N_2206,N_2957);
nand U3912 (N_3912,N_2757,N_2880);
nor U3913 (N_3913,N_2803,N_2411);
nand U3914 (N_3914,N_2830,N_2920);
nor U3915 (N_3915,N_2146,N_2783);
or U3916 (N_3916,N_2788,N_2323);
or U3917 (N_3917,N_2722,N_2785);
xnor U3918 (N_3918,N_2489,N_2021);
nand U3919 (N_3919,N_2688,N_2631);
nand U3920 (N_3920,N_2141,N_2870);
nand U3921 (N_3921,N_2593,N_2219);
xor U3922 (N_3922,N_2016,N_2480);
nor U3923 (N_3923,N_2413,N_2452);
and U3924 (N_3924,N_2373,N_2903);
and U3925 (N_3925,N_2175,N_2905);
and U3926 (N_3926,N_2835,N_2771);
or U3927 (N_3927,N_2099,N_2848);
nand U3928 (N_3928,N_2623,N_2341);
nand U3929 (N_3929,N_2981,N_2453);
nand U3930 (N_3930,N_2364,N_2260);
nand U3931 (N_3931,N_2992,N_2309);
nor U3932 (N_3932,N_2372,N_2773);
nand U3933 (N_3933,N_2129,N_2012);
or U3934 (N_3934,N_2966,N_2211);
or U3935 (N_3935,N_2780,N_2028);
nor U3936 (N_3936,N_2049,N_2376);
nor U3937 (N_3937,N_2613,N_2571);
or U3938 (N_3938,N_2389,N_2794);
nand U3939 (N_3939,N_2511,N_2549);
or U3940 (N_3940,N_2419,N_2474);
nand U3941 (N_3941,N_2609,N_2478);
xor U3942 (N_3942,N_2486,N_2271);
or U3943 (N_3943,N_2226,N_2450);
nor U3944 (N_3944,N_2805,N_2328);
xor U3945 (N_3945,N_2347,N_2091);
or U3946 (N_3946,N_2993,N_2833);
nand U3947 (N_3947,N_2460,N_2507);
nand U3948 (N_3948,N_2683,N_2285);
xor U3949 (N_3949,N_2154,N_2730);
and U3950 (N_3950,N_2215,N_2638);
xor U3951 (N_3951,N_2713,N_2290);
nor U3952 (N_3952,N_2296,N_2946);
nor U3953 (N_3953,N_2391,N_2111);
or U3954 (N_3954,N_2030,N_2816);
xor U3955 (N_3955,N_2458,N_2266);
xor U3956 (N_3956,N_2922,N_2703);
nand U3957 (N_3957,N_2779,N_2805);
and U3958 (N_3958,N_2088,N_2729);
xnor U3959 (N_3959,N_2979,N_2930);
nand U3960 (N_3960,N_2709,N_2600);
and U3961 (N_3961,N_2506,N_2837);
nand U3962 (N_3962,N_2440,N_2816);
nor U3963 (N_3963,N_2697,N_2663);
nor U3964 (N_3964,N_2452,N_2669);
and U3965 (N_3965,N_2100,N_2810);
nor U3966 (N_3966,N_2915,N_2413);
nor U3967 (N_3967,N_2041,N_2381);
and U3968 (N_3968,N_2405,N_2012);
or U3969 (N_3969,N_2991,N_2982);
nor U3970 (N_3970,N_2205,N_2418);
xor U3971 (N_3971,N_2236,N_2743);
xor U3972 (N_3972,N_2679,N_2471);
nand U3973 (N_3973,N_2550,N_2542);
nor U3974 (N_3974,N_2049,N_2337);
xor U3975 (N_3975,N_2329,N_2336);
or U3976 (N_3976,N_2130,N_2554);
and U3977 (N_3977,N_2747,N_2883);
xor U3978 (N_3978,N_2327,N_2448);
xor U3979 (N_3979,N_2453,N_2339);
nor U3980 (N_3980,N_2464,N_2546);
xnor U3981 (N_3981,N_2423,N_2470);
nand U3982 (N_3982,N_2974,N_2522);
and U3983 (N_3983,N_2729,N_2286);
or U3984 (N_3984,N_2411,N_2007);
nor U3985 (N_3985,N_2662,N_2483);
nand U3986 (N_3986,N_2343,N_2657);
xor U3987 (N_3987,N_2443,N_2713);
and U3988 (N_3988,N_2757,N_2952);
or U3989 (N_3989,N_2001,N_2959);
nor U3990 (N_3990,N_2779,N_2532);
or U3991 (N_3991,N_2126,N_2331);
nand U3992 (N_3992,N_2648,N_2820);
or U3993 (N_3993,N_2111,N_2871);
and U3994 (N_3994,N_2922,N_2787);
nand U3995 (N_3995,N_2895,N_2745);
nor U3996 (N_3996,N_2519,N_2132);
nor U3997 (N_3997,N_2501,N_2347);
and U3998 (N_3998,N_2523,N_2855);
nor U3999 (N_3999,N_2447,N_2283);
nor U4000 (N_4000,N_3214,N_3219);
or U4001 (N_4001,N_3687,N_3993);
nand U4002 (N_4002,N_3288,N_3978);
or U4003 (N_4003,N_3135,N_3611);
and U4004 (N_4004,N_3195,N_3765);
or U4005 (N_4005,N_3380,N_3351);
or U4006 (N_4006,N_3273,N_3137);
and U4007 (N_4007,N_3524,N_3951);
nand U4008 (N_4008,N_3349,N_3182);
xor U4009 (N_4009,N_3651,N_3234);
and U4010 (N_4010,N_3863,N_3431);
and U4011 (N_4011,N_3790,N_3718);
nand U4012 (N_4012,N_3448,N_3064);
nor U4013 (N_4013,N_3659,N_3079);
xnor U4014 (N_4014,N_3158,N_3539);
xor U4015 (N_4015,N_3062,N_3484);
xor U4016 (N_4016,N_3245,N_3266);
nand U4017 (N_4017,N_3289,N_3996);
and U4018 (N_4018,N_3468,N_3056);
nand U4019 (N_4019,N_3393,N_3053);
xnor U4020 (N_4020,N_3039,N_3426);
or U4021 (N_4021,N_3155,N_3577);
xor U4022 (N_4022,N_3824,N_3196);
and U4023 (N_4023,N_3989,N_3973);
nor U4024 (N_4024,N_3004,N_3507);
nor U4025 (N_4025,N_3425,N_3136);
xnor U4026 (N_4026,N_3419,N_3726);
or U4027 (N_4027,N_3304,N_3040);
xor U4028 (N_4028,N_3164,N_3736);
xnor U4029 (N_4029,N_3814,N_3059);
nor U4030 (N_4030,N_3140,N_3959);
xnor U4031 (N_4031,N_3485,N_3202);
xor U4032 (N_4032,N_3506,N_3181);
xor U4033 (N_4033,N_3027,N_3057);
nor U4034 (N_4034,N_3638,N_3386);
nand U4035 (N_4035,N_3769,N_3329);
or U4036 (N_4036,N_3678,N_3646);
xor U4037 (N_4037,N_3543,N_3576);
nor U4038 (N_4038,N_3744,N_3738);
nand U4039 (N_4039,N_3885,N_3003);
and U4040 (N_4040,N_3836,N_3120);
or U4041 (N_4041,N_3067,N_3495);
xnor U4042 (N_4042,N_3110,N_3170);
and U4043 (N_4043,N_3821,N_3267);
or U4044 (N_4044,N_3392,N_3982);
nor U4045 (N_4045,N_3190,N_3819);
nor U4046 (N_4046,N_3389,N_3369);
and U4047 (N_4047,N_3604,N_3911);
xnor U4048 (N_4048,N_3566,N_3330);
or U4049 (N_4049,N_3966,N_3893);
xor U4050 (N_4050,N_3034,N_3250);
xor U4051 (N_4051,N_3331,N_3674);
nor U4052 (N_4052,N_3068,N_3645);
and U4053 (N_4053,N_3222,N_3071);
and U4054 (N_4054,N_3035,N_3435);
xor U4055 (N_4055,N_3969,N_3152);
nor U4056 (N_4056,N_3588,N_3513);
or U4057 (N_4057,N_3694,N_3984);
nor U4058 (N_4058,N_3860,N_3256);
nand U4059 (N_4059,N_3361,N_3009);
nand U4060 (N_4060,N_3381,N_3442);
or U4061 (N_4061,N_3301,N_3953);
nand U4062 (N_4062,N_3342,N_3773);
xnor U4063 (N_4063,N_3391,N_3334);
and U4064 (N_4064,N_3707,N_3394);
nor U4065 (N_4065,N_3755,N_3218);
nor U4066 (N_4066,N_3197,N_3227);
and U4067 (N_4067,N_3698,N_3584);
and U4068 (N_4068,N_3449,N_3208);
nor U4069 (N_4069,N_3859,N_3985);
nand U4070 (N_4070,N_3261,N_3931);
xor U4071 (N_4071,N_3338,N_3173);
and U4072 (N_4072,N_3591,N_3574);
nor U4073 (N_4073,N_3141,N_3221);
xnor U4074 (N_4074,N_3533,N_3921);
nand U4075 (N_4075,N_3917,N_3127);
nand U4076 (N_4076,N_3815,N_3326);
xor U4077 (N_4077,N_3630,N_3060);
nor U4078 (N_4078,N_3168,N_3232);
xor U4079 (N_4079,N_3246,N_3474);
and U4080 (N_4080,N_3555,N_3276);
or U4081 (N_4081,N_3797,N_3876);
xor U4082 (N_4082,N_3470,N_3480);
nand U4083 (N_4083,N_3534,N_3831);
nor U4084 (N_4084,N_3722,N_3999);
nor U4085 (N_4085,N_3800,N_3430);
and U4086 (N_4086,N_3567,N_3293);
nand U4087 (N_4087,N_3725,N_3306);
xor U4088 (N_4088,N_3408,N_3240);
or U4089 (N_4089,N_3749,N_3496);
or U4090 (N_4090,N_3285,N_3469);
xor U4091 (N_4091,N_3241,N_3945);
and U4092 (N_4092,N_3211,N_3699);
nor U4093 (N_4093,N_3016,N_3479);
nand U4094 (N_4094,N_3820,N_3542);
xor U4095 (N_4095,N_3676,N_3954);
nor U4096 (N_4096,N_3807,N_3090);
or U4097 (N_4097,N_3925,N_3082);
xor U4098 (N_4098,N_3462,N_3296);
nand U4099 (N_4099,N_3081,N_3672);
and U4100 (N_4100,N_3353,N_3465);
nor U4101 (N_4101,N_3872,N_3509);
nor U4102 (N_4102,N_3437,N_3541);
xnor U4103 (N_4103,N_3383,N_3160);
nand U4104 (N_4104,N_3049,N_3176);
nor U4105 (N_4105,N_3943,N_3179);
and U4106 (N_4106,N_3839,N_3500);
or U4107 (N_4107,N_3995,N_3157);
and U4108 (N_4108,N_3516,N_3663);
nand U4109 (N_4109,N_3786,N_3990);
nor U4110 (N_4110,N_3362,N_3230);
nor U4111 (N_4111,N_3713,N_3705);
nand U4112 (N_4112,N_3554,N_3680);
xor U4113 (N_4113,N_3413,N_3048);
and U4114 (N_4114,N_3602,N_3434);
and U4115 (N_4115,N_3387,N_3411);
nand U4116 (N_4116,N_3036,N_3545);
xor U4117 (N_4117,N_3011,N_3601);
xor U4118 (N_4118,N_3624,N_3249);
or U4119 (N_4119,N_3758,N_3453);
or U4120 (N_4120,N_3668,N_3318);
nand U4121 (N_4121,N_3855,N_3649);
nand U4122 (N_4122,N_3111,N_3108);
and U4123 (N_4123,N_3540,N_3258);
nand U4124 (N_4124,N_3089,N_3078);
xnor U4125 (N_4125,N_3028,N_3882);
or U4126 (N_4126,N_3096,N_3637);
xor U4127 (N_4127,N_3086,N_3756);
nand U4128 (N_4128,N_3263,N_3433);
xnor U4129 (N_4129,N_3374,N_3851);
nor U4130 (N_4130,N_3432,N_3766);
nor U4131 (N_4131,N_3950,N_3400);
and U4132 (N_4132,N_3847,N_3948);
or U4133 (N_4133,N_3771,N_3938);
or U4134 (N_4134,N_3279,N_3018);
xor U4135 (N_4135,N_3906,N_3148);
nor U4136 (N_4136,N_3956,N_3916);
xnor U4137 (N_4137,N_3551,N_3890);
nand U4138 (N_4138,N_3874,N_3185);
and U4139 (N_4139,N_3311,N_3023);
xnor U4140 (N_4140,N_3000,N_3941);
or U4141 (N_4141,N_3401,N_3706);
nand U4142 (N_4142,N_3104,N_3147);
or U4143 (N_4143,N_3026,N_3073);
or U4144 (N_4144,N_3428,N_3121);
and U4145 (N_4145,N_3704,N_3372);
and U4146 (N_4146,N_3243,N_3528);
nand U4147 (N_4147,N_3128,N_3379);
xnor U4148 (N_4148,N_3849,N_3535);
xnor U4149 (N_4149,N_3325,N_3633);
nor U4150 (N_4150,N_3805,N_3050);
xor U4151 (N_4151,N_3677,N_3970);
nor U4152 (N_4152,N_3563,N_3124);
and U4153 (N_4153,N_3344,N_3452);
and U4154 (N_4154,N_3614,N_3251);
nor U4155 (N_4155,N_3536,N_3519);
nand U4156 (N_4156,N_3711,N_3366);
nand U4157 (N_4157,N_3730,N_3998);
xnor U4158 (N_4158,N_3910,N_3122);
or U4159 (N_4159,N_3787,N_3627);
or U4160 (N_4160,N_3686,N_3986);
nor U4161 (N_4161,N_3742,N_3348);
nor U4162 (N_4162,N_3568,N_3459);
nor U4163 (N_4163,N_3504,N_3570);
nand U4164 (N_4164,N_3940,N_3826);
and U4165 (N_4165,N_3818,N_3076);
and U4166 (N_4166,N_3467,N_3530);
and U4167 (N_4167,N_3572,N_3414);
nor U4168 (N_4168,N_3134,N_3088);
or U4169 (N_4169,N_3520,N_3537);
nand U4170 (N_4170,N_3547,N_3006);
and U4171 (N_4171,N_3092,N_3345);
or U4172 (N_4172,N_3697,N_3192);
or U4173 (N_4173,N_3375,N_3102);
nand U4174 (N_4174,N_3650,N_3517);
xor U4175 (N_4175,N_3239,N_3721);
and U4176 (N_4176,N_3660,N_3903);
and U4177 (N_4177,N_3981,N_3367);
xnor U4178 (N_4178,N_3901,N_3904);
nor U4179 (N_4179,N_3983,N_3729);
xnor U4180 (N_4180,N_3487,N_3852);
xnor U4181 (N_4181,N_3866,N_3184);
or U4182 (N_4182,N_3052,N_3175);
nand U4183 (N_4183,N_3363,N_3264);
nand U4184 (N_4184,N_3189,N_3094);
and U4185 (N_4185,N_3475,N_3946);
xor U4186 (N_4186,N_3673,N_3199);
and U4187 (N_4187,N_3881,N_3731);
xor U4188 (N_4188,N_3991,N_3955);
or U4189 (N_4189,N_3287,N_3971);
or U4190 (N_4190,N_3317,N_3780);
or U4191 (N_4191,N_3489,N_3277);
or U4192 (N_4192,N_3868,N_3690);
or U4193 (N_4193,N_3908,N_3929);
and U4194 (N_4194,N_3488,N_3320);
nand U4195 (N_4195,N_3324,N_3976);
nor U4196 (N_4196,N_3212,N_3781);
or U4197 (N_4197,N_3074,N_3303);
nor U4198 (N_4198,N_3887,N_3935);
or U4199 (N_4199,N_3870,N_3753);
or U4200 (N_4200,N_3119,N_3666);
xor U4201 (N_4201,N_3217,N_3879);
xnor U4202 (N_4202,N_3354,N_3132);
nor U4203 (N_4203,N_3912,N_3974);
or U4204 (N_4204,N_3445,N_3880);
or U4205 (N_4205,N_3799,N_3857);
and U4206 (N_4206,N_3965,N_3612);
or U4207 (N_4207,N_3639,N_3924);
nor U4208 (N_4208,N_3675,N_3759);
or U4209 (N_4209,N_3305,N_3272);
nor U4210 (N_4210,N_3606,N_3531);
xor U4211 (N_4211,N_3806,N_3733);
nand U4212 (N_4212,N_3429,N_3888);
nand U4213 (N_4213,N_3741,N_3194);
xnor U4214 (N_4214,N_3145,N_3077);
or U4215 (N_4215,N_3117,N_3237);
or U4216 (N_4216,N_3636,N_3174);
or U4217 (N_4217,N_3662,N_3171);
xnor U4218 (N_4218,N_3020,N_3936);
and U4219 (N_4219,N_3928,N_3803);
nor U4220 (N_4220,N_3198,N_3980);
nand U4221 (N_4221,N_3510,N_3270);
and U4222 (N_4222,N_3365,N_3856);
xor U4223 (N_4223,N_3746,N_3332);
and U4224 (N_4224,N_3385,N_3891);
nand U4225 (N_4225,N_3858,N_3492);
or U4226 (N_4226,N_3720,N_3456);
nand U4227 (N_4227,N_3233,N_3556);
or U4228 (N_4228,N_3752,N_3934);
nor U4229 (N_4229,N_3292,N_3669);
and U4230 (N_4230,N_3865,N_3631);
or U4231 (N_4231,N_3031,N_3047);
or U4232 (N_4232,N_3390,N_3407);
xnor U4233 (N_4233,N_3446,N_3255);
nor U4234 (N_4234,N_3187,N_3295);
xnor U4235 (N_4235,N_3244,N_3837);
nor U4236 (N_4236,N_3364,N_3963);
nor U4237 (N_4237,N_3768,N_3165);
and U4238 (N_4238,N_3822,N_3493);
nand U4239 (N_4239,N_3024,N_3905);
xnor U4240 (N_4240,N_3420,N_3626);
or U4241 (N_4241,N_3617,N_3335);
nand U4242 (N_4242,N_3550,N_3439);
nand U4243 (N_4243,N_3037,N_3825);
nor U4244 (N_4244,N_3791,N_3377);
or U4245 (N_4245,N_3754,N_3061);
and U4246 (N_4246,N_3415,N_3511);
xor U4247 (N_4247,N_3340,N_3281);
and U4248 (N_4248,N_3840,N_3902);
nor U4249 (N_4249,N_3247,N_3975);
or U4250 (N_4250,N_3346,N_3914);
and U4251 (N_4251,N_3191,N_3892);
nor U4252 (N_4252,N_3564,N_3274);
nor U4253 (N_4253,N_3640,N_3615);
nand U4254 (N_4254,N_3087,N_3162);
or U4255 (N_4255,N_3313,N_3327);
nand U4256 (N_4256,N_3231,N_3853);
nor U4257 (N_4257,N_3683,N_3664);
or U4258 (N_4258,N_3682,N_3038);
nor U4259 (N_4259,N_3220,N_3977);
nand U4260 (N_4260,N_3154,N_3114);
nand U4261 (N_4261,N_3498,N_3225);
nor U4262 (N_4262,N_3322,N_3804);
xnor U4263 (N_4263,N_3412,N_3656);
xor U4264 (N_4264,N_3900,N_3581);
or U4265 (N_4265,N_3029,N_3850);
nor U4266 (N_4266,N_3228,N_3538);
nand U4267 (N_4267,N_3491,N_3188);
or U4268 (N_4268,N_3817,N_3101);
and U4269 (N_4269,N_3552,N_3599);
and U4270 (N_4270,N_3632,N_3253);
nor U4271 (N_4271,N_3607,N_3942);
or U4272 (N_4272,N_3869,N_3186);
nand U4273 (N_4273,N_3571,N_3129);
and U4274 (N_4274,N_3823,N_3947);
and U4275 (N_4275,N_3205,N_3788);
or U4276 (N_4276,N_3012,N_3514);
or U4277 (N_4277,N_3693,N_3590);
nand U4278 (N_4278,N_3871,N_3418);
and U4279 (N_4279,N_3080,N_3441);
or U4280 (N_4280,N_3569,N_3580);
nand U4281 (N_4281,N_3033,N_3177);
or U4282 (N_4282,N_3319,N_3298);
nand U4283 (N_4283,N_3629,N_3620);
nand U4284 (N_4284,N_3001,N_3653);
nand U4285 (N_4285,N_3703,N_3779);
nand U4286 (N_4286,N_3310,N_3490);
or U4287 (N_4287,N_3792,N_3183);
and U4288 (N_4288,N_3213,N_3200);
or U4289 (N_4289,N_3356,N_3565);
nor U4290 (N_4290,N_3688,N_3597);
or U4291 (N_4291,N_3618,N_3378);
or U4292 (N_4292,N_3045,N_3333);
xor U4293 (N_4293,N_3957,N_3770);
or U4294 (N_4294,N_3404,N_3579);
nand U4295 (N_4295,N_3151,N_3671);
xor U4296 (N_4296,N_3695,N_3696);
nor U4297 (N_4297,N_3605,N_3403);
and U4298 (N_4298,N_3907,N_3314);
nand U4299 (N_4299,N_3795,N_3278);
and U4300 (N_4300,N_3641,N_3161);
or U4301 (N_4301,N_3939,N_3778);
nand U4302 (N_4302,N_3523,N_3613);
nand U4303 (N_4303,N_3300,N_3979);
nor U4304 (N_4304,N_3867,N_3149);
nand U4305 (N_4305,N_3455,N_3497);
xor U4306 (N_4306,N_3458,N_3417);
or U4307 (N_4307,N_3472,N_3422);
or U4308 (N_4308,N_3229,N_3058);
nand U4309 (N_4309,N_3501,N_3784);
and U4310 (N_4310,N_3710,N_3235);
xnor U4311 (N_4311,N_3447,N_3041);
nor U4312 (N_4312,N_3546,N_3763);
and U4313 (N_4313,N_3384,N_3809);
and U4314 (N_4314,N_3846,N_3884);
xnor U4315 (N_4315,N_3421,N_3685);
nor U4316 (N_4316,N_3410,N_3125);
xor U4317 (N_4317,N_3548,N_3723);
nand U4318 (N_4318,N_3156,N_3084);
nor U4319 (N_4319,N_3665,N_3679);
or U4320 (N_4320,N_3962,N_3337);
xor U4321 (N_4321,N_3302,N_3451);
nand U4322 (N_4322,N_3987,N_3734);
xor U4323 (N_4323,N_3098,N_3883);
nand U4324 (N_4324,N_3248,N_3402);
nor U4325 (N_4325,N_3309,N_3864);
or U4326 (N_4326,N_3312,N_3926);
nand U4327 (N_4327,N_3476,N_3623);
or U4328 (N_4328,N_3262,N_3294);
nand U4329 (N_4329,N_3268,N_3478);
and U4330 (N_4330,N_3223,N_3586);
or U4331 (N_4331,N_3396,N_3575);
and U4332 (N_4332,N_3283,N_3359);
or U4333 (N_4333,N_3054,N_3163);
nand U4334 (N_4334,N_3347,N_3416);
xnor U4335 (N_4335,N_3600,N_3635);
nand U4336 (N_4336,N_3997,N_3099);
nand U4337 (N_4337,N_3700,N_3065);
nand U4338 (N_4338,N_3915,N_3242);
or U4339 (N_4339,N_3518,N_3178);
nand U4340 (N_4340,N_3502,N_3144);
nand U4341 (N_4341,N_3505,N_3106);
and U4342 (N_4342,N_3757,N_3275);
nor U4343 (N_4343,N_3561,N_3323);
nor U4344 (N_4344,N_3648,N_3461);
and U4345 (N_4345,N_3014,N_3861);
and U4346 (N_4346,N_3833,N_3463);
and U4347 (N_4347,N_3794,N_3595);
xor U4348 (N_4348,N_3097,N_3282);
nor U4349 (N_4349,N_3789,N_3207);
nor U4350 (N_4350,N_3260,N_3343);
nor U4351 (N_4351,N_3010,N_3109);
nor U4352 (N_4352,N_3002,N_3043);
nand U4353 (N_4353,N_3336,N_3589);
xnor U4354 (N_4354,N_3203,N_3745);
nand U4355 (N_4355,N_3471,N_3661);
nand U4356 (N_4356,N_3271,N_3886);
nor U4357 (N_4357,N_3210,N_3644);
and U4358 (N_4358,N_3952,N_3712);
and U4359 (N_4359,N_3832,N_3810);
nor U4360 (N_4360,N_3559,N_3438);
nand U4361 (N_4361,N_3069,N_3257);
nand U4362 (N_4362,N_3717,N_3732);
and U4363 (N_4363,N_3019,N_3215);
xor U4364 (N_4364,N_3499,N_3843);
nand U4365 (N_4365,N_3159,N_3521);
nand U4366 (N_4366,N_3008,N_3423);
or U4367 (N_4367,N_3044,N_3388);
nor U4368 (N_4368,N_3503,N_3206);
and U4369 (N_4369,N_3553,N_3055);
and U4370 (N_4370,N_3667,N_3204);
nand U4371 (N_4371,N_3582,N_3436);
and U4372 (N_4372,N_3767,N_3596);
nand U4373 (N_4373,N_3670,N_3005);
or U4374 (N_4374,N_3328,N_3922);
and U4375 (N_4375,N_3923,N_3297);
or U4376 (N_4376,N_3875,N_3284);
nand U4377 (N_4377,N_3466,N_3619);
or U4378 (N_4378,N_3838,N_3592);
and U4379 (N_4379,N_3025,N_3709);
nand U4380 (N_4380,N_3030,N_3444);
nand U4381 (N_4381,N_3142,N_3918);
or U4382 (N_4382,N_3116,N_3719);
xor U4383 (N_4383,N_3180,N_3046);
or U4384 (N_4384,N_3355,N_3813);
and U4385 (N_4385,N_3811,N_3269);
nand U4386 (N_4386,N_3842,N_3209);
or U4387 (N_4387,N_3793,N_3167);
nand U4388 (N_4388,N_3933,N_3802);
or U4389 (N_4389,N_3616,N_3944);
and U4390 (N_4390,N_3105,N_3932);
or U4391 (N_4391,N_3032,N_3238);
or U4392 (N_4392,N_3007,N_3796);
and U4393 (N_4393,N_3265,N_3315);
xnor U4394 (N_4394,N_3123,N_3558);
and U4395 (N_4395,N_3308,N_3015);
nand U4396 (N_4396,N_3608,N_3897);
nor U4397 (N_4397,N_3405,N_3424);
nand U4398 (N_4398,N_3785,N_3443);
xor U4399 (N_4399,N_3739,N_3621);
and U4400 (N_4400,N_3894,N_3481);
and U4401 (N_4401,N_3835,N_3828);
and U4402 (N_4402,N_3399,N_3406);
and U4403 (N_4403,N_3483,N_3370);
xnor U4404 (N_4404,N_3578,N_3095);
xnor U4405 (N_4405,N_3103,N_3013);
nor U4406 (N_4406,N_3172,N_3748);
nand U4407 (N_4407,N_3350,N_3913);
nor U4408 (N_4408,N_3681,N_3236);
nand U4409 (N_4409,N_3750,N_3609);
or U4410 (N_4410,N_3958,N_3658);
and U4411 (N_4411,N_3515,N_3702);
nand U4412 (N_4412,N_3358,N_3634);
nor U4413 (N_4413,N_3139,N_3085);
nand U4414 (N_4414,N_3512,N_3460);
or U4415 (N_4415,N_3532,N_3737);
or U4416 (N_4416,N_3728,N_3091);
nor U4417 (N_4417,N_3286,N_3150);
or U4418 (N_4418,N_3657,N_3307);
nor U4419 (N_4419,N_3066,N_3774);
xor U4420 (N_4420,N_3395,N_3254);
or U4421 (N_4421,N_3625,N_3642);
xor U4422 (N_4422,N_3964,N_3368);
nand U4423 (N_4423,N_3834,N_3259);
xnor U4424 (N_4424,N_3133,N_3409);
nand U4425 (N_4425,N_3854,N_3949);
and U4426 (N_4426,N_3454,N_3593);
nor U4427 (N_4427,N_3937,N_3961);
nand U4428 (N_4428,N_3022,N_3844);
nand U4429 (N_4429,N_3093,N_3341);
or U4430 (N_4430,N_3316,N_3761);
xnor U4431 (N_4431,N_3021,N_3777);
nand U4432 (N_4432,N_3126,N_3585);
and U4433 (N_4433,N_3226,N_3841);
xor U4434 (N_4434,N_3486,N_3689);
nor U4435 (N_4435,N_3224,N_3877);
or U4436 (N_4436,N_3587,N_3072);
nand U4437 (N_4437,N_3772,N_3115);
nand U4438 (N_4438,N_3549,N_3583);
and U4439 (N_4439,N_3622,N_3708);
xor U4440 (N_4440,N_3994,N_3930);
and U4441 (N_4441,N_3560,N_3684);
or U4442 (N_4442,N_3440,N_3830);
nor U4443 (N_4443,N_3113,N_3594);
nor U4444 (N_4444,N_3743,N_3715);
or U4445 (N_4445,N_3701,N_3130);
and U4446 (N_4446,N_3692,N_3373);
nand U4447 (N_4447,N_3522,N_3562);
and U4448 (N_4448,N_3654,N_3112);
nor U4449 (N_4449,N_3714,N_3398);
nor U4450 (N_4450,N_3357,N_3557);
nand U4451 (N_4451,N_3827,N_3727);
or U4452 (N_4452,N_3376,N_3339);
nor U4453 (N_4453,N_3967,N_3464);
xnor U4454 (N_4454,N_3482,N_3131);
or U4455 (N_4455,N_3927,N_3427);
nand U4456 (N_4456,N_3878,N_3473);
nand U4457 (N_4457,N_3138,N_3107);
nand U4458 (N_4458,N_3735,N_3808);
xor U4459 (N_4459,N_3382,N_3042);
and U4460 (N_4460,N_3166,N_3895);
nand U4461 (N_4461,N_3968,N_3747);
or U4462 (N_4462,N_3146,N_3873);
nor U4463 (N_4463,N_3252,N_3610);
nand U4464 (N_4464,N_3889,N_3691);
nand U4465 (N_4465,N_3760,N_3628);
xor U4466 (N_4466,N_3525,N_3494);
nand U4467 (N_4467,N_3816,N_3216);
or U4468 (N_4468,N_3193,N_3153);
and U4469 (N_4469,N_3201,N_3751);
nor U4470 (N_4470,N_3801,N_3477);
or U4471 (N_4471,N_3899,N_3764);
nor U4472 (N_4472,N_3291,N_3573);
xnor U4473 (N_4473,N_3508,N_3972);
nor U4474 (N_4474,N_3371,N_3299);
and U4475 (N_4475,N_3083,N_3526);
and U4476 (N_4476,N_3643,N_3775);
xor U4477 (N_4477,N_3598,N_3848);
or U4478 (N_4478,N_3100,N_3017);
xor U4479 (N_4479,N_3321,N_3740);
xnor U4480 (N_4480,N_3450,N_3070);
or U4481 (N_4481,N_3782,N_3920);
nand U4482 (N_4482,N_3724,N_3169);
or U4483 (N_4483,N_3960,N_3783);
nor U4484 (N_4484,N_3527,N_3352);
nor U4485 (N_4485,N_3812,N_3360);
nand U4486 (N_4486,N_3280,N_3397);
nand U4487 (N_4487,N_3063,N_3051);
xor U4488 (N_4488,N_3647,N_3988);
xor U4489 (N_4489,N_3798,N_3862);
or U4490 (N_4490,N_3919,N_3762);
and U4491 (N_4491,N_3143,N_3457);
or U4492 (N_4492,N_3716,N_3845);
and U4493 (N_4493,N_3829,N_3898);
nor U4494 (N_4494,N_3118,N_3776);
nor U4495 (N_4495,N_3529,N_3896);
nor U4496 (N_4496,N_3909,N_3603);
and U4497 (N_4497,N_3290,N_3655);
nand U4498 (N_4498,N_3544,N_3075);
nor U4499 (N_4499,N_3652,N_3992);
nand U4500 (N_4500,N_3308,N_3842);
and U4501 (N_4501,N_3291,N_3947);
nand U4502 (N_4502,N_3018,N_3546);
nand U4503 (N_4503,N_3945,N_3198);
nor U4504 (N_4504,N_3236,N_3241);
or U4505 (N_4505,N_3878,N_3800);
xor U4506 (N_4506,N_3552,N_3428);
nand U4507 (N_4507,N_3370,N_3059);
xor U4508 (N_4508,N_3158,N_3551);
xor U4509 (N_4509,N_3561,N_3775);
xor U4510 (N_4510,N_3813,N_3000);
xnor U4511 (N_4511,N_3449,N_3120);
nor U4512 (N_4512,N_3093,N_3495);
nor U4513 (N_4513,N_3991,N_3937);
and U4514 (N_4514,N_3772,N_3770);
xnor U4515 (N_4515,N_3357,N_3384);
and U4516 (N_4516,N_3484,N_3523);
or U4517 (N_4517,N_3781,N_3497);
and U4518 (N_4518,N_3424,N_3221);
or U4519 (N_4519,N_3511,N_3501);
nand U4520 (N_4520,N_3864,N_3983);
xnor U4521 (N_4521,N_3682,N_3710);
nand U4522 (N_4522,N_3887,N_3931);
and U4523 (N_4523,N_3641,N_3442);
xnor U4524 (N_4524,N_3506,N_3794);
xor U4525 (N_4525,N_3926,N_3795);
and U4526 (N_4526,N_3788,N_3488);
or U4527 (N_4527,N_3710,N_3050);
nor U4528 (N_4528,N_3144,N_3199);
and U4529 (N_4529,N_3719,N_3840);
and U4530 (N_4530,N_3044,N_3974);
xnor U4531 (N_4531,N_3462,N_3884);
xor U4532 (N_4532,N_3889,N_3747);
or U4533 (N_4533,N_3267,N_3120);
nand U4534 (N_4534,N_3713,N_3537);
nand U4535 (N_4535,N_3698,N_3192);
nor U4536 (N_4536,N_3001,N_3122);
nand U4537 (N_4537,N_3162,N_3118);
or U4538 (N_4538,N_3955,N_3387);
nand U4539 (N_4539,N_3995,N_3335);
and U4540 (N_4540,N_3232,N_3986);
xor U4541 (N_4541,N_3485,N_3399);
nor U4542 (N_4542,N_3280,N_3820);
nor U4543 (N_4543,N_3058,N_3035);
nor U4544 (N_4544,N_3251,N_3926);
xnor U4545 (N_4545,N_3659,N_3455);
and U4546 (N_4546,N_3251,N_3041);
or U4547 (N_4547,N_3947,N_3616);
or U4548 (N_4548,N_3292,N_3576);
or U4549 (N_4549,N_3705,N_3883);
or U4550 (N_4550,N_3336,N_3431);
xor U4551 (N_4551,N_3375,N_3206);
nand U4552 (N_4552,N_3796,N_3584);
nand U4553 (N_4553,N_3873,N_3159);
nand U4554 (N_4554,N_3211,N_3565);
nor U4555 (N_4555,N_3709,N_3846);
or U4556 (N_4556,N_3715,N_3180);
xor U4557 (N_4557,N_3944,N_3870);
nor U4558 (N_4558,N_3451,N_3307);
and U4559 (N_4559,N_3745,N_3711);
or U4560 (N_4560,N_3914,N_3220);
or U4561 (N_4561,N_3083,N_3620);
nand U4562 (N_4562,N_3919,N_3336);
nand U4563 (N_4563,N_3743,N_3644);
nor U4564 (N_4564,N_3849,N_3605);
and U4565 (N_4565,N_3212,N_3560);
nor U4566 (N_4566,N_3842,N_3175);
nand U4567 (N_4567,N_3918,N_3406);
nand U4568 (N_4568,N_3847,N_3300);
or U4569 (N_4569,N_3462,N_3694);
nor U4570 (N_4570,N_3380,N_3622);
nor U4571 (N_4571,N_3969,N_3185);
xnor U4572 (N_4572,N_3208,N_3458);
xor U4573 (N_4573,N_3037,N_3694);
or U4574 (N_4574,N_3639,N_3027);
and U4575 (N_4575,N_3792,N_3340);
nand U4576 (N_4576,N_3394,N_3855);
or U4577 (N_4577,N_3421,N_3176);
nor U4578 (N_4578,N_3105,N_3121);
nor U4579 (N_4579,N_3910,N_3094);
xnor U4580 (N_4580,N_3006,N_3958);
nand U4581 (N_4581,N_3058,N_3125);
or U4582 (N_4582,N_3147,N_3341);
and U4583 (N_4583,N_3458,N_3999);
xnor U4584 (N_4584,N_3563,N_3178);
or U4585 (N_4585,N_3800,N_3324);
and U4586 (N_4586,N_3134,N_3813);
xnor U4587 (N_4587,N_3448,N_3089);
nor U4588 (N_4588,N_3114,N_3442);
and U4589 (N_4589,N_3641,N_3814);
nor U4590 (N_4590,N_3340,N_3505);
xor U4591 (N_4591,N_3514,N_3596);
and U4592 (N_4592,N_3323,N_3175);
xor U4593 (N_4593,N_3025,N_3712);
xor U4594 (N_4594,N_3364,N_3999);
nand U4595 (N_4595,N_3549,N_3332);
nand U4596 (N_4596,N_3878,N_3198);
or U4597 (N_4597,N_3314,N_3179);
nand U4598 (N_4598,N_3367,N_3637);
nand U4599 (N_4599,N_3757,N_3772);
nand U4600 (N_4600,N_3424,N_3438);
nand U4601 (N_4601,N_3419,N_3356);
nor U4602 (N_4602,N_3444,N_3447);
and U4603 (N_4603,N_3503,N_3040);
nor U4604 (N_4604,N_3634,N_3911);
and U4605 (N_4605,N_3087,N_3880);
or U4606 (N_4606,N_3541,N_3401);
xor U4607 (N_4607,N_3859,N_3101);
or U4608 (N_4608,N_3656,N_3797);
xor U4609 (N_4609,N_3095,N_3907);
or U4610 (N_4610,N_3444,N_3286);
xor U4611 (N_4611,N_3899,N_3121);
or U4612 (N_4612,N_3688,N_3905);
xor U4613 (N_4613,N_3943,N_3125);
nand U4614 (N_4614,N_3033,N_3806);
or U4615 (N_4615,N_3607,N_3395);
nand U4616 (N_4616,N_3545,N_3138);
xnor U4617 (N_4617,N_3877,N_3527);
and U4618 (N_4618,N_3391,N_3375);
and U4619 (N_4619,N_3264,N_3710);
nor U4620 (N_4620,N_3809,N_3882);
nand U4621 (N_4621,N_3640,N_3759);
xor U4622 (N_4622,N_3402,N_3182);
or U4623 (N_4623,N_3417,N_3625);
or U4624 (N_4624,N_3589,N_3229);
xor U4625 (N_4625,N_3933,N_3964);
nand U4626 (N_4626,N_3258,N_3867);
xor U4627 (N_4627,N_3497,N_3126);
and U4628 (N_4628,N_3170,N_3863);
nand U4629 (N_4629,N_3041,N_3450);
nor U4630 (N_4630,N_3324,N_3957);
and U4631 (N_4631,N_3667,N_3838);
xor U4632 (N_4632,N_3137,N_3347);
or U4633 (N_4633,N_3222,N_3369);
nor U4634 (N_4634,N_3100,N_3248);
nand U4635 (N_4635,N_3432,N_3922);
nand U4636 (N_4636,N_3907,N_3925);
xnor U4637 (N_4637,N_3105,N_3084);
xor U4638 (N_4638,N_3173,N_3054);
and U4639 (N_4639,N_3532,N_3326);
xnor U4640 (N_4640,N_3330,N_3486);
nor U4641 (N_4641,N_3882,N_3969);
or U4642 (N_4642,N_3276,N_3855);
xnor U4643 (N_4643,N_3172,N_3154);
and U4644 (N_4644,N_3526,N_3918);
nor U4645 (N_4645,N_3145,N_3053);
and U4646 (N_4646,N_3941,N_3457);
and U4647 (N_4647,N_3284,N_3991);
nor U4648 (N_4648,N_3409,N_3121);
nor U4649 (N_4649,N_3516,N_3662);
or U4650 (N_4650,N_3104,N_3664);
nor U4651 (N_4651,N_3069,N_3336);
nor U4652 (N_4652,N_3245,N_3335);
and U4653 (N_4653,N_3284,N_3207);
nor U4654 (N_4654,N_3876,N_3855);
or U4655 (N_4655,N_3550,N_3284);
xnor U4656 (N_4656,N_3448,N_3046);
nor U4657 (N_4657,N_3299,N_3796);
or U4658 (N_4658,N_3300,N_3776);
and U4659 (N_4659,N_3312,N_3068);
and U4660 (N_4660,N_3522,N_3249);
nand U4661 (N_4661,N_3381,N_3402);
nor U4662 (N_4662,N_3161,N_3333);
and U4663 (N_4663,N_3163,N_3805);
xnor U4664 (N_4664,N_3583,N_3700);
nand U4665 (N_4665,N_3732,N_3908);
and U4666 (N_4666,N_3823,N_3591);
nor U4667 (N_4667,N_3060,N_3315);
or U4668 (N_4668,N_3090,N_3066);
nand U4669 (N_4669,N_3849,N_3012);
nand U4670 (N_4670,N_3436,N_3480);
and U4671 (N_4671,N_3431,N_3528);
or U4672 (N_4672,N_3081,N_3949);
or U4673 (N_4673,N_3726,N_3343);
xnor U4674 (N_4674,N_3782,N_3256);
nand U4675 (N_4675,N_3343,N_3604);
or U4676 (N_4676,N_3434,N_3195);
or U4677 (N_4677,N_3934,N_3062);
nor U4678 (N_4678,N_3762,N_3284);
nor U4679 (N_4679,N_3610,N_3793);
or U4680 (N_4680,N_3251,N_3915);
and U4681 (N_4681,N_3658,N_3435);
nand U4682 (N_4682,N_3804,N_3660);
and U4683 (N_4683,N_3737,N_3522);
and U4684 (N_4684,N_3672,N_3034);
nor U4685 (N_4685,N_3676,N_3130);
and U4686 (N_4686,N_3893,N_3774);
nor U4687 (N_4687,N_3694,N_3689);
nand U4688 (N_4688,N_3691,N_3607);
nor U4689 (N_4689,N_3246,N_3348);
or U4690 (N_4690,N_3207,N_3281);
nand U4691 (N_4691,N_3202,N_3836);
nor U4692 (N_4692,N_3676,N_3410);
and U4693 (N_4693,N_3122,N_3181);
nand U4694 (N_4694,N_3740,N_3713);
xnor U4695 (N_4695,N_3538,N_3607);
xor U4696 (N_4696,N_3820,N_3655);
nor U4697 (N_4697,N_3787,N_3983);
xnor U4698 (N_4698,N_3281,N_3886);
and U4699 (N_4699,N_3923,N_3501);
nand U4700 (N_4700,N_3429,N_3332);
xnor U4701 (N_4701,N_3758,N_3332);
xnor U4702 (N_4702,N_3598,N_3478);
or U4703 (N_4703,N_3967,N_3994);
and U4704 (N_4704,N_3279,N_3658);
nand U4705 (N_4705,N_3589,N_3328);
nor U4706 (N_4706,N_3216,N_3931);
or U4707 (N_4707,N_3939,N_3051);
and U4708 (N_4708,N_3732,N_3750);
nor U4709 (N_4709,N_3264,N_3856);
and U4710 (N_4710,N_3204,N_3933);
and U4711 (N_4711,N_3049,N_3194);
nand U4712 (N_4712,N_3074,N_3497);
xor U4713 (N_4713,N_3594,N_3697);
nand U4714 (N_4714,N_3773,N_3097);
and U4715 (N_4715,N_3291,N_3850);
nor U4716 (N_4716,N_3931,N_3935);
nor U4717 (N_4717,N_3697,N_3072);
nor U4718 (N_4718,N_3021,N_3231);
nand U4719 (N_4719,N_3363,N_3215);
or U4720 (N_4720,N_3743,N_3336);
or U4721 (N_4721,N_3100,N_3899);
nor U4722 (N_4722,N_3938,N_3088);
nor U4723 (N_4723,N_3992,N_3705);
nand U4724 (N_4724,N_3297,N_3083);
xor U4725 (N_4725,N_3947,N_3994);
and U4726 (N_4726,N_3722,N_3958);
or U4727 (N_4727,N_3171,N_3129);
and U4728 (N_4728,N_3030,N_3476);
nand U4729 (N_4729,N_3925,N_3093);
nand U4730 (N_4730,N_3982,N_3779);
xnor U4731 (N_4731,N_3575,N_3700);
xnor U4732 (N_4732,N_3195,N_3176);
nand U4733 (N_4733,N_3369,N_3571);
and U4734 (N_4734,N_3146,N_3115);
xnor U4735 (N_4735,N_3503,N_3539);
nor U4736 (N_4736,N_3959,N_3724);
or U4737 (N_4737,N_3216,N_3099);
or U4738 (N_4738,N_3748,N_3460);
and U4739 (N_4739,N_3280,N_3465);
and U4740 (N_4740,N_3020,N_3959);
nand U4741 (N_4741,N_3131,N_3913);
nand U4742 (N_4742,N_3633,N_3069);
nor U4743 (N_4743,N_3122,N_3311);
or U4744 (N_4744,N_3280,N_3590);
nand U4745 (N_4745,N_3548,N_3576);
or U4746 (N_4746,N_3767,N_3466);
or U4747 (N_4747,N_3725,N_3943);
or U4748 (N_4748,N_3882,N_3646);
nor U4749 (N_4749,N_3382,N_3389);
or U4750 (N_4750,N_3226,N_3350);
nand U4751 (N_4751,N_3839,N_3592);
or U4752 (N_4752,N_3820,N_3498);
nor U4753 (N_4753,N_3179,N_3449);
nand U4754 (N_4754,N_3887,N_3116);
or U4755 (N_4755,N_3618,N_3697);
nand U4756 (N_4756,N_3450,N_3016);
nor U4757 (N_4757,N_3594,N_3312);
and U4758 (N_4758,N_3783,N_3232);
nor U4759 (N_4759,N_3519,N_3963);
or U4760 (N_4760,N_3886,N_3216);
nor U4761 (N_4761,N_3121,N_3511);
xor U4762 (N_4762,N_3078,N_3957);
or U4763 (N_4763,N_3618,N_3929);
xnor U4764 (N_4764,N_3206,N_3149);
nand U4765 (N_4765,N_3353,N_3718);
or U4766 (N_4766,N_3314,N_3277);
xor U4767 (N_4767,N_3460,N_3527);
and U4768 (N_4768,N_3331,N_3531);
nand U4769 (N_4769,N_3655,N_3895);
and U4770 (N_4770,N_3540,N_3640);
nand U4771 (N_4771,N_3815,N_3873);
or U4772 (N_4772,N_3815,N_3443);
nand U4773 (N_4773,N_3164,N_3817);
and U4774 (N_4774,N_3237,N_3803);
or U4775 (N_4775,N_3304,N_3401);
or U4776 (N_4776,N_3042,N_3298);
and U4777 (N_4777,N_3053,N_3142);
xnor U4778 (N_4778,N_3171,N_3941);
nand U4779 (N_4779,N_3178,N_3299);
or U4780 (N_4780,N_3403,N_3125);
nand U4781 (N_4781,N_3441,N_3600);
xnor U4782 (N_4782,N_3516,N_3266);
xor U4783 (N_4783,N_3790,N_3688);
nor U4784 (N_4784,N_3512,N_3629);
or U4785 (N_4785,N_3911,N_3092);
nor U4786 (N_4786,N_3993,N_3898);
nor U4787 (N_4787,N_3320,N_3753);
or U4788 (N_4788,N_3667,N_3958);
or U4789 (N_4789,N_3118,N_3889);
and U4790 (N_4790,N_3332,N_3061);
nor U4791 (N_4791,N_3460,N_3113);
nor U4792 (N_4792,N_3719,N_3596);
or U4793 (N_4793,N_3626,N_3576);
and U4794 (N_4794,N_3636,N_3338);
nor U4795 (N_4795,N_3062,N_3734);
or U4796 (N_4796,N_3724,N_3825);
and U4797 (N_4797,N_3057,N_3534);
or U4798 (N_4798,N_3208,N_3761);
nand U4799 (N_4799,N_3109,N_3431);
nor U4800 (N_4800,N_3634,N_3153);
and U4801 (N_4801,N_3715,N_3203);
xor U4802 (N_4802,N_3460,N_3819);
and U4803 (N_4803,N_3096,N_3006);
or U4804 (N_4804,N_3709,N_3877);
nor U4805 (N_4805,N_3651,N_3871);
or U4806 (N_4806,N_3181,N_3165);
xor U4807 (N_4807,N_3622,N_3738);
xnor U4808 (N_4808,N_3200,N_3006);
and U4809 (N_4809,N_3024,N_3242);
xnor U4810 (N_4810,N_3804,N_3406);
nand U4811 (N_4811,N_3669,N_3895);
or U4812 (N_4812,N_3691,N_3137);
nor U4813 (N_4813,N_3101,N_3422);
or U4814 (N_4814,N_3537,N_3673);
nor U4815 (N_4815,N_3183,N_3738);
xor U4816 (N_4816,N_3462,N_3322);
nor U4817 (N_4817,N_3785,N_3923);
nor U4818 (N_4818,N_3607,N_3369);
nor U4819 (N_4819,N_3766,N_3735);
xor U4820 (N_4820,N_3985,N_3606);
nor U4821 (N_4821,N_3698,N_3605);
and U4822 (N_4822,N_3437,N_3145);
or U4823 (N_4823,N_3322,N_3723);
or U4824 (N_4824,N_3231,N_3581);
nand U4825 (N_4825,N_3370,N_3623);
nand U4826 (N_4826,N_3238,N_3754);
xor U4827 (N_4827,N_3852,N_3610);
and U4828 (N_4828,N_3569,N_3751);
nor U4829 (N_4829,N_3810,N_3697);
and U4830 (N_4830,N_3289,N_3942);
nand U4831 (N_4831,N_3558,N_3130);
and U4832 (N_4832,N_3773,N_3636);
nand U4833 (N_4833,N_3784,N_3293);
nand U4834 (N_4834,N_3132,N_3224);
nor U4835 (N_4835,N_3731,N_3326);
and U4836 (N_4836,N_3498,N_3456);
nor U4837 (N_4837,N_3922,N_3081);
or U4838 (N_4838,N_3765,N_3745);
and U4839 (N_4839,N_3970,N_3456);
nor U4840 (N_4840,N_3777,N_3686);
or U4841 (N_4841,N_3394,N_3249);
or U4842 (N_4842,N_3472,N_3659);
xor U4843 (N_4843,N_3666,N_3016);
xor U4844 (N_4844,N_3650,N_3617);
xor U4845 (N_4845,N_3943,N_3554);
xnor U4846 (N_4846,N_3891,N_3992);
and U4847 (N_4847,N_3688,N_3737);
and U4848 (N_4848,N_3365,N_3780);
nand U4849 (N_4849,N_3618,N_3934);
nor U4850 (N_4850,N_3643,N_3543);
xnor U4851 (N_4851,N_3909,N_3780);
xnor U4852 (N_4852,N_3908,N_3449);
nor U4853 (N_4853,N_3492,N_3159);
nor U4854 (N_4854,N_3232,N_3566);
or U4855 (N_4855,N_3305,N_3899);
nand U4856 (N_4856,N_3638,N_3741);
and U4857 (N_4857,N_3123,N_3393);
xor U4858 (N_4858,N_3040,N_3542);
or U4859 (N_4859,N_3344,N_3108);
and U4860 (N_4860,N_3179,N_3273);
nand U4861 (N_4861,N_3180,N_3697);
nor U4862 (N_4862,N_3626,N_3128);
nor U4863 (N_4863,N_3617,N_3313);
nor U4864 (N_4864,N_3061,N_3240);
or U4865 (N_4865,N_3311,N_3212);
xnor U4866 (N_4866,N_3473,N_3284);
xnor U4867 (N_4867,N_3920,N_3207);
nor U4868 (N_4868,N_3659,N_3490);
or U4869 (N_4869,N_3133,N_3769);
or U4870 (N_4870,N_3884,N_3741);
and U4871 (N_4871,N_3627,N_3573);
or U4872 (N_4872,N_3332,N_3246);
xnor U4873 (N_4873,N_3376,N_3503);
and U4874 (N_4874,N_3461,N_3817);
nor U4875 (N_4875,N_3638,N_3050);
or U4876 (N_4876,N_3928,N_3469);
or U4877 (N_4877,N_3339,N_3194);
nand U4878 (N_4878,N_3043,N_3565);
nand U4879 (N_4879,N_3057,N_3483);
nor U4880 (N_4880,N_3827,N_3577);
nor U4881 (N_4881,N_3392,N_3112);
nand U4882 (N_4882,N_3922,N_3181);
nor U4883 (N_4883,N_3881,N_3699);
nand U4884 (N_4884,N_3654,N_3146);
or U4885 (N_4885,N_3730,N_3194);
xnor U4886 (N_4886,N_3380,N_3115);
xor U4887 (N_4887,N_3031,N_3073);
and U4888 (N_4888,N_3311,N_3741);
and U4889 (N_4889,N_3624,N_3753);
and U4890 (N_4890,N_3524,N_3745);
nor U4891 (N_4891,N_3108,N_3002);
nor U4892 (N_4892,N_3723,N_3297);
and U4893 (N_4893,N_3727,N_3281);
or U4894 (N_4894,N_3664,N_3871);
or U4895 (N_4895,N_3325,N_3242);
or U4896 (N_4896,N_3513,N_3392);
nand U4897 (N_4897,N_3312,N_3210);
and U4898 (N_4898,N_3432,N_3169);
nor U4899 (N_4899,N_3355,N_3399);
nand U4900 (N_4900,N_3400,N_3030);
and U4901 (N_4901,N_3350,N_3316);
and U4902 (N_4902,N_3854,N_3993);
and U4903 (N_4903,N_3110,N_3893);
xor U4904 (N_4904,N_3740,N_3562);
nor U4905 (N_4905,N_3432,N_3775);
nand U4906 (N_4906,N_3495,N_3801);
and U4907 (N_4907,N_3109,N_3985);
nand U4908 (N_4908,N_3924,N_3567);
and U4909 (N_4909,N_3926,N_3045);
and U4910 (N_4910,N_3366,N_3753);
or U4911 (N_4911,N_3848,N_3933);
or U4912 (N_4912,N_3724,N_3614);
xnor U4913 (N_4913,N_3150,N_3561);
nor U4914 (N_4914,N_3439,N_3507);
xor U4915 (N_4915,N_3248,N_3304);
xnor U4916 (N_4916,N_3906,N_3267);
or U4917 (N_4917,N_3447,N_3385);
nor U4918 (N_4918,N_3644,N_3083);
or U4919 (N_4919,N_3062,N_3698);
and U4920 (N_4920,N_3623,N_3070);
xnor U4921 (N_4921,N_3109,N_3631);
nand U4922 (N_4922,N_3447,N_3635);
nand U4923 (N_4923,N_3201,N_3278);
or U4924 (N_4924,N_3716,N_3134);
xor U4925 (N_4925,N_3502,N_3372);
and U4926 (N_4926,N_3281,N_3714);
nor U4927 (N_4927,N_3983,N_3723);
nand U4928 (N_4928,N_3663,N_3136);
and U4929 (N_4929,N_3148,N_3336);
and U4930 (N_4930,N_3743,N_3944);
nor U4931 (N_4931,N_3203,N_3919);
and U4932 (N_4932,N_3127,N_3779);
xor U4933 (N_4933,N_3557,N_3754);
nor U4934 (N_4934,N_3500,N_3977);
or U4935 (N_4935,N_3528,N_3134);
or U4936 (N_4936,N_3865,N_3225);
or U4937 (N_4937,N_3386,N_3996);
nand U4938 (N_4938,N_3061,N_3150);
nor U4939 (N_4939,N_3166,N_3897);
and U4940 (N_4940,N_3555,N_3094);
or U4941 (N_4941,N_3205,N_3048);
or U4942 (N_4942,N_3990,N_3983);
nand U4943 (N_4943,N_3675,N_3955);
nor U4944 (N_4944,N_3033,N_3508);
xnor U4945 (N_4945,N_3155,N_3815);
and U4946 (N_4946,N_3131,N_3989);
and U4947 (N_4947,N_3256,N_3294);
or U4948 (N_4948,N_3757,N_3763);
or U4949 (N_4949,N_3310,N_3560);
nor U4950 (N_4950,N_3102,N_3702);
or U4951 (N_4951,N_3420,N_3744);
nor U4952 (N_4952,N_3024,N_3061);
xnor U4953 (N_4953,N_3198,N_3856);
nand U4954 (N_4954,N_3873,N_3543);
nor U4955 (N_4955,N_3431,N_3593);
nand U4956 (N_4956,N_3912,N_3083);
xnor U4957 (N_4957,N_3170,N_3235);
or U4958 (N_4958,N_3980,N_3742);
nor U4959 (N_4959,N_3788,N_3750);
xnor U4960 (N_4960,N_3400,N_3446);
or U4961 (N_4961,N_3954,N_3725);
nor U4962 (N_4962,N_3874,N_3403);
nand U4963 (N_4963,N_3700,N_3102);
nor U4964 (N_4964,N_3241,N_3365);
nand U4965 (N_4965,N_3156,N_3476);
nand U4966 (N_4966,N_3873,N_3798);
or U4967 (N_4967,N_3396,N_3842);
and U4968 (N_4968,N_3774,N_3306);
and U4969 (N_4969,N_3369,N_3289);
or U4970 (N_4970,N_3161,N_3738);
nand U4971 (N_4971,N_3329,N_3482);
or U4972 (N_4972,N_3841,N_3779);
xor U4973 (N_4973,N_3007,N_3228);
nor U4974 (N_4974,N_3902,N_3936);
nand U4975 (N_4975,N_3616,N_3308);
xor U4976 (N_4976,N_3495,N_3664);
nand U4977 (N_4977,N_3767,N_3299);
nand U4978 (N_4978,N_3268,N_3744);
nor U4979 (N_4979,N_3432,N_3429);
nor U4980 (N_4980,N_3844,N_3886);
nor U4981 (N_4981,N_3226,N_3081);
nor U4982 (N_4982,N_3651,N_3992);
and U4983 (N_4983,N_3950,N_3051);
and U4984 (N_4984,N_3998,N_3358);
xnor U4985 (N_4985,N_3275,N_3649);
or U4986 (N_4986,N_3803,N_3337);
xnor U4987 (N_4987,N_3418,N_3684);
and U4988 (N_4988,N_3229,N_3626);
nor U4989 (N_4989,N_3625,N_3671);
and U4990 (N_4990,N_3611,N_3197);
and U4991 (N_4991,N_3901,N_3707);
nor U4992 (N_4992,N_3848,N_3475);
nor U4993 (N_4993,N_3963,N_3865);
xor U4994 (N_4994,N_3782,N_3996);
nor U4995 (N_4995,N_3549,N_3703);
nor U4996 (N_4996,N_3439,N_3045);
or U4997 (N_4997,N_3673,N_3103);
xnor U4998 (N_4998,N_3401,N_3176);
nor U4999 (N_4999,N_3151,N_3946);
or U5000 (N_5000,N_4994,N_4435);
and U5001 (N_5001,N_4491,N_4863);
nor U5002 (N_5002,N_4497,N_4219);
xor U5003 (N_5003,N_4932,N_4006);
or U5004 (N_5004,N_4022,N_4878);
nand U5005 (N_5005,N_4028,N_4152);
xnor U5006 (N_5006,N_4218,N_4430);
nand U5007 (N_5007,N_4766,N_4475);
and U5008 (N_5008,N_4266,N_4903);
and U5009 (N_5009,N_4482,N_4990);
or U5010 (N_5010,N_4551,N_4904);
or U5011 (N_5011,N_4993,N_4421);
and U5012 (N_5012,N_4592,N_4817);
and U5013 (N_5013,N_4397,N_4331);
nor U5014 (N_5014,N_4630,N_4829);
or U5015 (N_5015,N_4850,N_4853);
nand U5016 (N_5016,N_4691,N_4857);
nand U5017 (N_5017,N_4207,N_4263);
xnor U5018 (N_5018,N_4976,N_4543);
xor U5019 (N_5019,N_4610,N_4957);
or U5020 (N_5020,N_4872,N_4443);
xnor U5021 (N_5021,N_4777,N_4288);
nor U5022 (N_5022,N_4518,N_4341);
nor U5023 (N_5023,N_4647,N_4333);
nand U5024 (N_5024,N_4859,N_4371);
xnor U5025 (N_5025,N_4786,N_4665);
xor U5026 (N_5026,N_4529,N_4827);
nand U5027 (N_5027,N_4548,N_4368);
and U5028 (N_5028,N_4703,N_4009);
and U5029 (N_5029,N_4605,N_4729);
xnor U5030 (N_5030,N_4923,N_4113);
nand U5031 (N_5031,N_4235,N_4176);
nor U5032 (N_5032,N_4492,N_4226);
nor U5033 (N_5033,N_4267,N_4713);
nor U5034 (N_5034,N_4940,N_4626);
xor U5035 (N_5035,N_4110,N_4483);
or U5036 (N_5036,N_4897,N_4679);
or U5037 (N_5037,N_4458,N_4404);
and U5038 (N_5038,N_4956,N_4547);
xor U5039 (N_5039,N_4600,N_4025);
or U5040 (N_5040,N_4507,N_4415);
and U5041 (N_5041,N_4583,N_4667);
nand U5042 (N_5042,N_4374,N_4012);
or U5043 (N_5043,N_4389,N_4325);
xnor U5044 (N_5044,N_4047,N_4385);
nand U5045 (N_5045,N_4178,N_4841);
or U5046 (N_5046,N_4702,N_4517);
xor U5047 (N_5047,N_4171,N_4106);
and U5048 (N_5048,N_4314,N_4925);
nand U5049 (N_5049,N_4063,N_4305);
and U5050 (N_5050,N_4036,N_4464);
xor U5051 (N_5051,N_4370,N_4005);
nand U5052 (N_5052,N_4060,N_4865);
or U5053 (N_5053,N_4274,N_4780);
nand U5054 (N_5054,N_4715,N_4920);
and U5055 (N_5055,N_4864,N_4882);
xnor U5056 (N_5056,N_4455,N_4130);
and U5057 (N_5057,N_4177,N_4574);
nand U5058 (N_5058,N_4030,N_4582);
and U5059 (N_5059,N_4253,N_4092);
and U5060 (N_5060,N_4871,N_4500);
and U5061 (N_5061,N_4624,N_4898);
and U5062 (N_5062,N_4425,N_4011);
nor U5063 (N_5063,N_4390,N_4714);
nand U5064 (N_5064,N_4296,N_4162);
nand U5065 (N_5065,N_4919,N_4079);
or U5066 (N_5066,N_4540,N_4654);
or U5067 (N_5067,N_4800,N_4391);
or U5068 (N_5068,N_4159,N_4280);
or U5069 (N_5069,N_4446,N_4598);
or U5070 (N_5070,N_4489,N_4151);
and U5071 (N_5071,N_4292,N_4620);
or U5072 (N_5072,N_4604,N_4033);
xnor U5073 (N_5073,N_4143,N_4965);
nor U5074 (N_5074,N_4375,N_4740);
or U5075 (N_5075,N_4186,N_4129);
xnor U5076 (N_5076,N_4462,N_4877);
xor U5077 (N_5077,N_4788,N_4660);
and U5078 (N_5078,N_4613,N_4680);
xnor U5079 (N_5079,N_4319,N_4429);
and U5080 (N_5080,N_4245,N_4222);
xor U5081 (N_5081,N_4479,N_4422);
nor U5082 (N_5082,N_4811,N_4456);
nor U5083 (N_5083,N_4577,N_4173);
nor U5084 (N_5084,N_4289,N_4705);
nand U5085 (N_5085,N_4791,N_4732);
or U5086 (N_5086,N_4142,N_4234);
and U5087 (N_5087,N_4444,N_4073);
or U5088 (N_5088,N_4531,N_4460);
and U5089 (N_5089,N_4363,N_4868);
or U5090 (N_5090,N_4513,N_4861);
xor U5091 (N_5091,N_4706,N_4646);
nor U5092 (N_5092,N_4787,N_4830);
nand U5093 (N_5093,N_4587,N_4942);
or U5094 (N_5094,N_4306,N_4217);
nand U5095 (N_5095,N_4287,N_4744);
and U5096 (N_5096,N_4156,N_4040);
and U5097 (N_5097,N_4140,N_4221);
nand U5098 (N_5098,N_4818,N_4992);
and U5099 (N_5099,N_4031,N_4843);
xnor U5100 (N_5100,N_4104,N_4242);
nand U5101 (N_5101,N_4378,N_4670);
and U5102 (N_5102,N_4058,N_4137);
nand U5103 (N_5103,N_4498,N_4769);
nand U5104 (N_5104,N_4180,N_4983);
or U5105 (N_5105,N_4188,N_4803);
nor U5106 (N_5106,N_4000,N_4027);
and U5107 (N_5107,N_4912,N_4407);
or U5108 (N_5108,N_4096,N_4192);
and U5109 (N_5109,N_4884,N_4959);
xnor U5110 (N_5110,N_4399,N_4820);
or U5111 (N_5111,N_4915,N_4150);
nor U5112 (N_5112,N_4534,N_4449);
nor U5113 (N_5113,N_4053,N_4308);
nand U5114 (N_5114,N_4121,N_4324);
or U5115 (N_5115,N_4332,N_4614);
and U5116 (N_5116,N_4494,N_4189);
or U5117 (N_5117,N_4916,N_4974);
and U5118 (N_5118,N_4725,N_4765);
and U5119 (N_5119,N_4286,N_4808);
nand U5120 (N_5120,N_4282,N_4776);
nor U5121 (N_5121,N_4416,N_4612);
nor U5122 (N_5122,N_4511,N_4487);
or U5123 (N_5123,N_4730,N_4366);
nor U5124 (N_5124,N_4671,N_4380);
nand U5125 (N_5125,N_4495,N_4484);
nor U5126 (N_5126,N_4069,N_4508);
nor U5127 (N_5127,N_4578,N_4989);
or U5128 (N_5128,N_4571,N_4295);
xor U5129 (N_5129,N_4533,N_4938);
xnor U5130 (N_5130,N_4210,N_4886);
nor U5131 (N_5131,N_4465,N_4386);
and U5132 (N_5132,N_4828,N_4698);
and U5133 (N_5133,N_4812,N_4418);
or U5134 (N_5134,N_4962,N_4690);
nand U5135 (N_5135,N_4401,N_4239);
nor U5136 (N_5136,N_4781,N_4269);
nor U5137 (N_5137,N_4199,N_4569);
or U5138 (N_5138,N_4590,N_4634);
nand U5139 (N_5139,N_4819,N_4082);
nor U5140 (N_5140,N_4064,N_4168);
nand U5141 (N_5141,N_4656,N_4419);
nand U5142 (N_5142,N_4695,N_4034);
or U5143 (N_5143,N_4050,N_4591);
or U5144 (N_5144,N_4666,N_4521);
nor U5145 (N_5145,N_4773,N_4493);
nor U5146 (N_5146,N_4616,N_4166);
nor U5147 (N_5147,N_4147,N_4985);
and U5148 (N_5148,N_4258,N_4016);
xnor U5149 (N_5149,N_4561,N_4453);
nor U5150 (N_5150,N_4738,N_4799);
and U5151 (N_5151,N_4327,N_4621);
or U5152 (N_5152,N_4760,N_4541);
nand U5153 (N_5153,N_4070,N_4170);
xor U5154 (N_5154,N_4095,N_4035);
or U5155 (N_5155,N_4608,N_4109);
nand U5156 (N_5156,N_4987,N_4899);
or U5157 (N_5157,N_4681,N_4554);
nor U5158 (N_5158,N_4148,N_4595);
nor U5159 (N_5159,N_4984,N_4383);
and U5160 (N_5160,N_4094,N_4270);
or U5161 (N_5161,N_4439,N_4568);
and U5162 (N_5162,N_4699,N_4051);
or U5163 (N_5163,N_4074,N_4284);
or U5164 (N_5164,N_4914,N_4833);
xor U5165 (N_5165,N_4798,N_4944);
or U5166 (N_5166,N_4523,N_4960);
nor U5167 (N_5167,N_4516,N_4043);
or U5168 (N_5168,N_4657,N_4570);
nand U5169 (N_5169,N_4860,N_4741);
nor U5170 (N_5170,N_4157,N_4467);
xor U5171 (N_5171,N_4562,N_4349);
and U5172 (N_5172,N_4640,N_4215);
xor U5173 (N_5173,N_4139,N_4054);
xnor U5174 (N_5174,N_4623,N_4015);
xor U5175 (N_5175,N_4975,N_4122);
nor U5176 (N_5176,N_4254,N_4686);
nor U5177 (N_5177,N_4238,N_4806);
nand U5178 (N_5178,N_4565,N_4514);
and U5179 (N_5179,N_4486,N_4816);
and U5180 (N_5180,N_4795,N_4801);
nand U5181 (N_5181,N_4427,N_4936);
nand U5182 (N_5182,N_4711,N_4745);
nor U5183 (N_5183,N_4361,N_4021);
xnor U5184 (N_5184,N_4826,N_4892);
nor U5185 (N_5185,N_4126,N_4302);
or U5186 (N_5186,N_4986,N_4161);
nand U5187 (N_5187,N_4653,N_4585);
nand U5188 (N_5188,N_4727,N_4472);
nor U5189 (N_5189,N_4154,N_4204);
and U5190 (N_5190,N_4717,N_4155);
nor U5191 (N_5191,N_4880,N_4510);
and U5192 (N_5192,N_4278,N_4693);
or U5193 (N_5193,N_4503,N_4169);
and U5194 (N_5194,N_4952,N_4979);
or U5195 (N_5195,N_4961,N_4538);
and U5196 (N_5196,N_4488,N_4356);
nor U5197 (N_5197,N_4659,N_4902);
and U5198 (N_5198,N_4193,N_4596);
or U5199 (N_5199,N_4573,N_4719);
xor U5200 (N_5200,N_4707,N_4271);
nand U5201 (N_5201,N_4118,N_4526);
or U5202 (N_5202,N_4567,N_4650);
or U5203 (N_5203,N_4953,N_4645);
nor U5204 (N_5204,N_4572,N_4772);
and U5205 (N_5205,N_4447,N_4704);
nand U5206 (N_5206,N_4255,N_4236);
and U5207 (N_5207,N_4739,N_4782);
or U5208 (N_5208,N_4874,N_4347);
nand U5209 (N_5209,N_4996,N_4307);
or U5210 (N_5210,N_4683,N_4196);
nand U5211 (N_5211,N_4553,N_4606);
nand U5212 (N_5212,N_4933,N_4243);
or U5213 (N_5213,N_4875,N_4209);
xnor U5214 (N_5214,N_4097,N_4206);
nor U5215 (N_5215,N_4297,N_4889);
or U5216 (N_5216,N_4358,N_4756);
nand U5217 (N_5217,N_4794,N_4726);
nand U5218 (N_5218,N_4580,N_4869);
or U5219 (N_5219,N_4758,N_4083);
or U5220 (N_5220,N_4136,N_4790);
nor U5221 (N_5221,N_4928,N_4682);
xor U5222 (N_5222,N_4748,N_4937);
xor U5223 (N_5223,N_4125,N_4339);
xor U5224 (N_5224,N_4203,N_4259);
xnor U5225 (N_5225,N_4550,N_4963);
and U5226 (N_5226,N_4087,N_4335);
or U5227 (N_5227,N_4958,N_4838);
nor U5228 (N_5228,N_4576,N_4895);
or U5229 (N_5229,N_4098,N_4537);
nand U5230 (N_5230,N_4896,N_4918);
nor U5231 (N_5231,N_4056,N_4135);
and U5232 (N_5232,N_4246,N_4870);
nor U5233 (N_5233,N_4948,N_4014);
or U5234 (N_5234,N_4228,N_4466);
xor U5235 (N_5235,N_4348,N_4910);
nand U5236 (N_5236,N_4619,N_4075);
and U5237 (N_5237,N_4424,N_4888);
nor U5238 (N_5238,N_4190,N_4736);
xor U5239 (N_5239,N_4310,N_4622);
or U5240 (N_5240,N_4793,N_4778);
or U5241 (N_5241,N_4119,N_4103);
and U5242 (N_5242,N_4013,N_4972);
nand U5243 (N_5243,N_4607,N_4856);
or U5244 (N_5244,N_4149,N_4586);
nor U5245 (N_5245,N_4542,N_4107);
and U5246 (N_5246,N_4771,N_4644);
or U5247 (N_5247,N_4977,N_4412);
nand U5248 (N_5248,N_4476,N_4629);
nand U5249 (N_5249,N_4692,N_4779);
nand U5250 (N_5250,N_4805,N_4968);
nor U5251 (N_5251,N_4409,N_4611);
and U5252 (N_5252,N_4244,N_4661);
or U5253 (N_5253,N_4250,N_4597);
or U5254 (N_5254,N_4480,N_4164);
nand U5255 (N_5255,N_4746,N_4291);
xor U5256 (N_5256,N_4594,N_4367);
nor U5257 (N_5257,N_4685,N_4544);
and U5258 (N_5258,N_4473,N_4023);
nor U5259 (N_5259,N_4546,N_4195);
nand U5260 (N_5260,N_4459,N_4539);
or U5261 (N_5261,N_4909,N_4396);
xnor U5262 (N_5262,N_4501,N_4873);
xnor U5263 (N_5263,N_4340,N_4810);
nor U5264 (N_5264,N_4978,N_4728);
nor U5265 (N_5265,N_4436,N_4825);
nor U5266 (N_5266,N_4426,N_4858);
or U5267 (N_5267,N_4499,N_4277);
or U5268 (N_5268,N_4609,N_4628);
nor U5269 (N_5269,N_4062,N_4232);
and U5270 (N_5270,N_4837,N_4675);
nor U5271 (N_5271,N_4835,N_4262);
nand U5272 (N_5272,N_4617,N_4381);
xnor U5273 (N_5273,N_4839,N_4247);
xnor U5274 (N_5274,N_4527,N_4988);
nand U5275 (N_5275,N_4018,N_4579);
or U5276 (N_5276,N_4849,N_4764);
nand U5277 (N_5277,N_4792,N_4301);
nor U5278 (N_5278,N_4328,N_4470);
nor U5279 (N_5279,N_4824,N_4545);
or U5280 (N_5280,N_4322,N_4048);
or U5281 (N_5281,N_4144,N_4663);
nor U5282 (N_5282,N_4212,N_4007);
xor U5283 (N_5283,N_4934,N_4900);
nand U5284 (N_5284,N_4982,N_4532);
nor U5285 (N_5285,N_4002,N_4638);
or U5286 (N_5286,N_4844,N_4907);
or U5287 (N_5287,N_4338,N_4796);
xnor U5288 (N_5288,N_4851,N_4105);
xor U5289 (N_5289,N_4452,N_4395);
nor U5290 (N_5290,N_4632,N_4566);
xor U5291 (N_5291,N_4505,N_4197);
xnor U5292 (N_5292,N_4211,N_4133);
nand U5293 (N_5293,N_4478,N_4750);
xor U5294 (N_5294,N_4037,N_4949);
xor U5295 (N_5295,N_4905,N_4172);
nor U5296 (N_5296,N_4408,N_4346);
or U5297 (N_5297,N_4722,N_4530);
or U5298 (N_5298,N_4929,N_4615);
nor U5299 (N_5299,N_4879,N_4260);
xor U5300 (N_5300,N_4194,N_4834);
or U5301 (N_5301,N_4261,N_4981);
or U5302 (N_5302,N_4101,N_4442);
or U5303 (N_5303,N_4716,N_4102);
xor U5304 (N_5304,N_4032,N_4184);
nor U5305 (N_5305,N_4669,N_4405);
nand U5306 (N_5306,N_4004,N_4970);
nand U5307 (N_5307,N_4709,N_4969);
and U5308 (N_5308,N_4127,N_4496);
nor U5309 (N_5309,N_4635,N_4676);
nand U5310 (N_5310,N_4939,N_4373);
or U5311 (N_5311,N_4490,N_4814);
nand U5312 (N_5312,N_4557,N_4298);
or U5313 (N_5313,N_4894,N_4823);
xnor U5314 (N_5314,N_4890,N_4272);
and U5315 (N_5315,N_4017,N_4697);
or U5316 (N_5316,N_4563,N_4230);
nor U5317 (N_5317,N_4668,N_4461);
or U5318 (N_5318,N_4352,N_4710);
nor U5319 (N_5319,N_4290,N_4625);
and U5320 (N_5320,N_4931,N_4636);
or U5321 (N_5321,N_4081,N_4268);
xor U5322 (N_5322,N_4807,N_4767);
and U5323 (N_5323,N_4078,N_4524);
xor U5324 (N_5324,N_4181,N_4967);
nand U5325 (N_5325,N_4128,N_4564);
nor U5326 (N_5326,N_4330,N_4862);
nand U5327 (N_5327,N_4584,N_4627);
or U5328 (N_5328,N_4132,N_4995);
xnor U5329 (N_5329,N_4019,N_4317);
nor U5330 (N_5330,N_4088,N_4588);
xor U5331 (N_5331,N_4202,N_4108);
and U5332 (N_5332,N_4420,N_4735);
or U5333 (N_5333,N_4227,N_4065);
and U5334 (N_5334,N_4343,N_4163);
nand U5335 (N_5335,N_4672,N_4351);
xnor U5336 (N_5336,N_4283,N_4631);
nand U5337 (N_5337,N_4689,N_4575);
xnor U5338 (N_5338,N_4930,N_4237);
nor U5339 (N_5339,N_4721,N_4309);
xnor U5340 (N_5340,N_4633,N_4355);
nor U5341 (N_5341,N_4813,N_4337);
or U5342 (N_5342,N_4887,N_4294);
and U5343 (N_5343,N_4362,N_4755);
or U5344 (N_5344,N_4240,N_4311);
xnor U5345 (N_5345,N_4326,N_4205);
xor U5346 (N_5346,N_4376,N_4091);
and U5347 (N_5347,N_4469,N_4922);
nand U5348 (N_5348,N_4775,N_4747);
or U5349 (N_5349,N_4304,N_4077);
nor U5350 (N_5350,N_4751,N_4846);
or U5351 (N_5351,N_4350,N_4279);
nor U5352 (N_5352,N_4251,N_4413);
nor U5353 (N_5353,N_4481,N_4115);
nand U5354 (N_5354,N_4881,N_4124);
xor U5355 (N_5355,N_4997,N_4753);
and U5356 (N_5356,N_4379,N_4049);
or U5357 (N_5357,N_4067,N_4917);
xor U5358 (N_5358,N_4201,N_4457);
and U5359 (N_5359,N_4520,N_4648);
xnor U5360 (N_5360,N_4734,N_4141);
and U5361 (N_5361,N_4602,N_4336);
and U5362 (N_5362,N_4403,N_4752);
nand U5363 (N_5363,N_4411,N_4276);
and U5364 (N_5364,N_4001,N_4123);
nand U5365 (N_5365,N_4885,N_4662);
or U5366 (N_5366,N_4468,N_4559);
or U5367 (N_5367,N_4382,N_4131);
xnor U5368 (N_5368,N_4973,N_4655);
nor U5369 (N_5369,N_4208,N_4761);
nor U5370 (N_5370,N_4980,N_4175);
or U5371 (N_5371,N_4770,N_4463);
and U5372 (N_5372,N_4146,N_4353);
and U5373 (N_5373,N_4406,N_4099);
nor U5374 (N_5374,N_4804,N_4743);
nor U5375 (N_5375,N_4059,N_4893);
xor U5376 (N_5376,N_4512,N_4964);
nor U5377 (N_5377,N_4854,N_4313);
or U5378 (N_5378,N_4618,N_4883);
nand U5379 (N_5379,N_4999,N_4428);
nand U5380 (N_5380,N_4364,N_4111);
xor U5381 (N_5381,N_4599,N_4300);
nor U5382 (N_5382,N_4112,N_4345);
nor U5383 (N_5383,N_4182,N_4966);
nor U5384 (N_5384,N_4684,N_4536);
nand U5385 (N_5385,N_4248,N_4089);
nor U5386 (N_5386,N_4822,N_4593);
or U5387 (N_5387,N_4410,N_4998);
or U5388 (N_5388,N_4876,N_4072);
or U5389 (N_5389,N_4673,N_4233);
nand U5390 (N_5390,N_4637,N_4522);
xnor U5391 (N_5391,N_4431,N_4008);
or U5392 (N_5392,N_4924,N_4055);
or U5393 (N_5393,N_4066,N_4252);
nand U5394 (N_5394,N_4560,N_4045);
or U5395 (N_5395,N_4951,N_4312);
and U5396 (N_5396,N_4320,N_4400);
or U5397 (N_5397,N_4589,N_4555);
or U5398 (N_5398,N_4445,N_4774);
xnor U5399 (N_5399,N_4954,N_4941);
xor U5400 (N_5400,N_4901,N_4165);
or U5401 (N_5401,N_4502,N_4116);
nand U5402 (N_5402,N_4652,N_4388);
or U5403 (N_5403,N_4093,N_4789);
nor U5404 (N_5404,N_4076,N_4768);
xor U5405 (N_5405,N_4438,N_4947);
nand U5406 (N_5406,N_4815,N_4090);
nand U5407 (N_5407,N_4100,N_4010);
nand U5408 (N_5408,N_4504,N_4387);
and U5409 (N_5409,N_4448,N_4138);
and U5410 (N_5410,N_4264,N_4913);
nor U5411 (N_5411,N_4649,N_4708);
nand U5412 (N_5412,N_4414,N_4257);
xor U5413 (N_5413,N_4836,N_4318);
or U5414 (N_5414,N_4214,N_4519);
and U5415 (N_5415,N_4114,N_4249);
nand U5416 (N_5416,N_4733,N_4334);
nand U5417 (N_5417,N_4299,N_4677);
nand U5418 (N_5418,N_4394,N_4955);
xor U5419 (N_5419,N_4971,N_4134);
or U5420 (N_5420,N_4821,N_4831);
xor U5421 (N_5421,N_4052,N_4285);
nand U5422 (N_5422,N_4344,N_4256);
xnor U5423 (N_5423,N_4342,N_4057);
nand U5424 (N_5424,N_4041,N_4506);
nor U5425 (N_5425,N_4525,N_4200);
nor U5426 (N_5426,N_4754,N_4509);
and U5427 (N_5427,N_4762,N_4039);
nand U5428 (N_5428,N_4866,N_4674);
nor U5429 (N_5429,N_4042,N_4701);
xor U5430 (N_5430,N_4450,N_4664);
xor U5431 (N_5431,N_4360,N_4474);
xnor U5432 (N_5432,N_4029,N_4688);
nand U5433 (N_5433,N_4784,N_4485);
nor U5434 (N_5434,N_4145,N_4323);
and U5435 (N_5435,N_4086,N_4847);
nor U5436 (N_5436,N_4026,N_4024);
nor U5437 (N_5437,N_4158,N_4737);
or U5438 (N_5438,N_4581,N_4265);
xor U5439 (N_5439,N_4840,N_4549);
nor U5440 (N_5440,N_4432,N_4417);
and U5441 (N_5441,N_4643,N_4187);
nand U5442 (N_5442,N_4068,N_4639);
nor U5443 (N_5443,N_4908,N_4451);
and U5444 (N_5444,N_4696,N_4183);
and U5445 (N_5445,N_4398,N_4678);
or U5446 (N_5446,N_4950,N_4921);
and U5447 (N_5447,N_4225,N_4393);
nand U5448 (N_5448,N_4515,N_4354);
xor U5449 (N_5449,N_4003,N_4229);
nand U5450 (N_5450,N_4372,N_4384);
xnor U5451 (N_5451,N_4434,N_4528);
nand U5452 (N_5452,N_4071,N_4061);
nor U5453 (N_5453,N_4044,N_4437);
and U5454 (N_5454,N_4185,N_4757);
xor U5455 (N_5455,N_4315,N_4556);
nand U5456 (N_5456,N_4216,N_4117);
nor U5457 (N_5457,N_4759,N_4321);
xor U5458 (N_5458,N_4832,N_4433);
nand U5459 (N_5459,N_4160,N_4891);
nor U5460 (N_5460,N_4369,N_4783);
nand U5461 (N_5461,N_4046,N_4224);
and U5462 (N_5462,N_4153,N_4651);
nand U5463 (N_5463,N_4848,N_4694);
nor U5464 (N_5464,N_4991,N_4392);
and U5465 (N_5465,N_4293,N_4085);
and U5466 (N_5466,N_4911,N_4723);
nor U5467 (N_5467,N_4720,N_4471);
and U5468 (N_5468,N_4231,N_4809);
and U5469 (N_5469,N_4167,N_4601);
xnor U5470 (N_5470,N_4926,N_4852);
and U5471 (N_5471,N_4174,N_4552);
and U5472 (N_5472,N_4281,N_4658);
and U5473 (N_5473,N_4377,N_4213);
nand U5474 (N_5474,N_4275,N_4687);
xnor U5475 (N_5475,N_4441,N_4329);
and U5476 (N_5476,N_4724,N_4241);
nand U5477 (N_5477,N_4731,N_4935);
xnor U5478 (N_5478,N_4303,N_4946);
nor U5479 (N_5479,N_4641,N_4220);
and U5480 (N_5480,N_4423,N_4316);
or U5481 (N_5481,N_4454,N_4179);
or U5482 (N_5482,N_4797,N_4558);
or U5483 (N_5483,N_4223,N_4927);
and U5484 (N_5484,N_4120,N_4802);
xnor U5485 (N_5485,N_4742,N_4718);
xor U5486 (N_5486,N_4365,N_4080);
or U5487 (N_5487,N_4273,N_4359);
or U5488 (N_5488,N_4855,N_4477);
and U5489 (N_5489,N_4845,N_4842);
xnor U5490 (N_5490,N_4357,N_4785);
and U5491 (N_5491,N_4712,N_4603);
xnor U5492 (N_5492,N_4763,N_4945);
nor U5493 (N_5493,N_4906,N_4198);
nand U5494 (N_5494,N_4084,N_4700);
or U5495 (N_5495,N_4038,N_4642);
and U5496 (N_5496,N_4440,N_4191);
and U5497 (N_5497,N_4749,N_4943);
nor U5498 (N_5498,N_4535,N_4402);
and U5499 (N_5499,N_4020,N_4867);
and U5500 (N_5500,N_4552,N_4589);
nand U5501 (N_5501,N_4515,N_4954);
or U5502 (N_5502,N_4971,N_4255);
nor U5503 (N_5503,N_4782,N_4674);
nand U5504 (N_5504,N_4722,N_4038);
or U5505 (N_5505,N_4038,N_4980);
nand U5506 (N_5506,N_4062,N_4423);
and U5507 (N_5507,N_4177,N_4780);
nand U5508 (N_5508,N_4969,N_4976);
and U5509 (N_5509,N_4221,N_4718);
or U5510 (N_5510,N_4761,N_4319);
xnor U5511 (N_5511,N_4645,N_4529);
nand U5512 (N_5512,N_4010,N_4060);
or U5513 (N_5513,N_4594,N_4400);
xnor U5514 (N_5514,N_4469,N_4254);
nor U5515 (N_5515,N_4827,N_4957);
and U5516 (N_5516,N_4774,N_4489);
or U5517 (N_5517,N_4213,N_4800);
nor U5518 (N_5518,N_4654,N_4269);
or U5519 (N_5519,N_4161,N_4548);
or U5520 (N_5520,N_4387,N_4108);
xnor U5521 (N_5521,N_4557,N_4584);
or U5522 (N_5522,N_4068,N_4025);
nor U5523 (N_5523,N_4063,N_4537);
and U5524 (N_5524,N_4844,N_4738);
or U5525 (N_5525,N_4933,N_4936);
nor U5526 (N_5526,N_4831,N_4427);
or U5527 (N_5527,N_4541,N_4595);
xnor U5528 (N_5528,N_4387,N_4699);
and U5529 (N_5529,N_4174,N_4838);
or U5530 (N_5530,N_4441,N_4124);
nand U5531 (N_5531,N_4538,N_4966);
xnor U5532 (N_5532,N_4450,N_4931);
or U5533 (N_5533,N_4003,N_4846);
or U5534 (N_5534,N_4330,N_4591);
xor U5535 (N_5535,N_4982,N_4067);
nand U5536 (N_5536,N_4189,N_4995);
nor U5537 (N_5537,N_4533,N_4307);
nand U5538 (N_5538,N_4326,N_4802);
xnor U5539 (N_5539,N_4295,N_4818);
xnor U5540 (N_5540,N_4235,N_4693);
xor U5541 (N_5541,N_4938,N_4267);
nand U5542 (N_5542,N_4350,N_4755);
nand U5543 (N_5543,N_4756,N_4846);
nor U5544 (N_5544,N_4674,N_4427);
or U5545 (N_5545,N_4340,N_4789);
nand U5546 (N_5546,N_4490,N_4285);
nor U5547 (N_5547,N_4500,N_4483);
xor U5548 (N_5548,N_4288,N_4757);
xor U5549 (N_5549,N_4608,N_4691);
nor U5550 (N_5550,N_4773,N_4974);
xnor U5551 (N_5551,N_4971,N_4026);
and U5552 (N_5552,N_4200,N_4488);
nand U5553 (N_5553,N_4335,N_4014);
xnor U5554 (N_5554,N_4106,N_4466);
and U5555 (N_5555,N_4021,N_4807);
and U5556 (N_5556,N_4471,N_4537);
xor U5557 (N_5557,N_4369,N_4832);
xor U5558 (N_5558,N_4615,N_4981);
xnor U5559 (N_5559,N_4630,N_4889);
xor U5560 (N_5560,N_4190,N_4372);
nor U5561 (N_5561,N_4921,N_4250);
nand U5562 (N_5562,N_4237,N_4860);
or U5563 (N_5563,N_4734,N_4911);
xnor U5564 (N_5564,N_4471,N_4738);
or U5565 (N_5565,N_4340,N_4138);
nor U5566 (N_5566,N_4521,N_4287);
or U5567 (N_5567,N_4288,N_4560);
nand U5568 (N_5568,N_4932,N_4801);
xor U5569 (N_5569,N_4128,N_4884);
nand U5570 (N_5570,N_4993,N_4061);
or U5571 (N_5571,N_4160,N_4768);
nor U5572 (N_5572,N_4937,N_4248);
or U5573 (N_5573,N_4579,N_4668);
and U5574 (N_5574,N_4158,N_4236);
and U5575 (N_5575,N_4157,N_4937);
and U5576 (N_5576,N_4303,N_4707);
xor U5577 (N_5577,N_4028,N_4835);
nand U5578 (N_5578,N_4191,N_4115);
or U5579 (N_5579,N_4938,N_4465);
and U5580 (N_5580,N_4054,N_4899);
or U5581 (N_5581,N_4688,N_4654);
or U5582 (N_5582,N_4054,N_4071);
xor U5583 (N_5583,N_4856,N_4524);
or U5584 (N_5584,N_4977,N_4459);
nand U5585 (N_5585,N_4518,N_4435);
nand U5586 (N_5586,N_4511,N_4288);
xor U5587 (N_5587,N_4861,N_4079);
or U5588 (N_5588,N_4095,N_4064);
and U5589 (N_5589,N_4653,N_4416);
and U5590 (N_5590,N_4012,N_4799);
nand U5591 (N_5591,N_4813,N_4224);
xor U5592 (N_5592,N_4331,N_4441);
nand U5593 (N_5593,N_4319,N_4647);
nand U5594 (N_5594,N_4138,N_4552);
nor U5595 (N_5595,N_4791,N_4215);
nor U5596 (N_5596,N_4015,N_4231);
nand U5597 (N_5597,N_4232,N_4858);
or U5598 (N_5598,N_4368,N_4397);
nor U5599 (N_5599,N_4445,N_4519);
or U5600 (N_5600,N_4893,N_4215);
xor U5601 (N_5601,N_4672,N_4280);
xor U5602 (N_5602,N_4471,N_4222);
nand U5603 (N_5603,N_4376,N_4834);
nor U5604 (N_5604,N_4327,N_4220);
and U5605 (N_5605,N_4785,N_4247);
nor U5606 (N_5606,N_4085,N_4549);
nand U5607 (N_5607,N_4044,N_4686);
or U5608 (N_5608,N_4509,N_4769);
xor U5609 (N_5609,N_4663,N_4871);
nand U5610 (N_5610,N_4441,N_4280);
nand U5611 (N_5611,N_4446,N_4493);
or U5612 (N_5612,N_4900,N_4541);
nor U5613 (N_5613,N_4229,N_4779);
xor U5614 (N_5614,N_4828,N_4847);
nor U5615 (N_5615,N_4446,N_4436);
nor U5616 (N_5616,N_4023,N_4667);
nor U5617 (N_5617,N_4269,N_4681);
nand U5618 (N_5618,N_4975,N_4865);
or U5619 (N_5619,N_4221,N_4445);
and U5620 (N_5620,N_4916,N_4686);
nor U5621 (N_5621,N_4561,N_4386);
or U5622 (N_5622,N_4594,N_4991);
nor U5623 (N_5623,N_4371,N_4411);
nand U5624 (N_5624,N_4812,N_4700);
or U5625 (N_5625,N_4453,N_4687);
xnor U5626 (N_5626,N_4232,N_4412);
or U5627 (N_5627,N_4632,N_4686);
and U5628 (N_5628,N_4552,N_4409);
or U5629 (N_5629,N_4333,N_4896);
nand U5630 (N_5630,N_4583,N_4545);
nand U5631 (N_5631,N_4918,N_4866);
and U5632 (N_5632,N_4036,N_4708);
nand U5633 (N_5633,N_4298,N_4174);
xnor U5634 (N_5634,N_4025,N_4716);
or U5635 (N_5635,N_4832,N_4319);
xor U5636 (N_5636,N_4522,N_4727);
or U5637 (N_5637,N_4766,N_4374);
xnor U5638 (N_5638,N_4256,N_4031);
nand U5639 (N_5639,N_4743,N_4012);
nand U5640 (N_5640,N_4599,N_4199);
or U5641 (N_5641,N_4553,N_4493);
and U5642 (N_5642,N_4232,N_4969);
nand U5643 (N_5643,N_4629,N_4876);
or U5644 (N_5644,N_4645,N_4523);
and U5645 (N_5645,N_4364,N_4604);
nand U5646 (N_5646,N_4289,N_4708);
and U5647 (N_5647,N_4482,N_4011);
and U5648 (N_5648,N_4267,N_4602);
and U5649 (N_5649,N_4026,N_4934);
xnor U5650 (N_5650,N_4379,N_4411);
nor U5651 (N_5651,N_4823,N_4860);
and U5652 (N_5652,N_4950,N_4225);
and U5653 (N_5653,N_4191,N_4396);
or U5654 (N_5654,N_4075,N_4141);
or U5655 (N_5655,N_4298,N_4985);
nor U5656 (N_5656,N_4329,N_4960);
or U5657 (N_5657,N_4466,N_4980);
xnor U5658 (N_5658,N_4791,N_4517);
nor U5659 (N_5659,N_4466,N_4809);
nand U5660 (N_5660,N_4503,N_4769);
xor U5661 (N_5661,N_4988,N_4075);
nand U5662 (N_5662,N_4368,N_4262);
or U5663 (N_5663,N_4071,N_4029);
xor U5664 (N_5664,N_4862,N_4241);
nand U5665 (N_5665,N_4476,N_4412);
and U5666 (N_5666,N_4744,N_4805);
xnor U5667 (N_5667,N_4148,N_4241);
nor U5668 (N_5668,N_4154,N_4158);
nand U5669 (N_5669,N_4423,N_4123);
xor U5670 (N_5670,N_4512,N_4852);
xor U5671 (N_5671,N_4286,N_4008);
nor U5672 (N_5672,N_4589,N_4292);
nand U5673 (N_5673,N_4038,N_4840);
nand U5674 (N_5674,N_4084,N_4937);
nor U5675 (N_5675,N_4025,N_4806);
nor U5676 (N_5676,N_4593,N_4968);
nand U5677 (N_5677,N_4307,N_4957);
nand U5678 (N_5678,N_4303,N_4343);
nand U5679 (N_5679,N_4024,N_4342);
or U5680 (N_5680,N_4668,N_4693);
or U5681 (N_5681,N_4828,N_4254);
nor U5682 (N_5682,N_4750,N_4796);
or U5683 (N_5683,N_4232,N_4510);
xor U5684 (N_5684,N_4249,N_4772);
and U5685 (N_5685,N_4379,N_4211);
nand U5686 (N_5686,N_4881,N_4871);
nand U5687 (N_5687,N_4116,N_4108);
and U5688 (N_5688,N_4463,N_4889);
xor U5689 (N_5689,N_4185,N_4360);
xnor U5690 (N_5690,N_4900,N_4490);
xnor U5691 (N_5691,N_4874,N_4609);
and U5692 (N_5692,N_4209,N_4601);
nor U5693 (N_5693,N_4947,N_4009);
nor U5694 (N_5694,N_4759,N_4276);
nor U5695 (N_5695,N_4270,N_4166);
xnor U5696 (N_5696,N_4304,N_4687);
or U5697 (N_5697,N_4591,N_4266);
nor U5698 (N_5698,N_4717,N_4888);
nor U5699 (N_5699,N_4736,N_4305);
nand U5700 (N_5700,N_4401,N_4048);
and U5701 (N_5701,N_4840,N_4428);
or U5702 (N_5702,N_4795,N_4426);
xor U5703 (N_5703,N_4773,N_4050);
and U5704 (N_5704,N_4238,N_4092);
and U5705 (N_5705,N_4172,N_4122);
and U5706 (N_5706,N_4100,N_4458);
nand U5707 (N_5707,N_4270,N_4146);
or U5708 (N_5708,N_4221,N_4328);
nand U5709 (N_5709,N_4246,N_4178);
and U5710 (N_5710,N_4739,N_4863);
xnor U5711 (N_5711,N_4453,N_4059);
or U5712 (N_5712,N_4585,N_4147);
or U5713 (N_5713,N_4465,N_4404);
nand U5714 (N_5714,N_4478,N_4299);
nor U5715 (N_5715,N_4772,N_4118);
and U5716 (N_5716,N_4958,N_4039);
and U5717 (N_5717,N_4403,N_4191);
xor U5718 (N_5718,N_4791,N_4027);
or U5719 (N_5719,N_4010,N_4297);
nor U5720 (N_5720,N_4296,N_4370);
xnor U5721 (N_5721,N_4834,N_4805);
and U5722 (N_5722,N_4321,N_4761);
nor U5723 (N_5723,N_4036,N_4349);
nand U5724 (N_5724,N_4416,N_4542);
and U5725 (N_5725,N_4443,N_4957);
nor U5726 (N_5726,N_4435,N_4166);
xor U5727 (N_5727,N_4675,N_4249);
or U5728 (N_5728,N_4351,N_4457);
and U5729 (N_5729,N_4430,N_4261);
or U5730 (N_5730,N_4718,N_4935);
nor U5731 (N_5731,N_4509,N_4578);
nor U5732 (N_5732,N_4416,N_4861);
nand U5733 (N_5733,N_4955,N_4227);
or U5734 (N_5734,N_4916,N_4575);
and U5735 (N_5735,N_4264,N_4765);
and U5736 (N_5736,N_4250,N_4961);
nor U5737 (N_5737,N_4161,N_4969);
or U5738 (N_5738,N_4997,N_4986);
and U5739 (N_5739,N_4589,N_4627);
xor U5740 (N_5740,N_4110,N_4533);
and U5741 (N_5741,N_4536,N_4583);
xnor U5742 (N_5742,N_4156,N_4395);
nand U5743 (N_5743,N_4435,N_4533);
and U5744 (N_5744,N_4223,N_4632);
and U5745 (N_5745,N_4759,N_4863);
or U5746 (N_5746,N_4472,N_4242);
nand U5747 (N_5747,N_4135,N_4826);
or U5748 (N_5748,N_4642,N_4824);
and U5749 (N_5749,N_4397,N_4206);
and U5750 (N_5750,N_4213,N_4538);
nor U5751 (N_5751,N_4672,N_4702);
or U5752 (N_5752,N_4766,N_4380);
xnor U5753 (N_5753,N_4217,N_4512);
xnor U5754 (N_5754,N_4179,N_4617);
nor U5755 (N_5755,N_4718,N_4649);
or U5756 (N_5756,N_4797,N_4416);
nand U5757 (N_5757,N_4686,N_4478);
xnor U5758 (N_5758,N_4362,N_4719);
nor U5759 (N_5759,N_4500,N_4617);
xnor U5760 (N_5760,N_4961,N_4356);
and U5761 (N_5761,N_4095,N_4138);
xnor U5762 (N_5762,N_4398,N_4600);
nand U5763 (N_5763,N_4477,N_4600);
or U5764 (N_5764,N_4517,N_4189);
nand U5765 (N_5765,N_4900,N_4651);
xnor U5766 (N_5766,N_4146,N_4213);
or U5767 (N_5767,N_4848,N_4979);
nor U5768 (N_5768,N_4740,N_4176);
and U5769 (N_5769,N_4836,N_4269);
or U5770 (N_5770,N_4737,N_4196);
nor U5771 (N_5771,N_4622,N_4798);
and U5772 (N_5772,N_4089,N_4573);
and U5773 (N_5773,N_4005,N_4581);
nor U5774 (N_5774,N_4690,N_4112);
or U5775 (N_5775,N_4237,N_4290);
nand U5776 (N_5776,N_4471,N_4983);
xnor U5777 (N_5777,N_4562,N_4515);
xnor U5778 (N_5778,N_4489,N_4632);
xnor U5779 (N_5779,N_4480,N_4107);
nand U5780 (N_5780,N_4247,N_4451);
nand U5781 (N_5781,N_4062,N_4632);
or U5782 (N_5782,N_4194,N_4447);
xor U5783 (N_5783,N_4000,N_4735);
or U5784 (N_5784,N_4634,N_4635);
nand U5785 (N_5785,N_4780,N_4193);
nor U5786 (N_5786,N_4918,N_4470);
nor U5787 (N_5787,N_4077,N_4893);
nor U5788 (N_5788,N_4221,N_4251);
or U5789 (N_5789,N_4356,N_4661);
xnor U5790 (N_5790,N_4471,N_4913);
nand U5791 (N_5791,N_4033,N_4665);
xnor U5792 (N_5792,N_4209,N_4232);
nand U5793 (N_5793,N_4854,N_4329);
and U5794 (N_5794,N_4652,N_4174);
xnor U5795 (N_5795,N_4431,N_4682);
nand U5796 (N_5796,N_4712,N_4390);
xor U5797 (N_5797,N_4619,N_4388);
nor U5798 (N_5798,N_4326,N_4400);
or U5799 (N_5799,N_4970,N_4289);
xor U5800 (N_5800,N_4340,N_4210);
nor U5801 (N_5801,N_4264,N_4705);
nor U5802 (N_5802,N_4510,N_4587);
nor U5803 (N_5803,N_4146,N_4385);
and U5804 (N_5804,N_4252,N_4485);
nor U5805 (N_5805,N_4906,N_4274);
and U5806 (N_5806,N_4973,N_4287);
and U5807 (N_5807,N_4689,N_4692);
nor U5808 (N_5808,N_4299,N_4562);
nand U5809 (N_5809,N_4206,N_4693);
nand U5810 (N_5810,N_4960,N_4095);
nor U5811 (N_5811,N_4930,N_4657);
xor U5812 (N_5812,N_4073,N_4491);
and U5813 (N_5813,N_4377,N_4868);
and U5814 (N_5814,N_4371,N_4660);
and U5815 (N_5815,N_4335,N_4374);
and U5816 (N_5816,N_4194,N_4848);
xnor U5817 (N_5817,N_4667,N_4876);
or U5818 (N_5818,N_4083,N_4590);
nand U5819 (N_5819,N_4545,N_4633);
xnor U5820 (N_5820,N_4554,N_4397);
xnor U5821 (N_5821,N_4283,N_4471);
nor U5822 (N_5822,N_4421,N_4949);
or U5823 (N_5823,N_4258,N_4142);
nand U5824 (N_5824,N_4256,N_4726);
xnor U5825 (N_5825,N_4832,N_4896);
xnor U5826 (N_5826,N_4829,N_4386);
xor U5827 (N_5827,N_4837,N_4261);
and U5828 (N_5828,N_4785,N_4897);
or U5829 (N_5829,N_4293,N_4789);
xor U5830 (N_5830,N_4496,N_4121);
nand U5831 (N_5831,N_4329,N_4031);
or U5832 (N_5832,N_4001,N_4280);
or U5833 (N_5833,N_4921,N_4805);
nand U5834 (N_5834,N_4769,N_4483);
nand U5835 (N_5835,N_4338,N_4420);
nand U5836 (N_5836,N_4607,N_4113);
nand U5837 (N_5837,N_4363,N_4988);
and U5838 (N_5838,N_4885,N_4844);
or U5839 (N_5839,N_4583,N_4051);
nor U5840 (N_5840,N_4553,N_4682);
and U5841 (N_5841,N_4838,N_4474);
nor U5842 (N_5842,N_4489,N_4129);
nand U5843 (N_5843,N_4367,N_4906);
or U5844 (N_5844,N_4366,N_4564);
and U5845 (N_5845,N_4426,N_4565);
xor U5846 (N_5846,N_4505,N_4361);
xnor U5847 (N_5847,N_4753,N_4862);
nand U5848 (N_5848,N_4198,N_4320);
nand U5849 (N_5849,N_4649,N_4120);
nand U5850 (N_5850,N_4793,N_4940);
xor U5851 (N_5851,N_4060,N_4148);
nand U5852 (N_5852,N_4170,N_4250);
nor U5853 (N_5853,N_4366,N_4195);
and U5854 (N_5854,N_4387,N_4893);
and U5855 (N_5855,N_4553,N_4657);
xor U5856 (N_5856,N_4400,N_4229);
or U5857 (N_5857,N_4547,N_4221);
nor U5858 (N_5858,N_4423,N_4346);
nor U5859 (N_5859,N_4161,N_4009);
and U5860 (N_5860,N_4500,N_4149);
nand U5861 (N_5861,N_4213,N_4584);
nand U5862 (N_5862,N_4415,N_4951);
or U5863 (N_5863,N_4139,N_4396);
or U5864 (N_5864,N_4835,N_4487);
or U5865 (N_5865,N_4602,N_4392);
xnor U5866 (N_5866,N_4240,N_4107);
nor U5867 (N_5867,N_4655,N_4106);
nor U5868 (N_5868,N_4737,N_4286);
nand U5869 (N_5869,N_4817,N_4336);
nor U5870 (N_5870,N_4546,N_4948);
nand U5871 (N_5871,N_4749,N_4166);
or U5872 (N_5872,N_4533,N_4463);
nand U5873 (N_5873,N_4286,N_4383);
xnor U5874 (N_5874,N_4780,N_4043);
or U5875 (N_5875,N_4984,N_4039);
or U5876 (N_5876,N_4598,N_4632);
nand U5877 (N_5877,N_4086,N_4345);
or U5878 (N_5878,N_4953,N_4534);
xor U5879 (N_5879,N_4400,N_4102);
or U5880 (N_5880,N_4168,N_4077);
nor U5881 (N_5881,N_4812,N_4161);
and U5882 (N_5882,N_4291,N_4290);
nand U5883 (N_5883,N_4388,N_4978);
nand U5884 (N_5884,N_4084,N_4262);
or U5885 (N_5885,N_4733,N_4076);
nand U5886 (N_5886,N_4897,N_4215);
nor U5887 (N_5887,N_4731,N_4178);
or U5888 (N_5888,N_4125,N_4858);
xor U5889 (N_5889,N_4846,N_4344);
and U5890 (N_5890,N_4397,N_4624);
xor U5891 (N_5891,N_4803,N_4009);
nor U5892 (N_5892,N_4348,N_4965);
xor U5893 (N_5893,N_4964,N_4931);
and U5894 (N_5894,N_4422,N_4099);
and U5895 (N_5895,N_4142,N_4890);
nor U5896 (N_5896,N_4907,N_4183);
xor U5897 (N_5897,N_4993,N_4191);
xnor U5898 (N_5898,N_4217,N_4061);
or U5899 (N_5899,N_4511,N_4680);
or U5900 (N_5900,N_4336,N_4250);
xnor U5901 (N_5901,N_4845,N_4169);
xor U5902 (N_5902,N_4126,N_4958);
nor U5903 (N_5903,N_4788,N_4952);
and U5904 (N_5904,N_4646,N_4741);
and U5905 (N_5905,N_4939,N_4497);
or U5906 (N_5906,N_4640,N_4908);
nand U5907 (N_5907,N_4009,N_4623);
xor U5908 (N_5908,N_4576,N_4211);
or U5909 (N_5909,N_4348,N_4251);
or U5910 (N_5910,N_4792,N_4849);
xnor U5911 (N_5911,N_4336,N_4507);
nand U5912 (N_5912,N_4622,N_4650);
nor U5913 (N_5913,N_4273,N_4468);
xnor U5914 (N_5914,N_4138,N_4051);
and U5915 (N_5915,N_4929,N_4906);
nand U5916 (N_5916,N_4903,N_4956);
or U5917 (N_5917,N_4870,N_4707);
xnor U5918 (N_5918,N_4367,N_4399);
and U5919 (N_5919,N_4422,N_4019);
or U5920 (N_5920,N_4404,N_4645);
xor U5921 (N_5921,N_4554,N_4822);
xor U5922 (N_5922,N_4130,N_4213);
xor U5923 (N_5923,N_4917,N_4780);
nor U5924 (N_5924,N_4675,N_4662);
or U5925 (N_5925,N_4194,N_4654);
or U5926 (N_5926,N_4300,N_4194);
nor U5927 (N_5927,N_4341,N_4720);
nand U5928 (N_5928,N_4739,N_4718);
nand U5929 (N_5929,N_4151,N_4902);
xor U5930 (N_5930,N_4928,N_4872);
nor U5931 (N_5931,N_4694,N_4947);
or U5932 (N_5932,N_4530,N_4557);
xnor U5933 (N_5933,N_4681,N_4718);
nor U5934 (N_5934,N_4339,N_4479);
and U5935 (N_5935,N_4995,N_4225);
and U5936 (N_5936,N_4457,N_4250);
nand U5937 (N_5937,N_4362,N_4311);
or U5938 (N_5938,N_4165,N_4921);
or U5939 (N_5939,N_4255,N_4051);
and U5940 (N_5940,N_4109,N_4102);
or U5941 (N_5941,N_4206,N_4652);
xor U5942 (N_5942,N_4082,N_4242);
nand U5943 (N_5943,N_4025,N_4305);
nand U5944 (N_5944,N_4710,N_4842);
and U5945 (N_5945,N_4912,N_4224);
or U5946 (N_5946,N_4738,N_4913);
or U5947 (N_5947,N_4602,N_4769);
nor U5948 (N_5948,N_4271,N_4579);
xnor U5949 (N_5949,N_4550,N_4690);
xnor U5950 (N_5950,N_4716,N_4180);
nand U5951 (N_5951,N_4435,N_4806);
and U5952 (N_5952,N_4207,N_4400);
nor U5953 (N_5953,N_4171,N_4098);
nand U5954 (N_5954,N_4682,N_4346);
nand U5955 (N_5955,N_4903,N_4752);
or U5956 (N_5956,N_4740,N_4386);
and U5957 (N_5957,N_4343,N_4498);
or U5958 (N_5958,N_4193,N_4409);
and U5959 (N_5959,N_4167,N_4765);
xor U5960 (N_5960,N_4814,N_4205);
or U5961 (N_5961,N_4256,N_4373);
nand U5962 (N_5962,N_4601,N_4249);
nand U5963 (N_5963,N_4281,N_4456);
and U5964 (N_5964,N_4057,N_4106);
or U5965 (N_5965,N_4411,N_4855);
xor U5966 (N_5966,N_4929,N_4142);
nand U5967 (N_5967,N_4027,N_4405);
xor U5968 (N_5968,N_4072,N_4897);
or U5969 (N_5969,N_4258,N_4338);
and U5970 (N_5970,N_4407,N_4693);
xnor U5971 (N_5971,N_4321,N_4157);
and U5972 (N_5972,N_4640,N_4923);
nor U5973 (N_5973,N_4466,N_4340);
or U5974 (N_5974,N_4377,N_4301);
xor U5975 (N_5975,N_4399,N_4985);
or U5976 (N_5976,N_4186,N_4233);
xnor U5977 (N_5977,N_4232,N_4761);
and U5978 (N_5978,N_4114,N_4698);
nand U5979 (N_5979,N_4312,N_4535);
nor U5980 (N_5980,N_4865,N_4866);
and U5981 (N_5981,N_4330,N_4518);
and U5982 (N_5982,N_4860,N_4774);
or U5983 (N_5983,N_4750,N_4240);
and U5984 (N_5984,N_4035,N_4633);
or U5985 (N_5985,N_4322,N_4402);
nand U5986 (N_5986,N_4990,N_4458);
nand U5987 (N_5987,N_4735,N_4002);
or U5988 (N_5988,N_4755,N_4215);
nor U5989 (N_5989,N_4650,N_4201);
and U5990 (N_5990,N_4531,N_4555);
and U5991 (N_5991,N_4365,N_4793);
and U5992 (N_5992,N_4333,N_4780);
and U5993 (N_5993,N_4628,N_4444);
nand U5994 (N_5994,N_4693,N_4681);
nor U5995 (N_5995,N_4552,N_4511);
or U5996 (N_5996,N_4595,N_4275);
and U5997 (N_5997,N_4459,N_4751);
nor U5998 (N_5998,N_4396,N_4675);
nor U5999 (N_5999,N_4611,N_4947);
xor U6000 (N_6000,N_5289,N_5993);
nor U6001 (N_6001,N_5334,N_5271);
xor U6002 (N_6002,N_5957,N_5238);
or U6003 (N_6003,N_5021,N_5306);
and U6004 (N_6004,N_5883,N_5694);
nor U6005 (N_6005,N_5661,N_5761);
nand U6006 (N_6006,N_5374,N_5878);
and U6007 (N_6007,N_5132,N_5783);
nand U6008 (N_6008,N_5253,N_5862);
and U6009 (N_6009,N_5102,N_5699);
and U6010 (N_6010,N_5764,N_5674);
nor U6011 (N_6011,N_5397,N_5656);
xor U6012 (N_6012,N_5398,N_5851);
xor U6013 (N_6013,N_5503,N_5210);
nand U6014 (N_6014,N_5229,N_5137);
nand U6015 (N_6015,N_5975,N_5319);
nor U6016 (N_6016,N_5314,N_5358);
and U6017 (N_6017,N_5574,N_5205);
and U6018 (N_6018,N_5537,N_5390);
nor U6019 (N_6019,N_5618,N_5192);
xnor U6020 (N_6020,N_5668,N_5465);
and U6021 (N_6021,N_5447,N_5295);
xor U6022 (N_6022,N_5258,N_5597);
and U6023 (N_6023,N_5990,N_5435);
xnor U6024 (N_6024,N_5810,N_5728);
and U6025 (N_6025,N_5543,N_5903);
nand U6026 (N_6026,N_5542,N_5348);
nor U6027 (N_6027,N_5167,N_5235);
or U6028 (N_6028,N_5785,N_5058);
xor U6029 (N_6029,N_5995,N_5458);
nor U6030 (N_6030,N_5377,N_5015);
xor U6031 (N_6031,N_5584,N_5480);
or U6032 (N_6032,N_5301,N_5476);
nand U6033 (N_6033,N_5557,N_5628);
or U6034 (N_6034,N_5240,N_5298);
nor U6035 (N_6035,N_5988,N_5360);
xor U6036 (N_6036,N_5259,N_5687);
xnor U6037 (N_6037,N_5912,N_5863);
or U6038 (N_6038,N_5572,N_5974);
nand U6039 (N_6039,N_5573,N_5620);
and U6040 (N_6040,N_5006,N_5925);
or U6041 (N_6041,N_5731,N_5062);
or U6042 (N_6042,N_5324,N_5945);
nor U6043 (N_6043,N_5412,N_5272);
xor U6044 (N_6044,N_5418,N_5855);
nand U6045 (N_6045,N_5313,N_5844);
nor U6046 (N_6046,N_5293,N_5742);
nand U6047 (N_6047,N_5588,N_5905);
nand U6048 (N_6048,N_5886,N_5089);
nand U6049 (N_6049,N_5485,N_5890);
and U6050 (N_6050,N_5926,N_5305);
or U6051 (N_6051,N_5516,N_5660);
or U6052 (N_6052,N_5913,N_5497);
nor U6053 (N_6053,N_5194,N_5378);
nor U6054 (N_6054,N_5868,N_5663);
nor U6055 (N_6055,N_5749,N_5532);
xnor U6056 (N_6056,N_5530,N_5416);
xnor U6057 (N_6057,N_5682,N_5357);
or U6058 (N_6058,N_5023,N_5985);
or U6059 (N_6059,N_5239,N_5846);
nand U6060 (N_6060,N_5018,N_5548);
or U6061 (N_6061,N_5819,N_5153);
nand U6062 (N_6062,N_5488,N_5747);
nor U6063 (N_6063,N_5343,N_5828);
nor U6064 (N_6064,N_5796,N_5623);
and U6065 (N_6065,N_5202,N_5437);
nor U6066 (N_6066,N_5899,N_5406);
nand U6067 (N_6067,N_5347,N_5440);
xnor U6068 (N_6068,N_5336,N_5333);
nor U6069 (N_6069,N_5723,N_5382);
nand U6070 (N_6070,N_5311,N_5455);
or U6071 (N_6071,N_5637,N_5754);
nand U6072 (N_6072,N_5188,N_5466);
or U6073 (N_6073,N_5748,N_5320);
xor U6074 (N_6074,N_5967,N_5185);
nand U6075 (N_6075,N_5951,N_5136);
or U6076 (N_6076,N_5077,N_5780);
and U6077 (N_6077,N_5395,N_5091);
nand U6078 (N_6078,N_5602,N_5627);
nand U6079 (N_6079,N_5198,N_5586);
or U6080 (N_6080,N_5702,N_5231);
nor U6081 (N_6081,N_5340,N_5156);
nor U6082 (N_6082,N_5902,N_5095);
or U6083 (N_6083,N_5714,N_5287);
and U6084 (N_6084,N_5415,N_5987);
and U6085 (N_6085,N_5977,N_5171);
xnor U6086 (N_6086,N_5473,N_5732);
and U6087 (N_6087,N_5138,N_5381);
nor U6088 (N_6088,N_5545,N_5341);
nand U6089 (N_6089,N_5809,N_5789);
nand U6090 (N_6090,N_5757,N_5936);
nand U6091 (N_6091,N_5034,N_5647);
nor U6092 (N_6092,N_5982,N_5587);
xnor U6093 (N_6093,N_5759,N_5555);
nand U6094 (N_6094,N_5017,N_5529);
xor U6095 (N_6095,N_5216,N_5133);
and U6096 (N_6096,N_5619,N_5818);
xor U6097 (N_6097,N_5048,N_5280);
or U6098 (N_6098,N_5436,N_5218);
nand U6099 (N_6099,N_5921,N_5459);
nor U6100 (N_6100,N_5019,N_5870);
or U6101 (N_6101,N_5472,N_5711);
or U6102 (N_6102,N_5965,N_5369);
or U6103 (N_6103,N_5014,N_5389);
nand U6104 (N_6104,N_5877,N_5182);
xnor U6105 (N_6105,N_5139,N_5332);
and U6106 (N_6106,N_5283,N_5431);
or U6107 (N_6107,N_5743,N_5492);
nand U6108 (N_6108,N_5859,N_5986);
xor U6109 (N_6109,N_5380,N_5786);
and U6110 (N_6110,N_5898,N_5676);
nor U6111 (N_6111,N_5457,N_5103);
nor U6112 (N_6112,N_5452,N_5801);
or U6113 (N_6113,N_5197,N_5422);
or U6114 (N_6114,N_5595,N_5356);
nand U6115 (N_6115,N_5693,N_5312);
nor U6116 (N_6116,N_5610,N_5812);
xor U6117 (N_6117,N_5657,N_5330);
xnor U6118 (N_6118,N_5142,N_5439);
and U6119 (N_6119,N_5716,N_5104);
nand U6120 (N_6120,N_5424,N_5566);
and U6121 (N_6121,N_5125,N_5063);
nand U6122 (N_6122,N_5551,N_5164);
and U6123 (N_6123,N_5052,N_5463);
nor U6124 (N_6124,N_5213,N_5897);
nor U6125 (N_6125,N_5950,N_5384);
or U6126 (N_6126,N_5867,N_5547);
nor U6127 (N_6127,N_5730,N_5546);
xnor U6128 (N_6128,N_5604,N_5001);
nor U6129 (N_6129,N_5413,N_5371);
or U6130 (N_6130,N_5710,N_5487);
nor U6131 (N_6131,N_5462,N_5166);
xnor U6132 (N_6132,N_5729,N_5174);
xor U6133 (N_6133,N_5746,N_5217);
xor U6134 (N_6134,N_5518,N_5854);
and U6135 (N_6135,N_5051,N_5172);
xnor U6136 (N_6136,N_5069,N_5454);
nand U6137 (N_6137,N_5740,N_5214);
xnor U6138 (N_6138,N_5425,N_5733);
xnor U6139 (N_6139,N_5300,N_5848);
xor U6140 (N_6140,N_5820,N_5549);
nand U6141 (N_6141,N_5328,N_5071);
nor U6142 (N_6142,N_5112,N_5852);
nand U6143 (N_6143,N_5046,N_5923);
or U6144 (N_6144,N_5241,N_5351);
nand U6145 (N_6145,N_5495,N_5885);
xnor U6146 (N_6146,N_5024,N_5326);
nor U6147 (N_6147,N_5725,N_5621);
xor U6148 (N_6148,N_5499,N_5858);
or U6149 (N_6149,N_5653,N_5344);
and U6150 (N_6150,N_5232,N_5254);
nor U6151 (N_6151,N_5101,N_5304);
and U6152 (N_6152,N_5163,N_5683);
and U6153 (N_6153,N_5813,N_5411);
nor U6154 (N_6154,N_5004,N_5949);
nor U6155 (N_6155,N_5094,N_5270);
and U6156 (N_6156,N_5582,N_5806);
nand U6157 (N_6157,N_5726,N_5294);
and U6158 (N_6158,N_5989,N_5449);
xnor U6159 (N_6159,N_5141,N_5636);
xnor U6160 (N_6160,N_5744,N_5453);
nand U6161 (N_6161,N_5028,N_5790);
or U6162 (N_6162,N_5792,N_5505);
and U6163 (N_6163,N_5494,N_5408);
nand U6164 (N_6164,N_5734,N_5802);
or U6165 (N_6165,N_5130,N_5622);
nand U6166 (N_6166,N_5044,N_5266);
and U6167 (N_6167,N_5978,N_5822);
nor U6168 (N_6168,N_5331,N_5521);
nand U6169 (N_6169,N_5670,N_5310);
nor U6170 (N_6170,N_5121,N_5207);
xor U6171 (N_6171,N_5404,N_5948);
nand U6172 (N_6172,N_5834,N_5168);
xor U6173 (N_6173,N_5662,N_5376);
xor U6174 (N_6174,N_5980,N_5025);
nor U6175 (N_6175,N_5659,N_5970);
and U6176 (N_6176,N_5506,N_5409);
or U6177 (N_6177,N_5955,N_5160);
or U6178 (N_6178,N_5379,N_5692);
xor U6179 (N_6179,N_5013,N_5771);
nand U6180 (N_6180,N_5486,N_5803);
and U6181 (N_6181,N_5154,N_5029);
xor U6182 (N_6182,N_5924,N_5918);
or U6183 (N_6183,N_5307,N_5644);
or U6184 (N_6184,N_5383,N_5276);
or U6185 (N_6185,N_5741,N_5129);
nor U6186 (N_6186,N_5143,N_5664);
nor U6187 (N_6187,N_5109,N_5027);
or U6188 (N_6188,N_5170,N_5118);
and U6189 (N_6189,N_5928,N_5673);
and U6190 (N_6190,N_5262,N_5072);
nand U6191 (N_6191,N_5609,N_5220);
nand U6192 (N_6192,N_5189,N_5954);
xor U6193 (N_6193,N_5501,N_5541);
or U6194 (N_6194,N_5632,N_5538);
nand U6195 (N_6195,N_5932,N_5115);
nor U6196 (N_6196,N_5147,N_5322);
and U6197 (N_6197,N_5490,N_5784);
nand U6198 (N_6198,N_5626,N_5433);
xnor U6199 (N_6199,N_5349,N_5895);
xnor U6200 (N_6200,N_5646,N_5116);
or U6201 (N_6201,N_5215,N_5363);
nand U6202 (N_6202,N_5561,N_5208);
or U6203 (N_6203,N_5066,N_5942);
or U6204 (N_6204,N_5688,N_5169);
or U6205 (N_6205,N_5624,N_5098);
or U6206 (N_6206,N_5339,N_5593);
nor U6207 (N_6207,N_5756,N_5869);
and U6208 (N_6208,N_5887,N_5434);
and U6209 (N_6209,N_5427,N_5900);
nand U6210 (N_6210,N_5005,N_5735);
and U6211 (N_6211,N_5944,N_5087);
and U6212 (N_6212,N_5522,N_5601);
and U6213 (N_6213,N_5346,N_5826);
and U6214 (N_6214,N_5697,N_5829);
nand U6215 (N_6215,N_5658,N_5464);
xor U6216 (N_6216,N_5263,N_5362);
nor U6217 (N_6217,N_5976,N_5365);
nor U6218 (N_6218,N_5387,N_5888);
nand U6219 (N_6219,N_5559,N_5686);
or U6220 (N_6220,N_5669,N_5583);
xnor U6221 (N_6221,N_5173,N_5817);
xnor U6222 (N_6222,N_5196,N_5513);
nor U6223 (N_6223,N_5691,N_5643);
xnor U6224 (N_6224,N_5477,N_5816);
nand U6225 (N_6225,N_5934,N_5782);
or U6226 (N_6226,N_5614,N_5078);
or U6227 (N_6227,N_5850,N_5874);
nand U6228 (N_6228,N_5605,N_5909);
nor U6229 (N_6229,N_5649,N_5893);
xnor U6230 (N_6230,N_5396,N_5685);
nor U6231 (N_6231,N_5251,N_5640);
xor U6232 (N_6232,N_5766,N_5318);
and U6233 (N_6233,N_5760,N_5002);
and U6234 (N_6234,N_5811,N_5080);
nand U6235 (N_6235,N_5842,N_5832);
or U6236 (N_6236,N_5243,N_5041);
xnor U6237 (N_6237,N_5500,N_5372);
or U6238 (N_6238,N_5625,N_5752);
or U6239 (N_6239,N_5474,N_5865);
or U6240 (N_6240,N_5630,N_5979);
and U6241 (N_6241,N_5290,N_5645);
or U6242 (N_6242,N_5966,N_5158);
nand U6243 (N_6243,N_5335,N_5338);
xor U6244 (N_6244,N_5600,N_5421);
nor U6245 (N_6245,N_5799,N_5099);
nand U6246 (N_6246,N_5068,N_5468);
or U6247 (N_6247,N_5991,N_5345);
and U6248 (N_6248,N_5519,N_5193);
and U6249 (N_6249,N_5680,N_5391);
nand U6250 (N_6250,N_5327,N_5157);
and U6251 (N_6251,N_5833,N_5525);
or U6252 (N_6252,N_5581,N_5149);
nand U6253 (N_6253,N_5718,N_5352);
nor U6254 (N_6254,N_5892,N_5508);
nor U6255 (N_6255,N_5469,N_5234);
nor U6256 (N_6256,N_5140,N_5835);
xnor U6257 (N_6257,N_5994,N_5767);
and U6258 (N_6258,N_5727,N_5775);
and U6259 (N_6259,N_5076,N_5373);
or U6260 (N_6260,N_5315,N_5049);
nand U6261 (N_6261,N_5788,N_5800);
nor U6262 (N_6262,N_5984,N_5633);
nor U6263 (N_6263,N_5405,N_5032);
nor U6264 (N_6264,N_5221,N_5146);
xnor U6265 (N_6265,N_5613,N_5774);
nor U6266 (N_6266,N_5642,N_5755);
nor U6267 (N_6267,N_5438,N_5444);
xor U6268 (N_6268,N_5126,N_5779);
xnor U6269 (N_6269,N_5776,N_5941);
or U6270 (N_6270,N_5033,N_5407);
nand U6271 (N_6271,N_5496,N_5317);
or U6272 (N_6272,N_5915,N_5297);
or U6273 (N_6273,N_5079,N_5947);
nand U6274 (N_6274,N_5589,N_5219);
and U6275 (N_6275,N_5222,N_5178);
xor U6276 (N_6276,N_5471,N_5249);
nand U6277 (N_6277,N_5629,N_5399);
nor U6278 (N_6278,N_5187,N_5113);
and U6279 (N_6279,N_5678,N_5961);
or U6280 (N_6280,N_5707,N_5873);
nor U6281 (N_6281,N_5814,N_5599);
xnor U6282 (N_6282,N_5291,N_5212);
and U6283 (N_6283,N_5666,N_5108);
or U6284 (N_6284,N_5969,N_5000);
and U6285 (N_6285,N_5914,N_5651);
nand U6286 (N_6286,N_5768,N_5594);
nand U6287 (N_6287,N_5491,N_5361);
and U6288 (N_6288,N_5681,N_5715);
or U6289 (N_6289,N_5511,N_5482);
and U6290 (N_6290,N_5917,N_5264);
nor U6291 (N_6291,N_5807,N_5540);
or U6292 (N_6292,N_5105,N_5539);
or U6293 (N_6293,N_5962,N_5042);
nand U6294 (N_6294,N_5904,N_5073);
or U6295 (N_6295,N_5823,N_5889);
or U6296 (N_6296,N_5713,N_5571);
xor U6297 (N_6297,N_5035,N_5781);
and U6298 (N_6298,N_5866,N_5879);
nor U6299 (N_6299,N_5751,N_5534);
nand U6300 (N_6300,N_5181,N_5908);
nor U6301 (N_6301,N_5916,N_5445);
nand U6302 (N_6302,N_5467,N_5203);
and U6303 (N_6303,N_5804,N_5920);
nand U6304 (N_6304,N_5708,N_5242);
nand U6305 (N_6305,N_5825,N_5576);
or U6306 (N_6306,N_5145,N_5689);
nor U6307 (N_6307,N_5403,N_5281);
nor U6308 (N_6308,N_5054,N_5872);
nor U6309 (N_6309,N_5608,N_5763);
and U6310 (N_6310,N_5321,N_5225);
and U6311 (N_6311,N_5736,N_5648);
or U6312 (N_6312,N_5086,N_5388);
nor U6313 (N_6313,N_5296,N_5798);
nor U6314 (N_6314,N_5512,N_5400);
or U6315 (N_6315,N_5690,N_5498);
nor U6316 (N_6316,N_5151,N_5841);
and U6317 (N_6317,N_5745,N_5123);
nand U6318 (N_6318,N_5180,N_5053);
or U6319 (N_6319,N_5550,N_5638);
or U6320 (N_6320,N_5162,N_5876);
or U6321 (N_6321,N_5010,N_5122);
and U6322 (N_6322,N_5256,N_5420);
nor U6323 (N_6323,N_5223,N_5364);
xnor U6324 (N_6324,N_5161,N_5808);
nor U6325 (N_6325,N_5769,N_5617);
xnor U6326 (N_6326,N_5045,N_5758);
and U6327 (N_6327,N_5201,N_5284);
or U6328 (N_6328,N_5943,N_5450);
or U6329 (N_6329,N_5937,N_5737);
nor U6330 (N_6330,N_5773,N_5679);
nand U6331 (N_6331,N_5698,N_5930);
nand U6332 (N_6332,N_5960,N_5037);
and U6333 (N_6333,N_5940,N_5939);
and U6334 (N_6334,N_5704,N_5131);
nor U6335 (N_6335,N_5836,N_5533);
and U6336 (N_6336,N_5938,N_5128);
nand U6337 (N_6337,N_5393,N_5631);
nand U6338 (N_6338,N_5199,N_5815);
and U6339 (N_6339,N_5502,N_5777);
nor U6340 (N_6340,N_5721,N_5209);
and U6341 (N_6341,N_5176,N_5120);
nand U6342 (N_6342,N_5585,N_5910);
xnor U6343 (N_6343,N_5047,N_5523);
nor U6344 (N_6344,N_5111,N_5838);
xor U6345 (N_6345,N_5857,N_5448);
nand U6346 (N_6346,N_5119,N_5368);
nor U6347 (N_6347,N_5303,N_5088);
nand U6348 (N_6348,N_5275,N_5059);
and U6349 (N_6349,N_5515,N_5267);
nor U6350 (N_6350,N_5709,N_5370);
nand U6351 (N_6351,N_5478,N_5881);
xnor U6352 (N_6352,N_5580,N_5292);
and U6353 (N_6353,N_5402,N_5279);
nand U6354 (N_6354,N_5607,N_5061);
nor U6355 (N_6355,N_5853,N_5135);
and U6356 (N_6356,N_5165,N_5972);
nand U6357 (N_6357,N_5355,N_5639);
nand U6358 (N_6358,N_5206,N_5724);
nand U6359 (N_6359,N_5544,N_5750);
and U6360 (N_6360,N_5514,N_5959);
or U6361 (N_6361,N_5675,N_5536);
and U6362 (N_6362,N_5483,N_5410);
xor U6363 (N_6363,N_5252,N_5030);
xor U6364 (N_6364,N_5057,N_5845);
xor U6365 (N_6365,N_5762,N_5884);
nor U6366 (N_6366,N_5155,N_5008);
or U6367 (N_6367,N_5430,N_5020);
nor U6368 (N_6368,N_5998,N_5067);
nor U6369 (N_6369,N_5794,N_5861);
or U6370 (N_6370,N_5106,N_5983);
nand U6371 (N_6371,N_5075,N_5230);
nand U6372 (N_6372,N_5428,N_5302);
and U6373 (N_6373,N_5520,N_5596);
and U6374 (N_6374,N_5824,N_5246);
nand U6375 (N_6375,N_5720,N_5083);
or U6376 (N_6376,N_5097,N_5671);
and U6377 (N_6377,N_5860,N_5765);
nor U6378 (N_6378,N_5696,N_5074);
xor U6379 (N_6379,N_5906,N_5772);
xnor U6380 (N_6380,N_5489,N_5186);
nand U6381 (N_6381,N_5493,N_5827);
and U6382 (N_6382,N_5929,N_5871);
and U6383 (N_6383,N_5717,N_5064);
nand U6384 (N_6384,N_5901,N_5244);
nor U6385 (N_6385,N_5026,N_5070);
nand U6386 (N_6386,N_5839,N_5875);
and U6387 (N_6387,N_5654,N_5864);
xor U6388 (N_6388,N_5956,N_5350);
nand U6389 (N_6389,N_5738,N_5159);
nand U6390 (N_6390,N_5933,N_5288);
and U6391 (N_6391,N_5795,N_5110);
xor U6392 (N_6392,N_5770,N_5635);
nor U6393 (N_6393,N_5931,N_5560);
nor U6394 (N_6394,N_5039,N_5981);
and U6395 (N_6395,N_5655,N_5245);
nor U6396 (N_6396,N_5968,N_5261);
xnor U6397 (N_6397,N_5255,N_5308);
nor U6398 (N_6398,N_5429,N_5553);
nor U6399 (N_6399,N_5700,N_5797);
and U6400 (N_6400,N_5484,N_5265);
nor U6401 (N_6401,N_5831,N_5992);
and U6402 (N_6402,N_5837,N_5843);
and U6403 (N_6403,N_5190,N_5060);
xnor U6404 (N_6404,N_5442,N_5233);
nor U6405 (N_6405,N_5590,N_5260);
nand U6406 (N_6406,N_5003,N_5847);
nand U6407 (N_6407,N_5591,N_5152);
nor U6408 (N_6408,N_5179,N_5507);
or U6409 (N_6409,N_5652,N_5882);
nand U6410 (N_6410,N_5082,N_5563);
nor U6411 (N_6411,N_5568,N_5703);
nand U6412 (N_6412,N_5050,N_5107);
or U6413 (N_6413,N_5394,N_5793);
nor U6414 (N_6414,N_5269,N_5556);
and U6415 (N_6415,N_5672,N_5558);
or U6416 (N_6416,N_5354,N_5144);
xnor U6417 (N_6417,N_5641,N_5554);
and U6418 (N_6418,N_5224,N_5856);
xor U6419 (N_6419,N_5247,N_5479);
xnor U6420 (N_6420,N_5117,N_5650);
or U6421 (N_6421,N_5701,N_5342);
nand U6422 (N_6422,N_5329,N_5150);
or U6423 (N_6423,N_5038,N_5090);
or U6424 (N_6424,N_5056,N_5577);
or U6425 (N_6425,N_5419,N_5603);
and U6426 (N_6426,N_5712,N_5470);
xnor U6427 (N_6427,N_5007,N_5677);
or U6428 (N_6428,N_5840,N_5092);
and U6429 (N_6429,N_5787,N_5191);
nor U6430 (N_6430,N_5093,N_5461);
xor U6431 (N_6431,N_5615,N_5528);
xnor U6432 (N_6432,N_5285,N_5043);
nor U6433 (N_6433,N_5031,N_5432);
nand U6434 (N_6434,N_5753,N_5228);
nand U6435 (N_6435,N_5184,N_5606);
xor U6436 (N_6436,N_5274,N_5236);
xnor U6437 (N_6437,N_5999,N_5973);
xor U6438 (N_6438,N_5927,N_5392);
and U6439 (N_6439,N_5527,N_5611);
nor U6440 (N_6440,N_5414,N_5526);
or U6441 (N_6441,N_5684,N_5719);
xor U6442 (N_6442,N_5722,N_5821);
xor U6443 (N_6443,N_5401,N_5706);
xor U6444 (N_6444,N_5971,N_5575);
or U6445 (N_6445,N_5919,N_5570);
xnor U6446 (N_6446,N_5273,N_5922);
nor U6447 (N_6447,N_5084,N_5616);
or U6448 (N_6448,N_5148,N_5124);
xor U6449 (N_6449,N_5227,N_5460);
xor U6450 (N_6450,N_5011,N_5299);
nand U6451 (N_6451,N_5705,N_5085);
nand U6452 (N_6452,N_5446,N_5114);
xnor U6453 (N_6453,N_5323,N_5366);
nand U6454 (N_6454,N_5204,N_5451);
xnor U6455 (N_6455,N_5237,N_5665);
nor U6456 (N_6456,N_5894,N_5531);
xnor U6457 (N_6457,N_5562,N_5036);
xnor U6458 (N_6458,N_5282,N_5598);
xnor U6459 (N_6459,N_5055,N_5022);
xnor U6460 (N_6460,N_5426,N_5353);
and U6461 (N_6461,N_5423,N_5012);
nand U6462 (N_6462,N_5564,N_5367);
nor U6463 (N_6463,N_5907,N_5278);
nand U6464 (N_6464,N_5535,N_5524);
and U6465 (N_6465,N_5849,N_5248);
and U6466 (N_6466,N_5805,N_5891);
and U6467 (N_6467,N_5226,N_5385);
xor U6468 (N_6468,N_5257,N_5183);
and U6469 (N_6469,N_5441,N_5475);
or U6470 (N_6470,N_5309,N_5456);
xor U6471 (N_6471,N_5579,N_5946);
nand U6472 (N_6472,N_5200,N_5578);
nor U6473 (N_6473,N_5964,N_5337);
or U6474 (N_6474,N_5359,N_5592);
nand U6475 (N_6475,N_5195,N_5375);
or U6476 (N_6476,N_5695,N_5935);
and U6477 (N_6477,N_5211,N_5250);
or U6478 (N_6478,N_5096,N_5667);
nand U6479 (N_6479,N_5958,N_5016);
xor U6480 (N_6480,N_5739,N_5634);
nor U6481 (N_6481,N_5567,N_5175);
xnor U6482 (N_6482,N_5778,N_5100);
xor U6483 (N_6483,N_5127,N_5517);
and U6484 (N_6484,N_5552,N_5510);
xor U6485 (N_6485,N_5569,N_5277);
and U6486 (N_6486,N_5963,N_5481);
nand U6487 (N_6487,N_5009,N_5286);
xnor U6488 (N_6488,N_5896,N_5325);
or U6489 (N_6489,N_5417,N_5081);
nor U6490 (N_6490,N_5065,N_5177);
or U6491 (N_6491,N_5911,N_5386);
xor U6492 (N_6492,N_5791,N_5443);
or U6493 (N_6493,N_5565,N_5612);
and U6494 (N_6494,N_5880,N_5504);
nand U6495 (N_6495,N_5953,N_5509);
nand U6496 (N_6496,N_5040,N_5134);
nand U6497 (N_6497,N_5996,N_5316);
nand U6498 (N_6498,N_5268,N_5952);
or U6499 (N_6499,N_5830,N_5997);
or U6500 (N_6500,N_5017,N_5042);
nand U6501 (N_6501,N_5631,N_5492);
nor U6502 (N_6502,N_5045,N_5020);
or U6503 (N_6503,N_5960,N_5354);
nand U6504 (N_6504,N_5485,N_5577);
and U6505 (N_6505,N_5531,N_5549);
nor U6506 (N_6506,N_5427,N_5097);
or U6507 (N_6507,N_5190,N_5088);
and U6508 (N_6508,N_5915,N_5291);
and U6509 (N_6509,N_5977,N_5795);
xnor U6510 (N_6510,N_5873,N_5171);
nand U6511 (N_6511,N_5381,N_5990);
and U6512 (N_6512,N_5835,N_5418);
nand U6513 (N_6513,N_5172,N_5662);
xor U6514 (N_6514,N_5300,N_5541);
nand U6515 (N_6515,N_5277,N_5870);
and U6516 (N_6516,N_5239,N_5002);
and U6517 (N_6517,N_5330,N_5943);
or U6518 (N_6518,N_5180,N_5700);
and U6519 (N_6519,N_5005,N_5255);
or U6520 (N_6520,N_5581,N_5092);
xnor U6521 (N_6521,N_5198,N_5406);
nor U6522 (N_6522,N_5999,N_5694);
xor U6523 (N_6523,N_5774,N_5776);
and U6524 (N_6524,N_5723,N_5644);
xor U6525 (N_6525,N_5612,N_5621);
and U6526 (N_6526,N_5695,N_5353);
and U6527 (N_6527,N_5403,N_5698);
and U6528 (N_6528,N_5331,N_5843);
and U6529 (N_6529,N_5553,N_5819);
or U6530 (N_6530,N_5405,N_5005);
nor U6531 (N_6531,N_5381,N_5056);
nand U6532 (N_6532,N_5494,N_5257);
and U6533 (N_6533,N_5521,N_5132);
nor U6534 (N_6534,N_5105,N_5829);
nor U6535 (N_6535,N_5876,N_5911);
or U6536 (N_6536,N_5744,N_5401);
nor U6537 (N_6537,N_5582,N_5082);
xor U6538 (N_6538,N_5408,N_5551);
xor U6539 (N_6539,N_5218,N_5383);
nor U6540 (N_6540,N_5312,N_5148);
xnor U6541 (N_6541,N_5408,N_5292);
nand U6542 (N_6542,N_5327,N_5429);
or U6543 (N_6543,N_5720,N_5586);
nand U6544 (N_6544,N_5641,N_5617);
or U6545 (N_6545,N_5671,N_5288);
nand U6546 (N_6546,N_5895,N_5878);
xor U6547 (N_6547,N_5924,N_5393);
and U6548 (N_6548,N_5631,N_5837);
and U6549 (N_6549,N_5744,N_5570);
and U6550 (N_6550,N_5688,N_5893);
xor U6551 (N_6551,N_5959,N_5673);
or U6552 (N_6552,N_5494,N_5421);
nor U6553 (N_6553,N_5321,N_5143);
and U6554 (N_6554,N_5132,N_5544);
nor U6555 (N_6555,N_5518,N_5371);
or U6556 (N_6556,N_5575,N_5449);
nand U6557 (N_6557,N_5397,N_5265);
and U6558 (N_6558,N_5935,N_5350);
and U6559 (N_6559,N_5308,N_5873);
xnor U6560 (N_6560,N_5961,N_5537);
and U6561 (N_6561,N_5491,N_5716);
xnor U6562 (N_6562,N_5332,N_5472);
nor U6563 (N_6563,N_5044,N_5105);
and U6564 (N_6564,N_5631,N_5003);
nand U6565 (N_6565,N_5966,N_5967);
xor U6566 (N_6566,N_5360,N_5959);
nand U6567 (N_6567,N_5452,N_5729);
or U6568 (N_6568,N_5851,N_5237);
or U6569 (N_6569,N_5452,N_5450);
xnor U6570 (N_6570,N_5233,N_5764);
nand U6571 (N_6571,N_5371,N_5310);
nand U6572 (N_6572,N_5679,N_5580);
or U6573 (N_6573,N_5871,N_5440);
nand U6574 (N_6574,N_5604,N_5023);
nand U6575 (N_6575,N_5559,N_5122);
xor U6576 (N_6576,N_5944,N_5341);
xor U6577 (N_6577,N_5416,N_5418);
or U6578 (N_6578,N_5043,N_5538);
xor U6579 (N_6579,N_5124,N_5686);
nor U6580 (N_6580,N_5889,N_5701);
or U6581 (N_6581,N_5368,N_5257);
nand U6582 (N_6582,N_5128,N_5280);
nor U6583 (N_6583,N_5754,N_5435);
nor U6584 (N_6584,N_5670,N_5289);
nor U6585 (N_6585,N_5725,N_5201);
xor U6586 (N_6586,N_5179,N_5338);
or U6587 (N_6587,N_5563,N_5077);
nand U6588 (N_6588,N_5338,N_5540);
nand U6589 (N_6589,N_5321,N_5525);
xor U6590 (N_6590,N_5346,N_5739);
nand U6591 (N_6591,N_5409,N_5617);
nor U6592 (N_6592,N_5374,N_5208);
or U6593 (N_6593,N_5836,N_5221);
or U6594 (N_6594,N_5502,N_5474);
or U6595 (N_6595,N_5229,N_5907);
or U6596 (N_6596,N_5572,N_5667);
nand U6597 (N_6597,N_5193,N_5683);
nand U6598 (N_6598,N_5971,N_5975);
nand U6599 (N_6599,N_5210,N_5091);
and U6600 (N_6600,N_5456,N_5672);
or U6601 (N_6601,N_5560,N_5637);
nand U6602 (N_6602,N_5399,N_5043);
and U6603 (N_6603,N_5656,N_5500);
or U6604 (N_6604,N_5628,N_5530);
nor U6605 (N_6605,N_5826,N_5610);
xor U6606 (N_6606,N_5165,N_5097);
xnor U6607 (N_6607,N_5577,N_5429);
or U6608 (N_6608,N_5319,N_5155);
xnor U6609 (N_6609,N_5925,N_5080);
or U6610 (N_6610,N_5310,N_5219);
or U6611 (N_6611,N_5788,N_5379);
or U6612 (N_6612,N_5301,N_5079);
xnor U6613 (N_6613,N_5897,N_5549);
or U6614 (N_6614,N_5329,N_5539);
xor U6615 (N_6615,N_5834,N_5277);
or U6616 (N_6616,N_5069,N_5421);
or U6617 (N_6617,N_5992,N_5630);
or U6618 (N_6618,N_5676,N_5296);
nand U6619 (N_6619,N_5552,N_5010);
or U6620 (N_6620,N_5630,N_5757);
xnor U6621 (N_6621,N_5274,N_5983);
nor U6622 (N_6622,N_5782,N_5516);
and U6623 (N_6623,N_5392,N_5366);
xnor U6624 (N_6624,N_5217,N_5820);
nand U6625 (N_6625,N_5716,N_5837);
nand U6626 (N_6626,N_5279,N_5192);
and U6627 (N_6627,N_5760,N_5227);
xor U6628 (N_6628,N_5863,N_5498);
and U6629 (N_6629,N_5884,N_5289);
nand U6630 (N_6630,N_5507,N_5643);
and U6631 (N_6631,N_5481,N_5578);
or U6632 (N_6632,N_5018,N_5557);
nand U6633 (N_6633,N_5741,N_5727);
and U6634 (N_6634,N_5838,N_5340);
or U6635 (N_6635,N_5137,N_5850);
xor U6636 (N_6636,N_5415,N_5980);
and U6637 (N_6637,N_5597,N_5222);
nand U6638 (N_6638,N_5834,N_5795);
nor U6639 (N_6639,N_5601,N_5343);
or U6640 (N_6640,N_5193,N_5194);
nor U6641 (N_6641,N_5383,N_5673);
nor U6642 (N_6642,N_5934,N_5817);
or U6643 (N_6643,N_5709,N_5689);
nor U6644 (N_6644,N_5469,N_5934);
or U6645 (N_6645,N_5327,N_5739);
nand U6646 (N_6646,N_5092,N_5249);
nor U6647 (N_6647,N_5829,N_5045);
or U6648 (N_6648,N_5384,N_5939);
xnor U6649 (N_6649,N_5193,N_5083);
and U6650 (N_6650,N_5355,N_5423);
and U6651 (N_6651,N_5360,N_5965);
and U6652 (N_6652,N_5660,N_5506);
xnor U6653 (N_6653,N_5430,N_5121);
nand U6654 (N_6654,N_5314,N_5796);
and U6655 (N_6655,N_5582,N_5235);
nor U6656 (N_6656,N_5218,N_5591);
nor U6657 (N_6657,N_5140,N_5447);
and U6658 (N_6658,N_5484,N_5422);
and U6659 (N_6659,N_5528,N_5963);
or U6660 (N_6660,N_5697,N_5244);
xor U6661 (N_6661,N_5364,N_5412);
nor U6662 (N_6662,N_5256,N_5277);
xnor U6663 (N_6663,N_5149,N_5860);
xor U6664 (N_6664,N_5518,N_5880);
or U6665 (N_6665,N_5156,N_5738);
nand U6666 (N_6666,N_5669,N_5255);
and U6667 (N_6667,N_5100,N_5568);
nor U6668 (N_6668,N_5169,N_5473);
and U6669 (N_6669,N_5519,N_5030);
nor U6670 (N_6670,N_5185,N_5717);
nand U6671 (N_6671,N_5064,N_5189);
xnor U6672 (N_6672,N_5226,N_5296);
nand U6673 (N_6673,N_5980,N_5165);
nor U6674 (N_6674,N_5512,N_5730);
or U6675 (N_6675,N_5240,N_5776);
and U6676 (N_6676,N_5796,N_5042);
or U6677 (N_6677,N_5725,N_5727);
nor U6678 (N_6678,N_5084,N_5351);
and U6679 (N_6679,N_5869,N_5946);
nand U6680 (N_6680,N_5212,N_5528);
or U6681 (N_6681,N_5270,N_5138);
nand U6682 (N_6682,N_5313,N_5155);
nor U6683 (N_6683,N_5688,N_5064);
and U6684 (N_6684,N_5187,N_5097);
nor U6685 (N_6685,N_5871,N_5591);
nand U6686 (N_6686,N_5082,N_5360);
or U6687 (N_6687,N_5491,N_5287);
nor U6688 (N_6688,N_5253,N_5355);
nor U6689 (N_6689,N_5154,N_5837);
nor U6690 (N_6690,N_5487,N_5694);
xor U6691 (N_6691,N_5191,N_5348);
and U6692 (N_6692,N_5476,N_5527);
nand U6693 (N_6693,N_5686,N_5685);
or U6694 (N_6694,N_5088,N_5019);
and U6695 (N_6695,N_5312,N_5977);
and U6696 (N_6696,N_5596,N_5105);
nand U6697 (N_6697,N_5072,N_5480);
or U6698 (N_6698,N_5688,N_5236);
nor U6699 (N_6699,N_5039,N_5422);
nor U6700 (N_6700,N_5022,N_5794);
nor U6701 (N_6701,N_5194,N_5451);
xor U6702 (N_6702,N_5269,N_5628);
xnor U6703 (N_6703,N_5110,N_5302);
and U6704 (N_6704,N_5225,N_5315);
nand U6705 (N_6705,N_5339,N_5051);
and U6706 (N_6706,N_5901,N_5889);
xnor U6707 (N_6707,N_5178,N_5616);
or U6708 (N_6708,N_5210,N_5012);
nand U6709 (N_6709,N_5094,N_5370);
xnor U6710 (N_6710,N_5563,N_5967);
or U6711 (N_6711,N_5005,N_5726);
and U6712 (N_6712,N_5828,N_5867);
nor U6713 (N_6713,N_5326,N_5031);
or U6714 (N_6714,N_5730,N_5715);
xor U6715 (N_6715,N_5371,N_5354);
or U6716 (N_6716,N_5536,N_5201);
and U6717 (N_6717,N_5600,N_5104);
nand U6718 (N_6718,N_5483,N_5637);
nor U6719 (N_6719,N_5501,N_5021);
and U6720 (N_6720,N_5724,N_5397);
or U6721 (N_6721,N_5576,N_5474);
xor U6722 (N_6722,N_5875,N_5791);
nand U6723 (N_6723,N_5312,N_5770);
nor U6724 (N_6724,N_5817,N_5973);
and U6725 (N_6725,N_5912,N_5295);
and U6726 (N_6726,N_5390,N_5196);
nand U6727 (N_6727,N_5858,N_5961);
or U6728 (N_6728,N_5206,N_5516);
and U6729 (N_6729,N_5936,N_5873);
nand U6730 (N_6730,N_5431,N_5873);
xor U6731 (N_6731,N_5327,N_5470);
nand U6732 (N_6732,N_5038,N_5344);
xor U6733 (N_6733,N_5054,N_5079);
xnor U6734 (N_6734,N_5463,N_5810);
nor U6735 (N_6735,N_5425,N_5500);
or U6736 (N_6736,N_5614,N_5817);
nand U6737 (N_6737,N_5529,N_5090);
nand U6738 (N_6738,N_5582,N_5483);
nor U6739 (N_6739,N_5223,N_5213);
xor U6740 (N_6740,N_5968,N_5849);
and U6741 (N_6741,N_5031,N_5668);
xor U6742 (N_6742,N_5450,N_5011);
xor U6743 (N_6743,N_5804,N_5722);
xor U6744 (N_6744,N_5713,N_5577);
and U6745 (N_6745,N_5490,N_5729);
nand U6746 (N_6746,N_5693,N_5894);
and U6747 (N_6747,N_5522,N_5215);
and U6748 (N_6748,N_5096,N_5378);
nor U6749 (N_6749,N_5018,N_5370);
and U6750 (N_6750,N_5598,N_5680);
nor U6751 (N_6751,N_5770,N_5024);
xnor U6752 (N_6752,N_5830,N_5909);
and U6753 (N_6753,N_5969,N_5672);
nand U6754 (N_6754,N_5182,N_5625);
xnor U6755 (N_6755,N_5040,N_5277);
nor U6756 (N_6756,N_5511,N_5807);
or U6757 (N_6757,N_5741,N_5127);
xor U6758 (N_6758,N_5775,N_5210);
xor U6759 (N_6759,N_5703,N_5203);
nor U6760 (N_6760,N_5056,N_5800);
xor U6761 (N_6761,N_5430,N_5378);
or U6762 (N_6762,N_5798,N_5965);
nor U6763 (N_6763,N_5700,N_5625);
xnor U6764 (N_6764,N_5399,N_5766);
and U6765 (N_6765,N_5463,N_5836);
nor U6766 (N_6766,N_5185,N_5315);
nor U6767 (N_6767,N_5273,N_5786);
nor U6768 (N_6768,N_5953,N_5142);
and U6769 (N_6769,N_5830,N_5829);
xnor U6770 (N_6770,N_5682,N_5136);
and U6771 (N_6771,N_5844,N_5716);
nand U6772 (N_6772,N_5221,N_5649);
nor U6773 (N_6773,N_5850,N_5297);
nand U6774 (N_6774,N_5799,N_5578);
or U6775 (N_6775,N_5346,N_5555);
nor U6776 (N_6776,N_5169,N_5384);
or U6777 (N_6777,N_5950,N_5421);
or U6778 (N_6778,N_5290,N_5535);
or U6779 (N_6779,N_5891,N_5346);
or U6780 (N_6780,N_5027,N_5407);
xor U6781 (N_6781,N_5957,N_5306);
xnor U6782 (N_6782,N_5511,N_5169);
and U6783 (N_6783,N_5400,N_5232);
or U6784 (N_6784,N_5602,N_5274);
nor U6785 (N_6785,N_5120,N_5808);
or U6786 (N_6786,N_5619,N_5053);
xnor U6787 (N_6787,N_5836,N_5250);
or U6788 (N_6788,N_5895,N_5091);
nand U6789 (N_6789,N_5804,N_5545);
nand U6790 (N_6790,N_5406,N_5029);
and U6791 (N_6791,N_5373,N_5558);
xnor U6792 (N_6792,N_5256,N_5824);
nand U6793 (N_6793,N_5684,N_5355);
or U6794 (N_6794,N_5241,N_5619);
nand U6795 (N_6795,N_5080,N_5403);
nand U6796 (N_6796,N_5257,N_5598);
or U6797 (N_6797,N_5710,N_5518);
xor U6798 (N_6798,N_5876,N_5968);
nor U6799 (N_6799,N_5070,N_5778);
xnor U6800 (N_6800,N_5542,N_5964);
nor U6801 (N_6801,N_5369,N_5143);
nor U6802 (N_6802,N_5001,N_5251);
nand U6803 (N_6803,N_5651,N_5172);
nor U6804 (N_6804,N_5342,N_5504);
nor U6805 (N_6805,N_5921,N_5096);
or U6806 (N_6806,N_5670,N_5526);
or U6807 (N_6807,N_5147,N_5016);
nand U6808 (N_6808,N_5755,N_5497);
and U6809 (N_6809,N_5047,N_5817);
nor U6810 (N_6810,N_5290,N_5705);
xnor U6811 (N_6811,N_5967,N_5425);
nor U6812 (N_6812,N_5810,N_5900);
nand U6813 (N_6813,N_5245,N_5602);
or U6814 (N_6814,N_5295,N_5206);
nor U6815 (N_6815,N_5160,N_5011);
xor U6816 (N_6816,N_5462,N_5163);
nor U6817 (N_6817,N_5104,N_5012);
or U6818 (N_6818,N_5785,N_5697);
nor U6819 (N_6819,N_5572,N_5442);
nor U6820 (N_6820,N_5292,N_5853);
nor U6821 (N_6821,N_5710,N_5558);
nor U6822 (N_6822,N_5573,N_5793);
or U6823 (N_6823,N_5356,N_5556);
xnor U6824 (N_6824,N_5335,N_5574);
and U6825 (N_6825,N_5748,N_5451);
xnor U6826 (N_6826,N_5837,N_5289);
and U6827 (N_6827,N_5626,N_5603);
nand U6828 (N_6828,N_5621,N_5427);
nor U6829 (N_6829,N_5848,N_5104);
and U6830 (N_6830,N_5617,N_5381);
nor U6831 (N_6831,N_5656,N_5649);
xnor U6832 (N_6832,N_5769,N_5224);
nand U6833 (N_6833,N_5931,N_5874);
and U6834 (N_6834,N_5180,N_5976);
xor U6835 (N_6835,N_5735,N_5618);
or U6836 (N_6836,N_5544,N_5892);
and U6837 (N_6837,N_5799,N_5310);
xor U6838 (N_6838,N_5142,N_5709);
xnor U6839 (N_6839,N_5990,N_5517);
or U6840 (N_6840,N_5631,N_5817);
and U6841 (N_6841,N_5110,N_5867);
and U6842 (N_6842,N_5326,N_5367);
nor U6843 (N_6843,N_5714,N_5001);
and U6844 (N_6844,N_5657,N_5573);
or U6845 (N_6845,N_5891,N_5916);
nor U6846 (N_6846,N_5134,N_5971);
nand U6847 (N_6847,N_5833,N_5178);
and U6848 (N_6848,N_5123,N_5350);
or U6849 (N_6849,N_5038,N_5258);
xnor U6850 (N_6850,N_5690,N_5253);
nand U6851 (N_6851,N_5743,N_5863);
or U6852 (N_6852,N_5100,N_5384);
and U6853 (N_6853,N_5435,N_5020);
nand U6854 (N_6854,N_5394,N_5611);
or U6855 (N_6855,N_5102,N_5216);
nand U6856 (N_6856,N_5302,N_5469);
nand U6857 (N_6857,N_5280,N_5331);
or U6858 (N_6858,N_5048,N_5203);
and U6859 (N_6859,N_5821,N_5923);
and U6860 (N_6860,N_5456,N_5618);
xnor U6861 (N_6861,N_5833,N_5383);
xor U6862 (N_6862,N_5027,N_5750);
xnor U6863 (N_6863,N_5379,N_5389);
xnor U6864 (N_6864,N_5528,N_5884);
xnor U6865 (N_6865,N_5243,N_5935);
nor U6866 (N_6866,N_5738,N_5579);
nand U6867 (N_6867,N_5195,N_5509);
xor U6868 (N_6868,N_5798,N_5703);
nand U6869 (N_6869,N_5737,N_5221);
nor U6870 (N_6870,N_5940,N_5921);
and U6871 (N_6871,N_5063,N_5390);
or U6872 (N_6872,N_5406,N_5037);
or U6873 (N_6873,N_5517,N_5266);
nor U6874 (N_6874,N_5389,N_5711);
nand U6875 (N_6875,N_5878,N_5935);
and U6876 (N_6876,N_5593,N_5685);
or U6877 (N_6877,N_5521,N_5397);
nand U6878 (N_6878,N_5840,N_5344);
xnor U6879 (N_6879,N_5375,N_5334);
and U6880 (N_6880,N_5992,N_5394);
or U6881 (N_6881,N_5931,N_5451);
or U6882 (N_6882,N_5252,N_5775);
xnor U6883 (N_6883,N_5652,N_5813);
or U6884 (N_6884,N_5210,N_5303);
xor U6885 (N_6885,N_5094,N_5313);
and U6886 (N_6886,N_5370,N_5750);
xor U6887 (N_6887,N_5687,N_5945);
and U6888 (N_6888,N_5896,N_5195);
and U6889 (N_6889,N_5547,N_5055);
xnor U6890 (N_6890,N_5479,N_5926);
nor U6891 (N_6891,N_5389,N_5497);
nor U6892 (N_6892,N_5651,N_5729);
xnor U6893 (N_6893,N_5884,N_5545);
nand U6894 (N_6894,N_5937,N_5597);
xnor U6895 (N_6895,N_5340,N_5278);
or U6896 (N_6896,N_5974,N_5682);
xnor U6897 (N_6897,N_5264,N_5981);
or U6898 (N_6898,N_5000,N_5489);
xor U6899 (N_6899,N_5422,N_5217);
nand U6900 (N_6900,N_5509,N_5153);
and U6901 (N_6901,N_5121,N_5199);
xnor U6902 (N_6902,N_5951,N_5793);
xor U6903 (N_6903,N_5703,N_5877);
xor U6904 (N_6904,N_5445,N_5516);
and U6905 (N_6905,N_5442,N_5507);
nand U6906 (N_6906,N_5459,N_5814);
and U6907 (N_6907,N_5987,N_5409);
or U6908 (N_6908,N_5463,N_5491);
and U6909 (N_6909,N_5077,N_5801);
or U6910 (N_6910,N_5415,N_5217);
xnor U6911 (N_6911,N_5960,N_5368);
xor U6912 (N_6912,N_5809,N_5642);
and U6913 (N_6913,N_5003,N_5428);
xor U6914 (N_6914,N_5247,N_5230);
nor U6915 (N_6915,N_5794,N_5081);
xnor U6916 (N_6916,N_5969,N_5923);
xor U6917 (N_6917,N_5384,N_5246);
nand U6918 (N_6918,N_5520,N_5366);
nand U6919 (N_6919,N_5155,N_5844);
xor U6920 (N_6920,N_5198,N_5303);
nor U6921 (N_6921,N_5468,N_5587);
and U6922 (N_6922,N_5131,N_5865);
nand U6923 (N_6923,N_5554,N_5210);
nand U6924 (N_6924,N_5634,N_5424);
nor U6925 (N_6925,N_5774,N_5937);
nand U6926 (N_6926,N_5341,N_5941);
and U6927 (N_6927,N_5631,N_5958);
and U6928 (N_6928,N_5924,N_5036);
or U6929 (N_6929,N_5267,N_5107);
and U6930 (N_6930,N_5987,N_5323);
xnor U6931 (N_6931,N_5637,N_5854);
xor U6932 (N_6932,N_5283,N_5773);
and U6933 (N_6933,N_5358,N_5200);
nand U6934 (N_6934,N_5211,N_5433);
or U6935 (N_6935,N_5502,N_5045);
or U6936 (N_6936,N_5642,N_5036);
and U6937 (N_6937,N_5438,N_5848);
nand U6938 (N_6938,N_5695,N_5728);
and U6939 (N_6939,N_5605,N_5905);
and U6940 (N_6940,N_5838,N_5962);
nand U6941 (N_6941,N_5374,N_5528);
or U6942 (N_6942,N_5162,N_5173);
nor U6943 (N_6943,N_5127,N_5049);
nand U6944 (N_6944,N_5084,N_5875);
xnor U6945 (N_6945,N_5289,N_5172);
nand U6946 (N_6946,N_5255,N_5578);
nand U6947 (N_6947,N_5042,N_5018);
and U6948 (N_6948,N_5997,N_5508);
xnor U6949 (N_6949,N_5940,N_5526);
nand U6950 (N_6950,N_5133,N_5627);
and U6951 (N_6951,N_5474,N_5465);
nor U6952 (N_6952,N_5827,N_5914);
xor U6953 (N_6953,N_5918,N_5830);
nor U6954 (N_6954,N_5145,N_5032);
nand U6955 (N_6955,N_5094,N_5645);
nand U6956 (N_6956,N_5882,N_5530);
xnor U6957 (N_6957,N_5162,N_5287);
nand U6958 (N_6958,N_5312,N_5537);
xnor U6959 (N_6959,N_5402,N_5525);
nand U6960 (N_6960,N_5054,N_5783);
or U6961 (N_6961,N_5395,N_5161);
and U6962 (N_6962,N_5015,N_5484);
nor U6963 (N_6963,N_5268,N_5871);
nand U6964 (N_6964,N_5894,N_5895);
xnor U6965 (N_6965,N_5371,N_5304);
nor U6966 (N_6966,N_5756,N_5264);
nor U6967 (N_6967,N_5583,N_5579);
nand U6968 (N_6968,N_5451,N_5567);
nand U6969 (N_6969,N_5146,N_5759);
xnor U6970 (N_6970,N_5373,N_5772);
nand U6971 (N_6971,N_5252,N_5990);
xnor U6972 (N_6972,N_5535,N_5087);
and U6973 (N_6973,N_5298,N_5400);
or U6974 (N_6974,N_5835,N_5946);
xor U6975 (N_6975,N_5346,N_5055);
or U6976 (N_6976,N_5910,N_5877);
or U6977 (N_6977,N_5209,N_5763);
nor U6978 (N_6978,N_5955,N_5210);
and U6979 (N_6979,N_5974,N_5578);
nand U6980 (N_6980,N_5780,N_5855);
and U6981 (N_6981,N_5701,N_5508);
nand U6982 (N_6982,N_5594,N_5527);
and U6983 (N_6983,N_5762,N_5557);
nor U6984 (N_6984,N_5099,N_5365);
nand U6985 (N_6985,N_5199,N_5652);
nor U6986 (N_6986,N_5711,N_5414);
xnor U6987 (N_6987,N_5828,N_5777);
xnor U6988 (N_6988,N_5219,N_5761);
and U6989 (N_6989,N_5155,N_5935);
xor U6990 (N_6990,N_5319,N_5440);
nand U6991 (N_6991,N_5295,N_5790);
or U6992 (N_6992,N_5159,N_5322);
or U6993 (N_6993,N_5681,N_5210);
or U6994 (N_6994,N_5445,N_5232);
nor U6995 (N_6995,N_5533,N_5081);
nor U6996 (N_6996,N_5814,N_5710);
nand U6997 (N_6997,N_5819,N_5301);
nand U6998 (N_6998,N_5665,N_5612);
nand U6999 (N_6999,N_5840,N_5949);
nand U7000 (N_7000,N_6550,N_6421);
nor U7001 (N_7001,N_6457,N_6608);
and U7002 (N_7002,N_6861,N_6908);
nor U7003 (N_7003,N_6751,N_6972);
nand U7004 (N_7004,N_6577,N_6310);
and U7005 (N_7005,N_6785,N_6396);
xor U7006 (N_7006,N_6215,N_6145);
nand U7007 (N_7007,N_6249,N_6174);
or U7008 (N_7008,N_6453,N_6901);
nor U7009 (N_7009,N_6938,N_6078);
xnor U7010 (N_7010,N_6038,N_6849);
and U7011 (N_7011,N_6259,N_6842);
xor U7012 (N_7012,N_6882,N_6462);
and U7013 (N_7013,N_6322,N_6479);
nor U7014 (N_7014,N_6728,N_6300);
nor U7015 (N_7015,N_6353,N_6979);
nand U7016 (N_7016,N_6970,N_6508);
or U7017 (N_7017,N_6250,N_6359);
nand U7018 (N_7018,N_6127,N_6212);
nor U7019 (N_7019,N_6167,N_6092);
xnor U7020 (N_7020,N_6893,N_6292);
and U7021 (N_7021,N_6976,N_6990);
nor U7022 (N_7022,N_6819,N_6470);
nand U7023 (N_7023,N_6389,N_6746);
xor U7024 (N_7024,N_6811,N_6697);
and U7025 (N_7025,N_6758,N_6579);
xor U7026 (N_7026,N_6646,N_6190);
nand U7027 (N_7027,N_6948,N_6983);
nor U7028 (N_7028,N_6563,N_6253);
xnor U7029 (N_7029,N_6308,N_6841);
or U7030 (N_7030,N_6641,N_6772);
and U7031 (N_7031,N_6536,N_6111);
nor U7032 (N_7032,N_6110,N_6930);
nand U7033 (N_7033,N_6251,N_6007);
nor U7034 (N_7034,N_6714,N_6160);
nor U7035 (N_7035,N_6175,N_6583);
and U7036 (N_7036,N_6791,N_6923);
nand U7037 (N_7037,N_6906,N_6875);
nor U7038 (N_7038,N_6917,N_6414);
nand U7039 (N_7039,N_6822,N_6594);
xor U7040 (N_7040,N_6416,N_6890);
nand U7041 (N_7041,N_6054,N_6341);
xor U7042 (N_7042,N_6080,N_6449);
and U7043 (N_7043,N_6737,N_6124);
nand U7044 (N_7044,N_6812,N_6753);
xnor U7045 (N_7045,N_6866,N_6115);
nand U7046 (N_7046,N_6671,N_6522);
nand U7047 (N_7047,N_6411,N_6944);
nor U7048 (N_7048,N_6719,N_6884);
nand U7049 (N_7049,N_6996,N_6014);
xor U7050 (N_7050,N_6126,N_6180);
or U7051 (N_7051,N_6278,N_6987);
or U7052 (N_7052,N_6897,N_6108);
nand U7053 (N_7053,N_6535,N_6178);
nand U7054 (N_7054,N_6258,N_6327);
nand U7055 (N_7055,N_6339,N_6821);
xor U7056 (N_7056,N_6869,N_6472);
nand U7057 (N_7057,N_6723,N_6920);
or U7058 (N_7058,N_6418,N_6189);
and U7059 (N_7059,N_6325,N_6372);
and U7060 (N_7060,N_6843,N_6801);
and U7061 (N_7061,N_6552,N_6686);
and U7062 (N_7062,N_6514,N_6820);
and U7063 (N_7063,N_6147,N_6570);
xor U7064 (N_7064,N_6048,N_6314);
and U7065 (N_7065,N_6564,N_6815);
and U7066 (N_7066,N_6613,N_6391);
and U7067 (N_7067,N_6778,N_6307);
nand U7068 (N_7068,N_6735,N_6363);
or U7069 (N_7069,N_6012,N_6531);
nor U7070 (N_7070,N_6280,N_6086);
nand U7071 (N_7071,N_6155,N_6103);
nand U7072 (N_7072,N_6705,N_6524);
xor U7073 (N_7073,N_6210,N_6852);
and U7074 (N_7074,N_6900,N_6943);
xnor U7075 (N_7075,N_6360,N_6766);
or U7076 (N_7076,N_6988,N_6222);
xor U7077 (N_7077,N_6960,N_6779);
xnor U7078 (N_7078,N_6729,N_6836);
nand U7079 (N_7079,N_6196,N_6713);
nand U7080 (N_7080,N_6847,N_6000);
and U7081 (N_7081,N_6755,N_6503);
and U7082 (N_7082,N_6030,N_6914);
nand U7083 (N_7083,N_6351,N_6208);
nor U7084 (N_7084,N_6216,N_6932);
nand U7085 (N_7085,N_6084,N_6828);
and U7086 (N_7086,N_6956,N_6984);
and U7087 (N_7087,N_6247,N_6478);
nand U7088 (N_7088,N_6853,N_6358);
or U7089 (N_7089,N_6218,N_6643);
or U7090 (N_7090,N_6826,N_6015);
xor U7091 (N_7091,N_6087,N_6112);
nor U7092 (N_7092,N_6448,N_6120);
and U7093 (N_7093,N_6637,N_6443);
xor U7094 (N_7094,N_6879,N_6378);
nor U7095 (N_7095,N_6761,N_6371);
and U7096 (N_7096,N_6625,N_6241);
and U7097 (N_7097,N_6818,N_6343);
nor U7098 (N_7098,N_6333,N_6904);
xnor U7099 (N_7099,N_6556,N_6878);
xnor U7100 (N_7100,N_6295,N_6540);
nor U7101 (N_7101,N_6927,N_6061);
nor U7102 (N_7102,N_6966,N_6848);
and U7103 (N_7103,N_6373,N_6635);
nand U7104 (N_7104,N_6480,N_6829);
and U7105 (N_7105,N_6808,N_6370);
xnor U7106 (N_7106,N_6867,N_6139);
xnor U7107 (N_7107,N_6079,N_6040);
xnor U7108 (N_7108,N_6626,N_6864);
and U7109 (N_7109,N_6315,N_6582);
nor U7110 (N_7110,N_6043,N_6033);
xor U7111 (N_7111,N_6885,N_6907);
xnor U7112 (N_7112,N_6961,N_6316);
xnor U7113 (N_7113,N_6876,N_6188);
nand U7114 (N_7114,N_6129,N_6454);
nand U7115 (N_7115,N_6279,N_6365);
or U7116 (N_7116,N_6660,N_6607);
nor U7117 (N_7117,N_6498,N_6616);
and U7118 (N_7118,N_6787,N_6986);
or U7119 (N_7119,N_6862,N_6130);
or U7120 (N_7120,N_6539,N_6614);
xor U7121 (N_7121,N_6615,N_6011);
nand U7122 (N_7122,N_6688,N_6924);
nand U7123 (N_7123,N_6534,N_6994);
nor U7124 (N_7124,N_6777,N_6747);
or U7125 (N_7125,N_6732,N_6285);
nor U7126 (N_7126,N_6991,N_6311);
and U7127 (N_7127,N_6549,N_6042);
xor U7128 (N_7128,N_6571,N_6148);
or U7129 (N_7129,N_6973,N_6967);
and U7130 (N_7130,N_6255,N_6335);
nand U7131 (N_7131,N_6515,N_6659);
or U7132 (N_7132,N_6050,N_6759);
nor U7133 (N_7133,N_6022,N_6098);
and U7134 (N_7134,N_6368,N_6382);
xnor U7135 (N_7135,N_6918,N_6790);
and U7136 (N_7136,N_6262,N_6168);
or U7137 (N_7137,N_6827,N_6995);
or U7138 (N_7138,N_6588,N_6533);
nand U7139 (N_7139,N_6150,N_6611);
nor U7140 (N_7140,N_6407,N_6282);
xor U7141 (N_7141,N_6450,N_6902);
or U7142 (N_7142,N_6634,N_6297);
nor U7143 (N_7143,N_6628,N_6679);
nor U7144 (N_7144,N_6565,N_6546);
nor U7145 (N_7145,N_6799,N_6949);
nand U7146 (N_7146,N_6667,N_6794);
nand U7147 (N_7147,N_6451,N_6206);
or U7148 (N_7148,N_6695,N_6870);
nand U7149 (N_7149,N_6655,N_6248);
nand U7150 (N_7150,N_6348,N_6832);
xnor U7151 (N_7151,N_6313,N_6653);
and U7152 (N_7152,N_6813,N_6865);
nand U7153 (N_7153,N_6543,N_6463);
xnor U7154 (N_7154,N_6274,N_6136);
or U7155 (N_7155,N_6393,N_6326);
or U7156 (N_7156,N_6545,N_6730);
xnor U7157 (N_7157,N_6648,N_6041);
and U7158 (N_7158,N_6770,N_6107);
xor U7159 (N_7159,N_6946,N_6551);
nor U7160 (N_7160,N_6817,N_6639);
and U7161 (N_7161,N_6525,N_6026);
and U7162 (N_7162,N_6789,N_6569);
nor U7163 (N_7163,N_6101,N_6925);
nor U7164 (N_7164,N_6992,N_6225);
nor U7165 (N_7165,N_6195,N_6741);
xnor U7166 (N_7166,N_6203,N_6141);
or U7167 (N_7167,N_6010,N_6270);
xor U7168 (N_7168,N_6654,N_6433);
and U7169 (N_7169,N_6538,N_6937);
xnor U7170 (N_7170,N_6383,N_6873);
and U7171 (N_7171,N_6511,N_6459);
nor U7172 (N_7172,N_6572,N_6420);
xnor U7173 (N_7173,N_6555,N_6762);
xor U7174 (N_7174,N_6431,N_6413);
and U7175 (N_7175,N_6760,N_6649);
and U7176 (N_7176,N_6709,N_6803);
or U7177 (N_7177,N_6501,N_6122);
nor U7178 (N_7178,N_6739,N_6939);
or U7179 (N_7179,N_6224,N_6717);
or U7180 (N_7180,N_6055,N_6580);
and U7181 (N_7181,N_6361,N_6073);
and U7182 (N_7182,N_6858,N_6272);
and U7183 (N_7183,N_6690,N_6461);
nand U7184 (N_7184,N_6936,N_6436);
nor U7185 (N_7185,N_6722,N_6476);
nor U7186 (N_7186,N_6602,N_6680);
nand U7187 (N_7187,N_6483,N_6256);
and U7188 (N_7188,N_6125,N_6512);
and U7189 (N_7189,N_6229,N_6574);
nand U7190 (N_7190,N_6355,N_6330);
xnor U7191 (N_7191,N_6887,N_6140);
nor U7192 (N_7192,N_6075,N_6342);
nor U7193 (N_7193,N_6119,N_6689);
nor U7194 (N_7194,N_6469,N_6752);
and U7195 (N_7195,N_6622,N_6261);
nand U7196 (N_7196,N_6985,N_6035);
nor U7197 (N_7197,N_6640,N_6143);
nand U7198 (N_7198,N_6299,N_6673);
xor U7199 (N_7199,N_6656,N_6381);
or U7200 (N_7200,N_6591,N_6687);
xnor U7201 (N_7201,N_6404,N_6593);
nand U7202 (N_7202,N_6781,N_6977);
xor U7203 (N_7203,N_6644,N_6627);
and U7204 (N_7204,N_6909,N_6156);
nor U7205 (N_7205,N_6810,N_6899);
nor U7206 (N_7206,N_6502,N_6645);
nand U7207 (N_7207,N_6070,N_6675);
nand U7208 (N_7208,N_6052,N_6047);
and U7209 (N_7209,N_6039,N_6312);
or U7210 (N_7210,N_6484,N_6441);
and U7211 (N_7211,N_6495,N_6856);
and U7212 (N_7212,N_6223,N_6239);
or U7213 (N_7213,N_6494,N_6064);
xnor U7214 (N_7214,N_6284,N_6093);
nand U7215 (N_7215,N_6186,N_6517);
or U7216 (N_7216,N_6481,N_6390);
and U7217 (N_7217,N_6194,N_6444);
nor U7218 (N_7218,N_6409,N_6490);
nor U7219 (N_7219,N_6402,N_6037);
nand U7220 (N_7220,N_6756,N_6850);
xor U7221 (N_7221,N_6488,N_6809);
or U7222 (N_7222,N_6768,N_6321);
nor U7223 (N_7223,N_6513,N_6013);
xnor U7224 (N_7224,N_6291,N_6521);
and U7225 (N_7225,N_6354,N_6375);
and U7226 (N_7226,N_6710,N_6068);
and U7227 (N_7227,N_6271,N_6796);
xnor U7228 (N_7228,N_6706,N_6116);
xor U7229 (N_7229,N_6780,N_6123);
or U7230 (N_7230,N_6769,N_6336);
xnor U7231 (N_7231,N_6135,N_6231);
or U7232 (N_7232,N_6001,N_6090);
nand U7233 (N_7233,N_6429,N_6164);
xnor U7234 (N_7234,N_6304,N_6587);
xnor U7235 (N_7235,N_6426,N_6004);
and U7236 (N_7236,N_6590,N_6027);
or U7237 (N_7237,N_6497,N_6095);
and U7238 (N_7238,N_6559,N_6993);
nor U7239 (N_7239,N_6105,N_6149);
or U7240 (N_7240,N_6317,N_6072);
nand U7241 (N_7241,N_6185,N_6699);
and U7242 (N_7242,N_6097,N_6388);
nor U7243 (N_7243,N_6672,N_6214);
nand U7244 (N_7244,N_6405,N_6474);
nand U7245 (N_7245,N_6731,N_6652);
nor U7246 (N_7246,N_6704,N_6056);
or U7247 (N_7247,N_6855,N_6267);
xor U7248 (N_7248,N_6106,N_6176);
nor U7249 (N_7249,N_6684,N_6945);
xor U7250 (N_7250,N_6379,N_6963);
or U7251 (N_7251,N_6621,N_6319);
nand U7252 (N_7252,N_6083,N_6493);
xnor U7253 (N_7253,N_6209,N_6465);
and U7254 (N_7254,N_6573,N_6169);
xnor U7255 (N_7255,N_6179,N_6076);
nor U7256 (N_7256,N_6506,N_6800);
xor U7257 (N_7257,N_6532,N_6666);
or U7258 (N_7258,N_6471,N_6837);
xnor U7259 (N_7259,N_6584,N_6578);
and U7260 (N_7260,N_6171,N_6200);
and U7261 (N_7261,N_6332,N_6109);
xnor U7262 (N_7262,N_6548,N_6219);
and U7263 (N_7263,N_6252,N_6889);
or U7264 (N_7264,N_6269,N_6903);
xor U7265 (N_7265,N_6942,N_6099);
and U7266 (N_7266,N_6157,N_6034);
xnor U7267 (N_7267,N_6374,N_6142);
xnor U7268 (N_7268,N_6959,N_6346);
and U7269 (N_7269,N_6558,N_6566);
xnor U7270 (N_7270,N_6238,N_6046);
or U7271 (N_7271,N_6446,N_6286);
xnor U7272 (N_7272,N_6430,N_6951);
nor U7273 (N_7273,N_6630,N_6337);
xnor U7274 (N_7274,N_6133,N_6211);
xor U7275 (N_7275,N_6019,N_6757);
xor U7276 (N_7276,N_6387,N_6468);
nor U7277 (N_7277,N_6165,N_6662);
or U7278 (N_7278,N_6151,N_6260);
nor U7279 (N_7279,N_6344,N_6568);
nand U7280 (N_7280,N_6542,N_6537);
xor U7281 (N_7281,N_6916,N_6331);
or U7282 (N_7282,N_6999,N_6170);
nand U7283 (N_7283,N_6971,N_6857);
nor U7284 (N_7284,N_6257,N_6029);
and U7285 (N_7285,N_6246,N_6096);
xor U7286 (N_7286,N_6919,N_6377);
xor U7287 (N_7287,N_6892,N_6561);
nor U7288 (N_7288,N_6094,N_6400);
or U7289 (N_7289,N_6036,N_6415);
xor U7290 (N_7290,N_6477,N_6466);
nor U7291 (N_7291,N_6896,N_6357);
or U7292 (N_7292,N_6191,N_6144);
or U7293 (N_7293,N_6700,N_6989);
nor U7294 (N_7294,N_6242,N_6386);
nor U7295 (N_7295,N_6871,N_6456);
nor U7296 (N_7296,N_6166,N_6698);
nand U7297 (N_7297,N_6118,N_6277);
nor U7298 (N_7298,N_6432,N_6349);
or U7299 (N_7299,N_6872,N_6067);
xnor U7300 (N_7300,N_6236,N_6044);
nand U7301 (N_7301,N_6807,N_6428);
and U7302 (N_7302,N_6589,N_6338);
xnor U7303 (N_7303,N_6773,N_6736);
nor U7304 (N_7304,N_6499,N_6162);
nor U7305 (N_7305,N_6121,N_6057);
nor U7306 (N_7306,N_6302,N_6283);
nor U7307 (N_7307,N_6604,N_6199);
xnor U7308 (N_7308,N_6399,N_6205);
xor U7309 (N_7309,N_6289,N_6691);
nor U7310 (N_7310,N_6005,N_6510);
nor U7311 (N_7311,N_6926,N_6347);
and U7312 (N_7312,N_6173,N_6676);
or U7313 (N_7313,N_6213,N_6629);
nor U7314 (N_7314,N_6711,N_6771);
xnor U7315 (N_7315,N_6567,N_6738);
nand U7316 (N_7316,N_6177,N_6955);
or U7317 (N_7317,N_6293,N_6838);
or U7318 (N_7318,N_6233,N_6599);
and U7319 (N_7319,N_6806,N_6703);
nand U7320 (N_7320,N_6782,N_6235);
nor U7321 (N_7321,N_6006,N_6650);
nor U7322 (N_7322,N_6306,N_6886);
nand U7323 (N_7323,N_6802,N_6245);
and U7324 (N_7324,N_6929,N_6586);
nor U7325 (N_7325,N_6793,N_6702);
xor U7326 (N_7326,N_6217,N_6795);
nand U7327 (N_7327,N_6172,N_6744);
nand U7328 (N_7328,N_6424,N_6071);
xnor U7329 (N_7329,N_6788,N_6184);
and U7330 (N_7330,N_6309,N_6017);
or U7331 (N_7331,N_6275,N_6859);
or U7332 (N_7332,N_6824,N_6018);
xor U7333 (N_7333,N_6104,N_6500);
nand U7334 (N_7334,N_6395,N_6597);
or U7335 (N_7335,N_6519,N_6187);
nand U7336 (N_7336,N_6576,N_6727);
xor U7337 (N_7337,N_6619,N_6268);
or U7338 (N_7338,N_6114,N_6633);
nand U7339 (N_7339,N_6254,N_6489);
or U7340 (N_7340,N_6137,N_6520);
xnor U7341 (N_7341,N_6058,N_6053);
xor U7342 (N_7342,N_6423,N_6792);
nor U7343 (N_7343,N_6526,N_6894);
and U7344 (N_7344,N_6968,N_6915);
xor U7345 (N_7345,N_6401,N_6804);
or U7346 (N_7346,N_6775,N_6008);
and U7347 (N_7347,N_6045,N_6301);
and U7348 (N_7348,N_6529,N_6965);
nand U7349 (N_7349,N_6715,N_6692);
nor U7350 (N_7350,N_6609,N_6560);
nand U7351 (N_7351,N_6835,N_6581);
nand U7352 (N_7352,N_6074,N_6077);
xor U7353 (N_7353,N_6933,N_6273);
nand U7354 (N_7354,N_6834,N_6784);
nand U7355 (N_7355,N_6204,N_6718);
and U7356 (N_7356,N_6696,N_6726);
nand U7357 (N_7357,N_6658,N_6868);
and U7358 (N_7358,N_6003,N_6763);
or U7359 (N_7359,N_6340,N_6606);
xnor U7360 (N_7360,N_6911,N_6197);
or U7361 (N_7361,N_6765,N_6716);
nor U7362 (N_7362,N_6910,N_6362);
nor U7363 (N_7363,N_6631,N_6922);
nor U7364 (N_7364,N_6482,N_6610);
and U7365 (N_7365,N_6437,N_6230);
and U7366 (N_7366,N_6394,N_6921);
xor U7367 (N_7367,N_6243,N_6888);
and U7368 (N_7368,N_6419,N_6846);
xnor U7369 (N_7369,N_6051,N_6953);
nor U7370 (N_7370,N_6860,N_6682);
nor U7371 (N_7371,N_6507,N_6783);
or U7372 (N_7372,N_6678,N_6647);
nand U7373 (N_7373,N_6603,N_6158);
xnor U7374 (N_7374,N_6733,N_6681);
xnor U7375 (N_7375,N_6016,N_6592);
or U7376 (N_7376,N_6069,N_6276);
and U7377 (N_7377,N_6324,N_6748);
and U7378 (N_7378,N_6288,N_6427);
xor U7379 (N_7379,N_6237,N_6234);
nand U7380 (N_7380,N_6674,N_6617);
and U7381 (N_7381,N_6701,N_6369);
nor U7382 (N_7382,N_6940,N_6367);
and U7383 (N_7383,N_6623,N_6452);
xor U7384 (N_7384,N_6575,N_6303);
nor U7385 (N_7385,N_6934,N_6670);
nor U7386 (N_7386,N_6181,N_6159);
xnor U7387 (N_7387,N_6998,N_6392);
and U7388 (N_7388,N_6417,N_6146);
nor U7389 (N_7389,N_6975,N_6439);
or U7390 (N_7390,N_6060,N_6683);
nand U7391 (N_7391,N_6596,N_6023);
xnor U7392 (N_7392,N_6406,N_6296);
xor U7393 (N_7393,N_6509,N_6740);
and U7394 (N_7394,N_6364,N_6002);
nand U7395 (N_7395,N_6618,N_6089);
xnor U7396 (N_7396,N_6677,N_6202);
nand U7397 (N_7397,N_6749,N_6183);
nor U7398 (N_7398,N_6874,N_6950);
xor U7399 (N_7399,N_6009,N_6877);
and U7400 (N_7400,N_6473,N_6438);
or U7401 (N_7401,N_6764,N_6774);
xor U7402 (N_7402,N_6962,N_6957);
nand U7403 (N_7403,N_6412,N_6969);
or U7404 (N_7404,N_6434,N_6062);
nand U7405 (N_7405,N_6504,N_6460);
or U7406 (N_7406,N_6486,N_6066);
or U7407 (N_7407,N_6435,N_6624);
nand U7408 (N_7408,N_6440,N_6638);
xnor U7409 (N_7409,N_6668,N_6193);
and U7410 (N_7410,N_6725,N_6028);
or U7411 (N_7411,N_6265,N_6883);
xor U7412 (N_7412,N_6153,N_6952);
nand U7413 (N_7413,N_6323,N_6492);
nor U7414 (N_7414,N_6328,N_6797);
nand U7415 (N_7415,N_6458,N_6201);
or U7416 (N_7416,N_6408,N_6163);
nand U7417 (N_7417,N_6805,N_6290);
nor U7418 (N_7418,N_6651,N_6021);
nor U7419 (N_7419,N_6221,N_6974);
xnor U7420 (N_7420,N_6661,N_6954);
nand U7421 (N_7421,N_6562,N_6287);
nand U7422 (N_7422,N_6958,N_6505);
nand U7423 (N_7423,N_6665,N_6032);
nor U7424 (N_7424,N_6088,N_6669);
nand U7425 (N_7425,N_6786,N_6356);
nand U7426 (N_7426,N_6693,N_6854);
nor U7427 (N_7427,N_6754,N_6712);
or U7428 (N_7428,N_6935,N_6663);
and U7429 (N_7429,N_6601,N_6541);
nand U7430 (N_7430,N_6266,N_6380);
xnor U7431 (N_7431,N_6298,N_6825);
nand U7432 (N_7432,N_6707,N_6487);
nor U7433 (N_7433,N_6947,N_6422);
and U7434 (N_7434,N_6823,N_6294);
and U7435 (N_7435,N_6844,N_6403);
nand U7436 (N_7436,N_6742,N_6720);
nand U7437 (N_7437,N_6694,N_6384);
and U7438 (N_7438,N_6117,N_6318);
nand U7439 (N_7439,N_6220,N_6059);
nand U7440 (N_7440,N_6544,N_6928);
nor U7441 (N_7441,N_6049,N_6598);
or U7442 (N_7442,N_6964,N_6516);
xor U7443 (N_7443,N_6445,N_6750);
and U7444 (N_7444,N_6743,N_6152);
xor U7445 (N_7445,N_6776,N_6345);
or U7446 (N_7446,N_6527,N_6814);
and U7447 (N_7447,N_6227,N_6664);
nand U7448 (N_7448,N_6425,N_6831);
and U7449 (N_7449,N_6350,N_6085);
nand U7450 (N_7450,N_6547,N_6132);
xor U7451 (N_7451,N_6620,N_6554);
and U7452 (N_7452,N_6518,N_6100);
and U7453 (N_7453,N_6207,N_6891);
or U7454 (N_7454,N_6240,N_6798);
xor U7455 (N_7455,N_6352,N_6182);
and U7456 (N_7456,N_6025,N_6113);
nand U7457 (N_7457,N_6980,N_6997);
nor U7458 (N_7458,N_6845,N_6161);
nor U7459 (N_7459,N_6881,N_6024);
nor U7460 (N_7460,N_6981,N_6467);
nand U7461 (N_7461,N_6898,N_6455);
and U7462 (N_7462,N_6131,N_6496);
nand U7463 (N_7463,N_6385,N_6708);
xor U7464 (N_7464,N_6232,N_6734);
nor U7465 (N_7465,N_6192,N_6198);
nor U7466 (N_7466,N_6082,N_6931);
nand U7467 (N_7467,N_6636,N_6905);
xnor U7468 (N_7468,N_6816,N_6397);
xor U7469 (N_7469,N_6657,N_6102);
xor U7470 (N_7470,N_6642,N_6134);
nand U7471 (N_7471,N_6063,N_6447);
xnor U7472 (N_7472,N_6031,N_6913);
or U7473 (N_7473,N_6263,N_6376);
or U7474 (N_7474,N_6895,N_6833);
nor U7475 (N_7475,N_6226,N_6264);
and U7476 (N_7476,N_6138,N_6523);
or U7477 (N_7477,N_6595,N_6081);
nand U7478 (N_7478,N_6978,N_6410);
nor U7479 (N_7479,N_6557,N_6228);
nor U7480 (N_7480,N_6334,N_6528);
or U7481 (N_7481,N_6840,N_6600);
and U7482 (N_7482,N_6154,N_6128);
nor U7483 (N_7483,N_6020,N_6485);
nand U7484 (N_7484,N_6830,N_6632);
or U7485 (N_7485,N_6982,N_6912);
or U7486 (N_7486,N_6065,N_6851);
and U7487 (N_7487,N_6721,N_6553);
nor U7488 (N_7488,N_6839,N_6724);
nor U7489 (N_7489,N_6863,N_6475);
or U7490 (N_7490,N_6442,N_6491);
and U7491 (N_7491,N_6281,N_6530);
nand U7492 (N_7492,N_6685,N_6320);
xor U7493 (N_7493,N_6767,N_6585);
nor U7494 (N_7494,N_6745,N_6398);
or U7495 (N_7495,N_6366,N_6464);
nor U7496 (N_7496,N_6880,N_6091);
nor U7497 (N_7497,N_6244,N_6605);
or U7498 (N_7498,N_6305,N_6612);
nand U7499 (N_7499,N_6941,N_6329);
xnor U7500 (N_7500,N_6701,N_6048);
nor U7501 (N_7501,N_6781,N_6596);
or U7502 (N_7502,N_6457,N_6349);
xnor U7503 (N_7503,N_6657,N_6094);
nor U7504 (N_7504,N_6541,N_6573);
or U7505 (N_7505,N_6824,N_6583);
xnor U7506 (N_7506,N_6469,N_6334);
nand U7507 (N_7507,N_6965,N_6144);
nand U7508 (N_7508,N_6657,N_6991);
and U7509 (N_7509,N_6852,N_6630);
and U7510 (N_7510,N_6322,N_6907);
nand U7511 (N_7511,N_6353,N_6017);
and U7512 (N_7512,N_6758,N_6625);
nand U7513 (N_7513,N_6356,N_6237);
xor U7514 (N_7514,N_6877,N_6922);
and U7515 (N_7515,N_6975,N_6758);
nand U7516 (N_7516,N_6751,N_6346);
nor U7517 (N_7517,N_6595,N_6537);
or U7518 (N_7518,N_6583,N_6248);
or U7519 (N_7519,N_6353,N_6499);
nor U7520 (N_7520,N_6648,N_6407);
or U7521 (N_7521,N_6295,N_6403);
or U7522 (N_7522,N_6375,N_6999);
nand U7523 (N_7523,N_6319,N_6120);
and U7524 (N_7524,N_6239,N_6607);
nor U7525 (N_7525,N_6416,N_6014);
and U7526 (N_7526,N_6848,N_6684);
nand U7527 (N_7527,N_6022,N_6236);
and U7528 (N_7528,N_6258,N_6371);
nor U7529 (N_7529,N_6300,N_6105);
or U7530 (N_7530,N_6405,N_6630);
and U7531 (N_7531,N_6214,N_6687);
or U7532 (N_7532,N_6719,N_6078);
and U7533 (N_7533,N_6936,N_6797);
nand U7534 (N_7534,N_6919,N_6123);
or U7535 (N_7535,N_6595,N_6171);
nor U7536 (N_7536,N_6765,N_6522);
nand U7537 (N_7537,N_6810,N_6399);
nand U7538 (N_7538,N_6141,N_6983);
xor U7539 (N_7539,N_6029,N_6097);
nand U7540 (N_7540,N_6279,N_6152);
or U7541 (N_7541,N_6575,N_6789);
nand U7542 (N_7542,N_6621,N_6627);
nor U7543 (N_7543,N_6066,N_6751);
or U7544 (N_7544,N_6125,N_6092);
nand U7545 (N_7545,N_6523,N_6241);
nand U7546 (N_7546,N_6756,N_6294);
nand U7547 (N_7547,N_6485,N_6926);
xnor U7548 (N_7548,N_6339,N_6203);
nor U7549 (N_7549,N_6050,N_6989);
and U7550 (N_7550,N_6983,N_6768);
and U7551 (N_7551,N_6511,N_6243);
or U7552 (N_7552,N_6065,N_6620);
xor U7553 (N_7553,N_6123,N_6700);
or U7554 (N_7554,N_6007,N_6792);
xnor U7555 (N_7555,N_6135,N_6045);
nor U7556 (N_7556,N_6413,N_6545);
and U7557 (N_7557,N_6708,N_6876);
nor U7558 (N_7558,N_6633,N_6764);
and U7559 (N_7559,N_6402,N_6866);
nand U7560 (N_7560,N_6732,N_6489);
and U7561 (N_7561,N_6430,N_6814);
nand U7562 (N_7562,N_6286,N_6291);
nor U7563 (N_7563,N_6023,N_6485);
or U7564 (N_7564,N_6199,N_6183);
nor U7565 (N_7565,N_6958,N_6137);
and U7566 (N_7566,N_6510,N_6610);
or U7567 (N_7567,N_6800,N_6053);
nand U7568 (N_7568,N_6574,N_6184);
nand U7569 (N_7569,N_6542,N_6061);
nand U7570 (N_7570,N_6036,N_6433);
nor U7571 (N_7571,N_6785,N_6118);
or U7572 (N_7572,N_6432,N_6394);
xor U7573 (N_7573,N_6431,N_6055);
nand U7574 (N_7574,N_6555,N_6899);
nand U7575 (N_7575,N_6965,N_6013);
and U7576 (N_7576,N_6591,N_6384);
nand U7577 (N_7577,N_6956,N_6472);
nor U7578 (N_7578,N_6532,N_6350);
or U7579 (N_7579,N_6413,N_6451);
xnor U7580 (N_7580,N_6735,N_6334);
xnor U7581 (N_7581,N_6062,N_6864);
nor U7582 (N_7582,N_6037,N_6936);
or U7583 (N_7583,N_6509,N_6895);
xnor U7584 (N_7584,N_6494,N_6750);
nor U7585 (N_7585,N_6486,N_6820);
nor U7586 (N_7586,N_6158,N_6081);
nand U7587 (N_7587,N_6413,N_6004);
nand U7588 (N_7588,N_6983,N_6223);
nor U7589 (N_7589,N_6825,N_6755);
nand U7590 (N_7590,N_6747,N_6270);
nand U7591 (N_7591,N_6302,N_6735);
nor U7592 (N_7592,N_6318,N_6548);
xor U7593 (N_7593,N_6429,N_6980);
nor U7594 (N_7594,N_6524,N_6471);
nor U7595 (N_7595,N_6651,N_6315);
and U7596 (N_7596,N_6660,N_6720);
or U7597 (N_7597,N_6541,N_6494);
nand U7598 (N_7598,N_6778,N_6273);
nand U7599 (N_7599,N_6360,N_6010);
xor U7600 (N_7600,N_6715,N_6025);
nand U7601 (N_7601,N_6382,N_6799);
and U7602 (N_7602,N_6457,N_6959);
or U7603 (N_7603,N_6188,N_6873);
nand U7604 (N_7604,N_6488,N_6404);
and U7605 (N_7605,N_6882,N_6590);
or U7606 (N_7606,N_6921,N_6854);
nand U7607 (N_7607,N_6860,N_6611);
nand U7608 (N_7608,N_6287,N_6658);
nand U7609 (N_7609,N_6960,N_6603);
xnor U7610 (N_7610,N_6947,N_6653);
nor U7611 (N_7611,N_6725,N_6534);
and U7612 (N_7612,N_6960,N_6513);
nand U7613 (N_7613,N_6025,N_6828);
nor U7614 (N_7614,N_6273,N_6929);
nor U7615 (N_7615,N_6584,N_6102);
or U7616 (N_7616,N_6711,N_6243);
or U7617 (N_7617,N_6786,N_6658);
xnor U7618 (N_7618,N_6541,N_6994);
and U7619 (N_7619,N_6549,N_6217);
and U7620 (N_7620,N_6323,N_6112);
nor U7621 (N_7621,N_6553,N_6299);
nand U7622 (N_7622,N_6109,N_6719);
xnor U7623 (N_7623,N_6373,N_6594);
nor U7624 (N_7624,N_6946,N_6007);
nor U7625 (N_7625,N_6754,N_6199);
xnor U7626 (N_7626,N_6882,N_6207);
nor U7627 (N_7627,N_6703,N_6246);
and U7628 (N_7628,N_6908,N_6000);
xnor U7629 (N_7629,N_6840,N_6489);
nand U7630 (N_7630,N_6893,N_6895);
nor U7631 (N_7631,N_6102,N_6735);
and U7632 (N_7632,N_6534,N_6699);
and U7633 (N_7633,N_6550,N_6705);
xnor U7634 (N_7634,N_6673,N_6910);
nor U7635 (N_7635,N_6010,N_6751);
nand U7636 (N_7636,N_6840,N_6480);
nand U7637 (N_7637,N_6112,N_6593);
nand U7638 (N_7638,N_6807,N_6607);
and U7639 (N_7639,N_6951,N_6529);
and U7640 (N_7640,N_6496,N_6626);
nor U7641 (N_7641,N_6121,N_6799);
and U7642 (N_7642,N_6254,N_6891);
nor U7643 (N_7643,N_6980,N_6935);
and U7644 (N_7644,N_6657,N_6649);
and U7645 (N_7645,N_6499,N_6315);
xor U7646 (N_7646,N_6343,N_6477);
nand U7647 (N_7647,N_6802,N_6543);
nor U7648 (N_7648,N_6102,N_6153);
or U7649 (N_7649,N_6028,N_6147);
nand U7650 (N_7650,N_6465,N_6513);
or U7651 (N_7651,N_6797,N_6848);
and U7652 (N_7652,N_6740,N_6029);
nand U7653 (N_7653,N_6709,N_6913);
nand U7654 (N_7654,N_6307,N_6338);
xnor U7655 (N_7655,N_6578,N_6735);
xnor U7656 (N_7656,N_6303,N_6309);
nand U7657 (N_7657,N_6375,N_6776);
and U7658 (N_7658,N_6242,N_6955);
and U7659 (N_7659,N_6935,N_6149);
xor U7660 (N_7660,N_6481,N_6136);
xor U7661 (N_7661,N_6145,N_6650);
nor U7662 (N_7662,N_6612,N_6811);
nand U7663 (N_7663,N_6097,N_6837);
nand U7664 (N_7664,N_6265,N_6768);
and U7665 (N_7665,N_6162,N_6188);
nand U7666 (N_7666,N_6338,N_6385);
and U7667 (N_7667,N_6840,N_6712);
nor U7668 (N_7668,N_6161,N_6859);
xor U7669 (N_7669,N_6913,N_6887);
and U7670 (N_7670,N_6995,N_6781);
xor U7671 (N_7671,N_6018,N_6024);
xor U7672 (N_7672,N_6340,N_6479);
or U7673 (N_7673,N_6573,N_6083);
nor U7674 (N_7674,N_6173,N_6300);
xnor U7675 (N_7675,N_6458,N_6891);
nand U7676 (N_7676,N_6339,N_6158);
nor U7677 (N_7677,N_6008,N_6093);
nor U7678 (N_7678,N_6580,N_6802);
xnor U7679 (N_7679,N_6276,N_6090);
or U7680 (N_7680,N_6977,N_6356);
nand U7681 (N_7681,N_6024,N_6250);
xor U7682 (N_7682,N_6889,N_6081);
or U7683 (N_7683,N_6446,N_6702);
and U7684 (N_7684,N_6439,N_6758);
nand U7685 (N_7685,N_6731,N_6076);
or U7686 (N_7686,N_6372,N_6757);
or U7687 (N_7687,N_6098,N_6902);
or U7688 (N_7688,N_6299,N_6028);
and U7689 (N_7689,N_6234,N_6447);
nand U7690 (N_7690,N_6363,N_6595);
or U7691 (N_7691,N_6809,N_6203);
nand U7692 (N_7692,N_6672,N_6976);
or U7693 (N_7693,N_6431,N_6737);
or U7694 (N_7694,N_6201,N_6205);
xnor U7695 (N_7695,N_6814,N_6886);
and U7696 (N_7696,N_6116,N_6778);
and U7697 (N_7697,N_6779,N_6763);
and U7698 (N_7698,N_6673,N_6205);
xor U7699 (N_7699,N_6340,N_6964);
or U7700 (N_7700,N_6553,N_6691);
nor U7701 (N_7701,N_6723,N_6954);
xnor U7702 (N_7702,N_6316,N_6308);
xor U7703 (N_7703,N_6861,N_6232);
xnor U7704 (N_7704,N_6528,N_6392);
nor U7705 (N_7705,N_6710,N_6412);
xor U7706 (N_7706,N_6584,N_6060);
and U7707 (N_7707,N_6671,N_6547);
nand U7708 (N_7708,N_6735,N_6491);
or U7709 (N_7709,N_6605,N_6594);
xor U7710 (N_7710,N_6260,N_6138);
and U7711 (N_7711,N_6077,N_6397);
xnor U7712 (N_7712,N_6858,N_6646);
or U7713 (N_7713,N_6110,N_6026);
nor U7714 (N_7714,N_6915,N_6294);
or U7715 (N_7715,N_6706,N_6996);
or U7716 (N_7716,N_6985,N_6403);
or U7717 (N_7717,N_6988,N_6438);
nand U7718 (N_7718,N_6418,N_6229);
and U7719 (N_7719,N_6462,N_6734);
or U7720 (N_7720,N_6784,N_6986);
nor U7721 (N_7721,N_6088,N_6423);
nor U7722 (N_7722,N_6343,N_6315);
or U7723 (N_7723,N_6074,N_6314);
or U7724 (N_7724,N_6921,N_6251);
xnor U7725 (N_7725,N_6266,N_6888);
xnor U7726 (N_7726,N_6480,N_6738);
or U7727 (N_7727,N_6433,N_6447);
xor U7728 (N_7728,N_6691,N_6207);
nor U7729 (N_7729,N_6486,N_6733);
or U7730 (N_7730,N_6813,N_6245);
nor U7731 (N_7731,N_6918,N_6530);
and U7732 (N_7732,N_6241,N_6184);
nand U7733 (N_7733,N_6354,N_6513);
nor U7734 (N_7734,N_6052,N_6077);
and U7735 (N_7735,N_6565,N_6800);
or U7736 (N_7736,N_6308,N_6718);
nor U7737 (N_7737,N_6802,N_6578);
nand U7738 (N_7738,N_6648,N_6698);
nand U7739 (N_7739,N_6188,N_6661);
nand U7740 (N_7740,N_6446,N_6019);
nand U7741 (N_7741,N_6834,N_6994);
or U7742 (N_7742,N_6250,N_6452);
or U7743 (N_7743,N_6281,N_6566);
or U7744 (N_7744,N_6946,N_6051);
or U7745 (N_7745,N_6402,N_6992);
and U7746 (N_7746,N_6016,N_6810);
nor U7747 (N_7747,N_6442,N_6959);
or U7748 (N_7748,N_6634,N_6875);
nor U7749 (N_7749,N_6473,N_6948);
xnor U7750 (N_7750,N_6788,N_6210);
xnor U7751 (N_7751,N_6146,N_6136);
xnor U7752 (N_7752,N_6752,N_6169);
or U7753 (N_7753,N_6777,N_6882);
or U7754 (N_7754,N_6700,N_6340);
xnor U7755 (N_7755,N_6403,N_6193);
or U7756 (N_7756,N_6577,N_6194);
xnor U7757 (N_7757,N_6989,N_6800);
xnor U7758 (N_7758,N_6797,N_6074);
nor U7759 (N_7759,N_6993,N_6894);
nor U7760 (N_7760,N_6596,N_6527);
nand U7761 (N_7761,N_6699,N_6333);
or U7762 (N_7762,N_6065,N_6307);
and U7763 (N_7763,N_6245,N_6499);
nor U7764 (N_7764,N_6186,N_6735);
nor U7765 (N_7765,N_6128,N_6823);
and U7766 (N_7766,N_6131,N_6550);
or U7767 (N_7767,N_6181,N_6124);
or U7768 (N_7768,N_6244,N_6934);
and U7769 (N_7769,N_6085,N_6057);
xnor U7770 (N_7770,N_6910,N_6942);
xor U7771 (N_7771,N_6409,N_6237);
nor U7772 (N_7772,N_6954,N_6039);
nor U7773 (N_7773,N_6050,N_6553);
and U7774 (N_7774,N_6706,N_6968);
or U7775 (N_7775,N_6931,N_6120);
and U7776 (N_7776,N_6512,N_6279);
nor U7777 (N_7777,N_6170,N_6051);
and U7778 (N_7778,N_6295,N_6454);
xnor U7779 (N_7779,N_6746,N_6436);
nand U7780 (N_7780,N_6189,N_6837);
and U7781 (N_7781,N_6327,N_6147);
nor U7782 (N_7782,N_6556,N_6190);
xnor U7783 (N_7783,N_6097,N_6080);
nor U7784 (N_7784,N_6837,N_6197);
and U7785 (N_7785,N_6208,N_6784);
xor U7786 (N_7786,N_6778,N_6877);
nand U7787 (N_7787,N_6155,N_6120);
xnor U7788 (N_7788,N_6326,N_6714);
nand U7789 (N_7789,N_6194,N_6890);
nand U7790 (N_7790,N_6837,N_6264);
or U7791 (N_7791,N_6956,N_6619);
or U7792 (N_7792,N_6092,N_6776);
or U7793 (N_7793,N_6725,N_6708);
or U7794 (N_7794,N_6662,N_6740);
or U7795 (N_7795,N_6708,N_6334);
xor U7796 (N_7796,N_6483,N_6979);
nand U7797 (N_7797,N_6415,N_6429);
nand U7798 (N_7798,N_6495,N_6612);
and U7799 (N_7799,N_6493,N_6171);
or U7800 (N_7800,N_6994,N_6172);
nand U7801 (N_7801,N_6945,N_6577);
nand U7802 (N_7802,N_6386,N_6036);
and U7803 (N_7803,N_6678,N_6577);
and U7804 (N_7804,N_6424,N_6193);
and U7805 (N_7805,N_6260,N_6591);
or U7806 (N_7806,N_6999,N_6507);
xor U7807 (N_7807,N_6582,N_6999);
and U7808 (N_7808,N_6940,N_6144);
nor U7809 (N_7809,N_6844,N_6768);
nand U7810 (N_7810,N_6411,N_6492);
xnor U7811 (N_7811,N_6131,N_6487);
or U7812 (N_7812,N_6315,N_6123);
nor U7813 (N_7813,N_6975,N_6901);
or U7814 (N_7814,N_6026,N_6201);
and U7815 (N_7815,N_6056,N_6362);
or U7816 (N_7816,N_6729,N_6465);
and U7817 (N_7817,N_6092,N_6174);
nor U7818 (N_7818,N_6295,N_6770);
and U7819 (N_7819,N_6730,N_6567);
or U7820 (N_7820,N_6517,N_6344);
or U7821 (N_7821,N_6739,N_6224);
xor U7822 (N_7822,N_6572,N_6871);
and U7823 (N_7823,N_6339,N_6192);
or U7824 (N_7824,N_6925,N_6206);
nor U7825 (N_7825,N_6446,N_6189);
or U7826 (N_7826,N_6825,N_6922);
nand U7827 (N_7827,N_6859,N_6058);
xor U7828 (N_7828,N_6259,N_6147);
nand U7829 (N_7829,N_6280,N_6131);
xnor U7830 (N_7830,N_6191,N_6271);
nand U7831 (N_7831,N_6325,N_6121);
nand U7832 (N_7832,N_6423,N_6801);
and U7833 (N_7833,N_6001,N_6217);
or U7834 (N_7834,N_6052,N_6569);
xor U7835 (N_7835,N_6627,N_6218);
or U7836 (N_7836,N_6007,N_6623);
nor U7837 (N_7837,N_6712,N_6422);
xnor U7838 (N_7838,N_6435,N_6604);
nand U7839 (N_7839,N_6192,N_6718);
and U7840 (N_7840,N_6381,N_6622);
nor U7841 (N_7841,N_6575,N_6744);
xnor U7842 (N_7842,N_6591,N_6677);
and U7843 (N_7843,N_6539,N_6006);
nand U7844 (N_7844,N_6249,N_6106);
nor U7845 (N_7845,N_6665,N_6445);
nand U7846 (N_7846,N_6577,N_6660);
nor U7847 (N_7847,N_6820,N_6805);
nand U7848 (N_7848,N_6846,N_6731);
nor U7849 (N_7849,N_6904,N_6652);
nand U7850 (N_7850,N_6375,N_6155);
or U7851 (N_7851,N_6864,N_6358);
nor U7852 (N_7852,N_6062,N_6586);
xnor U7853 (N_7853,N_6078,N_6159);
xor U7854 (N_7854,N_6732,N_6021);
xor U7855 (N_7855,N_6982,N_6650);
or U7856 (N_7856,N_6353,N_6681);
and U7857 (N_7857,N_6822,N_6794);
or U7858 (N_7858,N_6968,N_6634);
nor U7859 (N_7859,N_6314,N_6911);
xnor U7860 (N_7860,N_6758,N_6870);
nand U7861 (N_7861,N_6696,N_6169);
xor U7862 (N_7862,N_6581,N_6565);
and U7863 (N_7863,N_6401,N_6039);
nor U7864 (N_7864,N_6511,N_6526);
xor U7865 (N_7865,N_6820,N_6030);
nand U7866 (N_7866,N_6519,N_6448);
and U7867 (N_7867,N_6349,N_6678);
or U7868 (N_7868,N_6089,N_6578);
and U7869 (N_7869,N_6003,N_6924);
or U7870 (N_7870,N_6518,N_6339);
xor U7871 (N_7871,N_6291,N_6621);
nand U7872 (N_7872,N_6405,N_6080);
and U7873 (N_7873,N_6937,N_6725);
nor U7874 (N_7874,N_6599,N_6981);
nand U7875 (N_7875,N_6117,N_6680);
nand U7876 (N_7876,N_6677,N_6436);
xnor U7877 (N_7877,N_6329,N_6559);
nor U7878 (N_7878,N_6924,N_6596);
and U7879 (N_7879,N_6518,N_6163);
nand U7880 (N_7880,N_6352,N_6997);
xnor U7881 (N_7881,N_6022,N_6324);
and U7882 (N_7882,N_6955,N_6506);
and U7883 (N_7883,N_6001,N_6444);
or U7884 (N_7884,N_6721,N_6277);
or U7885 (N_7885,N_6650,N_6586);
or U7886 (N_7886,N_6643,N_6270);
or U7887 (N_7887,N_6862,N_6501);
nand U7888 (N_7888,N_6861,N_6164);
xnor U7889 (N_7889,N_6433,N_6749);
nand U7890 (N_7890,N_6163,N_6697);
or U7891 (N_7891,N_6980,N_6035);
nor U7892 (N_7892,N_6429,N_6189);
and U7893 (N_7893,N_6725,N_6910);
nand U7894 (N_7894,N_6223,N_6921);
xnor U7895 (N_7895,N_6706,N_6067);
xor U7896 (N_7896,N_6108,N_6819);
or U7897 (N_7897,N_6775,N_6465);
or U7898 (N_7898,N_6239,N_6099);
and U7899 (N_7899,N_6982,N_6450);
nor U7900 (N_7900,N_6084,N_6981);
xor U7901 (N_7901,N_6737,N_6896);
and U7902 (N_7902,N_6419,N_6614);
and U7903 (N_7903,N_6264,N_6369);
xor U7904 (N_7904,N_6431,N_6969);
or U7905 (N_7905,N_6459,N_6017);
and U7906 (N_7906,N_6225,N_6407);
or U7907 (N_7907,N_6362,N_6781);
nand U7908 (N_7908,N_6469,N_6330);
or U7909 (N_7909,N_6340,N_6154);
nand U7910 (N_7910,N_6538,N_6675);
nor U7911 (N_7911,N_6944,N_6365);
or U7912 (N_7912,N_6473,N_6926);
nand U7913 (N_7913,N_6798,N_6927);
and U7914 (N_7914,N_6325,N_6626);
or U7915 (N_7915,N_6469,N_6481);
xor U7916 (N_7916,N_6862,N_6269);
nand U7917 (N_7917,N_6046,N_6826);
or U7918 (N_7918,N_6129,N_6038);
xnor U7919 (N_7919,N_6646,N_6157);
and U7920 (N_7920,N_6223,N_6595);
nor U7921 (N_7921,N_6046,N_6441);
or U7922 (N_7922,N_6296,N_6747);
xor U7923 (N_7923,N_6648,N_6065);
xnor U7924 (N_7924,N_6698,N_6241);
nand U7925 (N_7925,N_6969,N_6708);
nor U7926 (N_7926,N_6385,N_6575);
and U7927 (N_7927,N_6373,N_6112);
nand U7928 (N_7928,N_6788,N_6144);
xnor U7929 (N_7929,N_6831,N_6119);
nand U7930 (N_7930,N_6343,N_6225);
nand U7931 (N_7931,N_6000,N_6645);
xnor U7932 (N_7932,N_6354,N_6092);
nor U7933 (N_7933,N_6184,N_6600);
xnor U7934 (N_7934,N_6499,N_6747);
nor U7935 (N_7935,N_6244,N_6758);
or U7936 (N_7936,N_6842,N_6213);
xnor U7937 (N_7937,N_6873,N_6291);
nand U7938 (N_7938,N_6897,N_6339);
or U7939 (N_7939,N_6508,N_6203);
xor U7940 (N_7940,N_6610,N_6156);
or U7941 (N_7941,N_6758,N_6960);
and U7942 (N_7942,N_6041,N_6823);
nand U7943 (N_7943,N_6914,N_6931);
or U7944 (N_7944,N_6187,N_6224);
xor U7945 (N_7945,N_6136,N_6964);
and U7946 (N_7946,N_6049,N_6902);
xnor U7947 (N_7947,N_6913,N_6994);
xor U7948 (N_7948,N_6208,N_6116);
or U7949 (N_7949,N_6457,N_6124);
or U7950 (N_7950,N_6067,N_6349);
xor U7951 (N_7951,N_6152,N_6816);
and U7952 (N_7952,N_6175,N_6372);
or U7953 (N_7953,N_6390,N_6557);
nor U7954 (N_7954,N_6553,N_6794);
and U7955 (N_7955,N_6679,N_6884);
xnor U7956 (N_7956,N_6626,N_6631);
xor U7957 (N_7957,N_6232,N_6592);
nor U7958 (N_7958,N_6548,N_6600);
nor U7959 (N_7959,N_6193,N_6029);
nand U7960 (N_7960,N_6803,N_6915);
or U7961 (N_7961,N_6862,N_6487);
nor U7962 (N_7962,N_6573,N_6991);
or U7963 (N_7963,N_6980,N_6189);
nor U7964 (N_7964,N_6465,N_6904);
nand U7965 (N_7965,N_6711,N_6802);
or U7966 (N_7966,N_6043,N_6278);
nor U7967 (N_7967,N_6921,N_6509);
or U7968 (N_7968,N_6503,N_6556);
nand U7969 (N_7969,N_6215,N_6316);
nor U7970 (N_7970,N_6125,N_6825);
nor U7971 (N_7971,N_6264,N_6326);
and U7972 (N_7972,N_6654,N_6943);
nand U7973 (N_7973,N_6401,N_6428);
or U7974 (N_7974,N_6986,N_6857);
xor U7975 (N_7975,N_6435,N_6913);
nor U7976 (N_7976,N_6144,N_6526);
or U7977 (N_7977,N_6084,N_6363);
or U7978 (N_7978,N_6032,N_6551);
nor U7979 (N_7979,N_6322,N_6765);
xor U7980 (N_7980,N_6541,N_6234);
nor U7981 (N_7981,N_6382,N_6171);
xor U7982 (N_7982,N_6502,N_6228);
nor U7983 (N_7983,N_6727,N_6954);
or U7984 (N_7984,N_6747,N_6167);
and U7985 (N_7985,N_6197,N_6365);
nand U7986 (N_7986,N_6223,N_6865);
nand U7987 (N_7987,N_6241,N_6565);
xnor U7988 (N_7988,N_6241,N_6276);
nor U7989 (N_7989,N_6415,N_6249);
or U7990 (N_7990,N_6274,N_6916);
nand U7991 (N_7991,N_6404,N_6164);
and U7992 (N_7992,N_6956,N_6813);
and U7993 (N_7993,N_6319,N_6961);
and U7994 (N_7994,N_6511,N_6597);
nand U7995 (N_7995,N_6683,N_6180);
nand U7996 (N_7996,N_6121,N_6495);
and U7997 (N_7997,N_6093,N_6604);
nand U7998 (N_7998,N_6092,N_6951);
and U7999 (N_7999,N_6359,N_6161);
and U8000 (N_8000,N_7866,N_7926);
and U8001 (N_8001,N_7968,N_7376);
or U8002 (N_8002,N_7411,N_7166);
and U8003 (N_8003,N_7727,N_7980);
xor U8004 (N_8004,N_7536,N_7995);
nor U8005 (N_8005,N_7712,N_7885);
nor U8006 (N_8006,N_7976,N_7513);
xnor U8007 (N_8007,N_7650,N_7342);
nor U8008 (N_8008,N_7941,N_7842);
nand U8009 (N_8009,N_7231,N_7948);
or U8010 (N_8010,N_7073,N_7213);
nor U8011 (N_8011,N_7293,N_7200);
xnor U8012 (N_8012,N_7978,N_7544);
nand U8013 (N_8013,N_7330,N_7349);
nand U8014 (N_8014,N_7253,N_7701);
or U8015 (N_8015,N_7967,N_7657);
or U8016 (N_8016,N_7945,N_7923);
or U8017 (N_8017,N_7837,N_7327);
or U8018 (N_8018,N_7595,N_7529);
nand U8019 (N_8019,N_7101,N_7408);
and U8020 (N_8020,N_7805,N_7568);
nand U8021 (N_8021,N_7096,N_7173);
xor U8022 (N_8022,N_7074,N_7791);
nor U8023 (N_8023,N_7737,N_7675);
and U8024 (N_8024,N_7627,N_7548);
nand U8025 (N_8025,N_7754,N_7400);
nand U8026 (N_8026,N_7619,N_7746);
nor U8027 (N_8027,N_7933,N_7680);
nor U8028 (N_8028,N_7849,N_7134);
xor U8029 (N_8029,N_7394,N_7336);
and U8030 (N_8030,N_7181,N_7296);
nand U8031 (N_8031,N_7000,N_7566);
and U8032 (N_8032,N_7884,N_7080);
or U8033 (N_8033,N_7780,N_7749);
nand U8034 (N_8034,N_7028,N_7475);
or U8035 (N_8035,N_7035,N_7130);
xnor U8036 (N_8036,N_7441,N_7076);
nand U8037 (N_8037,N_7894,N_7869);
or U8038 (N_8038,N_7397,N_7452);
xor U8039 (N_8039,N_7410,N_7267);
nand U8040 (N_8040,N_7579,N_7072);
xor U8041 (N_8041,N_7345,N_7565);
or U8042 (N_8042,N_7038,N_7915);
nor U8043 (N_8043,N_7422,N_7956);
nor U8044 (N_8044,N_7703,N_7402);
or U8045 (N_8045,N_7347,N_7370);
nor U8046 (N_8046,N_7390,N_7716);
xor U8047 (N_8047,N_7199,N_7026);
nor U8048 (N_8048,N_7818,N_7725);
or U8049 (N_8049,N_7556,N_7042);
xnor U8050 (N_8050,N_7799,N_7205);
and U8051 (N_8051,N_7584,N_7647);
and U8052 (N_8052,N_7501,N_7547);
and U8053 (N_8053,N_7508,N_7460);
and U8054 (N_8054,N_7616,N_7116);
and U8055 (N_8055,N_7520,N_7624);
and U8056 (N_8056,N_7263,N_7734);
nand U8057 (N_8057,N_7141,N_7132);
or U8058 (N_8058,N_7399,N_7832);
nand U8059 (N_8059,N_7273,N_7490);
and U8060 (N_8060,N_7123,N_7722);
nand U8061 (N_8061,N_7021,N_7011);
nand U8062 (N_8062,N_7241,N_7449);
nand U8063 (N_8063,N_7121,N_7177);
xnor U8064 (N_8064,N_7808,N_7672);
and U8065 (N_8065,N_7900,N_7685);
xor U8066 (N_8066,N_7360,N_7835);
nand U8067 (N_8067,N_7748,N_7505);
xor U8068 (N_8068,N_7937,N_7502);
nor U8069 (N_8069,N_7631,N_7554);
nand U8070 (N_8070,N_7796,N_7625);
nand U8071 (N_8071,N_7588,N_7389);
xor U8072 (N_8072,N_7645,N_7421);
nor U8073 (N_8073,N_7939,N_7215);
xnor U8074 (N_8074,N_7474,N_7683);
nand U8075 (N_8075,N_7087,N_7462);
nor U8076 (N_8076,N_7227,N_7740);
or U8077 (N_8077,N_7160,N_7829);
or U8078 (N_8078,N_7586,N_7320);
xor U8079 (N_8079,N_7644,N_7498);
nand U8080 (N_8080,N_7735,N_7664);
nor U8081 (N_8081,N_7391,N_7515);
or U8082 (N_8082,N_7761,N_7052);
or U8083 (N_8083,N_7783,N_7585);
and U8084 (N_8084,N_7507,N_7797);
xnor U8085 (N_8085,N_7610,N_7274);
xnor U8086 (N_8086,N_7518,N_7673);
and U8087 (N_8087,N_7363,N_7299);
nand U8088 (N_8088,N_7744,N_7487);
and U8089 (N_8089,N_7867,N_7353);
xnor U8090 (N_8090,N_7942,N_7691);
nand U8091 (N_8091,N_7925,N_7162);
or U8092 (N_8092,N_7553,N_7886);
or U8093 (N_8093,N_7247,N_7341);
nand U8094 (N_8094,N_7752,N_7214);
nand U8095 (N_8095,N_7872,N_7146);
or U8096 (N_8096,N_7949,N_7036);
and U8097 (N_8097,N_7029,N_7033);
and U8098 (N_8098,N_7030,N_7233);
xor U8099 (N_8099,N_7950,N_7031);
nor U8100 (N_8100,N_7965,N_7963);
nor U8101 (N_8101,N_7527,N_7732);
nand U8102 (N_8102,N_7420,N_7534);
nor U8103 (N_8103,N_7469,N_7789);
nor U8104 (N_8104,N_7383,N_7537);
and U8105 (N_8105,N_7380,N_7929);
or U8106 (N_8106,N_7984,N_7180);
nor U8107 (N_8107,N_7179,N_7377);
or U8108 (N_8108,N_7632,N_7742);
or U8109 (N_8109,N_7739,N_7064);
nor U8110 (N_8110,N_7897,N_7438);
or U8111 (N_8111,N_7541,N_7145);
nand U8112 (N_8112,N_7670,N_7510);
or U8113 (N_8113,N_7993,N_7889);
and U8114 (N_8114,N_7830,N_7238);
and U8115 (N_8115,N_7729,N_7539);
nand U8116 (N_8116,N_7086,N_7395);
or U8117 (N_8117,N_7615,N_7335);
or U8118 (N_8118,N_7663,N_7398);
or U8119 (N_8119,N_7388,N_7458);
and U8120 (N_8120,N_7059,N_7065);
nand U8121 (N_8121,N_7142,N_7094);
nor U8122 (N_8122,N_7165,N_7099);
xor U8123 (N_8123,N_7300,N_7730);
nand U8124 (N_8124,N_7229,N_7150);
or U8125 (N_8125,N_7479,N_7283);
nand U8126 (N_8126,N_7882,N_7759);
and U8127 (N_8127,N_7480,N_7082);
or U8128 (N_8128,N_7062,N_7843);
nand U8129 (N_8129,N_7856,N_7540);
nand U8130 (N_8130,N_7662,N_7887);
and U8131 (N_8131,N_7545,N_7079);
xnor U8132 (N_8132,N_7551,N_7039);
and U8133 (N_8133,N_7317,N_7138);
nor U8134 (N_8134,N_7671,N_7940);
or U8135 (N_8135,N_7590,N_7677);
nor U8136 (N_8136,N_7111,N_7450);
or U8137 (N_8137,N_7324,N_7599);
nor U8138 (N_8138,N_7307,N_7212);
and U8139 (N_8139,N_7055,N_7758);
nand U8140 (N_8140,N_7118,N_7374);
and U8141 (N_8141,N_7580,N_7931);
nand U8142 (N_8142,N_7041,N_7120);
nand U8143 (N_8143,N_7668,N_7092);
and U8144 (N_8144,N_7239,N_7523);
nor U8145 (N_8145,N_7351,N_7543);
nand U8146 (N_8146,N_7218,N_7291);
and U8147 (N_8147,N_7305,N_7877);
nor U8148 (N_8148,N_7252,N_7718);
and U8149 (N_8149,N_7917,N_7892);
xnor U8150 (N_8150,N_7436,N_7924);
xor U8151 (N_8151,N_7025,N_7051);
nor U8152 (N_8152,N_7382,N_7425);
xor U8153 (N_8153,N_7004,N_7655);
nand U8154 (N_8154,N_7969,N_7847);
nor U8155 (N_8155,N_7578,N_7868);
nor U8156 (N_8156,N_7741,N_7432);
nor U8157 (N_8157,N_7192,N_7198);
nor U8158 (N_8158,N_7699,N_7017);
xnor U8159 (N_8159,N_7640,N_7093);
xnor U8160 (N_8160,N_7652,N_7778);
nor U8161 (N_8161,N_7827,N_7187);
or U8162 (N_8162,N_7107,N_7356);
or U8163 (N_8163,N_7012,N_7817);
nor U8164 (N_8164,N_7986,N_7295);
and U8165 (N_8165,N_7128,N_7174);
or U8166 (N_8166,N_7801,N_7069);
and U8167 (N_8167,N_7800,N_7254);
nand U8168 (N_8168,N_7845,N_7463);
and U8169 (N_8169,N_7521,N_7044);
nor U8170 (N_8170,N_7085,N_7522);
nand U8171 (N_8171,N_7635,N_7137);
nor U8172 (N_8172,N_7560,N_7824);
nand U8173 (N_8173,N_7467,N_7598);
and U8174 (N_8174,N_7806,N_7169);
and U8175 (N_8175,N_7176,N_7256);
xnor U8176 (N_8176,N_7709,N_7228);
and U8177 (N_8177,N_7157,N_7952);
nor U8178 (N_8178,N_7765,N_7098);
nor U8179 (N_8179,N_7015,N_7045);
or U8180 (N_8180,N_7442,N_7981);
and U8181 (N_8181,N_7816,N_7184);
nor U8182 (N_8182,N_7495,N_7183);
or U8183 (N_8183,N_7569,N_7953);
nand U8184 (N_8184,N_7155,N_7589);
xnor U8185 (N_8185,N_7710,N_7282);
xor U8186 (N_8186,N_7998,N_7958);
and U8187 (N_8187,N_7607,N_7182);
or U8188 (N_8188,N_7606,N_7658);
or U8189 (N_8189,N_7384,N_7678);
or U8190 (N_8190,N_7996,N_7839);
nand U8191 (N_8191,N_7368,N_7704);
xor U8192 (N_8192,N_7144,N_7831);
nand U8193 (N_8193,N_7403,N_7911);
nand U8194 (N_8194,N_7100,N_7466);
and U8195 (N_8195,N_7339,N_7990);
xnor U8196 (N_8196,N_7129,N_7001);
and U8197 (N_8197,N_7999,N_7433);
nor U8198 (N_8198,N_7623,N_7104);
nor U8199 (N_8199,N_7891,N_7190);
nor U8200 (N_8200,N_7208,N_7840);
and U8201 (N_8201,N_7636,N_7524);
nand U8202 (N_8202,N_7637,N_7426);
or U8203 (N_8203,N_7440,N_7938);
nor U8204 (N_8204,N_7914,N_7966);
and U8205 (N_8205,N_7626,N_7535);
nor U8206 (N_8206,N_7642,N_7696);
xor U8207 (N_8207,N_7620,N_7597);
and U8208 (N_8208,N_7930,N_7406);
nand U8209 (N_8209,N_7189,N_7465);
nand U8210 (N_8210,N_7812,N_7878);
or U8211 (N_8211,N_7147,N_7552);
nor U8212 (N_8212,N_7898,N_7334);
and U8213 (N_8213,N_7201,N_7024);
nor U8214 (N_8214,N_7815,N_7684);
or U8215 (N_8215,N_7769,N_7312);
xnor U8216 (N_8216,N_7301,N_7081);
nor U8217 (N_8217,N_7210,N_7514);
or U8218 (N_8218,N_7804,N_7387);
and U8219 (N_8219,N_7875,N_7302);
xor U8220 (N_8220,N_7982,N_7451);
nand U8221 (N_8221,N_7946,N_7193);
or U8222 (N_8222,N_7723,N_7570);
xnor U8223 (N_8223,N_7861,N_7496);
nor U8224 (N_8224,N_7902,N_7666);
xor U8225 (N_8225,N_7279,N_7161);
and U8226 (N_8226,N_7373,N_7023);
nor U8227 (N_8227,N_7826,N_7484);
and U8228 (N_8228,N_7857,N_7220);
xnor U8229 (N_8229,N_7124,N_7136);
or U8230 (N_8230,N_7054,N_7656);
nor U8231 (N_8231,N_7516,N_7057);
nand U8232 (N_8232,N_7795,N_7242);
or U8233 (N_8233,N_7821,N_7468);
nor U8234 (N_8234,N_7272,N_7600);
nand U8235 (N_8235,N_7550,N_7932);
nand U8236 (N_8236,N_7910,N_7255);
nor U8237 (N_8237,N_7077,N_7720);
xor U8238 (N_8238,N_7794,N_7083);
nor U8239 (N_8239,N_7018,N_7890);
xnor U8240 (N_8240,N_7280,N_7322);
or U8241 (N_8241,N_7027,N_7776);
xor U8242 (N_8242,N_7439,N_7454);
or U8243 (N_8243,N_7191,N_7158);
and U8244 (N_8244,N_7862,N_7010);
xor U8245 (N_8245,N_7332,N_7604);
nand U8246 (N_8246,N_7261,N_7594);
nor U8247 (N_8247,N_7067,N_7807);
nand U8248 (N_8248,N_7477,N_7893);
nand U8249 (N_8249,N_7367,N_7489);
and U8250 (N_8250,N_7037,N_7206);
nand U8251 (N_8251,N_7316,N_7298);
nor U8252 (N_8252,N_7908,N_7943);
nor U8253 (N_8253,N_7154,N_7097);
xnor U8254 (N_8254,N_7770,N_7500);
xor U8255 (N_8255,N_7721,N_7309);
or U8256 (N_8256,N_7863,N_7369);
nand U8257 (N_8257,N_7413,N_7230);
or U8258 (N_8258,N_7575,N_7582);
nand U8259 (N_8259,N_7983,N_7738);
and U8260 (N_8260,N_7549,N_7592);
nand U8261 (N_8261,N_7921,N_7927);
xor U8262 (N_8262,N_7936,N_7194);
nor U8263 (N_8263,N_7424,N_7702);
xnor U8264 (N_8264,N_7412,N_7131);
nor U8265 (N_8265,N_7453,N_7728);
or U8266 (N_8266,N_7667,N_7630);
nor U8267 (N_8267,N_7928,N_7841);
or U8268 (N_8268,N_7782,N_7343);
or U8269 (N_8269,N_7517,N_7538);
nand U8270 (N_8270,N_7622,N_7577);
xnor U8271 (N_8271,N_7511,N_7143);
or U8272 (N_8272,N_7651,N_7994);
nand U8273 (N_8273,N_7276,N_7971);
nor U8274 (N_8274,N_7638,N_7557);
nor U8275 (N_8275,N_7119,N_7314);
xor U8276 (N_8276,N_7961,N_7409);
xor U8277 (N_8277,N_7488,N_7234);
or U8278 (N_8278,N_7755,N_7034);
and U8279 (N_8279,N_7944,N_7331);
and U8280 (N_8280,N_7763,N_7355);
and U8281 (N_8281,N_7661,N_7281);
and U8282 (N_8282,N_7504,N_7957);
xnor U8283 (N_8283,N_7879,N_7286);
and U8284 (N_8284,N_7243,N_7292);
or U8285 (N_8285,N_7698,N_7266);
nor U8286 (N_8286,N_7581,N_7471);
nand U8287 (N_8287,N_7546,N_7591);
nand U8288 (N_8288,N_7270,N_7905);
xnor U8289 (N_8289,N_7009,N_7649);
xnor U8290 (N_8290,N_7972,N_7526);
nor U8291 (N_8291,N_7559,N_7906);
xor U8292 (N_8292,N_7692,N_7583);
xnor U8293 (N_8293,N_7563,N_7310);
nand U8294 (N_8294,N_7779,N_7365);
xnor U8295 (N_8295,N_7753,N_7386);
or U8296 (N_8296,N_7315,N_7311);
and U8297 (N_8297,N_7020,N_7895);
xor U8298 (N_8298,N_7864,N_7003);
xor U8299 (N_8299,N_7714,N_7974);
or U8300 (N_8300,N_7275,N_7955);
nor U8301 (N_8301,N_7108,N_7002);
or U8302 (N_8302,N_7113,N_7777);
nor U8303 (N_8303,N_7987,N_7991);
xor U8304 (N_8304,N_7329,N_7428);
nand U8305 (N_8305,N_7171,N_7676);
xor U8306 (N_8306,N_7114,N_7525);
or U8307 (N_8307,N_7809,N_7935);
nor U8308 (N_8308,N_7013,N_7985);
nand U8309 (N_8309,N_7854,N_7874);
or U8310 (N_8310,N_7660,N_7139);
or U8311 (N_8311,N_7919,N_7870);
xnor U8312 (N_8312,N_7325,N_7481);
and U8313 (N_8313,N_7418,N_7697);
and U8314 (N_8314,N_7750,N_7688);
nand U8315 (N_8315,N_7690,N_7032);
xor U8316 (N_8316,N_7609,N_7532);
and U8317 (N_8317,N_7122,N_7531);
and U8318 (N_8318,N_7603,N_7608);
and U8319 (N_8319,N_7922,N_7308);
nor U8320 (N_8320,N_7357,N_7485);
nand U8321 (N_8321,N_7512,N_7235);
and U8322 (N_8322,N_7061,N_7639);
xor U8323 (N_8323,N_7416,N_7681);
nand U8324 (N_8324,N_7979,N_7249);
and U8325 (N_8325,N_7593,N_7125);
xor U8326 (N_8326,N_7708,N_7197);
or U8327 (N_8327,N_7833,N_7088);
and U8328 (N_8328,N_7558,N_7223);
xnor U8329 (N_8329,N_7112,N_7430);
nor U8330 (N_8330,N_7359,N_7989);
xnor U8331 (N_8331,N_7686,N_7682);
and U8332 (N_8332,N_7068,N_7792);
xnor U8333 (N_8333,N_7509,N_7251);
or U8334 (N_8334,N_7070,N_7448);
nor U8335 (N_8335,N_7934,N_7572);
xor U8336 (N_8336,N_7762,N_7617);
nor U8337 (N_8337,N_7419,N_7287);
nand U8338 (N_8338,N_7333,N_7457);
xor U8339 (N_8339,N_7225,N_7271);
and U8340 (N_8340,N_7156,N_7056);
nand U8341 (N_8341,N_7602,N_7019);
and U8342 (N_8342,N_7423,N_7605);
nand U8343 (N_8343,N_7715,N_7354);
nor U8344 (N_8344,N_7711,N_7674);
and U8345 (N_8345,N_7110,N_7385);
nand U8346 (N_8346,N_7836,N_7918);
or U8347 (N_8347,N_7016,N_7071);
nand U8348 (N_8348,N_7008,N_7264);
and U8349 (N_8349,N_7084,N_7445);
or U8350 (N_8350,N_7811,N_7294);
nor U8351 (N_8351,N_7043,N_7596);
nor U8352 (N_8352,N_7170,N_7319);
or U8353 (N_8353,N_7903,N_7050);
nand U8354 (N_8354,N_7066,N_7262);
nand U8355 (N_8355,N_7105,N_7289);
or U8356 (N_8356,N_7375,N_7216);
nand U8357 (N_8357,N_7973,N_7834);
nand U8358 (N_8358,N_7211,N_7063);
nand U8359 (N_8359,N_7571,N_7899);
or U8360 (N_8360,N_7858,N_7250);
nor U8361 (N_8361,N_7371,N_7876);
xor U8362 (N_8362,N_7773,N_7148);
or U8363 (N_8363,N_7259,N_7172);
or U8364 (N_8364,N_7846,N_7920);
nand U8365 (N_8365,N_7186,N_7562);
nand U8366 (N_8366,N_7163,N_7290);
xnor U8367 (N_8367,N_7694,N_7951);
nor U8368 (N_8368,N_7786,N_7323);
nor U8369 (N_8369,N_7232,N_7724);
nor U8370 (N_8370,N_7153,N_7313);
xor U8371 (N_8371,N_7258,N_7352);
or U8372 (N_8372,N_7326,N_7306);
xnor U8373 (N_8373,N_7407,N_7446);
xnor U8374 (N_8374,N_7321,N_7106);
or U8375 (N_8375,N_7404,N_7528);
nand U8376 (N_8376,N_7530,N_7366);
xor U8377 (N_8377,N_7135,N_7246);
xnor U8378 (N_8378,N_7771,N_7459);
or U8379 (N_8379,N_7344,N_7090);
nand U8380 (N_8380,N_7859,N_7493);
or U8381 (N_8381,N_7431,N_7444);
nor U8382 (N_8382,N_7822,N_7049);
or U8383 (N_8383,N_7237,N_7358);
xor U8384 (N_8384,N_7954,N_7178);
or U8385 (N_8385,N_7717,N_7047);
or U8386 (N_8386,N_7888,N_7005);
nand U8387 (N_8387,N_7964,N_7587);
nor U8388 (N_8388,N_7614,N_7519);
nor U8389 (N_8389,N_7303,N_7719);
or U8390 (N_8390,N_7629,N_7643);
or U8391 (N_8391,N_7401,N_7909);
and U8392 (N_8392,N_7494,N_7803);
nor U8393 (N_8393,N_7379,N_7288);
or U8394 (N_8394,N_7217,N_7304);
xnor U8395 (N_8395,N_7533,N_7185);
nand U8396 (N_8396,N_7126,N_7297);
xor U8397 (N_8397,N_7764,N_7415);
nand U8398 (N_8398,N_7766,N_7574);
and U8399 (N_8399,N_7871,N_7434);
nand U8400 (N_8400,N_7492,N_7464);
xor U8401 (N_8401,N_7959,N_7634);
xor U8402 (N_8402,N_7705,N_7784);
and U8403 (N_8403,N_7700,N_7679);
nand U8404 (N_8404,N_7695,N_7053);
and U8405 (N_8405,N_7346,N_7167);
nor U8406 (N_8406,N_7209,N_7621);
or U8407 (N_8407,N_7455,N_7855);
xor U8408 (N_8408,N_7653,N_7499);
nor U8409 (N_8409,N_7881,N_7244);
nand U8410 (N_8410,N_7022,N_7736);
nor U8411 (N_8411,N_7497,N_7338);
and U8412 (N_8412,N_7473,N_7798);
or U8413 (N_8413,N_7788,N_7693);
nor U8414 (N_8414,N_7149,N_7058);
and U8415 (N_8415,N_7476,N_7561);
xnor U8416 (N_8416,N_7601,N_7103);
and U8417 (N_8417,N_7853,N_7248);
xor U8418 (N_8418,N_7665,N_7977);
or U8419 (N_8419,N_7745,N_7506);
nor U8420 (N_8420,N_7767,N_7960);
or U8421 (N_8421,N_7361,N_7268);
xnor U8422 (N_8422,N_7912,N_7350);
nor U8423 (N_8423,N_7486,N_7414);
xor U8424 (N_8424,N_7221,N_7285);
nand U8425 (N_8425,N_7151,N_7706);
or U8426 (N_8426,N_7204,N_7751);
and U8427 (N_8427,N_7277,N_7340);
and U8428 (N_8428,N_7427,N_7947);
nand U8429 (N_8429,N_7393,N_7040);
nor U8430 (N_8430,N_7284,N_7417);
xor U8431 (N_8431,N_7195,N_7362);
or U8432 (N_8432,N_7896,N_7447);
nand U8433 (N_8433,N_7318,N_7916);
nor U8434 (N_8434,N_7175,N_7851);
nor U8435 (N_8435,N_7774,N_7203);
nor U8436 (N_8436,N_7823,N_7726);
and U8437 (N_8437,N_7852,N_7348);
and U8438 (N_8438,N_7873,N_7226);
nand U8439 (N_8439,N_7628,N_7269);
or U8440 (N_8440,N_7848,N_7785);
and U8441 (N_8441,N_7265,N_7975);
xnor U8442 (N_8442,N_7461,N_7611);
xor U8443 (N_8443,N_7865,N_7819);
and U8444 (N_8444,N_7278,N_7483);
xnor U8445 (N_8445,N_7641,N_7901);
nand U8446 (N_8446,N_7396,N_7372);
nand U8447 (N_8447,N_7775,N_7364);
and U8448 (N_8448,N_7613,N_7576);
xnor U8449 (N_8449,N_7236,N_7102);
or U8450 (N_8450,N_7659,N_7109);
or U8451 (N_8451,N_7757,N_7988);
or U8452 (N_8452,N_7612,N_7810);
or U8453 (N_8453,N_7075,N_7707);
and U8454 (N_8454,N_7542,N_7224);
nor U8455 (N_8455,N_7207,N_7140);
xor U8456 (N_8456,N_7007,N_7095);
or U8457 (N_8457,N_7115,N_7825);
xor U8458 (N_8458,N_7733,N_7772);
or U8459 (N_8459,N_7219,N_7913);
or U8460 (N_8460,N_7970,N_7567);
xor U8461 (N_8461,N_7159,N_7743);
nor U8462 (N_8462,N_7202,N_7731);
xnor U8463 (N_8463,N_7669,N_7907);
and U8464 (N_8464,N_7337,N_7747);
or U8465 (N_8465,N_7381,N_7117);
nand U8466 (N_8466,N_7850,N_7756);
or U8467 (N_8467,N_7048,N_7222);
nand U8468 (N_8468,N_7618,N_7482);
nor U8469 (N_8469,N_7188,N_7646);
nor U8470 (N_8470,N_7687,N_7491);
nor U8471 (N_8471,N_7573,N_7880);
and U8472 (N_8472,N_7014,N_7713);
or U8473 (N_8473,N_7760,N_7820);
and U8474 (N_8474,N_7429,N_7470);
nand U8475 (N_8475,N_7790,N_7555);
xor U8476 (N_8476,N_7443,N_7883);
and U8477 (N_8477,N_7472,N_7392);
nand U8478 (N_8478,N_7240,N_7564);
nand U8479 (N_8479,N_7787,N_7127);
or U8480 (N_8480,N_7405,N_7328);
nor U8481 (N_8481,N_7828,N_7152);
nor U8482 (N_8482,N_7793,N_7904);
nor U8483 (N_8483,N_7814,N_7633);
nor U8484 (N_8484,N_7078,N_7456);
nor U8485 (N_8485,N_7245,N_7435);
and U8486 (N_8486,N_7133,N_7844);
nand U8487 (N_8487,N_7997,N_7768);
and U8488 (N_8488,N_7437,N_7654);
xnor U8489 (N_8489,N_7838,N_7164);
or U8490 (N_8490,N_7802,N_7091);
and U8491 (N_8491,N_7257,N_7378);
nor U8492 (N_8492,N_7478,N_7689);
xnor U8493 (N_8493,N_7196,N_7781);
nand U8494 (N_8494,N_7006,N_7089);
or U8495 (N_8495,N_7992,N_7046);
nor U8496 (N_8496,N_7060,N_7860);
nand U8497 (N_8497,N_7648,N_7168);
xor U8498 (N_8498,N_7813,N_7260);
and U8499 (N_8499,N_7503,N_7962);
nor U8500 (N_8500,N_7818,N_7364);
nor U8501 (N_8501,N_7504,N_7616);
nand U8502 (N_8502,N_7656,N_7997);
and U8503 (N_8503,N_7801,N_7601);
and U8504 (N_8504,N_7991,N_7164);
nand U8505 (N_8505,N_7828,N_7374);
nor U8506 (N_8506,N_7598,N_7995);
nand U8507 (N_8507,N_7839,N_7051);
and U8508 (N_8508,N_7771,N_7740);
xnor U8509 (N_8509,N_7748,N_7076);
or U8510 (N_8510,N_7173,N_7247);
and U8511 (N_8511,N_7579,N_7578);
xor U8512 (N_8512,N_7665,N_7283);
and U8513 (N_8513,N_7000,N_7221);
and U8514 (N_8514,N_7296,N_7673);
xor U8515 (N_8515,N_7735,N_7959);
or U8516 (N_8516,N_7934,N_7433);
nand U8517 (N_8517,N_7706,N_7245);
nand U8518 (N_8518,N_7813,N_7575);
and U8519 (N_8519,N_7840,N_7864);
and U8520 (N_8520,N_7665,N_7732);
and U8521 (N_8521,N_7665,N_7205);
nor U8522 (N_8522,N_7888,N_7012);
and U8523 (N_8523,N_7512,N_7350);
and U8524 (N_8524,N_7984,N_7216);
and U8525 (N_8525,N_7472,N_7665);
xor U8526 (N_8526,N_7575,N_7324);
nand U8527 (N_8527,N_7752,N_7024);
nand U8528 (N_8528,N_7947,N_7492);
nand U8529 (N_8529,N_7613,N_7091);
and U8530 (N_8530,N_7784,N_7412);
nor U8531 (N_8531,N_7056,N_7885);
or U8532 (N_8532,N_7235,N_7092);
nor U8533 (N_8533,N_7561,N_7236);
or U8534 (N_8534,N_7133,N_7460);
and U8535 (N_8535,N_7968,N_7199);
nand U8536 (N_8536,N_7917,N_7457);
and U8537 (N_8537,N_7631,N_7144);
nor U8538 (N_8538,N_7767,N_7029);
nand U8539 (N_8539,N_7149,N_7388);
and U8540 (N_8540,N_7887,N_7820);
nand U8541 (N_8541,N_7766,N_7226);
nand U8542 (N_8542,N_7811,N_7258);
nor U8543 (N_8543,N_7097,N_7492);
or U8544 (N_8544,N_7200,N_7295);
nor U8545 (N_8545,N_7370,N_7562);
nand U8546 (N_8546,N_7686,N_7054);
nand U8547 (N_8547,N_7093,N_7983);
and U8548 (N_8548,N_7105,N_7870);
or U8549 (N_8549,N_7876,N_7331);
xnor U8550 (N_8550,N_7100,N_7943);
and U8551 (N_8551,N_7459,N_7451);
and U8552 (N_8552,N_7706,N_7662);
nor U8553 (N_8553,N_7730,N_7108);
or U8554 (N_8554,N_7000,N_7070);
xnor U8555 (N_8555,N_7485,N_7319);
or U8556 (N_8556,N_7378,N_7724);
and U8557 (N_8557,N_7247,N_7085);
and U8558 (N_8558,N_7202,N_7915);
xnor U8559 (N_8559,N_7604,N_7475);
nor U8560 (N_8560,N_7082,N_7829);
and U8561 (N_8561,N_7445,N_7623);
nand U8562 (N_8562,N_7545,N_7975);
and U8563 (N_8563,N_7759,N_7143);
nand U8564 (N_8564,N_7345,N_7907);
and U8565 (N_8565,N_7367,N_7530);
nor U8566 (N_8566,N_7400,N_7278);
and U8567 (N_8567,N_7515,N_7689);
and U8568 (N_8568,N_7781,N_7489);
xor U8569 (N_8569,N_7824,N_7245);
nor U8570 (N_8570,N_7470,N_7220);
xor U8571 (N_8571,N_7226,N_7457);
or U8572 (N_8572,N_7562,N_7844);
nand U8573 (N_8573,N_7882,N_7498);
xnor U8574 (N_8574,N_7054,N_7590);
nor U8575 (N_8575,N_7054,N_7516);
and U8576 (N_8576,N_7000,N_7309);
nor U8577 (N_8577,N_7667,N_7144);
and U8578 (N_8578,N_7576,N_7775);
and U8579 (N_8579,N_7023,N_7889);
or U8580 (N_8580,N_7437,N_7256);
and U8581 (N_8581,N_7751,N_7697);
xor U8582 (N_8582,N_7868,N_7645);
nor U8583 (N_8583,N_7531,N_7628);
and U8584 (N_8584,N_7177,N_7045);
xnor U8585 (N_8585,N_7283,N_7174);
and U8586 (N_8586,N_7710,N_7774);
xnor U8587 (N_8587,N_7362,N_7209);
or U8588 (N_8588,N_7553,N_7707);
or U8589 (N_8589,N_7636,N_7771);
nand U8590 (N_8590,N_7833,N_7139);
or U8591 (N_8591,N_7188,N_7984);
and U8592 (N_8592,N_7563,N_7989);
nor U8593 (N_8593,N_7892,N_7912);
and U8594 (N_8594,N_7394,N_7311);
or U8595 (N_8595,N_7849,N_7223);
xnor U8596 (N_8596,N_7161,N_7774);
nor U8597 (N_8597,N_7729,N_7097);
nor U8598 (N_8598,N_7247,N_7263);
nor U8599 (N_8599,N_7669,N_7993);
nor U8600 (N_8600,N_7445,N_7945);
nand U8601 (N_8601,N_7909,N_7852);
and U8602 (N_8602,N_7941,N_7160);
nor U8603 (N_8603,N_7024,N_7156);
nor U8604 (N_8604,N_7105,N_7563);
and U8605 (N_8605,N_7921,N_7737);
nand U8606 (N_8606,N_7271,N_7953);
xnor U8607 (N_8607,N_7095,N_7934);
nand U8608 (N_8608,N_7017,N_7228);
xnor U8609 (N_8609,N_7568,N_7717);
nor U8610 (N_8610,N_7134,N_7946);
or U8611 (N_8611,N_7273,N_7981);
nor U8612 (N_8612,N_7808,N_7471);
nor U8613 (N_8613,N_7062,N_7718);
xor U8614 (N_8614,N_7005,N_7412);
nand U8615 (N_8615,N_7565,N_7321);
nor U8616 (N_8616,N_7648,N_7748);
nand U8617 (N_8617,N_7546,N_7924);
nand U8618 (N_8618,N_7386,N_7313);
nand U8619 (N_8619,N_7566,N_7005);
xnor U8620 (N_8620,N_7668,N_7581);
or U8621 (N_8621,N_7819,N_7334);
and U8622 (N_8622,N_7786,N_7238);
or U8623 (N_8623,N_7514,N_7551);
or U8624 (N_8624,N_7890,N_7784);
nor U8625 (N_8625,N_7360,N_7198);
or U8626 (N_8626,N_7177,N_7531);
nand U8627 (N_8627,N_7709,N_7245);
or U8628 (N_8628,N_7767,N_7659);
nand U8629 (N_8629,N_7135,N_7617);
nor U8630 (N_8630,N_7783,N_7498);
nand U8631 (N_8631,N_7719,N_7217);
or U8632 (N_8632,N_7642,N_7261);
and U8633 (N_8633,N_7478,N_7123);
or U8634 (N_8634,N_7409,N_7603);
xnor U8635 (N_8635,N_7115,N_7054);
xnor U8636 (N_8636,N_7756,N_7357);
and U8637 (N_8637,N_7811,N_7647);
nor U8638 (N_8638,N_7147,N_7722);
xnor U8639 (N_8639,N_7912,N_7990);
nor U8640 (N_8640,N_7165,N_7215);
nor U8641 (N_8641,N_7056,N_7763);
xor U8642 (N_8642,N_7681,N_7717);
and U8643 (N_8643,N_7048,N_7399);
nor U8644 (N_8644,N_7395,N_7855);
and U8645 (N_8645,N_7929,N_7925);
or U8646 (N_8646,N_7056,N_7316);
nand U8647 (N_8647,N_7710,N_7215);
xnor U8648 (N_8648,N_7041,N_7487);
and U8649 (N_8649,N_7143,N_7001);
nor U8650 (N_8650,N_7545,N_7638);
or U8651 (N_8651,N_7580,N_7699);
nand U8652 (N_8652,N_7393,N_7096);
and U8653 (N_8653,N_7414,N_7750);
nand U8654 (N_8654,N_7377,N_7650);
and U8655 (N_8655,N_7005,N_7282);
nor U8656 (N_8656,N_7921,N_7408);
nand U8657 (N_8657,N_7385,N_7820);
nor U8658 (N_8658,N_7293,N_7232);
xnor U8659 (N_8659,N_7836,N_7371);
nor U8660 (N_8660,N_7907,N_7459);
xnor U8661 (N_8661,N_7806,N_7695);
nor U8662 (N_8662,N_7720,N_7820);
nor U8663 (N_8663,N_7702,N_7039);
nor U8664 (N_8664,N_7465,N_7498);
or U8665 (N_8665,N_7809,N_7002);
nor U8666 (N_8666,N_7367,N_7272);
xnor U8667 (N_8667,N_7841,N_7628);
nor U8668 (N_8668,N_7541,N_7242);
xnor U8669 (N_8669,N_7971,N_7697);
and U8670 (N_8670,N_7847,N_7391);
xnor U8671 (N_8671,N_7505,N_7772);
and U8672 (N_8672,N_7737,N_7097);
and U8673 (N_8673,N_7305,N_7214);
nor U8674 (N_8674,N_7030,N_7749);
or U8675 (N_8675,N_7544,N_7393);
or U8676 (N_8676,N_7049,N_7934);
and U8677 (N_8677,N_7760,N_7482);
nor U8678 (N_8678,N_7223,N_7693);
xnor U8679 (N_8679,N_7243,N_7104);
and U8680 (N_8680,N_7119,N_7671);
or U8681 (N_8681,N_7318,N_7799);
nand U8682 (N_8682,N_7787,N_7210);
or U8683 (N_8683,N_7031,N_7019);
or U8684 (N_8684,N_7510,N_7944);
or U8685 (N_8685,N_7433,N_7693);
or U8686 (N_8686,N_7580,N_7942);
nor U8687 (N_8687,N_7904,N_7115);
nor U8688 (N_8688,N_7850,N_7277);
or U8689 (N_8689,N_7700,N_7067);
and U8690 (N_8690,N_7111,N_7073);
nand U8691 (N_8691,N_7128,N_7125);
nand U8692 (N_8692,N_7733,N_7469);
nand U8693 (N_8693,N_7880,N_7451);
nor U8694 (N_8694,N_7140,N_7898);
xor U8695 (N_8695,N_7567,N_7505);
and U8696 (N_8696,N_7454,N_7203);
or U8697 (N_8697,N_7599,N_7094);
nor U8698 (N_8698,N_7637,N_7059);
xnor U8699 (N_8699,N_7174,N_7447);
or U8700 (N_8700,N_7312,N_7436);
nand U8701 (N_8701,N_7193,N_7578);
xnor U8702 (N_8702,N_7685,N_7391);
nor U8703 (N_8703,N_7015,N_7226);
nand U8704 (N_8704,N_7520,N_7121);
xor U8705 (N_8705,N_7359,N_7748);
nor U8706 (N_8706,N_7862,N_7318);
nor U8707 (N_8707,N_7667,N_7200);
xor U8708 (N_8708,N_7033,N_7025);
nand U8709 (N_8709,N_7528,N_7122);
xor U8710 (N_8710,N_7608,N_7249);
nand U8711 (N_8711,N_7368,N_7645);
xor U8712 (N_8712,N_7240,N_7419);
xor U8713 (N_8713,N_7151,N_7516);
nor U8714 (N_8714,N_7701,N_7914);
and U8715 (N_8715,N_7463,N_7917);
and U8716 (N_8716,N_7107,N_7565);
xor U8717 (N_8717,N_7817,N_7520);
and U8718 (N_8718,N_7695,N_7158);
xor U8719 (N_8719,N_7111,N_7696);
nand U8720 (N_8720,N_7990,N_7083);
and U8721 (N_8721,N_7864,N_7219);
xor U8722 (N_8722,N_7514,N_7592);
or U8723 (N_8723,N_7547,N_7131);
xor U8724 (N_8724,N_7140,N_7341);
or U8725 (N_8725,N_7610,N_7422);
xnor U8726 (N_8726,N_7683,N_7732);
or U8727 (N_8727,N_7315,N_7962);
nor U8728 (N_8728,N_7692,N_7809);
nor U8729 (N_8729,N_7831,N_7310);
nor U8730 (N_8730,N_7820,N_7963);
nor U8731 (N_8731,N_7999,N_7833);
nand U8732 (N_8732,N_7508,N_7163);
nor U8733 (N_8733,N_7573,N_7871);
nor U8734 (N_8734,N_7253,N_7863);
nor U8735 (N_8735,N_7383,N_7645);
nor U8736 (N_8736,N_7035,N_7698);
nor U8737 (N_8737,N_7358,N_7118);
and U8738 (N_8738,N_7864,N_7937);
nor U8739 (N_8739,N_7244,N_7691);
or U8740 (N_8740,N_7885,N_7585);
nand U8741 (N_8741,N_7179,N_7309);
and U8742 (N_8742,N_7060,N_7388);
or U8743 (N_8743,N_7984,N_7288);
nand U8744 (N_8744,N_7549,N_7203);
xnor U8745 (N_8745,N_7867,N_7547);
xor U8746 (N_8746,N_7885,N_7170);
or U8747 (N_8747,N_7356,N_7345);
and U8748 (N_8748,N_7450,N_7384);
nor U8749 (N_8749,N_7571,N_7412);
xor U8750 (N_8750,N_7777,N_7529);
and U8751 (N_8751,N_7930,N_7071);
nor U8752 (N_8752,N_7636,N_7708);
or U8753 (N_8753,N_7591,N_7544);
xnor U8754 (N_8754,N_7812,N_7724);
nand U8755 (N_8755,N_7334,N_7737);
nand U8756 (N_8756,N_7136,N_7554);
and U8757 (N_8757,N_7455,N_7669);
xor U8758 (N_8758,N_7646,N_7450);
and U8759 (N_8759,N_7979,N_7422);
xor U8760 (N_8760,N_7390,N_7695);
and U8761 (N_8761,N_7335,N_7939);
or U8762 (N_8762,N_7405,N_7846);
xnor U8763 (N_8763,N_7321,N_7306);
nor U8764 (N_8764,N_7910,N_7936);
nand U8765 (N_8765,N_7184,N_7654);
nand U8766 (N_8766,N_7363,N_7865);
or U8767 (N_8767,N_7599,N_7739);
xnor U8768 (N_8768,N_7815,N_7449);
xnor U8769 (N_8769,N_7602,N_7645);
nor U8770 (N_8770,N_7105,N_7741);
nand U8771 (N_8771,N_7144,N_7813);
nand U8772 (N_8772,N_7574,N_7477);
nor U8773 (N_8773,N_7779,N_7833);
xor U8774 (N_8774,N_7825,N_7405);
xor U8775 (N_8775,N_7885,N_7815);
nor U8776 (N_8776,N_7430,N_7356);
xnor U8777 (N_8777,N_7876,N_7614);
nand U8778 (N_8778,N_7779,N_7703);
and U8779 (N_8779,N_7306,N_7099);
and U8780 (N_8780,N_7798,N_7383);
xor U8781 (N_8781,N_7723,N_7708);
nor U8782 (N_8782,N_7105,N_7301);
nor U8783 (N_8783,N_7181,N_7816);
nor U8784 (N_8784,N_7892,N_7776);
nand U8785 (N_8785,N_7335,N_7284);
nor U8786 (N_8786,N_7967,N_7342);
xnor U8787 (N_8787,N_7192,N_7759);
nand U8788 (N_8788,N_7469,N_7426);
and U8789 (N_8789,N_7116,N_7192);
xnor U8790 (N_8790,N_7137,N_7640);
and U8791 (N_8791,N_7059,N_7616);
nand U8792 (N_8792,N_7161,N_7731);
nand U8793 (N_8793,N_7274,N_7470);
and U8794 (N_8794,N_7173,N_7866);
nor U8795 (N_8795,N_7416,N_7554);
and U8796 (N_8796,N_7194,N_7507);
xnor U8797 (N_8797,N_7391,N_7667);
nand U8798 (N_8798,N_7883,N_7495);
and U8799 (N_8799,N_7238,N_7499);
xor U8800 (N_8800,N_7351,N_7560);
xnor U8801 (N_8801,N_7457,N_7194);
xnor U8802 (N_8802,N_7934,N_7091);
nand U8803 (N_8803,N_7339,N_7401);
nor U8804 (N_8804,N_7879,N_7243);
or U8805 (N_8805,N_7426,N_7427);
nand U8806 (N_8806,N_7062,N_7532);
nor U8807 (N_8807,N_7958,N_7638);
or U8808 (N_8808,N_7219,N_7185);
nand U8809 (N_8809,N_7780,N_7587);
and U8810 (N_8810,N_7877,N_7824);
nand U8811 (N_8811,N_7556,N_7856);
nand U8812 (N_8812,N_7895,N_7953);
nor U8813 (N_8813,N_7059,N_7656);
xnor U8814 (N_8814,N_7410,N_7806);
or U8815 (N_8815,N_7522,N_7158);
or U8816 (N_8816,N_7350,N_7199);
xnor U8817 (N_8817,N_7225,N_7186);
nor U8818 (N_8818,N_7674,N_7278);
nor U8819 (N_8819,N_7695,N_7428);
nor U8820 (N_8820,N_7605,N_7582);
and U8821 (N_8821,N_7482,N_7275);
and U8822 (N_8822,N_7884,N_7256);
and U8823 (N_8823,N_7428,N_7762);
or U8824 (N_8824,N_7753,N_7518);
nor U8825 (N_8825,N_7277,N_7432);
nand U8826 (N_8826,N_7525,N_7958);
nand U8827 (N_8827,N_7499,N_7846);
nand U8828 (N_8828,N_7231,N_7781);
nor U8829 (N_8829,N_7080,N_7343);
or U8830 (N_8830,N_7023,N_7303);
xnor U8831 (N_8831,N_7308,N_7968);
or U8832 (N_8832,N_7815,N_7936);
nor U8833 (N_8833,N_7527,N_7574);
nand U8834 (N_8834,N_7932,N_7936);
nor U8835 (N_8835,N_7459,N_7939);
and U8836 (N_8836,N_7090,N_7212);
nor U8837 (N_8837,N_7495,N_7533);
nand U8838 (N_8838,N_7384,N_7709);
nand U8839 (N_8839,N_7667,N_7879);
and U8840 (N_8840,N_7641,N_7018);
xor U8841 (N_8841,N_7060,N_7179);
and U8842 (N_8842,N_7014,N_7560);
nand U8843 (N_8843,N_7245,N_7861);
nor U8844 (N_8844,N_7911,N_7028);
nand U8845 (N_8845,N_7796,N_7159);
nand U8846 (N_8846,N_7286,N_7835);
xnor U8847 (N_8847,N_7998,N_7907);
xor U8848 (N_8848,N_7960,N_7557);
nor U8849 (N_8849,N_7287,N_7411);
nand U8850 (N_8850,N_7846,N_7863);
nor U8851 (N_8851,N_7880,N_7513);
nand U8852 (N_8852,N_7500,N_7727);
xnor U8853 (N_8853,N_7148,N_7879);
nand U8854 (N_8854,N_7737,N_7336);
nand U8855 (N_8855,N_7570,N_7345);
nand U8856 (N_8856,N_7763,N_7378);
and U8857 (N_8857,N_7522,N_7998);
nor U8858 (N_8858,N_7076,N_7762);
or U8859 (N_8859,N_7884,N_7020);
and U8860 (N_8860,N_7637,N_7108);
nor U8861 (N_8861,N_7524,N_7335);
nor U8862 (N_8862,N_7057,N_7291);
nand U8863 (N_8863,N_7306,N_7042);
nor U8864 (N_8864,N_7112,N_7061);
and U8865 (N_8865,N_7012,N_7401);
and U8866 (N_8866,N_7164,N_7167);
nand U8867 (N_8867,N_7210,N_7434);
and U8868 (N_8868,N_7075,N_7220);
nor U8869 (N_8869,N_7167,N_7105);
nor U8870 (N_8870,N_7258,N_7992);
nand U8871 (N_8871,N_7077,N_7153);
nor U8872 (N_8872,N_7258,N_7779);
nand U8873 (N_8873,N_7549,N_7406);
nor U8874 (N_8874,N_7774,N_7275);
nor U8875 (N_8875,N_7474,N_7481);
xor U8876 (N_8876,N_7980,N_7394);
nand U8877 (N_8877,N_7216,N_7526);
xnor U8878 (N_8878,N_7269,N_7808);
nor U8879 (N_8879,N_7632,N_7737);
nor U8880 (N_8880,N_7830,N_7364);
or U8881 (N_8881,N_7225,N_7922);
or U8882 (N_8882,N_7747,N_7756);
xor U8883 (N_8883,N_7132,N_7400);
and U8884 (N_8884,N_7012,N_7959);
nand U8885 (N_8885,N_7868,N_7148);
nor U8886 (N_8886,N_7380,N_7060);
or U8887 (N_8887,N_7025,N_7308);
nor U8888 (N_8888,N_7891,N_7313);
and U8889 (N_8889,N_7315,N_7460);
nor U8890 (N_8890,N_7205,N_7618);
nor U8891 (N_8891,N_7596,N_7404);
xor U8892 (N_8892,N_7572,N_7371);
or U8893 (N_8893,N_7515,N_7434);
or U8894 (N_8894,N_7479,N_7033);
or U8895 (N_8895,N_7980,N_7502);
xnor U8896 (N_8896,N_7791,N_7599);
nor U8897 (N_8897,N_7706,N_7262);
and U8898 (N_8898,N_7623,N_7834);
nand U8899 (N_8899,N_7011,N_7335);
xnor U8900 (N_8900,N_7646,N_7125);
nand U8901 (N_8901,N_7392,N_7581);
nand U8902 (N_8902,N_7892,N_7535);
nor U8903 (N_8903,N_7707,N_7818);
xor U8904 (N_8904,N_7268,N_7385);
or U8905 (N_8905,N_7523,N_7141);
or U8906 (N_8906,N_7500,N_7390);
nor U8907 (N_8907,N_7920,N_7168);
xor U8908 (N_8908,N_7201,N_7853);
or U8909 (N_8909,N_7381,N_7611);
nand U8910 (N_8910,N_7063,N_7939);
xor U8911 (N_8911,N_7284,N_7691);
or U8912 (N_8912,N_7148,N_7074);
and U8913 (N_8913,N_7452,N_7900);
and U8914 (N_8914,N_7763,N_7157);
or U8915 (N_8915,N_7285,N_7859);
nor U8916 (N_8916,N_7219,N_7038);
nor U8917 (N_8917,N_7722,N_7527);
nor U8918 (N_8918,N_7407,N_7685);
xnor U8919 (N_8919,N_7853,N_7077);
xor U8920 (N_8920,N_7351,N_7885);
or U8921 (N_8921,N_7400,N_7752);
and U8922 (N_8922,N_7613,N_7827);
nor U8923 (N_8923,N_7173,N_7964);
nor U8924 (N_8924,N_7446,N_7382);
and U8925 (N_8925,N_7790,N_7127);
or U8926 (N_8926,N_7934,N_7148);
nor U8927 (N_8927,N_7616,N_7371);
nand U8928 (N_8928,N_7785,N_7262);
or U8929 (N_8929,N_7458,N_7959);
nor U8930 (N_8930,N_7784,N_7946);
xnor U8931 (N_8931,N_7201,N_7547);
or U8932 (N_8932,N_7051,N_7091);
or U8933 (N_8933,N_7899,N_7718);
nor U8934 (N_8934,N_7172,N_7834);
or U8935 (N_8935,N_7590,N_7152);
nand U8936 (N_8936,N_7218,N_7601);
nor U8937 (N_8937,N_7634,N_7994);
nor U8938 (N_8938,N_7580,N_7121);
nand U8939 (N_8939,N_7538,N_7529);
and U8940 (N_8940,N_7153,N_7367);
and U8941 (N_8941,N_7380,N_7569);
and U8942 (N_8942,N_7852,N_7663);
nand U8943 (N_8943,N_7985,N_7065);
or U8944 (N_8944,N_7366,N_7140);
and U8945 (N_8945,N_7192,N_7207);
xor U8946 (N_8946,N_7653,N_7759);
xor U8947 (N_8947,N_7685,N_7237);
xnor U8948 (N_8948,N_7596,N_7926);
nand U8949 (N_8949,N_7675,N_7986);
nand U8950 (N_8950,N_7167,N_7607);
nor U8951 (N_8951,N_7565,N_7444);
nand U8952 (N_8952,N_7374,N_7317);
or U8953 (N_8953,N_7898,N_7506);
nand U8954 (N_8954,N_7774,N_7869);
and U8955 (N_8955,N_7479,N_7620);
and U8956 (N_8956,N_7109,N_7765);
and U8957 (N_8957,N_7324,N_7649);
nor U8958 (N_8958,N_7421,N_7981);
nor U8959 (N_8959,N_7377,N_7135);
or U8960 (N_8960,N_7812,N_7509);
and U8961 (N_8961,N_7661,N_7532);
nor U8962 (N_8962,N_7947,N_7059);
or U8963 (N_8963,N_7444,N_7710);
nor U8964 (N_8964,N_7700,N_7172);
nand U8965 (N_8965,N_7849,N_7139);
nand U8966 (N_8966,N_7638,N_7210);
xor U8967 (N_8967,N_7174,N_7592);
or U8968 (N_8968,N_7244,N_7697);
xnor U8969 (N_8969,N_7693,N_7589);
and U8970 (N_8970,N_7017,N_7549);
and U8971 (N_8971,N_7372,N_7724);
xnor U8972 (N_8972,N_7558,N_7688);
nor U8973 (N_8973,N_7555,N_7310);
nand U8974 (N_8974,N_7603,N_7184);
nand U8975 (N_8975,N_7592,N_7355);
xor U8976 (N_8976,N_7478,N_7701);
nand U8977 (N_8977,N_7973,N_7137);
nand U8978 (N_8978,N_7856,N_7377);
xor U8979 (N_8979,N_7716,N_7857);
nor U8980 (N_8980,N_7396,N_7761);
nand U8981 (N_8981,N_7809,N_7861);
xor U8982 (N_8982,N_7819,N_7258);
nor U8983 (N_8983,N_7103,N_7162);
and U8984 (N_8984,N_7651,N_7294);
nand U8985 (N_8985,N_7303,N_7767);
and U8986 (N_8986,N_7555,N_7755);
nor U8987 (N_8987,N_7859,N_7118);
nand U8988 (N_8988,N_7106,N_7466);
xnor U8989 (N_8989,N_7557,N_7964);
nor U8990 (N_8990,N_7941,N_7024);
or U8991 (N_8991,N_7408,N_7816);
nand U8992 (N_8992,N_7601,N_7759);
or U8993 (N_8993,N_7476,N_7970);
or U8994 (N_8994,N_7969,N_7624);
or U8995 (N_8995,N_7503,N_7780);
and U8996 (N_8996,N_7086,N_7861);
xnor U8997 (N_8997,N_7111,N_7206);
xnor U8998 (N_8998,N_7486,N_7741);
and U8999 (N_8999,N_7070,N_7487);
nand U9000 (N_9000,N_8597,N_8116);
xnor U9001 (N_9001,N_8888,N_8881);
or U9002 (N_9002,N_8882,N_8914);
xnor U9003 (N_9003,N_8331,N_8978);
xor U9004 (N_9004,N_8101,N_8968);
nand U9005 (N_9005,N_8863,N_8641);
xnor U9006 (N_9006,N_8056,N_8012);
or U9007 (N_9007,N_8994,N_8281);
xor U9008 (N_9008,N_8538,N_8670);
nand U9009 (N_9009,N_8645,N_8232);
and U9010 (N_9010,N_8296,N_8775);
and U9011 (N_9011,N_8284,N_8586);
or U9012 (N_9012,N_8457,N_8467);
and U9013 (N_9013,N_8529,N_8515);
or U9014 (N_9014,N_8769,N_8736);
nor U9015 (N_9015,N_8040,N_8032);
nand U9016 (N_9016,N_8157,N_8916);
or U9017 (N_9017,N_8452,N_8193);
xnor U9018 (N_9018,N_8733,N_8025);
and U9019 (N_9019,N_8265,N_8253);
xnor U9020 (N_9020,N_8725,N_8398);
nor U9021 (N_9021,N_8128,N_8635);
or U9022 (N_9022,N_8320,N_8828);
nand U9023 (N_9023,N_8010,N_8346);
xnor U9024 (N_9024,N_8506,N_8058);
or U9025 (N_9025,N_8435,N_8434);
and U9026 (N_9026,N_8546,N_8239);
nand U9027 (N_9027,N_8716,N_8865);
or U9028 (N_9028,N_8471,N_8577);
xor U9029 (N_9029,N_8785,N_8276);
nor U9030 (N_9030,N_8352,N_8942);
nor U9031 (N_9031,N_8723,N_8222);
nand U9032 (N_9032,N_8464,N_8244);
and U9033 (N_9033,N_8403,N_8172);
nor U9034 (N_9034,N_8406,N_8849);
nor U9035 (N_9035,N_8424,N_8742);
nor U9036 (N_9036,N_8724,N_8963);
and U9037 (N_9037,N_8607,N_8988);
and U9038 (N_9038,N_8905,N_8463);
and U9039 (N_9039,N_8788,N_8563);
and U9040 (N_9040,N_8878,N_8475);
and U9041 (N_9041,N_8686,N_8497);
nor U9042 (N_9042,N_8708,N_8349);
nor U9043 (N_9043,N_8521,N_8480);
or U9044 (N_9044,N_8114,N_8687);
nand U9045 (N_9045,N_8117,N_8889);
or U9046 (N_9046,N_8306,N_8353);
or U9047 (N_9047,N_8336,N_8564);
nand U9048 (N_9048,N_8808,N_8718);
xor U9049 (N_9049,N_8523,N_8519);
nor U9050 (N_9050,N_8400,N_8451);
or U9051 (N_9051,N_8355,N_8273);
or U9052 (N_9052,N_8777,N_8109);
and U9053 (N_9053,N_8933,N_8877);
or U9054 (N_9054,N_8998,N_8572);
nor U9055 (N_9055,N_8612,N_8062);
xor U9056 (N_9056,N_8105,N_8308);
nor U9057 (N_9057,N_8841,N_8805);
or U9058 (N_9058,N_8057,N_8330);
nor U9059 (N_9059,N_8162,N_8498);
or U9060 (N_9060,N_8035,N_8674);
nand U9061 (N_9061,N_8195,N_8554);
and U9062 (N_9062,N_8247,N_8111);
xnor U9063 (N_9063,N_8477,N_8379);
or U9064 (N_9064,N_8932,N_8217);
and U9065 (N_9065,N_8199,N_8999);
nand U9066 (N_9066,N_8527,N_8350);
nor U9067 (N_9067,N_8892,N_8219);
nand U9068 (N_9068,N_8649,N_8149);
nand U9069 (N_9069,N_8496,N_8950);
nand U9070 (N_9070,N_8692,N_8082);
and U9071 (N_9071,N_8928,N_8132);
nand U9072 (N_9072,N_8059,N_8587);
nor U9073 (N_9073,N_8404,N_8447);
or U9074 (N_9074,N_8163,N_8616);
or U9075 (N_9075,N_8039,N_8268);
and U9076 (N_9076,N_8569,N_8160);
and U9077 (N_9077,N_8154,N_8227);
nand U9078 (N_9078,N_8773,N_8593);
nor U9079 (N_9079,N_8858,N_8634);
nor U9080 (N_9080,N_8924,N_8257);
nor U9081 (N_9081,N_8310,N_8432);
nand U9082 (N_9082,N_8324,N_8259);
xnor U9083 (N_9083,N_8526,N_8995);
nand U9084 (N_9084,N_8976,N_8539);
nor U9085 (N_9085,N_8312,N_8703);
nor U9086 (N_9086,N_8840,N_8588);
and U9087 (N_9087,N_8817,N_8422);
nand U9088 (N_9088,N_8120,N_8943);
nor U9089 (N_9089,N_8748,N_8411);
or U9090 (N_9090,N_8390,N_8771);
nor U9091 (N_9091,N_8606,N_8739);
or U9092 (N_9092,N_8644,N_8333);
nor U9093 (N_9093,N_8959,N_8694);
or U9094 (N_9094,N_8318,N_8251);
nor U9095 (N_9095,N_8602,N_8412);
xor U9096 (N_9096,N_8441,N_8671);
and U9097 (N_9097,N_8949,N_8740);
nand U9098 (N_9098,N_8679,N_8704);
or U9099 (N_9099,N_8042,N_8054);
or U9100 (N_9100,N_8706,N_8046);
and U9101 (N_9101,N_8283,N_8946);
nor U9102 (N_9102,N_8125,N_8070);
and U9103 (N_9103,N_8798,N_8936);
or U9104 (N_9104,N_8838,N_8302);
nand U9105 (N_9105,N_8601,N_8233);
nand U9106 (N_9106,N_8776,N_8384);
nor U9107 (N_9107,N_8014,N_8800);
nor U9108 (N_9108,N_8181,N_8734);
and U9109 (N_9109,N_8919,N_8534);
nand U9110 (N_9110,N_8866,N_8565);
xor U9111 (N_9111,N_8381,N_8166);
nand U9112 (N_9112,N_8600,N_8632);
nor U9113 (N_9113,N_8875,N_8960);
nor U9114 (N_9114,N_8030,N_8009);
nor U9115 (N_9115,N_8551,N_8864);
nor U9116 (N_9116,N_8927,N_8610);
nor U9117 (N_9117,N_8338,N_8490);
or U9118 (N_9118,N_8374,N_8853);
and U9119 (N_9119,N_8126,N_8397);
or U9120 (N_9120,N_8002,N_8666);
nand U9121 (N_9121,N_8423,N_8510);
or U9122 (N_9122,N_8985,N_8197);
nand U9123 (N_9123,N_8474,N_8814);
xor U9124 (N_9124,N_8396,N_8782);
nor U9125 (N_9125,N_8886,N_8375);
and U9126 (N_9126,N_8815,N_8392);
nor U9127 (N_9127,N_8084,N_8683);
nor U9128 (N_9128,N_8696,N_8494);
nand U9129 (N_9129,N_8297,N_8603);
nor U9130 (N_9130,N_8034,N_8504);
nand U9131 (N_9131,N_8596,N_8891);
nor U9132 (N_9132,N_8314,N_8509);
or U9133 (N_9133,N_8263,N_8107);
nor U9134 (N_9134,N_8688,N_8407);
or U9135 (N_9135,N_8874,N_8461);
nor U9136 (N_9136,N_8388,N_8582);
or U9137 (N_9137,N_8419,N_8678);
nand U9138 (N_9138,N_8071,N_8409);
nand U9139 (N_9139,N_8174,N_8394);
xor U9140 (N_9140,N_8221,N_8448);
nor U9141 (N_9141,N_8072,N_8726);
xnor U9142 (N_9142,N_8668,N_8345);
or U9143 (N_9143,N_8656,N_8469);
or U9144 (N_9144,N_8052,N_8953);
nor U9145 (N_9145,N_8341,N_8140);
xor U9146 (N_9146,N_8541,N_8291);
xnor U9147 (N_9147,N_8011,N_8759);
xor U9148 (N_9148,N_8021,N_8013);
nand U9149 (N_9149,N_8608,N_8340);
nor U9150 (N_9150,N_8847,N_8611);
xnor U9151 (N_9151,N_8536,N_8727);
and U9152 (N_9152,N_8460,N_8488);
nand U9153 (N_9153,N_8544,N_8767);
or U9154 (N_9154,N_8661,N_8236);
nand U9155 (N_9155,N_8486,N_8074);
nor U9156 (N_9156,N_8749,N_8789);
or U9157 (N_9157,N_8286,N_8904);
nor U9158 (N_9158,N_8614,N_8391);
or U9159 (N_9159,N_8364,N_8231);
nor U9160 (N_9160,N_8556,N_8366);
and U9161 (N_9161,N_8387,N_8295);
nand U9162 (N_9162,N_8050,N_8619);
nand U9163 (N_9163,N_8848,N_8780);
xor U9164 (N_9164,N_8750,N_8473);
xnor U9165 (N_9165,N_8737,N_8643);
nor U9166 (N_9166,N_8762,N_8027);
nand U9167 (N_9167,N_8557,N_8684);
xor U9168 (N_9168,N_8026,N_8561);
and U9169 (N_9169,N_8187,N_8356);
or U9170 (N_9170,N_8063,N_8633);
or U9171 (N_9171,N_8520,N_8981);
xnor U9172 (N_9172,N_8278,N_8761);
nand U9173 (N_9173,N_8907,N_8260);
nor U9174 (N_9174,N_8478,N_8136);
or U9175 (N_9175,N_8745,N_8549);
or U9176 (N_9176,N_8617,N_8148);
or U9177 (N_9177,N_8813,N_8533);
or U9178 (N_9178,N_8972,N_8547);
xor U9179 (N_9179,N_8605,N_8906);
nor U9180 (N_9180,N_8592,N_8680);
xnor U9181 (N_9181,N_8279,N_8839);
xor U9182 (N_9182,N_8676,N_8855);
nand U9183 (N_9183,N_8426,N_8990);
or U9184 (N_9184,N_8235,N_8370);
nand U9185 (N_9185,N_8573,N_8272);
nor U9186 (N_9186,N_8941,N_8418);
or U9187 (N_9187,N_8112,N_8049);
or U9188 (N_9188,N_8885,N_8883);
and U9189 (N_9189,N_8127,N_8872);
or U9190 (N_9190,N_8413,N_8266);
nand U9191 (N_9191,N_8535,N_8873);
nand U9192 (N_9192,N_8884,N_8303);
xor U9193 (N_9193,N_8378,N_8137);
and U9194 (N_9194,N_8944,N_8442);
nand U9195 (N_9195,N_8399,N_8316);
nand U9196 (N_9196,N_8216,N_8335);
nor U9197 (N_9197,N_8568,N_8827);
or U9198 (N_9198,N_8122,N_8167);
nor U9199 (N_9199,N_8246,N_8772);
nor U9200 (N_9200,N_8648,N_8362);
xor U9201 (N_9201,N_8690,N_8096);
nand U9202 (N_9202,N_8934,N_8439);
nor U9203 (N_9203,N_8465,N_8756);
and U9204 (N_9204,N_8479,N_8323);
or U9205 (N_9205,N_8925,N_8626);
xnor U9206 (N_9206,N_8138,N_8511);
or U9207 (N_9207,N_8862,N_8859);
nand U9208 (N_9208,N_8093,N_8031);
nor U9209 (N_9209,N_8518,N_8240);
or U9210 (N_9210,N_8019,N_8898);
nand U9211 (N_9211,N_8225,N_8755);
nand U9212 (N_9212,N_8850,N_8468);
nand U9213 (N_9213,N_8639,N_8792);
nand U9214 (N_9214,N_8646,N_8747);
xnor U9215 (N_9215,N_8351,N_8214);
and U9216 (N_9216,N_8015,N_8757);
and U9217 (N_9217,N_8191,N_8092);
and U9218 (N_9218,N_8090,N_8657);
nor U9219 (N_9219,N_8682,N_8957);
and U9220 (N_9220,N_8438,N_8810);
xnor U9221 (N_9221,N_8437,N_8067);
and U9222 (N_9222,N_8583,N_8020);
nand U9223 (N_9223,N_8023,N_8570);
xnor U9224 (N_9224,N_8237,N_8408);
and U9225 (N_9225,N_8337,N_8580);
or U9226 (N_9226,N_8961,N_8833);
and U9227 (N_9227,N_8970,N_8594);
and U9228 (N_9228,N_8146,N_8618);
nor U9229 (N_9229,N_8028,N_8826);
nand U9230 (N_9230,N_8121,N_8098);
nor U9231 (N_9231,N_8425,N_8326);
and U9232 (N_9232,N_8879,N_8334);
or U9233 (N_9233,N_8818,N_8202);
nand U9234 (N_9234,N_8287,N_8578);
and U9235 (N_9235,N_8223,N_8017);
xor U9236 (N_9236,N_8804,N_8992);
or U9237 (N_9237,N_8512,N_8047);
nand U9238 (N_9238,N_8178,N_8053);
xor U9239 (N_9239,N_8207,N_8753);
nor U9240 (N_9240,N_8304,N_8104);
and U9241 (N_9241,N_8282,N_8651);
and U9242 (N_9242,N_8454,N_8410);
and U9243 (N_9243,N_8201,N_8728);
and U9244 (N_9244,N_8175,N_8076);
nand U9245 (N_9245,N_8658,N_8713);
nor U9246 (N_9246,N_8524,N_8576);
nor U9247 (N_9247,N_8363,N_8143);
nand U9248 (N_9248,N_8389,N_8667);
xor U9249 (N_9249,N_8779,N_8103);
nor U9250 (N_9250,N_8443,N_8190);
xnor U9251 (N_9251,N_8675,N_8514);
nand U9252 (N_9252,N_8760,N_8170);
and U9253 (N_9253,N_8880,N_8507);
nand U9254 (N_9254,N_8361,N_8824);
or U9255 (N_9255,N_8669,N_8856);
nor U9256 (N_9256,N_8313,N_8198);
nand U9257 (N_9257,N_8095,N_8086);
nor U9258 (N_9258,N_8079,N_8794);
or U9259 (N_9259,N_8061,N_8595);
and U9260 (N_9260,N_8258,N_8188);
nor U9261 (N_9261,N_8842,N_8134);
and U9262 (N_9262,N_8663,N_8900);
nand U9263 (N_9263,N_8077,N_8940);
nor U9264 (N_9264,N_8209,N_8652);
nand U9265 (N_9265,N_8180,N_8182);
nor U9266 (N_9266,N_8129,N_8380);
and U9267 (N_9267,N_8806,N_8786);
or U9268 (N_9268,N_8517,N_8493);
xor U9269 (N_9269,N_8693,N_8368);
nor U9270 (N_9270,N_8908,N_8930);
nand U9271 (N_9271,N_8861,N_8764);
nor U9272 (N_9272,N_8964,N_8912);
nor U9273 (N_9273,N_8405,N_8360);
nor U9274 (N_9274,N_8901,N_8401);
nand U9275 (N_9275,N_8395,N_8234);
or U9276 (N_9276,N_8613,N_8532);
xor U9277 (N_9277,N_8954,N_8068);
nor U9278 (N_9278,N_8489,N_8110);
nand U9279 (N_9279,N_8205,N_8483);
nor U9280 (N_9280,N_8774,N_8359);
and U9281 (N_9281,N_8189,N_8701);
or U9282 (N_9282,N_8069,N_8948);
nor U9283 (N_9283,N_8041,N_8719);
or U9284 (N_9284,N_8289,N_8887);
and U9285 (N_9285,N_8829,N_8659);
or U9286 (N_9286,N_8044,N_8746);
nand U9287 (N_9287,N_8825,N_8311);
xnor U9288 (N_9288,N_8835,N_8037);
xor U9289 (N_9289,N_8270,N_8073);
nor U9290 (N_9290,N_8436,N_8846);
or U9291 (N_9291,N_8735,N_8008);
nor U9292 (N_9292,N_8973,N_8870);
nand U9293 (N_9293,N_8857,N_8935);
nand U9294 (N_9294,N_8275,N_8256);
xor U9295 (N_9295,N_8629,N_8552);
nand U9296 (N_9296,N_8081,N_8444);
or U9297 (N_9297,N_8382,N_8620);
and U9298 (N_9298,N_8809,N_8357);
xor U9299 (N_9299,N_8791,N_8385);
or U9300 (N_9300,N_8665,N_8038);
nand U9301 (N_9301,N_8043,N_8902);
nor U9302 (N_9302,N_8503,N_8383);
xnor U9303 (N_9303,N_8758,N_8894);
nor U9304 (N_9304,N_8705,N_8540);
nor U9305 (N_9305,N_8300,N_8910);
and U9306 (N_9306,N_8691,N_8342);
xor U9307 (N_9307,N_8156,N_8522);
nand U9308 (N_9308,N_8989,N_8230);
or U9309 (N_9309,N_8937,N_8969);
nor U9310 (N_9310,N_8714,N_8599);
xnor U9311 (N_9311,N_8173,N_8179);
and U9312 (N_9312,N_8249,N_8458);
xnor U9313 (N_9313,N_8135,N_8784);
and U9314 (N_9314,N_8897,N_8367);
xor U9315 (N_9315,N_8650,N_8393);
or U9316 (N_9316,N_8144,N_8636);
or U9317 (N_9317,N_8196,N_8820);
nor U9318 (N_9318,N_8429,N_8783);
xnor U9319 (N_9319,N_8164,N_8832);
or U9320 (N_9320,N_8702,N_8006);
or U9321 (N_9321,N_8150,N_8358);
or U9322 (N_9322,N_8171,N_8860);
nor U9323 (N_9323,N_8446,N_8051);
and U9324 (N_9324,N_8699,N_8631);
xnor U9325 (N_9325,N_8274,N_8709);
or U9326 (N_9326,N_8184,N_8427);
and U9327 (N_9327,N_8194,N_8416);
xor U9328 (N_9328,N_8048,N_8955);
or U9329 (N_9329,N_8720,N_8248);
nand U9330 (N_9330,N_8119,N_8501);
or U9331 (N_9331,N_8781,N_8321);
xnor U9332 (N_9332,N_8807,N_8801);
nor U9333 (N_9333,N_8796,N_8655);
and U9334 (N_9334,N_8654,N_8770);
nand U9335 (N_9335,N_8224,N_8348);
or U9336 (N_9336,N_8915,N_8001);
and U9337 (N_9337,N_8124,N_8575);
and U9338 (N_9338,N_8951,N_8036);
or U9339 (N_9339,N_8228,N_8911);
nor U9340 (N_9340,N_8339,N_8567);
or U9341 (N_9341,N_8307,N_8868);
nand U9342 (N_9342,N_8371,N_8495);
or U9343 (N_9343,N_8545,N_8064);
and U9344 (N_9344,N_8876,N_8492);
and U9345 (N_9345,N_8269,N_8029);
nand U9346 (N_9346,N_8530,N_8243);
nand U9347 (N_9347,N_8799,N_8751);
and U9348 (N_9348,N_8369,N_8168);
nor U9349 (N_9349,N_8087,N_8695);
xor U9350 (N_9350,N_8455,N_8242);
or U9351 (N_9351,N_8255,N_8123);
nor U9352 (N_9352,N_8731,N_8212);
or U9353 (N_9353,N_8476,N_8491);
nand U9354 (N_9354,N_8262,N_8290);
nand U9355 (N_9355,N_8766,N_8823);
nor U9356 (N_9356,N_8177,N_8505);
and U9357 (N_9357,N_8500,N_8280);
nor U9358 (N_9358,N_8373,N_8045);
xnor U9359 (N_9359,N_8811,N_8627);
or U9360 (N_9360,N_8765,N_8956);
xor U9361 (N_9361,N_8837,N_8797);
xor U9362 (N_9362,N_8787,N_8113);
or U9363 (N_9363,N_8637,N_8200);
nor U9364 (N_9364,N_8845,N_8895);
or U9365 (N_9365,N_8974,N_8738);
and U9366 (N_9366,N_8965,N_8975);
nor U9367 (N_9367,N_8292,N_8803);
or U9368 (N_9368,N_8790,N_8741);
or U9369 (N_9369,N_8579,N_8918);
or U9370 (N_9370,N_8621,N_8947);
xnor U9371 (N_9371,N_8664,N_8913);
and U9372 (N_9372,N_8288,N_8834);
nor U9373 (N_9373,N_8867,N_8450);
xnor U9374 (N_9374,N_8075,N_8005);
nand U9375 (N_9375,N_8007,N_8903);
nor U9376 (N_9376,N_8241,N_8971);
or U9377 (N_9377,N_8459,N_8590);
or U9378 (N_9378,N_8097,N_8083);
nand U9379 (N_9379,N_8977,N_8309);
nor U9380 (N_9380,N_8929,N_8327);
nor U9381 (N_9381,N_8332,N_8712);
nand U9382 (N_9382,N_8264,N_8322);
and U9383 (N_9383,N_8206,N_8922);
and U9384 (N_9384,N_8100,N_8151);
nand U9385 (N_9385,N_8183,N_8991);
nand U9386 (N_9386,N_8250,N_8261);
xor U9387 (N_9387,N_8625,N_8923);
and U9388 (N_9388,N_8299,N_8528);
nand U9389 (N_9389,N_8768,N_8711);
xor U9390 (N_9390,N_8513,N_8537);
and U9391 (N_9391,N_8294,N_8743);
xnor U9392 (N_9392,N_8598,N_8722);
or U9393 (N_9393,N_8899,N_8213);
or U9394 (N_9394,N_8979,N_8099);
nor U9395 (N_9395,N_8729,N_8836);
or U9396 (N_9396,N_8980,N_8984);
nand U9397 (N_9397,N_8710,N_8317);
or U9398 (N_9398,N_8996,N_8456);
xnor U9399 (N_9399,N_8343,N_8548);
or U9400 (N_9400,N_8591,N_8372);
nor U9401 (N_9401,N_8319,N_8660);
xnor U9402 (N_9402,N_8793,N_8831);
and U9403 (N_9403,N_8016,N_8543);
nand U9404 (N_9404,N_8508,N_8153);
or U9405 (N_9405,N_8571,N_8516);
nor U9406 (N_9406,N_8133,N_8344);
or U9407 (N_9407,N_8685,N_8161);
and U9408 (N_9408,N_8589,N_8466);
and U9409 (N_9409,N_8677,N_8673);
nand U9410 (N_9410,N_8604,N_8893);
or U9411 (N_9411,N_8420,N_8108);
nand U9412 (N_9412,N_8821,N_8707);
xnor U9413 (N_9413,N_8118,N_8445);
nand U9414 (N_9414,N_8802,N_8615);
xor U9415 (N_9415,N_8698,N_8531);
and U9416 (N_9416,N_8271,N_8700);
xor U9417 (N_9417,N_8485,N_8525);
nand U9418 (N_9418,N_8653,N_8089);
nor U9419 (N_9419,N_8869,N_8624);
or U9420 (N_9420,N_8566,N_8204);
nand U9421 (N_9421,N_8159,N_8414);
or U9422 (N_9422,N_8628,N_8697);
or U9423 (N_9423,N_8890,N_8816);
or U9424 (N_9424,N_8022,N_8623);
nor U9425 (N_9425,N_8462,N_8744);
or U9426 (N_9426,N_8871,N_8328);
nand U9427 (N_9427,N_8453,N_8945);
nor U9428 (N_9428,N_8581,N_8920);
and U9429 (N_9429,N_8000,N_8630);
nand U9430 (N_9430,N_8142,N_8078);
and U9431 (N_9431,N_8732,N_8415);
and U9432 (N_9432,N_8066,N_8210);
nor U9433 (N_9433,N_8830,N_8553);
and U9434 (N_9434,N_8487,N_8962);
and U9435 (N_9435,N_8376,N_8647);
xnor U9436 (N_9436,N_8430,N_8851);
xor U9437 (N_9437,N_8131,N_8305);
xnor U9438 (N_9438,N_8421,N_8254);
nor U9439 (N_9439,N_8795,N_8208);
nor U9440 (N_9440,N_8844,N_8102);
or U9441 (N_9441,N_8939,N_8386);
nor U9442 (N_9442,N_8130,N_8428);
nor U9443 (N_9443,N_8298,N_8347);
nor U9444 (N_9444,N_8169,N_8285);
nor U9445 (N_9445,N_8754,N_8293);
and U9446 (N_9446,N_8987,N_8003);
or U9447 (N_9447,N_8185,N_8717);
nor U9448 (N_9448,N_8560,N_8917);
and U9449 (N_9449,N_8843,N_8481);
or U9450 (N_9450,N_8721,N_8417);
or U9451 (N_9451,N_8354,N_8176);
nand U9452 (N_9452,N_8672,N_8609);
and U9453 (N_9453,N_8449,N_8267);
or U9454 (N_9454,N_8730,N_8926);
or U9455 (N_9455,N_8115,N_8165);
nor U9456 (N_9456,N_8931,N_8763);
nor U9457 (N_9457,N_8574,N_8085);
nand U9458 (N_9458,N_8640,N_8986);
nand U9459 (N_9459,N_8715,N_8018);
and U9460 (N_9460,N_8982,N_8229);
and U9461 (N_9461,N_8689,N_8472);
nand U9462 (N_9462,N_8004,N_8080);
nor U9463 (N_9463,N_8315,N_8088);
or U9464 (N_9464,N_8301,N_8226);
xnor U9465 (N_9465,N_8203,N_8220);
and U9466 (N_9466,N_8211,N_8502);
xor U9467 (N_9467,N_8215,N_8139);
nand U9468 (N_9468,N_8681,N_8440);
and U9469 (N_9469,N_8060,N_8622);
nor U9470 (N_9470,N_8967,N_8952);
or U9471 (N_9471,N_8277,N_8033);
nor U9472 (N_9472,N_8218,N_8245);
xnor U9473 (N_9473,N_8812,N_8186);
xnor U9474 (N_9474,N_8854,N_8550);
and U9475 (N_9475,N_8482,N_8152);
nor U9476 (N_9476,N_8819,N_8147);
or U9477 (N_9477,N_8433,N_8106);
nor U9478 (N_9478,N_8938,N_8141);
xor U9479 (N_9479,N_8094,N_8993);
or U9480 (N_9480,N_8997,N_8752);
nand U9481 (N_9481,N_8921,N_8559);
and U9482 (N_9482,N_8958,N_8192);
or U9483 (N_9483,N_8558,N_8966);
and U9484 (N_9484,N_8562,N_8155);
nand U9485 (N_9485,N_8402,N_8065);
and U9486 (N_9486,N_8024,N_8091);
xor U9487 (N_9487,N_8377,N_8555);
nor U9488 (N_9488,N_8238,N_8584);
nor U9489 (N_9489,N_8158,N_8896);
nand U9490 (N_9490,N_8470,N_8778);
nand U9491 (N_9491,N_8431,N_8329);
or U9492 (N_9492,N_8252,N_8585);
xor U9493 (N_9493,N_8484,N_8365);
and U9494 (N_9494,N_8055,N_8852);
xnor U9495 (N_9495,N_8325,N_8822);
or U9496 (N_9496,N_8983,N_8909);
nor U9497 (N_9497,N_8642,N_8638);
or U9498 (N_9498,N_8662,N_8499);
nor U9499 (N_9499,N_8145,N_8542);
or U9500 (N_9500,N_8968,N_8230);
nor U9501 (N_9501,N_8655,N_8666);
and U9502 (N_9502,N_8683,N_8821);
xnor U9503 (N_9503,N_8600,N_8909);
xor U9504 (N_9504,N_8974,N_8613);
or U9505 (N_9505,N_8797,N_8706);
or U9506 (N_9506,N_8377,N_8994);
nor U9507 (N_9507,N_8917,N_8987);
nand U9508 (N_9508,N_8772,N_8704);
or U9509 (N_9509,N_8725,N_8652);
nand U9510 (N_9510,N_8336,N_8107);
or U9511 (N_9511,N_8592,N_8001);
nand U9512 (N_9512,N_8229,N_8100);
nand U9513 (N_9513,N_8678,N_8384);
or U9514 (N_9514,N_8466,N_8077);
and U9515 (N_9515,N_8518,N_8855);
nand U9516 (N_9516,N_8919,N_8922);
nor U9517 (N_9517,N_8038,N_8269);
nand U9518 (N_9518,N_8397,N_8823);
nor U9519 (N_9519,N_8963,N_8055);
nor U9520 (N_9520,N_8113,N_8488);
nor U9521 (N_9521,N_8973,N_8552);
or U9522 (N_9522,N_8634,N_8317);
nor U9523 (N_9523,N_8609,N_8502);
xor U9524 (N_9524,N_8209,N_8264);
nand U9525 (N_9525,N_8449,N_8140);
and U9526 (N_9526,N_8019,N_8581);
and U9527 (N_9527,N_8111,N_8115);
and U9528 (N_9528,N_8160,N_8429);
and U9529 (N_9529,N_8053,N_8800);
and U9530 (N_9530,N_8152,N_8192);
and U9531 (N_9531,N_8310,N_8087);
xnor U9532 (N_9532,N_8689,N_8644);
or U9533 (N_9533,N_8264,N_8481);
nor U9534 (N_9534,N_8167,N_8144);
and U9535 (N_9535,N_8310,N_8142);
nor U9536 (N_9536,N_8196,N_8345);
and U9537 (N_9537,N_8229,N_8546);
or U9538 (N_9538,N_8060,N_8373);
or U9539 (N_9539,N_8337,N_8359);
or U9540 (N_9540,N_8142,N_8627);
nand U9541 (N_9541,N_8354,N_8131);
nor U9542 (N_9542,N_8312,N_8908);
nor U9543 (N_9543,N_8043,N_8255);
nor U9544 (N_9544,N_8531,N_8721);
or U9545 (N_9545,N_8288,N_8171);
xnor U9546 (N_9546,N_8038,N_8580);
xnor U9547 (N_9547,N_8454,N_8950);
and U9548 (N_9548,N_8750,N_8822);
or U9549 (N_9549,N_8218,N_8605);
xnor U9550 (N_9550,N_8529,N_8633);
and U9551 (N_9551,N_8769,N_8084);
nand U9552 (N_9552,N_8473,N_8106);
nand U9553 (N_9553,N_8162,N_8047);
xor U9554 (N_9554,N_8992,N_8251);
or U9555 (N_9555,N_8322,N_8752);
and U9556 (N_9556,N_8074,N_8304);
nor U9557 (N_9557,N_8237,N_8630);
nand U9558 (N_9558,N_8271,N_8069);
or U9559 (N_9559,N_8096,N_8098);
or U9560 (N_9560,N_8794,N_8127);
nand U9561 (N_9561,N_8772,N_8558);
and U9562 (N_9562,N_8717,N_8125);
or U9563 (N_9563,N_8322,N_8123);
and U9564 (N_9564,N_8636,N_8025);
nand U9565 (N_9565,N_8677,N_8139);
nor U9566 (N_9566,N_8183,N_8313);
and U9567 (N_9567,N_8331,N_8334);
and U9568 (N_9568,N_8402,N_8070);
nor U9569 (N_9569,N_8834,N_8845);
and U9570 (N_9570,N_8290,N_8199);
and U9571 (N_9571,N_8518,N_8398);
xor U9572 (N_9572,N_8178,N_8663);
nand U9573 (N_9573,N_8541,N_8951);
and U9574 (N_9574,N_8523,N_8115);
nand U9575 (N_9575,N_8500,N_8916);
nor U9576 (N_9576,N_8479,N_8541);
or U9577 (N_9577,N_8258,N_8666);
nand U9578 (N_9578,N_8809,N_8558);
nor U9579 (N_9579,N_8670,N_8170);
or U9580 (N_9580,N_8191,N_8323);
nand U9581 (N_9581,N_8741,N_8280);
or U9582 (N_9582,N_8188,N_8356);
and U9583 (N_9583,N_8520,N_8006);
nor U9584 (N_9584,N_8235,N_8926);
nand U9585 (N_9585,N_8781,N_8583);
xnor U9586 (N_9586,N_8016,N_8897);
or U9587 (N_9587,N_8970,N_8451);
nor U9588 (N_9588,N_8997,N_8849);
xnor U9589 (N_9589,N_8343,N_8563);
xor U9590 (N_9590,N_8434,N_8937);
and U9591 (N_9591,N_8680,N_8917);
xor U9592 (N_9592,N_8527,N_8316);
nand U9593 (N_9593,N_8879,N_8312);
nand U9594 (N_9594,N_8245,N_8870);
or U9595 (N_9595,N_8038,N_8920);
xnor U9596 (N_9596,N_8358,N_8760);
or U9597 (N_9597,N_8671,N_8353);
xnor U9598 (N_9598,N_8930,N_8915);
nand U9599 (N_9599,N_8711,N_8949);
and U9600 (N_9600,N_8939,N_8911);
nor U9601 (N_9601,N_8733,N_8481);
xor U9602 (N_9602,N_8310,N_8459);
nand U9603 (N_9603,N_8155,N_8373);
and U9604 (N_9604,N_8098,N_8888);
nor U9605 (N_9605,N_8021,N_8215);
xor U9606 (N_9606,N_8255,N_8789);
xor U9607 (N_9607,N_8637,N_8449);
or U9608 (N_9608,N_8330,N_8753);
or U9609 (N_9609,N_8059,N_8001);
and U9610 (N_9610,N_8587,N_8248);
xnor U9611 (N_9611,N_8354,N_8274);
nor U9612 (N_9612,N_8500,N_8785);
or U9613 (N_9613,N_8285,N_8489);
and U9614 (N_9614,N_8746,N_8472);
nand U9615 (N_9615,N_8730,N_8201);
or U9616 (N_9616,N_8350,N_8522);
nand U9617 (N_9617,N_8590,N_8653);
nor U9618 (N_9618,N_8223,N_8529);
nand U9619 (N_9619,N_8934,N_8869);
or U9620 (N_9620,N_8410,N_8022);
or U9621 (N_9621,N_8171,N_8961);
nor U9622 (N_9622,N_8155,N_8463);
xnor U9623 (N_9623,N_8527,N_8355);
nor U9624 (N_9624,N_8824,N_8136);
nand U9625 (N_9625,N_8612,N_8572);
xor U9626 (N_9626,N_8403,N_8241);
nand U9627 (N_9627,N_8534,N_8805);
or U9628 (N_9628,N_8473,N_8807);
and U9629 (N_9629,N_8566,N_8705);
and U9630 (N_9630,N_8694,N_8999);
or U9631 (N_9631,N_8493,N_8196);
xnor U9632 (N_9632,N_8206,N_8066);
nand U9633 (N_9633,N_8220,N_8381);
or U9634 (N_9634,N_8686,N_8182);
and U9635 (N_9635,N_8313,N_8778);
xnor U9636 (N_9636,N_8974,N_8233);
and U9637 (N_9637,N_8202,N_8875);
xor U9638 (N_9638,N_8620,N_8163);
nand U9639 (N_9639,N_8622,N_8912);
xor U9640 (N_9640,N_8170,N_8498);
xnor U9641 (N_9641,N_8768,N_8098);
and U9642 (N_9642,N_8263,N_8406);
or U9643 (N_9643,N_8195,N_8258);
nand U9644 (N_9644,N_8982,N_8193);
nor U9645 (N_9645,N_8337,N_8216);
or U9646 (N_9646,N_8960,N_8982);
or U9647 (N_9647,N_8690,N_8598);
and U9648 (N_9648,N_8801,N_8438);
nand U9649 (N_9649,N_8815,N_8301);
and U9650 (N_9650,N_8842,N_8574);
nand U9651 (N_9651,N_8392,N_8659);
or U9652 (N_9652,N_8362,N_8695);
and U9653 (N_9653,N_8049,N_8819);
xor U9654 (N_9654,N_8862,N_8412);
xnor U9655 (N_9655,N_8478,N_8119);
xor U9656 (N_9656,N_8211,N_8729);
or U9657 (N_9657,N_8484,N_8125);
xor U9658 (N_9658,N_8014,N_8154);
and U9659 (N_9659,N_8264,N_8821);
or U9660 (N_9660,N_8130,N_8802);
nand U9661 (N_9661,N_8228,N_8746);
and U9662 (N_9662,N_8369,N_8150);
nor U9663 (N_9663,N_8940,N_8311);
or U9664 (N_9664,N_8739,N_8189);
nor U9665 (N_9665,N_8999,N_8405);
nand U9666 (N_9666,N_8765,N_8238);
or U9667 (N_9667,N_8279,N_8201);
nand U9668 (N_9668,N_8912,N_8055);
or U9669 (N_9669,N_8421,N_8075);
or U9670 (N_9670,N_8709,N_8409);
nand U9671 (N_9671,N_8241,N_8565);
and U9672 (N_9672,N_8982,N_8426);
or U9673 (N_9673,N_8643,N_8499);
nand U9674 (N_9674,N_8080,N_8961);
xor U9675 (N_9675,N_8096,N_8612);
nor U9676 (N_9676,N_8682,N_8409);
xor U9677 (N_9677,N_8273,N_8263);
xor U9678 (N_9678,N_8484,N_8811);
nor U9679 (N_9679,N_8434,N_8899);
xnor U9680 (N_9680,N_8935,N_8601);
xnor U9681 (N_9681,N_8810,N_8652);
nor U9682 (N_9682,N_8340,N_8417);
xnor U9683 (N_9683,N_8681,N_8530);
nor U9684 (N_9684,N_8322,N_8345);
nor U9685 (N_9685,N_8751,N_8126);
or U9686 (N_9686,N_8454,N_8134);
nand U9687 (N_9687,N_8730,N_8831);
or U9688 (N_9688,N_8962,N_8374);
xnor U9689 (N_9689,N_8937,N_8836);
or U9690 (N_9690,N_8788,N_8509);
xnor U9691 (N_9691,N_8199,N_8739);
or U9692 (N_9692,N_8802,N_8541);
or U9693 (N_9693,N_8529,N_8934);
and U9694 (N_9694,N_8166,N_8169);
nand U9695 (N_9695,N_8001,N_8753);
xor U9696 (N_9696,N_8897,N_8069);
nor U9697 (N_9697,N_8805,N_8654);
and U9698 (N_9698,N_8326,N_8714);
or U9699 (N_9699,N_8681,N_8032);
and U9700 (N_9700,N_8952,N_8931);
nor U9701 (N_9701,N_8981,N_8868);
nor U9702 (N_9702,N_8855,N_8239);
nand U9703 (N_9703,N_8385,N_8721);
nor U9704 (N_9704,N_8888,N_8736);
xor U9705 (N_9705,N_8439,N_8035);
xor U9706 (N_9706,N_8517,N_8782);
xnor U9707 (N_9707,N_8040,N_8330);
xnor U9708 (N_9708,N_8795,N_8180);
nor U9709 (N_9709,N_8018,N_8623);
xnor U9710 (N_9710,N_8386,N_8487);
nor U9711 (N_9711,N_8978,N_8933);
xnor U9712 (N_9712,N_8231,N_8978);
nor U9713 (N_9713,N_8099,N_8658);
nand U9714 (N_9714,N_8492,N_8085);
xnor U9715 (N_9715,N_8920,N_8982);
nand U9716 (N_9716,N_8986,N_8865);
nor U9717 (N_9717,N_8329,N_8081);
xnor U9718 (N_9718,N_8763,N_8648);
and U9719 (N_9719,N_8320,N_8707);
xnor U9720 (N_9720,N_8171,N_8202);
or U9721 (N_9721,N_8732,N_8850);
and U9722 (N_9722,N_8222,N_8918);
xor U9723 (N_9723,N_8467,N_8657);
xor U9724 (N_9724,N_8012,N_8457);
xor U9725 (N_9725,N_8291,N_8824);
xor U9726 (N_9726,N_8406,N_8028);
and U9727 (N_9727,N_8356,N_8746);
nor U9728 (N_9728,N_8747,N_8953);
or U9729 (N_9729,N_8095,N_8566);
xnor U9730 (N_9730,N_8671,N_8670);
nor U9731 (N_9731,N_8986,N_8743);
and U9732 (N_9732,N_8436,N_8088);
nor U9733 (N_9733,N_8680,N_8066);
nand U9734 (N_9734,N_8164,N_8245);
and U9735 (N_9735,N_8130,N_8736);
nand U9736 (N_9736,N_8275,N_8898);
nand U9737 (N_9737,N_8834,N_8521);
xnor U9738 (N_9738,N_8188,N_8995);
nor U9739 (N_9739,N_8353,N_8150);
and U9740 (N_9740,N_8055,N_8419);
xor U9741 (N_9741,N_8359,N_8737);
or U9742 (N_9742,N_8154,N_8348);
nand U9743 (N_9743,N_8743,N_8470);
or U9744 (N_9744,N_8793,N_8604);
or U9745 (N_9745,N_8112,N_8659);
xnor U9746 (N_9746,N_8057,N_8353);
or U9747 (N_9747,N_8836,N_8317);
nand U9748 (N_9748,N_8052,N_8288);
xor U9749 (N_9749,N_8740,N_8898);
and U9750 (N_9750,N_8834,N_8626);
nand U9751 (N_9751,N_8895,N_8165);
or U9752 (N_9752,N_8313,N_8363);
or U9753 (N_9753,N_8943,N_8661);
nor U9754 (N_9754,N_8303,N_8136);
or U9755 (N_9755,N_8608,N_8288);
nor U9756 (N_9756,N_8447,N_8703);
nand U9757 (N_9757,N_8842,N_8744);
xnor U9758 (N_9758,N_8318,N_8966);
nand U9759 (N_9759,N_8519,N_8614);
xor U9760 (N_9760,N_8272,N_8889);
nor U9761 (N_9761,N_8553,N_8985);
nand U9762 (N_9762,N_8173,N_8608);
and U9763 (N_9763,N_8233,N_8704);
xnor U9764 (N_9764,N_8833,N_8842);
xnor U9765 (N_9765,N_8991,N_8506);
nand U9766 (N_9766,N_8904,N_8221);
or U9767 (N_9767,N_8864,N_8242);
or U9768 (N_9768,N_8656,N_8265);
or U9769 (N_9769,N_8352,N_8688);
or U9770 (N_9770,N_8309,N_8433);
xor U9771 (N_9771,N_8590,N_8250);
nand U9772 (N_9772,N_8091,N_8029);
nor U9773 (N_9773,N_8946,N_8181);
xnor U9774 (N_9774,N_8728,N_8716);
xnor U9775 (N_9775,N_8973,N_8122);
nand U9776 (N_9776,N_8541,N_8292);
or U9777 (N_9777,N_8789,N_8167);
and U9778 (N_9778,N_8371,N_8575);
or U9779 (N_9779,N_8536,N_8280);
nand U9780 (N_9780,N_8330,N_8263);
nor U9781 (N_9781,N_8051,N_8254);
and U9782 (N_9782,N_8927,N_8249);
or U9783 (N_9783,N_8066,N_8265);
and U9784 (N_9784,N_8687,N_8469);
and U9785 (N_9785,N_8949,N_8495);
and U9786 (N_9786,N_8897,N_8892);
and U9787 (N_9787,N_8150,N_8895);
or U9788 (N_9788,N_8325,N_8688);
nand U9789 (N_9789,N_8384,N_8186);
nor U9790 (N_9790,N_8514,N_8134);
nand U9791 (N_9791,N_8299,N_8632);
xnor U9792 (N_9792,N_8754,N_8450);
nor U9793 (N_9793,N_8481,N_8420);
nor U9794 (N_9794,N_8383,N_8467);
nor U9795 (N_9795,N_8072,N_8194);
and U9796 (N_9796,N_8178,N_8845);
nand U9797 (N_9797,N_8360,N_8159);
nand U9798 (N_9798,N_8086,N_8605);
nand U9799 (N_9799,N_8874,N_8607);
and U9800 (N_9800,N_8479,N_8786);
and U9801 (N_9801,N_8381,N_8018);
and U9802 (N_9802,N_8105,N_8266);
nand U9803 (N_9803,N_8248,N_8321);
and U9804 (N_9804,N_8126,N_8598);
or U9805 (N_9805,N_8698,N_8584);
nor U9806 (N_9806,N_8424,N_8592);
and U9807 (N_9807,N_8092,N_8479);
and U9808 (N_9808,N_8854,N_8772);
or U9809 (N_9809,N_8207,N_8616);
or U9810 (N_9810,N_8476,N_8700);
and U9811 (N_9811,N_8870,N_8068);
and U9812 (N_9812,N_8498,N_8804);
and U9813 (N_9813,N_8271,N_8636);
nand U9814 (N_9814,N_8384,N_8090);
or U9815 (N_9815,N_8481,N_8551);
nor U9816 (N_9816,N_8432,N_8816);
nand U9817 (N_9817,N_8333,N_8579);
nand U9818 (N_9818,N_8249,N_8595);
or U9819 (N_9819,N_8343,N_8872);
and U9820 (N_9820,N_8259,N_8080);
nand U9821 (N_9821,N_8952,N_8262);
or U9822 (N_9822,N_8092,N_8653);
nand U9823 (N_9823,N_8588,N_8582);
or U9824 (N_9824,N_8872,N_8687);
nand U9825 (N_9825,N_8967,N_8121);
and U9826 (N_9826,N_8222,N_8552);
nor U9827 (N_9827,N_8259,N_8238);
nand U9828 (N_9828,N_8453,N_8319);
or U9829 (N_9829,N_8812,N_8751);
nand U9830 (N_9830,N_8324,N_8394);
or U9831 (N_9831,N_8381,N_8616);
nor U9832 (N_9832,N_8618,N_8067);
or U9833 (N_9833,N_8774,N_8004);
nand U9834 (N_9834,N_8137,N_8289);
nand U9835 (N_9835,N_8130,N_8929);
nand U9836 (N_9836,N_8891,N_8530);
or U9837 (N_9837,N_8542,N_8391);
nor U9838 (N_9838,N_8478,N_8868);
and U9839 (N_9839,N_8726,N_8139);
and U9840 (N_9840,N_8709,N_8293);
and U9841 (N_9841,N_8355,N_8308);
nor U9842 (N_9842,N_8744,N_8238);
or U9843 (N_9843,N_8990,N_8431);
nand U9844 (N_9844,N_8907,N_8834);
nor U9845 (N_9845,N_8687,N_8113);
nand U9846 (N_9846,N_8526,N_8355);
xor U9847 (N_9847,N_8769,N_8489);
nor U9848 (N_9848,N_8845,N_8160);
and U9849 (N_9849,N_8668,N_8831);
nor U9850 (N_9850,N_8086,N_8685);
xor U9851 (N_9851,N_8783,N_8051);
or U9852 (N_9852,N_8660,N_8189);
and U9853 (N_9853,N_8747,N_8981);
nor U9854 (N_9854,N_8101,N_8676);
or U9855 (N_9855,N_8143,N_8320);
xnor U9856 (N_9856,N_8866,N_8566);
nand U9857 (N_9857,N_8804,N_8522);
xor U9858 (N_9858,N_8341,N_8822);
nor U9859 (N_9859,N_8798,N_8864);
and U9860 (N_9860,N_8128,N_8076);
nor U9861 (N_9861,N_8965,N_8524);
nor U9862 (N_9862,N_8752,N_8285);
nand U9863 (N_9863,N_8508,N_8590);
xor U9864 (N_9864,N_8008,N_8582);
nor U9865 (N_9865,N_8583,N_8984);
or U9866 (N_9866,N_8224,N_8660);
xnor U9867 (N_9867,N_8702,N_8030);
nand U9868 (N_9868,N_8136,N_8110);
nor U9869 (N_9869,N_8214,N_8148);
xor U9870 (N_9870,N_8331,N_8332);
nand U9871 (N_9871,N_8932,N_8445);
nand U9872 (N_9872,N_8711,N_8306);
nand U9873 (N_9873,N_8351,N_8857);
or U9874 (N_9874,N_8849,N_8784);
and U9875 (N_9875,N_8946,N_8924);
xor U9876 (N_9876,N_8499,N_8412);
nand U9877 (N_9877,N_8721,N_8045);
nor U9878 (N_9878,N_8859,N_8698);
or U9879 (N_9879,N_8928,N_8402);
and U9880 (N_9880,N_8950,N_8191);
or U9881 (N_9881,N_8956,N_8973);
nand U9882 (N_9882,N_8324,N_8290);
nand U9883 (N_9883,N_8218,N_8435);
or U9884 (N_9884,N_8300,N_8125);
or U9885 (N_9885,N_8234,N_8196);
nand U9886 (N_9886,N_8444,N_8767);
xor U9887 (N_9887,N_8916,N_8294);
xor U9888 (N_9888,N_8406,N_8687);
or U9889 (N_9889,N_8199,N_8286);
or U9890 (N_9890,N_8586,N_8905);
and U9891 (N_9891,N_8963,N_8596);
nor U9892 (N_9892,N_8472,N_8753);
or U9893 (N_9893,N_8985,N_8218);
or U9894 (N_9894,N_8957,N_8473);
and U9895 (N_9895,N_8923,N_8220);
nor U9896 (N_9896,N_8255,N_8977);
nor U9897 (N_9897,N_8626,N_8812);
nor U9898 (N_9898,N_8187,N_8434);
nor U9899 (N_9899,N_8678,N_8600);
xor U9900 (N_9900,N_8222,N_8670);
nand U9901 (N_9901,N_8095,N_8788);
nand U9902 (N_9902,N_8316,N_8055);
nand U9903 (N_9903,N_8884,N_8632);
nand U9904 (N_9904,N_8447,N_8393);
xnor U9905 (N_9905,N_8462,N_8756);
and U9906 (N_9906,N_8072,N_8973);
xor U9907 (N_9907,N_8032,N_8310);
nand U9908 (N_9908,N_8355,N_8640);
xnor U9909 (N_9909,N_8574,N_8190);
xor U9910 (N_9910,N_8116,N_8025);
or U9911 (N_9911,N_8769,N_8667);
nor U9912 (N_9912,N_8483,N_8244);
xnor U9913 (N_9913,N_8831,N_8138);
or U9914 (N_9914,N_8657,N_8345);
or U9915 (N_9915,N_8607,N_8614);
nor U9916 (N_9916,N_8208,N_8760);
and U9917 (N_9917,N_8841,N_8061);
or U9918 (N_9918,N_8536,N_8007);
nor U9919 (N_9919,N_8834,N_8539);
nand U9920 (N_9920,N_8262,N_8539);
xor U9921 (N_9921,N_8800,N_8189);
or U9922 (N_9922,N_8332,N_8250);
or U9923 (N_9923,N_8099,N_8199);
nor U9924 (N_9924,N_8364,N_8202);
or U9925 (N_9925,N_8042,N_8494);
nor U9926 (N_9926,N_8430,N_8907);
nor U9927 (N_9927,N_8525,N_8913);
or U9928 (N_9928,N_8323,N_8311);
xor U9929 (N_9929,N_8093,N_8126);
and U9930 (N_9930,N_8430,N_8446);
nand U9931 (N_9931,N_8533,N_8432);
nand U9932 (N_9932,N_8792,N_8285);
and U9933 (N_9933,N_8922,N_8547);
or U9934 (N_9934,N_8568,N_8125);
xor U9935 (N_9935,N_8974,N_8821);
or U9936 (N_9936,N_8762,N_8367);
or U9937 (N_9937,N_8517,N_8208);
xnor U9938 (N_9938,N_8791,N_8806);
nor U9939 (N_9939,N_8892,N_8761);
xnor U9940 (N_9940,N_8427,N_8059);
nand U9941 (N_9941,N_8622,N_8312);
nand U9942 (N_9942,N_8860,N_8296);
xnor U9943 (N_9943,N_8445,N_8748);
nand U9944 (N_9944,N_8978,N_8908);
xnor U9945 (N_9945,N_8109,N_8420);
xnor U9946 (N_9946,N_8069,N_8132);
or U9947 (N_9947,N_8160,N_8593);
nor U9948 (N_9948,N_8616,N_8533);
and U9949 (N_9949,N_8143,N_8321);
nor U9950 (N_9950,N_8865,N_8233);
and U9951 (N_9951,N_8327,N_8092);
xor U9952 (N_9952,N_8106,N_8048);
or U9953 (N_9953,N_8061,N_8028);
nand U9954 (N_9954,N_8017,N_8327);
or U9955 (N_9955,N_8975,N_8982);
and U9956 (N_9956,N_8972,N_8384);
and U9957 (N_9957,N_8045,N_8717);
xnor U9958 (N_9958,N_8111,N_8066);
xnor U9959 (N_9959,N_8301,N_8543);
or U9960 (N_9960,N_8662,N_8987);
or U9961 (N_9961,N_8742,N_8002);
nand U9962 (N_9962,N_8634,N_8803);
nor U9963 (N_9963,N_8590,N_8668);
xnor U9964 (N_9964,N_8298,N_8984);
and U9965 (N_9965,N_8235,N_8778);
or U9966 (N_9966,N_8461,N_8643);
nand U9967 (N_9967,N_8058,N_8019);
or U9968 (N_9968,N_8503,N_8922);
nand U9969 (N_9969,N_8825,N_8136);
or U9970 (N_9970,N_8949,N_8894);
and U9971 (N_9971,N_8213,N_8301);
nor U9972 (N_9972,N_8095,N_8385);
nor U9973 (N_9973,N_8140,N_8310);
xnor U9974 (N_9974,N_8215,N_8361);
xor U9975 (N_9975,N_8632,N_8491);
nor U9976 (N_9976,N_8724,N_8781);
xor U9977 (N_9977,N_8046,N_8926);
and U9978 (N_9978,N_8826,N_8797);
nand U9979 (N_9979,N_8091,N_8415);
or U9980 (N_9980,N_8481,N_8427);
nand U9981 (N_9981,N_8482,N_8644);
nor U9982 (N_9982,N_8130,N_8481);
nand U9983 (N_9983,N_8139,N_8741);
nor U9984 (N_9984,N_8887,N_8514);
and U9985 (N_9985,N_8605,N_8206);
xor U9986 (N_9986,N_8728,N_8097);
xor U9987 (N_9987,N_8177,N_8558);
and U9988 (N_9988,N_8837,N_8117);
or U9989 (N_9989,N_8861,N_8771);
nand U9990 (N_9990,N_8587,N_8915);
nor U9991 (N_9991,N_8847,N_8656);
or U9992 (N_9992,N_8421,N_8566);
and U9993 (N_9993,N_8541,N_8628);
nand U9994 (N_9994,N_8716,N_8143);
or U9995 (N_9995,N_8108,N_8505);
xnor U9996 (N_9996,N_8008,N_8541);
nand U9997 (N_9997,N_8819,N_8216);
or U9998 (N_9998,N_8328,N_8609);
and U9999 (N_9999,N_8577,N_8707);
nand U10000 (N_10000,N_9401,N_9022);
and U10001 (N_10001,N_9934,N_9704);
nor U10002 (N_10002,N_9292,N_9363);
or U10003 (N_10003,N_9259,N_9491);
xnor U10004 (N_10004,N_9318,N_9312);
nand U10005 (N_10005,N_9624,N_9775);
or U10006 (N_10006,N_9416,N_9516);
nand U10007 (N_10007,N_9920,N_9229);
nor U10008 (N_10008,N_9531,N_9530);
or U10009 (N_10009,N_9771,N_9782);
or U10010 (N_10010,N_9099,N_9681);
nor U10011 (N_10011,N_9223,N_9371);
nor U10012 (N_10012,N_9072,N_9674);
xor U10013 (N_10013,N_9939,N_9859);
xor U10014 (N_10014,N_9694,N_9120);
xor U10015 (N_10015,N_9357,N_9869);
and U10016 (N_10016,N_9861,N_9595);
nor U10017 (N_10017,N_9776,N_9945);
xor U10018 (N_10018,N_9262,N_9266);
nand U10019 (N_10019,N_9239,N_9247);
nand U10020 (N_10020,N_9629,N_9333);
or U10021 (N_10021,N_9358,N_9592);
or U10022 (N_10022,N_9682,N_9524);
nor U10023 (N_10023,N_9575,N_9112);
nand U10024 (N_10024,N_9211,N_9482);
or U10025 (N_10025,N_9621,N_9314);
nor U10026 (N_10026,N_9744,N_9885);
nor U10027 (N_10027,N_9911,N_9634);
nor U10028 (N_10028,N_9620,N_9270);
nand U10029 (N_10029,N_9503,N_9253);
nand U10030 (N_10030,N_9369,N_9457);
nor U10031 (N_10031,N_9951,N_9053);
nor U10032 (N_10032,N_9195,N_9774);
nand U10033 (N_10033,N_9581,N_9930);
and U10034 (N_10034,N_9940,N_9403);
xnor U10035 (N_10035,N_9683,N_9556);
nand U10036 (N_10036,N_9111,N_9467);
and U10037 (N_10037,N_9721,N_9626);
xnor U10038 (N_10038,N_9608,N_9154);
or U10039 (N_10039,N_9660,N_9716);
and U10040 (N_10040,N_9236,N_9548);
nor U10041 (N_10041,N_9271,N_9156);
nand U10042 (N_10042,N_9280,N_9673);
nor U10043 (N_10043,N_9577,N_9559);
and U10044 (N_10044,N_9038,N_9442);
or U10045 (N_10045,N_9356,N_9695);
xnor U10046 (N_10046,N_9009,N_9452);
or U10047 (N_10047,N_9554,N_9488);
and U10048 (N_10048,N_9421,N_9670);
nand U10049 (N_10049,N_9545,N_9551);
nand U10050 (N_10050,N_9919,N_9272);
xnor U10051 (N_10051,N_9227,N_9470);
nand U10052 (N_10052,N_9522,N_9310);
nand U10053 (N_10053,N_9046,N_9102);
nand U10054 (N_10054,N_9769,N_9844);
xor U10055 (N_10055,N_9365,N_9364);
nand U10056 (N_10056,N_9507,N_9486);
nor U10057 (N_10057,N_9777,N_9607);
or U10058 (N_10058,N_9726,N_9792);
and U10059 (N_10059,N_9203,N_9068);
nand U10060 (N_10060,N_9468,N_9037);
nand U10061 (N_10061,N_9534,N_9164);
and U10062 (N_10062,N_9377,N_9886);
nand U10063 (N_10063,N_9205,N_9323);
and U10064 (N_10064,N_9331,N_9031);
and U10065 (N_10065,N_9754,N_9167);
or U10066 (N_10066,N_9857,N_9804);
or U10067 (N_10067,N_9100,N_9348);
nor U10068 (N_10068,N_9615,N_9131);
xnor U10069 (N_10069,N_9284,N_9512);
xor U10070 (N_10070,N_9678,N_9879);
nor U10071 (N_10071,N_9258,N_9207);
xnor U10072 (N_10072,N_9130,N_9995);
or U10073 (N_10073,N_9246,N_9648);
or U10074 (N_10074,N_9631,N_9872);
xnor U10075 (N_10075,N_9260,N_9090);
nor U10076 (N_10076,N_9394,N_9226);
nand U10077 (N_10077,N_9847,N_9813);
and U10078 (N_10078,N_9697,N_9650);
xnor U10079 (N_10079,N_9484,N_9293);
or U10080 (N_10080,N_9108,N_9836);
nand U10081 (N_10081,N_9501,N_9533);
nand U10082 (N_10082,N_9079,N_9557);
or U10083 (N_10083,N_9330,N_9301);
xor U10084 (N_10084,N_9839,N_9938);
nand U10085 (N_10085,N_9334,N_9448);
nor U10086 (N_10086,N_9181,N_9722);
and U10087 (N_10087,N_9909,N_9538);
or U10088 (N_10088,N_9180,N_9191);
or U10089 (N_10089,N_9671,N_9489);
and U10090 (N_10090,N_9360,N_9736);
nand U10091 (N_10091,N_9216,N_9101);
xnor U10092 (N_10092,N_9322,N_9587);
xnor U10093 (N_10093,N_9659,N_9997);
xor U10094 (N_10094,N_9431,N_9618);
and U10095 (N_10095,N_9989,N_9687);
and U10096 (N_10096,N_9441,N_9791);
nor U10097 (N_10097,N_9815,N_9640);
or U10098 (N_10098,N_9252,N_9908);
nor U10099 (N_10099,N_9917,N_9641);
or U10100 (N_10100,N_9460,N_9596);
nand U10101 (N_10101,N_9389,N_9235);
xnor U10102 (N_10102,N_9446,N_9213);
nor U10103 (N_10103,N_9838,N_9993);
nor U10104 (N_10104,N_9342,N_9927);
or U10105 (N_10105,N_9766,N_9924);
or U10106 (N_10106,N_9883,N_9829);
nor U10107 (N_10107,N_9513,N_9462);
xnor U10108 (N_10108,N_9669,N_9811);
nor U10109 (N_10109,N_9174,N_9854);
nor U10110 (N_10110,N_9657,N_9913);
nor U10111 (N_10111,N_9150,N_9426);
or U10112 (N_10112,N_9332,N_9921);
xnor U10113 (N_10113,N_9500,N_9043);
nand U10114 (N_10114,N_9477,N_9616);
and U10115 (N_10115,N_9047,N_9982);
xnor U10116 (N_10116,N_9395,N_9492);
xor U10117 (N_10117,N_9083,N_9054);
nand U10118 (N_10118,N_9667,N_9523);
and U10119 (N_10119,N_9555,N_9230);
or U10120 (N_10120,N_9619,N_9315);
xnor U10121 (N_10121,N_9187,N_9413);
or U10122 (N_10122,N_9455,N_9427);
nor U10123 (N_10123,N_9439,N_9851);
xor U10124 (N_10124,N_9042,N_9387);
xor U10125 (N_10125,N_9378,N_9081);
and U10126 (N_10126,N_9021,N_9093);
and U10127 (N_10127,N_9275,N_9625);
and U10128 (N_10128,N_9240,N_9349);
and U10129 (N_10129,N_9406,N_9677);
or U10130 (N_10130,N_9822,N_9429);
nand U10131 (N_10131,N_9296,N_9988);
nand U10132 (N_10132,N_9064,N_9162);
nor U10133 (N_10133,N_9140,N_9693);
xor U10134 (N_10134,N_9076,N_9169);
or U10135 (N_10135,N_9073,N_9243);
or U10136 (N_10136,N_9148,N_9380);
and U10137 (N_10137,N_9381,N_9008);
xor U10138 (N_10138,N_9033,N_9176);
nand U10139 (N_10139,N_9004,N_9092);
and U10140 (N_10140,N_9882,N_9566);
nor U10141 (N_10141,N_9341,N_9141);
xnor U10142 (N_10142,N_9316,N_9225);
xor U10143 (N_10143,N_9887,N_9637);
or U10144 (N_10144,N_9819,N_9599);
and U10145 (N_10145,N_9194,N_9104);
or U10146 (N_10146,N_9739,N_9543);
and U10147 (N_10147,N_9425,N_9606);
xor U10148 (N_10148,N_9490,N_9933);
xor U10149 (N_10149,N_9784,N_9653);
xor U10150 (N_10150,N_9755,N_9476);
xor U10151 (N_10151,N_9757,N_9837);
nand U10152 (N_10152,N_9153,N_9878);
and U10153 (N_10153,N_9807,N_9088);
xor U10154 (N_10154,N_9149,N_9967);
or U10155 (N_10155,N_9060,N_9422);
xor U10156 (N_10156,N_9294,N_9497);
nor U10157 (N_10157,N_9304,N_9485);
nor U10158 (N_10158,N_9443,N_9762);
or U10159 (N_10159,N_9864,N_9496);
nand U10160 (N_10160,N_9115,N_9015);
xnor U10161 (N_10161,N_9506,N_9165);
xor U10162 (N_10162,N_9445,N_9273);
or U10163 (N_10163,N_9086,N_9562);
and U10164 (N_10164,N_9466,N_9105);
nor U10165 (N_10165,N_9517,N_9898);
xor U10166 (N_10166,N_9990,N_9895);
xnor U10167 (N_10167,N_9151,N_9238);
xnor U10168 (N_10168,N_9688,N_9639);
nand U10169 (N_10169,N_9337,N_9818);
or U10170 (N_10170,N_9289,N_9125);
nor U10171 (N_10171,N_9998,N_9248);
and U10172 (N_10172,N_9579,N_9627);
and U10173 (N_10173,N_9904,N_9161);
or U10174 (N_10174,N_9221,N_9179);
nand U10175 (N_10175,N_9576,N_9094);
xor U10176 (N_10176,N_9986,N_9550);
and U10177 (N_10177,N_9824,N_9779);
nand U10178 (N_10178,N_9113,N_9372);
and U10179 (N_10179,N_9834,N_9668);
and U10180 (N_10180,N_9269,N_9144);
and U10181 (N_10181,N_9339,N_9728);
nand U10182 (N_10182,N_9831,N_9547);
nand U10183 (N_10183,N_9404,N_9944);
and U10184 (N_10184,N_9397,N_9114);
or U10185 (N_10185,N_9956,N_9758);
nor U10186 (N_10186,N_9584,N_9635);
nor U10187 (N_10187,N_9277,N_9096);
and U10188 (N_10188,N_9877,N_9655);
xnor U10189 (N_10189,N_9067,N_9256);
nor U10190 (N_10190,N_9850,N_9388);
or U10191 (N_10191,N_9706,N_9502);
nor U10192 (N_10192,N_9495,N_9400);
or U10193 (N_10193,N_9071,N_9707);
and U10194 (N_10194,N_9515,N_9261);
xor U10195 (N_10195,N_9536,N_9918);
nor U10196 (N_10196,N_9865,N_9355);
nor U10197 (N_10197,N_9080,N_9750);
or U10198 (N_10198,N_9061,N_9019);
and U10199 (N_10199,N_9329,N_9698);
xor U10200 (N_10200,N_9320,N_9578);
or U10201 (N_10201,N_9753,N_9799);
and U10202 (N_10202,N_9544,N_9741);
and U10203 (N_10203,N_9359,N_9107);
xor U10204 (N_10204,N_9402,N_9601);
or U10205 (N_10205,N_9288,N_9961);
and U10206 (N_10206,N_9307,N_9126);
or U10207 (N_10207,N_9175,N_9123);
nor U10208 (N_10208,N_9873,N_9035);
and U10209 (N_10209,N_9025,N_9379);
nor U10210 (N_10210,N_9202,N_9303);
and U10211 (N_10211,N_9712,N_9832);
nor U10212 (N_10212,N_9978,N_9219);
and U10213 (N_10213,N_9267,N_9353);
and U10214 (N_10214,N_9410,N_9504);
nand U10215 (N_10215,N_9800,N_9672);
nand U10216 (N_10216,N_9463,N_9969);
nand U10217 (N_10217,N_9833,N_9168);
nand U10218 (N_10218,N_9255,N_9862);
and U10219 (N_10219,N_9770,N_9910);
nand U10220 (N_10220,N_9013,N_9276);
or U10221 (N_10221,N_9806,N_9185);
and U10222 (N_10222,N_9208,N_9163);
nand U10223 (N_10223,N_9264,N_9214);
and U10224 (N_10224,N_9737,N_9423);
nand U10225 (N_10225,N_9604,N_9409);
or U10226 (N_10226,N_9717,N_9723);
nand U10227 (N_10227,N_9656,N_9237);
or U10228 (N_10228,N_9136,N_9350);
xnor U10229 (N_10229,N_9393,N_9302);
nand U10230 (N_10230,N_9487,N_9052);
or U10231 (N_10231,N_9049,N_9773);
nor U10232 (N_10232,N_9535,N_9705);
nand U10233 (N_10233,N_9166,N_9078);
and U10234 (N_10234,N_9138,N_9935);
or U10235 (N_10235,N_9328,N_9024);
nor U10236 (N_10236,N_9133,N_9265);
nand U10237 (N_10237,N_9868,N_9570);
xnor U10238 (N_10238,N_9417,N_9241);
xor U10239 (N_10239,N_9884,N_9875);
xor U10240 (N_10240,N_9937,N_9311);
and U10241 (N_10241,N_9709,N_9948);
nand U10242 (N_10242,N_9250,N_9305);
or U10243 (N_10243,N_9890,N_9768);
and U10244 (N_10244,N_9032,N_9563);
or U10245 (N_10245,N_9614,N_9399);
nand U10246 (N_10246,N_9891,N_9603);
nand U10247 (N_10247,N_9324,N_9980);
or U10248 (N_10248,N_9572,N_9147);
or U10249 (N_10249,N_9444,N_9647);
or U10250 (N_10250,N_9069,N_9075);
nand U10251 (N_10251,N_9597,N_9842);
xor U10252 (N_10252,N_9200,N_9374);
xnor U10253 (N_10253,N_9541,N_9765);
nor U10254 (N_10254,N_9903,N_9204);
nor U10255 (N_10255,N_9198,N_9006);
xor U10256 (N_10256,N_9233,N_9941);
nor U10257 (N_10257,N_9249,N_9011);
nand U10258 (N_10258,N_9040,N_9116);
xnor U10259 (N_10259,N_9415,N_9752);
nand U10260 (N_10260,N_9798,N_9830);
or U10261 (N_10261,N_9970,N_9244);
and U10262 (N_10262,N_9014,N_9343);
nand U10263 (N_10263,N_9591,N_9965);
or U10264 (N_10264,N_9866,N_9058);
xor U10265 (N_10265,N_9756,N_9222);
nand U10266 (N_10266,N_9007,N_9145);
nor U10267 (N_10267,N_9684,N_9821);
nand U10268 (N_10268,N_9835,N_9731);
xor U10269 (N_10269,N_9735,N_9772);
nor U10270 (N_10270,N_9055,N_9017);
nand U10271 (N_10271,N_9996,N_9118);
xor U10272 (N_10272,N_9636,N_9066);
and U10273 (N_10273,N_9880,N_9048);
or U10274 (N_10274,N_9451,N_9336);
nand U10275 (N_10275,N_9340,N_9793);
and U10276 (N_10276,N_9816,N_9494);
xnor U10277 (N_10277,N_9950,N_9178);
nand U10278 (N_10278,N_9291,N_9906);
nand U10279 (N_10279,N_9686,N_9027);
nor U10280 (N_10280,N_9170,N_9665);
nand U10281 (N_10281,N_9158,N_9801);
xor U10282 (N_10282,N_9142,N_9675);
nand U10283 (N_10283,N_9730,N_9893);
nand U10284 (N_10284,N_9991,N_9718);
and U10285 (N_10285,N_9438,N_9508);
or U10286 (N_10286,N_9041,N_9215);
xor U10287 (N_10287,N_9645,N_9110);
nor U10288 (N_10288,N_9790,N_9732);
xor U10289 (N_10289,N_9527,N_9525);
and U10290 (N_10290,N_9471,N_9977);
and U10291 (N_10291,N_9224,N_9609);
or U10292 (N_10292,N_9521,N_9385);
and U10293 (N_10293,N_9326,N_9984);
nand U10294 (N_10294,N_9119,N_9899);
and U10295 (N_10295,N_9710,N_9745);
or U10296 (N_10296,N_9802,N_9117);
and U10297 (N_10297,N_9720,N_9391);
and U10298 (N_10298,N_9796,N_9321);
xnor U10299 (N_10299,N_9568,N_9711);
or U10300 (N_10300,N_9905,N_9590);
nand U10301 (N_10301,N_9888,N_9560);
nor U10302 (N_10302,N_9795,N_9892);
xnor U10303 (N_10303,N_9407,N_9245);
nor U10304 (N_10304,N_9600,N_9605);
and U10305 (N_10305,N_9084,N_9440);
nor U10306 (N_10306,N_9912,N_9783);
xor U10307 (N_10307,N_9971,N_9499);
nand U10308 (N_10308,N_9430,N_9966);
and U10309 (N_10309,N_9580,N_9361);
nand U10310 (N_10310,N_9386,N_9690);
and U10311 (N_10311,N_9778,N_9519);
or U10312 (N_10312,N_9567,N_9797);
nand U10313 (N_10313,N_9747,N_9569);
nor U10314 (N_10314,N_9916,N_9201);
nand U10315 (N_10315,N_9992,N_9016);
or U10316 (N_10316,N_9952,N_9172);
xnor U10317 (N_10317,N_9708,N_9308);
nand U10318 (N_10318,N_9327,N_9498);
and U10319 (N_10319,N_9958,N_9623);
nand U10320 (N_10320,N_9373,N_9173);
or U10321 (N_10321,N_9999,N_9564);
nand U10322 (N_10322,N_9003,N_9433);
or U10323 (N_10323,N_9651,N_9351);
or U10324 (N_10324,N_9963,N_9594);
xor U10325 (N_10325,N_9074,N_9367);
or U10326 (N_10326,N_9109,N_9479);
nand U10327 (N_10327,N_9785,N_9692);
nor U10328 (N_10328,N_9091,N_9676);
nor U10329 (N_10329,N_9571,N_9309);
or U10330 (N_10330,N_9602,N_9345);
nor U10331 (N_10331,N_9860,N_9932);
nor U10332 (N_10332,N_9335,N_9132);
nand U10333 (N_10333,N_9023,N_9124);
xor U10334 (N_10334,N_9947,N_9474);
nor U10335 (N_10335,N_9155,N_9480);
nand U10336 (N_10336,N_9077,N_9632);
and U10337 (N_10337,N_9748,N_9464);
nand U10338 (N_10338,N_9082,N_9306);
or U10339 (N_10339,N_9146,N_9257);
or U10340 (N_10340,N_9549,N_9274);
or U10341 (N_10341,N_9781,N_9384);
nor U10342 (N_10342,N_9896,N_9696);
and U10343 (N_10343,N_9983,N_9539);
and U10344 (N_10344,N_9408,N_9218);
xor U10345 (N_10345,N_9719,N_9840);
or U10346 (N_10346,N_9232,N_9808);
or U10347 (N_10347,N_9955,N_9481);
nand U10348 (N_10348,N_9949,N_9699);
nor U10349 (N_10349,N_9810,N_9858);
xor U10350 (N_10350,N_9573,N_9788);
nand U10351 (N_10351,N_9652,N_9733);
or U10352 (N_10352,N_9186,N_9542);
or U10353 (N_10353,N_9742,N_9514);
nor U10354 (N_10354,N_9942,N_9610);
nor U10355 (N_10355,N_9354,N_9026);
and U10356 (N_10356,N_9925,N_9143);
or U10357 (N_10357,N_9209,N_9703);
nand U10358 (N_10358,N_9649,N_9411);
nand U10359 (N_10359,N_9628,N_9059);
nand U10360 (N_10360,N_9434,N_9435);
or U10361 (N_10361,N_9589,N_9290);
xnor U10362 (N_10362,N_9044,N_9190);
nand U10363 (N_10363,N_9552,N_9018);
nand U10364 (N_10364,N_9558,N_9450);
nand U10365 (N_10365,N_9680,N_9192);
or U10366 (N_10366,N_9030,N_9376);
or U10367 (N_10367,N_9749,N_9432);
and U10368 (N_10368,N_9282,N_9953);
or U10369 (N_10369,N_9994,N_9871);
nand U10370 (N_10370,N_9001,N_9390);
xnor U10371 (N_10371,N_9220,N_9894);
or U10372 (N_10372,N_9020,N_9085);
or U10373 (N_10373,N_9287,N_9812);
and U10374 (N_10374,N_9518,N_9157);
or U10375 (N_10375,N_9197,N_9297);
or U10376 (N_10376,N_9787,N_9565);
nand U10377 (N_10377,N_9537,N_9428);
xor U10378 (N_10378,N_9825,N_9405);
and U10379 (N_10379,N_9002,N_9122);
xor U10380 (N_10380,N_9613,N_9039);
nand U10381 (N_10381,N_9414,N_9964);
nand U10382 (N_10382,N_9729,N_9843);
or U10383 (N_10383,N_9889,N_9420);
nor U10384 (N_10384,N_9199,N_9398);
and U10385 (N_10385,N_9268,N_9317);
nor U10386 (N_10386,N_9593,N_9715);
nand U10387 (N_10387,N_9231,N_9658);
nor U10388 (N_10388,N_9846,N_9763);
xor U10389 (N_10389,N_9300,N_9897);
nor U10390 (N_10390,N_9689,N_9900);
nand U10391 (N_10391,N_9841,N_9612);
nand U10392 (N_10392,N_9483,N_9465);
and U10393 (N_10393,N_9574,N_9418);
and U10394 (N_10394,N_9098,N_9121);
xor U10395 (N_10395,N_9943,N_9702);
and U10396 (N_10396,N_9664,N_9051);
or U10397 (N_10397,N_9424,N_9127);
xnor U10398 (N_10398,N_9368,N_9701);
nor U10399 (N_10399,N_9976,N_9901);
nand U10400 (N_10400,N_9931,N_9028);
or U10401 (N_10401,N_9546,N_9848);
xor U10402 (N_10402,N_9902,N_9298);
nor U10403 (N_10403,N_9622,N_9396);
nor U10404 (N_10404,N_9975,N_9642);
and U10405 (N_10405,N_9461,N_9700);
nor U10406 (N_10406,N_9473,N_9981);
or U10407 (N_10407,N_9985,N_9855);
nand U10408 (N_10408,N_9299,N_9295);
xor U10409 (N_10409,N_9630,N_9805);
and U10410 (N_10410,N_9454,N_9979);
and U10411 (N_10411,N_9281,N_9863);
and U10412 (N_10412,N_9196,N_9876);
or U10413 (N_10413,N_9134,N_9057);
and U10414 (N_10414,N_9685,N_9325);
nor U10415 (N_10415,N_9820,N_9346);
nor U10416 (N_10416,N_9097,N_9193);
and U10417 (N_10417,N_9189,N_9646);
or U10418 (N_10418,N_9828,N_9780);
nand U10419 (N_10419,N_9845,N_9505);
and U10420 (N_10420,N_9743,N_9005);
or U10421 (N_10421,N_9973,N_9493);
and U10422 (N_10422,N_9050,N_9472);
nand U10423 (N_10423,N_9412,N_9638);
and U10424 (N_10424,N_9936,N_9313);
or U10425 (N_10425,N_9528,N_9987);
nand U10426 (N_10426,N_9907,N_9926);
or U10427 (N_10427,N_9714,N_9760);
or U10428 (N_10428,N_9437,N_9724);
or U10429 (N_10429,N_9852,N_9511);
nand U10430 (N_10430,N_9070,N_9914);
nor U10431 (N_10431,N_9087,N_9089);
or U10432 (N_10432,N_9242,N_9458);
nand U10433 (N_10433,N_9654,N_9974);
xor U10434 (N_10434,N_9475,N_9177);
and U10435 (N_10435,N_9362,N_9725);
or U10436 (N_10436,N_9526,N_9962);
nor U10437 (N_10437,N_9529,N_9449);
or U10438 (N_10438,N_9012,N_9746);
or U10439 (N_10439,N_9159,N_9010);
and U10440 (N_10440,N_9286,N_9585);
and U10441 (N_10441,N_9661,N_9234);
or U10442 (N_10442,N_9095,N_9520);
xor U10443 (N_10443,N_9767,N_9662);
nand U10444 (N_10444,N_9382,N_9817);
and U10445 (N_10445,N_9106,N_9338);
nor U10446 (N_10446,N_9056,N_9456);
xnor U10447 (N_10447,N_9751,N_9598);
nand U10448 (N_10448,N_9929,N_9188);
nor U10449 (N_10449,N_9922,N_9347);
and U10450 (N_10450,N_9870,N_9759);
and U10451 (N_10451,N_9786,N_9459);
xor U10452 (N_10452,N_9643,N_9065);
and U10453 (N_10453,N_9254,N_9972);
xnor U10454 (N_10454,N_9915,N_9469);
and U10455 (N_10455,N_9128,N_9881);
and U10456 (N_10456,N_9928,N_9960);
nor U10457 (N_10457,N_9849,N_9063);
xnor U10458 (N_10458,N_9867,N_9583);
xnor U10459 (N_10459,N_9135,N_9212);
or U10460 (N_10460,N_9182,N_9727);
and U10461 (N_10461,N_9814,N_9713);
xor U10462 (N_10462,N_9803,N_9352);
xor U10463 (N_10463,N_9137,N_9045);
or U10464 (N_10464,N_9509,N_9278);
nand U10465 (N_10465,N_9319,N_9954);
nand U10466 (N_10466,N_9366,N_9532);
nand U10467 (N_10467,N_9823,N_9375);
nor U10468 (N_10468,N_9738,N_9761);
or U10469 (N_10469,N_9184,N_9171);
nand U10470 (N_10470,N_9478,N_9586);
nor U10471 (N_10471,N_9827,N_9436);
nor U10472 (N_10472,N_9826,N_9553);
nor U10473 (N_10473,N_9874,N_9764);
xnor U10474 (N_10474,N_9447,N_9968);
and U10475 (N_10475,N_9959,N_9617);
nor U10476 (N_10476,N_9062,N_9383);
and U10477 (N_10477,N_9279,N_9856);
xnor U10478 (N_10478,N_9210,N_9789);
nor U10479 (N_10479,N_9183,N_9663);
and U10480 (N_10480,N_9370,N_9103);
or U10481 (N_10481,N_9263,N_9582);
xnor U10482 (N_10482,N_9679,N_9228);
nand U10483 (N_10483,N_9034,N_9160);
or U10484 (N_10484,N_9344,N_9285);
or U10485 (N_10485,N_9139,N_9217);
or U10486 (N_10486,N_9666,N_9691);
or U10487 (N_10487,N_9510,N_9152);
or U10488 (N_10488,N_9734,N_9206);
and U10489 (N_10489,N_9251,N_9000);
nor U10490 (N_10490,N_9419,N_9611);
nor U10491 (N_10491,N_9453,N_9392);
and U10492 (N_10492,N_9561,N_9794);
nand U10493 (N_10493,N_9036,N_9633);
xor U10494 (N_10494,N_9809,N_9129);
xnor U10495 (N_10495,N_9946,N_9923);
nor U10496 (N_10496,N_9853,N_9283);
and U10497 (N_10497,N_9957,N_9540);
nand U10498 (N_10498,N_9588,N_9029);
xnor U10499 (N_10499,N_9740,N_9644);
xor U10500 (N_10500,N_9468,N_9611);
nand U10501 (N_10501,N_9955,N_9658);
or U10502 (N_10502,N_9690,N_9188);
or U10503 (N_10503,N_9423,N_9252);
and U10504 (N_10504,N_9159,N_9795);
or U10505 (N_10505,N_9430,N_9261);
xor U10506 (N_10506,N_9289,N_9507);
or U10507 (N_10507,N_9432,N_9418);
and U10508 (N_10508,N_9489,N_9203);
or U10509 (N_10509,N_9358,N_9000);
and U10510 (N_10510,N_9464,N_9015);
nor U10511 (N_10511,N_9932,N_9799);
xnor U10512 (N_10512,N_9714,N_9062);
nor U10513 (N_10513,N_9450,N_9879);
xnor U10514 (N_10514,N_9115,N_9248);
xnor U10515 (N_10515,N_9747,N_9154);
or U10516 (N_10516,N_9548,N_9863);
nor U10517 (N_10517,N_9428,N_9060);
nand U10518 (N_10518,N_9737,N_9398);
nand U10519 (N_10519,N_9536,N_9958);
xor U10520 (N_10520,N_9093,N_9774);
or U10521 (N_10521,N_9100,N_9168);
nand U10522 (N_10522,N_9984,N_9023);
nor U10523 (N_10523,N_9894,N_9911);
or U10524 (N_10524,N_9637,N_9449);
nand U10525 (N_10525,N_9287,N_9403);
and U10526 (N_10526,N_9614,N_9224);
or U10527 (N_10527,N_9660,N_9856);
xor U10528 (N_10528,N_9177,N_9200);
xor U10529 (N_10529,N_9101,N_9554);
and U10530 (N_10530,N_9645,N_9809);
or U10531 (N_10531,N_9215,N_9846);
xor U10532 (N_10532,N_9131,N_9864);
or U10533 (N_10533,N_9063,N_9622);
and U10534 (N_10534,N_9024,N_9281);
nor U10535 (N_10535,N_9714,N_9810);
and U10536 (N_10536,N_9855,N_9310);
nand U10537 (N_10537,N_9210,N_9919);
or U10538 (N_10538,N_9637,N_9092);
or U10539 (N_10539,N_9270,N_9520);
xor U10540 (N_10540,N_9442,N_9048);
or U10541 (N_10541,N_9206,N_9160);
and U10542 (N_10542,N_9542,N_9824);
nor U10543 (N_10543,N_9309,N_9046);
xnor U10544 (N_10544,N_9783,N_9609);
and U10545 (N_10545,N_9767,N_9513);
or U10546 (N_10546,N_9522,N_9606);
nor U10547 (N_10547,N_9933,N_9022);
or U10548 (N_10548,N_9258,N_9626);
and U10549 (N_10549,N_9733,N_9070);
nor U10550 (N_10550,N_9357,N_9196);
nor U10551 (N_10551,N_9741,N_9332);
and U10552 (N_10552,N_9372,N_9974);
nand U10553 (N_10553,N_9766,N_9037);
or U10554 (N_10554,N_9474,N_9208);
or U10555 (N_10555,N_9860,N_9590);
and U10556 (N_10556,N_9261,N_9435);
and U10557 (N_10557,N_9492,N_9941);
or U10558 (N_10558,N_9287,N_9011);
xor U10559 (N_10559,N_9295,N_9517);
nor U10560 (N_10560,N_9621,N_9390);
or U10561 (N_10561,N_9210,N_9528);
and U10562 (N_10562,N_9258,N_9426);
or U10563 (N_10563,N_9670,N_9870);
xor U10564 (N_10564,N_9447,N_9245);
nand U10565 (N_10565,N_9168,N_9056);
nand U10566 (N_10566,N_9085,N_9121);
or U10567 (N_10567,N_9493,N_9172);
nor U10568 (N_10568,N_9594,N_9791);
nand U10569 (N_10569,N_9258,N_9296);
or U10570 (N_10570,N_9502,N_9483);
nor U10571 (N_10571,N_9796,N_9432);
nand U10572 (N_10572,N_9826,N_9283);
and U10573 (N_10573,N_9245,N_9130);
or U10574 (N_10574,N_9091,N_9668);
nand U10575 (N_10575,N_9514,N_9583);
xor U10576 (N_10576,N_9165,N_9692);
nor U10577 (N_10577,N_9523,N_9059);
xnor U10578 (N_10578,N_9679,N_9224);
nand U10579 (N_10579,N_9135,N_9327);
and U10580 (N_10580,N_9692,N_9615);
and U10581 (N_10581,N_9232,N_9746);
or U10582 (N_10582,N_9240,N_9031);
nor U10583 (N_10583,N_9455,N_9270);
and U10584 (N_10584,N_9070,N_9560);
nand U10585 (N_10585,N_9663,N_9698);
xnor U10586 (N_10586,N_9822,N_9444);
nor U10587 (N_10587,N_9585,N_9740);
or U10588 (N_10588,N_9123,N_9034);
xor U10589 (N_10589,N_9648,N_9195);
or U10590 (N_10590,N_9968,N_9695);
nor U10591 (N_10591,N_9623,N_9955);
nand U10592 (N_10592,N_9276,N_9122);
and U10593 (N_10593,N_9342,N_9609);
xnor U10594 (N_10594,N_9347,N_9862);
nand U10595 (N_10595,N_9956,N_9049);
or U10596 (N_10596,N_9610,N_9853);
or U10597 (N_10597,N_9363,N_9996);
and U10598 (N_10598,N_9630,N_9170);
or U10599 (N_10599,N_9389,N_9572);
nor U10600 (N_10600,N_9613,N_9917);
xor U10601 (N_10601,N_9802,N_9390);
and U10602 (N_10602,N_9410,N_9952);
and U10603 (N_10603,N_9631,N_9044);
xor U10604 (N_10604,N_9535,N_9580);
nor U10605 (N_10605,N_9579,N_9348);
nand U10606 (N_10606,N_9952,N_9751);
xnor U10607 (N_10607,N_9269,N_9100);
nor U10608 (N_10608,N_9801,N_9232);
nand U10609 (N_10609,N_9311,N_9314);
or U10610 (N_10610,N_9479,N_9679);
and U10611 (N_10611,N_9355,N_9320);
or U10612 (N_10612,N_9164,N_9203);
xnor U10613 (N_10613,N_9002,N_9019);
xor U10614 (N_10614,N_9903,N_9194);
xnor U10615 (N_10615,N_9887,N_9511);
and U10616 (N_10616,N_9705,N_9237);
xnor U10617 (N_10617,N_9551,N_9860);
and U10618 (N_10618,N_9882,N_9953);
nor U10619 (N_10619,N_9925,N_9157);
or U10620 (N_10620,N_9492,N_9713);
nor U10621 (N_10621,N_9241,N_9178);
nor U10622 (N_10622,N_9801,N_9013);
or U10623 (N_10623,N_9232,N_9053);
and U10624 (N_10624,N_9082,N_9133);
nor U10625 (N_10625,N_9905,N_9143);
nor U10626 (N_10626,N_9380,N_9489);
nor U10627 (N_10627,N_9989,N_9223);
nand U10628 (N_10628,N_9030,N_9535);
nor U10629 (N_10629,N_9617,N_9449);
nand U10630 (N_10630,N_9788,N_9104);
and U10631 (N_10631,N_9862,N_9065);
nor U10632 (N_10632,N_9256,N_9469);
or U10633 (N_10633,N_9317,N_9865);
nor U10634 (N_10634,N_9623,N_9789);
or U10635 (N_10635,N_9607,N_9871);
nor U10636 (N_10636,N_9633,N_9075);
nand U10637 (N_10637,N_9201,N_9816);
xnor U10638 (N_10638,N_9799,N_9052);
or U10639 (N_10639,N_9914,N_9186);
nand U10640 (N_10640,N_9481,N_9193);
nand U10641 (N_10641,N_9029,N_9349);
and U10642 (N_10642,N_9113,N_9244);
nand U10643 (N_10643,N_9041,N_9557);
or U10644 (N_10644,N_9951,N_9397);
nand U10645 (N_10645,N_9097,N_9473);
or U10646 (N_10646,N_9547,N_9389);
nand U10647 (N_10647,N_9850,N_9875);
nand U10648 (N_10648,N_9036,N_9790);
and U10649 (N_10649,N_9069,N_9741);
or U10650 (N_10650,N_9453,N_9510);
and U10651 (N_10651,N_9026,N_9650);
nor U10652 (N_10652,N_9451,N_9351);
nand U10653 (N_10653,N_9803,N_9616);
and U10654 (N_10654,N_9902,N_9827);
and U10655 (N_10655,N_9431,N_9453);
xor U10656 (N_10656,N_9794,N_9935);
and U10657 (N_10657,N_9453,N_9607);
or U10658 (N_10658,N_9792,N_9670);
nand U10659 (N_10659,N_9056,N_9043);
and U10660 (N_10660,N_9834,N_9930);
and U10661 (N_10661,N_9960,N_9887);
nand U10662 (N_10662,N_9898,N_9514);
xnor U10663 (N_10663,N_9626,N_9411);
and U10664 (N_10664,N_9206,N_9240);
nor U10665 (N_10665,N_9965,N_9534);
nor U10666 (N_10666,N_9586,N_9353);
xor U10667 (N_10667,N_9964,N_9042);
nand U10668 (N_10668,N_9421,N_9817);
and U10669 (N_10669,N_9082,N_9564);
nor U10670 (N_10670,N_9924,N_9200);
nand U10671 (N_10671,N_9792,N_9215);
and U10672 (N_10672,N_9828,N_9667);
xnor U10673 (N_10673,N_9970,N_9472);
xor U10674 (N_10674,N_9441,N_9917);
xor U10675 (N_10675,N_9281,N_9442);
and U10676 (N_10676,N_9741,N_9013);
nor U10677 (N_10677,N_9924,N_9109);
and U10678 (N_10678,N_9721,N_9357);
and U10679 (N_10679,N_9169,N_9267);
nand U10680 (N_10680,N_9700,N_9595);
or U10681 (N_10681,N_9057,N_9029);
and U10682 (N_10682,N_9992,N_9653);
nor U10683 (N_10683,N_9604,N_9501);
xnor U10684 (N_10684,N_9380,N_9647);
nor U10685 (N_10685,N_9265,N_9344);
nand U10686 (N_10686,N_9471,N_9179);
or U10687 (N_10687,N_9603,N_9576);
and U10688 (N_10688,N_9526,N_9609);
nand U10689 (N_10689,N_9648,N_9454);
xnor U10690 (N_10690,N_9711,N_9375);
nor U10691 (N_10691,N_9361,N_9607);
and U10692 (N_10692,N_9010,N_9098);
or U10693 (N_10693,N_9665,N_9563);
nor U10694 (N_10694,N_9523,N_9570);
or U10695 (N_10695,N_9675,N_9484);
or U10696 (N_10696,N_9977,N_9540);
xnor U10697 (N_10697,N_9739,N_9571);
nor U10698 (N_10698,N_9431,N_9911);
or U10699 (N_10699,N_9111,N_9854);
nor U10700 (N_10700,N_9022,N_9019);
nand U10701 (N_10701,N_9555,N_9833);
xor U10702 (N_10702,N_9394,N_9096);
xnor U10703 (N_10703,N_9997,N_9208);
and U10704 (N_10704,N_9242,N_9162);
and U10705 (N_10705,N_9341,N_9784);
nand U10706 (N_10706,N_9636,N_9126);
nand U10707 (N_10707,N_9508,N_9891);
nand U10708 (N_10708,N_9536,N_9935);
nor U10709 (N_10709,N_9772,N_9669);
nor U10710 (N_10710,N_9675,N_9188);
nand U10711 (N_10711,N_9412,N_9155);
xor U10712 (N_10712,N_9683,N_9098);
xnor U10713 (N_10713,N_9991,N_9297);
nand U10714 (N_10714,N_9218,N_9844);
nor U10715 (N_10715,N_9929,N_9620);
or U10716 (N_10716,N_9052,N_9442);
nand U10717 (N_10717,N_9773,N_9879);
and U10718 (N_10718,N_9606,N_9472);
xnor U10719 (N_10719,N_9791,N_9549);
and U10720 (N_10720,N_9127,N_9262);
xnor U10721 (N_10721,N_9242,N_9867);
or U10722 (N_10722,N_9203,N_9356);
nor U10723 (N_10723,N_9077,N_9651);
nand U10724 (N_10724,N_9310,N_9931);
nor U10725 (N_10725,N_9027,N_9824);
nor U10726 (N_10726,N_9954,N_9761);
or U10727 (N_10727,N_9105,N_9993);
xnor U10728 (N_10728,N_9517,N_9881);
nor U10729 (N_10729,N_9645,N_9610);
or U10730 (N_10730,N_9068,N_9593);
nand U10731 (N_10731,N_9565,N_9719);
or U10732 (N_10732,N_9386,N_9459);
xnor U10733 (N_10733,N_9879,N_9250);
nor U10734 (N_10734,N_9992,N_9809);
xor U10735 (N_10735,N_9117,N_9914);
nand U10736 (N_10736,N_9789,N_9312);
xnor U10737 (N_10737,N_9275,N_9998);
or U10738 (N_10738,N_9966,N_9380);
xnor U10739 (N_10739,N_9627,N_9735);
and U10740 (N_10740,N_9485,N_9272);
and U10741 (N_10741,N_9521,N_9917);
xnor U10742 (N_10742,N_9087,N_9110);
xor U10743 (N_10743,N_9418,N_9795);
nor U10744 (N_10744,N_9562,N_9736);
or U10745 (N_10745,N_9864,N_9121);
or U10746 (N_10746,N_9520,N_9412);
and U10747 (N_10747,N_9670,N_9635);
or U10748 (N_10748,N_9614,N_9635);
nand U10749 (N_10749,N_9147,N_9777);
or U10750 (N_10750,N_9770,N_9254);
and U10751 (N_10751,N_9264,N_9756);
nand U10752 (N_10752,N_9814,N_9560);
nor U10753 (N_10753,N_9217,N_9832);
nor U10754 (N_10754,N_9182,N_9206);
nand U10755 (N_10755,N_9431,N_9482);
or U10756 (N_10756,N_9093,N_9692);
nor U10757 (N_10757,N_9533,N_9843);
and U10758 (N_10758,N_9650,N_9800);
nor U10759 (N_10759,N_9024,N_9286);
nor U10760 (N_10760,N_9074,N_9315);
or U10761 (N_10761,N_9847,N_9374);
and U10762 (N_10762,N_9761,N_9640);
and U10763 (N_10763,N_9098,N_9802);
xor U10764 (N_10764,N_9102,N_9352);
or U10765 (N_10765,N_9479,N_9595);
nand U10766 (N_10766,N_9235,N_9988);
xnor U10767 (N_10767,N_9787,N_9603);
and U10768 (N_10768,N_9600,N_9938);
and U10769 (N_10769,N_9370,N_9234);
nor U10770 (N_10770,N_9553,N_9452);
xnor U10771 (N_10771,N_9167,N_9649);
nand U10772 (N_10772,N_9393,N_9146);
and U10773 (N_10773,N_9794,N_9070);
nor U10774 (N_10774,N_9570,N_9314);
xnor U10775 (N_10775,N_9764,N_9173);
xor U10776 (N_10776,N_9236,N_9115);
and U10777 (N_10777,N_9459,N_9741);
xor U10778 (N_10778,N_9580,N_9420);
xor U10779 (N_10779,N_9329,N_9191);
and U10780 (N_10780,N_9143,N_9829);
or U10781 (N_10781,N_9179,N_9325);
or U10782 (N_10782,N_9696,N_9415);
xnor U10783 (N_10783,N_9465,N_9216);
xnor U10784 (N_10784,N_9066,N_9259);
and U10785 (N_10785,N_9712,N_9897);
or U10786 (N_10786,N_9916,N_9750);
nor U10787 (N_10787,N_9095,N_9293);
or U10788 (N_10788,N_9457,N_9363);
or U10789 (N_10789,N_9360,N_9160);
nor U10790 (N_10790,N_9789,N_9062);
and U10791 (N_10791,N_9541,N_9660);
and U10792 (N_10792,N_9145,N_9390);
nor U10793 (N_10793,N_9324,N_9457);
or U10794 (N_10794,N_9257,N_9166);
xor U10795 (N_10795,N_9846,N_9488);
xnor U10796 (N_10796,N_9439,N_9622);
nor U10797 (N_10797,N_9328,N_9323);
nor U10798 (N_10798,N_9093,N_9015);
nand U10799 (N_10799,N_9920,N_9327);
nand U10800 (N_10800,N_9388,N_9727);
and U10801 (N_10801,N_9497,N_9706);
nand U10802 (N_10802,N_9686,N_9424);
and U10803 (N_10803,N_9588,N_9227);
xor U10804 (N_10804,N_9727,N_9192);
and U10805 (N_10805,N_9231,N_9928);
nand U10806 (N_10806,N_9262,N_9975);
nand U10807 (N_10807,N_9688,N_9935);
nor U10808 (N_10808,N_9345,N_9914);
and U10809 (N_10809,N_9557,N_9176);
and U10810 (N_10810,N_9519,N_9514);
and U10811 (N_10811,N_9317,N_9193);
nor U10812 (N_10812,N_9538,N_9831);
and U10813 (N_10813,N_9050,N_9812);
or U10814 (N_10814,N_9925,N_9161);
nand U10815 (N_10815,N_9513,N_9010);
xor U10816 (N_10816,N_9072,N_9820);
nor U10817 (N_10817,N_9935,N_9382);
and U10818 (N_10818,N_9820,N_9590);
xnor U10819 (N_10819,N_9982,N_9419);
nand U10820 (N_10820,N_9189,N_9463);
and U10821 (N_10821,N_9157,N_9336);
xor U10822 (N_10822,N_9523,N_9900);
and U10823 (N_10823,N_9122,N_9129);
nand U10824 (N_10824,N_9365,N_9540);
xnor U10825 (N_10825,N_9869,N_9366);
xor U10826 (N_10826,N_9054,N_9475);
or U10827 (N_10827,N_9892,N_9440);
nor U10828 (N_10828,N_9450,N_9689);
or U10829 (N_10829,N_9031,N_9369);
xnor U10830 (N_10830,N_9793,N_9816);
nor U10831 (N_10831,N_9604,N_9020);
and U10832 (N_10832,N_9431,N_9104);
xor U10833 (N_10833,N_9312,N_9023);
nor U10834 (N_10834,N_9125,N_9282);
xnor U10835 (N_10835,N_9955,N_9451);
and U10836 (N_10836,N_9570,N_9344);
nor U10837 (N_10837,N_9035,N_9413);
nand U10838 (N_10838,N_9791,N_9028);
or U10839 (N_10839,N_9950,N_9800);
nand U10840 (N_10840,N_9857,N_9148);
and U10841 (N_10841,N_9971,N_9326);
or U10842 (N_10842,N_9597,N_9192);
nor U10843 (N_10843,N_9087,N_9120);
or U10844 (N_10844,N_9020,N_9116);
xor U10845 (N_10845,N_9155,N_9630);
or U10846 (N_10846,N_9089,N_9791);
nor U10847 (N_10847,N_9071,N_9232);
nand U10848 (N_10848,N_9260,N_9536);
xnor U10849 (N_10849,N_9533,N_9566);
nor U10850 (N_10850,N_9452,N_9237);
or U10851 (N_10851,N_9687,N_9629);
xor U10852 (N_10852,N_9240,N_9171);
xnor U10853 (N_10853,N_9368,N_9639);
nor U10854 (N_10854,N_9621,N_9160);
nor U10855 (N_10855,N_9846,N_9930);
nand U10856 (N_10856,N_9259,N_9542);
nand U10857 (N_10857,N_9244,N_9945);
xor U10858 (N_10858,N_9245,N_9453);
xnor U10859 (N_10859,N_9818,N_9788);
nor U10860 (N_10860,N_9618,N_9695);
or U10861 (N_10861,N_9095,N_9909);
and U10862 (N_10862,N_9299,N_9846);
and U10863 (N_10863,N_9894,N_9298);
and U10864 (N_10864,N_9683,N_9590);
and U10865 (N_10865,N_9043,N_9480);
and U10866 (N_10866,N_9055,N_9635);
and U10867 (N_10867,N_9389,N_9858);
xor U10868 (N_10868,N_9853,N_9665);
xor U10869 (N_10869,N_9285,N_9917);
nor U10870 (N_10870,N_9501,N_9280);
or U10871 (N_10871,N_9626,N_9279);
xor U10872 (N_10872,N_9763,N_9739);
and U10873 (N_10873,N_9311,N_9565);
or U10874 (N_10874,N_9596,N_9725);
nand U10875 (N_10875,N_9460,N_9160);
nand U10876 (N_10876,N_9016,N_9247);
nand U10877 (N_10877,N_9696,N_9428);
nand U10878 (N_10878,N_9625,N_9953);
xor U10879 (N_10879,N_9144,N_9587);
nand U10880 (N_10880,N_9595,N_9488);
nand U10881 (N_10881,N_9175,N_9416);
xnor U10882 (N_10882,N_9814,N_9073);
or U10883 (N_10883,N_9382,N_9455);
or U10884 (N_10884,N_9395,N_9574);
nand U10885 (N_10885,N_9257,N_9691);
and U10886 (N_10886,N_9606,N_9718);
or U10887 (N_10887,N_9383,N_9044);
xnor U10888 (N_10888,N_9263,N_9763);
nand U10889 (N_10889,N_9587,N_9505);
nor U10890 (N_10890,N_9396,N_9649);
nor U10891 (N_10891,N_9976,N_9503);
nand U10892 (N_10892,N_9715,N_9490);
nand U10893 (N_10893,N_9869,N_9938);
xor U10894 (N_10894,N_9412,N_9369);
nor U10895 (N_10895,N_9363,N_9598);
xnor U10896 (N_10896,N_9760,N_9428);
nand U10897 (N_10897,N_9091,N_9749);
nor U10898 (N_10898,N_9602,N_9654);
nand U10899 (N_10899,N_9469,N_9889);
and U10900 (N_10900,N_9458,N_9797);
or U10901 (N_10901,N_9069,N_9868);
xnor U10902 (N_10902,N_9871,N_9225);
nand U10903 (N_10903,N_9617,N_9764);
nor U10904 (N_10904,N_9078,N_9396);
or U10905 (N_10905,N_9993,N_9162);
or U10906 (N_10906,N_9062,N_9658);
nor U10907 (N_10907,N_9367,N_9592);
and U10908 (N_10908,N_9501,N_9883);
nand U10909 (N_10909,N_9195,N_9555);
or U10910 (N_10910,N_9249,N_9184);
nand U10911 (N_10911,N_9826,N_9420);
nor U10912 (N_10912,N_9173,N_9137);
xnor U10913 (N_10913,N_9711,N_9333);
or U10914 (N_10914,N_9295,N_9030);
or U10915 (N_10915,N_9745,N_9306);
nand U10916 (N_10916,N_9372,N_9160);
nand U10917 (N_10917,N_9271,N_9486);
nor U10918 (N_10918,N_9745,N_9809);
nor U10919 (N_10919,N_9194,N_9875);
and U10920 (N_10920,N_9092,N_9233);
or U10921 (N_10921,N_9137,N_9121);
or U10922 (N_10922,N_9395,N_9124);
nor U10923 (N_10923,N_9329,N_9076);
xor U10924 (N_10924,N_9288,N_9075);
or U10925 (N_10925,N_9804,N_9596);
or U10926 (N_10926,N_9257,N_9633);
nand U10927 (N_10927,N_9087,N_9015);
and U10928 (N_10928,N_9615,N_9604);
xnor U10929 (N_10929,N_9339,N_9691);
or U10930 (N_10930,N_9827,N_9799);
xor U10931 (N_10931,N_9740,N_9346);
xor U10932 (N_10932,N_9140,N_9586);
nor U10933 (N_10933,N_9780,N_9696);
and U10934 (N_10934,N_9090,N_9813);
nand U10935 (N_10935,N_9570,N_9425);
nand U10936 (N_10936,N_9835,N_9259);
or U10937 (N_10937,N_9542,N_9610);
nand U10938 (N_10938,N_9208,N_9465);
xnor U10939 (N_10939,N_9451,N_9761);
and U10940 (N_10940,N_9966,N_9289);
nor U10941 (N_10941,N_9738,N_9836);
and U10942 (N_10942,N_9289,N_9462);
and U10943 (N_10943,N_9841,N_9443);
xnor U10944 (N_10944,N_9036,N_9429);
and U10945 (N_10945,N_9656,N_9937);
or U10946 (N_10946,N_9313,N_9390);
or U10947 (N_10947,N_9491,N_9622);
xor U10948 (N_10948,N_9963,N_9823);
nand U10949 (N_10949,N_9663,N_9704);
and U10950 (N_10950,N_9485,N_9576);
nor U10951 (N_10951,N_9457,N_9736);
and U10952 (N_10952,N_9032,N_9508);
and U10953 (N_10953,N_9195,N_9690);
and U10954 (N_10954,N_9853,N_9765);
or U10955 (N_10955,N_9873,N_9920);
xnor U10956 (N_10956,N_9478,N_9370);
nand U10957 (N_10957,N_9053,N_9561);
nor U10958 (N_10958,N_9619,N_9162);
nand U10959 (N_10959,N_9559,N_9898);
xnor U10960 (N_10960,N_9546,N_9675);
nand U10961 (N_10961,N_9094,N_9780);
and U10962 (N_10962,N_9533,N_9850);
xnor U10963 (N_10963,N_9317,N_9310);
xnor U10964 (N_10964,N_9488,N_9354);
nand U10965 (N_10965,N_9791,N_9978);
xor U10966 (N_10966,N_9658,N_9305);
or U10967 (N_10967,N_9659,N_9844);
xor U10968 (N_10968,N_9309,N_9293);
or U10969 (N_10969,N_9906,N_9093);
xor U10970 (N_10970,N_9075,N_9039);
nand U10971 (N_10971,N_9731,N_9638);
xor U10972 (N_10972,N_9248,N_9591);
and U10973 (N_10973,N_9262,N_9077);
nand U10974 (N_10974,N_9352,N_9781);
nand U10975 (N_10975,N_9799,N_9342);
nor U10976 (N_10976,N_9860,N_9012);
nand U10977 (N_10977,N_9646,N_9923);
nor U10978 (N_10978,N_9738,N_9742);
xnor U10979 (N_10979,N_9911,N_9153);
xnor U10980 (N_10980,N_9311,N_9135);
nand U10981 (N_10981,N_9803,N_9642);
nand U10982 (N_10982,N_9670,N_9315);
xnor U10983 (N_10983,N_9157,N_9864);
or U10984 (N_10984,N_9994,N_9051);
xnor U10985 (N_10985,N_9446,N_9842);
xnor U10986 (N_10986,N_9128,N_9750);
or U10987 (N_10987,N_9617,N_9167);
nand U10988 (N_10988,N_9720,N_9431);
xor U10989 (N_10989,N_9838,N_9958);
nand U10990 (N_10990,N_9814,N_9140);
xor U10991 (N_10991,N_9380,N_9236);
or U10992 (N_10992,N_9483,N_9826);
or U10993 (N_10993,N_9408,N_9311);
and U10994 (N_10994,N_9410,N_9225);
or U10995 (N_10995,N_9562,N_9519);
and U10996 (N_10996,N_9803,N_9584);
and U10997 (N_10997,N_9499,N_9990);
or U10998 (N_10998,N_9017,N_9485);
nand U10999 (N_10999,N_9086,N_9377);
nor U11000 (N_11000,N_10406,N_10095);
nand U11001 (N_11001,N_10690,N_10976);
and U11002 (N_11002,N_10045,N_10570);
nand U11003 (N_11003,N_10751,N_10325);
nand U11004 (N_11004,N_10285,N_10730);
xor U11005 (N_11005,N_10000,N_10146);
and U11006 (N_11006,N_10495,N_10858);
nor U11007 (N_11007,N_10636,N_10100);
or U11008 (N_11008,N_10800,N_10519);
nor U11009 (N_11009,N_10958,N_10318);
nor U11010 (N_11010,N_10569,N_10719);
xor U11011 (N_11011,N_10423,N_10142);
xor U11012 (N_11012,N_10249,N_10979);
nor U11013 (N_11013,N_10471,N_10481);
nand U11014 (N_11014,N_10524,N_10301);
and U11015 (N_11015,N_10252,N_10606);
nor U11016 (N_11016,N_10724,N_10357);
or U11017 (N_11017,N_10314,N_10411);
or U11018 (N_11018,N_10040,N_10974);
nand U11019 (N_11019,N_10163,N_10205);
nand U11020 (N_11020,N_10176,N_10831);
xor U11021 (N_11021,N_10064,N_10628);
nor U11022 (N_11022,N_10919,N_10910);
or U11023 (N_11023,N_10257,N_10386);
or U11024 (N_11024,N_10713,N_10230);
nand U11025 (N_11025,N_10262,N_10487);
xor U11026 (N_11026,N_10592,N_10439);
xor U11027 (N_11027,N_10180,N_10246);
and U11028 (N_11028,N_10173,N_10295);
nand U11029 (N_11029,N_10920,N_10110);
or U11030 (N_11030,N_10348,N_10824);
or U11031 (N_11031,N_10984,N_10201);
or U11032 (N_11032,N_10617,N_10154);
or U11033 (N_11033,N_10827,N_10161);
xor U11034 (N_11034,N_10632,N_10311);
nor U11035 (N_11035,N_10897,N_10305);
and U11036 (N_11036,N_10403,N_10344);
xor U11037 (N_11037,N_10714,N_10964);
nor U11038 (N_11038,N_10150,N_10124);
nand U11039 (N_11039,N_10275,N_10589);
and U11040 (N_11040,N_10613,N_10598);
nand U11041 (N_11041,N_10806,N_10511);
nand U11042 (N_11042,N_10611,N_10351);
and U11043 (N_11043,N_10336,N_10343);
xor U11044 (N_11044,N_10122,N_10946);
nor U11045 (N_11045,N_10623,N_10172);
nor U11046 (N_11046,N_10650,N_10680);
and U11047 (N_11047,N_10737,N_10326);
and U11048 (N_11048,N_10260,N_10629);
xnor U11049 (N_11049,N_10833,N_10277);
xnor U11050 (N_11050,N_10312,N_10470);
nand U11051 (N_11051,N_10459,N_10744);
xor U11052 (N_11052,N_10716,N_10004);
and U11053 (N_11053,N_10847,N_10079);
and U11054 (N_11054,N_10171,N_10672);
and U11055 (N_11055,N_10290,N_10155);
xnor U11056 (N_11056,N_10681,N_10178);
or U11057 (N_11057,N_10810,N_10400);
xor U11058 (N_11058,N_10783,N_10540);
or U11059 (N_11059,N_10300,N_10030);
xnor U11060 (N_11060,N_10961,N_10039);
xor U11061 (N_11061,N_10588,N_10826);
or U11062 (N_11062,N_10885,N_10691);
nand U11063 (N_11063,N_10354,N_10864);
xor U11064 (N_11064,N_10571,N_10269);
xnor U11065 (N_11065,N_10157,N_10425);
and U11066 (N_11066,N_10838,N_10693);
or U11067 (N_11067,N_10056,N_10368);
and U11068 (N_11068,N_10767,N_10947);
nor U11069 (N_11069,N_10139,N_10073);
nor U11070 (N_11070,N_10355,N_10208);
xnor U11071 (N_11071,N_10795,N_10328);
or U11072 (N_11072,N_10408,N_10583);
or U11073 (N_11073,N_10273,N_10983);
and U11074 (N_11074,N_10772,N_10720);
nand U11075 (N_11075,N_10440,N_10447);
and U11076 (N_11076,N_10182,N_10526);
or U11077 (N_11077,N_10652,N_10130);
nand U11078 (N_11078,N_10011,N_10010);
nand U11079 (N_11079,N_10705,N_10510);
xor U11080 (N_11080,N_10552,N_10942);
nand U11081 (N_11081,N_10229,N_10528);
nor U11082 (N_11082,N_10417,N_10683);
or U11083 (N_11083,N_10508,N_10771);
nor U11084 (N_11084,N_10382,N_10203);
nor U11085 (N_11085,N_10574,N_10840);
nor U11086 (N_11086,N_10981,N_10245);
xnor U11087 (N_11087,N_10754,N_10679);
nor U11088 (N_11088,N_10472,N_10414);
nor U11089 (N_11089,N_10206,N_10333);
and U11090 (N_11090,N_10863,N_10215);
nor U11091 (N_11091,N_10279,N_10909);
or U11092 (N_11092,N_10190,N_10120);
nand U11093 (N_11093,N_10950,N_10373);
and U11094 (N_11094,N_10189,N_10776);
or U11095 (N_11095,N_10980,N_10107);
and U11096 (N_11096,N_10993,N_10389);
nor U11097 (N_11097,N_10242,N_10653);
and U11098 (N_11098,N_10620,N_10894);
or U11099 (N_11099,N_10335,N_10835);
xnor U11100 (N_11100,N_10594,N_10543);
or U11101 (N_11101,N_10216,N_10538);
xor U11102 (N_11102,N_10012,N_10953);
and U11103 (N_11103,N_10119,N_10480);
or U11104 (N_11104,N_10711,N_10868);
and U11105 (N_11105,N_10449,N_10627);
nor U11106 (N_11106,N_10019,N_10654);
and U11107 (N_11107,N_10086,N_10071);
xnor U11108 (N_11108,N_10427,N_10151);
or U11109 (N_11109,N_10126,N_10074);
xnor U11110 (N_11110,N_10226,N_10371);
or U11111 (N_11111,N_10225,N_10726);
or U11112 (N_11112,N_10531,N_10936);
xor U11113 (N_11113,N_10890,N_10084);
or U11114 (N_11114,N_10456,N_10322);
nor U11115 (N_11115,N_10873,N_10133);
xor U11116 (N_11116,N_10689,N_10550);
nor U11117 (N_11117,N_10584,N_10553);
nand U11118 (N_11118,N_10777,N_10548);
or U11119 (N_11119,N_10736,N_10916);
xor U11120 (N_11120,N_10972,N_10391);
nand U11121 (N_11121,N_10198,N_10413);
nand U11122 (N_11122,N_10419,N_10676);
nor U11123 (N_11123,N_10259,N_10340);
nand U11124 (N_11124,N_10903,N_10963);
nor U11125 (N_11125,N_10310,N_10365);
xor U11126 (N_11126,N_10687,N_10763);
nand U11127 (N_11127,N_10135,N_10614);
and U11128 (N_11128,N_10610,N_10888);
xor U11129 (N_11129,N_10153,N_10655);
nor U11130 (N_11130,N_10970,N_10102);
and U11131 (N_11131,N_10374,N_10227);
nor U11132 (N_11132,N_10127,N_10814);
xnor U11133 (N_11133,N_10448,N_10590);
nand U11134 (N_11134,N_10765,N_10708);
or U11135 (N_11135,N_10179,N_10609);
and U11136 (N_11136,N_10812,N_10501);
nor U11137 (N_11137,N_10643,N_10458);
nor U11138 (N_11138,N_10282,N_10394);
or U11139 (N_11139,N_10067,N_10433);
and U11140 (N_11140,N_10346,N_10364);
and U11141 (N_11141,N_10671,N_10383);
xnor U11142 (N_11142,N_10995,N_10410);
nand U11143 (N_11143,N_10384,N_10641);
nand U11144 (N_11144,N_10843,N_10759);
nor U11145 (N_11145,N_10867,N_10851);
xnor U11146 (N_11146,N_10774,N_10522);
nor U11147 (N_11147,N_10529,N_10779);
nor U11148 (N_11148,N_10061,N_10962);
nor U11149 (N_11149,N_10017,N_10234);
nor U11150 (N_11150,N_10829,N_10455);
or U11151 (N_11151,N_10306,N_10619);
xnor U11152 (N_11152,N_10228,N_10175);
and U11153 (N_11153,N_10323,N_10985);
nor U11154 (N_11154,N_10006,N_10339);
xor U11155 (N_11155,N_10872,N_10461);
xor U11156 (N_11156,N_10880,N_10618);
xor U11157 (N_11157,N_10463,N_10784);
nand U11158 (N_11158,N_10760,N_10802);
nand U11159 (N_11159,N_10454,N_10482);
nor U11160 (N_11160,N_10442,N_10268);
nor U11161 (N_11161,N_10565,N_10852);
nor U11162 (N_11162,N_10005,N_10334);
and U11163 (N_11163,N_10430,N_10659);
or U11164 (N_11164,N_10089,N_10352);
and U11165 (N_11165,N_10445,N_10794);
nor U11166 (N_11166,N_10140,N_10360);
and U11167 (N_11167,N_10008,N_10068);
nand U11168 (N_11168,N_10533,N_10256);
xor U11169 (N_11169,N_10271,N_10184);
and U11170 (N_11170,N_10299,N_10270);
nand U11171 (N_11171,N_10399,N_10181);
and U11172 (N_11172,N_10546,N_10350);
nor U11173 (N_11173,N_10707,N_10786);
xor U11174 (N_11174,N_10202,N_10992);
xor U11175 (N_11175,N_10839,N_10670);
nand U11176 (N_11176,N_10889,N_10881);
and U11177 (N_11177,N_10093,N_10506);
nand U11178 (N_11178,N_10212,N_10823);
or U11179 (N_11179,N_10302,N_10345);
nand U11180 (N_11180,N_10072,N_10063);
and U11181 (N_11181,N_10393,N_10315);
xnor U11182 (N_11182,N_10168,N_10855);
and U11183 (N_11183,N_10421,N_10809);
nor U11184 (N_11184,N_10044,N_10735);
and U11185 (N_11185,N_10258,N_10453);
or U11186 (N_11186,N_10948,N_10284);
xnor U11187 (N_11187,N_10832,N_10055);
or U11188 (N_11188,N_10576,N_10324);
or U11189 (N_11189,N_10604,N_10341);
or U11190 (N_11190,N_10090,N_10381);
nor U11191 (N_11191,N_10804,N_10537);
xnor U11192 (N_11192,N_10267,N_10597);
xnor U11193 (N_11193,N_10605,N_10177);
nand U11194 (N_11194,N_10541,N_10775);
or U11195 (N_11195,N_10990,N_10952);
or U11196 (N_11196,N_10684,N_10498);
or U11197 (N_11197,N_10291,N_10549);
nor U11198 (N_11198,N_10485,N_10050);
or U11199 (N_11199,N_10036,N_10398);
nand U11200 (N_11200,N_10435,N_10704);
xor U11201 (N_11201,N_10596,N_10927);
nor U11202 (N_11202,N_10288,N_10327);
or U11203 (N_11203,N_10758,N_10562);
xnor U11204 (N_11204,N_10642,N_10977);
nand U11205 (N_11205,N_10307,N_10219);
xor U11206 (N_11206,N_10145,N_10276);
xor U11207 (N_11207,N_10504,N_10418);
or U11208 (N_11208,N_10075,N_10821);
nor U11209 (N_11209,N_10356,N_10287);
nand U11210 (N_11210,N_10105,N_10768);
nand U11211 (N_11211,N_10038,N_10217);
nor U11212 (N_11212,N_10791,N_10536);
nand U11213 (N_11213,N_10298,N_10405);
or U11214 (N_11214,N_10465,N_10018);
nand U11215 (N_11215,N_10696,N_10164);
xor U11216 (N_11216,N_10294,N_10507);
or U11217 (N_11217,N_10026,N_10196);
xor U11218 (N_11218,N_10853,N_10372);
nor U11219 (N_11219,N_10192,N_10367);
nand U11220 (N_11220,N_10998,N_10525);
or U11221 (N_11221,N_10865,N_10033);
nor U11222 (N_11222,N_10437,N_10043);
or U11223 (N_11223,N_10928,N_10875);
and U11224 (N_11224,N_10789,N_10624);
nand U11225 (N_11225,N_10505,N_10692);
nand U11226 (N_11226,N_10057,N_10370);
or U11227 (N_11227,N_10466,N_10631);
and U11228 (N_11228,N_10931,N_10296);
nand U11229 (N_11229,N_10429,N_10003);
and U11230 (N_11230,N_10994,N_10309);
and U11231 (N_11231,N_10669,N_10160);
and U11232 (N_11232,N_10109,N_10441);
nand U11233 (N_11233,N_10493,N_10673);
nand U11234 (N_11234,N_10224,N_10113);
or U11235 (N_11235,N_10599,N_10630);
xor U11236 (N_11236,N_10921,N_10479);
xnor U11237 (N_11237,N_10392,N_10603);
and U11238 (N_11238,N_10060,N_10143);
xor U11239 (N_11239,N_10283,N_10042);
xor U11240 (N_11240,N_10884,N_10460);
nand U11241 (N_11241,N_10407,N_10059);
xnor U11242 (N_11242,N_10527,N_10280);
or U11243 (N_11243,N_10940,N_10462);
or U11244 (N_11244,N_10807,N_10420);
xor U11245 (N_11245,N_10165,N_10330);
or U11246 (N_11246,N_10424,N_10578);
or U11247 (N_11247,N_10523,N_10248);
nor U11248 (N_11248,N_10490,N_10475);
nor U11249 (N_11249,N_10697,N_10808);
xnor U11250 (N_11250,N_10752,N_10729);
and U11251 (N_11251,N_10634,N_10366);
and U11252 (N_11252,N_10024,N_10710);
and U11253 (N_11253,N_10762,N_10907);
nand U11254 (N_11254,N_10815,N_10937);
xor U11255 (N_11255,N_10223,N_10787);
and U11256 (N_11256,N_10728,N_10349);
nand U11257 (N_11257,N_10002,N_10415);
xnor U11258 (N_11258,N_10949,N_10148);
xnor U11259 (N_11259,N_10938,N_10987);
xor U11260 (N_11260,N_10092,N_10635);
xnor U11261 (N_11261,N_10069,N_10542);
or U11262 (N_11262,N_10944,N_10723);
xnor U11263 (N_11263,N_10664,N_10138);
nor U11264 (N_11264,N_10820,N_10401);
xor U11265 (N_11265,N_10685,N_10021);
nor U11266 (N_11266,N_10756,N_10099);
nand U11267 (N_11267,N_10222,N_10796);
and U11268 (N_11268,N_10207,N_10123);
xnor U11269 (N_11269,N_10982,N_10934);
xnor U11270 (N_11270,N_10845,N_10753);
nand U11271 (N_11271,N_10112,N_10286);
nor U11272 (N_11272,N_10353,N_10313);
or U11273 (N_11273,N_10239,N_10563);
or U11274 (N_11274,N_10811,N_10255);
or U11275 (N_11275,N_10149,N_10443);
xor U11276 (N_11276,N_10929,N_10377);
or U11277 (N_11277,N_10049,N_10051);
nor U11278 (N_11278,N_10261,N_10699);
nor U11279 (N_11279,N_10925,N_10639);
nor U11280 (N_11280,N_10106,N_10220);
and U11281 (N_11281,N_10695,N_10530);
nor U11282 (N_11282,N_10798,N_10830);
nor U11283 (N_11283,N_10098,N_10478);
xor U11284 (N_11284,N_10854,N_10491);
nor U11285 (N_11285,N_10877,N_10602);
nand U11286 (N_11286,N_10745,N_10580);
xor U11287 (N_11287,N_10272,N_10361);
nor U11288 (N_11288,N_10973,N_10819);
nor U11289 (N_11289,N_10083,N_10503);
xnor U11290 (N_11290,N_10121,N_10954);
nand U11291 (N_11291,N_10579,N_10878);
nor U11292 (N_11292,N_10734,N_10144);
or U11293 (N_11293,N_10933,N_10882);
or U11294 (N_11294,N_10379,N_10500);
nor U11295 (N_11295,N_10476,N_10134);
xor U11296 (N_11296,N_10675,N_10761);
and U11297 (N_11297,N_10651,N_10790);
nand U11298 (N_11298,N_10674,N_10887);
and U11299 (N_11299,N_10721,N_10496);
or U11300 (N_11300,N_10081,N_10387);
xnor U11301 (N_11301,N_10231,N_10788);
xor U11302 (N_11302,N_10846,N_10125);
and U11303 (N_11303,N_10514,N_10739);
nand U11304 (N_11304,N_10428,N_10661);
nor U11305 (N_11305,N_10186,N_10844);
xor U11306 (N_11306,N_10557,N_10930);
nor U11307 (N_11307,N_10725,N_10905);
nand U11308 (N_11308,N_10660,N_10015);
and U11309 (N_11309,N_10385,N_10515);
nor U11310 (N_11310,N_10715,N_10782);
xor U11311 (N_11311,N_10263,N_10922);
nand U11312 (N_11312,N_10822,N_10971);
xor U11313 (N_11313,N_10091,N_10532);
or U11314 (N_11314,N_10321,N_10567);
or U11315 (N_11315,N_10062,N_10156);
and U11316 (N_11316,N_10213,N_10132);
nand U11317 (N_11317,N_10438,N_10862);
nor U11318 (N_11318,N_10170,N_10240);
nand U11319 (N_11319,N_10935,N_10101);
xnor U11320 (N_11320,N_10757,N_10876);
or U11321 (N_11321,N_10332,N_10347);
xnor U11322 (N_11322,N_10913,N_10253);
xnor U11323 (N_11323,N_10717,N_10362);
or U11324 (N_11324,N_10022,N_10577);
nand U11325 (N_11325,N_10899,N_10615);
xor U11326 (N_11326,N_10009,N_10238);
nand U11327 (N_11327,N_10568,N_10686);
or U11328 (N_11328,N_10559,N_10870);
and U11329 (N_11329,N_10886,N_10191);
or U11330 (N_11330,N_10509,N_10402);
nand U11331 (N_11331,N_10077,N_10426);
or U11332 (N_11332,N_10581,N_10035);
nor U11333 (N_11333,N_10195,N_10029);
nand U11334 (N_11334,N_10965,N_10116);
or U11335 (N_11335,N_10545,N_10896);
or U11336 (N_11336,N_10560,N_10197);
nor U11337 (N_11337,N_10633,N_10939);
nor U11338 (N_11338,N_10743,N_10956);
nand U11339 (N_11339,N_10989,N_10667);
nand U11340 (N_11340,N_10945,N_10128);
and U11341 (N_11341,N_10103,N_10169);
xnor U11342 (N_11342,N_10593,N_10600);
nand U11343 (N_11343,N_10975,N_10432);
xnor U11344 (N_11344,N_10444,N_10078);
nor U11345 (N_11345,N_10801,N_10250);
or U11346 (N_11346,N_10741,N_10167);
or U11347 (N_11347,N_10712,N_10988);
xnor U11348 (N_11348,N_10917,N_10718);
and U11349 (N_11349,N_10722,N_10278);
nor U11350 (N_11350,N_10467,N_10727);
and U11351 (N_11351,N_10129,N_10037);
nand U11352 (N_11352,N_10678,N_10337);
and U11353 (N_11353,N_10085,N_10236);
and U11354 (N_11354,N_10117,N_10521);
and U11355 (N_11355,N_10211,N_10625);
nand U11356 (N_11356,N_10047,N_10969);
nor U11357 (N_11357,N_10986,N_10233);
xnor U11358 (N_11358,N_10999,N_10032);
nor U11359 (N_11359,N_10702,N_10422);
xnor U11360 (N_11360,N_10070,N_10014);
and U11361 (N_11361,N_10204,N_10094);
or U11362 (N_11362,N_10595,N_10484);
nor U11363 (N_11363,N_10662,N_10648);
nand U11364 (N_11364,N_10547,N_10968);
and U11365 (N_11365,N_10647,N_10572);
or U11366 (N_11366,N_10573,N_10621);
nor U11367 (N_11367,N_10665,N_10740);
or U11368 (N_11368,N_10911,N_10668);
and U11369 (N_11369,N_10781,N_10477);
xnor U11370 (N_11370,N_10817,N_10380);
and U11371 (N_11371,N_10450,N_10431);
or U11372 (N_11372,N_10320,N_10612);
and U11373 (N_11373,N_10778,N_10898);
xnor U11374 (N_11374,N_10108,N_10409);
nand U11375 (N_11375,N_10793,N_10601);
nor U11376 (N_11376,N_10825,N_10001);
or U11377 (N_11377,N_10303,N_10805);
and U11378 (N_11378,N_10656,N_10369);
and U11379 (N_11379,N_10906,N_10141);
nor U11380 (N_11380,N_10749,N_10046);
and U11381 (N_11381,N_10908,N_10193);
nand U11382 (N_11382,N_10658,N_10232);
or U11383 (N_11383,N_10304,N_10358);
and U11384 (N_11384,N_10857,N_10566);
xnor U11385 (N_11385,N_10111,N_10816);
and U11386 (N_11386,N_10616,N_10048);
and U11387 (N_11387,N_10732,N_10554);
nand U11388 (N_11388,N_10096,N_10978);
xnor U11389 (N_11389,N_10516,N_10706);
or U11390 (N_11390,N_10766,N_10166);
xor U11391 (N_11391,N_10640,N_10649);
nor U11392 (N_11392,N_10136,N_10194);
nand U11393 (N_11393,N_10866,N_10746);
and U11394 (N_11394,N_10742,N_10188);
xor U11395 (N_11395,N_10152,N_10359);
nor U11396 (N_11396,N_10066,N_10274);
and U11397 (N_11397,N_10265,N_10183);
nand U11398 (N_11398,N_10915,N_10464);
and U11399 (N_11399,N_10446,N_10874);
and U11400 (N_11400,N_10199,N_10544);
xor U11401 (N_11401,N_10850,N_10058);
xor U11402 (N_11402,N_10375,N_10137);
nand U11403 (N_11403,N_10813,N_10308);
or U11404 (N_11404,N_10007,N_10241);
nor U11405 (N_11405,N_10488,N_10991);
and U11406 (N_11406,N_10243,N_10080);
xnor U11407 (N_11407,N_10281,N_10967);
nor U11408 (N_11408,N_10837,N_10396);
or U11409 (N_11409,N_10709,N_10034);
or U11410 (N_11410,N_10682,N_10292);
or U11411 (N_11411,N_10088,N_10028);
nor U11412 (N_11412,N_10518,N_10914);
or U11413 (N_11413,N_10904,N_10703);
nand U11414 (N_11414,N_10895,N_10586);
xor U11415 (N_11415,N_10097,N_10918);
and U11416 (N_11416,N_10317,N_10645);
xor U11417 (N_11417,N_10780,N_10483);
xnor U11418 (N_11418,N_10390,N_10582);
or U11419 (N_11419,N_10893,N_10297);
xnor U11420 (N_11420,N_10688,N_10966);
nor U11421 (N_11421,N_10797,N_10803);
nand U11422 (N_11422,N_10879,N_10535);
nand U11423 (N_11423,N_10841,N_10053);
nand U11424 (N_11424,N_10502,N_10955);
nand U11425 (N_11425,N_10395,N_10943);
xor U11426 (N_11426,N_10869,N_10264);
xnor U11427 (N_11427,N_10469,N_10836);
and U11428 (N_11428,N_10118,N_10701);
or U11429 (N_11429,N_10926,N_10663);
or U11430 (N_11430,N_10247,N_10738);
nor U11431 (N_11431,N_10200,N_10534);
xor U11432 (N_11432,N_10266,N_10316);
nor U11433 (N_11433,N_10251,N_10891);
nor U11434 (N_11434,N_10082,N_10923);
or U11435 (N_11435,N_10871,N_10932);
nand U11436 (N_11436,N_10210,N_10436);
nand U11437 (N_11437,N_10342,N_10158);
and U11438 (N_11438,N_10025,N_10564);
and U11439 (N_11439,N_10052,N_10900);
xnor U11440 (N_11440,N_10376,N_10329);
and U11441 (N_11441,N_10856,N_10187);
and U11442 (N_11442,N_10677,N_10997);
nor U11443 (N_11443,N_10770,N_10700);
and U11444 (N_11444,N_10289,N_10551);
xnor U11445 (N_11445,N_10027,N_10497);
nand U11446 (N_11446,N_10792,N_10486);
nand U11447 (N_11447,N_10363,N_10147);
xnor U11448 (N_11448,N_10218,N_10694);
and U11449 (N_11449,N_10698,N_10912);
or U11450 (N_11450,N_10799,N_10941);
or U11451 (N_11451,N_10115,N_10773);
xnor U11452 (N_11452,N_10638,N_10474);
and U11453 (N_11453,N_10861,N_10517);
nor U11454 (N_11454,N_10499,N_10556);
nor U11455 (N_11455,N_10214,N_10404);
or U11456 (N_11456,N_10159,N_10860);
or U11457 (N_11457,N_10733,N_10416);
xnor U11458 (N_11458,N_10104,N_10608);
nor U11459 (N_11459,N_10031,N_10622);
nand U11460 (N_11460,N_10020,N_10492);
xor U11461 (N_11461,N_10174,N_10512);
or U11462 (N_11462,N_10254,N_10114);
nand U11463 (N_11463,N_10054,N_10644);
or U11464 (N_11464,N_10468,N_10646);
nor U11465 (N_11465,N_10747,N_10587);
and U11466 (N_11466,N_10087,N_10957);
nand U11467 (N_11467,N_10666,N_10293);
and U11468 (N_11468,N_10607,N_10657);
or U11469 (N_11469,N_10016,N_10473);
or U11470 (N_11470,N_10539,N_10065);
nand U11471 (N_11471,N_10818,N_10489);
and U11472 (N_11472,N_10828,N_10378);
and U11473 (N_11473,N_10023,N_10013);
nor U11474 (N_11474,N_10388,N_10842);
or U11475 (N_11475,N_10131,N_10561);
nand U11476 (N_11476,N_10750,N_10494);
xor U11477 (N_11477,N_10951,N_10331);
nor U11478 (N_11478,N_10235,N_10319);
xnor U11479 (N_11479,N_10626,N_10834);
nor U11480 (N_11480,N_10892,N_10769);
or U11481 (N_11481,N_10901,N_10185);
and U11482 (N_11482,N_10591,N_10076);
and U11483 (N_11483,N_10555,N_10520);
nand U11484 (N_11484,N_10960,N_10209);
nand U11485 (N_11485,N_10237,N_10451);
xnor U11486 (N_11486,N_10883,N_10755);
nand U11487 (N_11487,N_10513,N_10637);
nor U11488 (N_11488,N_10412,N_10558);
and U11489 (N_11489,N_10221,N_10434);
nand U11490 (N_11490,N_10748,N_10731);
and U11491 (N_11491,N_10924,N_10457);
nor U11492 (N_11492,N_10849,N_10575);
xnor U11493 (N_11493,N_10338,N_10162);
xor U11494 (N_11494,N_10902,N_10785);
nand U11495 (N_11495,N_10041,N_10996);
and U11496 (N_11496,N_10959,N_10859);
or U11497 (N_11497,N_10244,N_10764);
nand U11498 (N_11498,N_10585,N_10848);
xnor U11499 (N_11499,N_10452,N_10397);
and U11500 (N_11500,N_10933,N_10114);
and U11501 (N_11501,N_10380,N_10969);
xor U11502 (N_11502,N_10322,N_10833);
nand U11503 (N_11503,N_10604,N_10590);
nand U11504 (N_11504,N_10778,N_10215);
and U11505 (N_11505,N_10234,N_10719);
or U11506 (N_11506,N_10556,N_10352);
nor U11507 (N_11507,N_10406,N_10612);
xor U11508 (N_11508,N_10619,N_10339);
nor U11509 (N_11509,N_10399,N_10584);
xnor U11510 (N_11510,N_10015,N_10645);
or U11511 (N_11511,N_10234,N_10358);
and U11512 (N_11512,N_10973,N_10780);
nand U11513 (N_11513,N_10878,N_10002);
and U11514 (N_11514,N_10112,N_10029);
xnor U11515 (N_11515,N_10875,N_10003);
and U11516 (N_11516,N_10411,N_10187);
or U11517 (N_11517,N_10209,N_10313);
or U11518 (N_11518,N_10970,N_10701);
nand U11519 (N_11519,N_10999,N_10956);
nor U11520 (N_11520,N_10884,N_10644);
xor U11521 (N_11521,N_10555,N_10932);
or U11522 (N_11522,N_10411,N_10354);
nand U11523 (N_11523,N_10999,N_10587);
nand U11524 (N_11524,N_10777,N_10013);
or U11525 (N_11525,N_10702,N_10452);
xor U11526 (N_11526,N_10699,N_10563);
or U11527 (N_11527,N_10200,N_10023);
nand U11528 (N_11528,N_10523,N_10002);
and U11529 (N_11529,N_10498,N_10465);
or U11530 (N_11530,N_10086,N_10813);
or U11531 (N_11531,N_10550,N_10832);
nand U11532 (N_11532,N_10692,N_10611);
nor U11533 (N_11533,N_10759,N_10595);
and U11534 (N_11534,N_10008,N_10860);
and U11535 (N_11535,N_10199,N_10777);
or U11536 (N_11536,N_10321,N_10394);
nand U11537 (N_11537,N_10315,N_10301);
or U11538 (N_11538,N_10168,N_10784);
xnor U11539 (N_11539,N_10917,N_10318);
nand U11540 (N_11540,N_10395,N_10526);
xor U11541 (N_11541,N_10269,N_10716);
or U11542 (N_11542,N_10557,N_10236);
nor U11543 (N_11543,N_10530,N_10073);
nand U11544 (N_11544,N_10913,N_10040);
or U11545 (N_11545,N_10066,N_10131);
nand U11546 (N_11546,N_10590,N_10632);
and U11547 (N_11547,N_10546,N_10301);
or U11548 (N_11548,N_10665,N_10189);
nand U11549 (N_11549,N_10393,N_10510);
or U11550 (N_11550,N_10781,N_10279);
or U11551 (N_11551,N_10934,N_10830);
xor U11552 (N_11552,N_10341,N_10464);
xnor U11553 (N_11553,N_10011,N_10788);
and U11554 (N_11554,N_10225,N_10099);
and U11555 (N_11555,N_10915,N_10436);
xnor U11556 (N_11556,N_10187,N_10062);
and U11557 (N_11557,N_10609,N_10039);
nor U11558 (N_11558,N_10837,N_10548);
nor U11559 (N_11559,N_10604,N_10457);
xnor U11560 (N_11560,N_10031,N_10416);
and U11561 (N_11561,N_10060,N_10675);
nor U11562 (N_11562,N_10405,N_10333);
nand U11563 (N_11563,N_10199,N_10731);
nand U11564 (N_11564,N_10370,N_10082);
nand U11565 (N_11565,N_10399,N_10496);
xor U11566 (N_11566,N_10628,N_10363);
nor U11567 (N_11567,N_10463,N_10247);
xor U11568 (N_11568,N_10770,N_10008);
nor U11569 (N_11569,N_10160,N_10208);
and U11570 (N_11570,N_10808,N_10225);
xnor U11571 (N_11571,N_10163,N_10854);
or U11572 (N_11572,N_10854,N_10507);
nand U11573 (N_11573,N_10640,N_10473);
nand U11574 (N_11574,N_10270,N_10008);
xnor U11575 (N_11575,N_10555,N_10327);
or U11576 (N_11576,N_10667,N_10904);
nor U11577 (N_11577,N_10633,N_10509);
nor U11578 (N_11578,N_10352,N_10898);
xor U11579 (N_11579,N_10975,N_10266);
or U11580 (N_11580,N_10359,N_10791);
xor U11581 (N_11581,N_10620,N_10035);
and U11582 (N_11582,N_10637,N_10975);
nor U11583 (N_11583,N_10418,N_10980);
xnor U11584 (N_11584,N_10084,N_10437);
and U11585 (N_11585,N_10360,N_10805);
nand U11586 (N_11586,N_10239,N_10973);
or U11587 (N_11587,N_10335,N_10146);
nor U11588 (N_11588,N_10418,N_10829);
and U11589 (N_11589,N_10495,N_10173);
nor U11590 (N_11590,N_10528,N_10396);
nand U11591 (N_11591,N_10985,N_10724);
nor U11592 (N_11592,N_10578,N_10405);
xor U11593 (N_11593,N_10784,N_10966);
xor U11594 (N_11594,N_10609,N_10937);
xnor U11595 (N_11595,N_10368,N_10355);
and U11596 (N_11596,N_10062,N_10706);
nor U11597 (N_11597,N_10871,N_10839);
xnor U11598 (N_11598,N_10502,N_10052);
nand U11599 (N_11599,N_10684,N_10522);
nor U11600 (N_11600,N_10359,N_10952);
and U11601 (N_11601,N_10357,N_10747);
nor U11602 (N_11602,N_10804,N_10753);
xnor U11603 (N_11603,N_10413,N_10113);
and U11604 (N_11604,N_10363,N_10092);
or U11605 (N_11605,N_10512,N_10780);
nand U11606 (N_11606,N_10457,N_10705);
nand U11607 (N_11607,N_10822,N_10379);
or U11608 (N_11608,N_10716,N_10279);
nand U11609 (N_11609,N_10466,N_10739);
or U11610 (N_11610,N_10327,N_10600);
and U11611 (N_11611,N_10530,N_10379);
nand U11612 (N_11612,N_10858,N_10801);
nor U11613 (N_11613,N_10548,N_10009);
nor U11614 (N_11614,N_10225,N_10874);
nor U11615 (N_11615,N_10266,N_10403);
nor U11616 (N_11616,N_10957,N_10896);
xor U11617 (N_11617,N_10272,N_10112);
or U11618 (N_11618,N_10530,N_10130);
xor U11619 (N_11619,N_10140,N_10423);
nor U11620 (N_11620,N_10671,N_10973);
nor U11621 (N_11621,N_10127,N_10347);
and U11622 (N_11622,N_10598,N_10564);
nor U11623 (N_11623,N_10150,N_10278);
nor U11624 (N_11624,N_10379,N_10886);
or U11625 (N_11625,N_10917,N_10489);
nand U11626 (N_11626,N_10257,N_10913);
xnor U11627 (N_11627,N_10137,N_10395);
nor U11628 (N_11628,N_10607,N_10595);
or U11629 (N_11629,N_10114,N_10623);
nand U11630 (N_11630,N_10849,N_10271);
xnor U11631 (N_11631,N_10827,N_10124);
xor U11632 (N_11632,N_10191,N_10221);
nor U11633 (N_11633,N_10527,N_10535);
nand U11634 (N_11634,N_10112,N_10402);
xnor U11635 (N_11635,N_10855,N_10921);
xnor U11636 (N_11636,N_10968,N_10089);
and U11637 (N_11637,N_10559,N_10817);
nand U11638 (N_11638,N_10072,N_10008);
xor U11639 (N_11639,N_10976,N_10423);
xnor U11640 (N_11640,N_10639,N_10128);
nor U11641 (N_11641,N_10535,N_10433);
and U11642 (N_11642,N_10412,N_10022);
nor U11643 (N_11643,N_10705,N_10342);
nand U11644 (N_11644,N_10614,N_10928);
or U11645 (N_11645,N_10171,N_10358);
nand U11646 (N_11646,N_10177,N_10119);
xnor U11647 (N_11647,N_10320,N_10628);
xnor U11648 (N_11648,N_10964,N_10776);
xor U11649 (N_11649,N_10828,N_10191);
and U11650 (N_11650,N_10754,N_10254);
xnor U11651 (N_11651,N_10043,N_10853);
or U11652 (N_11652,N_10670,N_10359);
nor U11653 (N_11653,N_10772,N_10300);
nand U11654 (N_11654,N_10935,N_10860);
nand U11655 (N_11655,N_10927,N_10206);
or U11656 (N_11656,N_10474,N_10675);
xnor U11657 (N_11657,N_10216,N_10966);
nor U11658 (N_11658,N_10628,N_10197);
nand U11659 (N_11659,N_10806,N_10103);
xnor U11660 (N_11660,N_10590,N_10843);
nor U11661 (N_11661,N_10513,N_10924);
nand U11662 (N_11662,N_10802,N_10700);
nand U11663 (N_11663,N_10929,N_10512);
xor U11664 (N_11664,N_10058,N_10164);
nand U11665 (N_11665,N_10552,N_10492);
nand U11666 (N_11666,N_10558,N_10722);
or U11667 (N_11667,N_10400,N_10333);
xnor U11668 (N_11668,N_10428,N_10273);
nor U11669 (N_11669,N_10791,N_10465);
and U11670 (N_11670,N_10210,N_10843);
and U11671 (N_11671,N_10360,N_10923);
and U11672 (N_11672,N_10541,N_10999);
nand U11673 (N_11673,N_10407,N_10536);
or U11674 (N_11674,N_10331,N_10534);
xor U11675 (N_11675,N_10506,N_10713);
nand U11676 (N_11676,N_10505,N_10033);
nand U11677 (N_11677,N_10322,N_10898);
nand U11678 (N_11678,N_10873,N_10751);
xnor U11679 (N_11679,N_10098,N_10744);
nand U11680 (N_11680,N_10867,N_10336);
xnor U11681 (N_11681,N_10268,N_10348);
nand U11682 (N_11682,N_10122,N_10701);
or U11683 (N_11683,N_10659,N_10008);
nand U11684 (N_11684,N_10226,N_10140);
xnor U11685 (N_11685,N_10486,N_10964);
xnor U11686 (N_11686,N_10220,N_10636);
or U11687 (N_11687,N_10834,N_10907);
and U11688 (N_11688,N_10352,N_10348);
nand U11689 (N_11689,N_10233,N_10864);
xor U11690 (N_11690,N_10858,N_10766);
nor U11691 (N_11691,N_10881,N_10647);
and U11692 (N_11692,N_10016,N_10176);
xor U11693 (N_11693,N_10317,N_10162);
or U11694 (N_11694,N_10301,N_10466);
nand U11695 (N_11695,N_10954,N_10050);
xnor U11696 (N_11696,N_10924,N_10781);
nand U11697 (N_11697,N_10907,N_10949);
or U11698 (N_11698,N_10662,N_10639);
nor U11699 (N_11699,N_10249,N_10176);
xor U11700 (N_11700,N_10295,N_10999);
and U11701 (N_11701,N_10984,N_10963);
xor U11702 (N_11702,N_10863,N_10569);
nand U11703 (N_11703,N_10557,N_10069);
and U11704 (N_11704,N_10251,N_10127);
and U11705 (N_11705,N_10318,N_10530);
xnor U11706 (N_11706,N_10988,N_10674);
and U11707 (N_11707,N_10641,N_10962);
nand U11708 (N_11708,N_10856,N_10929);
nor U11709 (N_11709,N_10691,N_10686);
nand U11710 (N_11710,N_10552,N_10413);
or U11711 (N_11711,N_10485,N_10489);
xnor U11712 (N_11712,N_10066,N_10861);
nand U11713 (N_11713,N_10856,N_10688);
nor U11714 (N_11714,N_10776,N_10360);
or U11715 (N_11715,N_10182,N_10437);
and U11716 (N_11716,N_10723,N_10114);
or U11717 (N_11717,N_10149,N_10635);
xor U11718 (N_11718,N_10141,N_10558);
nor U11719 (N_11719,N_10758,N_10347);
xor U11720 (N_11720,N_10809,N_10001);
xor U11721 (N_11721,N_10121,N_10682);
nand U11722 (N_11722,N_10679,N_10315);
nor U11723 (N_11723,N_10478,N_10629);
or U11724 (N_11724,N_10108,N_10365);
nand U11725 (N_11725,N_10290,N_10594);
and U11726 (N_11726,N_10161,N_10426);
nand U11727 (N_11727,N_10422,N_10719);
or U11728 (N_11728,N_10983,N_10178);
or U11729 (N_11729,N_10387,N_10238);
and U11730 (N_11730,N_10047,N_10353);
and U11731 (N_11731,N_10883,N_10354);
xnor U11732 (N_11732,N_10898,N_10009);
nor U11733 (N_11733,N_10878,N_10265);
xnor U11734 (N_11734,N_10710,N_10651);
and U11735 (N_11735,N_10727,N_10693);
and U11736 (N_11736,N_10405,N_10618);
xnor U11737 (N_11737,N_10115,N_10599);
or U11738 (N_11738,N_10016,N_10584);
xnor U11739 (N_11739,N_10205,N_10517);
and U11740 (N_11740,N_10729,N_10911);
and U11741 (N_11741,N_10562,N_10170);
nand U11742 (N_11742,N_10796,N_10427);
xor U11743 (N_11743,N_10799,N_10249);
and U11744 (N_11744,N_10541,N_10314);
or U11745 (N_11745,N_10649,N_10972);
nor U11746 (N_11746,N_10291,N_10795);
xor U11747 (N_11747,N_10274,N_10797);
or U11748 (N_11748,N_10470,N_10466);
or U11749 (N_11749,N_10389,N_10093);
nor U11750 (N_11750,N_10560,N_10855);
xor U11751 (N_11751,N_10001,N_10564);
nand U11752 (N_11752,N_10197,N_10790);
nor U11753 (N_11753,N_10287,N_10887);
nor U11754 (N_11754,N_10859,N_10419);
nand U11755 (N_11755,N_10831,N_10951);
or U11756 (N_11756,N_10196,N_10986);
or U11757 (N_11757,N_10802,N_10068);
or U11758 (N_11758,N_10826,N_10468);
nand U11759 (N_11759,N_10709,N_10288);
and U11760 (N_11760,N_10722,N_10997);
nand U11761 (N_11761,N_10750,N_10094);
and U11762 (N_11762,N_10263,N_10763);
xor U11763 (N_11763,N_10951,N_10177);
and U11764 (N_11764,N_10788,N_10853);
xor U11765 (N_11765,N_10845,N_10267);
and U11766 (N_11766,N_10684,N_10255);
nand U11767 (N_11767,N_10635,N_10697);
nor U11768 (N_11768,N_10426,N_10167);
nor U11769 (N_11769,N_10722,N_10584);
nand U11770 (N_11770,N_10540,N_10388);
xnor U11771 (N_11771,N_10273,N_10386);
nand U11772 (N_11772,N_10887,N_10720);
xnor U11773 (N_11773,N_10420,N_10043);
nor U11774 (N_11774,N_10744,N_10087);
nand U11775 (N_11775,N_10920,N_10271);
nand U11776 (N_11776,N_10362,N_10970);
xnor U11777 (N_11777,N_10707,N_10458);
xor U11778 (N_11778,N_10647,N_10292);
or U11779 (N_11779,N_10468,N_10539);
xnor U11780 (N_11780,N_10700,N_10047);
nand U11781 (N_11781,N_10403,N_10684);
xnor U11782 (N_11782,N_10415,N_10907);
and U11783 (N_11783,N_10215,N_10577);
nor U11784 (N_11784,N_10669,N_10950);
nand U11785 (N_11785,N_10654,N_10791);
and U11786 (N_11786,N_10277,N_10805);
or U11787 (N_11787,N_10583,N_10927);
nand U11788 (N_11788,N_10652,N_10547);
nor U11789 (N_11789,N_10477,N_10894);
nor U11790 (N_11790,N_10815,N_10367);
or U11791 (N_11791,N_10603,N_10207);
or U11792 (N_11792,N_10422,N_10802);
nor U11793 (N_11793,N_10008,N_10537);
and U11794 (N_11794,N_10701,N_10312);
nor U11795 (N_11795,N_10284,N_10240);
nor U11796 (N_11796,N_10677,N_10015);
and U11797 (N_11797,N_10815,N_10644);
or U11798 (N_11798,N_10701,N_10328);
nand U11799 (N_11799,N_10928,N_10209);
and U11800 (N_11800,N_10430,N_10326);
and U11801 (N_11801,N_10450,N_10731);
or U11802 (N_11802,N_10607,N_10502);
nand U11803 (N_11803,N_10578,N_10921);
or U11804 (N_11804,N_10764,N_10310);
xnor U11805 (N_11805,N_10686,N_10875);
nor U11806 (N_11806,N_10236,N_10782);
nand U11807 (N_11807,N_10916,N_10073);
or U11808 (N_11808,N_10791,N_10161);
xor U11809 (N_11809,N_10049,N_10210);
xnor U11810 (N_11810,N_10093,N_10558);
and U11811 (N_11811,N_10332,N_10441);
and U11812 (N_11812,N_10110,N_10087);
nand U11813 (N_11813,N_10785,N_10030);
nor U11814 (N_11814,N_10876,N_10234);
nand U11815 (N_11815,N_10561,N_10271);
and U11816 (N_11816,N_10123,N_10842);
and U11817 (N_11817,N_10873,N_10884);
nand U11818 (N_11818,N_10526,N_10728);
and U11819 (N_11819,N_10246,N_10504);
nor U11820 (N_11820,N_10912,N_10034);
nor U11821 (N_11821,N_10233,N_10801);
nand U11822 (N_11822,N_10709,N_10061);
xnor U11823 (N_11823,N_10455,N_10987);
or U11824 (N_11824,N_10850,N_10993);
nand U11825 (N_11825,N_10240,N_10462);
nor U11826 (N_11826,N_10693,N_10114);
and U11827 (N_11827,N_10912,N_10500);
nand U11828 (N_11828,N_10957,N_10898);
nand U11829 (N_11829,N_10312,N_10505);
nor U11830 (N_11830,N_10184,N_10195);
nand U11831 (N_11831,N_10061,N_10893);
nand U11832 (N_11832,N_10059,N_10760);
and U11833 (N_11833,N_10591,N_10030);
or U11834 (N_11834,N_10563,N_10555);
xor U11835 (N_11835,N_10502,N_10074);
or U11836 (N_11836,N_10016,N_10153);
or U11837 (N_11837,N_10331,N_10683);
and U11838 (N_11838,N_10522,N_10596);
xor U11839 (N_11839,N_10174,N_10574);
and U11840 (N_11840,N_10719,N_10683);
nor U11841 (N_11841,N_10649,N_10351);
xnor U11842 (N_11842,N_10593,N_10134);
and U11843 (N_11843,N_10507,N_10518);
xnor U11844 (N_11844,N_10971,N_10926);
or U11845 (N_11845,N_10796,N_10343);
xor U11846 (N_11846,N_10225,N_10923);
and U11847 (N_11847,N_10047,N_10668);
or U11848 (N_11848,N_10425,N_10790);
nor U11849 (N_11849,N_10252,N_10571);
xor U11850 (N_11850,N_10255,N_10327);
nand U11851 (N_11851,N_10823,N_10414);
nand U11852 (N_11852,N_10787,N_10925);
and U11853 (N_11853,N_10283,N_10549);
nand U11854 (N_11854,N_10379,N_10197);
or U11855 (N_11855,N_10000,N_10551);
xor U11856 (N_11856,N_10764,N_10473);
and U11857 (N_11857,N_10143,N_10850);
or U11858 (N_11858,N_10999,N_10746);
nor U11859 (N_11859,N_10546,N_10314);
nor U11860 (N_11860,N_10844,N_10837);
xor U11861 (N_11861,N_10904,N_10785);
xnor U11862 (N_11862,N_10091,N_10551);
xnor U11863 (N_11863,N_10816,N_10568);
nand U11864 (N_11864,N_10413,N_10350);
or U11865 (N_11865,N_10368,N_10537);
nor U11866 (N_11866,N_10610,N_10801);
or U11867 (N_11867,N_10784,N_10531);
xnor U11868 (N_11868,N_10364,N_10197);
or U11869 (N_11869,N_10893,N_10127);
xnor U11870 (N_11870,N_10790,N_10349);
nor U11871 (N_11871,N_10229,N_10690);
and U11872 (N_11872,N_10042,N_10711);
nand U11873 (N_11873,N_10303,N_10975);
or U11874 (N_11874,N_10534,N_10427);
nand U11875 (N_11875,N_10234,N_10708);
nor U11876 (N_11876,N_10709,N_10243);
nor U11877 (N_11877,N_10668,N_10261);
xnor U11878 (N_11878,N_10523,N_10242);
and U11879 (N_11879,N_10030,N_10112);
nor U11880 (N_11880,N_10565,N_10119);
nor U11881 (N_11881,N_10957,N_10885);
nor U11882 (N_11882,N_10295,N_10762);
nand U11883 (N_11883,N_10836,N_10899);
xnor U11884 (N_11884,N_10573,N_10691);
and U11885 (N_11885,N_10485,N_10558);
and U11886 (N_11886,N_10836,N_10342);
xor U11887 (N_11887,N_10622,N_10953);
and U11888 (N_11888,N_10328,N_10481);
xor U11889 (N_11889,N_10451,N_10523);
and U11890 (N_11890,N_10161,N_10688);
or U11891 (N_11891,N_10778,N_10524);
nor U11892 (N_11892,N_10172,N_10297);
or U11893 (N_11893,N_10291,N_10804);
nor U11894 (N_11894,N_10985,N_10755);
nor U11895 (N_11895,N_10691,N_10034);
nand U11896 (N_11896,N_10191,N_10291);
nand U11897 (N_11897,N_10865,N_10075);
nand U11898 (N_11898,N_10777,N_10212);
or U11899 (N_11899,N_10330,N_10485);
nor U11900 (N_11900,N_10885,N_10743);
xor U11901 (N_11901,N_10411,N_10168);
or U11902 (N_11902,N_10798,N_10891);
or U11903 (N_11903,N_10995,N_10262);
nor U11904 (N_11904,N_10247,N_10908);
nor U11905 (N_11905,N_10443,N_10103);
xor U11906 (N_11906,N_10460,N_10389);
nor U11907 (N_11907,N_10680,N_10952);
or U11908 (N_11908,N_10274,N_10203);
and U11909 (N_11909,N_10879,N_10708);
and U11910 (N_11910,N_10728,N_10838);
nor U11911 (N_11911,N_10134,N_10737);
and U11912 (N_11912,N_10478,N_10555);
xnor U11913 (N_11913,N_10695,N_10440);
or U11914 (N_11914,N_10449,N_10880);
xnor U11915 (N_11915,N_10682,N_10540);
nor U11916 (N_11916,N_10931,N_10763);
or U11917 (N_11917,N_10844,N_10528);
nor U11918 (N_11918,N_10779,N_10158);
nand U11919 (N_11919,N_10702,N_10527);
nand U11920 (N_11920,N_10229,N_10649);
xor U11921 (N_11921,N_10873,N_10896);
or U11922 (N_11922,N_10331,N_10587);
nand U11923 (N_11923,N_10462,N_10877);
or U11924 (N_11924,N_10975,N_10217);
or U11925 (N_11925,N_10221,N_10324);
nor U11926 (N_11926,N_10182,N_10920);
nor U11927 (N_11927,N_10749,N_10908);
nand U11928 (N_11928,N_10883,N_10612);
or U11929 (N_11929,N_10715,N_10295);
or U11930 (N_11930,N_10218,N_10133);
nor U11931 (N_11931,N_10965,N_10033);
and U11932 (N_11932,N_10159,N_10271);
and U11933 (N_11933,N_10019,N_10343);
xor U11934 (N_11934,N_10810,N_10858);
xnor U11935 (N_11935,N_10532,N_10690);
or U11936 (N_11936,N_10123,N_10448);
nor U11937 (N_11937,N_10736,N_10958);
xor U11938 (N_11938,N_10783,N_10344);
nor U11939 (N_11939,N_10086,N_10403);
nand U11940 (N_11940,N_10602,N_10239);
nand U11941 (N_11941,N_10073,N_10876);
nor U11942 (N_11942,N_10320,N_10075);
nand U11943 (N_11943,N_10546,N_10083);
nand U11944 (N_11944,N_10329,N_10602);
or U11945 (N_11945,N_10275,N_10482);
or U11946 (N_11946,N_10175,N_10230);
and U11947 (N_11947,N_10693,N_10375);
xor U11948 (N_11948,N_10061,N_10695);
and U11949 (N_11949,N_10866,N_10417);
nor U11950 (N_11950,N_10958,N_10822);
and U11951 (N_11951,N_10597,N_10540);
or U11952 (N_11952,N_10700,N_10889);
xor U11953 (N_11953,N_10448,N_10230);
and U11954 (N_11954,N_10149,N_10366);
nor U11955 (N_11955,N_10620,N_10362);
nand U11956 (N_11956,N_10938,N_10252);
or U11957 (N_11957,N_10561,N_10846);
or U11958 (N_11958,N_10939,N_10634);
and U11959 (N_11959,N_10314,N_10934);
and U11960 (N_11960,N_10326,N_10684);
and U11961 (N_11961,N_10545,N_10465);
and U11962 (N_11962,N_10199,N_10000);
nand U11963 (N_11963,N_10607,N_10483);
nor U11964 (N_11964,N_10091,N_10754);
and U11965 (N_11965,N_10120,N_10025);
xor U11966 (N_11966,N_10454,N_10103);
and U11967 (N_11967,N_10648,N_10901);
nor U11968 (N_11968,N_10404,N_10695);
xor U11969 (N_11969,N_10997,N_10312);
nand U11970 (N_11970,N_10933,N_10695);
xnor U11971 (N_11971,N_10940,N_10965);
xor U11972 (N_11972,N_10551,N_10893);
xor U11973 (N_11973,N_10870,N_10524);
nand U11974 (N_11974,N_10252,N_10438);
nand U11975 (N_11975,N_10212,N_10473);
nor U11976 (N_11976,N_10359,N_10963);
xnor U11977 (N_11977,N_10292,N_10988);
xor U11978 (N_11978,N_10018,N_10008);
xnor U11979 (N_11979,N_10368,N_10311);
nand U11980 (N_11980,N_10769,N_10015);
xnor U11981 (N_11981,N_10728,N_10098);
or U11982 (N_11982,N_10341,N_10355);
or U11983 (N_11983,N_10334,N_10627);
and U11984 (N_11984,N_10415,N_10570);
nand U11985 (N_11985,N_10459,N_10076);
and U11986 (N_11986,N_10175,N_10400);
and U11987 (N_11987,N_10231,N_10809);
and U11988 (N_11988,N_10474,N_10486);
or U11989 (N_11989,N_10552,N_10050);
and U11990 (N_11990,N_10903,N_10286);
nor U11991 (N_11991,N_10681,N_10088);
nor U11992 (N_11992,N_10577,N_10091);
and U11993 (N_11993,N_10219,N_10837);
and U11994 (N_11994,N_10276,N_10421);
xor U11995 (N_11995,N_10551,N_10439);
or U11996 (N_11996,N_10017,N_10927);
nor U11997 (N_11997,N_10144,N_10041);
or U11998 (N_11998,N_10069,N_10602);
xnor U11999 (N_11999,N_10247,N_10024);
nor U12000 (N_12000,N_11518,N_11373);
xor U12001 (N_12001,N_11659,N_11288);
or U12002 (N_12002,N_11245,N_11845);
or U12003 (N_12003,N_11131,N_11662);
nor U12004 (N_12004,N_11834,N_11752);
nand U12005 (N_12005,N_11593,N_11560);
nand U12006 (N_12006,N_11940,N_11857);
and U12007 (N_12007,N_11991,N_11666);
nor U12008 (N_12008,N_11559,N_11856);
nand U12009 (N_12009,N_11722,N_11434);
nor U12010 (N_12010,N_11459,N_11596);
nand U12011 (N_12011,N_11212,N_11744);
xnor U12012 (N_12012,N_11531,N_11925);
nand U12013 (N_12013,N_11619,N_11575);
and U12014 (N_12014,N_11658,N_11720);
or U12015 (N_12015,N_11092,N_11929);
nor U12016 (N_12016,N_11431,N_11352);
and U12017 (N_12017,N_11934,N_11819);
nor U12018 (N_12018,N_11533,N_11871);
xnor U12019 (N_12019,N_11050,N_11168);
or U12020 (N_12020,N_11591,N_11792);
xnor U12021 (N_12021,N_11319,N_11858);
or U12022 (N_12022,N_11699,N_11051);
nand U12023 (N_12023,N_11182,N_11877);
xor U12024 (N_12024,N_11972,N_11968);
xnor U12025 (N_12025,N_11625,N_11414);
nand U12026 (N_12026,N_11797,N_11290);
nand U12027 (N_12027,N_11519,N_11029);
or U12028 (N_12028,N_11975,N_11402);
nand U12029 (N_12029,N_11813,N_11043);
and U12030 (N_12030,N_11692,N_11399);
and U12031 (N_12031,N_11375,N_11580);
nand U12032 (N_12032,N_11473,N_11527);
xnor U12033 (N_12033,N_11392,N_11380);
or U12034 (N_12034,N_11607,N_11757);
nand U12035 (N_12035,N_11472,N_11111);
nand U12036 (N_12036,N_11070,N_11069);
and U12037 (N_12037,N_11852,N_11046);
xnor U12038 (N_12038,N_11740,N_11210);
nand U12039 (N_12039,N_11851,N_11880);
or U12040 (N_12040,N_11027,N_11170);
or U12041 (N_12041,N_11995,N_11389);
xor U12042 (N_12042,N_11407,N_11208);
and U12043 (N_12043,N_11774,N_11983);
nand U12044 (N_12044,N_11644,N_11003);
nor U12045 (N_12045,N_11578,N_11935);
xor U12046 (N_12046,N_11450,N_11759);
and U12047 (N_12047,N_11861,N_11725);
and U12048 (N_12048,N_11639,N_11984);
or U12049 (N_12049,N_11259,N_11491);
xor U12050 (N_12050,N_11201,N_11299);
nor U12051 (N_12051,N_11276,N_11787);
xnor U12052 (N_12052,N_11839,N_11000);
or U12053 (N_12053,N_11501,N_11687);
or U12054 (N_12054,N_11180,N_11647);
nand U12055 (N_12055,N_11967,N_11097);
xor U12056 (N_12056,N_11040,N_11869);
or U12057 (N_12057,N_11715,N_11469);
xor U12058 (N_12058,N_11285,N_11360);
or U12059 (N_12059,N_11919,N_11308);
or U12060 (N_12060,N_11179,N_11166);
and U12061 (N_12061,N_11325,N_11635);
xor U12062 (N_12062,N_11783,N_11548);
nor U12063 (N_12063,N_11035,N_11994);
and U12064 (N_12064,N_11340,N_11897);
xnor U12065 (N_12065,N_11221,N_11159);
or U12066 (N_12066,N_11749,N_11911);
nor U12067 (N_12067,N_11028,N_11086);
nor U12068 (N_12068,N_11495,N_11354);
nor U12069 (N_12069,N_11363,N_11146);
nand U12070 (N_12070,N_11913,N_11423);
xnor U12071 (N_12071,N_11950,N_11653);
xnor U12072 (N_12072,N_11569,N_11095);
xnor U12073 (N_12073,N_11253,N_11899);
or U12074 (N_12074,N_11753,N_11160);
or U12075 (N_12075,N_11781,N_11885);
nand U12076 (N_12076,N_11891,N_11550);
nand U12077 (N_12077,N_11395,N_11551);
and U12078 (N_12078,N_11650,N_11597);
nor U12079 (N_12079,N_11264,N_11816);
or U12080 (N_12080,N_11741,N_11016);
nor U12081 (N_12081,N_11500,N_11280);
or U12082 (N_12082,N_11056,N_11019);
nor U12083 (N_12083,N_11467,N_11920);
xor U12084 (N_12084,N_11445,N_11075);
xor U12085 (N_12085,N_11694,N_11162);
or U12086 (N_12086,N_11383,N_11430);
xnor U12087 (N_12087,N_11735,N_11353);
xor U12088 (N_12088,N_11987,N_11145);
nand U12089 (N_12089,N_11704,N_11476);
nand U12090 (N_12090,N_11444,N_11368);
nor U12091 (N_12091,N_11660,N_11009);
or U12092 (N_12092,N_11717,N_11274);
and U12093 (N_12093,N_11388,N_11778);
or U12094 (N_12094,N_11125,N_11656);
xnor U12095 (N_12095,N_11840,N_11760);
or U12096 (N_12096,N_11788,N_11102);
or U12097 (N_12097,N_11679,N_11214);
and U12098 (N_12098,N_11317,N_11083);
and U12099 (N_12099,N_11942,N_11055);
xor U12100 (N_12100,N_11808,N_11232);
xnor U12101 (N_12101,N_11732,N_11057);
nor U12102 (N_12102,N_11693,N_11498);
and U12103 (N_12103,N_11215,N_11297);
nor U12104 (N_12104,N_11543,N_11842);
and U12105 (N_12105,N_11439,N_11361);
nand U12106 (N_12106,N_11119,N_11148);
and U12107 (N_12107,N_11268,N_11198);
and U12108 (N_12108,N_11990,N_11698);
nand U12109 (N_12109,N_11870,N_11697);
xor U12110 (N_12110,N_11184,N_11396);
and U12111 (N_12111,N_11526,N_11628);
nand U12112 (N_12112,N_11511,N_11785);
and U12113 (N_12113,N_11981,N_11709);
xnor U12114 (N_12114,N_11194,N_11178);
or U12115 (N_12115,N_11626,N_11806);
or U12116 (N_12116,N_11138,N_11471);
or U12117 (N_12117,N_11298,N_11181);
or U12118 (N_12118,N_11237,N_11553);
xnor U12119 (N_12119,N_11962,N_11712);
and U12120 (N_12120,N_11229,N_11376);
xor U12121 (N_12121,N_11961,N_11608);
xor U12122 (N_12122,N_11209,N_11127);
nand U12123 (N_12123,N_11505,N_11770);
nor U12124 (N_12124,N_11828,N_11204);
nand U12125 (N_12125,N_11163,N_11651);
or U12126 (N_12126,N_11943,N_11134);
xor U12127 (N_12127,N_11572,N_11969);
nor U12128 (N_12128,N_11584,N_11826);
nor U12129 (N_12129,N_11391,N_11303);
xnor U12130 (N_12130,N_11794,N_11520);
xnor U12131 (N_12131,N_11989,N_11137);
nand U12132 (N_12132,N_11780,N_11283);
and U12133 (N_12133,N_11509,N_11453);
and U12134 (N_12134,N_11873,N_11664);
and U12135 (N_12135,N_11507,N_11408);
nand U12136 (N_12136,N_11177,N_11084);
nand U12137 (N_12137,N_11986,N_11811);
nor U12138 (N_12138,N_11648,N_11410);
or U12139 (N_12139,N_11535,N_11196);
nand U12140 (N_12140,N_11844,N_11627);
nor U12141 (N_12141,N_11676,N_11827);
nor U12142 (N_12142,N_11490,N_11571);
and U12143 (N_12143,N_11203,N_11218);
and U12144 (N_12144,N_11510,N_11566);
nand U12145 (N_12145,N_11767,N_11089);
nand U12146 (N_12146,N_11066,N_11295);
or U12147 (N_12147,N_11678,N_11404);
nor U12148 (N_12148,N_11413,N_11405);
or U12149 (N_12149,N_11002,N_11073);
nor U12150 (N_12150,N_11104,N_11789);
or U12151 (N_12151,N_11773,N_11233);
or U12152 (N_12152,N_11377,N_11023);
xnor U12153 (N_12153,N_11928,N_11988);
or U12154 (N_12154,N_11492,N_11546);
nand U12155 (N_12155,N_11106,N_11195);
or U12156 (N_12156,N_11384,N_11764);
xor U12157 (N_12157,N_11949,N_11805);
and U12158 (N_12158,N_11031,N_11985);
or U12159 (N_12159,N_11085,N_11107);
xnor U12160 (N_12160,N_11174,N_11401);
and U12161 (N_12161,N_11830,N_11310);
xor U12162 (N_12162,N_11955,N_11927);
or U12163 (N_12163,N_11386,N_11745);
and U12164 (N_12164,N_11549,N_11618);
and U12165 (N_12165,N_11406,N_11677);
and U12166 (N_12166,N_11818,N_11153);
and U12167 (N_12167,N_11048,N_11442);
and U12168 (N_12168,N_11337,N_11585);
nand U12169 (N_12169,N_11613,N_11385);
nor U12170 (N_12170,N_11926,N_11393);
nand U12171 (N_12171,N_11436,N_11887);
xor U12172 (N_12172,N_11750,N_11790);
and U12173 (N_12173,N_11091,N_11358);
xor U12174 (N_12174,N_11640,N_11979);
or U12175 (N_12175,N_11341,N_11320);
nor U12176 (N_12176,N_11912,N_11165);
nand U12177 (N_12177,N_11971,N_11965);
and U12178 (N_12178,N_11631,N_11428);
or U12179 (N_12179,N_11344,N_11803);
nor U12180 (N_12180,N_11630,N_11945);
nor U12181 (N_12181,N_11737,N_11817);
nand U12182 (N_12182,N_11525,N_11530);
nor U12183 (N_12183,N_11485,N_11683);
nand U12184 (N_12184,N_11604,N_11192);
nor U12185 (N_12185,N_11700,N_11799);
and U12186 (N_12186,N_11742,N_11561);
xnor U12187 (N_12187,N_11282,N_11052);
and U12188 (N_12188,N_11641,N_11831);
nor U12189 (N_12189,N_11800,N_11574);
xnor U12190 (N_12190,N_11843,N_11915);
nor U12191 (N_12191,N_11123,N_11727);
xnor U12192 (N_12192,N_11802,N_11458);
and U12193 (N_12193,N_11503,N_11022);
and U12194 (N_12194,N_11748,N_11502);
nor U12195 (N_12195,N_11425,N_11364);
or U12196 (N_12196,N_11464,N_11810);
xor U12197 (N_12197,N_11959,N_11812);
and U12198 (N_12198,N_11768,N_11594);
xor U12199 (N_12199,N_11652,N_11848);
xnor U12200 (N_12200,N_11494,N_11415);
nand U12201 (N_12201,N_11226,N_11225);
or U12202 (N_12202,N_11815,N_11256);
nand U12203 (N_12203,N_11909,N_11087);
and U12204 (N_12204,N_11980,N_11524);
or U12205 (N_12205,N_11449,N_11854);
and U12206 (N_12206,N_11381,N_11433);
nor U12207 (N_12207,N_11036,N_11207);
nor U12208 (N_12208,N_11684,N_11875);
nor U12209 (N_12209,N_11907,N_11038);
and U12210 (N_12210,N_11080,N_11582);
xnor U12211 (N_12211,N_11305,N_11825);
or U12212 (N_12212,N_11211,N_11782);
nand U12213 (N_12213,N_11323,N_11882);
nor U12214 (N_12214,N_11217,N_11903);
nor U12215 (N_12215,N_11595,N_11188);
xor U12216 (N_12216,N_11853,N_11366);
nor U12217 (N_12217,N_11872,N_11251);
nand U12218 (N_12218,N_11292,N_11465);
nor U12219 (N_12219,N_11175,N_11371);
nand U12220 (N_12220,N_11629,N_11776);
nor U12221 (N_12221,N_11878,N_11623);
or U12222 (N_12222,N_11937,N_11820);
nand U12223 (N_12223,N_11821,N_11103);
xor U12224 (N_12224,N_11197,N_11426);
xor U12225 (N_12225,N_11420,N_11592);
or U12226 (N_12226,N_11416,N_11952);
xor U12227 (N_12227,N_11866,N_11904);
nand U12228 (N_12228,N_11015,N_11126);
or U12229 (N_12229,N_11468,N_11916);
or U12230 (N_12230,N_11387,N_11568);
and U12231 (N_12231,N_11523,N_11541);
nor U12232 (N_12232,N_11017,N_11814);
or U12233 (N_12233,N_11633,N_11124);
nor U12234 (N_12234,N_11099,N_11172);
xor U12235 (N_12235,N_11155,N_11260);
nor U12236 (N_12236,N_11456,N_11287);
and U12237 (N_12237,N_11564,N_11661);
or U12238 (N_12238,N_11176,N_11369);
nor U12239 (N_12239,N_11304,N_11222);
nand U12240 (N_12240,N_11382,N_11101);
and U12241 (N_12241,N_11183,N_11605);
and U12242 (N_12242,N_11532,N_11963);
xor U12243 (N_12243,N_11890,N_11761);
nand U12244 (N_12244,N_11847,N_11506);
nor U12245 (N_12245,N_11242,N_11786);
and U12246 (N_12246,N_11589,N_11311);
or U12247 (N_12247,N_11889,N_11266);
xnor U12248 (N_12248,N_11824,N_11616);
and U12249 (N_12249,N_11809,N_11689);
xor U12250 (N_12250,N_11432,N_11440);
and U12251 (N_12251,N_11258,N_11335);
or U12252 (N_12252,N_11944,N_11946);
nand U12253 (N_12253,N_11484,N_11504);
and U12254 (N_12254,N_11795,N_11508);
and U12255 (N_12255,N_11976,N_11941);
nor U12256 (N_12256,N_11567,N_11970);
or U12257 (N_12257,N_11673,N_11721);
or U12258 (N_12258,N_11427,N_11681);
or U12259 (N_12259,N_11837,N_11865);
nand U12260 (N_12260,N_11874,N_11977);
xnor U12261 (N_12261,N_11695,N_11517);
or U12262 (N_12262,N_11013,N_11193);
nand U12263 (N_12263,N_11054,N_11823);
or U12264 (N_12264,N_11252,N_11973);
or U12265 (N_12265,N_11832,N_11041);
and U12266 (N_12266,N_11478,N_11948);
or U12267 (N_12267,N_11634,N_11483);
and U12268 (N_12268,N_11703,N_11884);
or U12269 (N_12269,N_11096,N_11108);
and U12270 (N_12270,N_11200,N_11112);
or U12271 (N_12271,N_11236,N_11910);
xnor U12272 (N_12272,N_11284,N_11090);
nand U12273 (N_12273,N_11958,N_11331);
xor U12274 (N_12274,N_11636,N_11999);
and U12275 (N_12275,N_11348,N_11719);
nor U12276 (N_12276,N_11932,N_11893);
nand U12277 (N_12277,N_11014,N_11862);
or U12278 (N_12278,N_11012,N_11997);
nor U12279 (N_12279,N_11321,N_11424);
nor U12280 (N_12280,N_11374,N_11632);
or U12281 (N_12281,N_11152,N_11164);
or U12282 (N_12282,N_11024,N_11637);
nand U12283 (N_12283,N_11723,N_11867);
nand U12284 (N_12284,N_11615,N_11528);
and U12285 (N_12285,N_11074,N_11105);
nand U12286 (N_12286,N_11349,N_11960);
nor U12287 (N_12287,N_11908,N_11860);
nand U12288 (N_12288,N_11100,N_11545);
xnor U12289 (N_12289,N_11068,N_11685);
nor U12290 (N_12290,N_11230,N_11586);
nand U12291 (N_12291,N_11144,N_11924);
or U12292 (N_12292,N_11536,N_11058);
xor U12293 (N_12293,N_11006,N_11294);
nor U12294 (N_12294,N_11351,N_11281);
nor U12295 (N_12295,N_11255,N_11900);
xnor U12296 (N_12296,N_11045,N_11185);
or U12297 (N_12297,N_11334,N_11898);
and U12298 (N_12298,N_11846,N_11173);
xor U12299 (N_12299,N_11906,N_11515);
nand U12300 (N_12300,N_11115,N_11610);
nor U12301 (N_12301,N_11435,N_11931);
nor U12302 (N_12302,N_11008,N_11047);
and U12303 (N_12303,N_11964,N_11982);
and U12304 (N_12304,N_11669,N_11347);
or U12305 (N_12305,N_11822,N_11249);
and U12306 (N_12306,N_11939,N_11611);
xor U12307 (N_12307,N_11079,N_11094);
and U12308 (N_12308,N_11728,N_11451);
or U12309 (N_12309,N_11110,N_11726);
nor U12310 (N_12310,N_11359,N_11390);
nor U12311 (N_12311,N_11250,N_11579);
nor U12312 (N_12312,N_11231,N_11338);
nor U12313 (N_12313,N_11565,N_11033);
and U12314 (N_12314,N_11346,N_11326);
nand U12315 (N_12315,N_11438,N_11365);
or U12316 (N_12316,N_11171,N_11542);
xor U12317 (N_12317,N_11324,N_11482);
and U12318 (N_12318,N_11062,N_11098);
nand U12319 (N_12319,N_11690,N_11602);
nand U12320 (N_12320,N_11018,N_11053);
or U12321 (N_12321,N_11227,N_11777);
and U12322 (N_12322,N_11779,N_11674);
and U12323 (N_12323,N_11267,N_11668);
or U12324 (N_12324,N_11060,N_11187);
nand U12325 (N_12325,N_11265,N_11448);
nor U12326 (N_12326,N_11718,N_11254);
nor U12327 (N_12327,N_11841,N_11167);
xor U12328 (N_12328,N_11544,N_11731);
nor U12329 (N_12329,N_11496,N_11974);
and U12330 (N_12330,N_11771,N_11158);
xor U12331 (N_12331,N_11953,N_11128);
nand U12332 (N_12332,N_11672,N_11784);
xnor U12333 (N_12333,N_11142,N_11191);
or U12334 (N_12334,N_11838,N_11763);
or U12335 (N_12335,N_11886,N_11883);
nand U12336 (N_12336,N_11149,N_11470);
or U12337 (N_12337,N_11923,N_11499);
or U12338 (N_12338,N_11315,N_11020);
nor U12339 (N_12339,N_11670,N_11443);
xor U12340 (N_12340,N_11758,N_11905);
nand U12341 (N_12341,N_11936,N_11409);
or U12342 (N_12342,N_11216,N_11751);
nand U12343 (N_12343,N_11421,N_11730);
and U12344 (N_12344,N_11362,N_11739);
or U12345 (N_12345,N_11244,N_11901);
nand U12346 (N_12346,N_11954,N_11996);
or U12347 (N_12347,N_11859,N_11279);
xor U12348 (N_12348,N_11474,N_11654);
xnor U12349 (N_12349,N_11855,N_11696);
or U12350 (N_12350,N_11322,N_11796);
or U12351 (N_12351,N_11756,N_11863);
nor U12352 (N_12352,N_11570,N_11261);
and U12353 (N_12353,N_11601,N_11555);
nor U12354 (N_12354,N_11356,N_11190);
xnor U12355 (N_12355,N_11289,N_11733);
xor U12356 (N_12356,N_11117,N_11301);
nand U12357 (N_12357,N_11686,N_11563);
or U12358 (N_12358,N_11804,N_11011);
or U12359 (N_12359,N_11093,N_11269);
xnor U12360 (N_12360,N_11835,N_11378);
nand U12361 (N_12361,N_11034,N_11461);
xor U12362 (N_12362,N_11135,N_11643);
and U12363 (N_12363,N_11705,N_11671);
and U12364 (N_12364,N_11622,N_11021);
xor U12365 (N_12365,N_11042,N_11275);
and U12366 (N_12366,N_11688,N_11113);
xnor U12367 (N_12367,N_11538,N_11609);
and U12368 (N_12368,N_11577,N_11587);
nand U12369 (N_12369,N_11379,N_11558);
nand U12370 (N_12370,N_11966,N_11262);
nand U12371 (N_12371,N_11447,N_11136);
nor U12372 (N_12372,N_11930,N_11746);
or U12373 (N_12373,N_11707,N_11228);
or U12374 (N_12374,N_11239,N_11223);
or U12375 (N_12375,N_11143,N_11599);
nor U12376 (N_12376,N_11938,N_11460);
or U12377 (N_12377,N_11150,N_11243);
nand U12378 (N_12378,N_11624,N_11114);
xor U12379 (N_12379,N_11411,N_11552);
and U12380 (N_12380,N_11133,N_11488);
nand U12381 (N_12381,N_11129,N_11762);
and U12382 (N_12382,N_11598,N_11077);
and U12383 (N_12383,N_11706,N_11522);
and U12384 (N_12384,N_11071,N_11333);
xnor U12385 (N_12385,N_11240,N_11154);
xor U12386 (N_12386,N_11708,N_11088);
nand U12387 (N_12387,N_11486,N_11296);
and U12388 (N_12388,N_11475,N_11049);
and U12389 (N_12389,N_11682,N_11947);
or U12390 (N_12390,N_11355,N_11477);
nand U12391 (N_12391,N_11219,N_11547);
or U12392 (N_12392,N_11202,N_11339);
or U12393 (N_12393,N_11082,N_11199);
and U12394 (N_12394,N_11122,N_11109);
or U12395 (N_12395,N_11454,N_11557);
xnor U12396 (N_12396,N_11026,N_11076);
or U12397 (N_12397,N_11064,N_11316);
nor U12398 (N_12398,N_11791,N_11367);
nor U12399 (N_12399,N_11612,N_11213);
nor U12400 (N_12400,N_11272,N_11291);
nor U12401 (N_12401,N_11829,N_11657);
nand U12402 (N_12402,N_11330,N_11663);
nand U12403 (N_12403,N_11896,N_11513);
xnor U12404 (N_12404,N_11329,N_11417);
xor U12405 (N_12405,N_11480,N_11743);
nor U12406 (N_12406,N_11271,N_11141);
nand U12407 (N_12407,N_11734,N_11914);
nor U12408 (N_12408,N_11581,N_11922);
or U12409 (N_12409,N_11554,N_11116);
xor U12410 (N_12410,N_11234,N_11037);
nor U12411 (N_12411,N_11418,N_11205);
xor U12412 (N_12412,N_11701,N_11801);
xor U12413 (N_12413,N_11881,N_11702);
xnor U12414 (N_12414,N_11336,N_11463);
nand U12415 (N_12415,N_11876,N_11775);
xor U12416 (N_12416,N_11868,N_11481);
xnor U12417 (N_12417,N_11529,N_11850);
nand U12418 (N_12418,N_11497,N_11446);
nand U12419 (N_12419,N_11429,N_11314);
nand U12420 (N_12420,N_11273,N_11992);
nor U12421 (N_12421,N_11590,N_11993);
and U12422 (N_12422,N_11309,N_11278);
xor U12423 (N_12423,N_11489,N_11642);
xor U12424 (N_12424,N_11892,N_11614);
and U12425 (N_12425,N_11139,N_11479);
and U12426 (N_12426,N_11956,N_11422);
or U12427 (N_12427,N_11754,N_11729);
nor U12428 (N_12428,N_11044,N_11516);
xnor U12429 (N_12429,N_11833,N_11001);
xnor U12430 (N_12430,N_11132,N_11151);
or U12431 (N_12431,N_11186,N_11078);
nor U12432 (N_12432,N_11638,N_11452);
xnor U12433 (N_12433,N_11998,N_11765);
xor U12434 (N_12434,N_11562,N_11241);
and U12435 (N_12435,N_11005,N_11072);
xnor U12436 (N_12436,N_11007,N_11206);
nand U12437 (N_12437,N_11798,N_11372);
and U12438 (N_12438,N_11120,N_11300);
or U12439 (N_12439,N_11307,N_11894);
or U12440 (N_12440,N_11514,N_11238);
and U12441 (N_12441,N_11665,N_11157);
nand U12442 (N_12442,N_11649,N_11724);
nand U12443 (N_12443,N_11063,N_11606);
nor U12444 (N_12444,N_11716,N_11646);
nand U12445 (N_12445,N_11680,N_11318);
nand U12446 (N_12446,N_11957,N_11888);
nand U12447 (N_12447,N_11394,N_11902);
and U12448 (N_12448,N_11539,N_11772);
and U12449 (N_12449,N_11419,N_11345);
and U12450 (N_12450,N_11747,N_11667);
nand U12451 (N_12451,N_11343,N_11437);
nor U12452 (N_12452,N_11655,N_11327);
or U12453 (N_12453,N_11067,N_11370);
xnor U12454 (N_12454,N_11357,N_11576);
nor U12455 (N_12455,N_11917,N_11065);
nor U12456 (N_12456,N_11487,N_11248);
nor U12457 (N_12457,N_11061,N_11918);
and U12458 (N_12458,N_11030,N_11711);
or U12459 (N_12459,N_11573,N_11600);
xor U12460 (N_12460,N_11895,N_11556);
nor U12461 (N_12461,N_11189,N_11583);
nor U12462 (N_12462,N_11224,N_11161);
and U12463 (N_12463,N_11864,N_11738);
nor U12464 (N_12464,N_11147,N_11466);
nor U12465 (N_12465,N_11313,N_11645);
xor U12466 (N_12466,N_11140,N_11412);
nand U12467 (N_12467,N_11603,N_11769);
or U12468 (N_12468,N_11534,N_11620);
xor U12469 (N_12469,N_11257,N_11766);
nor U12470 (N_12470,N_11879,N_11521);
nand U12471 (N_12471,N_11312,N_11059);
nor U12472 (N_12472,N_11457,N_11286);
or U12473 (N_12473,N_11328,N_11032);
and U12474 (N_12474,N_11118,N_11441);
and U12475 (N_12475,N_11537,N_11130);
nand U12476 (N_12476,N_11235,N_11978);
and U12477 (N_12477,N_11293,N_11302);
and U12478 (N_12478,N_11621,N_11793);
or U12479 (N_12479,N_11691,N_11220);
and U12480 (N_12480,N_11081,N_11951);
or U12481 (N_12481,N_11617,N_11755);
or U12482 (N_12482,N_11714,N_11493);
and U12483 (N_12483,N_11263,N_11921);
xor U12484 (N_12484,N_11713,N_11121);
xnor U12485 (N_12485,N_11350,N_11736);
nor U12486 (N_12486,N_11306,N_11455);
or U12487 (N_12487,N_11462,N_11398);
nand U12488 (N_12488,N_11512,N_11025);
or U12489 (N_12489,N_11588,N_11710);
or U12490 (N_12490,N_11675,N_11403);
nand U12491 (N_12491,N_11247,N_11400);
xnor U12492 (N_12492,N_11246,N_11169);
or U12493 (N_12493,N_11004,N_11342);
and U12494 (N_12494,N_11039,N_11270);
nand U12495 (N_12495,N_11807,N_11010);
and U12496 (N_12496,N_11540,N_11332);
xnor U12497 (N_12497,N_11277,N_11836);
xor U12498 (N_12498,N_11156,N_11849);
and U12499 (N_12499,N_11933,N_11397);
or U12500 (N_12500,N_11247,N_11956);
nor U12501 (N_12501,N_11928,N_11500);
xnor U12502 (N_12502,N_11845,N_11787);
and U12503 (N_12503,N_11835,N_11133);
and U12504 (N_12504,N_11577,N_11664);
or U12505 (N_12505,N_11982,N_11381);
or U12506 (N_12506,N_11473,N_11270);
nor U12507 (N_12507,N_11192,N_11594);
and U12508 (N_12508,N_11041,N_11748);
nor U12509 (N_12509,N_11301,N_11130);
and U12510 (N_12510,N_11956,N_11065);
or U12511 (N_12511,N_11190,N_11019);
nand U12512 (N_12512,N_11025,N_11285);
or U12513 (N_12513,N_11792,N_11160);
or U12514 (N_12514,N_11672,N_11162);
xnor U12515 (N_12515,N_11884,N_11607);
or U12516 (N_12516,N_11224,N_11615);
nand U12517 (N_12517,N_11309,N_11368);
nor U12518 (N_12518,N_11473,N_11551);
xnor U12519 (N_12519,N_11420,N_11192);
nand U12520 (N_12520,N_11114,N_11997);
nor U12521 (N_12521,N_11855,N_11595);
or U12522 (N_12522,N_11650,N_11766);
nand U12523 (N_12523,N_11013,N_11797);
and U12524 (N_12524,N_11974,N_11649);
nor U12525 (N_12525,N_11263,N_11282);
nor U12526 (N_12526,N_11415,N_11440);
or U12527 (N_12527,N_11708,N_11120);
and U12528 (N_12528,N_11415,N_11739);
nor U12529 (N_12529,N_11326,N_11151);
xnor U12530 (N_12530,N_11556,N_11864);
nand U12531 (N_12531,N_11848,N_11184);
nor U12532 (N_12532,N_11893,N_11377);
nand U12533 (N_12533,N_11781,N_11867);
nand U12534 (N_12534,N_11451,N_11742);
xnor U12535 (N_12535,N_11466,N_11067);
and U12536 (N_12536,N_11915,N_11569);
nand U12537 (N_12537,N_11757,N_11242);
nand U12538 (N_12538,N_11409,N_11004);
xor U12539 (N_12539,N_11606,N_11818);
and U12540 (N_12540,N_11405,N_11271);
nand U12541 (N_12541,N_11653,N_11137);
and U12542 (N_12542,N_11125,N_11757);
nand U12543 (N_12543,N_11538,N_11976);
and U12544 (N_12544,N_11028,N_11751);
xnor U12545 (N_12545,N_11215,N_11167);
nor U12546 (N_12546,N_11611,N_11871);
or U12547 (N_12547,N_11910,N_11802);
nor U12548 (N_12548,N_11622,N_11443);
nand U12549 (N_12549,N_11216,N_11588);
and U12550 (N_12550,N_11390,N_11069);
xnor U12551 (N_12551,N_11173,N_11308);
nand U12552 (N_12552,N_11119,N_11478);
xor U12553 (N_12553,N_11490,N_11933);
or U12554 (N_12554,N_11300,N_11940);
nand U12555 (N_12555,N_11570,N_11785);
nor U12556 (N_12556,N_11693,N_11606);
nor U12557 (N_12557,N_11741,N_11640);
or U12558 (N_12558,N_11512,N_11343);
nand U12559 (N_12559,N_11684,N_11478);
nand U12560 (N_12560,N_11975,N_11061);
xor U12561 (N_12561,N_11450,N_11908);
and U12562 (N_12562,N_11801,N_11360);
nor U12563 (N_12563,N_11972,N_11379);
nor U12564 (N_12564,N_11850,N_11894);
or U12565 (N_12565,N_11332,N_11819);
nor U12566 (N_12566,N_11168,N_11350);
nand U12567 (N_12567,N_11283,N_11876);
and U12568 (N_12568,N_11246,N_11513);
nor U12569 (N_12569,N_11328,N_11475);
and U12570 (N_12570,N_11455,N_11600);
nand U12571 (N_12571,N_11830,N_11242);
nand U12572 (N_12572,N_11563,N_11261);
or U12573 (N_12573,N_11889,N_11656);
nand U12574 (N_12574,N_11179,N_11387);
and U12575 (N_12575,N_11396,N_11823);
nor U12576 (N_12576,N_11461,N_11595);
or U12577 (N_12577,N_11010,N_11176);
nand U12578 (N_12578,N_11525,N_11756);
and U12579 (N_12579,N_11948,N_11808);
xnor U12580 (N_12580,N_11511,N_11891);
xnor U12581 (N_12581,N_11478,N_11603);
or U12582 (N_12582,N_11554,N_11603);
nor U12583 (N_12583,N_11715,N_11071);
and U12584 (N_12584,N_11653,N_11556);
nand U12585 (N_12585,N_11901,N_11548);
and U12586 (N_12586,N_11969,N_11598);
and U12587 (N_12587,N_11984,N_11501);
xor U12588 (N_12588,N_11845,N_11627);
or U12589 (N_12589,N_11811,N_11473);
and U12590 (N_12590,N_11121,N_11550);
and U12591 (N_12591,N_11387,N_11585);
xnor U12592 (N_12592,N_11603,N_11579);
nor U12593 (N_12593,N_11408,N_11268);
nor U12594 (N_12594,N_11946,N_11469);
nand U12595 (N_12595,N_11265,N_11348);
nor U12596 (N_12596,N_11074,N_11462);
nand U12597 (N_12597,N_11680,N_11207);
or U12598 (N_12598,N_11181,N_11617);
and U12599 (N_12599,N_11954,N_11592);
or U12600 (N_12600,N_11404,N_11844);
and U12601 (N_12601,N_11969,N_11305);
xnor U12602 (N_12602,N_11889,N_11967);
nor U12603 (N_12603,N_11871,N_11579);
and U12604 (N_12604,N_11101,N_11979);
xor U12605 (N_12605,N_11041,N_11579);
nand U12606 (N_12606,N_11891,N_11857);
nor U12607 (N_12607,N_11121,N_11454);
xor U12608 (N_12608,N_11121,N_11139);
nor U12609 (N_12609,N_11757,N_11470);
nor U12610 (N_12610,N_11016,N_11267);
nand U12611 (N_12611,N_11657,N_11675);
nand U12612 (N_12612,N_11663,N_11481);
nor U12613 (N_12613,N_11161,N_11381);
or U12614 (N_12614,N_11949,N_11936);
nand U12615 (N_12615,N_11936,N_11707);
or U12616 (N_12616,N_11459,N_11956);
nor U12617 (N_12617,N_11895,N_11231);
nor U12618 (N_12618,N_11081,N_11436);
nor U12619 (N_12619,N_11605,N_11768);
and U12620 (N_12620,N_11639,N_11081);
nor U12621 (N_12621,N_11828,N_11384);
nand U12622 (N_12622,N_11735,N_11773);
nor U12623 (N_12623,N_11426,N_11725);
nor U12624 (N_12624,N_11939,N_11882);
nor U12625 (N_12625,N_11154,N_11443);
or U12626 (N_12626,N_11182,N_11605);
or U12627 (N_12627,N_11972,N_11429);
xor U12628 (N_12628,N_11236,N_11013);
nor U12629 (N_12629,N_11392,N_11939);
and U12630 (N_12630,N_11909,N_11666);
xor U12631 (N_12631,N_11916,N_11708);
nor U12632 (N_12632,N_11954,N_11934);
and U12633 (N_12633,N_11482,N_11789);
xnor U12634 (N_12634,N_11103,N_11461);
or U12635 (N_12635,N_11990,N_11221);
xor U12636 (N_12636,N_11884,N_11311);
xnor U12637 (N_12637,N_11095,N_11789);
or U12638 (N_12638,N_11692,N_11763);
xor U12639 (N_12639,N_11341,N_11867);
nand U12640 (N_12640,N_11822,N_11768);
nand U12641 (N_12641,N_11025,N_11536);
nand U12642 (N_12642,N_11287,N_11682);
and U12643 (N_12643,N_11355,N_11156);
or U12644 (N_12644,N_11155,N_11306);
nor U12645 (N_12645,N_11031,N_11187);
xnor U12646 (N_12646,N_11199,N_11405);
nand U12647 (N_12647,N_11241,N_11131);
or U12648 (N_12648,N_11385,N_11348);
xor U12649 (N_12649,N_11928,N_11611);
nand U12650 (N_12650,N_11789,N_11609);
nand U12651 (N_12651,N_11953,N_11227);
and U12652 (N_12652,N_11422,N_11094);
or U12653 (N_12653,N_11536,N_11155);
nand U12654 (N_12654,N_11185,N_11150);
or U12655 (N_12655,N_11443,N_11755);
nand U12656 (N_12656,N_11988,N_11275);
nor U12657 (N_12657,N_11906,N_11031);
nand U12658 (N_12658,N_11891,N_11884);
nor U12659 (N_12659,N_11102,N_11392);
nand U12660 (N_12660,N_11146,N_11489);
nor U12661 (N_12661,N_11388,N_11433);
nand U12662 (N_12662,N_11066,N_11237);
nand U12663 (N_12663,N_11138,N_11373);
or U12664 (N_12664,N_11273,N_11577);
xor U12665 (N_12665,N_11940,N_11641);
or U12666 (N_12666,N_11470,N_11628);
or U12667 (N_12667,N_11960,N_11655);
nor U12668 (N_12668,N_11151,N_11529);
nor U12669 (N_12669,N_11933,N_11489);
or U12670 (N_12670,N_11971,N_11548);
and U12671 (N_12671,N_11257,N_11516);
xor U12672 (N_12672,N_11853,N_11264);
or U12673 (N_12673,N_11462,N_11513);
or U12674 (N_12674,N_11623,N_11593);
and U12675 (N_12675,N_11219,N_11104);
or U12676 (N_12676,N_11019,N_11245);
nand U12677 (N_12677,N_11297,N_11380);
xor U12678 (N_12678,N_11837,N_11244);
xnor U12679 (N_12679,N_11748,N_11393);
or U12680 (N_12680,N_11818,N_11754);
and U12681 (N_12681,N_11672,N_11028);
and U12682 (N_12682,N_11417,N_11184);
nor U12683 (N_12683,N_11322,N_11348);
or U12684 (N_12684,N_11434,N_11939);
and U12685 (N_12685,N_11255,N_11540);
or U12686 (N_12686,N_11863,N_11741);
or U12687 (N_12687,N_11889,N_11649);
nor U12688 (N_12688,N_11570,N_11043);
and U12689 (N_12689,N_11613,N_11897);
nand U12690 (N_12690,N_11790,N_11248);
nor U12691 (N_12691,N_11890,N_11453);
nor U12692 (N_12692,N_11912,N_11861);
nor U12693 (N_12693,N_11392,N_11142);
nand U12694 (N_12694,N_11546,N_11837);
xor U12695 (N_12695,N_11942,N_11507);
nand U12696 (N_12696,N_11601,N_11533);
nand U12697 (N_12697,N_11383,N_11907);
nor U12698 (N_12698,N_11941,N_11743);
or U12699 (N_12699,N_11522,N_11193);
nor U12700 (N_12700,N_11397,N_11730);
nor U12701 (N_12701,N_11788,N_11582);
or U12702 (N_12702,N_11545,N_11302);
and U12703 (N_12703,N_11597,N_11705);
and U12704 (N_12704,N_11495,N_11199);
xnor U12705 (N_12705,N_11774,N_11482);
nand U12706 (N_12706,N_11053,N_11292);
nand U12707 (N_12707,N_11354,N_11125);
nand U12708 (N_12708,N_11065,N_11868);
and U12709 (N_12709,N_11258,N_11508);
and U12710 (N_12710,N_11797,N_11752);
nor U12711 (N_12711,N_11030,N_11049);
nand U12712 (N_12712,N_11378,N_11381);
and U12713 (N_12713,N_11343,N_11476);
nor U12714 (N_12714,N_11353,N_11328);
xor U12715 (N_12715,N_11508,N_11593);
nand U12716 (N_12716,N_11487,N_11604);
or U12717 (N_12717,N_11707,N_11677);
nor U12718 (N_12718,N_11424,N_11536);
or U12719 (N_12719,N_11056,N_11533);
nand U12720 (N_12720,N_11376,N_11151);
xnor U12721 (N_12721,N_11051,N_11547);
xnor U12722 (N_12722,N_11729,N_11709);
or U12723 (N_12723,N_11621,N_11664);
xnor U12724 (N_12724,N_11702,N_11315);
and U12725 (N_12725,N_11785,N_11091);
and U12726 (N_12726,N_11933,N_11213);
or U12727 (N_12727,N_11046,N_11182);
nor U12728 (N_12728,N_11365,N_11329);
or U12729 (N_12729,N_11349,N_11228);
nand U12730 (N_12730,N_11387,N_11468);
and U12731 (N_12731,N_11428,N_11404);
and U12732 (N_12732,N_11869,N_11507);
xor U12733 (N_12733,N_11904,N_11447);
and U12734 (N_12734,N_11543,N_11904);
nor U12735 (N_12735,N_11764,N_11024);
xnor U12736 (N_12736,N_11051,N_11898);
or U12737 (N_12737,N_11931,N_11296);
or U12738 (N_12738,N_11352,N_11928);
or U12739 (N_12739,N_11842,N_11642);
nand U12740 (N_12740,N_11428,N_11497);
and U12741 (N_12741,N_11188,N_11123);
xor U12742 (N_12742,N_11364,N_11176);
nor U12743 (N_12743,N_11581,N_11212);
and U12744 (N_12744,N_11171,N_11624);
nor U12745 (N_12745,N_11108,N_11774);
nor U12746 (N_12746,N_11378,N_11087);
nand U12747 (N_12747,N_11113,N_11085);
xnor U12748 (N_12748,N_11653,N_11654);
and U12749 (N_12749,N_11979,N_11966);
and U12750 (N_12750,N_11079,N_11219);
and U12751 (N_12751,N_11403,N_11912);
or U12752 (N_12752,N_11187,N_11433);
nand U12753 (N_12753,N_11839,N_11311);
xor U12754 (N_12754,N_11948,N_11093);
or U12755 (N_12755,N_11308,N_11114);
or U12756 (N_12756,N_11489,N_11483);
and U12757 (N_12757,N_11265,N_11687);
nor U12758 (N_12758,N_11378,N_11108);
nor U12759 (N_12759,N_11235,N_11390);
nand U12760 (N_12760,N_11807,N_11716);
nand U12761 (N_12761,N_11527,N_11484);
nand U12762 (N_12762,N_11188,N_11748);
and U12763 (N_12763,N_11992,N_11536);
nand U12764 (N_12764,N_11776,N_11386);
nand U12765 (N_12765,N_11988,N_11173);
and U12766 (N_12766,N_11124,N_11693);
xnor U12767 (N_12767,N_11393,N_11657);
xnor U12768 (N_12768,N_11569,N_11294);
or U12769 (N_12769,N_11158,N_11166);
nand U12770 (N_12770,N_11436,N_11874);
nand U12771 (N_12771,N_11127,N_11606);
nor U12772 (N_12772,N_11548,N_11607);
xor U12773 (N_12773,N_11897,N_11620);
nor U12774 (N_12774,N_11450,N_11640);
nand U12775 (N_12775,N_11133,N_11550);
nor U12776 (N_12776,N_11295,N_11241);
nand U12777 (N_12777,N_11544,N_11814);
xnor U12778 (N_12778,N_11831,N_11378);
xor U12779 (N_12779,N_11854,N_11087);
nand U12780 (N_12780,N_11335,N_11729);
nand U12781 (N_12781,N_11355,N_11944);
nor U12782 (N_12782,N_11073,N_11233);
nand U12783 (N_12783,N_11028,N_11928);
and U12784 (N_12784,N_11053,N_11534);
or U12785 (N_12785,N_11258,N_11102);
xor U12786 (N_12786,N_11828,N_11621);
and U12787 (N_12787,N_11919,N_11712);
and U12788 (N_12788,N_11298,N_11471);
xor U12789 (N_12789,N_11780,N_11540);
xnor U12790 (N_12790,N_11201,N_11106);
nand U12791 (N_12791,N_11259,N_11312);
and U12792 (N_12792,N_11015,N_11680);
and U12793 (N_12793,N_11015,N_11429);
and U12794 (N_12794,N_11271,N_11726);
and U12795 (N_12795,N_11596,N_11067);
xnor U12796 (N_12796,N_11210,N_11122);
nor U12797 (N_12797,N_11400,N_11629);
xnor U12798 (N_12798,N_11362,N_11864);
or U12799 (N_12799,N_11604,N_11701);
and U12800 (N_12800,N_11674,N_11819);
or U12801 (N_12801,N_11880,N_11400);
xnor U12802 (N_12802,N_11683,N_11132);
or U12803 (N_12803,N_11981,N_11896);
nand U12804 (N_12804,N_11588,N_11574);
xnor U12805 (N_12805,N_11307,N_11473);
xnor U12806 (N_12806,N_11980,N_11845);
nand U12807 (N_12807,N_11342,N_11753);
nor U12808 (N_12808,N_11955,N_11658);
nand U12809 (N_12809,N_11847,N_11038);
or U12810 (N_12810,N_11183,N_11464);
xnor U12811 (N_12811,N_11763,N_11452);
or U12812 (N_12812,N_11218,N_11096);
nand U12813 (N_12813,N_11078,N_11667);
nor U12814 (N_12814,N_11724,N_11080);
or U12815 (N_12815,N_11130,N_11004);
nor U12816 (N_12816,N_11751,N_11001);
xor U12817 (N_12817,N_11059,N_11384);
and U12818 (N_12818,N_11374,N_11171);
nor U12819 (N_12819,N_11203,N_11317);
xnor U12820 (N_12820,N_11872,N_11965);
nor U12821 (N_12821,N_11674,N_11821);
nand U12822 (N_12822,N_11793,N_11895);
and U12823 (N_12823,N_11618,N_11239);
nor U12824 (N_12824,N_11965,N_11159);
nor U12825 (N_12825,N_11503,N_11245);
xnor U12826 (N_12826,N_11291,N_11128);
or U12827 (N_12827,N_11758,N_11122);
and U12828 (N_12828,N_11159,N_11500);
and U12829 (N_12829,N_11574,N_11120);
nor U12830 (N_12830,N_11934,N_11689);
xnor U12831 (N_12831,N_11712,N_11470);
nor U12832 (N_12832,N_11376,N_11456);
or U12833 (N_12833,N_11118,N_11502);
or U12834 (N_12834,N_11468,N_11274);
xor U12835 (N_12835,N_11075,N_11091);
or U12836 (N_12836,N_11634,N_11969);
xor U12837 (N_12837,N_11243,N_11453);
nand U12838 (N_12838,N_11559,N_11392);
or U12839 (N_12839,N_11899,N_11060);
nand U12840 (N_12840,N_11838,N_11871);
or U12841 (N_12841,N_11175,N_11321);
xnor U12842 (N_12842,N_11887,N_11199);
xor U12843 (N_12843,N_11215,N_11287);
nand U12844 (N_12844,N_11533,N_11313);
and U12845 (N_12845,N_11639,N_11990);
or U12846 (N_12846,N_11745,N_11328);
xnor U12847 (N_12847,N_11813,N_11465);
and U12848 (N_12848,N_11606,N_11504);
and U12849 (N_12849,N_11145,N_11113);
xor U12850 (N_12850,N_11498,N_11686);
and U12851 (N_12851,N_11678,N_11454);
or U12852 (N_12852,N_11384,N_11707);
nand U12853 (N_12853,N_11780,N_11322);
or U12854 (N_12854,N_11660,N_11415);
nor U12855 (N_12855,N_11040,N_11999);
nor U12856 (N_12856,N_11057,N_11784);
xor U12857 (N_12857,N_11038,N_11087);
xor U12858 (N_12858,N_11789,N_11235);
or U12859 (N_12859,N_11506,N_11009);
and U12860 (N_12860,N_11947,N_11684);
nor U12861 (N_12861,N_11601,N_11559);
or U12862 (N_12862,N_11617,N_11679);
or U12863 (N_12863,N_11170,N_11586);
xor U12864 (N_12864,N_11989,N_11702);
nor U12865 (N_12865,N_11133,N_11066);
and U12866 (N_12866,N_11953,N_11465);
or U12867 (N_12867,N_11053,N_11453);
nor U12868 (N_12868,N_11652,N_11003);
and U12869 (N_12869,N_11943,N_11343);
nor U12870 (N_12870,N_11305,N_11739);
or U12871 (N_12871,N_11355,N_11613);
and U12872 (N_12872,N_11570,N_11054);
and U12873 (N_12873,N_11669,N_11796);
or U12874 (N_12874,N_11471,N_11627);
or U12875 (N_12875,N_11451,N_11767);
xnor U12876 (N_12876,N_11913,N_11164);
and U12877 (N_12877,N_11712,N_11748);
nand U12878 (N_12878,N_11536,N_11371);
xnor U12879 (N_12879,N_11488,N_11639);
or U12880 (N_12880,N_11620,N_11323);
and U12881 (N_12881,N_11219,N_11179);
nor U12882 (N_12882,N_11578,N_11340);
and U12883 (N_12883,N_11517,N_11255);
or U12884 (N_12884,N_11309,N_11634);
xor U12885 (N_12885,N_11787,N_11508);
nand U12886 (N_12886,N_11030,N_11408);
nand U12887 (N_12887,N_11773,N_11090);
xnor U12888 (N_12888,N_11466,N_11691);
nor U12889 (N_12889,N_11140,N_11556);
nand U12890 (N_12890,N_11637,N_11030);
nor U12891 (N_12891,N_11783,N_11419);
nand U12892 (N_12892,N_11568,N_11556);
nand U12893 (N_12893,N_11780,N_11304);
nor U12894 (N_12894,N_11263,N_11812);
xnor U12895 (N_12895,N_11321,N_11488);
xnor U12896 (N_12896,N_11148,N_11768);
xnor U12897 (N_12897,N_11308,N_11435);
and U12898 (N_12898,N_11564,N_11144);
nor U12899 (N_12899,N_11231,N_11273);
nand U12900 (N_12900,N_11028,N_11342);
nand U12901 (N_12901,N_11279,N_11758);
xor U12902 (N_12902,N_11443,N_11913);
xor U12903 (N_12903,N_11715,N_11827);
or U12904 (N_12904,N_11266,N_11144);
nand U12905 (N_12905,N_11978,N_11156);
xor U12906 (N_12906,N_11896,N_11342);
nand U12907 (N_12907,N_11527,N_11258);
and U12908 (N_12908,N_11353,N_11443);
nand U12909 (N_12909,N_11726,N_11060);
xor U12910 (N_12910,N_11535,N_11623);
and U12911 (N_12911,N_11004,N_11792);
or U12912 (N_12912,N_11413,N_11170);
and U12913 (N_12913,N_11397,N_11472);
or U12914 (N_12914,N_11659,N_11163);
or U12915 (N_12915,N_11705,N_11383);
and U12916 (N_12916,N_11482,N_11277);
nand U12917 (N_12917,N_11029,N_11015);
nand U12918 (N_12918,N_11047,N_11114);
nand U12919 (N_12919,N_11433,N_11710);
or U12920 (N_12920,N_11236,N_11540);
or U12921 (N_12921,N_11225,N_11477);
nor U12922 (N_12922,N_11773,N_11602);
xnor U12923 (N_12923,N_11571,N_11196);
xor U12924 (N_12924,N_11265,N_11452);
nand U12925 (N_12925,N_11919,N_11799);
xor U12926 (N_12926,N_11650,N_11172);
or U12927 (N_12927,N_11610,N_11948);
and U12928 (N_12928,N_11084,N_11060);
or U12929 (N_12929,N_11107,N_11989);
xnor U12930 (N_12930,N_11758,N_11248);
nor U12931 (N_12931,N_11575,N_11508);
or U12932 (N_12932,N_11569,N_11058);
nor U12933 (N_12933,N_11387,N_11293);
and U12934 (N_12934,N_11576,N_11684);
nor U12935 (N_12935,N_11210,N_11852);
or U12936 (N_12936,N_11732,N_11440);
or U12937 (N_12937,N_11832,N_11049);
nand U12938 (N_12938,N_11758,N_11995);
nand U12939 (N_12939,N_11942,N_11856);
nand U12940 (N_12940,N_11298,N_11053);
and U12941 (N_12941,N_11052,N_11879);
and U12942 (N_12942,N_11620,N_11597);
xnor U12943 (N_12943,N_11633,N_11959);
nand U12944 (N_12944,N_11539,N_11752);
or U12945 (N_12945,N_11424,N_11002);
nand U12946 (N_12946,N_11214,N_11774);
or U12947 (N_12947,N_11203,N_11584);
or U12948 (N_12948,N_11591,N_11254);
nand U12949 (N_12949,N_11390,N_11024);
nand U12950 (N_12950,N_11529,N_11437);
nor U12951 (N_12951,N_11904,N_11991);
nand U12952 (N_12952,N_11818,N_11147);
xor U12953 (N_12953,N_11004,N_11659);
nor U12954 (N_12954,N_11187,N_11936);
nand U12955 (N_12955,N_11101,N_11466);
or U12956 (N_12956,N_11877,N_11550);
or U12957 (N_12957,N_11586,N_11250);
or U12958 (N_12958,N_11838,N_11418);
xnor U12959 (N_12959,N_11711,N_11258);
xnor U12960 (N_12960,N_11850,N_11405);
xnor U12961 (N_12961,N_11077,N_11421);
or U12962 (N_12962,N_11477,N_11714);
nor U12963 (N_12963,N_11734,N_11957);
or U12964 (N_12964,N_11715,N_11160);
and U12965 (N_12965,N_11840,N_11264);
nand U12966 (N_12966,N_11160,N_11556);
and U12967 (N_12967,N_11057,N_11564);
nor U12968 (N_12968,N_11502,N_11945);
nand U12969 (N_12969,N_11156,N_11250);
or U12970 (N_12970,N_11538,N_11088);
nor U12971 (N_12971,N_11164,N_11419);
and U12972 (N_12972,N_11371,N_11111);
or U12973 (N_12973,N_11132,N_11653);
nand U12974 (N_12974,N_11602,N_11812);
xnor U12975 (N_12975,N_11036,N_11275);
nor U12976 (N_12976,N_11363,N_11233);
and U12977 (N_12977,N_11514,N_11529);
xor U12978 (N_12978,N_11248,N_11034);
xor U12979 (N_12979,N_11469,N_11356);
or U12980 (N_12980,N_11661,N_11088);
or U12981 (N_12981,N_11469,N_11264);
xnor U12982 (N_12982,N_11381,N_11867);
nor U12983 (N_12983,N_11063,N_11289);
nor U12984 (N_12984,N_11098,N_11962);
or U12985 (N_12985,N_11215,N_11246);
or U12986 (N_12986,N_11000,N_11537);
or U12987 (N_12987,N_11469,N_11140);
nor U12988 (N_12988,N_11039,N_11392);
xor U12989 (N_12989,N_11961,N_11522);
or U12990 (N_12990,N_11046,N_11511);
xor U12991 (N_12991,N_11916,N_11027);
or U12992 (N_12992,N_11552,N_11829);
or U12993 (N_12993,N_11640,N_11797);
xnor U12994 (N_12994,N_11863,N_11020);
xnor U12995 (N_12995,N_11538,N_11185);
and U12996 (N_12996,N_11017,N_11373);
and U12997 (N_12997,N_11973,N_11032);
xor U12998 (N_12998,N_11597,N_11747);
xor U12999 (N_12999,N_11380,N_11735);
and U13000 (N_13000,N_12578,N_12449);
and U13001 (N_13001,N_12158,N_12344);
xnor U13002 (N_13002,N_12435,N_12661);
or U13003 (N_13003,N_12123,N_12525);
and U13004 (N_13004,N_12125,N_12469);
xnor U13005 (N_13005,N_12777,N_12984);
xor U13006 (N_13006,N_12851,N_12061);
or U13007 (N_13007,N_12737,N_12729);
xor U13008 (N_13008,N_12367,N_12756);
nand U13009 (N_13009,N_12467,N_12269);
and U13010 (N_13010,N_12214,N_12021);
or U13011 (N_13011,N_12529,N_12447);
nor U13012 (N_13012,N_12673,N_12423);
or U13013 (N_13013,N_12657,N_12677);
xnor U13014 (N_13014,N_12891,N_12372);
nor U13015 (N_13015,N_12281,N_12478);
nor U13016 (N_13016,N_12468,N_12514);
nor U13017 (N_13017,N_12609,N_12622);
xor U13018 (N_13018,N_12180,N_12111);
and U13019 (N_13019,N_12297,N_12414);
xnor U13020 (N_13020,N_12588,N_12678);
and U13021 (N_13021,N_12858,N_12191);
or U13022 (N_13022,N_12473,N_12133);
nand U13023 (N_13023,N_12538,N_12542);
or U13024 (N_13024,N_12357,N_12752);
and U13025 (N_13025,N_12863,N_12878);
nor U13026 (N_13026,N_12034,N_12759);
and U13027 (N_13027,N_12896,N_12639);
or U13028 (N_13028,N_12662,N_12483);
and U13029 (N_13029,N_12574,N_12193);
nand U13030 (N_13030,N_12317,N_12341);
nand U13031 (N_13031,N_12727,N_12918);
nor U13032 (N_13032,N_12807,N_12088);
nor U13033 (N_13033,N_12565,N_12108);
xor U13034 (N_13034,N_12746,N_12175);
nor U13035 (N_13035,N_12054,N_12448);
nor U13036 (N_13036,N_12121,N_12608);
nand U13037 (N_13037,N_12779,N_12131);
and U13038 (N_13038,N_12065,N_12235);
or U13039 (N_13039,N_12633,N_12917);
nor U13040 (N_13040,N_12390,N_12489);
nor U13041 (N_13041,N_12496,N_12391);
and U13042 (N_13042,N_12028,N_12450);
nand U13043 (N_13043,N_12969,N_12647);
and U13044 (N_13044,N_12910,N_12534);
or U13045 (N_13045,N_12334,N_12310);
or U13046 (N_13046,N_12646,N_12706);
xor U13047 (N_13047,N_12069,N_12063);
or U13048 (N_13048,N_12362,N_12796);
nor U13049 (N_13049,N_12000,N_12008);
nand U13050 (N_13050,N_12804,N_12707);
or U13051 (N_13051,N_12651,N_12562);
and U13052 (N_13052,N_12200,N_12304);
nor U13053 (N_13053,N_12217,N_12300);
and U13054 (N_13054,N_12479,N_12905);
nand U13055 (N_13055,N_12396,N_12454);
or U13056 (N_13056,N_12726,N_12405);
xor U13057 (N_13057,N_12937,N_12728);
nand U13058 (N_13058,N_12914,N_12603);
xnor U13059 (N_13059,N_12406,N_12455);
and U13060 (N_13060,N_12812,N_12619);
or U13061 (N_13061,N_12890,N_12652);
or U13062 (N_13062,N_12120,N_12747);
and U13063 (N_13063,N_12009,N_12501);
and U13064 (N_13064,N_12822,N_12995);
nand U13065 (N_13065,N_12254,N_12273);
or U13066 (N_13066,N_12466,N_12554);
or U13067 (N_13067,N_12295,N_12583);
nand U13068 (N_13068,N_12048,N_12664);
or U13069 (N_13069,N_12572,N_12909);
xor U13070 (N_13070,N_12298,N_12241);
or U13071 (N_13071,N_12083,N_12660);
nor U13072 (N_13072,N_12921,N_12550);
nand U13073 (N_13073,N_12680,N_12764);
xnor U13074 (N_13074,N_12844,N_12480);
and U13075 (N_13075,N_12799,N_12347);
nand U13076 (N_13076,N_12611,N_12685);
or U13077 (N_13077,N_12732,N_12027);
xnor U13078 (N_13078,N_12860,N_12306);
xor U13079 (N_13079,N_12838,N_12519);
nand U13080 (N_13080,N_12580,N_12547);
or U13081 (N_13081,N_12323,N_12990);
nor U13082 (N_13082,N_12490,N_12723);
nor U13083 (N_13083,N_12943,N_12299);
xnor U13084 (N_13084,N_12442,N_12753);
nor U13085 (N_13085,N_12950,N_12109);
xor U13086 (N_13086,N_12776,N_12687);
xor U13087 (N_13087,N_12928,N_12849);
nand U13088 (N_13088,N_12203,N_12958);
nand U13089 (N_13089,N_12865,N_12630);
or U13090 (N_13090,N_12744,N_12915);
or U13091 (N_13091,N_12020,N_12399);
or U13092 (N_13092,N_12135,N_12268);
nand U13093 (N_13093,N_12640,N_12183);
xor U13094 (N_13094,N_12582,N_12825);
nor U13095 (N_13095,N_12107,N_12612);
and U13096 (N_13096,N_12495,N_12951);
nand U13097 (N_13097,N_12102,N_12023);
and U13098 (N_13098,N_12335,N_12568);
nand U13099 (N_13099,N_12637,N_12190);
or U13100 (N_13100,N_12348,N_12907);
and U13101 (N_13101,N_12709,N_12518);
xnor U13102 (N_13102,N_12936,N_12079);
or U13103 (N_13103,N_12232,N_12174);
or U13104 (N_13104,N_12940,N_12982);
or U13105 (N_13105,N_12245,N_12201);
nor U13106 (N_13106,N_12381,N_12931);
xnor U13107 (N_13107,N_12618,N_12354);
or U13108 (N_13108,N_12096,N_12005);
and U13109 (N_13109,N_12117,N_12824);
or U13110 (N_13110,N_12368,N_12902);
or U13111 (N_13111,N_12531,N_12981);
nor U13112 (N_13112,N_12977,N_12826);
nor U13113 (N_13113,N_12967,N_12136);
nor U13114 (N_13114,N_12521,N_12654);
nand U13115 (N_13115,N_12409,N_12927);
nor U13116 (N_13116,N_12352,N_12702);
nand U13117 (N_13117,N_12094,N_12598);
nor U13118 (N_13118,N_12997,N_12557);
or U13119 (N_13119,N_12590,N_12388);
or U13120 (N_13120,N_12929,N_12146);
xor U13121 (N_13121,N_12333,N_12077);
and U13122 (N_13122,N_12867,N_12427);
xnor U13123 (N_13123,N_12340,N_12095);
and U13124 (N_13124,N_12041,N_12284);
or U13125 (N_13125,N_12326,N_12974);
xnor U13126 (N_13126,N_12104,N_12968);
nand U13127 (N_13127,N_12877,N_12179);
and U13128 (N_13128,N_12091,N_12738);
and U13129 (N_13129,N_12144,N_12266);
nor U13130 (N_13130,N_12426,N_12806);
xnor U13131 (N_13131,N_12003,N_12762);
and U13132 (N_13132,N_12563,N_12605);
nand U13133 (N_13133,N_12332,N_12591);
nand U13134 (N_13134,N_12274,N_12081);
or U13135 (N_13135,N_12503,N_12161);
or U13136 (N_13136,N_12827,N_12187);
or U13137 (N_13137,N_12432,N_12606);
xnor U13138 (N_13138,N_12551,N_12165);
and U13139 (N_13139,N_12404,N_12952);
nor U13140 (N_13140,N_12624,N_12528);
nand U13141 (N_13141,N_12830,N_12197);
nor U13142 (N_13142,N_12810,N_12443);
nand U13143 (N_13143,N_12820,N_12745);
or U13144 (N_13144,N_12780,N_12577);
and U13145 (N_13145,N_12434,N_12832);
xor U13146 (N_13146,N_12789,N_12979);
nand U13147 (N_13147,N_12567,N_12290);
or U13148 (N_13148,N_12586,N_12794);
and U13149 (N_13149,N_12893,N_12142);
or U13150 (N_13150,N_12944,N_12072);
xnor U13151 (N_13151,N_12970,N_12631);
nor U13152 (N_13152,N_12342,N_12512);
nor U13153 (N_13153,N_12036,N_12584);
nand U13154 (N_13154,N_12267,N_12697);
xnor U13155 (N_13155,N_12033,N_12437);
and U13156 (N_13156,N_12206,N_12643);
xnor U13157 (N_13157,N_12705,N_12155);
and U13158 (N_13158,N_12209,N_12996);
and U13159 (N_13159,N_12097,N_12634);
or U13160 (N_13160,N_12422,N_12338);
or U13161 (N_13161,N_12198,N_12387);
or U13162 (N_13162,N_12420,N_12162);
or U13163 (N_13163,N_12594,N_12684);
nand U13164 (N_13164,N_12171,N_12485);
or U13165 (N_13165,N_12258,N_12527);
nor U13166 (N_13166,N_12614,N_12576);
or U13167 (N_13167,N_12236,N_12213);
xor U13168 (N_13168,N_12816,N_12260);
xor U13169 (N_13169,N_12901,N_12540);
xnor U13170 (N_13170,N_12847,N_12470);
xnor U13171 (N_13171,N_12879,N_12708);
or U13172 (N_13172,N_12132,N_12163);
xnor U13173 (N_13173,N_12623,N_12526);
xor U13174 (N_13174,N_12415,N_12278);
or U13175 (N_13175,N_12945,N_12075);
nor U13176 (N_13176,N_12430,N_12872);
xor U13177 (N_13177,N_12785,N_12949);
nor U13178 (N_13178,N_12765,N_12148);
and U13179 (N_13179,N_12736,N_12895);
nand U13180 (N_13180,N_12889,N_12211);
nand U13181 (N_13181,N_12143,N_12972);
nand U13182 (N_13182,N_12749,N_12456);
nor U13183 (N_13183,N_12965,N_12441);
nor U13184 (N_13184,N_12989,N_12818);
nor U13185 (N_13185,N_12924,N_12755);
or U13186 (N_13186,N_12581,N_12038);
nor U13187 (N_13187,N_12821,N_12597);
nand U13188 (N_13188,N_12051,N_12181);
or U13189 (N_13189,N_12817,N_12313);
nor U13190 (N_13190,N_12815,N_12600);
and U13191 (N_13191,N_12057,N_12182);
xnor U13192 (N_13192,N_12463,N_12172);
or U13193 (N_13193,N_12122,N_12499);
nor U13194 (N_13194,N_12280,N_12115);
nor U13195 (N_13195,N_12641,N_12253);
nor U13196 (N_13196,N_12429,N_12316);
nand U13197 (N_13197,N_12164,N_12301);
or U13198 (N_13198,N_12841,N_12482);
nor U13199 (N_13199,N_12919,N_12243);
nand U13200 (N_13200,N_12963,N_12150);
nand U13201 (N_13201,N_12375,N_12536);
nor U13202 (N_13202,N_12668,N_12460);
and U13203 (N_13203,N_12411,N_12419);
and U13204 (N_13204,N_12066,N_12007);
nor U13205 (N_13205,N_12371,N_12322);
xnor U13206 (N_13206,N_12595,N_12792);
xor U13207 (N_13207,N_12226,N_12991);
xnor U13208 (N_13208,N_12119,N_12801);
xor U13209 (N_13209,N_12436,N_12740);
xnor U13210 (N_13210,N_12558,N_12229);
nand U13211 (N_13211,N_12032,N_12711);
nand U13212 (N_13212,N_12575,N_12186);
nor U13213 (N_13213,N_12899,N_12541);
xor U13214 (N_13214,N_12741,N_12089);
xnor U13215 (N_13215,N_12569,N_12848);
nor U13216 (N_13216,N_12683,N_12410);
and U13217 (N_13217,N_12670,N_12282);
and U13218 (N_13218,N_12380,N_12166);
nand U13219 (N_13219,N_12843,N_12870);
xor U13220 (N_13220,N_12461,N_12855);
and U13221 (N_13221,N_12486,N_12625);
and U13222 (N_13222,N_12800,N_12758);
nand U13223 (N_13223,N_12398,N_12768);
nor U13224 (N_13224,N_12658,N_12445);
xor U13225 (N_13225,N_12085,N_12386);
or U13226 (N_13226,N_12986,N_12644);
or U13227 (N_13227,N_12733,N_12249);
and U13228 (N_13228,N_12339,N_12189);
nor U13229 (N_13229,N_12735,N_12355);
and U13230 (N_13230,N_12270,N_12067);
nand U13231 (N_13231,N_12882,N_12472);
nor U13232 (N_13232,N_12070,N_12681);
and U13233 (N_13233,N_12731,N_12192);
or U13234 (N_13234,N_12345,N_12234);
nor U13235 (N_13235,N_12864,N_12215);
and U13236 (N_13236,N_12916,N_12655);
nand U13237 (N_13237,N_12045,N_12359);
nand U13238 (N_13238,N_12845,N_12992);
nor U13239 (N_13239,N_12857,N_12022);
nand U13240 (N_13240,N_12440,N_12154);
nor U13241 (N_13241,N_12138,N_12418);
nand U13242 (N_13242,N_12932,N_12648);
xnor U13243 (N_13243,N_12856,N_12327);
xor U13244 (N_13244,N_12767,N_12058);
or U13245 (N_13245,N_12823,N_12199);
nand U13246 (N_13246,N_12987,N_12859);
nor U13247 (N_13247,N_12365,N_12725);
and U13248 (N_13248,N_12465,N_12052);
nand U13249 (N_13249,N_12993,N_12178);
and U13250 (N_13250,N_12222,N_12311);
xor U13251 (N_13251,N_12659,N_12185);
nor U13252 (N_13252,N_12261,N_12988);
nand U13253 (N_13253,N_12113,N_12263);
or U13254 (N_13254,N_12530,N_12378);
nand U13255 (N_13255,N_12701,N_12498);
or U13256 (N_13256,N_12137,N_12960);
nand U13257 (N_13257,N_12720,N_12509);
nand U13258 (N_13258,N_12044,N_12888);
or U13259 (N_13259,N_12686,N_12975);
nor U13260 (N_13260,N_12934,N_12803);
or U13261 (N_13261,N_12385,N_12082);
nand U13262 (N_13262,N_12477,N_12956);
or U13263 (N_13263,N_12688,N_12016);
xor U13264 (N_13264,N_12307,N_12237);
and U13265 (N_13265,N_12862,N_12961);
xnor U13266 (N_13266,N_12769,N_12560);
nor U13267 (N_13267,N_12129,N_12152);
xnor U13268 (N_13268,N_12204,N_12689);
or U13269 (N_13269,N_12238,N_12556);
and U13270 (N_13270,N_12101,N_12971);
xnor U13271 (N_13271,N_12959,N_12431);
or U13272 (N_13272,N_12805,N_12656);
or U13273 (N_13273,N_12004,N_12632);
and U13274 (N_13274,N_12545,N_12840);
nor U13275 (N_13275,N_12739,N_12302);
xor U13276 (N_13276,N_12105,N_12885);
and U13277 (N_13277,N_12369,N_12231);
nand U13278 (N_13278,N_12839,N_12087);
and U13279 (N_13279,N_12698,N_12046);
nor U13280 (N_13280,N_12771,N_12283);
nand U13281 (N_13281,N_12544,N_12195);
nand U13282 (N_13282,N_12176,N_12694);
and U13283 (N_13283,N_12602,N_12252);
xor U13284 (N_13284,N_12080,N_12124);
nor U13285 (N_13285,N_12230,N_12444);
or U13286 (N_13286,N_12853,N_12886);
nor U13287 (N_13287,N_12086,N_12566);
nand U13288 (N_13288,N_12358,N_12285);
nand U13289 (N_13289,N_12911,N_12118);
xnor U13290 (N_13290,N_12819,N_12715);
or U13291 (N_13291,N_12320,N_12695);
xnor U13292 (N_13292,N_12106,N_12828);
nand U13293 (N_13293,N_12255,N_12220);
and U13294 (N_13294,N_12050,N_12887);
or U13295 (N_13295,N_12246,N_12130);
xor U13296 (N_13296,N_12787,N_12056);
nand U13297 (N_13297,N_12103,N_12766);
or U13298 (N_13298,N_12312,N_12535);
xor U13299 (N_13299,N_12294,N_12939);
or U13300 (N_13300,N_12453,N_12025);
xor U13301 (N_13301,N_12247,N_12601);
and U13302 (N_13302,N_12330,N_12329);
nor U13303 (N_13303,N_12791,N_12265);
or U13304 (N_13304,N_12999,N_12653);
and U13305 (N_13305,N_12168,N_12754);
nor U13306 (N_13306,N_12693,N_12328);
and U13307 (N_13307,N_12589,N_12868);
nor U13308 (N_13308,N_12402,N_12510);
nand U13309 (N_13309,N_12424,N_12153);
xor U13310 (N_13310,N_12484,N_12059);
or U13311 (N_13311,N_12403,N_12876);
or U13312 (N_13312,N_12718,N_12880);
or U13313 (N_13313,N_12256,N_12384);
xnor U13314 (N_13314,N_12691,N_12679);
nand U13315 (N_13315,N_12833,N_12373);
and U13316 (N_13316,N_12098,N_12325);
nor U13317 (N_13317,N_12305,N_12781);
xor U13318 (N_13318,N_12721,N_12356);
nand U13319 (N_13319,N_12464,N_12704);
and U13320 (N_13320,N_12599,N_12293);
nand U13321 (N_13321,N_12628,N_12433);
nor U13322 (N_13322,N_12713,N_12957);
xor U13323 (N_13323,N_12128,N_12397);
or U13324 (N_13324,N_12846,N_12092);
or U13325 (N_13325,N_12935,N_12053);
xnor U13326 (N_13326,N_12922,N_12714);
or U13327 (N_13327,N_12829,N_12157);
or U13328 (N_13328,N_12134,N_12401);
nand U13329 (N_13329,N_12763,N_12446);
nand U13330 (N_13330,N_12458,N_12552);
nor U13331 (N_13331,N_12474,N_12425);
nor U13332 (N_13332,N_12983,N_12699);
xnor U13333 (N_13333,N_12438,N_12978);
or U13334 (N_13334,N_12497,N_12607);
and U13335 (N_13335,N_12672,N_12126);
or U13336 (N_13336,N_12795,N_12170);
or U13337 (N_13337,N_12507,N_12522);
and U13338 (N_13338,N_12227,N_12884);
and U13339 (N_13339,N_12516,N_12636);
nor U13340 (N_13340,N_12060,N_12913);
nor U13341 (N_13341,N_12296,N_12188);
and U13342 (N_13342,N_12629,N_12650);
xor U13343 (N_13343,N_12850,N_12871);
nor U13344 (N_13344,N_12012,N_12084);
nand U13345 (N_13345,N_12376,N_12233);
xor U13346 (N_13346,N_12015,N_12842);
and U13347 (N_13347,N_12955,N_12116);
and U13348 (N_13348,N_12515,N_12364);
nor U13349 (N_13349,N_12292,N_12757);
or U13350 (N_13350,N_12585,N_12035);
and U13351 (N_13351,N_12377,N_12219);
and U13352 (N_13352,N_12750,N_12579);
or U13353 (N_13353,N_12620,N_12156);
or U13354 (N_13354,N_12331,N_12546);
nand U13355 (N_13355,N_12775,N_12537);
nor U13356 (N_13356,N_12147,N_12047);
nand U13357 (N_13357,N_12271,N_12571);
or U13358 (N_13358,N_12360,N_12114);
xnor U13359 (N_13359,N_12221,N_12242);
nand U13360 (N_13360,N_12941,N_12523);
and U13361 (N_13361,N_12517,N_12006);
xnor U13362 (N_13362,N_12262,N_12548);
xnor U13363 (N_13363,N_12883,N_12553);
xor U13364 (N_13364,N_12346,N_12774);
xnor U13365 (N_13365,N_12488,N_12017);
or U13366 (N_13366,N_12064,N_12370);
and U13367 (N_13367,N_12835,N_12898);
nor U13368 (N_13368,N_12866,N_12288);
nor U13369 (N_13369,N_12742,N_12207);
or U13370 (N_13370,N_12511,N_12014);
nand U13371 (N_13371,N_12225,N_12149);
and U13372 (N_13372,N_12451,N_12013);
nand U13373 (N_13373,N_12493,N_12475);
and U13374 (N_13374,N_12502,N_12194);
nand U13375 (N_13375,N_12904,N_12861);
xnor U13376 (N_13376,N_12994,N_12169);
nor U13377 (N_13377,N_12457,N_12324);
nor U13378 (N_13378,N_12090,N_12491);
nor U13379 (N_13379,N_12287,N_12786);
or U13380 (N_13380,N_12894,N_12039);
and U13381 (N_13381,N_12412,N_12773);
and U13382 (N_13382,N_12793,N_12349);
or U13383 (N_13383,N_12321,N_12788);
nor U13384 (N_13384,N_12966,N_12615);
or U13385 (N_13385,N_12906,N_12948);
nor U13386 (N_13386,N_12112,N_12802);
nand U13387 (N_13387,N_12223,N_12811);
or U13388 (N_13388,N_12923,N_12462);
nor U13389 (N_13389,N_12782,N_12407);
nor U13390 (N_13390,N_12145,N_12814);
and U13391 (N_13391,N_12210,N_12635);
xnor U13392 (N_13392,N_12073,N_12587);
or U13393 (N_13393,N_12953,N_12690);
and U13394 (N_13394,N_12055,N_12353);
nand U13395 (N_13395,N_12383,N_12874);
nand U13396 (N_13396,N_12596,N_12205);
and U13397 (N_13397,N_12881,N_12665);
nor U13398 (N_13398,N_12734,N_12616);
or U13399 (N_13399,N_12314,N_12676);
nand U13400 (N_13400,N_12318,N_12366);
and U13401 (N_13401,N_12703,N_12627);
and U13402 (N_13402,N_12001,N_12029);
or U13403 (N_13403,N_12513,N_12748);
xor U13404 (N_13404,N_12700,N_12421);
nand U13405 (N_13405,N_12024,N_12291);
or U13406 (N_13406,N_12184,N_12533);
xnor U13407 (N_13407,N_12277,N_12481);
nor U13408 (N_13408,N_12239,N_12011);
nand U13409 (N_13409,N_12177,N_12492);
and U13410 (N_13410,N_12696,N_12869);
xor U13411 (N_13411,N_12716,N_12408);
nand U13412 (N_13412,N_12250,N_12671);
or U13413 (N_13413,N_12240,N_12854);
nand U13414 (N_13414,N_12962,N_12040);
and U13415 (N_13415,N_12675,N_12487);
nor U13416 (N_13416,N_12626,N_12520);
nand U13417 (N_13417,N_12980,N_12062);
or U13418 (N_13418,N_12140,N_12836);
and U13419 (N_13419,N_12667,N_12770);
nand U13420 (N_13420,N_12760,N_12573);
xor U13421 (N_13421,N_12272,N_12010);
nand U13422 (N_13422,N_12724,N_12363);
xor U13423 (N_13423,N_12798,N_12617);
nand U13424 (N_13424,N_12336,N_12043);
nand U13425 (N_13425,N_12279,N_12722);
xor U13426 (N_13426,N_12208,N_12337);
or U13427 (N_13427,N_12524,N_12784);
and U13428 (N_13428,N_12315,N_12400);
xnor U13429 (N_13429,N_12613,N_12167);
or U13430 (N_13430,N_12351,N_12938);
xnor U13431 (N_13431,N_12797,N_12710);
and U13432 (N_13432,N_12099,N_12417);
and U13433 (N_13433,N_12674,N_12031);
nand U13434 (N_13434,N_12834,N_12561);
nor U13435 (N_13435,N_12439,N_12508);
nor U13436 (N_13436,N_12663,N_12808);
or U13437 (N_13437,N_12309,N_12692);
nor U13438 (N_13438,N_12549,N_12218);
and U13439 (N_13439,N_12151,N_12160);
nor U13440 (N_13440,N_12393,N_12505);
xor U13441 (N_13441,N_12139,N_12778);
and U13442 (N_13442,N_12303,N_12998);
or U13443 (N_13443,N_12539,N_12264);
or U13444 (N_13444,N_12946,N_12942);
xnor U13445 (N_13445,N_12244,N_12228);
nor U13446 (N_13446,N_12382,N_12248);
and U13447 (N_13447,N_12413,N_12873);
xor U13448 (N_13448,N_12428,N_12964);
nand U13449 (N_13449,N_12761,N_12350);
nor U13450 (N_13450,N_12621,N_12892);
xor U13451 (N_13451,N_12730,N_12173);
nor U13452 (N_13452,N_12379,N_12071);
nand U13453 (N_13453,N_12259,N_12093);
nor U13454 (N_13454,N_12500,N_12912);
xnor U13455 (N_13455,N_12343,N_12389);
nand U13456 (N_13456,N_12049,N_12926);
xor U13457 (N_13457,N_12308,N_12459);
and U13458 (N_13458,N_12159,N_12592);
nor U13459 (N_13459,N_12212,N_12319);
nand U13460 (N_13460,N_12875,N_12026);
xnor U13461 (N_13461,N_12908,N_12374);
nand U13462 (N_13462,N_12019,N_12018);
and U13463 (N_13463,N_12669,N_12506);
or U13464 (N_13464,N_12361,N_12638);
nand U13465 (N_13465,N_12666,N_12604);
and U13466 (N_13466,N_12719,N_12790);
or U13467 (N_13467,N_12559,N_12743);
nand U13468 (N_13468,N_12394,N_12930);
xor U13469 (N_13469,N_12471,N_12494);
or U13470 (N_13470,N_12476,N_12074);
xnor U13471 (N_13471,N_12078,N_12395);
nor U13472 (N_13472,N_12831,N_12985);
and U13473 (N_13473,N_12202,N_12593);
nor U13474 (N_13474,N_12717,N_12852);
nand U13475 (N_13475,N_12682,N_12837);
and U13476 (N_13476,N_12076,N_12555);
nand U13477 (N_13477,N_12042,N_12954);
or U13478 (N_13478,N_12925,N_12286);
nand U13479 (N_13479,N_12452,N_12276);
or U13480 (N_13480,N_12610,N_12543);
xor U13481 (N_13481,N_12037,N_12645);
and U13482 (N_13482,N_12224,N_12897);
and U13483 (N_13483,N_12532,N_12642);
nor U13484 (N_13484,N_12416,N_12947);
xnor U13485 (N_13485,N_12289,N_12920);
nor U13486 (N_13486,N_12504,N_12649);
xnor U13487 (N_13487,N_12216,N_12251);
nor U13488 (N_13488,N_12712,N_12141);
or U13489 (N_13489,N_12002,N_12275);
nor U13490 (N_13490,N_12030,N_12392);
nand U13491 (N_13491,N_12257,N_12783);
or U13492 (N_13492,N_12903,N_12933);
or U13493 (N_13493,N_12976,N_12813);
and U13494 (N_13494,N_12196,N_12772);
and U13495 (N_13495,N_12127,N_12570);
xor U13496 (N_13496,N_12564,N_12110);
and U13497 (N_13497,N_12973,N_12809);
nand U13498 (N_13498,N_12751,N_12100);
xor U13499 (N_13499,N_12068,N_12900);
or U13500 (N_13500,N_12902,N_12037);
nand U13501 (N_13501,N_12715,N_12931);
nor U13502 (N_13502,N_12550,N_12272);
xnor U13503 (N_13503,N_12342,N_12093);
and U13504 (N_13504,N_12424,N_12653);
or U13505 (N_13505,N_12567,N_12376);
or U13506 (N_13506,N_12074,N_12934);
and U13507 (N_13507,N_12041,N_12617);
nor U13508 (N_13508,N_12896,N_12470);
nand U13509 (N_13509,N_12983,N_12819);
xnor U13510 (N_13510,N_12878,N_12555);
and U13511 (N_13511,N_12333,N_12136);
and U13512 (N_13512,N_12317,N_12601);
nor U13513 (N_13513,N_12248,N_12921);
xor U13514 (N_13514,N_12346,N_12813);
nand U13515 (N_13515,N_12616,N_12533);
xor U13516 (N_13516,N_12099,N_12936);
or U13517 (N_13517,N_12037,N_12434);
nand U13518 (N_13518,N_12150,N_12951);
nand U13519 (N_13519,N_12490,N_12032);
xor U13520 (N_13520,N_12803,N_12328);
xor U13521 (N_13521,N_12103,N_12414);
nand U13522 (N_13522,N_12068,N_12401);
and U13523 (N_13523,N_12098,N_12480);
xor U13524 (N_13524,N_12871,N_12598);
xor U13525 (N_13525,N_12812,N_12589);
and U13526 (N_13526,N_12353,N_12712);
or U13527 (N_13527,N_12140,N_12859);
xor U13528 (N_13528,N_12582,N_12804);
or U13529 (N_13529,N_12229,N_12131);
xor U13530 (N_13530,N_12574,N_12256);
or U13531 (N_13531,N_12754,N_12904);
xor U13532 (N_13532,N_12981,N_12471);
and U13533 (N_13533,N_12409,N_12416);
nor U13534 (N_13534,N_12724,N_12581);
nor U13535 (N_13535,N_12759,N_12906);
nor U13536 (N_13536,N_12816,N_12030);
nand U13537 (N_13537,N_12650,N_12215);
nand U13538 (N_13538,N_12013,N_12314);
nand U13539 (N_13539,N_12287,N_12710);
xnor U13540 (N_13540,N_12630,N_12390);
nor U13541 (N_13541,N_12889,N_12759);
xnor U13542 (N_13542,N_12869,N_12268);
nand U13543 (N_13543,N_12875,N_12286);
nor U13544 (N_13544,N_12058,N_12620);
xnor U13545 (N_13545,N_12179,N_12144);
and U13546 (N_13546,N_12066,N_12868);
nand U13547 (N_13547,N_12162,N_12964);
and U13548 (N_13548,N_12457,N_12705);
or U13549 (N_13549,N_12609,N_12469);
and U13550 (N_13550,N_12080,N_12445);
nor U13551 (N_13551,N_12036,N_12429);
nand U13552 (N_13552,N_12172,N_12254);
or U13553 (N_13553,N_12583,N_12344);
or U13554 (N_13554,N_12393,N_12030);
xnor U13555 (N_13555,N_12698,N_12454);
and U13556 (N_13556,N_12990,N_12689);
nor U13557 (N_13557,N_12381,N_12707);
and U13558 (N_13558,N_12443,N_12556);
xnor U13559 (N_13559,N_12445,N_12179);
nand U13560 (N_13560,N_12942,N_12913);
or U13561 (N_13561,N_12379,N_12359);
nor U13562 (N_13562,N_12563,N_12083);
or U13563 (N_13563,N_12276,N_12919);
nand U13564 (N_13564,N_12397,N_12313);
or U13565 (N_13565,N_12533,N_12001);
nand U13566 (N_13566,N_12843,N_12138);
or U13567 (N_13567,N_12565,N_12538);
and U13568 (N_13568,N_12291,N_12636);
nor U13569 (N_13569,N_12502,N_12861);
xor U13570 (N_13570,N_12106,N_12207);
and U13571 (N_13571,N_12134,N_12525);
xor U13572 (N_13572,N_12975,N_12190);
nand U13573 (N_13573,N_12735,N_12902);
nand U13574 (N_13574,N_12241,N_12254);
xnor U13575 (N_13575,N_12834,N_12478);
xnor U13576 (N_13576,N_12792,N_12227);
nor U13577 (N_13577,N_12262,N_12170);
and U13578 (N_13578,N_12178,N_12845);
nand U13579 (N_13579,N_12322,N_12011);
xnor U13580 (N_13580,N_12597,N_12591);
nand U13581 (N_13581,N_12661,N_12090);
xnor U13582 (N_13582,N_12307,N_12113);
xor U13583 (N_13583,N_12877,N_12191);
and U13584 (N_13584,N_12839,N_12346);
and U13585 (N_13585,N_12675,N_12127);
xor U13586 (N_13586,N_12115,N_12294);
xnor U13587 (N_13587,N_12528,N_12902);
xor U13588 (N_13588,N_12615,N_12891);
nand U13589 (N_13589,N_12798,N_12765);
and U13590 (N_13590,N_12074,N_12616);
xnor U13591 (N_13591,N_12983,N_12576);
nor U13592 (N_13592,N_12251,N_12794);
and U13593 (N_13593,N_12036,N_12006);
or U13594 (N_13594,N_12048,N_12582);
xor U13595 (N_13595,N_12629,N_12432);
xnor U13596 (N_13596,N_12008,N_12431);
nand U13597 (N_13597,N_12318,N_12861);
xnor U13598 (N_13598,N_12732,N_12883);
and U13599 (N_13599,N_12106,N_12842);
and U13600 (N_13600,N_12792,N_12000);
or U13601 (N_13601,N_12879,N_12433);
xnor U13602 (N_13602,N_12584,N_12753);
nand U13603 (N_13603,N_12969,N_12797);
and U13604 (N_13604,N_12750,N_12289);
nand U13605 (N_13605,N_12011,N_12136);
nand U13606 (N_13606,N_12095,N_12060);
nand U13607 (N_13607,N_12374,N_12128);
nand U13608 (N_13608,N_12321,N_12323);
nand U13609 (N_13609,N_12448,N_12987);
and U13610 (N_13610,N_12278,N_12717);
nor U13611 (N_13611,N_12402,N_12399);
nor U13612 (N_13612,N_12134,N_12097);
nand U13613 (N_13613,N_12813,N_12043);
nor U13614 (N_13614,N_12781,N_12522);
xor U13615 (N_13615,N_12310,N_12320);
and U13616 (N_13616,N_12014,N_12980);
or U13617 (N_13617,N_12178,N_12352);
xor U13618 (N_13618,N_12192,N_12299);
nor U13619 (N_13619,N_12494,N_12891);
nor U13620 (N_13620,N_12070,N_12355);
nor U13621 (N_13621,N_12722,N_12247);
xor U13622 (N_13622,N_12947,N_12127);
nor U13623 (N_13623,N_12689,N_12742);
nand U13624 (N_13624,N_12778,N_12651);
nor U13625 (N_13625,N_12373,N_12505);
nor U13626 (N_13626,N_12132,N_12495);
or U13627 (N_13627,N_12815,N_12345);
nand U13628 (N_13628,N_12660,N_12246);
and U13629 (N_13629,N_12876,N_12455);
or U13630 (N_13630,N_12584,N_12811);
and U13631 (N_13631,N_12988,N_12064);
or U13632 (N_13632,N_12055,N_12826);
nand U13633 (N_13633,N_12807,N_12122);
nand U13634 (N_13634,N_12086,N_12677);
nor U13635 (N_13635,N_12338,N_12598);
nand U13636 (N_13636,N_12130,N_12610);
xnor U13637 (N_13637,N_12383,N_12038);
nand U13638 (N_13638,N_12885,N_12614);
or U13639 (N_13639,N_12898,N_12663);
xnor U13640 (N_13640,N_12720,N_12688);
nor U13641 (N_13641,N_12963,N_12394);
and U13642 (N_13642,N_12498,N_12740);
nor U13643 (N_13643,N_12510,N_12015);
xor U13644 (N_13644,N_12524,N_12442);
or U13645 (N_13645,N_12500,N_12010);
and U13646 (N_13646,N_12214,N_12097);
nor U13647 (N_13647,N_12694,N_12937);
or U13648 (N_13648,N_12339,N_12080);
nand U13649 (N_13649,N_12618,N_12920);
xnor U13650 (N_13650,N_12085,N_12509);
and U13651 (N_13651,N_12605,N_12192);
or U13652 (N_13652,N_12242,N_12136);
or U13653 (N_13653,N_12350,N_12777);
xor U13654 (N_13654,N_12094,N_12398);
nand U13655 (N_13655,N_12804,N_12477);
xnor U13656 (N_13656,N_12252,N_12528);
nor U13657 (N_13657,N_12882,N_12718);
nand U13658 (N_13658,N_12405,N_12677);
nor U13659 (N_13659,N_12887,N_12117);
or U13660 (N_13660,N_12668,N_12101);
or U13661 (N_13661,N_12729,N_12433);
or U13662 (N_13662,N_12658,N_12209);
nor U13663 (N_13663,N_12120,N_12410);
and U13664 (N_13664,N_12836,N_12389);
nand U13665 (N_13665,N_12440,N_12216);
nand U13666 (N_13666,N_12627,N_12096);
and U13667 (N_13667,N_12522,N_12893);
xor U13668 (N_13668,N_12986,N_12409);
nand U13669 (N_13669,N_12906,N_12453);
nor U13670 (N_13670,N_12147,N_12503);
and U13671 (N_13671,N_12324,N_12727);
and U13672 (N_13672,N_12866,N_12647);
nor U13673 (N_13673,N_12747,N_12483);
nor U13674 (N_13674,N_12232,N_12392);
xnor U13675 (N_13675,N_12271,N_12724);
and U13676 (N_13676,N_12601,N_12584);
xnor U13677 (N_13677,N_12544,N_12987);
nand U13678 (N_13678,N_12242,N_12022);
and U13679 (N_13679,N_12169,N_12084);
nand U13680 (N_13680,N_12706,N_12592);
nand U13681 (N_13681,N_12050,N_12288);
and U13682 (N_13682,N_12328,N_12261);
nor U13683 (N_13683,N_12748,N_12862);
nor U13684 (N_13684,N_12152,N_12734);
nand U13685 (N_13685,N_12631,N_12607);
and U13686 (N_13686,N_12613,N_12585);
and U13687 (N_13687,N_12223,N_12260);
or U13688 (N_13688,N_12540,N_12814);
or U13689 (N_13689,N_12789,N_12191);
nand U13690 (N_13690,N_12995,N_12427);
and U13691 (N_13691,N_12149,N_12083);
xnor U13692 (N_13692,N_12736,N_12910);
nor U13693 (N_13693,N_12768,N_12548);
xor U13694 (N_13694,N_12442,N_12329);
nand U13695 (N_13695,N_12701,N_12111);
nor U13696 (N_13696,N_12379,N_12836);
nor U13697 (N_13697,N_12315,N_12655);
nor U13698 (N_13698,N_12605,N_12277);
and U13699 (N_13699,N_12915,N_12900);
nor U13700 (N_13700,N_12608,N_12088);
or U13701 (N_13701,N_12911,N_12447);
xor U13702 (N_13702,N_12436,N_12524);
nand U13703 (N_13703,N_12302,N_12692);
nor U13704 (N_13704,N_12311,N_12834);
nand U13705 (N_13705,N_12188,N_12706);
nand U13706 (N_13706,N_12901,N_12763);
xor U13707 (N_13707,N_12596,N_12120);
nor U13708 (N_13708,N_12657,N_12558);
nand U13709 (N_13709,N_12284,N_12713);
nand U13710 (N_13710,N_12182,N_12561);
xnor U13711 (N_13711,N_12909,N_12831);
nand U13712 (N_13712,N_12872,N_12146);
xnor U13713 (N_13713,N_12688,N_12088);
nor U13714 (N_13714,N_12864,N_12169);
nor U13715 (N_13715,N_12149,N_12577);
nor U13716 (N_13716,N_12178,N_12535);
nand U13717 (N_13717,N_12058,N_12112);
nor U13718 (N_13718,N_12682,N_12468);
and U13719 (N_13719,N_12630,N_12146);
or U13720 (N_13720,N_12674,N_12645);
nor U13721 (N_13721,N_12102,N_12613);
nor U13722 (N_13722,N_12018,N_12357);
nor U13723 (N_13723,N_12424,N_12374);
xor U13724 (N_13724,N_12419,N_12821);
xnor U13725 (N_13725,N_12389,N_12096);
and U13726 (N_13726,N_12166,N_12560);
nor U13727 (N_13727,N_12798,N_12847);
or U13728 (N_13728,N_12993,N_12553);
xor U13729 (N_13729,N_12173,N_12472);
nand U13730 (N_13730,N_12492,N_12939);
or U13731 (N_13731,N_12646,N_12361);
and U13732 (N_13732,N_12305,N_12678);
or U13733 (N_13733,N_12107,N_12161);
or U13734 (N_13734,N_12276,N_12468);
nand U13735 (N_13735,N_12990,N_12700);
or U13736 (N_13736,N_12114,N_12418);
nor U13737 (N_13737,N_12025,N_12663);
and U13738 (N_13738,N_12737,N_12628);
nand U13739 (N_13739,N_12665,N_12228);
and U13740 (N_13740,N_12870,N_12494);
nand U13741 (N_13741,N_12488,N_12117);
xnor U13742 (N_13742,N_12284,N_12130);
nand U13743 (N_13743,N_12586,N_12131);
and U13744 (N_13744,N_12722,N_12486);
xor U13745 (N_13745,N_12493,N_12000);
nor U13746 (N_13746,N_12326,N_12503);
nor U13747 (N_13747,N_12450,N_12608);
xor U13748 (N_13748,N_12752,N_12107);
nand U13749 (N_13749,N_12823,N_12995);
nor U13750 (N_13750,N_12451,N_12599);
nor U13751 (N_13751,N_12313,N_12188);
xnor U13752 (N_13752,N_12059,N_12912);
and U13753 (N_13753,N_12494,N_12962);
and U13754 (N_13754,N_12965,N_12533);
nor U13755 (N_13755,N_12382,N_12315);
xor U13756 (N_13756,N_12172,N_12239);
xnor U13757 (N_13757,N_12391,N_12477);
nor U13758 (N_13758,N_12553,N_12047);
nand U13759 (N_13759,N_12786,N_12983);
nor U13760 (N_13760,N_12553,N_12363);
nor U13761 (N_13761,N_12072,N_12910);
or U13762 (N_13762,N_12139,N_12999);
nor U13763 (N_13763,N_12747,N_12693);
nand U13764 (N_13764,N_12130,N_12538);
nand U13765 (N_13765,N_12120,N_12191);
nand U13766 (N_13766,N_12012,N_12248);
nand U13767 (N_13767,N_12418,N_12071);
or U13768 (N_13768,N_12550,N_12378);
xnor U13769 (N_13769,N_12614,N_12998);
and U13770 (N_13770,N_12364,N_12528);
nand U13771 (N_13771,N_12834,N_12993);
xor U13772 (N_13772,N_12007,N_12137);
xor U13773 (N_13773,N_12036,N_12578);
or U13774 (N_13774,N_12889,N_12616);
nand U13775 (N_13775,N_12167,N_12929);
nor U13776 (N_13776,N_12751,N_12972);
xor U13777 (N_13777,N_12680,N_12035);
or U13778 (N_13778,N_12187,N_12136);
and U13779 (N_13779,N_12847,N_12833);
xor U13780 (N_13780,N_12269,N_12077);
and U13781 (N_13781,N_12647,N_12045);
xor U13782 (N_13782,N_12759,N_12903);
or U13783 (N_13783,N_12646,N_12955);
and U13784 (N_13784,N_12915,N_12138);
or U13785 (N_13785,N_12852,N_12458);
or U13786 (N_13786,N_12804,N_12833);
nor U13787 (N_13787,N_12826,N_12137);
and U13788 (N_13788,N_12657,N_12394);
xnor U13789 (N_13789,N_12194,N_12256);
and U13790 (N_13790,N_12750,N_12801);
and U13791 (N_13791,N_12666,N_12696);
nor U13792 (N_13792,N_12604,N_12063);
and U13793 (N_13793,N_12703,N_12571);
nand U13794 (N_13794,N_12068,N_12542);
or U13795 (N_13795,N_12371,N_12283);
and U13796 (N_13796,N_12798,N_12233);
or U13797 (N_13797,N_12443,N_12095);
or U13798 (N_13798,N_12260,N_12192);
and U13799 (N_13799,N_12917,N_12687);
nand U13800 (N_13800,N_12390,N_12948);
xnor U13801 (N_13801,N_12366,N_12247);
or U13802 (N_13802,N_12095,N_12994);
or U13803 (N_13803,N_12844,N_12132);
nand U13804 (N_13804,N_12477,N_12309);
nand U13805 (N_13805,N_12096,N_12399);
nor U13806 (N_13806,N_12531,N_12927);
nand U13807 (N_13807,N_12457,N_12279);
and U13808 (N_13808,N_12680,N_12650);
and U13809 (N_13809,N_12593,N_12901);
nor U13810 (N_13810,N_12836,N_12818);
and U13811 (N_13811,N_12363,N_12012);
and U13812 (N_13812,N_12055,N_12091);
or U13813 (N_13813,N_12020,N_12281);
or U13814 (N_13814,N_12428,N_12890);
and U13815 (N_13815,N_12858,N_12568);
or U13816 (N_13816,N_12672,N_12881);
or U13817 (N_13817,N_12862,N_12559);
and U13818 (N_13818,N_12558,N_12782);
xor U13819 (N_13819,N_12681,N_12127);
nand U13820 (N_13820,N_12237,N_12377);
and U13821 (N_13821,N_12133,N_12517);
nor U13822 (N_13822,N_12229,N_12582);
xnor U13823 (N_13823,N_12781,N_12158);
and U13824 (N_13824,N_12576,N_12414);
or U13825 (N_13825,N_12202,N_12061);
nand U13826 (N_13826,N_12333,N_12682);
or U13827 (N_13827,N_12318,N_12929);
and U13828 (N_13828,N_12258,N_12597);
nand U13829 (N_13829,N_12794,N_12615);
nor U13830 (N_13830,N_12119,N_12813);
and U13831 (N_13831,N_12396,N_12546);
or U13832 (N_13832,N_12541,N_12573);
xnor U13833 (N_13833,N_12500,N_12457);
nand U13834 (N_13834,N_12106,N_12185);
or U13835 (N_13835,N_12786,N_12242);
nor U13836 (N_13836,N_12627,N_12763);
and U13837 (N_13837,N_12924,N_12124);
xor U13838 (N_13838,N_12170,N_12099);
nand U13839 (N_13839,N_12575,N_12481);
nand U13840 (N_13840,N_12138,N_12571);
and U13841 (N_13841,N_12674,N_12091);
nor U13842 (N_13842,N_12217,N_12388);
xor U13843 (N_13843,N_12666,N_12770);
nand U13844 (N_13844,N_12014,N_12434);
nor U13845 (N_13845,N_12257,N_12397);
or U13846 (N_13846,N_12460,N_12880);
or U13847 (N_13847,N_12649,N_12840);
and U13848 (N_13848,N_12566,N_12028);
nand U13849 (N_13849,N_12532,N_12796);
xor U13850 (N_13850,N_12433,N_12382);
or U13851 (N_13851,N_12538,N_12783);
nand U13852 (N_13852,N_12239,N_12129);
and U13853 (N_13853,N_12746,N_12110);
and U13854 (N_13854,N_12006,N_12211);
nand U13855 (N_13855,N_12011,N_12170);
and U13856 (N_13856,N_12762,N_12937);
xnor U13857 (N_13857,N_12369,N_12451);
and U13858 (N_13858,N_12597,N_12743);
xnor U13859 (N_13859,N_12308,N_12391);
xor U13860 (N_13860,N_12007,N_12256);
and U13861 (N_13861,N_12021,N_12219);
nor U13862 (N_13862,N_12708,N_12548);
xor U13863 (N_13863,N_12072,N_12510);
xnor U13864 (N_13864,N_12781,N_12871);
or U13865 (N_13865,N_12871,N_12525);
nand U13866 (N_13866,N_12208,N_12486);
or U13867 (N_13867,N_12140,N_12877);
xor U13868 (N_13868,N_12871,N_12227);
nor U13869 (N_13869,N_12240,N_12820);
xor U13870 (N_13870,N_12637,N_12571);
or U13871 (N_13871,N_12714,N_12394);
nor U13872 (N_13872,N_12553,N_12665);
nor U13873 (N_13873,N_12382,N_12337);
xnor U13874 (N_13874,N_12110,N_12524);
and U13875 (N_13875,N_12366,N_12388);
and U13876 (N_13876,N_12578,N_12938);
nor U13877 (N_13877,N_12240,N_12719);
nand U13878 (N_13878,N_12583,N_12250);
and U13879 (N_13879,N_12591,N_12672);
nand U13880 (N_13880,N_12380,N_12117);
or U13881 (N_13881,N_12332,N_12984);
nor U13882 (N_13882,N_12646,N_12082);
or U13883 (N_13883,N_12821,N_12477);
nor U13884 (N_13884,N_12571,N_12870);
xor U13885 (N_13885,N_12225,N_12667);
xor U13886 (N_13886,N_12432,N_12845);
or U13887 (N_13887,N_12761,N_12736);
nand U13888 (N_13888,N_12418,N_12066);
or U13889 (N_13889,N_12734,N_12815);
nor U13890 (N_13890,N_12094,N_12766);
xnor U13891 (N_13891,N_12163,N_12174);
and U13892 (N_13892,N_12488,N_12532);
or U13893 (N_13893,N_12809,N_12833);
xnor U13894 (N_13894,N_12914,N_12135);
or U13895 (N_13895,N_12192,N_12914);
xnor U13896 (N_13896,N_12277,N_12765);
or U13897 (N_13897,N_12830,N_12492);
or U13898 (N_13898,N_12580,N_12270);
and U13899 (N_13899,N_12160,N_12063);
xnor U13900 (N_13900,N_12763,N_12665);
xor U13901 (N_13901,N_12500,N_12538);
and U13902 (N_13902,N_12409,N_12082);
or U13903 (N_13903,N_12510,N_12382);
nand U13904 (N_13904,N_12635,N_12683);
and U13905 (N_13905,N_12895,N_12430);
xnor U13906 (N_13906,N_12199,N_12899);
or U13907 (N_13907,N_12353,N_12486);
xor U13908 (N_13908,N_12092,N_12329);
xor U13909 (N_13909,N_12829,N_12959);
nand U13910 (N_13910,N_12196,N_12828);
nand U13911 (N_13911,N_12801,N_12707);
and U13912 (N_13912,N_12737,N_12305);
and U13913 (N_13913,N_12574,N_12845);
nand U13914 (N_13914,N_12500,N_12023);
xnor U13915 (N_13915,N_12436,N_12017);
xor U13916 (N_13916,N_12330,N_12524);
nand U13917 (N_13917,N_12071,N_12008);
nand U13918 (N_13918,N_12846,N_12172);
or U13919 (N_13919,N_12973,N_12053);
xnor U13920 (N_13920,N_12755,N_12995);
nor U13921 (N_13921,N_12334,N_12539);
xor U13922 (N_13922,N_12388,N_12910);
nand U13923 (N_13923,N_12332,N_12085);
nand U13924 (N_13924,N_12904,N_12134);
nor U13925 (N_13925,N_12673,N_12814);
nand U13926 (N_13926,N_12315,N_12761);
nor U13927 (N_13927,N_12192,N_12705);
or U13928 (N_13928,N_12902,N_12005);
or U13929 (N_13929,N_12439,N_12891);
nor U13930 (N_13930,N_12355,N_12476);
nand U13931 (N_13931,N_12522,N_12924);
nand U13932 (N_13932,N_12386,N_12726);
or U13933 (N_13933,N_12566,N_12811);
and U13934 (N_13934,N_12962,N_12461);
and U13935 (N_13935,N_12721,N_12954);
and U13936 (N_13936,N_12735,N_12839);
and U13937 (N_13937,N_12599,N_12560);
and U13938 (N_13938,N_12888,N_12240);
nand U13939 (N_13939,N_12779,N_12542);
nor U13940 (N_13940,N_12697,N_12525);
nor U13941 (N_13941,N_12407,N_12140);
nand U13942 (N_13942,N_12406,N_12422);
or U13943 (N_13943,N_12553,N_12413);
nand U13944 (N_13944,N_12221,N_12301);
nand U13945 (N_13945,N_12446,N_12342);
or U13946 (N_13946,N_12871,N_12349);
or U13947 (N_13947,N_12639,N_12563);
nand U13948 (N_13948,N_12559,N_12270);
xnor U13949 (N_13949,N_12797,N_12890);
nor U13950 (N_13950,N_12741,N_12523);
nor U13951 (N_13951,N_12649,N_12500);
xor U13952 (N_13952,N_12726,N_12185);
xnor U13953 (N_13953,N_12976,N_12397);
nor U13954 (N_13954,N_12803,N_12382);
nand U13955 (N_13955,N_12590,N_12837);
nor U13956 (N_13956,N_12868,N_12233);
and U13957 (N_13957,N_12360,N_12365);
nor U13958 (N_13958,N_12423,N_12974);
or U13959 (N_13959,N_12508,N_12797);
nor U13960 (N_13960,N_12885,N_12777);
or U13961 (N_13961,N_12800,N_12955);
nor U13962 (N_13962,N_12132,N_12652);
nand U13963 (N_13963,N_12811,N_12745);
or U13964 (N_13964,N_12908,N_12019);
and U13965 (N_13965,N_12444,N_12993);
and U13966 (N_13966,N_12882,N_12118);
or U13967 (N_13967,N_12653,N_12199);
nor U13968 (N_13968,N_12868,N_12293);
or U13969 (N_13969,N_12419,N_12606);
nor U13970 (N_13970,N_12086,N_12285);
xnor U13971 (N_13971,N_12643,N_12271);
nor U13972 (N_13972,N_12253,N_12472);
or U13973 (N_13973,N_12784,N_12542);
or U13974 (N_13974,N_12687,N_12651);
nand U13975 (N_13975,N_12883,N_12804);
or U13976 (N_13976,N_12551,N_12080);
xnor U13977 (N_13977,N_12292,N_12382);
nor U13978 (N_13978,N_12896,N_12201);
nand U13979 (N_13979,N_12873,N_12339);
xnor U13980 (N_13980,N_12779,N_12849);
and U13981 (N_13981,N_12715,N_12434);
and U13982 (N_13982,N_12581,N_12355);
nand U13983 (N_13983,N_12249,N_12147);
nand U13984 (N_13984,N_12471,N_12187);
nor U13985 (N_13985,N_12859,N_12581);
nor U13986 (N_13986,N_12776,N_12825);
nor U13987 (N_13987,N_12018,N_12016);
nor U13988 (N_13988,N_12032,N_12201);
or U13989 (N_13989,N_12246,N_12823);
xor U13990 (N_13990,N_12458,N_12875);
nor U13991 (N_13991,N_12615,N_12880);
nor U13992 (N_13992,N_12832,N_12371);
nor U13993 (N_13993,N_12445,N_12394);
xor U13994 (N_13994,N_12837,N_12447);
xnor U13995 (N_13995,N_12521,N_12500);
nor U13996 (N_13996,N_12609,N_12369);
or U13997 (N_13997,N_12284,N_12359);
and U13998 (N_13998,N_12983,N_12568);
and U13999 (N_13999,N_12156,N_12921);
nand U14000 (N_14000,N_13548,N_13821);
or U14001 (N_14001,N_13423,N_13169);
xor U14002 (N_14002,N_13659,N_13135);
nor U14003 (N_14003,N_13830,N_13287);
nor U14004 (N_14004,N_13337,N_13476);
and U14005 (N_14005,N_13353,N_13240);
nor U14006 (N_14006,N_13433,N_13801);
nand U14007 (N_14007,N_13612,N_13194);
xnor U14008 (N_14008,N_13113,N_13211);
or U14009 (N_14009,N_13691,N_13846);
nor U14010 (N_14010,N_13312,N_13876);
or U14011 (N_14011,N_13982,N_13740);
nand U14012 (N_14012,N_13653,N_13416);
nand U14013 (N_14013,N_13391,N_13276);
xnor U14014 (N_14014,N_13804,N_13989);
nand U14015 (N_14015,N_13731,N_13803);
and U14016 (N_14016,N_13481,N_13511);
nand U14017 (N_14017,N_13586,N_13522);
nor U14018 (N_14018,N_13361,N_13131);
and U14019 (N_14019,N_13026,N_13692);
or U14020 (N_14020,N_13616,N_13623);
nand U14021 (N_14021,N_13806,N_13634);
nand U14022 (N_14022,N_13293,N_13921);
nor U14023 (N_14023,N_13122,N_13350);
nand U14024 (N_14024,N_13894,N_13392);
xor U14025 (N_14025,N_13782,N_13385);
xnor U14026 (N_14026,N_13075,N_13333);
nor U14027 (N_14027,N_13095,N_13638);
or U14028 (N_14028,N_13329,N_13282);
nand U14029 (N_14029,N_13307,N_13195);
or U14030 (N_14030,N_13327,N_13648);
and U14031 (N_14031,N_13847,N_13184);
xnor U14032 (N_14032,N_13726,N_13457);
xor U14033 (N_14033,N_13364,N_13158);
nand U14034 (N_14034,N_13837,N_13802);
and U14035 (N_14035,N_13465,N_13508);
and U14036 (N_14036,N_13605,N_13566);
and U14037 (N_14037,N_13761,N_13315);
xnor U14038 (N_14038,N_13763,N_13179);
nor U14039 (N_14039,N_13979,N_13028);
or U14040 (N_14040,N_13303,N_13469);
or U14041 (N_14041,N_13020,N_13283);
and U14042 (N_14042,N_13112,N_13973);
and U14043 (N_14043,N_13063,N_13816);
nor U14044 (N_14044,N_13372,N_13064);
or U14045 (N_14045,N_13954,N_13785);
and U14046 (N_14046,N_13765,N_13927);
and U14047 (N_14047,N_13222,N_13013);
and U14048 (N_14048,N_13844,N_13811);
and U14049 (N_14049,N_13067,N_13794);
nand U14050 (N_14050,N_13498,N_13658);
nor U14051 (N_14051,N_13243,N_13996);
nand U14052 (N_14052,N_13902,N_13983);
or U14053 (N_14053,N_13219,N_13775);
and U14054 (N_14054,N_13091,N_13199);
xnor U14055 (N_14055,N_13736,N_13300);
nand U14056 (N_14056,N_13474,N_13723);
xnor U14057 (N_14057,N_13912,N_13880);
or U14058 (N_14058,N_13126,N_13396);
and U14059 (N_14059,N_13602,N_13881);
and U14060 (N_14060,N_13629,N_13621);
nand U14061 (N_14061,N_13237,N_13681);
or U14062 (N_14062,N_13482,N_13796);
nor U14063 (N_14063,N_13210,N_13836);
xnor U14064 (N_14064,N_13878,N_13571);
xnor U14065 (N_14065,N_13226,N_13551);
and U14066 (N_14066,N_13850,N_13684);
and U14067 (N_14067,N_13727,N_13228);
xnor U14068 (N_14068,N_13932,N_13149);
xnor U14069 (N_14069,N_13784,N_13077);
xor U14070 (N_14070,N_13948,N_13008);
nor U14071 (N_14071,N_13885,N_13102);
or U14072 (N_14072,N_13165,N_13001);
and U14073 (N_14073,N_13834,N_13640);
and U14074 (N_14074,N_13872,N_13710);
and U14075 (N_14075,N_13084,N_13233);
xnor U14076 (N_14076,N_13456,N_13892);
nor U14077 (N_14077,N_13600,N_13576);
nor U14078 (N_14078,N_13851,N_13060);
and U14079 (N_14079,N_13815,N_13764);
nor U14080 (N_14080,N_13752,N_13206);
xor U14081 (N_14081,N_13715,N_13514);
or U14082 (N_14082,N_13120,N_13048);
or U14083 (N_14083,N_13073,N_13485);
xnor U14084 (N_14084,N_13769,N_13045);
xor U14085 (N_14085,N_13907,N_13117);
and U14086 (N_14086,N_13827,N_13929);
or U14087 (N_14087,N_13947,N_13682);
and U14088 (N_14088,N_13147,N_13177);
nor U14089 (N_14089,N_13032,N_13491);
nand U14090 (N_14090,N_13411,N_13635);
xor U14091 (N_14091,N_13035,N_13777);
nand U14092 (N_14092,N_13232,N_13589);
xor U14093 (N_14093,N_13384,N_13415);
nand U14094 (N_14094,N_13029,N_13565);
nor U14095 (N_14095,N_13760,N_13478);
nor U14096 (N_14096,N_13351,N_13175);
nand U14097 (N_14097,N_13757,N_13579);
nand U14098 (N_14098,N_13578,N_13173);
xnor U14099 (N_14099,N_13537,N_13201);
or U14100 (N_14100,N_13399,N_13408);
and U14101 (N_14101,N_13146,N_13431);
or U14102 (N_14102,N_13231,N_13174);
nor U14103 (N_14103,N_13119,N_13156);
or U14104 (N_14104,N_13883,N_13202);
xnor U14105 (N_14105,N_13945,N_13022);
nor U14106 (N_14106,N_13607,N_13272);
and U14107 (N_14107,N_13034,N_13845);
nand U14108 (N_14108,N_13182,N_13019);
xnor U14109 (N_14109,N_13627,N_13573);
and U14110 (N_14110,N_13288,N_13963);
xnor U14111 (N_14111,N_13314,N_13234);
or U14112 (N_14112,N_13459,N_13289);
and U14113 (N_14113,N_13848,N_13434);
nand U14114 (N_14114,N_13745,N_13855);
nand U14115 (N_14115,N_13114,N_13323);
and U14116 (N_14116,N_13393,N_13426);
and U14117 (N_14117,N_13338,N_13654);
nand U14118 (N_14118,N_13718,N_13357);
and U14119 (N_14119,N_13525,N_13488);
and U14120 (N_14120,N_13517,N_13859);
xnor U14121 (N_14121,N_13613,N_13557);
nand U14122 (N_14122,N_13800,N_13441);
and U14123 (N_14123,N_13500,N_13563);
and U14124 (N_14124,N_13261,N_13269);
nand U14125 (N_14125,N_13931,N_13667);
nor U14126 (N_14126,N_13220,N_13241);
xor U14127 (N_14127,N_13383,N_13780);
or U14128 (N_14128,N_13196,N_13247);
nand U14129 (N_14129,N_13879,N_13510);
or U14130 (N_14130,N_13424,N_13754);
or U14131 (N_14131,N_13601,N_13055);
nand U14132 (N_14132,N_13734,N_13406);
xnor U14133 (N_14133,N_13208,N_13593);
and U14134 (N_14134,N_13239,N_13388);
and U14135 (N_14135,N_13330,N_13334);
and U14136 (N_14136,N_13292,N_13581);
nor U14137 (N_14137,N_13504,N_13301);
and U14138 (N_14138,N_13935,N_13884);
nor U14139 (N_14139,N_13628,N_13153);
nand U14140 (N_14140,N_13286,N_13753);
nor U14141 (N_14141,N_13118,N_13311);
nor U14142 (N_14142,N_13087,N_13322);
and U14143 (N_14143,N_13524,N_13365);
nand U14144 (N_14144,N_13000,N_13052);
xor U14145 (N_14145,N_13766,N_13253);
and U14146 (N_14146,N_13660,N_13093);
nor U14147 (N_14147,N_13904,N_13747);
nand U14148 (N_14148,N_13866,N_13911);
and U14149 (N_14149,N_13622,N_13987);
nand U14150 (N_14150,N_13890,N_13442);
xnor U14151 (N_14151,N_13405,N_13922);
and U14152 (N_14152,N_13939,N_13676);
xnor U14153 (N_14153,N_13422,N_13893);
or U14154 (N_14154,N_13507,N_13549);
xnor U14155 (N_14155,N_13097,N_13750);
nand U14156 (N_14156,N_13428,N_13965);
and U14157 (N_14157,N_13429,N_13273);
nand U14158 (N_14158,N_13995,N_13502);
nor U14159 (N_14159,N_13271,N_13448);
and U14160 (N_14160,N_13799,N_13709);
and U14161 (N_14161,N_13244,N_13661);
nor U14162 (N_14162,N_13284,N_13224);
and U14163 (N_14163,N_13460,N_13853);
and U14164 (N_14164,N_13187,N_13523);
nand U14165 (N_14165,N_13266,N_13212);
nor U14166 (N_14166,N_13778,N_13076);
nand U14167 (N_14167,N_13221,N_13347);
nand U14168 (N_14168,N_13795,N_13235);
or U14169 (N_14169,N_13908,N_13438);
nor U14170 (N_14170,N_13376,N_13695);
nand U14171 (N_14171,N_13157,N_13547);
nor U14172 (N_14172,N_13310,N_13620);
nor U14173 (N_14173,N_13352,N_13011);
and U14174 (N_14174,N_13756,N_13567);
xor U14175 (N_14175,N_13545,N_13340);
and U14176 (N_14176,N_13839,N_13767);
nor U14177 (N_14177,N_13749,N_13991);
and U14178 (N_14178,N_13479,N_13952);
or U14179 (N_14179,N_13400,N_13722);
nand U14180 (N_14180,N_13900,N_13069);
nor U14181 (N_14181,N_13694,N_13185);
or U14182 (N_14182,N_13964,N_13192);
xor U14183 (N_14183,N_13650,N_13527);
and U14184 (N_14184,N_13216,N_13043);
nor U14185 (N_14185,N_13572,N_13395);
xnor U14186 (N_14186,N_13025,N_13103);
xnor U14187 (N_14187,N_13402,N_13444);
nand U14188 (N_14188,N_13713,N_13798);
xor U14189 (N_14189,N_13919,N_13701);
nand U14190 (N_14190,N_13379,N_13615);
or U14191 (N_14191,N_13840,N_13430);
nand U14192 (N_14192,N_13298,N_13018);
nor U14193 (N_14193,N_13611,N_13374);
nor U14194 (N_14194,N_13373,N_13637);
nor U14195 (N_14195,N_13492,N_13814);
nor U14196 (N_14196,N_13462,N_13590);
and U14197 (N_14197,N_13100,N_13976);
and U14198 (N_14198,N_13506,N_13528);
nor U14199 (N_14199,N_13992,N_13010);
nor U14200 (N_14200,N_13267,N_13789);
nor U14201 (N_14201,N_13852,N_13369);
nand U14202 (N_14202,N_13386,N_13550);
xor U14203 (N_14203,N_13015,N_13421);
or U14204 (N_14204,N_13874,N_13223);
and U14205 (N_14205,N_13132,N_13154);
nand U14206 (N_14206,N_13541,N_13082);
xor U14207 (N_14207,N_13030,N_13464);
and U14208 (N_14208,N_13309,N_13978);
nand U14209 (N_14209,N_13320,N_13822);
or U14210 (N_14210,N_13348,N_13959);
nor U14211 (N_14211,N_13072,N_13435);
nor U14212 (N_14212,N_13042,N_13554);
and U14213 (N_14213,N_13703,N_13940);
and U14214 (N_14214,N_13407,N_13728);
xnor U14215 (N_14215,N_13362,N_13066);
and U14216 (N_14216,N_13170,N_13378);
nand U14217 (N_14217,N_13652,N_13920);
nand U14218 (N_14218,N_13059,N_13553);
nor U14219 (N_14219,N_13249,N_13213);
xor U14220 (N_14220,N_13630,N_13138);
nand U14221 (N_14221,N_13040,N_13257);
nor U14222 (N_14222,N_13439,N_13229);
nand U14223 (N_14223,N_13260,N_13746);
and U14224 (N_14224,N_13918,N_13655);
nor U14225 (N_14225,N_13044,N_13748);
nor U14226 (N_14226,N_13535,N_13265);
and U14227 (N_14227,N_13227,N_13955);
or U14228 (N_14228,N_13242,N_13090);
xor U14229 (N_14229,N_13606,N_13735);
and U14230 (N_14230,N_13555,N_13826);
nand U14231 (N_14231,N_13246,N_13024);
xor U14232 (N_14232,N_13644,N_13259);
nand U14233 (N_14233,N_13302,N_13036);
nand U14234 (N_14234,N_13843,N_13033);
and U14235 (N_14235,N_13452,N_13558);
or U14236 (N_14236,N_13057,N_13588);
and U14237 (N_14237,N_13544,N_13009);
and U14238 (N_14238,N_13109,N_13639);
nand U14239 (N_14239,N_13985,N_13533);
and U14240 (N_14240,N_13693,N_13285);
nand U14241 (N_14241,N_13598,N_13556);
nand U14242 (N_14242,N_13121,N_13704);
or U14243 (N_14243,N_13536,N_13451);
xnor U14244 (N_14244,N_13074,N_13349);
and U14245 (N_14245,N_13290,N_13123);
nand U14246 (N_14246,N_13688,N_13531);
nor U14247 (N_14247,N_13862,N_13092);
nand U14248 (N_14248,N_13546,N_13262);
xnor U14249 (N_14249,N_13994,N_13129);
and U14250 (N_14250,N_13200,N_13432);
xnor U14251 (N_14251,N_13171,N_13291);
or U14252 (N_14252,N_13145,N_13743);
xor U14253 (N_14253,N_13662,N_13418);
and U14254 (N_14254,N_13998,N_13007);
or U14255 (N_14255,N_13294,N_13868);
xor U14256 (N_14256,N_13410,N_13732);
xnor U14257 (N_14257,N_13958,N_13197);
xor U14258 (N_14258,N_13759,N_13779);
or U14259 (N_14259,N_13136,N_13670);
xnor U14260 (N_14260,N_13336,N_13509);
and U14261 (N_14261,N_13079,N_13455);
xor U14262 (N_14262,N_13651,N_13552);
nor U14263 (N_14263,N_13513,N_13377);
and U14264 (N_14264,N_13833,N_13130);
xor U14265 (N_14265,N_13966,N_13813);
xor U14266 (N_14266,N_13215,N_13248);
nor U14267 (N_14267,N_13081,N_13990);
xor U14268 (N_14268,N_13915,N_13207);
nand U14269 (N_14269,N_13398,N_13768);
and U14270 (N_14270,N_13111,N_13168);
and U14271 (N_14271,N_13217,N_13596);
nand U14272 (N_14272,N_13316,N_13863);
or U14273 (N_14273,N_13870,N_13755);
or U14274 (N_14274,N_13762,N_13645);
nor U14275 (N_14275,N_13610,N_13751);
nor U14276 (N_14276,N_13071,N_13970);
or U14277 (N_14277,N_13618,N_13281);
nor U14278 (N_14278,N_13949,N_13706);
xor U14279 (N_14279,N_13115,N_13162);
or U14280 (N_14280,N_13062,N_13370);
and U14281 (N_14281,N_13274,N_13313);
or U14282 (N_14282,N_13716,N_13397);
xnor U14283 (N_14283,N_13561,N_13086);
nor U14284 (N_14284,N_13923,N_13188);
nand U14285 (N_14285,N_13236,N_13986);
nor U14286 (N_14286,N_13065,N_13520);
nor U14287 (N_14287,N_13897,N_13980);
nor U14288 (N_14288,N_13413,N_13205);
and U14289 (N_14289,N_13142,N_13968);
and U14290 (N_14290,N_13591,N_13582);
and U14291 (N_14291,N_13898,N_13595);
xnor U14292 (N_14292,N_13542,N_13512);
xnor U14293 (N_14293,N_13790,N_13070);
or U14294 (N_14294,N_13449,N_13487);
nor U14295 (N_14295,N_13166,N_13463);
and U14296 (N_14296,N_13818,N_13258);
or U14297 (N_14297,N_13608,N_13574);
or U14298 (N_14298,N_13854,N_13308);
or U14299 (N_14299,N_13360,N_13559);
nand U14300 (N_14300,N_13331,N_13698);
or U14301 (N_14301,N_13819,N_13675);
or U14302 (N_14302,N_13039,N_13975);
xnor U14303 (N_14303,N_13403,N_13251);
nor U14304 (N_14304,N_13832,N_13930);
nand U14305 (N_14305,N_13678,N_13673);
nor U14306 (N_14306,N_13471,N_13677);
or U14307 (N_14307,N_13592,N_13705);
xnor U14308 (N_14308,N_13381,N_13758);
nand U14309 (N_14309,N_13160,N_13599);
nor U14310 (N_14310,N_13860,N_13354);
nand U14311 (N_14311,N_13027,N_13058);
nand U14312 (N_14312,N_13943,N_13218);
or U14313 (N_14313,N_13882,N_13647);
or U14314 (N_14314,N_13917,N_13903);
xnor U14315 (N_14315,N_13107,N_13324);
and U14316 (N_14316,N_13961,N_13341);
nand U14317 (N_14317,N_13106,N_13937);
or U14318 (N_14318,N_13280,N_13409);
and U14319 (N_14319,N_13203,N_13906);
nor U14320 (N_14320,N_13910,N_13049);
and U14321 (N_14321,N_13928,N_13702);
nor U14322 (N_14322,N_13642,N_13152);
nand U14323 (N_14323,N_13105,N_13375);
xor U14324 (N_14324,N_13717,N_13962);
xor U14325 (N_14325,N_13950,N_13969);
and U14326 (N_14326,N_13913,N_13946);
nor U14327 (N_14327,N_13101,N_13663);
or U14328 (N_14328,N_13742,N_13299);
nor U14329 (N_14329,N_13787,N_13916);
nor U14330 (N_14330,N_13808,N_13161);
nand U14331 (N_14331,N_13807,N_13128);
xnor U14332 (N_14332,N_13467,N_13458);
or U14333 (N_14333,N_13080,N_13888);
or U14334 (N_14334,N_13971,N_13696);
xor U14335 (N_14335,N_13538,N_13425);
xor U14336 (N_14336,N_13490,N_13841);
nand U14337 (N_14337,N_13047,N_13321);
and U14338 (N_14338,N_13172,N_13875);
or U14339 (N_14339,N_13669,N_13214);
or U14340 (N_14340,N_13690,N_13636);
nand U14341 (N_14341,N_13560,N_13575);
and U14342 (N_14342,N_13012,N_13021);
or U14343 (N_14343,N_13417,N_13346);
xnor U14344 (N_14344,N_13339,N_13526);
or U14345 (N_14345,N_13603,N_13108);
nor U14346 (N_14346,N_13404,N_13252);
xnor U14347 (N_14347,N_13484,N_13190);
or U14348 (N_14348,N_13116,N_13094);
xnor U14349 (N_14349,N_13163,N_13486);
or U14350 (N_14350,N_13981,N_13499);
nor U14351 (N_14351,N_13141,N_13016);
xor U14352 (N_14352,N_13318,N_13817);
or U14353 (N_14353,N_13583,N_13797);
xnor U14354 (N_14354,N_13665,N_13617);
and U14355 (N_14355,N_13711,N_13225);
or U14356 (N_14356,N_13858,N_13356);
nand U14357 (N_14357,N_13686,N_13264);
nand U14358 (N_14358,N_13230,N_13689);
nor U14359 (N_14359,N_13577,N_13137);
xor U14360 (N_14360,N_13865,N_13401);
xor U14361 (N_14361,N_13304,N_13914);
and U14362 (N_14362,N_13366,N_13532);
and U14363 (N_14363,N_13104,N_13873);
or U14364 (N_14364,N_13041,N_13295);
and U14365 (N_14365,N_13905,N_13887);
or U14366 (N_14366,N_13176,N_13445);
nand U14367 (N_14367,N_13580,N_13326);
nor U14368 (N_14368,N_13632,N_13984);
or U14369 (N_14369,N_13614,N_13254);
nand U14370 (N_14370,N_13842,N_13772);
and U14371 (N_14371,N_13359,N_13186);
or U14372 (N_14372,N_13503,N_13389);
nand U14373 (N_14373,N_13098,N_13150);
nor U14374 (N_14374,N_13719,N_13960);
and U14375 (N_14375,N_13125,N_13899);
and U14376 (N_14376,N_13771,N_13999);
or U14377 (N_14377,N_13367,N_13006);
xnor U14378 (N_14378,N_13744,N_13355);
nand U14379 (N_14379,N_13901,N_13468);
nor U14380 (N_14380,N_13148,N_13414);
nand U14381 (N_14381,N_13387,N_13530);
nor U14382 (N_14382,N_13515,N_13671);
nor U14383 (N_14383,N_13518,N_13909);
nand U14384 (N_14384,N_13721,N_13562);
and U14385 (N_14385,N_13869,N_13683);
xor U14386 (N_14386,N_13088,N_13933);
nand U14387 (N_14387,N_13427,N_13604);
nor U14388 (N_14388,N_13877,N_13972);
xor U14389 (N_14389,N_13685,N_13788);
nand U14390 (N_14390,N_13720,N_13134);
and U14391 (N_14391,N_13809,N_13521);
or U14392 (N_14392,N_13997,N_13594);
nand U14393 (N_14393,N_13891,N_13089);
nand U14394 (N_14394,N_13133,N_13825);
nor U14395 (N_14395,N_13781,N_13495);
nand U14396 (N_14396,N_13159,N_13317);
or U14397 (N_14397,N_13124,N_13003);
or U14398 (N_14398,N_13540,N_13569);
nor U14399 (N_14399,N_13679,N_13489);
nor U14400 (N_14400,N_13505,N_13956);
nand U14401 (N_14401,N_13680,N_13256);
and U14402 (N_14402,N_13023,N_13483);
or U14403 (N_14403,N_13708,N_13649);
nor U14404 (N_14404,N_13061,N_13741);
xor U14405 (N_14405,N_13443,N_13516);
or U14406 (N_14406,N_13934,N_13178);
nand U14407 (N_14407,N_13856,N_13493);
nand U14408 (N_14408,N_13279,N_13419);
nand U14409 (N_14409,N_13829,N_13774);
nand U14410 (N_14410,N_13861,N_13151);
nor U14411 (N_14411,N_13164,N_13739);
or U14412 (N_14412,N_13371,N_13953);
nor U14413 (N_14413,N_13770,N_13564);
nand U14414 (N_14414,N_13420,N_13519);
or U14415 (N_14415,N_13344,N_13193);
nand U14416 (N_14416,N_13730,N_13453);
nand U14417 (N_14417,N_13472,N_13597);
nand U14418 (N_14418,N_13306,N_13944);
xor U14419 (N_14419,N_13738,N_13167);
and U14420 (N_14420,N_13776,N_13926);
nand U14421 (N_14421,N_13886,N_13864);
and U14422 (N_14422,N_13773,N_13181);
nor U14423 (N_14423,N_13823,N_13051);
nor U14424 (N_14424,N_13277,N_13390);
xnor U14425 (N_14425,N_13031,N_13440);
or U14426 (N_14426,N_13450,N_13002);
nand U14427 (N_14427,N_13786,N_13496);
nand U14428 (N_14428,N_13646,N_13724);
xor U14429 (N_14429,N_13977,N_13038);
nand U14430 (N_14430,N_13143,N_13951);
nor U14431 (N_14431,N_13127,N_13305);
or U14432 (N_14432,N_13480,N_13729);
xnor U14433 (N_14433,N_13672,N_13810);
and U14434 (N_14434,N_13828,N_13657);
xor U14435 (N_14435,N_13447,N_13204);
nor U14436 (N_14436,N_13099,N_13957);
and U14437 (N_14437,N_13096,N_13633);
and U14438 (N_14438,N_13941,N_13570);
nor U14439 (N_14439,N_13068,N_13466);
and U14440 (N_14440,N_13144,N_13626);
nor U14441 (N_14441,N_13725,N_13005);
nor U14442 (N_14442,N_13473,N_13587);
nor U14443 (N_14443,N_13278,N_13446);
xnor U14444 (N_14444,N_13270,N_13643);
nand U14445 (N_14445,N_13475,N_13189);
nand U14446 (N_14446,N_13477,N_13568);
and U14447 (N_14447,N_13412,N_13664);
xnor U14448 (N_14448,N_13319,N_13831);
nor U14449 (N_14449,N_13342,N_13820);
and U14450 (N_14450,N_13394,N_13053);
or U14451 (N_14451,N_13534,N_13687);
or U14452 (N_14452,N_13363,N_13641);
or U14453 (N_14453,N_13824,N_13792);
and U14454 (N_14454,N_13180,N_13942);
and U14455 (N_14455,N_13714,N_13245);
xor U14456 (N_14456,N_13014,N_13297);
nand U14457 (N_14457,N_13494,N_13791);
nor U14458 (N_14458,N_13268,N_13631);
or U14459 (N_14459,N_13335,N_13078);
or U14460 (N_14460,N_13083,N_13110);
nor U14461 (N_14461,N_13343,N_13993);
nand U14462 (N_14462,N_13275,N_13017);
xnor U14463 (N_14463,N_13624,N_13889);
nand U14464 (N_14464,N_13436,N_13835);
nand U14465 (N_14465,N_13805,N_13332);
nor U14466 (N_14466,N_13967,N_13250);
and U14467 (N_14467,N_13296,N_13707);
and U14468 (N_14468,N_13461,N_13263);
xnor U14469 (N_14469,N_13470,N_13974);
nor U14470 (N_14470,N_13382,N_13699);
xor U14471 (N_14471,N_13238,N_13697);
nor U14472 (N_14472,N_13619,N_13857);
nand U14473 (N_14473,N_13004,N_13871);
and U14474 (N_14474,N_13925,N_13345);
nand U14475 (N_14475,N_13838,N_13895);
nand U14476 (N_14476,N_13255,N_13529);
xor U14477 (N_14477,N_13501,N_13584);
and U14478 (N_14478,N_13358,N_13368);
xnor U14479 (N_14479,N_13812,N_13056);
or U14480 (N_14480,N_13037,N_13938);
and U14481 (N_14481,N_13497,N_13209);
or U14482 (N_14482,N_13539,N_13793);
and U14483 (N_14483,N_13712,N_13737);
nor U14484 (N_14484,N_13988,N_13139);
nor U14485 (N_14485,N_13140,N_13183);
xor U14486 (N_14486,N_13454,N_13050);
and U14487 (N_14487,N_13849,N_13625);
or U14488 (N_14488,N_13198,N_13674);
nor U14489 (N_14489,N_13085,N_13543);
nor U14490 (N_14490,N_13609,N_13328);
nor U14491 (N_14491,N_13325,N_13046);
and U14492 (N_14492,N_13054,N_13585);
nor U14493 (N_14493,N_13924,N_13191);
or U14494 (N_14494,N_13936,N_13656);
nand U14495 (N_14495,N_13700,N_13896);
nand U14496 (N_14496,N_13155,N_13666);
xor U14497 (N_14497,N_13867,N_13783);
or U14498 (N_14498,N_13380,N_13668);
nor U14499 (N_14499,N_13733,N_13437);
xor U14500 (N_14500,N_13404,N_13443);
xor U14501 (N_14501,N_13129,N_13639);
and U14502 (N_14502,N_13669,N_13386);
or U14503 (N_14503,N_13586,N_13124);
and U14504 (N_14504,N_13628,N_13800);
nand U14505 (N_14505,N_13215,N_13330);
or U14506 (N_14506,N_13458,N_13212);
nor U14507 (N_14507,N_13733,N_13051);
and U14508 (N_14508,N_13797,N_13859);
and U14509 (N_14509,N_13931,N_13182);
nor U14510 (N_14510,N_13333,N_13355);
xor U14511 (N_14511,N_13463,N_13372);
nand U14512 (N_14512,N_13042,N_13736);
or U14513 (N_14513,N_13424,N_13444);
nand U14514 (N_14514,N_13999,N_13895);
nor U14515 (N_14515,N_13963,N_13408);
and U14516 (N_14516,N_13880,N_13341);
nor U14517 (N_14517,N_13342,N_13078);
or U14518 (N_14518,N_13799,N_13801);
xor U14519 (N_14519,N_13306,N_13801);
and U14520 (N_14520,N_13874,N_13175);
xnor U14521 (N_14521,N_13586,N_13335);
nand U14522 (N_14522,N_13823,N_13154);
and U14523 (N_14523,N_13672,N_13917);
xnor U14524 (N_14524,N_13028,N_13644);
xnor U14525 (N_14525,N_13314,N_13197);
xor U14526 (N_14526,N_13309,N_13914);
nand U14527 (N_14527,N_13600,N_13569);
xor U14528 (N_14528,N_13783,N_13762);
and U14529 (N_14529,N_13585,N_13395);
and U14530 (N_14530,N_13427,N_13495);
nor U14531 (N_14531,N_13606,N_13094);
xor U14532 (N_14532,N_13010,N_13168);
xnor U14533 (N_14533,N_13616,N_13892);
nor U14534 (N_14534,N_13395,N_13180);
nor U14535 (N_14535,N_13424,N_13021);
nand U14536 (N_14536,N_13210,N_13594);
or U14537 (N_14537,N_13141,N_13594);
nand U14538 (N_14538,N_13542,N_13560);
or U14539 (N_14539,N_13907,N_13966);
xor U14540 (N_14540,N_13641,N_13670);
xnor U14541 (N_14541,N_13983,N_13424);
nand U14542 (N_14542,N_13045,N_13019);
and U14543 (N_14543,N_13859,N_13553);
or U14544 (N_14544,N_13289,N_13747);
or U14545 (N_14545,N_13551,N_13264);
nand U14546 (N_14546,N_13126,N_13888);
nor U14547 (N_14547,N_13815,N_13246);
xnor U14548 (N_14548,N_13555,N_13101);
and U14549 (N_14549,N_13038,N_13866);
and U14550 (N_14550,N_13264,N_13986);
or U14551 (N_14551,N_13252,N_13155);
xnor U14552 (N_14552,N_13949,N_13281);
and U14553 (N_14553,N_13049,N_13323);
nor U14554 (N_14554,N_13274,N_13736);
or U14555 (N_14555,N_13611,N_13688);
and U14556 (N_14556,N_13526,N_13432);
or U14557 (N_14557,N_13785,N_13454);
xor U14558 (N_14558,N_13531,N_13446);
nor U14559 (N_14559,N_13582,N_13611);
xor U14560 (N_14560,N_13323,N_13989);
nand U14561 (N_14561,N_13656,N_13897);
xnor U14562 (N_14562,N_13176,N_13753);
xor U14563 (N_14563,N_13652,N_13714);
nor U14564 (N_14564,N_13806,N_13195);
and U14565 (N_14565,N_13591,N_13546);
and U14566 (N_14566,N_13185,N_13823);
nand U14567 (N_14567,N_13079,N_13558);
xor U14568 (N_14568,N_13322,N_13101);
xnor U14569 (N_14569,N_13166,N_13836);
nand U14570 (N_14570,N_13004,N_13249);
nand U14571 (N_14571,N_13517,N_13298);
nand U14572 (N_14572,N_13923,N_13572);
xor U14573 (N_14573,N_13936,N_13336);
or U14574 (N_14574,N_13258,N_13661);
and U14575 (N_14575,N_13268,N_13244);
nand U14576 (N_14576,N_13195,N_13965);
nand U14577 (N_14577,N_13283,N_13420);
or U14578 (N_14578,N_13815,N_13515);
xnor U14579 (N_14579,N_13197,N_13528);
and U14580 (N_14580,N_13769,N_13801);
and U14581 (N_14581,N_13784,N_13301);
or U14582 (N_14582,N_13414,N_13837);
or U14583 (N_14583,N_13669,N_13539);
nor U14584 (N_14584,N_13661,N_13755);
and U14585 (N_14585,N_13274,N_13283);
xor U14586 (N_14586,N_13133,N_13924);
or U14587 (N_14587,N_13206,N_13553);
nand U14588 (N_14588,N_13019,N_13601);
and U14589 (N_14589,N_13505,N_13201);
and U14590 (N_14590,N_13300,N_13243);
xnor U14591 (N_14591,N_13020,N_13917);
nor U14592 (N_14592,N_13150,N_13073);
nor U14593 (N_14593,N_13315,N_13568);
or U14594 (N_14594,N_13877,N_13093);
nand U14595 (N_14595,N_13403,N_13312);
xor U14596 (N_14596,N_13691,N_13913);
and U14597 (N_14597,N_13008,N_13238);
or U14598 (N_14598,N_13598,N_13267);
nand U14599 (N_14599,N_13444,N_13592);
nor U14600 (N_14600,N_13642,N_13680);
xnor U14601 (N_14601,N_13982,N_13107);
nor U14602 (N_14602,N_13318,N_13540);
and U14603 (N_14603,N_13652,N_13322);
xnor U14604 (N_14604,N_13042,N_13561);
or U14605 (N_14605,N_13648,N_13848);
nor U14606 (N_14606,N_13452,N_13621);
or U14607 (N_14607,N_13565,N_13818);
nor U14608 (N_14608,N_13421,N_13453);
xnor U14609 (N_14609,N_13445,N_13374);
or U14610 (N_14610,N_13075,N_13162);
or U14611 (N_14611,N_13659,N_13905);
xor U14612 (N_14612,N_13798,N_13667);
xnor U14613 (N_14613,N_13744,N_13050);
nand U14614 (N_14614,N_13906,N_13543);
nor U14615 (N_14615,N_13608,N_13946);
xnor U14616 (N_14616,N_13145,N_13151);
or U14617 (N_14617,N_13750,N_13893);
nand U14618 (N_14618,N_13215,N_13746);
or U14619 (N_14619,N_13495,N_13893);
or U14620 (N_14620,N_13075,N_13638);
xor U14621 (N_14621,N_13838,N_13392);
or U14622 (N_14622,N_13014,N_13738);
and U14623 (N_14623,N_13686,N_13975);
xnor U14624 (N_14624,N_13801,N_13804);
or U14625 (N_14625,N_13833,N_13895);
nor U14626 (N_14626,N_13069,N_13912);
xnor U14627 (N_14627,N_13125,N_13638);
nor U14628 (N_14628,N_13475,N_13461);
xnor U14629 (N_14629,N_13991,N_13806);
nand U14630 (N_14630,N_13686,N_13226);
or U14631 (N_14631,N_13265,N_13629);
nor U14632 (N_14632,N_13433,N_13303);
or U14633 (N_14633,N_13697,N_13675);
nor U14634 (N_14634,N_13599,N_13832);
and U14635 (N_14635,N_13658,N_13292);
nor U14636 (N_14636,N_13874,N_13901);
xnor U14637 (N_14637,N_13458,N_13546);
or U14638 (N_14638,N_13499,N_13378);
or U14639 (N_14639,N_13011,N_13177);
nand U14640 (N_14640,N_13252,N_13842);
nand U14641 (N_14641,N_13230,N_13059);
or U14642 (N_14642,N_13610,N_13028);
nor U14643 (N_14643,N_13323,N_13454);
nand U14644 (N_14644,N_13090,N_13948);
nand U14645 (N_14645,N_13061,N_13802);
xnor U14646 (N_14646,N_13398,N_13525);
nor U14647 (N_14647,N_13111,N_13183);
xor U14648 (N_14648,N_13969,N_13170);
and U14649 (N_14649,N_13419,N_13249);
nor U14650 (N_14650,N_13989,N_13108);
or U14651 (N_14651,N_13266,N_13619);
xnor U14652 (N_14652,N_13158,N_13408);
nand U14653 (N_14653,N_13975,N_13995);
and U14654 (N_14654,N_13825,N_13417);
nor U14655 (N_14655,N_13942,N_13890);
xor U14656 (N_14656,N_13919,N_13901);
nor U14657 (N_14657,N_13407,N_13113);
nand U14658 (N_14658,N_13182,N_13156);
xnor U14659 (N_14659,N_13625,N_13699);
and U14660 (N_14660,N_13928,N_13617);
and U14661 (N_14661,N_13194,N_13825);
nand U14662 (N_14662,N_13750,N_13785);
and U14663 (N_14663,N_13451,N_13613);
nor U14664 (N_14664,N_13527,N_13311);
and U14665 (N_14665,N_13614,N_13065);
or U14666 (N_14666,N_13718,N_13523);
and U14667 (N_14667,N_13293,N_13346);
or U14668 (N_14668,N_13331,N_13959);
xnor U14669 (N_14669,N_13322,N_13826);
and U14670 (N_14670,N_13684,N_13352);
or U14671 (N_14671,N_13768,N_13162);
xor U14672 (N_14672,N_13548,N_13134);
nand U14673 (N_14673,N_13124,N_13715);
nand U14674 (N_14674,N_13038,N_13161);
and U14675 (N_14675,N_13123,N_13902);
nand U14676 (N_14676,N_13946,N_13382);
xor U14677 (N_14677,N_13740,N_13357);
nor U14678 (N_14678,N_13596,N_13391);
xor U14679 (N_14679,N_13157,N_13303);
nand U14680 (N_14680,N_13657,N_13608);
nor U14681 (N_14681,N_13797,N_13504);
nor U14682 (N_14682,N_13752,N_13258);
and U14683 (N_14683,N_13459,N_13909);
nand U14684 (N_14684,N_13574,N_13388);
and U14685 (N_14685,N_13417,N_13984);
or U14686 (N_14686,N_13158,N_13145);
xor U14687 (N_14687,N_13244,N_13048);
nor U14688 (N_14688,N_13362,N_13851);
nor U14689 (N_14689,N_13581,N_13260);
xnor U14690 (N_14690,N_13699,N_13258);
xnor U14691 (N_14691,N_13572,N_13682);
xor U14692 (N_14692,N_13875,N_13647);
xor U14693 (N_14693,N_13911,N_13148);
and U14694 (N_14694,N_13832,N_13584);
xor U14695 (N_14695,N_13441,N_13682);
nor U14696 (N_14696,N_13761,N_13786);
or U14697 (N_14697,N_13098,N_13108);
nand U14698 (N_14698,N_13315,N_13305);
or U14699 (N_14699,N_13118,N_13901);
nor U14700 (N_14700,N_13758,N_13528);
or U14701 (N_14701,N_13386,N_13795);
nand U14702 (N_14702,N_13991,N_13889);
nand U14703 (N_14703,N_13551,N_13020);
xor U14704 (N_14704,N_13788,N_13547);
nand U14705 (N_14705,N_13788,N_13269);
or U14706 (N_14706,N_13176,N_13464);
and U14707 (N_14707,N_13626,N_13056);
nor U14708 (N_14708,N_13822,N_13254);
and U14709 (N_14709,N_13267,N_13944);
nand U14710 (N_14710,N_13019,N_13126);
nand U14711 (N_14711,N_13729,N_13533);
nor U14712 (N_14712,N_13613,N_13794);
nand U14713 (N_14713,N_13698,N_13629);
nor U14714 (N_14714,N_13400,N_13846);
nor U14715 (N_14715,N_13066,N_13517);
nand U14716 (N_14716,N_13474,N_13869);
or U14717 (N_14717,N_13444,N_13667);
or U14718 (N_14718,N_13030,N_13467);
or U14719 (N_14719,N_13687,N_13313);
nand U14720 (N_14720,N_13640,N_13048);
nor U14721 (N_14721,N_13737,N_13002);
or U14722 (N_14722,N_13089,N_13845);
nand U14723 (N_14723,N_13337,N_13815);
nor U14724 (N_14724,N_13923,N_13332);
nor U14725 (N_14725,N_13120,N_13219);
nor U14726 (N_14726,N_13800,N_13028);
xnor U14727 (N_14727,N_13930,N_13686);
or U14728 (N_14728,N_13550,N_13195);
or U14729 (N_14729,N_13026,N_13545);
or U14730 (N_14730,N_13944,N_13157);
or U14731 (N_14731,N_13271,N_13943);
or U14732 (N_14732,N_13703,N_13882);
or U14733 (N_14733,N_13996,N_13036);
and U14734 (N_14734,N_13072,N_13795);
or U14735 (N_14735,N_13376,N_13716);
and U14736 (N_14736,N_13815,N_13581);
nor U14737 (N_14737,N_13265,N_13965);
nand U14738 (N_14738,N_13053,N_13257);
nor U14739 (N_14739,N_13809,N_13629);
xnor U14740 (N_14740,N_13015,N_13349);
nor U14741 (N_14741,N_13865,N_13746);
and U14742 (N_14742,N_13057,N_13847);
or U14743 (N_14743,N_13289,N_13999);
nor U14744 (N_14744,N_13834,N_13503);
nand U14745 (N_14745,N_13575,N_13833);
nand U14746 (N_14746,N_13753,N_13835);
xor U14747 (N_14747,N_13279,N_13826);
nor U14748 (N_14748,N_13500,N_13746);
and U14749 (N_14749,N_13584,N_13997);
xor U14750 (N_14750,N_13521,N_13122);
nor U14751 (N_14751,N_13063,N_13768);
nor U14752 (N_14752,N_13894,N_13958);
xnor U14753 (N_14753,N_13351,N_13572);
nor U14754 (N_14754,N_13100,N_13603);
nor U14755 (N_14755,N_13757,N_13848);
and U14756 (N_14756,N_13583,N_13632);
and U14757 (N_14757,N_13776,N_13061);
and U14758 (N_14758,N_13694,N_13438);
nand U14759 (N_14759,N_13738,N_13432);
xor U14760 (N_14760,N_13365,N_13181);
and U14761 (N_14761,N_13584,N_13144);
nor U14762 (N_14762,N_13305,N_13833);
nor U14763 (N_14763,N_13089,N_13203);
xor U14764 (N_14764,N_13132,N_13765);
xnor U14765 (N_14765,N_13462,N_13925);
or U14766 (N_14766,N_13107,N_13047);
nand U14767 (N_14767,N_13287,N_13006);
or U14768 (N_14768,N_13944,N_13304);
xnor U14769 (N_14769,N_13199,N_13994);
xor U14770 (N_14770,N_13855,N_13020);
nor U14771 (N_14771,N_13581,N_13548);
nand U14772 (N_14772,N_13819,N_13663);
nand U14773 (N_14773,N_13333,N_13271);
nor U14774 (N_14774,N_13415,N_13823);
xnor U14775 (N_14775,N_13133,N_13128);
nand U14776 (N_14776,N_13771,N_13065);
nor U14777 (N_14777,N_13368,N_13824);
xnor U14778 (N_14778,N_13020,N_13397);
nand U14779 (N_14779,N_13341,N_13311);
xnor U14780 (N_14780,N_13980,N_13224);
or U14781 (N_14781,N_13324,N_13357);
xor U14782 (N_14782,N_13228,N_13458);
xnor U14783 (N_14783,N_13576,N_13618);
xor U14784 (N_14784,N_13848,N_13803);
nor U14785 (N_14785,N_13660,N_13480);
nand U14786 (N_14786,N_13696,N_13504);
nand U14787 (N_14787,N_13909,N_13284);
or U14788 (N_14788,N_13778,N_13907);
nor U14789 (N_14789,N_13698,N_13898);
and U14790 (N_14790,N_13694,N_13906);
nor U14791 (N_14791,N_13840,N_13792);
nand U14792 (N_14792,N_13934,N_13397);
and U14793 (N_14793,N_13658,N_13240);
or U14794 (N_14794,N_13071,N_13278);
xnor U14795 (N_14795,N_13526,N_13855);
nand U14796 (N_14796,N_13269,N_13231);
nand U14797 (N_14797,N_13206,N_13049);
nor U14798 (N_14798,N_13964,N_13302);
xnor U14799 (N_14799,N_13931,N_13468);
nor U14800 (N_14800,N_13784,N_13448);
xnor U14801 (N_14801,N_13770,N_13001);
nand U14802 (N_14802,N_13100,N_13351);
or U14803 (N_14803,N_13014,N_13876);
nand U14804 (N_14804,N_13118,N_13580);
nor U14805 (N_14805,N_13182,N_13502);
or U14806 (N_14806,N_13907,N_13603);
or U14807 (N_14807,N_13646,N_13863);
nand U14808 (N_14808,N_13887,N_13881);
xor U14809 (N_14809,N_13438,N_13716);
nand U14810 (N_14810,N_13384,N_13165);
or U14811 (N_14811,N_13463,N_13428);
xnor U14812 (N_14812,N_13897,N_13842);
xnor U14813 (N_14813,N_13403,N_13043);
xnor U14814 (N_14814,N_13140,N_13137);
nand U14815 (N_14815,N_13172,N_13339);
nand U14816 (N_14816,N_13127,N_13191);
nand U14817 (N_14817,N_13555,N_13000);
and U14818 (N_14818,N_13496,N_13431);
nor U14819 (N_14819,N_13691,N_13578);
xnor U14820 (N_14820,N_13927,N_13842);
nand U14821 (N_14821,N_13847,N_13882);
nand U14822 (N_14822,N_13874,N_13102);
and U14823 (N_14823,N_13115,N_13961);
nand U14824 (N_14824,N_13952,N_13659);
nor U14825 (N_14825,N_13805,N_13703);
nand U14826 (N_14826,N_13495,N_13606);
and U14827 (N_14827,N_13249,N_13234);
xnor U14828 (N_14828,N_13110,N_13193);
nor U14829 (N_14829,N_13171,N_13490);
and U14830 (N_14830,N_13010,N_13414);
or U14831 (N_14831,N_13928,N_13648);
nand U14832 (N_14832,N_13913,N_13933);
nor U14833 (N_14833,N_13358,N_13114);
xor U14834 (N_14834,N_13902,N_13086);
xor U14835 (N_14835,N_13332,N_13538);
and U14836 (N_14836,N_13453,N_13707);
and U14837 (N_14837,N_13695,N_13375);
and U14838 (N_14838,N_13796,N_13624);
nor U14839 (N_14839,N_13970,N_13779);
xnor U14840 (N_14840,N_13556,N_13178);
and U14841 (N_14841,N_13037,N_13013);
nor U14842 (N_14842,N_13393,N_13424);
nor U14843 (N_14843,N_13533,N_13187);
or U14844 (N_14844,N_13005,N_13960);
or U14845 (N_14845,N_13771,N_13798);
xor U14846 (N_14846,N_13488,N_13103);
nor U14847 (N_14847,N_13076,N_13436);
nand U14848 (N_14848,N_13086,N_13361);
nor U14849 (N_14849,N_13707,N_13638);
and U14850 (N_14850,N_13246,N_13147);
nand U14851 (N_14851,N_13429,N_13328);
nand U14852 (N_14852,N_13884,N_13641);
and U14853 (N_14853,N_13429,N_13422);
or U14854 (N_14854,N_13428,N_13493);
or U14855 (N_14855,N_13838,N_13702);
xnor U14856 (N_14856,N_13180,N_13330);
or U14857 (N_14857,N_13211,N_13177);
nand U14858 (N_14858,N_13362,N_13108);
nor U14859 (N_14859,N_13951,N_13494);
xnor U14860 (N_14860,N_13505,N_13126);
nand U14861 (N_14861,N_13128,N_13372);
xnor U14862 (N_14862,N_13260,N_13938);
or U14863 (N_14863,N_13982,N_13183);
and U14864 (N_14864,N_13698,N_13539);
xnor U14865 (N_14865,N_13189,N_13693);
or U14866 (N_14866,N_13575,N_13351);
xnor U14867 (N_14867,N_13477,N_13216);
nor U14868 (N_14868,N_13764,N_13564);
nand U14869 (N_14869,N_13319,N_13460);
nand U14870 (N_14870,N_13640,N_13327);
xor U14871 (N_14871,N_13363,N_13565);
xor U14872 (N_14872,N_13722,N_13265);
or U14873 (N_14873,N_13226,N_13775);
and U14874 (N_14874,N_13986,N_13235);
or U14875 (N_14875,N_13434,N_13859);
and U14876 (N_14876,N_13707,N_13748);
nand U14877 (N_14877,N_13655,N_13215);
nand U14878 (N_14878,N_13242,N_13868);
xnor U14879 (N_14879,N_13147,N_13773);
xor U14880 (N_14880,N_13801,N_13910);
and U14881 (N_14881,N_13906,N_13505);
and U14882 (N_14882,N_13735,N_13692);
nand U14883 (N_14883,N_13757,N_13405);
nor U14884 (N_14884,N_13471,N_13357);
and U14885 (N_14885,N_13123,N_13407);
xor U14886 (N_14886,N_13955,N_13767);
nand U14887 (N_14887,N_13830,N_13061);
and U14888 (N_14888,N_13517,N_13206);
nand U14889 (N_14889,N_13034,N_13918);
nand U14890 (N_14890,N_13988,N_13079);
xor U14891 (N_14891,N_13410,N_13841);
nand U14892 (N_14892,N_13442,N_13268);
or U14893 (N_14893,N_13808,N_13329);
nor U14894 (N_14894,N_13361,N_13861);
nor U14895 (N_14895,N_13358,N_13658);
and U14896 (N_14896,N_13685,N_13926);
nand U14897 (N_14897,N_13317,N_13810);
nand U14898 (N_14898,N_13295,N_13140);
or U14899 (N_14899,N_13078,N_13083);
nand U14900 (N_14900,N_13865,N_13222);
xor U14901 (N_14901,N_13745,N_13987);
nor U14902 (N_14902,N_13621,N_13574);
and U14903 (N_14903,N_13298,N_13983);
xor U14904 (N_14904,N_13248,N_13169);
nor U14905 (N_14905,N_13096,N_13168);
nand U14906 (N_14906,N_13136,N_13390);
nor U14907 (N_14907,N_13181,N_13487);
nand U14908 (N_14908,N_13011,N_13993);
and U14909 (N_14909,N_13792,N_13099);
or U14910 (N_14910,N_13186,N_13466);
xnor U14911 (N_14911,N_13847,N_13648);
or U14912 (N_14912,N_13647,N_13124);
nor U14913 (N_14913,N_13840,N_13264);
and U14914 (N_14914,N_13269,N_13568);
and U14915 (N_14915,N_13732,N_13181);
or U14916 (N_14916,N_13517,N_13340);
and U14917 (N_14917,N_13376,N_13064);
xor U14918 (N_14918,N_13238,N_13263);
nor U14919 (N_14919,N_13836,N_13693);
nand U14920 (N_14920,N_13320,N_13971);
nor U14921 (N_14921,N_13560,N_13002);
nand U14922 (N_14922,N_13883,N_13495);
or U14923 (N_14923,N_13333,N_13487);
nand U14924 (N_14924,N_13095,N_13394);
or U14925 (N_14925,N_13556,N_13073);
nor U14926 (N_14926,N_13314,N_13726);
and U14927 (N_14927,N_13597,N_13919);
xnor U14928 (N_14928,N_13541,N_13128);
nor U14929 (N_14929,N_13358,N_13283);
nor U14930 (N_14930,N_13740,N_13456);
and U14931 (N_14931,N_13075,N_13580);
nor U14932 (N_14932,N_13666,N_13288);
nand U14933 (N_14933,N_13328,N_13599);
nand U14934 (N_14934,N_13333,N_13346);
or U14935 (N_14935,N_13735,N_13948);
or U14936 (N_14936,N_13236,N_13995);
nor U14937 (N_14937,N_13181,N_13050);
xor U14938 (N_14938,N_13413,N_13103);
and U14939 (N_14939,N_13196,N_13754);
and U14940 (N_14940,N_13907,N_13762);
and U14941 (N_14941,N_13068,N_13661);
xnor U14942 (N_14942,N_13931,N_13508);
xor U14943 (N_14943,N_13563,N_13255);
nand U14944 (N_14944,N_13904,N_13032);
or U14945 (N_14945,N_13860,N_13605);
xnor U14946 (N_14946,N_13073,N_13727);
nor U14947 (N_14947,N_13410,N_13904);
nor U14948 (N_14948,N_13159,N_13026);
nor U14949 (N_14949,N_13116,N_13869);
xor U14950 (N_14950,N_13516,N_13217);
nor U14951 (N_14951,N_13619,N_13523);
and U14952 (N_14952,N_13810,N_13635);
nand U14953 (N_14953,N_13456,N_13226);
nor U14954 (N_14954,N_13207,N_13478);
or U14955 (N_14955,N_13120,N_13170);
or U14956 (N_14956,N_13028,N_13690);
xor U14957 (N_14957,N_13421,N_13981);
nor U14958 (N_14958,N_13825,N_13622);
xnor U14959 (N_14959,N_13538,N_13799);
or U14960 (N_14960,N_13055,N_13609);
nand U14961 (N_14961,N_13136,N_13018);
nor U14962 (N_14962,N_13267,N_13398);
and U14963 (N_14963,N_13552,N_13860);
xnor U14964 (N_14964,N_13439,N_13046);
nor U14965 (N_14965,N_13552,N_13640);
or U14966 (N_14966,N_13392,N_13654);
or U14967 (N_14967,N_13305,N_13028);
nand U14968 (N_14968,N_13566,N_13998);
or U14969 (N_14969,N_13923,N_13774);
and U14970 (N_14970,N_13187,N_13225);
or U14971 (N_14971,N_13714,N_13962);
nor U14972 (N_14972,N_13387,N_13007);
nor U14973 (N_14973,N_13008,N_13049);
xor U14974 (N_14974,N_13484,N_13538);
xor U14975 (N_14975,N_13914,N_13594);
xor U14976 (N_14976,N_13097,N_13426);
nor U14977 (N_14977,N_13635,N_13415);
and U14978 (N_14978,N_13036,N_13618);
nand U14979 (N_14979,N_13319,N_13306);
nor U14980 (N_14980,N_13459,N_13070);
nor U14981 (N_14981,N_13800,N_13419);
nand U14982 (N_14982,N_13550,N_13008);
nand U14983 (N_14983,N_13352,N_13206);
xor U14984 (N_14984,N_13058,N_13777);
nor U14985 (N_14985,N_13882,N_13237);
xor U14986 (N_14986,N_13122,N_13461);
nor U14987 (N_14987,N_13414,N_13900);
nor U14988 (N_14988,N_13107,N_13170);
nor U14989 (N_14989,N_13532,N_13661);
or U14990 (N_14990,N_13808,N_13921);
nor U14991 (N_14991,N_13372,N_13408);
xnor U14992 (N_14992,N_13955,N_13600);
nor U14993 (N_14993,N_13863,N_13454);
nand U14994 (N_14994,N_13872,N_13119);
and U14995 (N_14995,N_13718,N_13880);
xnor U14996 (N_14996,N_13894,N_13149);
and U14997 (N_14997,N_13528,N_13305);
nand U14998 (N_14998,N_13636,N_13157);
or U14999 (N_14999,N_13195,N_13199);
nor U15000 (N_15000,N_14422,N_14655);
nand U15001 (N_15001,N_14837,N_14957);
or U15002 (N_15002,N_14420,N_14930);
xnor U15003 (N_15003,N_14790,N_14924);
xor U15004 (N_15004,N_14405,N_14386);
nor U15005 (N_15005,N_14016,N_14952);
and U15006 (N_15006,N_14012,N_14281);
nor U15007 (N_15007,N_14528,N_14310);
nor U15008 (N_15008,N_14412,N_14081);
nand U15009 (N_15009,N_14292,N_14305);
nor U15010 (N_15010,N_14427,N_14443);
or U15011 (N_15011,N_14151,N_14185);
or U15012 (N_15012,N_14569,N_14168);
nor U15013 (N_15013,N_14426,N_14803);
or U15014 (N_15014,N_14255,N_14552);
xor U15015 (N_15015,N_14110,N_14159);
or U15016 (N_15016,N_14778,N_14440);
and U15017 (N_15017,N_14107,N_14647);
nand U15018 (N_15018,N_14774,N_14482);
and U15019 (N_15019,N_14002,N_14199);
nand U15020 (N_15020,N_14903,N_14222);
nor U15021 (N_15021,N_14008,N_14949);
xnor U15022 (N_15022,N_14969,N_14929);
nand U15023 (N_15023,N_14864,N_14925);
and U15024 (N_15024,N_14741,N_14200);
nor U15025 (N_15025,N_14376,N_14979);
nand U15026 (N_15026,N_14728,N_14772);
or U15027 (N_15027,N_14373,N_14831);
or U15028 (N_15028,N_14415,N_14001);
nor U15029 (N_15029,N_14239,N_14242);
xnor U15030 (N_15030,N_14411,N_14762);
or U15031 (N_15031,N_14437,N_14716);
nand U15032 (N_15032,N_14184,N_14073);
nand U15033 (N_15033,N_14320,N_14722);
xor U15034 (N_15034,N_14100,N_14613);
or U15035 (N_15035,N_14982,N_14156);
or U15036 (N_15036,N_14153,N_14919);
nand U15037 (N_15037,N_14082,N_14744);
nand U15038 (N_15038,N_14830,N_14083);
or U15039 (N_15039,N_14254,N_14959);
or U15040 (N_15040,N_14840,N_14948);
and U15041 (N_15041,N_14350,N_14288);
nand U15042 (N_15042,N_14692,N_14686);
xor U15043 (N_15043,N_14112,N_14869);
and U15044 (N_15044,N_14379,N_14021);
or U15045 (N_15045,N_14280,N_14032);
nand U15046 (N_15046,N_14985,N_14961);
xor U15047 (N_15047,N_14935,N_14230);
nor U15048 (N_15048,N_14413,N_14589);
and U15049 (N_15049,N_14912,N_14125);
nand U15050 (N_15050,N_14526,N_14852);
xnor U15051 (N_15051,N_14024,N_14534);
and U15052 (N_15052,N_14055,N_14127);
xor U15053 (N_15053,N_14245,N_14357);
xnor U15054 (N_15054,N_14780,N_14901);
and U15055 (N_15055,N_14515,N_14554);
or U15056 (N_15056,N_14769,N_14047);
nand U15057 (N_15057,N_14375,N_14543);
nor U15058 (N_15058,N_14755,N_14758);
nor U15059 (N_15059,N_14171,N_14071);
or U15060 (N_15060,N_14214,N_14459);
nand U15061 (N_15061,N_14216,N_14318);
nor U15062 (N_15062,N_14337,N_14966);
or U15063 (N_15063,N_14074,N_14696);
and U15064 (N_15064,N_14816,N_14968);
and U15065 (N_15065,N_14844,N_14117);
and U15066 (N_15066,N_14879,N_14224);
xnor U15067 (N_15067,N_14633,N_14329);
nand U15068 (N_15068,N_14548,N_14884);
nand U15069 (N_15069,N_14231,N_14389);
nor U15070 (N_15070,N_14394,N_14439);
xnor U15071 (N_15071,N_14701,N_14211);
nand U15072 (N_15072,N_14654,N_14436);
nand U15073 (N_15073,N_14496,N_14177);
and U15074 (N_15074,N_14084,N_14328);
or U15075 (N_15075,N_14981,N_14163);
or U15076 (N_15076,N_14457,N_14409);
xnor U15077 (N_15077,N_14445,N_14727);
xnor U15078 (N_15078,N_14547,N_14279);
or U15079 (N_15079,N_14527,N_14627);
or U15080 (N_15080,N_14616,N_14890);
and U15081 (N_15081,N_14519,N_14210);
or U15082 (N_15082,N_14619,N_14735);
nor U15083 (N_15083,N_14308,N_14581);
nor U15084 (N_15084,N_14804,N_14689);
xnor U15085 (N_15085,N_14808,N_14975);
or U15086 (N_15086,N_14060,N_14250);
xnor U15087 (N_15087,N_14994,N_14223);
xor U15088 (N_15088,N_14011,N_14247);
nor U15089 (N_15089,N_14867,N_14452);
and U15090 (N_15090,N_14567,N_14698);
and U15091 (N_15091,N_14212,N_14737);
or U15092 (N_15092,N_14368,N_14466);
or U15093 (N_15093,N_14046,N_14296);
xor U15094 (N_15094,N_14309,N_14313);
nand U15095 (N_15095,N_14556,N_14304);
and U15096 (N_15096,N_14285,N_14990);
and U15097 (N_15097,N_14180,N_14390);
nand U15098 (N_15098,N_14009,N_14160);
nand U15099 (N_15099,N_14781,N_14150);
xor U15100 (N_15100,N_14586,N_14623);
and U15101 (N_15101,N_14834,N_14612);
and U15102 (N_15102,N_14101,N_14307);
or U15103 (N_15103,N_14656,N_14022);
or U15104 (N_15104,N_14472,N_14905);
nand U15105 (N_15105,N_14723,N_14189);
and U15106 (N_15106,N_14677,N_14710);
nand U15107 (N_15107,N_14511,N_14049);
or U15108 (N_15108,N_14932,N_14766);
xor U15109 (N_15109,N_14020,N_14441);
nand U15110 (N_15110,N_14321,N_14907);
nand U15111 (N_15111,N_14704,N_14461);
or U15112 (N_15112,N_14040,N_14476);
or U15113 (N_15113,N_14237,N_14950);
or U15114 (N_15114,N_14683,N_14372);
nand U15115 (N_15115,N_14401,N_14504);
and U15116 (N_15116,N_14494,N_14743);
xor U15117 (N_15117,N_14585,N_14090);
or U15118 (N_15118,N_14684,N_14395);
xor U15119 (N_15119,N_14227,N_14339);
or U15120 (N_15120,N_14038,N_14518);
xnor U15121 (N_15121,N_14577,N_14617);
xnor U15122 (N_15122,N_14479,N_14871);
or U15123 (N_15123,N_14832,N_14489);
or U15124 (N_15124,N_14414,N_14603);
nand U15125 (N_15125,N_14668,N_14332);
nand U15126 (N_15126,N_14520,N_14785);
xor U15127 (N_15127,N_14103,N_14551);
xor U15128 (N_15128,N_14356,N_14849);
nand U15129 (N_15129,N_14067,N_14809);
nor U15130 (N_15130,N_14480,N_14165);
xnor U15131 (N_15131,N_14407,N_14497);
xnor U15132 (N_15132,N_14186,N_14746);
nor U15133 (N_15133,N_14674,N_14050);
nand U15134 (N_15134,N_14246,N_14642);
xnor U15135 (N_15135,N_14467,N_14039);
nand U15136 (N_15136,N_14017,N_14895);
xnor U15137 (N_15137,N_14815,N_14600);
and U15138 (N_15138,N_14399,N_14207);
or U15139 (N_15139,N_14796,N_14324);
and U15140 (N_15140,N_14491,N_14152);
xnor U15141 (N_15141,N_14665,N_14927);
nor U15142 (N_15142,N_14195,N_14444);
nand U15143 (N_15143,N_14027,N_14419);
nor U15144 (N_15144,N_14141,N_14418);
nor U15145 (N_15145,N_14433,N_14805);
and U15146 (N_15146,N_14825,N_14252);
nor U15147 (N_15147,N_14417,N_14605);
and U15148 (N_15148,N_14161,N_14889);
xor U15149 (N_15149,N_14777,N_14118);
or U15150 (N_15150,N_14971,N_14575);
nor U15151 (N_15151,N_14004,N_14749);
nand U15152 (N_15152,N_14240,N_14899);
or U15153 (N_15153,N_14123,N_14992);
and U15154 (N_15154,N_14828,N_14509);
nand U15155 (N_15155,N_14920,N_14383);
nand U15156 (N_15156,N_14524,N_14000);
nor U15157 (N_15157,N_14469,N_14824);
or U15158 (N_15158,N_14068,N_14505);
xor U15159 (N_15159,N_14611,N_14922);
xor U15160 (N_15160,N_14987,N_14911);
xor U15161 (N_15161,N_14064,N_14442);
or U15162 (N_15162,N_14253,N_14513);
xnor U15163 (N_15163,N_14106,N_14725);
nor U15164 (N_15164,N_14653,N_14814);
and U15165 (N_15165,N_14972,N_14503);
nand U15166 (N_15166,N_14779,N_14051);
and U15167 (N_15167,N_14640,N_14681);
or U15168 (N_15168,N_14388,N_14259);
and U15169 (N_15169,N_14536,N_14102);
or U15170 (N_15170,N_14980,N_14193);
and U15171 (N_15171,N_14198,N_14133);
xnor U15172 (N_15172,N_14649,N_14622);
nand U15173 (N_15173,N_14023,N_14268);
nand U15174 (N_15174,N_14996,N_14587);
or U15175 (N_15175,N_14984,N_14732);
nand U15176 (N_15176,N_14391,N_14063);
xnor U15177 (N_15177,N_14462,N_14842);
nand U15178 (N_15178,N_14841,N_14641);
or U15179 (N_15179,N_14946,N_14558);
and U15180 (N_15180,N_14770,N_14095);
xor U15181 (N_15181,N_14934,N_14178);
nand U15182 (N_15182,N_14345,N_14352);
and U15183 (N_15183,N_14893,N_14314);
nor U15184 (N_15184,N_14059,N_14348);
and U15185 (N_15185,N_14113,N_14977);
nand U15186 (N_15186,N_14187,N_14205);
and U15187 (N_15187,N_14079,N_14155);
nand U15188 (N_15188,N_14602,N_14970);
nand U15189 (N_15189,N_14340,N_14891);
nor U15190 (N_15190,N_14056,N_14578);
nand U15191 (N_15191,N_14190,N_14229);
nor U15192 (N_15192,N_14072,N_14499);
xnor U15193 (N_15193,N_14136,N_14298);
nor U15194 (N_15194,N_14643,N_14848);
nand U15195 (N_15195,N_14974,N_14637);
nor U15196 (N_15196,N_14037,N_14145);
and U15197 (N_15197,N_14069,N_14721);
xnor U15198 (N_15198,N_14300,N_14061);
nor U15199 (N_15199,N_14374,N_14960);
and U15200 (N_15200,N_14474,N_14752);
and U15201 (N_15201,N_14858,N_14546);
nor U15202 (N_15202,N_14826,N_14859);
and U15203 (N_15203,N_14204,N_14030);
xor U15204 (N_15204,N_14299,N_14498);
and U15205 (N_15205,N_14584,N_14460);
nand U15206 (N_15206,N_14438,N_14636);
nand U15207 (N_15207,N_14582,N_14835);
nor U15208 (N_15208,N_14349,N_14175);
nor U15209 (N_15209,N_14998,N_14302);
or U15210 (N_15210,N_14764,N_14776);
xnor U15211 (N_15211,N_14523,N_14731);
nor U15212 (N_15212,N_14219,N_14111);
xnor U15213 (N_15213,N_14691,N_14955);
xnor U15214 (N_15214,N_14688,N_14164);
nand U15215 (N_15215,N_14750,N_14410);
nand U15216 (N_15216,N_14166,N_14364);
xor U15217 (N_15217,N_14351,N_14167);
or U15218 (N_15218,N_14408,N_14289);
nor U15219 (N_15219,N_14392,N_14615);
or U15220 (N_15220,N_14471,N_14042);
or U15221 (N_15221,N_14817,N_14751);
nor U15222 (N_15222,N_14138,N_14316);
or U15223 (N_15223,N_14760,N_14652);
or U15224 (N_15224,N_14277,N_14506);
or U15225 (N_15225,N_14290,N_14286);
xor U15226 (N_15226,N_14666,N_14396);
nand U15227 (N_15227,N_14029,N_14365);
and U15228 (N_15228,N_14378,N_14812);
xor U15229 (N_15229,N_14108,N_14545);
and U15230 (N_15230,N_14174,N_14119);
or U15231 (N_15231,N_14791,N_14745);
or U15232 (N_15232,N_14644,N_14188);
xor U15233 (N_15233,N_14821,N_14789);
nor U15234 (N_15234,N_14624,N_14202);
xor U15235 (N_15235,N_14036,N_14311);
nand U15236 (N_15236,N_14382,N_14909);
or U15237 (N_15237,N_14483,N_14597);
xor U15238 (N_15238,N_14664,N_14659);
xor U15239 (N_15239,N_14713,N_14026);
and U15240 (N_15240,N_14099,N_14147);
or U15241 (N_15241,N_14135,N_14730);
xnor U15242 (N_15242,N_14926,N_14753);
nand U15243 (N_15243,N_14053,N_14724);
nand U15244 (N_15244,N_14976,N_14945);
xnor U15245 (N_15245,N_14048,N_14126);
nor U15246 (N_15246,N_14393,N_14341);
xnor U15247 (N_15247,N_14261,N_14882);
nor U15248 (N_15248,N_14260,N_14435);
and U15249 (N_15249,N_14599,N_14034);
or U15250 (N_15250,N_14986,N_14559);
nor U15251 (N_15251,N_14514,N_14967);
nand U15252 (N_15252,N_14729,N_14470);
xnor U15253 (N_15253,N_14667,N_14455);
or U15254 (N_15254,N_14404,N_14542);
xnor U15255 (N_15255,N_14428,N_14917);
or U15256 (N_15256,N_14784,N_14507);
nand U15257 (N_15257,N_14522,N_14423);
nor U15258 (N_15258,N_14525,N_14276);
nor U15259 (N_15259,N_14293,N_14819);
nor U15260 (N_15260,N_14544,N_14236);
and U15261 (N_15261,N_14645,N_14574);
nor U15262 (N_15262,N_14366,N_14733);
nand U15263 (N_15263,N_14041,N_14266);
or U15264 (N_15264,N_14576,N_14783);
nand U15265 (N_15265,N_14065,N_14275);
xnor U15266 (N_15266,N_14562,N_14323);
and U15267 (N_15267,N_14031,N_14887);
and U15268 (N_15268,N_14456,N_14263);
and U15269 (N_15269,N_14080,N_14402);
or U15270 (N_15270,N_14326,N_14233);
xor U15271 (N_15271,N_14464,N_14820);
nor U15272 (N_15272,N_14282,N_14923);
and U15273 (N_15273,N_14448,N_14468);
nand U15274 (N_15274,N_14991,N_14269);
xor U15275 (N_15275,N_14606,N_14715);
nand U15276 (N_15276,N_14257,N_14109);
xor U15277 (N_15277,N_14303,N_14885);
nand U15278 (N_15278,N_14669,N_14898);
or U15279 (N_15279,N_14788,N_14473);
nand U15280 (N_15280,N_14734,N_14857);
or U15281 (N_15281,N_14854,N_14806);
or U15282 (N_15282,N_14913,N_14104);
nor U15283 (N_15283,N_14873,N_14595);
nor U15284 (N_15284,N_14999,N_14888);
nand U15285 (N_15285,N_14315,N_14590);
and U15286 (N_15286,N_14294,N_14035);
nand U15287 (N_15287,N_14670,N_14897);
nor U15288 (N_15288,N_14580,N_14449);
nor U15289 (N_15289,N_14380,N_14333);
or U15290 (N_15290,N_14014,N_14549);
or U15291 (N_15291,N_14516,N_14880);
xor U15292 (N_15292,N_14338,N_14088);
or U15293 (N_15293,N_14144,N_14661);
nor U15294 (N_15294,N_14771,N_14711);
nor U15295 (N_15295,N_14093,N_14533);
nand U15296 (N_15296,N_14564,N_14209);
nand U15297 (N_15297,N_14902,N_14767);
nor U15298 (N_15298,N_14098,N_14553);
xor U15299 (N_15299,N_14610,N_14863);
nand U15300 (N_15300,N_14823,N_14005);
or U15301 (N_15301,N_14921,N_14192);
nor U15302 (N_15302,N_14134,N_14836);
nor U15303 (N_15303,N_14362,N_14007);
or U15304 (N_15304,N_14742,N_14928);
and U15305 (N_15305,N_14075,N_14856);
and U15306 (N_15306,N_14700,N_14931);
nand U15307 (N_15307,N_14517,N_14601);
nor U15308 (N_15308,N_14978,N_14853);
or U15309 (N_15309,N_14964,N_14572);
xor U15310 (N_15310,N_14381,N_14800);
nor U15311 (N_15311,N_14833,N_14942);
nor U15312 (N_15312,N_14130,N_14486);
and U15313 (N_15313,N_14176,N_14218);
and U15314 (N_15314,N_14400,N_14965);
xor U15315 (N_15315,N_14943,N_14416);
and U15316 (N_15316,N_14086,N_14360);
nand U15317 (N_15317,N_14937,N_14355);
or U15318 (N_15318,N_14620,N_14813);
nand U15319 (N_15319,N_14720,N_14810);
nand U15320 (N_15320,N_14787,N_14485);
and U15321 (N_15321,N_14058,N_14786);
nor U15322 (N_15322,N_14203,N_14262);
nor U15323 (N_15323,N_14874,N_14962);
nand U15324 (N_15324,N_14162,N_14487);
or U15325 (N_15325,N_14675,N_14284);
nand U15326 (N_15326,N_14488,N_14447);
nand U15327 (N_15327,N_14596,N_14588);
and U15328 (N_15328,N_14630,N_14657);
xnor U15329 (N_15329,N_14936,N_14226);
nand U15330 (N_15330,N_14658,N_14648);
and U15331 (N_15331,N_14097,N_14490);
and U15332 (N_15332,N_14274,N_14331);
and U15333 (N_15333,N_14747,N_14122);
nor U15334 (N_15334,N_14353,N_14306);
nor U15335 (N_15335,N_14709,N_14406);
nand U15336 (N_15336,N_14799,N_14561);
and U15337 (N_15337,N_14941,N_14361);
nor U15338 (N_15338,N_14748,N_14702);
nand U15339 (N_15339,N_14451,N_14283);
and U15340 (N_15340,N_14301,N_14217);
xor U15341 (N_15341,N_14078,N_14843);
xor U15342 (N_15342,N_14988,N_14384);
xnor U15343 (N_15343,N_14718,N_14773);
or U15344 (N_15344,N_14697,N_14775);
nor U15345 (N_15345,N_14196,N_14792);
and U15346 (N_15346,N_14215,N_14446);
nor U15347 (N_15347,N_14904,N_14638);
and U15348 (N_15348,N_14875,N_14019);
and U15349 (N_15349,N_14953,N_14827);
and U15350 (N_15350,N_14736,N_14385);
or U15351 (N_15351,N_14695,N_14573);
and U15352 (N_15352,N_14555,N_14956);
xnor U15353 (N_15353,N_14993,N_14765);
nand U15354 (N_15354,N_14502,N_14883);
nor U15355 (N_15355,N_14028,N_14421);
and U15356 (N_15356,N_14272,N_14591);
xnor U15357 (N_15357,N_14557,N_14862);
xnor U15358 (N_15358,N_14248,N_14344);
nor U15359 (N_15359,N_14651,N_14629);
and U15360 (N_15360,N_14132,N_14997);
nand U15361 (N_15361,N_14278,N_14940);
and U15362 (N_15362,N_14908,N_14430);
nor U15363 (N_15363,N_14173,N_14477);
and U15364 (N_15364,N_14481,N_14018);
xnor U15365 (N_15365,N_14954,N_14115);
nor U15366 (N_15366,N_14939,N_14244);
xor U15367 (N_15367,N_14626,N_14197);
and U15368 (N_15368,N_14951,N_14371);
or U15369 (N_15369,N_14521,N_14855);
or U15370 (N_15370,N_14270,N_14432);
nand U15371 (N_15371,N_14845,N_14425);
and U15372 (N_15372,N_14794,N_14592);
or U15373 (N_15373,N_14679,N_14944);
or U15374 (N_15374,N_14738,N_14608);
nand U15375 (N_15375,N_14571,N_14717);
or U15376 (N_15376,N_14094,N_14501);
nor U15377 (N_15377,N_14354,N_14057);
and U15378 (N_15378,N_14958,N_14838);
or U15379 (N_15379,N_14916,N_14708);
nand U15380 (N_15380,N_14662,N_14120);
or U15381 (N_15381,N_14714,N_14628);
nor U15382 (N_15382,N_14170,N_14822);
xor U15383 (N_15383,N_14878,N_14363);
nand U15384 (N_15384,N_14484,N_14811);
nand U15385 (N_15385,N_14369,N_14782);
or U15386 (N_15386,N_14087,N_14264);
xor U15387 (N_15387,N_14172,N_14297);
xor U15388 (N_15388,N_14317,N_14091);
nor U15389 (N_15389,N_14973,N_14033);
and U15390 (N_15390,N_14802,N_14131);
xor U15391 (N_15391,N_14918,N_14757);
xnor U15392 (N_15392,N_14148,N_14671);
nor U15393 (N_15393,N_14829,N_14273);
or U15394 (N_15394,N_14342,N_14876);
and U15395 (N_15395,N_14795,N_14495);
nand U15396 (N_15396,N_14535,N_14492);
and U15397 (N_15397,N_14015,N_14105);
or U15398 (N_15398,N_14798,N_14330);
and U15399 (N_15399,N_14687,N_14872);
nor U15400 (N_15400,N_14915,N_14707);
nor U15401 (N_15401,N_14359,N_14139);
xnor U15402 (N_15402,N_14539,N_14892);
and U15403 (N_15403,N_14847,N_14343);
nor U15404 (N_15404,N_14335,N_14678);
nor U15405 (N_15405,N_14910,N_14010);
xnor U15406 (N_15406,N_14194,N_14763);
nand U15407 (N_15407,N_14249,N_14676);
or U15408 (N_15408,N_14635,N_14672);
or U15409 (N_15409,N_14025,N_14900);
or U15410 (N_15410,N_14191,N_14625);
or U15411 (N_15411,N_14768,N_14705);
nand U15412 (N_15412,N_14756,N_14291);
nor U15413 (N_15413,N_14137,N_14614);
xnor U15414 (N_15414,N_14699,N_14066);
nor U15415 (N_15415,N_14006,N_14241);
xor U15416 (N_15416,N_14358,N_14158);
nand U15417 (N_15417,N_14693,N_14703);
and U15418 (N_15418,N_14225,N_14510);
and U15419 (N_15419,N_14801,N_14850);
nor U15420 (N_15420,N_14650,N_14938);
and U15421 (N_15421,N_14431,N_14865);
and U15422 (N_15422,N_14463,N_14881);
xor U15423 (N_15423,N_14740,N_14963);
and U15424 (N_15424,N_14013,N_14598);
and U15425 (N_15425,N_14673,N_14759);
nor U15426 (N_15426,N_14983,N_14450);
xor U15427 (N_15427,N_14347,N_14201);
or U15428 (N_15428,N_14846,N_14565);
or U15429 (N_15429,N_14243,N_14541);
or U15430 (N_15430,N_14312,N_14458);
or U15431 (N_15431,N_14140,N_14116);
nor U15432 (N_15432,N_14604,N_14726);
xnor U15433 (N_15433,N_14346,N_14256);
and U15434 (N_15434,N_14287,N_14076);
and U15435 (N_15435,N_14870,N_14124);
or U15436 (N_15436,N_14367,N_14807);
nand U15437 (N_15437,N_14114,N_14052);
nor U15438 (N_15438,N_14129,N_14868);
or U15439 (N_15439,N_14685,N_14690);
nor U15440 (N_15440,N_14995,N_14540);
and U15441 (N_15441,N_14866,N_14851);
nor U15442 (N_15442,N_14327,N_14621);
and U15443 (N_15443,N_14563,N_14531);
nor U15444 (N_15444,N_14560,N_14793);
and U15445 (N_15445,N_14706,N_14593);
and U15446 (N_15446,N_14906,N_14512);
xnor U15447 (N_15447,N_14877,N_14493);
nand U15448 (N_15448,N_14797,N_14336);
or U15449 (N_15449,N_14530,N_14054);
xor U15450 (N_15450,N_14478,N_14085);
nor U15451 (N_15451,N_14680,N_14181);
nand U15452 (N_15452,N_14398,N_14183);
xnor U15453 (N_15453,N_14570,N_14465);
nand U15454 (N_15454,N_14634,N_14295);
nand U15455 (N_15455,N_14712,N_14896);
and U15456 (N_15456,N_14894,N_14149);
or U15457 (N_15457,N_14251,N_14609);
and U15458 (N_15458,N_14267,N_14322);
nor U15459 (N_15459,N_14403,N_14397);
xor U15460 (N_15460,N_14377,N_14143);
or U15461 (N_15461,N_14429,N_14003);
and U15462 (N_15462,N_14325,N_14206);
and U15463 (N_15463,N_14594,N_14538);
nor U15464 (N_15464,N_14818,N_14682);
nor U15465 (N_15465,N_14583,N_14537);
and U15466 (N_15466,N_14146,N_14453);
or U15467 (N_15467,N_14089,N_14424);
xnor U15468 (N_15468,N_14265,N_14639);
or U15469 (N_15469,N_14434,N_14062);
nor U15470 (N_15470,N_14121,N_14719);
nand U15471 (N_15471,N_14070,N_14839);
or U15472 (N_15472,N_14500,N_14475);
and U15473 (N_15473,N_14096,N_14142);
xnor U15474 (N_15474,N_14694,N_14607);
nor U15475 (N_15475,N_14454,N_14387);
or U15476 (N_15476,N_14043,N_14234);
nor U15477 (N_15477,N_14213,N_14179);
nor U15478 (N_15478,N_14532,N_14660);
xor U15479 (N_15479,N_14157,N_14566);
and U15480 (N_15480,N_14128,N_14221);
xor U15481 (N_15481,N_14663,N_14860);
xor U15482 (N_15482,N_14319,N_14761);
nand U15483 (N_15483,N_14077,N_14258);
or U15484 (N_15484,N_14220,N_14914);
nor U15485 (N_15485,N_14045,N_14886);
xnor U15486 (N_15486,N_14754,N_14334);
nand U15487 (N_15487,N_14529,N_14208);
and U15488 (N_15488,N_14370,N_14861);
nand U15489 (N_15489,N_14154,N_14646);
nand U15490 (N_15490,N_14235,N_14579);
and U15491 (N_15491,N_14228,N_14989);
nor U15492 (N_15492,N_14933,N_14044);
nor U15493 (N_15493,N_14550,N_14169);
or U15494 (N_15494,N_14508,N_14618);
and U15495 (N_15495,N_14092,N_14739);
or U15496 (N_15496,N_14631,N_14238);
and U15497 (N_15497,N_14232,N_14947);
nand U15498 (N_15498,N_14568,N_14271);
nor U15499 (N_15499,N_14182,N_14632);
and U15500 (N_15500,N_14840,N_14195);
and U15501 (N_15501,N_14341,N_14420);
or U15502 (N_15502,N_14193,N_14639);
or U15503 (N_15503,N_14255,N_14479);
xnor U15504 (N_15504,N_14806,N_14061);
nand U15505 (N_15505,N_14485,N_14554);
or U15506 (N_15506,N_14290,N_14798);
and U15507 (N_15507,N_14904,N_14088);
nor U15508 (N_15508,N_14964,N_14045);
xnor U15509 (N_15509,N_14083,N_14046);
and U15510 (N_15510,N_14597,N_14530);
nor U15511 (N_15511,N_14008,N_14481);
nand U15512 (N_15512,N_14192,N_14684);
nor U15513 (N_15513,N_14670,N_14779);
nor U15514 (N_15514,N_14277,N_14751);
and U15515 (N_15515,N_14639,N_14434);
and U15516 (N_15516,N_14566,N_14470);
nor U15517 (N_15517,N_14944,N_14447);
nand U15518 (N_15518,N_14144,N_14918);
xor U15519 (N_15519,N_14005,N_14129);
xnor U15520 (N_15520,N_14627,N_14659);
nor U15521 (N_15521,N_14455,N_14821);
nor U15522 (N_15522,N_14977,N_14735);
nor U15523 (N_15523,N_14806,N_14762);
and U15524 (N_15524,N_14478,N_14266);
and U15525 (N_15525,N_14361,N_14338);
nor U15526 (N_15526,N_14489,N_14177);
nand U15527 (N_15527,N_14565,N_14288);
xnor U15528 (N_15528,N_14447,N_14773);
nand U15529 (N_15529,N_14527,N_14004);
and U15530 (N_15530,N_14476,N_14389);
xor U15531 (N_15531,N_14515,N_14149);
and U15532 (N_15532,N_14781,N_14461);
nand U15533 (N_15533,N_14256,N_14372);
nor U15534 (N_15534,N_14798,N_14968);
or U15535 (N_15535,N_14550,N_14283);
nand U15536 (N_15536,N_14420,N_14177);
and U15537 (N_15537,N_14202,N_14319);
nand U15538 (N_15538,N_14235,N_14947);
nand U15539 (N_15539,N_14854,N_14913);
and U15540 (N_15540,N_14107,N_14457);
xnor U15541 (N_15541,N_14211,N_14244);
nor U15542 (N_15542,N_14249,N_14239);
or U15543 (N_15543,N_14957,N_14373);
and U15544 (N_15544,N_14681,N_14902);
and U15545 (N_15545,N_14705,N_14555);
nand U15546 (N_15546,N_14199,N_14005);
xnor U15547 (N_15547,N_14151,N_14226);
nor U15548 (N_15548,N_14137,N_14939);
nor U15549 (N_15549,N_14354,N_14041);
or U15550 (N_15550,N_14654,N_14472);
xnor U15551 (N_15551,N_14345,N_14757);
and U15552 (N_15552,N_14288,N_14162);
or U15553 (N_15553,N_14048,N_14487);
or U15554 (N_15554,N_14779,N_14416);
xnor U15555 (N_15555,N_14410,N_14874);
nor U15556 (N_15556,N_14509,N_14737);
nand U15557 (N_15557,N_14441,N_14088);
and U15558 (N_15558,N_14991,N_14547);
nor U15559 (N_15559,N_14299,N_14155);
and U15560 (N_15560,N_14800,N_14974);
and U15561 (N_15561,N_14114,N_14851);
and U15562 (N_15562,N_14282,N_14048);
or U15563 (N_15563,N_14754,N_14551);
nor U15564 (N_15564,N_14011,N_14047);
xnor U15565 (N_15565,N_14744,N_14703);
or U15566 (N_15566,N_14851,N_14319);
nand U15567 (N_15567,N_14553,N_14170);
and U15568 (N_15568,N_14827,N_14030);
nand U15569 (N_15569,N_14158,N_14929);
xnor U15570 (N_15570,N_14450,N_14753);
nor U15571 (N_15571,N_14153,N_14197);
nor U15572 (N_15572,N_14653,N_14735);
nor U15573 (N_15573,N_14567,N_14959);
and U15574 (N_15574,N_14026,N_14679);
nand U15575 (N_15575,N_14469,N_14042);
nand U15576 (N_15576,N_14285,N_14725);
nor U15577 (N_15577,N_14813,N_14323);
nand U15578 (N_15578,N_14461,N_14652);
nor U15579 (N_15579,N_14685,N_14082);
or U15580 (N_15580,N_14909,N_14049);
or U15581 (N_15581,N_14455,N_14744);
and U15582 (N_15582,N_14018,N_14518);
nand U15583 (N_15583,N_14364,N_14708);
xnor U15584 (N_15584,N_14930,N_14159);
nand U15585 (N_15585,N_14491,N_14929);
xor U15586 (N_15586,N_14328,N_14670);
nor U15587 (N_15587,N_14361,N_14550);
or U15588 (N_15588,N_14530,N_14555);
nand U15589 (N_15589,N_14678,N_14635);
nor U15590 (N_15590,N_14057,N_14422);
nor U15591 (N_15591,N_14532,N_14264);
and U15592 (N_15592,N_14521,N_14036);
nand U15593 (N_15593,N_14331,N_14868);
or U15594 (N_15594,N_14228,N_14859);
nor U15595 (N_15595,N_14923,N_14894);
xor U15596 (N_15596,N_14407,N_14761);
nor U15597 (N_15597,N_14356,N_14298);
and U15598 (N_15598,N_14538,N_14688);
nor U15599 (N_15599,N_14835,N_14695);
nand U15600 (N_15600,N_14563,N_14106);
and U15601 (N_15601,N_14450,N_14170);
and U15602 (N_15602,N_14050,N_14904);
and U15603 (N_15603,N_14543,N_14814);
nand U15604 (N_15604,N_14325,N_14811);
nor U15605 (N_15605,N_14355,N_14834);
nor U15606 (N_15606,N_14635,N_14109);
nand U15607 (N_15607,N_14726,N_14622);
xnor U15608 (N_15608,N_14226,N_14380);
nor U15609 (N_15609,N_14606,N_14351);
or U15610 (N_15610,N_14948,N_14395);
nand U15611 (N_15611,N_14659,N_14616);
or U15612 (N_15612,N_14022,N_14300);
or U15613 (N_15613,N_14065,N_14468);
nor U15614 (N_15614,N_14296,N_14068);
nand U15615 (N_15615,N_14744,N_14182);
xor U15616 (N_15616,N_14229,N_14063);
nand U15617 (N_15617,N_14754,N_14310);
or U15618 (N_15618,N_14481,N_14594);
nor U15619 (N_15619,N_14932,N_14206);
and U15620 (N_15620,N_14895,N_14437);
or U15621 (N_15621,N_14983,N_14048);
or U15622 (N_15622,N_14534,N_14527);
and U15623 (N_15623,N_14074,N_14719);
or U15624 (N_15624,N_14008,N_14423);
nand U15625 (N_15625,N_14149,N_14730);
nand U15626 (N_15626,N_14652,N_14879);
nor U15627 (N_15627,N_14202,N_14051);
xor U15628 (N_15628,N_14461,N_14747);
and U15629 (N_15629,N_14779,N_14560);
and U15630 (N_15630,N_14378,N_14525);
nand U15631 (N_15631,N_14582,N_14011);
xor U15632 (N_15632,N_14555,N_14332);
nand U15633 (N_15633,N_14823,N_14203);
and U15634 (N_15634,N_14453,N_14590);
and U15635 (N_15635,N_14742,N_14776);
nor U15636 (N_15636,N_14360,N_14569);
and U15637 (N_15637,N_14813,N_14106);
and U15638 (N_15638,N_14873,N_14615);
nand U15639 (N_15639,N_14213,N_14122);
xor U15640 (N_15640,N_14238,N_14744);
or U15641 (N_15641,N_14152,N_14338);
or U15642 (N_15642,N_14725,N_14803);
xnor U15643 (N_15643,N_14650,N_14391);
nor U15644 (N_15644,N_14527,N_14613);
nor U15645 (N_15645,N_14015,N_14090);
nor U15646 (N_15646,N_14830,N_14117);
or U15647 (N_15647,N_14111,N_14863);
or U15648 (N_15648,N_14152,N_14981);
xor U15649 (N_15649,N_14975,N_14329);
xnor U15650 (N_15650,N_14557,N_14438);
or U15651 (N_15651,N_14355,N_14111);
or U15652 (N_15652,N_14584,N_14554);
nand U15653 (N_15653,N_14210,N_14380);
and U15654 (N_15654,N_14902,N_14051);
or U15655 (N_15655,N_14718,N_14213);
and U15656 (N_15656,N_14700,N_14651);
or U15657 (N_15657,N_14566,N_14207);
xnor U15658 (N_15658,N_14615,N_14918);
nand U15659 (N_15659,N_14480,N_14867);
and U15660 (N_15660,N_14700,N_14155);
nor U15661 (N_15661,N_14102,N_14425);
or U15662 (N_15662,N_14374,N_14362);
nor U15663 (N_15663,N_14432,N_14328);
nand U15664 (N_15664,N_14249,N_14255);
and U15665 (N_15665,N_14938,N_14863);
nand U15666 (N_15666,N_14156,N_14147);
and U15667 (N_15667,N_14996,N_14591);
nor U15668 (N_15668,N_14847,N_14635);
xnor U15669 (N_15669,N_14305,N_14274);
nand U15670 (N_15670,N_14828,N_14730);
nand U15671 (N_15671,N_14154,N_14533);
or U15672 (N_15672,N_14039,N_14999);
or U15673 (N_15673,N_14551,N_14467);
nor U15674 (N_15674,N_14094,N_14227);
and U15675 (N_15675,N_14163,N_14237);
xor U15676 (N_15676,N_14489,N_14844);
nand U15677 (N_15677,N_14192,N_14038);
xnor U15678 (N_15678,N_14317,N_14110);
or U15679 (N_15679,N_14842,N_14937);
nor U15680 (N_15680,N_14811,N_14384);
or U15681 (N_15681,N_14339,N_14154);
xor U15682 (N_15682,N_14303,N_14642);
xnor U15683 (N_15683,N_14987,N_14518);
nor U15684 (N_15684,N_14875,N_14066);
and U15685 (N_15685,N_14708,N_14700);
and U15686 (N_15686,N_14778,N_14349);
nand U15687 (N_15687,N_14079,N_14095);
and U15688 (N_15688,N_14720,N_14291);
and U15689 (N_15689,N_14692,N_14964);
and U15690 (N_15690,N_14343,N_14721);
nor U15691 (N_15691,N_14162,N_14181);
nand U15692 (N_15692,N_14327,N_14147);
nand U15693 (N_15693,N_14467,N_14465);
xnor U15694 (N_15694,N_14884,N_14271);
nand U15695 (N_15695,N_14668,N_14450);
xor U15696 (N_15696,N_14089,N_14358);
xor U15697 (N_15697,N_14849,N_14168);
and U15698 (N_15698,N_14171,N_14650);
or U15699 (N_15699,N_14197,N_14289);
nand U15700 (N_15700,N_14046,N_14718);
and U15701 (N_15701,N_14181,N_14362);
nand U15702 (N_15702,N_14121,N_14445);
xnor U15703 (N_15703,N_14610,N_14130);
or U15704 (N_15704,N_14883,N_14685);
nor U15705 (N_15705,N_14020,N_14427);
or U15706 (N_15706,N_14628,N_14890);
or U15707 (N_15707,N_14968,N_14850);
nor U15708 (N_15708,N_14204,N_14661);
nand U15709 (N_15709,N_14655,N_14970);
xor U15710 (N_15710,N_14266,N_14233);
nand U15711 (N_15711,N_14516,N_14787);
nor U15712 (N_15712,N_14597,N_14646);
nand U15713 (N_15713,N_14435,N_14387);
xnor U15714 (N_15714,N_14083,N_14713);
and U15715 (N_15715,N_14091,N_14602);
and U15716 (N_15716,N_14291,N_14039);
nand U15717 (N_15717,N_14759,N_14107);
or U15718 (N_15718,N_14564,N_14731);
xnor U15719 (N_15719,N_14752,N_14779);
nor U15720 (N_15720,N_14624,N_14258);
and U15721 (N_15721,N_14604,N_14570);
nand U15722 (N_15722,N_14405,N_14127);
xor U15723 (N_15723,N_14325,N_14676);
or U15724 (N_15724,N_14790,N_14946);
nand U15725 (N_15725,N_14939,N_14258);
and U15726 (N_15726,N_14347,N_14177);
or U15727 (N_15727,N_14145,N_14899);
nor U15728 (N_15728,N_14773,N_14590);
and U15729 (N_15729,N_14356,N_14719);
or U15730 (N_15730,N_14669,N_14445);
or U15731 (N_15731,N_14583,N_14784);
xnor U15732 (N_15732,N_14351,N_14811);
and U15733 (N_15733,N_14460,N_14388);
or U15734 (N_15734,N_14170,N_14929);
nor U15735 (N_15735,N_14124,N_14720);
nor U15736 (N_15736,N_14704,N_14221);
nor U15737 (N_15737,N_14389,N_14129);
nand U15738 (N_15738,N_14681,N_14358);
nand U15739 (N_15739,N_14360,N_14631);
xnor U15740 (N_15740,N_14792,N_14532);
and U15741 (N_15741,N_14623,N_14939);
nor U15742 (N_15742,N_14422,N_14417);
or U15743 (N_15743,N_14379,N_14283);
and U15744 (N_15744,N_14643,N_14313);
nand U15745 (N_15745,N_14439,N_14389);
or U15746 (N_15746,N_14124,N_14246);
nor U15747 (N_15747,N_14197,N_14622);
xor U15748 (N_15748,N_14753,N_14240);
nor U15749 (N_15749,N_14597,N_14684);
nand U15750 (N_15750,N_14980,N_14799);
and U15751 (N_15751,N_14350,N_14021);
nand U15752 (N_15752,N_14882,N_14720);
and U15753 (N_15753,N_14638,N_14047);
nand U15754 (N_15754,N_14908,N_14048);
and U15755 (N_15755,N_14677,N_14578);
nor U15756 (N_15756,N_14077,N_14057);
xor U15757 (N_15757,N_14434,N_14879);
nor U15758 (N_15758,N_14209,N_14633);
xor U15759 (N_15759,N_14493,N_14593);
nand U15760 (N_15760,N_14742,N_14146);
nand U15761 (N_15761,N_14813,N_14715);
xnor U15762 (N_15762,N_14498,N_14465);
nand U15763 (N_15763,N_14995,N_14381);
nor U15764 (N_15764,N_14043,N_14672);
xor U15765 (N_15765,N_14350,N_14116);
or U15766 (N_15766,N_14246,N_14269);
and U15767 (N_15767,N_14928,N_14598);
nor U15768 (N_15768,N_14363,N_14471);
nor U15769 (N_15769,N_14477,N_14669);
nand U15770 (N_15770,N_14395,N_14228);
and U15771 (N_15771,N_14119,N_14838);
nor U15772 (N_15772,N_14168,N_14236);
and U15773 (N_15773,N_14295,N_14863);
nor U15774 (N_15774,N_14032,N_14381);
nor U15775 (N_15775,N_14794,N_14912);
nor U15776 (N_15776,N_14600,N_14997);
nand U15777 (N_15777,N_14420,N_14655);
and U15778 (N_15778,N_14269,N_14025);
nor U15779 (N_15779,N_14587,N_14741);
nand U15780 (N_15780,N_14517,N_14491);
xor U15781 (N_15781,N_14274,N_14821);
nand U15782 (N_15782,N_14331,N_14103);
nand U15783 (N_15783,N_14002,N_14459);
or U15784 (N_15784,N_14425,N_14802);
or U15785 (N_15785,N_14636,N_14703);
nor U15786 (N_15786,N_14904,N_14812);
nand U15787 (N_15787,N_14021,N_14667);
and U15788 (N_15788,N_14242,N_14594);
nand U15789 (N_15789,N_14288,N_14776);
xor U15790 (N_15790,N_14176,N_14891);
or U15791 (N_15791,N_14643,N_14709);
nor U15792 (N_15792,N_14051,N_14460);
xnor U15793 (N_15793,N_14643,N_14952);
or U15794 (N_15794,N_14942,N_14730);
and U15795 (N_15795,N_14420,N_14191);
nand U15796 (N_15796,N_14157,N_14064);
or U15797 (N_15797,N_14155,N_14266);
nor U15798 (N_15798,N_14744,N_14053);
and U15799 (N_15799,N_14842,N_14945);
nand U15800 (N_15800,N_14839,N_14734);
nand U15801 (N_15801,N_14723,N_14857);
nor U15802 (N_15802,N_14582,N_14169);
and U15803 (N_15803,N_14293,N_14730);
or U15804 (N_15804,N_14620,N_14217);
and U15805 (N_15805,N_14702,N_14524);
and U15806 (N_15806,N_14472,N_14915);
or U15807 (N_15807,N_14063,N_14174);
nand U15808 (N_15808,N_14003,N_14525);
nor U15809 (N_15809,N_14637,N_14396);
and U15810 (N_15810,N_14080,N_14973);
or U15811 (N_15811,N_14094,N_14764);
nand U15812 (N_15812,N_14770,N_14156);
nor U15813 (N_15813,N_14762,N_14090);
xor U15814 (N_15814,N_14018,N_14447);
nand U15815 (N_15815,N_14168,N_14882);
and U15816 (N_15816,N_14260,N_14360);
nand U15817 (N_15817,N_14464,N_14998);
xor U15818 (N_15818,N_14811,N_14181);
nand U15819 (N_15819,N_14550,N_14955);
nor U15820 (N_15820,N_14018,N_14102);
nor U15821 (N_15821,N_14876,N_14243);
nand U15822 (N_15822,N_14571,N_14076);
nand U15823 (N_15823,N_14697,N_14258);
nor U15824 (N_15824,N_14523,N_14891);
and U15825 (N_15825,N_14958,N_14226);
nor U15826 (N_15826,N_14884,N_14979);
xnor U15827 (N_15827,N_14521,N_14181);
nor U15828 (N_15828,N_14093,N_14412);
or U15829 (N_15829,N_14963,N_14187);
nand U15830 (N_15830,N_14654,N_14506);
and U15831 (N_15831,N_14493,N_14893);
nor U15832 (N_15832,N_14324,N_14290);
and U15833 (N_15833,N_14938,N_14993);
nand U15834 (N_15834,N_14657,N_14398);
xor U15835 (N_15835,N_14270,N_14756);
or U15836 (N_15836,N_14973,N_14083);
or U15837 (N_15837,N_14881,N_14681);
and U15838 (N_15838,N_14381,N_14591);
nand U15839 (N_15839,N_14325,N_14860);
and U15840 (N_15840,N_14350,N_14323);
xnor U15841 (N_15841,N_14435,N_14868);
or U15842 (N_15842,N_14450,N_14224);
nand U15843 (N_15843,N_14765,N_14899);
nand U15844 (N_15844,N_14145,N_14435);
or U15845 (N_15845,N_14951,N_14139);
xnor U15846 (N_15846,N_14806,N_14923);
or U15847 (N_15847,N_14719,N_14061);
nand U15848 (N_15848,N_14918,N_14650);
nor U15849 (N_15849,N_14986,N_14228);
nand U15850 (N_15850,N_14877,N_14660);
xor U15851 (N_15851,N_14651,N_14474);
or U15852 (N_15852,N_14657,N_14991);
and U15853 (N_15853,N_14560,N_14762);
and U15854 (N_15854,N_14034,N_14635);
xnor U15855 (N_15855,N_14095,N_14234);
nor U15856 (N_15856,N_14840,N_14593);
and U15857 (N_15857,N_14741,N_14117);
and U15858 (N_15858,N_14260,N_14576);
nand U15859 (N_15859,N_14972,N_14058);
and U15860 (N_15860,N_14111,N_14597);
xnor U15861 (N_15861,N_14041,N_14173);
and U15862 (N_15862,N_14917,N_14670);
nand U15863 (N_15863,N_14333,N_14969);
xor U15864 (N_15864,N_14481,N_14443);
xnor U15865 (N_15865,N_14349,N_14036);
xor U15866 (N_15866,N_14148,N_14878);
and U15867 (N_15867,N_14678,N_14939);
and U15868 (N_15868,N_14922,N_14526);
or U15869 (N_15869,N_14380,N_14754);
or U15870 (N_15870,N_14967,N_14104);
xor U15871 (N_15871,N_14970,N_14977);
and U15872 (N_15872,N_14321,N_14658);
nand U15873 (N_15873,N_14069,N_14241);
xor U15874 (N_15874,N_14034,N_14025);
xnor U15875 (N_15875,N_14127,N_14275);
or U15876 (N_15876,N_14904,N_14124);
nand U15877 (N_15877,N_14243,N_14845);
or U15878 (N_15878,N_14759,N_14399);
and U15879 (N_15879,N_14585,N_14986);
or U15880 (N_15880,N_14561,N_14393);
or U15881 (N_15881,N_14808,N_14756);
or U15882 (N_15882,N_14712,N_14723);
nand U15883 (N_15883,N_14890,N_14604);
or U15884 (N_15884,N_14679,N_14190);
or U15885 (N_15885,N_14911,N_14582);
and U15886 (N_15886,N_14702,N_14043);
nor U15887 (N_15887,N_14454,N_14029);
and U15888 (N_15888,N_14907,N_14707);
and U15889 (N_15889,N_14802,N_14443);
xnor U15890 (N_15890,N_14785,N_14105);
nand U15891 (N_15891,N_14790,N_14110);
nand U15892 (N_15892,N_14184,N_14957);
nor U15893 (N_15893,N_14501,N_14310);
xnor U15894 (N_15894,N_14374,N_14323);
nand U15895 (N_15895,N_14785,N_14673);
xor U15896 (N_15896,N_14654,N_14014);
or U15897 (N_15897,N_14317,N_14491);
and U15898 (N_15898,N_14807,N_14737);
xor U15899 (N_15899,N_14389,N_14271);
nand U15900 (N_15900,N_14687,N_14576);
nand U15901 (N_15901,N_14043,N_14549);
nor U15902 (N_15902,N_14990,N_14346);
nor U15903 (N_15903,N_14665,N_14491);
nand U15904 (N_15904,N_14940,N_14527);
nor U15905 (N_15905,N_14613,N_14642);
nand U15906 (N_15906,N_14431,N_14854);
and U15907 (N_15907,N_14657,N_14641);
and U15908 (N_15908,N_14289,N_14990);
xor U15909 (N_15909,N_14073,N_14588);
or U15910 (N_15910,N_14462,N_14368);
nand U15911 (N_15911,N_14358,N_14822);
and U15912 (N_15912,N_14372,N_14919);
or U15913 (N_15913,N_14251,N_14134);
xnor U15914 (N_15914,N_14475,N_14523);
nand U15915 (N_15915,N_14320,N_14065);
and U15916 (N_15916,N_14989,N_14775);
xor U15917 (N_15917,N_14237,N_14132);
or U15918 (N_15918,N_14991,N_14406);
nor U15919 (N_15919,N_14678,N_14751);
or U15920 (N_15920,N_14664,N_14408);
and U15921 (N_15921,N_14915,N_14362);
nor U15922 (N_15922,N_14388,N_14474);
nand U15923 (N_15923,N_14757,N_14104);
nor U15924 (N_15924,N_14422,N_14538);
nand U15925 (N_15925,N_14307,N_14606);
and U15926 (N_15926,N_14592,N_14107);
nor U15927 (N_15927,N_14108,N_14529);
nor U15928 (N_15928,N_14176,N_14982);
nor U15929 (N_15929,N_14038,N_14189);
nor U15930 (N_15930,N_14170,N_14230);
nand U15931 (N_15931,N_14624,N_14557);
nand U15932 (N_15932,N_14743,N_14490);
and U15933 (N_15933,N_14356,N_14831);
nor U15934 (N_15934,N_14563,N_14464);
or U15935 (N_15935,N_14639,N_14819);
nand U15936 (N_15936,N_14404,N_14348);
and U15937 (N_15937,N_14644,N_14160);
nand U15938 (N_15938,N_14306,N_14474);
xnor U15939 (N_15939,N_14390,N_14284);
and U15940 (N_15940,N_14386,N_14665);
nor U15941 (N_15941,N_14054,N_14693);
nor U15942 (N_15942,N_14871,N_14949);
xor U15943 (N_15943,N_14914,N_14330);
nor U15944 (N_15944,N_14428,N_14570);
and U15945 (N_15945,N_14931,N_14958);
and U15946 (N_15946,N_14798,N_14584);
or U15947 (N_15947,N_14772,N_14024);
nor U15948 (N_15948,N_14209,N_14833);
nor U15949 (N_15949,N_14430,N_14229);
nand U15950 (N_15950,N_14166,N_14902);
and U15951 (N_15951,N_14143,N_14706);
and U15952 (N_15952,N_14238,N_14529);
or U15953 (N_15953,N_14552,N_14557);
or U15954 (N_15954,N_14394,N_14021);
or U15955 (N_15955,N_14727,N_14864);
and U15956 (N_15956,N_14994,N_14069);
xor U15957 (N_15957,N_14895,N_14105);
or U15958 (N_15958,N_14618,N_14652);
nand U15959 (N_15959,N_14322,N_14487);
and U15960 (N_15960,N_14246,N_14169);
nand U15961 (N_15961,N_14021,N_14148);
or U15962 (N_15962,N_14495,N_14104);
nand U15963 (N_15963,N_14719,N_14989);
nor U15964 (N_15964,N_14959,N_14350);
xnor U15965 (N_15965,N_14609,N_14005);
and U15966 (N_15966,N_14838,N_14303);
nand U15967 (N_15967,N_14182,N_14316);
xor U15968 (N_15968,N_14720,N_14460);
and U15969 (N_15969,N_14862,N_14555);
nand U15970 (N_15970,N_14194,N_14001);
nor U15971 (N_15971,N_14189,N_14389);
nand U15972 (N_15972,N_14651,N_14322);
xor U15973 (N_15973,N_14088,N_14882);
nand U15974 (N_15974,N_14105,N_14001);
and U15975 (N_15975,N_14194,N_14729);
nand U15976 (N_15976,N_14849,N_14301);
and U15977 (N_15977,N_14966,N_14011);
nor U15978 (N_15978,N_14112,N_14888);
xor U15979 (N_15979,N_14932,N_14577);
nor U15980 (N_15980,N_14805,N_14718);
xnor U15981 (N_15981,N_14817,N_14025);
nor U15982 (N_15982,N_14286,N_14912);
nand U15983 (N_15983,N_14301,N_14905);
nor U15984 (N_15984,N_14300,N_14923);
nor U15985 (N_15985,N_14138,N_14613);
nor U15986 (N_15986,N_14764,N_14760);
nand U15987 (N_15987,N_14972,N_14984);
or U15988 (N_15988,N_14540,N_14216);
or U15989 (N_15989,N_14652,N_14089);
or U15990 (N_15990,N_14853,N_14657);
nor U15991 (N_15991,N_14930,N_14627);
xnor U15992 (N_15992,N_14421,N_14979);
xor U15993 (N_15993,N_14777,N_14546);
nor U15994 (N_15994,N_14897,N_14823);
nor U15995 (N_15995,N_14814,N_14203);
and U15996 (N_15996,N_14454,N_14503);
nor U15997 (N_15997,N_14325,N_14804);
nand U15998 (N_15998,N_14081,N_14737);
xnor U15999 (N_15999,N_14841,N_14732);
nand U16000 (N_16000,N_15936,N_15209);
or U16001 (N_16001,N_15875,N_15431);
nand U16002 (N_16002,N_15592,N_15728);
nand U16003 (N_16003,N_15811,N_15471);
and U16004 (N_16004,N_15435,N_15814);
or U16005 (N_16005,N_15798,N_15323);
nand U16006 (N_16006,N_15862,N_15355);
nand U16007 (N_16007,N_15660,N_15681);
nor U16008 (N_16008,N_15813,N_15043);
nor U16009 (N_16009,N_15468,N_15670);
or U16010 (N_16010,N_15595,N_15159);
xor U16011 (N_16011,N_15881,N_15910);
xor U16012 (N_16012,N_15416,N_15509);
or U16013 (N_16013,N_15842,N_15917);
and U16014 (N_16014,N_15121,N_15089);
or U16015 (N_16015,N_15008,N_15408);
xor U16016 (N_16016,N_15107,N_15099);
nand U16017 (N_16017,N_15083,N_15488);
xor U16018 (N_16018,N_15604,N_15826);
xor U16019 (N_16019,N_15919,N_15596);
or U16020 (N_16020,N_15343,N_15432);
nor U16021 (N_16021,N_15791,N_15329);
nand U16022 (N_16022,N_15539,N_15401);
and U16023 (N_16023,N_15087,N_15244);
nor U16024 (N_16024,N_15508,N_15652);
nor U16025 (N_16025,N_15748,N_15450);
nor U16026 (N_16026,N_15672,N_15852);
nand U16027 (N_16027,N_15319,N_15016);
and U16028 (N_16028,N_15983,N_15800);
nor U16029 (N_16029,N_15196,N_15533);
nor U16030 (N_16030,N_15184,N_15033);
or U16031 (N_16031,N_15048,N_15760);
and U16032 (N_16032,N_15393,N_15040);
nor U16033 (N_16033,N_15897,N_15141);
xor U16034 (N_16034,N_15844,N_15402);
nor U16035 (N_16035,N_15603,N_15927);
nand U16036 (N_16036,N_15618,N_15258);
nand U16037 (N_16037,N_15105,N_15286);
nand U16038 (N_16038,N_15017,N_15893);
nand U16039 (N_16039,N_15808,N_15149);
nor U16040 (N_16040,N_15625,N_15487);
nand U16041 (N_16041,N_15536,N_15654);
or U16042 (N_16042,N_15578,N_15322);
nor U16043 (N_16043,N_15207,N_15552);
xnor U16044 (N_16044,N_15250,N_15366);
nor U16045 (N_16045,N_15839,N_15352);
and U16046 (N_16046,N_15550,N_15115);
or U16047 (N_16047,N_15002,N_15377);
or U16048 (N_16048,N_15986,N_15540);
xor U16049 (N_16049,N_15415,N_15441);
nand U16050 (N_16050,N_15980,N_15133);
nor U16051 (N_16051,N_15677,N_15421);
xnor U16052 (N_16052,N_15695,N_15277);
nor U16053 (N_16053,N_15104,N_15753);
nand U16054 (N_16054,N_15650,N_15489);
xor U16055 (N_16055,N_15890,N_15187);
nor U16056 (N_16056,N_15887,N_15920);
nor U16057 (N_16057,N_15111,N_15679);
xnor U16058 (N_16058,N_15264,N_15123);
xnor U16059 (N_16059,N_15263,N_15397);
and U16060 (N_16060,N_15470,N_15374);
or U16061 (N_16061,N_15417,N_15231);
nand U16062 (N_16062,N_15720,N_15195);
or U16063 (N_16063,N_15061,N_15546);
nand U16064 (N_16064,N_15460,N_15532);
or U16065 (N_16065,N_15392,N_15294);
or U16066 (N_16066,N_15062,N_15372);
or U16067 (N_16067,N_15100,N_15590);
or U16068 (N_16068,N_15032,N_15758);
nand U16069 (N_16069,N_15741,N_15621);
xor U16070 (N_16070,N_15136,N_15205);
and U16071 (N_16071,N_15406,N_15499);
or U16072 (N_16072,N_15714,N_15906);
xor U16073 (N_16073,N_15840,N_15075);
nor U16074 (N_16074,N_15426,N_15346);
xor U16075 (N_16075,N_15232,N_15481);
or U16076 (N_16076,N_15573,N_15663);
nand U16077 (N_16077,N_15365,N_15042);
or U16078 (N_16078,N_15360,N_15849);
nand U16079 (N_16079,N_15351,N_15742);
and U16080 (N_16080,N_15966,N_15480);
and U16081 (N_16081,N_15288,N_15127);
and U16082 (N_16082,N_15052,N_15262);
or U16083 (N_16083,N_15281,N_15916);
or U16084 (N_16084,N_15805,N_15193);
and U16085 (N_16085,N_15006,N_15519);
nand U16086 (N_16086,N_15307,N_15703);
xor U16087 (N_16087,N_15995,N_15167);
xnor U16088 (N_16088,N_15170,N_15518);
nand U16089 (N_16089,N_15582,N_15148);
and U16090 (N_16090,N_15420,N_15154);
and U16091 (N_16091,N_15345,N_15969);
nand U16092 (N_16092,N_15562,N_15283);
or U16093 (N_16093,N_15873,N_15845);
xnor U16094 (N_16094,N_15851,N_15561);
or U16095 (N_16095,N_15433,N_15461);
xnor U16096 (N_16096,N_15238,N_15825);
nor U16097 (N_16097,N_15338,N_15874);
and U16098 (N_16098,N_15600,N_15306);
nand U16099 (N_16099,N_15653,N_15587);
nor U16100 (N_16100,N_15453,N_15199);
xor U16101 (N_16101,N_15063,N_15185);
nor U16102 (N_16102,N_15144,N_15918);
xnor U16103 (N_16103,N_15191,N_15254);
or U16104 (N_16104,N_15516,N_15878);
and U16105 (N_16105,N_15449,N_15614);
or U16106 (N_16106,N_15999,N_15413);
nand U16107 (N_16107,N_15000,N_15529);
xor U16108 (N_16108,N_15029,N_15359);
and U16109 (N_16109,N_15216,N_15778);
xor U16110 (N_16110,N_15865,N_15451);
xor U16111 (N_16111,N_15977,N_15541);
nor U16112 (N_16112,N_15383,N_15394);
nand U16113 (N_16113,N_15130,N_15140);
nor U16114 (N_16114,N_15869,N_15841);
and U16115 (N_16115,N_15563,N_15882);
or U16116 (N_16116,N_15733,N_15945);
or U16117 (N_16117,N_15682,N_15382);
or U16118 (N_16118,N_15026,N_15092);
nor U16119 (N_16119,N_15796,N_15558);
nor U16120 (N_16120,N_15914,N_15217);
nand U16121 (N_16121,N_15308,N_15903);
and U16122 (N_16122,N_15086,N_15755);
and U16123 (N_16123,N_15014,N_15340);
nor U16124 (N_16124,N_15454,N_15937);
or U16125 (N_16125,N_15375,N_15613);
and U16126 (N_16126,N_15058,N_15990);
or U16127 (N_16127,N_15609,N_15472);
nor U16128 (N_16128,N_15166,N_15743);
nand U16129 (N_16129,N_15819,N_15907);
nor U16130 (N_16130,N_15267,N_15673);
xnor U16131 (N_16131,N_15924,N_15169);
nand U16132 (N_16132,N_15651,N_15896);
xor U16133 (N_16133,N_15786,N_15446);
nand U16134 (N_16134,N_15429,N_15309);
and U16135 (N_16135,N_15671,N_15566);
xor U16136 (N_16136,N_15456,N_15737);
nand U16137 (N_16137,N_15899,N_15291);
xor U16138 (N_16138,N_15165,N_15669);
nand U16139 (N_16139,N_15220,N_15353);
nand U16140 (N_16140,N_15895,N_15103);
nor U16141 (N_16141,N_15303,N_15877);
or U16142 (N_16142,N_15114,N_15337);
or U16143 (N_16143,N_15719,N_15611);
xnor U16144 (N_16144,N_15102,N_15381);
nand U16145 (N_16145,N_15172,N_15527);
or U16146 (N_16146,N_15560,N_15387);
and U16147 (N_16147,N_15601,N_15003);
and U16148 (N_16148,N_15135,N_15946);
xnor U16149 (N_16149,N_15789,N_15004);
xnor U16150 (N_16150,N_15665,N_15368);
and U16151 (N_16151,N_15339,N_15156);
or U16152 (N_16152,N_15608,N_15829);
and U16153 (N_16153,N_15153,N_15547);
and U16154 (N_16154,N_15271,N_15521);
xnor U16155 (N_16155,N_15632,N_15593);
nor U16156 (N_16156,N_15280,N_15523);
nor U16157 (N_16157,N_15820,N_15675);
nand U16158 (N_16158,N_15589,N_15510);
xnor U16159 (N_16159,N_15396,N_15973);
or U16160 (N_16160,N_15577,N_15506);
and U16161 (N_16161,N_15022,N_15953);
and U16162 (N_16162,N_15304,N_15357);
and U16163 (N_16163,N_15385,N_15188);
nand U16164 (N_16164,N_15316,N_15751);
nor U16165 (N_16165,N_15943,N_15078);
xor U16166 (N_16166,N_15705,N_15934);
or U16167 (N_16167,N_15300,N_15362);
nor U16168 (N_16168,N_15777,N_15350);
and U16169 (N_16169,N_15010,N_15443);
xor U16170 (N_16170,N_15635,N_15823);
and U16171 (N_16171,N_15740,N_15599);
and U16172 (N_16172,N_15074,N_15576);
xor U16173 (N_16173,N_15859,N_15567);
nor U16174 (N_16174,N_15968,N_15211);
and U16175 (N_16175,N_15011,N_15181);
nor U16176 (N_16176,N_15866,N_15627);
nand U16177 (N_16177,N_15607,N_15157);
or U16178 (N_16178,N_15584,N_15715);
nand U16179 (N_16179,N_15575,N_15568);
nor U16180 (N_16180,N_15994,N_15347);
nor U16181 (N_16181,N_15783,N_15356);
nand U16182 (N_16182,N_15828,N_15019);
or U16183 (N_16183,N_15249,N_15597);
nand U16184 (N_16184,N_15469,N_15296);
or U16185 (N_16185,N_15424,N_15399);
nand U16186 (N_16186,N_15838,N_15512);
and U16187 (N_16187,N_15116,N_15248);
xnor U16188 (N_16188,N_15380,N_15222);
or U16189 (N_16189,N_15015,N_15400);
and U16190 (N_16190,N_15348,N_15932);
nor U16191 (N_16191,N_15009,N_15886);
or U16192 (N_16192,N_15298,N_15046);
or U16193 (N_16193,N_15730,N_15491);
or U16194 (N_16194,N_15626,N_15206);
or U16195 (N_16195,N_15414,N_15437);
or U16196 (N_16196,N_15077,N_15332);
nand U16197 (N_16197,N_15500,N_15284);
xnor U16198 (N_16198,N_15987,N_15780);
xnor U16199 (N_16199,N_15405,N_15770);
or U16200 (N_16200,N_15687,N_15571);
nand U16201 (N_16201,N_15126,N_15428);
or U16202 (N_16202,N_15128,N_15749);
nand U16203 (N_16203,N_15554,N_15556);
and U16204 (N_16204,N_15678,N_15268);
or U16205 (N_16205,N_15879,N_15962);
or U16206 (N_16206,N_15623,N_15120);
and U16207 (N_16207,N_15649,N_15091);
nor U16208 (N_16208,N_15302,N_15422);
nand U16209 (N_16209,N_15711,N_15605);
or U16210 (N_16210,N_15542,N_15311);
nor U16211 (N_16211,N_15894,N_15767);
and U16212 (N_16212,N_15096,N_15984);
xor U16213 (N_16213,N_15688,N_15548);
or U16214 (N_16214,N_15900,N_15646);
xor U16215 (N_16215,N_15629,N_15069);
nand U16216 (N_16216,N_15132,N_15479);
nand U16217 (N_16217,N_15694,N_15620);
nand U16218 (N_16218,N_15949,N_15490);
nor U16219 (N_16219,N_15328,N_15664);
and U16220 (N_16220,N_15905,N_15790);
and U16221 (N_16221,N_15318,N_15961);
or U16222 (N_16222,N_15320,N_15638);
and U16223 (N_16223,N_15731,N_15967);
or U16224 (N_16224,N_15138,N_15938);
or U16225 (N_16225,N_15274,N_15950);
and U16226 (N_16226,N_15979,N_15389);
xor U16227 (N_16227,N_15423,N_15177);
nand U16228 (N_16228,N_15955,N_15971);
nor U16229 (N_16229,N_15657,N_15020);
and U16230 (N_16230,N_15139,N_15223);
nor U16231 (N_16231,N_15197,N_15704);
xor U16232 (N_16232,N_15239,N_15243);
nor U16233 (N_16233,N_15788,N_15301);
xnor U16234 (N_16234,N_15923,N_15827);
and U16235 (N_16235,N_15794,N_15978);
nand U16236 (N_16236,N_15993,N_15225);
xnor U16237 (N_16237,N_15390,N_15848);
and U16238 (N_16238,N_15963,N_15501);
or U16239 (N_16239,N_15067,N_15942);
nand U16240 (N_16240,N_15929,N_15985);
or U16241 (N_16241,N_15373,N_15053);
nand U16242 (N_16242,N_15717,N_15691);
nor U16243 (N_16243,N_15549,N_15425);
xnor U16244 (N_16244,N_15628,N_15391);
nand U16245 (N_16245,N_15513,N_15049);
nor U16246 (N_16246,N_15958,N_15598);
nor U16247 (N_16247,N_15427,N_15313);
nor U16248 (N_16248,N_15989,N_15492);
and U16249 (N_16249,N_15692,N_15774);
or U16250 (N_16250,N_15781,N_15683);
nand U16251 (N_16251,N_15333,N_15964);
nand U16252 (N_16252,N_15707,N_15059);
nand U16253 (N_16253,N_15176,N_15459);
nor U16254 (N_16254,N_15363,N_15537);
nor U16255 (N_16255,N_15684,N_15106);
xnor U16256 (N_16256,N_15018,N_15213);
xnor U16257 (N_16257,N_15384,N_15118);
nand U16258 (N_16258,N_15037,N_15754);
xor U16259 (N_16259,N_15543,N_15113);
and U16260 (N_16260,N_15021,N_15245);
nand U16261 (N_16261,N_15230,N_15700);
nand U16262 (N_16262,N_15855,N_15214);
or U16263 (N_16263,N_15066,N_15530);
nand U16264 (N_16264,N_15898,N_15622);
or U16265 (N_16265,N_15094,N_15030);
nor U16266 (N_16266,N_15708,N_15064);
xnor U16267 (N_16267,N_15334,N_15137);
xor U16268 (N_16268,N_15444,N_15716);
nand U16269 (N_16269,N_15484,N_15411);
xor U16270 (N_16270,N_15095,N_15610);
and U16271 (N_16271,N_15555,N_15504);
nand U16272 (N_16272,N_15644,N_15386);
nand U16273 (N_16273,N_15395,N_15602);
nor U16274 (N_16274,N_15119,N_15606);
xor U16275 (N_16275,N_15641,N_15806);
and U16276 (N_16276,N_15361,N_15572);
or U16277 (N_16277,N_15834,N_15194);
and U16278 (N_16278,N_15473,N_15434);
and U16279 (N_16279,N_15041,N_15583);
and U16280 (N_16280,N_15528,N_15146);
xnor U16281 (N_16281,N_15410,N_15976);
or U16282 (N_16282,N_15335,N_15926);
and U16283 (N_16283,N_15911,N_15772);
nor U16284 (N_16284,N_15336,N_15902);
nor U16285 (N_16285,N_15493,N_15520);
and U16286 (N_16286,N_15044,N_15880);
xor U16287 (N_16287,N_15407,N_15738);
and U16288 (N_16288,N_15068,N_15412);
nor U16289 (N_16289,N_15761,N_15732);
or U16290 (N_16290,N_15912,N_15221);
nor U16291 (N_16291,N_15656,N_15081);
nor U16292 (N_16292,N_15775,N_15981);
nand U16293 (N_16293,N_15988,N_15464);
or U16294 (N_16294,N_15358,N_15325);
nand U16295 (N_16295,N_15585,N_15082);
xnor U16296 (N_16296,N_15639,N_15270);
or U16297 (N_16297,N_15901,N_15642);
or U16298 (N_16298,N_15084,N_15734);
or U16299 (N_16299,N_15637,N_15570);
nor U16300 (N_16300,N_15112,N_15025);
xor U16301 (N_16301,N_15970,N_15726);
nor U16302 (N_16302,N_15233,N_15785);
and U16303 (N_16303,N_15371,N_15676);
nand U16304 (N_16304,N_15007,N_15455);
or U16305 (N_16305,N_15545,N_15474);
nand U16306 (N_16306,N_15699,N_15850);
or U16307 (N_16307,N_15252,N_15447);
nor U16308 (N_16308,N_15494,N_15312);
and U16309 (N_16309,N_15388,N_15178);
or U16310 (N_16310,N_15122,N_15466);
nand U16311 (N_16311,N_15616,N_15723);
or U16312 (N_16312,N_15835,N_15766);
nor U16313 (N_16313,N_15940,N_15045);
nand U16314 (N_16314,N_15776,N_15847);
nand U16315 (N_16315,N_15888,N_15739);
nand U16316 (N_16316,N_15485,N_15809);
nand U16317 (N_16317,N_15764,N_15522);
and U16318 (N_16318,N_15080,N_15242);
nor U16319 (N_16319,N_15941,N_15398);
or U16320 (N_16320,N_15151,N_15160);
nand U16321 (N_16321,N_15867,N_15369);
or U16322 (N_16322,N_15769,N_15615);
xor U16323 (N_16323,N_15051,N_15784);
nor U16324 (N_16324,N_15860,N_15965);
and U16325 (N_16325,N_15310,N_15257);
xor U16326 (N_16326,N_15957,N_15324);
nor U16327 (N_16327,N_15246,N_15354);
and U16328 (N_16328,N_15710,N_15183);
xnor U16329 (N_16329,N_15782,N_15580);
xnor U16330 (N_16330,N_15210,N_15192);
and U16331 (N_16331,N_15709,N_15735);
nor U16332 (N_16332,N_15908,N_15565);
xor U16333 (N_16333,N_15229,N_15885);
nand U16334 (N_16334,N_15027,N_15815);
and U16335 (N_16335,N_15846,N_15736);
nand U16336 (N_16336,N_15952,N_15174);
and U16337 (N_16337,N_15787,N_15931);
xnor U16338 (N_16338,N_15921,N_15282);
and U16339 (N_16339,N_15706,N_15236);
or U16340 (N_16340,N_15633,N_15727);
nand U16341 (N_16341,N_15863,N_15034);
nand U16342 (N_16342,N_15793,N_15190);
and U16343 (N_16343,N_15564,N_15293);
or U16344 (N_16344,N_15645,N_15698);
nor U16345 (N_16345,N_15463,N_15925);
or U16346 (N_16346,N_15314,N_15370);
xor U16347 (N_16347,N_15974,N_15960);
and U16348 (N_16348,N_15648,N_15680);
nand U16349 (N_16349,N_15531,N_15525);
nand U16350 (N_16350,N_15551,N_15810);
or U16351 (N_16351,N_15795,N_15036);
xor U16352 (N_16352,N_15515,N_15591);
nor U16353 (N_16353,N_15757,N_15180);
nor U16354 (N_16354,N_15559,N_15647);
and U16355 (N_16355,N_15904,N_15812);
and U16356 (N_16356,N_15718,N_15035);
xor U16357 (N_16357,N_15868,N_15497);
or U16358 (N_16358,N_15871,N_15054);
nor U16359 (N_16359,N_15452,N_15643);
nor U16360 (N_16360,N_15145,N_15418);
nor U16361 (N_16361,N_15667,N_15076);
xnor U16362 (N_16362,N_15574,N_15822);
or U16363 (N_16363,N_15079,N_15685);
and U16364 (N_16364,N_15124,N_15364);
and U16365 (N_16365,N_15891,N_15234);
xnor U16366 (N_16366,N_15476,N_15640);
or U16367 (N_16367,N_15771,N_15276);
or U16368 (N_16368,N_15305,N_15269);
xnor U16369 (N_16369,N_15486,N_15171);
xor U16370 (N_16370,N_15259,N_15055);
nand U16371 (N_16371,N_15266,N_15071);
or U16372 (N_16372,N_15803,N_15768);
or U16373 (N_16373,N_15330,N_15275);
or U16374 (N_16374,N_15168,N_15430);
xnor U16375 (N_16375,N_15038,N_15884);
or U16376 (N_16376,N_15458,N_15219);
nand U16377 (N_16377,N_15817,N_15870);
or U16378 (N_16378,N_15198,N_15744);
and U16379 (N_16379,N_15517,N_15093);
or U16380 (N_16380,N_15801,N_15797);
nand U16381 (N_16381,N_15227,N_15109);
nand U16382 (N_16382,N_15256,N_15403);
nor U16383 (N_16383,N_15147,N_15612);
or U16384 (N_16384,N_15889,N_15617);
nor U16385 (N_16385,N_15125,N_15448);
nand U16386 (N_16386,N_15872,N_15179);
xnor U16387 (N_16387,N_15260,N_15721);
nor U16388 (N_16388,N_15445,N_15404);
nand U16389 (N_16389,N_15696,N_15047);
or U16390 (N_16390,N_15379,N_15750);
nand U16391 (N_16391,N_15944,N_15658);
and U16392 (N_16392,N_15247,N_15224);
xnor U16393 (N_16393,N_15465,N_15892);
and U16394 (N_16394,N_15023,N_15503);
nand U16395 (N_16395,N_15948,N_15436);
nor U16396 (N_16396,N_15005,N_15655);
nor U16397 (N_16397,N_15502,N_15861);
nor U16398 (N_16398,N_15186,N_15746);
xnor U16399 (N_16399,N_15251,N_15070);
nor U16400 (N_16400,N_15440,N_15725);
xnor U16401 (N_16401,N_15297,N_15295);
nand U16402 (N_16402,N_15341,N_15327);
xnor U16403 (N_16403,N_15630,N_15557);
nor U16404 (N_16404,N_15951,N_15342);
xnor U16405 (N_16405,N_15482,N_15495);
nand U16406 (N_16406,N_15837,N_15241);
xnor U16407 (N_16407,N_15579,N_15535);
or U16408 (N_16408,N_15668,N_15594);
or U16409 (N_16409,N_15747,N_15854);
nand U16410 (N_16410,N_15514,N_15155);
nand U16411 (N_16411,N_15378,N_15544);
and U16412 (N_16412,N_15883,N_15235);
nor U16413 (N_16413,N_15765,N_15661);
xnor U16414 (N_16414,N_15853,N_15240);
or U16415 (N_16415,N_15279,N_15202);
nor U16416 (N_16416,N_15507,N_15317);
and U16417 (N_16417,N_15636,N_15175);
nand U16418 (N_16418,N_15255,N_15935);
and U16419 (N_16419,N_15913,N_15409);
nor U16420 (N_16420,N_15804,N_15056);
nand U16421 (N_16421,N_15662,N_15833);
nand U16422 (N_16422,N_15569,N_15992);
nor U16423 (N_16423,N_15659,N_15876);
xnor U16424 (N_16424,N_15321,N_15108);
or U16425 (N_16425,N_15581,N_15265);
nand U16426 (N_16426,N_15110,N_15215);
or U16427 (N_16427,N_15376,N_15060);
and U16428 (N_16428,N_15909,N_15228);
and U16429 (N_16429,N_15477,N_15701);
or U16430 (N_16430,N_15072,N_15956);
and U16431 (N_16431,N_15253,N_15686);
or U16432 (N_16432,N_15697,N_15930);
or U16433 (N_16433,N_15802,N_15152);
and U16434 (N_16434,N_15331,N_15818);
or U16435 (N_16435,N_15182,N_15586);
xor U16436 (N_16436,N_15050,N_15712);
nand U16437 (N_16437,N_15928,N_15161);
nor U16438 (N_16438,N_15773,N_15619);
nor U16439 (N_16439,N_15634,N_15203);
nand U16440 (N_16440,N_15439,N_15762);
nand U16441 (N_16441,N_15674,N_15001);
nor U16442 (N_16442,N_15997,N_15807);
or U16443 (N_16443,N_15101,N_15831);
and U16444 (N_16444,N_15836,N_15457);
and U16445 (N_16445,N_15085,N_15511);
xor U16446 (N_16446,N_15273,N_15028);
and U16447 (N_16447,N_15524,N_15024);
and U16448 (N_16448,N_15496,N_15013);
and U16449 (N_16449,N_15666,N_15039);
nor U16450 (N_16450,N_15745,N_15419);
xnor U16451 (N_16451,N_15729,N_15690);
xor U16452 (N_16452,N_15821,N_15857);
nand U16453 (N_16453,N_15204,N_15462);
and U16454 (N_16454,N_15693,N_15299);
nor U16455 (N_16455,N_15349,N_15689);
xor U16456 (N_16456,N_15189,N_15982);
nor U16457 (N_16457,N_15031,N_15588);
and U16458 (N_16458,N_15856,N_15799);
nor U16459 (N_16459,N_15830,N_15752);
and U16460 (N_16460,N_15915,N_15292);
xnor U16461 (N_16461,N_15998,N_15129);
nand U16462 (N_16462,N_15722,N_15098);
nor U16463 (N_16463,N_15290,N_15534);
nor U16464 (N_16464,N_15142,N_15285);
nand U16465 (N_16465,N_15483,N_15713);
nor U16466 (N_16466,N_15226,N_15922);
or U16467 (N_16467,N_15864,N_15261);
and U16468 (N_16468,N_15272,N_15012);
nor U16469 (N_16469,N_15702,N_15763);
nand U16470 (N_16470,N_15088,N_15779);
nand U16471 (N_16471,N_15218,N_15816);
or U16472 (N_16472,N_15208,N_15631);
xor U16473 (N_16473,N_15212,N_15538);
nand U16474 (N_16474,N_15824,N_15947);
and U16475 (N_16475,N_15158,N_15143);
or U16476 (N_16476,N_15164,N_15843);
or U16477 (N_16477,N_15475,N_15237);
xor U16478 (N_16478,N_15832,N_15478);
xor U16479 (N_16479,N_15759,N_15792);
or U16480 (N_16480,N_15201,N_15526);
nor U16481 (N_16481,N_15090,N_15150);
nand U16482 (N_16482,N_15438,N_15289);
nor U16483 (N_16483,N_15991,N_15065);
and U16484 (N_16484,N_15278,N_15442);
or U16485 (N_16485,N_15724,N_15117);
xor U16486 (N_16486,N_15097,N_15467);
nand U16487 (N_16487,N_15505,N_15326);
nand U16488 (N_16488,N_15553,N_15933);
nand U16489 (N_16489,N_15163,N_15756);
and U16490 (N_16490,N_15954,N_15162);
or U16491 (N_16491,N_15996,N_15200);
xnor U16492 (N_16492,N_15498,N_15073);
and U16493 (N_16493,N_15972,N_15344);
nor U16494 (N_16494,N_15173,N_15624);
or U16495 (N_16495,N_15975,N_15367);
nand U16496 (N_16496,N_15959,N_15287);
xnor U16497 (N_16497,N_15131,N_15858);
nand U16498 (N_16498,N_15134,N_15315);
nor U16499 (N_16499,N_15939,N_15057);
nor U16500 (N_16500,N_15021,N_15510);
xnor U16501 (N_16501,N_15137,N_15381);
nor U16502 (N_16502,N_15620,N_15335);
nor U16503 (N_16503,N_15655,N_15457);
and U16504 (N_16504,N_15699,N_15501);
and U16505 (N_16505,N_15817,N_15872);
nand U16506 (N_16506,N_15020,N_15387);
or U16507 (N_16507,N_15052,N_15963);
or U16508 (N_16508,N_15314,N_15380);
or U16509 (N_16509,N_15283,N_15710);
nor U16510 (N_16510,N_15017,N_15798);
nand U16511 (N_16511,N_15157,N_15085);
or U16512 (N_16512,N_15896,N_15442);
and U16513 (N_16513,N_15707,N_15971);
or U16514 (N_16514,N_15570,N_15817);
and U16515 (N_16515,N_15426,N_15270);
xnor U16516 (N_16516,N_15725,N_15252);
xor U16517 (N_16517,N_15311,N_15704);
xor U16518 (N_16518,N_15130,N_15115);
xnor U16519 (N_16519,N_15111,N_15981);
or U16520 (N_16520,N_15278,N_15558);
nor U16521 (N_16521,N_15235,N_15964);
and U16522 (N_16522,N_15751,N_15710);
nand U16523 (N_16523,N_15280,N_15159);
nand U16524 (N_16524,N_15574,N_15041);
xor U16525 (N_16525,N_15524,N_15796);
and U16526 (N_16526,N_15494,N_15784);
nor U16527 (N_16527,N_15755,N_15239);
xor U16528 (N_16528,N_15700,N_15344);
nor U16529 (N_16529,N_15127,N_15149);
or U16530 (N_16530,N_15946,N_15136);
nor U16531 (N_16531,N_15147,N_15902);
and U16532 (N_16532,N_15018,N_15737);
and U16533 (N_16533,N_15495,N_15679);
xor U16534 (N_16534,N_15422,N_15038);
and U16535 (N_16535,N_15578,N_15065);
nor U16536 (N_16536,N_15423,N_15430);
or U16537 (N_16537,N_15261,N_15536);
or U16538 (N_16538,N_15270,N_15305);
or U16539 (N_16539,N_15610,N_15391);
nor U16540 (N_16540,N_15861,N_15826);
xnor U16541 (N_16541,N_15717,N_15095);
nand U16542 (N_16542,N_15075,N_15662);
and U16543 (N_16543,N_15022,N_15393);
nor U16544 (N_16544,N_15859,N_15847);
nor U16545 (N_16545,N_15013,N_15202);
nand U16546 (N_16546,N_15750,N_15002);
and U16547 (N_16547,N_15952,N_15505);
xnor U16548 (N_16548,N_15474,N_15571);
xnor U16549 (N_16549,N_15797,N_15540);
or U16550 (N_16550,N_15341,N_15515);
nor U16551 (N_16551,N_15751,N_15813);
and U16552 (N_16552,N_15850,N_15440);
nor U16553 (N_16553,N_15019,N_15129);
or U16554 (N_16554,N_15023,N_15958);
xor U16555 (N_16555,N_15328,N_15748);
and U16556 (N_16556,N_15255,N_15627);
and U16557 (N_16557,N_15679,N_15951);
or U16558 (N_16558,N_15120,N_15129);
or U16559 (N_16559,N_15564,N_15558);
or U16560 (N_16560,N_15861,N_15026);
nor U16561 (N_16561,N_15490,N_15299);
xnor U16562 (N_16562,N_15536,N_15984);
nand U16563 (N_16563,N_15689,N_15432);
nor U16564 (N_16564,N_15409,N_15627);
xor U16565 (N_16565,N_15433,N_15665);
xor U16566 (N_16566,N_15514,N_15575);
or U16567 (N_16567,N_15417,N_15713);
and U16568 (N_16568,N_15420,N_15809);
nor U16569 (N_16569,N_15167,N_15375);
or U16570 (N_16570,N_15139,N_15731);
and U16571 (N_16571,N_15265,N_15816);
nand U16572 (N_16572,N_15774,N_15695);
nor U16573 (N_16573,N_15484,N_15850);
xnor U16574 (N_16574,N_15204,N_15807);
nor U16575 (N_16575,N_15656,N_15624);
nand U16576 (N_16576,N_15553,N_15845);
nand U16577 (N_16577,N_15978,N_15631);
or U16578 (N_16578,N_15652,N_15659);
xnor U16579 (N_16579,N_15294,N_15241);
and U16580 (N_16580,N_15421,N_15366);
or U16581 (N_16581,N_15859,N_15290);
and U16582 (N_16582,N_15650,N_15197);
nor U16583 (N_16583,N_15685,N_15141);
and U16584 (N_16584,N_15549,N_15357);
or U16585 (N_16585,N_15712,N_15804);
and U16586 (N_16586,N_15518,N_15602);
or U16587 (N_16587,N_15439,N_15446);
nand U16588 (N_16588,N_15298,N_15189);
and U16589 (N_16589,N_15648,N_15306);
nor U16590 (N_16590,N_15811,N_15955);
or U16591 (N_16591,N_15842,N_15896);
or U16592 (N_16592,N_15201,N_15194);
and U16593 (N_16593,N_15200,N_15537);
xnor U16594 (N_16594,N_15245,N_15285);
xor U16595 (N_16595,N_15074,N_15202);
and U16596 (N_16596,N_15201,N_15861);
xor U16597 (N_16597,N_15583,N_15161);
or U16598 (N_16598,N_15635,N_15455);
nor U16599 (N_16599,N_15507,N_15803);
or U16600 (N_16600,N_15291,N_15912);
or U16601 (N_16601,N_15521,N_15252);
xor U16602 (N_16602,N_15710,N_15967);
xor U16603 (N_16603,N_15286,N_15085);
or U16604 (N_16604,N_15336,N_15318);
xnor U16605 (N_16605,N_15033,N_15405);
or U16606 (N_16606,N_15773,N_15205);
nand U16607 (N_16607,N_15676,N_15966);
or U16608 (N_16608,N_15518,N_15669);
xnor U16609 (N_16609,N_15229,N_15681);
and U16610 (N_16610,N_15114,N_15409);
nand U16611 (N_16611,N_15155,N_15890);
xor U16612 (N_16612,N_15860,N_15872);
nor U16613 (N_16613,N_15047,N_15814);
nor U16614 (N_16614,N_15449,N_15099);
nor U16615 (N_16615,N_15299,N_15990);
xnor U16616 (N_16616,N_15259,N_15177);
or U16617 (N_16617,N_15356,N_15653);
and U16618 (N_16618,N_15587,N_15456);
or U16619 (N_16619,N_15406,N_15958);
nand U16620 (N_16620,N_15299,N_15621);
nand U16621 (N_16621,N_15687,N_15394);
and U16622 (N_16622,N_15780,N_15994);
xnor U16623 (N_16623,N_15187,N_15046);
nor U16624 (N_16624,N_15372,N_15312);
or U16625 (N_16625,N_15637,N_15217);
or U16626 (N_16626,N_15175,N_15614);
nand U16627 (N_16627,N_15251,N_15185);
nand U16628 (N_16628,N_15075,N_15210);
nor U16629 (N_16629,N_15677,N_15557);
nor U16630 (N_16630,N_15078,N_15106);
or U16631 (N_16631,N_15395,N_15648);
nand U16632 (N_16632,N_15397,N_15582);
nor U16633 (N_16633,N_15313,N_15019);
or U16634 (N_16634,N_15688,N_15582);
or U16635 (N_16635,N_15167,N_15416);
and U16636 (N_16636,N_15228,N_15453);
xor U16637 (N_16637,N_15675,N_15940);
nor U16638 (N_16638,N_15556,N_15474);
or U16639 (N_16639,N_15253,N_15734);
xor U16640 (N_16640,N_15826,N_15621);
xnor U16641 (N_16641,N_15473,N_15819);
nor U16642 (N_16642,N_15472,N_15219);
or U16643 (N_16643,N_15733,N_15149);
xor U16644 (N_16644,N_15700,N_15812);
xor U16645 (N_16645,N_15805,N_15512);
nand U16646 (N_16646,N_15883,N_15663);
or U16647 (N_16647,N_15456,N_15324);
or U16648 (N_16648,N_15661,N_15050);
and U16649 (N_16649,N_15029,N_15537);
nor U16650 (N_16650,N_15307,N_15451);
or U16651 (N_16651,N_15765,N_15154);
nor U16652 (N_16652,N_15074,N_15272);
nor U16653 (N_16653,N_15737,N_15483);
and U16654 (N_16654,N_15550,N_15809);
and U16655 (N_16655,N_15111,N_15227);
and U16656 (N_16656,N_15485,N_15004);
and U16657 (N_16657,N_15187,N_15145);
nand U16658 (N_16658,N_15945,N_15285);
or U16659 (N_16659,N_15564,N_15010);
and U16660 (N_16660,N_15362,N_15863);
xnor U16661 (N_16661,N_15621,N_15786);
nand U16662 (N_16662,N_15597,N_15822);
and U16663 (N_16663,N_15492,N_15223);
nand U16664 (N_16664,N_15701,N_15655);
xnor U16665 (N_16665,N_15698,N_15863);
and U16666 (N_16666,N_15836,N_15557);
or U16667 (N_16667,N_15039,N_15714);
or U16668 (N_16668,N_15539,N_15070);
nor U16669 (N_16669,N_15675,N_15988);
or U16670 (N_16670,N_15246,N_15969);
and U16671 (N_16671,N_15754,N_15237);
nand U16672 (N_16672,N_15538,N_15342);
nor U16673 (N_16673,N_15378,N_15614);
nand U16674 (N_16674,N_15022,N_15843);
and U16675 (N_16675,N_15824,N_15225);
and U16676 (N_16676,N_15766,N_15990);
nor U16677 (N_16677,N_15388,N_15529);
nand U16678 (N_16678,N_15724,N_15162);
and U16679 (N_16679,N_15724,N_15375);
xor U16680 (N_16680,N_15617,N_15098);
xor U16681 (N_16681,N_15093,N_15499);
and U16682 (N_16682,N_15503,N_15215);
nor U16683 (N_16683,N_15625,N_15447);
nand U16684 (N_16684,N_15409,N_15064);
and U16685 (N_16685,N_15175,N_15514);
or U16686 (N_16686,N_15636,N_15050);
or U16687 (N_16687,N_15227,N_15741);
nor U16688 (N_16688,N_15147,N_15171);
or U16689 (N_16689,N_15135,N_15348);
nor U16690 (N_16690,N_15470,N_15261);
nor U16691 (N_16691,N_15117,N_15328);
and U16692 (N_16692,N_15835,N_15728);
nor U16693 (N_16693,N_15245,N_15609);
nor U16694 (N_16694,N_15946,N_15316);
and U16695 (N_16695,N_15545,N_15986);
or U16696 (N_16696,N_15472,N_15923);
or U16697 (N_16697,N_15360,N_15757);
and U16698 (N_16698,N_15573,N_15265);
xor U16699 (N_16699,N_15525,N_15694);
and U16700 (N_16700,N_15660,N_15002);
nor U16701 (N_16701,N_15074,N_15332);
nand U16702 (N_16702,N_15219,N_15778);
and U16703 (N_16703,N_15541,N_15575);
or U16704 (N_16704,N_15152,N_15718);
nand U16705 (N_16705,N_15281,N_15141);
nand U16706 (N_16706,N_15881,N_15171);
or U16707 (N_16707,N_15223,N_15192);
nor U16708 (N_16708,N_15659,N_15358);
xnor U16709 (N_16709,N_15718,N_15142);
nor U16710 (N_16710,N_15274,N_15990);
nor U16711 (N_16711,N_15239,N_15365);
xnor U16712 (N_16712,N_15435,N_15515);
nor U16713 (N_16713,N_15832,N_15366);
nor U16714 (N_16714,N_15061,N_15211);
nor U16715 (N_16715,N_15079,N_15473);
and U16716 (N_16716,N_15476,N_15709);
xnor U16717 (N_16717,N_15872,N_15905);
nor U16718 (N_16718,N_15788,N_15364);
xor U16719 (N_16719,N_15452,N_15458);
nor U16720 (N_16720,N_15295,N_15316);
and U16721 (N_16721,N_15490,N_15784);
or U16722 (N_16722,N_15383,N_15145);
xnor U16723 (N_16723,N_15862,N_15056);
nand U16724 (N_16724,N_15651,N_15738);
xnor U16725 (N_16725,N_15140,N_15664);
or U16726 (N_16726,N_15403,N_15013);
nand U16727 (N_16727,N_15681,N_15748);
or U16728 (N_16728,N_15494,N_15276);
nor U16729 (N_16729,N_15001,N_15468);
nor U16730 (N_16730,N_15676,N_15688);
xnor U16731 (N_16731,N_15663,N_15014);
or U16732 (N_16732,N_15099,N_15306);
xnor U16733 (N_16733,N_15638,N_15411);
and U16734 (N_16734,N_15859,N_15564);
nor U16735 (N_16735,N_15662,N_15529);
xor U16736 (N_16736,N_15106,N_15745);
nand U16737 (N_16737,N_15042,N_15390);
nor U16738 (N_16738,N_15258,N_15668);
nand U16739 (N_16739,N_15867,N_15332);
and U16740 (N_16740,N_15015,N_15882);
xor U16741 (N_16741,N_15967,N_15356);
nor U16742 (N_16742,N_15626,N_15245);
nand U16743 (N_16743,N_15217,N_15510);
nand U16744 (N_16744,N_15787,N_15412);
nor U16745 (N_16745,N_15575,N_15516);
or U16746 (N_16746,N_15055,N_15607);
nor U16747 (N_16747,N_15112,N_15407);
nand U16748 (N_16748,N_15407,N_15477);
nor U16749 (N_16749,N_15462,N_15881);
xor U16750 (N_16750,N_15902,N_15864);
nand U16751 (N_16751,N_15000,N_15205);
nor U16752 (N_16752,N_15548,N_15433);
nand U16753 (N_16753,N_15425,N_15052);
xnor U16754 (N_16754,N_15502,N_15972);
nor U16755 (N_16755,N_15211,N_15489);
xnor U16756 (N_16756,N_15157,N_15987);
nand U16757 (N_16757,N_15561,N_15231);
or U16758 (N_16758,N_15447,N_15710);
nand U16759 (N_16759,N_15171,N_15391);
nor U16760 (N_16760,N_15618,N_15667);
and U16761 (N_16761,N_15363,N_15121);
nor U16762 (N_16762,N_15728,N_15102);
or U16763 (N_16763,N_15774,N_15167);
xor U16764 (N_16764,N_15334,N_15839);
nor U16765 (N_16765,N_15238,N_15532);
and U16766 (N_16766,N_15469,N_15581);
nor U16767 (N_16767,N_15424,N_15477);
nor U16768 (N_16768,N_15279,N_15334);
nor U16769 (N_16769,N_15836,N_15089);
or U16770 (N_16770,N_15051,N_15701);
nor U16771 (N_16771,N_15273,N_15158);
nand U16772 (N_16772,N_15778,N_15092);
nor U16773 (N_16773,N_15794,N_15158);
or U16774 (N_16774,N_15452,N_15719);
and U16775 (N_16775,N_15300,N_15094);
or U16776 (N_16776,N_15587,N_15123);
nor U16777 (N_16777,N_15192,N_15354);
xor U16778 (N_16778,N_15095,N_15831);
or U16779 (N_16779,N_15175,N_15441);
nand U16780 (N_16780,N_15378,N_15428);
or U16781 (N_16781,N_15396,N_15787);
xor U16782 (N_16782,N_15345,N_15455);
and U16783 (N_16783,N_15507,N_15702);
or U16784 (N_16784,N_15180,N_15080);
xor U16785 (N_16785,N_15386,N_15443);
nor U16786 (N_16786,N_15958,N_15765);
and U16787 (N_16787,N_15741,N_15179);
nand U16788 (N_16788,N_15001,N_15389);
xnor U16789 (N_16789,N_15095,N_15660);
or U16790 (N_16790,N_15944,N_15568);
nand U16791 (N_16791,N_15199,N_15539);
and U16792 (N_16792,N_15357,N_15873);
and U16793 (N_16793,N_15661,N_15666);
and U16794 (N_16794,N_15862,N_15388);
or U16795 (N_16795,N_15441,N_15923);
nor U16796 (N_16796,N_15238,N_15289);
nor U16797 (N_16797,N_15692,N_15277);
and U16798 (N_16798,N_15389,N_15568);
xnor U16799 (N_16799,N_15341,N_15633);
and U16800 (N_16800,N_15223,N_15630);
xor U16801 (N_16801,N_15766,N_15219);
nand U16802 (N_16802,N_15784,N_15748);
nand U16803 (N_16803,N_15016,N_15828);
nand U16804 (N_16804,N_15794,N_15257);
and U16805 (N_16805,N_15641,N_15003);
nand U16806 (N_16806,N_15647,N_15898);
nand U16807 (N_16807,N_15531,N_15564);
and U16808 (N_16808,N_15209,N_15869);
nand U16809 (N_16809,N_15789,N_15785);
or U16810 (N_16810,N_15564,N_15831);
nand U16811 (N_16811,N_15504,N_15921);
and U16812 (N_16812,N_15966,N_15164);
or U16813 (N_16813,N_15116,N_15207);
or U16814 (N_16814,N_15922,N_15713);
xnor U16815 (N_16815,N_15925,N_15025);
and U16816 (N_16816,N_15671,N_15894);
nor U16817 (N_16817,N_15403,N_15550);
or U16818 (N_16818,N_15706,N_15158);
nand U16819 (N_16819,N_15802,N_15121);
xnor U16820 (N_16820,N_15870,N_15044);
and U16821 (N_16821,N_15114,N_15295);
nor U16822 (N_16822,N_15260,N_15628);
and U16823 (N_16823,N_15391,N_15780);
or U16824 (N_16824,N_15269,N_15103);
nand U16825 (N_16825,N_15671,N_15722);
or U16826 (N_16826,N_15734,N_15539);
or U16827 (N_16827,N_15711,N_15806);
and U16828 (N_16828,N_15011,N_15807);
nor U16829 (N_16829,N_15184,N_15198);
nor U16830 (N_16830,N_15042,N_15470);
nor U16831 (N_16831,N_15292,N_15083);
nand U16832 (N_16832,N_15607,N_15392);
and U16833 (N_16833,N_15135,N_15858);
xnor U16834 (N_16834,N_15074,N_15556);
xnor U16835 (N_16835,N_15188,N_15068);
xnor U16836 (N_16836,N_15555,N_15747);
nor U16837 (N_16837,N_15823,N_15255);
or U16838 (N_16838,N_15773,N_15973);
or U16839 (N_16839,N_15234,N_15223);
and U16840 (N_16840,N_15896,N_15499);
nor U16841 (N_16841,N_15068,N_15562);
xnor U16842 (N_16842,N_15526,N_15752);
or U16843 (N_16843,N_15498,N_15521);
nand U16844 (N_16844,N_15791,N_15178);
or U16845 (N_16845,N_15410,N_15025);
nor U16846 (N_16846,N_15978,N_15840);
nor U16847 (N_16847,N_15131,N_15537);
nand U16848 (N_16848,N_15350,N_15461);
nor U16849 (N_16849,N_15115,N_15741);
nand U16850 (N_16850,N_15857,N_15279);
nor U16851 (N_16851,N_15046,N_15022);
nor U16852 (N_16852,N_15574,N_15807);
xor U16853 (N_16853,N_15214,N_15063);
xor U16854 (N_16854,N_15291,N_15865);
nor U16855 (N_16855,N_15575,N_15580);
xnor U16856 (N_16856,N_15865,N_15723);
xnor U16857 (N_16857,N_15311,N_15587);
or U16858 (N_16858,N_15520,N_15629);
nand U16859 (N_16859,N_15663,N_15980);
nand U16860 (N_16860,N_15154,N_15995);
nor U16861 (N_16861,N_15389,N_15749);
and U16862 (N_16862,N_15587,N_15818);
or U16863 (N_16863,N_15230,N_15696);
or U16864 (N_16864,N_15831,N_15038);
nand U16865 (N_16865,N_15022,N_15344);
xor U16866 (N_16866,N_15226,N_15527);
xor U16867 (N_16867,N_15238,N_15072);
xor U16868 (N_16868,N_15324,N_15453);
and U16869 (N_16869,N_15638,N_15327);
xnor U16870 (N_16870,N_15964,N_15827);
nand U16871 (N_16871,N_15954,N_15631);
nand U16872 (N_16872,N_15050,N_15167);
and U16873 (N_16873,N_15700,N_15134);
or U16874 (N_16874,N_15061,N_15380);
nor U16875 (N_16875,N_15889,N_15822);
nor U16876 (N_16876,N_15512,N_15545);
or U16877 (N_16877,N_15869,N_15105);
and U16878 (N_16878,N_15040,N_15656);
and U16879 (N_16879,N_15718,N_15432);
nor U16880 (N_16880,N_15494,N_15502);
nand U16881 (N_16881,N_15516,N_15378);
or U16882 (N_16882,N_15578,N_15178);
xnor U16883 (N_16883,N_15864,N_15921);
or U16884 (N_16884,N_15540,N_15519);
nor U16885 (N_16885,N_15419,N_15004);
and U16886 (N_16886,N_15803,N_15271);
and U16887 (N_16887,N_15373,N_15461);
and U16888 (N_16888,N_15326,N_15759);
nand U16889 (N_16889,N_15211,N_15729);
nand U16890 (N_16890,N_15126,N_15338);
nor U16891 (N_16891,N_15635,N_15459);
and U16892 (N_16892,N_15182,N_15602);
nand U16893 (N_16893,N_15314,N_15323);
nand U16894 (N_16894,N_15534,N_15609);
and U16895 (N_16895,N_15908,N_15650);
or U16896 (N_16896,N_15545,N_15802);
and U16897 (N_16897,N_15017,N_15331);
and U16898 (N_16898,N_15550,N_15979);
xnor U16899 (N_16899,N_15454,N_15585);
nor U16900 (N_16900,N_15759,N_15227);
or U16901 (N_16901,N_15626,N_15496);
xnor U16902 (N_16902,N_15204,N_15878);
or U16903 (N_16903,N_15918,N_15756);
and U16904 (N_16904,N_15386,N_15303);
xnor U16905 (N_16905,N_15931,N_15649);
and U16906 (N_16906,N_15078,N_15691);
nand U16907 (N_16907,N_15092,N_15949);
xnor U16908 (N_16908,N_15010,N_15053);
xor U16909 (N_16909,N_15795,N_15522);
nand U16910 (N_16910,N_15828,N_15224);
nand U16911 (N_16911,N_15882,N_15782);
nor U16912 (N_16912,N_15999,N_15861);
or U16913 (N_16913,N_15955,N_15617);
xnor U16914 (N_16914,N_15966,N_15256);
nor U16915 (N_16915,N_15148,N_15634);
and U16916 (N_16916,N_15539,N_15389);
nor U16917 (N_16917,N_15543,N_15841);
xnor U16918 (N_16918,N_15368,N_15158);
and U16919 (N_16919,N_15760,N_15244);
and U16920 (N_16920,N_15545,N_15580);
and U16921 (N_16921,N_15924,N_15552);
and U16922 (N_16922,N_15263,N_15304);
nand U16923 (N_16923,N_15561,N_15075);
and U16924 (N_16924,N_15013,N_15551);
xnor U16925 (N_16925,N_15044,N_15320);
nand U16926 (N_16926,N_15061,N_15397);
xor U16927 (N_16927,N_15303,N_15590);
nor U16928 (N_16928,N_15102,N_15346);
or U16929 (N_16929,N_15295,N_15739);
xor U16930 (N_16930,N_15001,N_15568);
nor U16931 (N_16931,N_15367,N_15069);
and U16932 (N_16932,N_15839,N_15335);
nor U16933 (N_16933,N_15963,N_15153);
nor U16934 (N_16934,N_15933,N_15673);
nor U16935 (N_16935,N_15879,N_15432);
and U16936 (N_16936,N_15182,N_15517);
and U16937 (N_16937,N_15204,N_15783);
nand U16938 (N_16938,N_15147,N_15627);
and U16939 (N_16939,N_15111,N_15213);
nand U16940 (N_16940,N_15293,N_15287);
nand U16941 (N_16941,N_15849,N_15931);
nor U16942 (N_16942,N_15021,N_15374);
and U16943 (N_16943,N_15584,N_15652);
xnor U16944 (N_16944,N_15970,N_15867);
or U16945 (N_16945,N_15500,N_15307);
nor U16946 (N_16946,N_15368,N_15610);
nand U16947 (N_16947,N_15555,N_15607);
nand U16948 (N_16948,N_15089,N_15062);
xor U16949 (N_16949,N_15750,N_15092);
and U16950 (N_16950,N_15340,N_15424);
or U16951 (N_16951,N_15958,N_15669);
and U16952 (N_16952,N_15433,N_15222);
or U16953 (N_16953,N_15463,N_15764);
nor U16954 (N_16954,N_15068,N_15482);
nor U16955 (N_16955,N_15999,N_15432);
nand U16956 (N_16956,N_15391,N_15179);
xor U16957 (N_16957,N_15413,N_15012);
and U16958 (N_16958,N_15875,N_15649);
and U16959 (N_16959,N_15253,N_15318);
nand U16960 (N_16960,N_15677,N_15426);
nand U16961 (N_16961,N_15481,N_15367);
and U16962 (N_16962,N_15884,N_15796);
and U16963 (N_16963,N_15032,N_15308);
nand U16964 (N_16964,N_15806,N_15938);
nor U16965 (N_16965,N_15314,N_15429);
xnor U16966 (N_16966,N_15515,N_15562);
nand U16967 (N_16967,N_15387,N_15338);
and U16968 (N_16968,N_15791,N_15471);
or U16969 (N_16969,N_15497,N_15199);
nor U16970 (N_16970,N_15111,N_15401);
or U16971 (N_16971,N_15371,N_15895);
and U16972 (N_16972,N_15992,N_15639);
nor U16973 (N_16973,N_15449,N_15299);
or U16974 (N_16974,N_15805,N_15188);
xor U16975 (N_16975,N_15118,N_15075);
xnor U16976 (N_16976,N_15776,N_15465);
or U16977 (N_16977,N_15613,N_15015);
xnor U16978 (N_16978,N_15041,N_15095);
or U16979 (N_16979,N_15798,N_15313);
nand U16980 (N_16980,N_15085,N_15397);
nand U16981 (N_16981,N_15966,N_15149);
and U16982 (N_16982,N_15265,N_15701);
and U16983 (N_16983,N_15417,N_15045);
or U16984 (N_16984,N_15894,N_15059);
xor U16985 (N_16985,N_15439,N_15258);
nand U16986 (N_16986,N_15296,N_15935);
nor U16987 (N_16987,N_15382,N_15361);
and U16988 (N_16988,N_15175,N_15201);
xor U16989 (N_16989,N_15240,N_15696);
nor U16990 (N_16990,N_15017,N_15834);
xor U16991 (N_16991,N_15048,N_15269);
nor U16992 (N_16992,N_15771,N_15776);
xor U16993 (N_16993,N_15806,N_15947);
and U16994 (N_16994,N_15147,N_15504);
xor U16995 (N_16995,N_15670,N_15328);
nor U16996 (N_16996,N_15520,N_15835);
or U16997 (N_16997,N_15996,N_15520);
and U16998 (N_16998,N_15686,N_15534);
and U16999 (N_16999,N_15383,N_15741);
nor U17000 (N_17000,N_16524,N_16089);
and U17001 (N_17001,N_16355,N_16767);
or U17002 (N_17002,N_16803,N_16742);
xnor U17003 (N_17003,N_16563,N_16979);
nand U17004 (N_17004,N_16005,N_16148);
nor U17005 (N_17005,N_16158,N_16987);
nor U17006 (N_17006,N_16991,N_16079);
xnor U17007 (N_17007,N_16077,N_16608);
and U17008 (N_17008,N_16229,N_16707);
nand U17009 (N_17009,N_16811,N_16364);
or U17010 (N_17010,N_16942,N_16051);
and U17011 (N_17011,N_16974,N_16163);
nor U17012 (N_17012,N_16497,N_16625);
or U17013 (N_17013,N_16753,N_16778);
or U17014 (N_17014,N_16142,N_16698);
and U17015 (N_17015,N_16349,N_16495);
nand U17016 (N_17016,N_16144,N_16078);
or U17017 (N_17017,N_16130,N_16779);
nor U17018 (N_17018,N_16222,N_16116);
xor U17019 (N_17019,N_16413,N_16145);
or U17020 (N_17020,N_16690,N_16387);
xor U17021 (N_17021,N_16194,N_16240);
xor U17022 (N_17022,N_16289,N_16352);
nand U17023 (N_17023,N_16214,N_16797);
or U17024 (N_17024,N_16265,N_16575);
or U17025 (N_17025,N_16584,N_16916);
and U17026 (N_17026,N_16607,N_16958);
xnor U17027 (N_17027,N_16191,N_16307);
or U17028 (N_17028,N_16316,N_16684);
nand U17029 (N_17029,N_16446,N_16800);
or U17030 (N_17030,N_16111,N_16311);
nand U17031 (N_17031,N_16697,N_16863);
xor U17032 (N_17032,N_16469,N_16131);
nand U17033 (N_17033,N_16490,N_16843);
nor U17034 (N_17034,N_16065,N_16948);
nor U17035 (N_17035,N_16225,N_16000);
nor U17036 (N_17036,N_16838,N_16712);
or U17037 (N_17037,N_16616,N_16795);
and U17038 (N_17038,N_16489,N_16199);
nand U17039 (N_17039,N_16571,N_16187);
nor U17040 (N_17040,N_16162,N_16688);
and U17041 (N_17041,N_16190,N_16211);
or U17042 (N_17042,N_16872,N_16132);
and U17043 (N_17043,N_16248,N_16787);
and U17044 (N_17044,N_16873,N_16754);
and U17045 (N_17045,N_16867,N_16839);
xor U17046 (N_17046,N_16444,N_16724);
nand U17047 (N_17047,N_16705,N_16911);
and U17048 (N_17048,N_16353,N_16431);
and U17049 (N_17049,N_16726,N_16391);
xnor U17050 (N_17050,N_16023,N_16700);
xor U17051 (N_17051,N_16953,N_16909);
or U17052 (N_17052,N_16224,N_16756);
nand U17053 (N_17053,N_16592,N_16128);
nor U17054 (N_17054,N_16852,N_16418);
or U17055 (N_17055,N_16792,N_16473);
or U17056 (N_17056,N_16530,N_16717);
and U17057 (N_17057,N_16918,N_16420);
nor U17058 (N_17058,N_16580,N_16462);
xor U17059 (N_17059,N_16663,N_16071);
or U17060 (N_17060,N_16458,N_16732);
xor U17061 (N_17061,N_16317,N_16041);
nor U17062 (N_17062,N_16939,N_16959);
nor U17063 (N_17063,N_16526,N_16227);
nand U17064 (N_17064,N_16842,N_16376);
nor U17065 (N_17065,N_16814,N_16239);
xor U17066 (N_17066,N_16955,N_16403);
nand U17067 (N_17067,N_16161,N_16525);
nand U17068 (N_17068,N_16609,N_16100);
or U17069 (N_17069,N_16416,N_16703);
xor U17070 (N_17070,N_16244,N_16306);
or U17071 (N_17071,N_16003,N_16113);
xnor U17072 (N_17072,N_16310,N_16589);
nand U17073 (N_17073,N_16174,N_16505);
nand U17074 (N_17074,N_16183,N_16381);
nor U17075 (N_17075,N_16831,N_16739);
nor U17076 (N_17076,N_16092,N_16247);
xor U17077 (N_17077,N_16196,N_16840);
or U17078 (N_17078,N_16876,N_16421);
nand U17079 (N_17079,N_16500,N_16336);
and U17080 (N_17080,N_16451,N_16629);
and U17081 (N_17081,N_16232,N_16817);
or U17082 (N_17082,N_16658,N_16371);
xnor U17083 (N_17083,N_16396,N_16321);
and U17084 (N_17084,N_16836,N_16338);
or U17085 (N_17085,N_16457,N_16896);
or U17086 (N_17086,N_16520,N_16279);
and U17087 (N_17087,N_16195,N_16346);
xor U17088 (N_17088,N_16819,N_16258);
nand U17089 (N_17089,N_16521,N_16374);
xor U17090 (N_17090,N_16782,N_16885);
and U17091 (N_17091,N_16203,N_16708);
or U17092 (N_17092,N_16822,N_16606);
nor U17093 (N_17093,N_16056,N_16670);
nand U17094 (N_17094,N_16808,N_16752);
nor U17095 (N_17095,N_16015,N_16082);
nand U17096 (N_17096,N_16004,N_16859);
nor U17097 (N_17097,N_16487,N_16680);
nor U17098 (N_17098,N_16133,N_16509);
or U17099 (N_17099,N_16108,N_16660);
nand U17100 (N_17100,N_16780,N_16043);
nor U17101 (N_17101,N_16242,N_16682);
or U17102 (N_17102,N_16810,N_16542);
or U17103 (N_17103,N_16491,N_16883);
nor U17104 (N_17104,N_16411,N_16801);
xor U17105 (N_17105,N_16764,N_16377);
and U17106 (N_17106,N_16408,N_16280);
or U17107 (N_17107,N_16315,N_16300);
xor U17108 (N_17108,N_16642,N_16611);
nor U17109 (N_17109,N_16328,N_16880);
xnor U17110 (N_17110,N_16012,N_16590);
or U17111 (N_17111,N_16140,N_16188);
nand U17112 (N_17112,N_16501,N_16298);
nand U17113 (N_17113,N_16744,N_16454);
or U17114 (N_17114,N_16647,N_16437);
nand U17115 (N_17115,N_16850,N_16983);
and U17116 (N_17116,N_16922,N_16054);
nor U17117 (N_17117,N_16910,N_16478);
xor U17118 (N_17118,N_16231,N_16498);
and U17119 (N_17119,N_16168,N_16924);
xnor U17120 (N_17120,N_16110,N_16706);
nand U17121 (N_17121,N_16479,N_16746);
or U17122 (N_17122,N_16933,N_16519);
nand U17123 (N_17123,N_16292,N_16516);
and U17124 (N_17124,N_16952,N_16855);
xnor U17125 (N_17125,N_16114,N_16623);
xnor U17126 (N_17126,N_16721,N_16370);
or U17127 (N_17127,N_16155,N_16638);
xnor U17128 (N_17128,N_16996,N_16379);
or U17129 (N_17129,N_16655,N_16157);
or U17130 (N_17130,N_16704,N_16973);
and U17131 (N_17131,N_16159,N_16686);
nand U17132 (N_17132,N_16319,N_16126);
nand U17133 (N_17133,N_16044,N_16031);
xor U17134 (N_17134,N_16599,N_16978);
xnor U17135 (N_17135,N_16105,N_16776);
xnor U17136 (N_17136,N_16601,N_16136);
nor U17137 (N_17137,N_16790,N_16785);
and U17138 (N_17138,N_16777,N_16694);
and U17139 (N_17139,N_16032,N_16283);
xor U17140 (N_17140,N_16674,N_16449);
nand U17141 (N_17141,N_16067,N_16947);
and U17142 (N_17142,N_16465,N_16982);
xnor U17143 (N_17143,N_16577,N_16255);
and U17144 (N_17144,N_16112,N_16944);
or U17145 (N_17145,N_16786,N_16197);
and U17146 (N_17146,N_16282,N_16406);
nor U17147 (N_17147,N_16578,N_16514);
or U17148 (N_17148,N_16361,N_16998);
or U17149 (N_17149,N_16603,N_16574);
xor U17150 (N_17150,N_16990,N_16927);
nor U17151 (N_17151,N_16511,N_16327);
nor U17152 (N_17152,N_16559,N_16014);
or U17153 (N_17153,N_16291,N_16201);
nor U17154 (N_17154,N_16124,N_16482);
xnor U17155 (N_17155,N_16646,N_16846);
nand U17156 (N_17156,N_16949,N_16597);
nor U17157 (N_17157,N_16486,N_16645);
and U17158 (N_17158,N_16560,N_16679);
and U17159 (N_17159,N_16167,N_16928);
or U17160 (N_17160,N_16453,N_16204);
xnor U17161 (N_17161,N_16877,N_16259);
nand U17162 (N_17162,N_16568,N_16083);
nor U17163 (N_17163,N_16305,N_16115);
nor U17164 (N_17164,N_16881,N_16585);
or U17165 (N_17165,N_16648,N_16354);
nand U17166 (N_17166,N_16615,N_16668);
and U17167 (N_17167,N_16141,N_16263);
xor U17168 (N_17168,N_16393,N_16011);
nand U17169 (N_17169,N_16804,N_16207);
or U17170 (N_17170,N_16308,N_16481);
nor U17171 (N_17171,N_16664,N_16281);
nand U17172 (N_17172,N_16864,N_16154);
nor U17173 (N_17173,N_16428,N_16313);
nor U17174 (N_17174,N_16433,N_16334);
nand U17175 (N_17175,N_16179,N_16172);
nor U17176 (N_17176,N_16860,N_16202);
nor U17177 (N_17177,N_16297,N_16543);
nor U17178 (N_17178,N_16920,N_16734);
nand U17179 (N_17179,N_16503,N_16039);
and U17180 (N_17180,N_16515,N_16314);
nand U17181 (N_17181,N_16731,N_16564);
nor U17182 (N_17182,N_16938,N_16774);
xor U17183 (N_17183,N_16824,N_16241);
nand U17184 (N_17184,N_16171,N_16369);
nor U17185 (N_17185,N_16692,N_16588);
nand U17186 (N_17186,N_16048,N_16081);
or U17187 (N_17187,N_16627,N_16320);
nand U17188 (N_17188,N_16820,N_16430);
nor U17189 (N_17189,N_16766,N_16326);
xnor U17190 (N_17190,N_16828,N_16340);
xnor U17191 (N_17191,N_16626,N_16441);
nand U17192 (N_17192,N_16788,N_16302);
or U17193 (N_17193,N_16076,N_16476);
and U17194 (N_17194,N_16122,N_16784);
nor U17195 (N_17195,N_16569,N_16866);
nor U17196 (N_17196,N_16793,N_16425);
nand U17197 (N_17197,N_16483,N_16384);
nor U17198 (N_17198,N_16095,N_16502);
and U17199 (N_17199,N_16266,N_16976);
and U17200 (N_17200,N_16743,N_16934);
xnor U17201 (N_17201,N_16026,N_16951);
and U17202 (N_17202,N_16254,N_16693);
or U17203 (N_17203,N_16558,N_16882);
xnor U17204 (N_17204,N_16557,N_16146);
xnor U17205 (N_17205,N_16901,N_16439);
or U17206 (N_17206,N_16600,N_16049);
or U17207 (N_17207,N_16986,N_16390);
nand U17208 (N_17208,N_16101,N_16965);
and U17209 (N_17209,N_16914,N_16166);
nor U17210 (N_17210,N_16691,N_16992);
nor U17211 (N_17211,N_16888,N_16718);
xor U17212 (N_17212,N_16274,N_16602);
nor U17213 (N_17213,N_16806,N_16593);
or U17214 (N_17214,N_16970,N_16541);
nor U17215 (N_17215,N_16977,N_16030);
or U17216 (N_17216,N_16488,N_16351);
nand U17217 (N_17217,N_16138,N_16392);
xor U17218 (N_17218,N_16714,N_16735);
and U17219 (N_17219,N_16999,N_16687);
or U17220 (N_17220,N_16737,N_16472);
nand U17221 (N_17221,N_16405,N_16156);
xnor U17222 (N_17222,N_16164,N_16250);
and U17223 (N_17223,N_16815,N_16654);
nor U17224 (N_17224,N_16285,N_16165);
and U17225 (N_17225,N_16286,N_16833);
or U17226 (N_17226,N_16093,N_16848);
nor U17227 (N_17227,N_16477,N_16980);
xor U17228 (N_17228,N_16905,N_16492);
xor U17229 (N_17229,N_16016,N_16937);
and U17230 (N_17230,N_16402,N_16740);
nor U17231 (N_17231,N_16343,N_16641);
or U17232 (N_17232,N_16565,N_16085);
nand U17233 (N_17233,N_16400,N_16365);
xnor U17234 (N_17234,N_16395,N_16745);
and U17235 (N_17235,N_16021,N_16531);
xnor U17236 (N_17236,N_16728,N_16218);
xnor U17237 (N_17237,N_16087,N_16290);
xnor U17238 (N_17238,N_16475,N_16323);
nand U17239 (N_17239,N_16741,N_16001);
and U17240 (N_17240,N_16696,N_16335);
nor U17241 (N_17241,N_16709,N_16635);
and U17242 (N_17242,N_16685,N_16208);
and U17243 (N_17243,N_16074,N_16926);
nor U17244 (N_17244,N_16825,N_16902);
xnor U17245 (N_17245,N_16964,N_16677);
or U17246 (N_17246,N_16052,N_16956);
xor U17247 (N_17247,N_16534,N_16632);
nor U17248 (N_17248,N_16125,N_16988);
xnor U17249 (N_17249,N_16997,N_16438);
or U17250 (N_17250,N_16858,N_16870);
nor U17251 (N_17251,N_16796,N_16650);
nor U17252 (N_17252,N_16018,N_16304);
xor U17253 (N_17253,N_16233,N_16002);
nand U17254 (N_17254,N_16567,N_16763);
nand U17255 (N_17255,N_16443,N_16669);
nor U17256 (N_17256,N_16634,N_16177);
nand U17257 (N_17257,N_16730,N_16761);
xnor U17258 (N_17258,N_16324,N_16925);
xor U17259 (N_17259,N_16221,N_16636);
or U17260 (N_17260,N_16591,N_16045);
or U17261 (N_17261,N_16807,N_16510);
and U17262 (N_17262,N_16061,N_16651);
xor U17263 (N_17263,N_16037,N_16385);
nor U17264 (N_17264,N_16529,N_16963);
xnor U17265 (N_17265,N_16228,N_16033);
and U17266 (N_17266,N_16410,N_16216);
and U17267 (N_17267,N_16419,N_16080);
or U17268 (N_17268,N_16331,N_16727);
and U17269 (N_17269,N_16871,N_16198);
and U17270 (N_17270,N_16103,N_16931);
xor U17271 (N_17271,N_16493,N_16388);
or U17272 (N_17272,N_16342,N_16212);
nand U17273 (N_17273,N_16672,N_16236);
nor U17274 (N_17274,N_16181,N_16849);
nand U17275 (N_17275,N_16649,N_16869);
nor U17276 (N_17276,N_16550,N_16484);
nand U17277 (N_17277,N_16414,N_16389);
or U17278 (N_17278,N_16234,N_16604);
or U17279 (N_17279,N_16546,N_16107);
and U17280 (N_17280,N_16573,N_16532);
nand U17281 (N_17281,N_16523,N_16772);
nor U17282 (N_17282,N_16192,N_16270);
and U17283 (N_17283,N_16506,N_16426);
or U17284 (N_17284,N_16826,N_16912);
xnor U17285 (N_17285,N_16832,N_16042);
xnor U17286 (N_17286,N_16710,N_16508);
xor U17287 (N_17287,N_16474,N_16264);
and U17288 (N_17288,N_16656,N_16455);
or U17289 (N_17289,N_16296,N_16072);
nand U17290 (N_17290,N_16943,N_16946);
and U17291 (N_17291,N_16630,N_16129);
nand U17292 (N_17292,N_16671,N_16967);
xnor U17293 (N_17293,N_16357,N_16442);
nor U17294 (N_17294,N_16865,N_16915);
nor U17295 (N_17295,N_16205,N_16605);
xor U17296 (N_17296,N_16711,N_16350);
xor U17297 (N_17297,N_16038,N_16587);
or U17298 (N_17298,N_16173,N_16223);
or U17299 (N_17299,N_16025,N_16090);
or U17300 (N_17300,N_16013,N_16213);
and U17301 (N_17301,N_16617,N_16637);
nand U17302 (N_17302,N_16440,N_16257);
and U17303 (N_17303,N_16681,N_16751);
or U17304 (N_17304,N_16884,N_16989);
or U17305 (N_17305,N_16835,N_16006);
or U17306 (N_17306,N_16427,N_16562);
or U17307 (N_17307,N_16322,N_16856);
and U17308 (N_17308,N_16152,N_16798);
nor U17309 (N_17309,N_16701,N_16903);
nand U17310 (N_17310,N_16237,N_16378);
and U17311 (N_17311,N_16360,N_16226);
and U17312 (N_17312,N_16422,N_16702);
nor U17313 (N_17313,N_16518,N_16193);
or U17314 (N_17314,N_16337,N_16347);
nand U17315 (N_17315,N_16341,N_16450);
or U17316 (N_17316,N_16661,N_16919);
or U17317 (N_17317,N_16556,N_16359);
or U17318 (N_17318,N_16358,N_16528);
or U17319 (N_17319,N_16275,N_16522);
and U17320 (N_17320,N_16612,N_16423);
or U17321 (N_17321,N_16086,N_16245);
nand U17322 (N_17322,N_16507,N_16667);
xor U17323 (N_17323,N_16513,N_16758);
xnor U17324 (N_17324,N_16809,N_16662);
and U17325 (N_17325,N_16215,N_16536);
nand U17326 (N_17326,N_16459,N_16941);
or U17327 (N_17327,N_16874,N_16084);
or U17328 (N_17328,N_16683,N_16401);
or U17329 (N_17329,N_16429,N_16366);
nand U17330 (N_17330,N_16109,N_16975);
nor U17331 (N_17331,N_16209,N_16397);
nand U17332 (N_17332,N_16613,N_16504);
and U17333 (N_17333,N_16723,N_16957);
xnor U17334 (N_17334,N_16252,N_16733);
nand U17335 (N_17335,N_16913,N_16028);
and U17336 (N_17336,N_16720,N_16945);
xnor U17337 (N_17337,N_16417,N_16539);
and U17338 (N_17338,N_16135,N_16719);
xor U17339 (N_17339,N_16123,N_16272);
and U17340 (N_17340,N_16059,N_16579);
or U17341 (N_17341,N_16748,N_16657);
nor U17342 (N_17342,N_16055,N_16180);
and U17343 (N_17343,N_16907,N_16027);
nand U17344 (N_17344,N_16050,N_16176);
or U17345 (N_17345,N_16935,N_16547);
nand U17346 (N_17346,N_16900,N_16586);
or U17347 (N_17347,N_16594,N_16678);
xor U17348 (N_17348,N_16102,N_16773);
and U17349 (N_17349,N_16120,N_16771);
or U17350 (N_17350,N_16435,N_16344);
xnor U17351 (N_17351,N_16596,N_16186);
xor U17352 (N_17352,N_16768,N_16512);
xnor U17353 (N_17353,N_16008,N_16595);
and U17354 (N_17354,N_16238,N_16348);
nor U17355 (N_17355,N_16496,N_16436);
or U17356 (N_17356,N_16019,N_16118);
and U17357 (N_17357,N_16862,N_16017);
and U17358 (N_17358,N_16269,N_16253);
nor U17359 (N_17359,N_16549,N_16972);
nor U17360 (N_17360,N_16699,N_16993);
nor U17361 (N_17361,N_16886,N_16689);
nor U17362 (N_17362,N_16598,N_16230);
or U17363 (N_17363,N_16251,N_16062);
or U17364 (N_17364,N_16398,N_16816);
or U17365 (N_17365,N_16545,N_16895);
and U17366 (N_17366,N_16759,N_16994);
or U17367 (N_17367,N_16007,N_16294);
and U17368 (N_17368,N_16046,N_16448);
nor U17369 (N_17369,N_16535,N_16261);
or U17370 (N_17370,N_16153,N_16640);
or U17371 (N_17371,N_16268,N_16749);
nor U17372 (N_17372,N_16332,N_16879);
xor U17373 (N_17373,N_16461,N_16295);
nand U17374 (N_17374,N_16057,N_16464);
or U17375 (N_17375,N_16729,N_16494);
nand U17376 (N_17376,N_16468,N_16182);
nor U17377 (N_17377,N_16470,N_16309);
xnor U17378 (N_17378,N_16666,N_16068);
nand U17379 (N_17379,N_16063,N_16217);
xnor U17380 (N_17380,N_16760,N_16375);
nand U17381 (N_17381,N_16106,N_16278);
xnor U17382 (N_17382,N_16614,N_16064);
nor U17383 (N_17383,N_16899,N_16908);
or U17384 (N_17384,N_16812,N_16452);
nand U17385 (N_17385,N_16287,N_16185);
nor U17386 (N_17386,N_16330,N_16932);
and U17387 (N_17387,N_16821,N_16367);
nor U17388 (N_17388,N_16151,N_16897);
nand U17389 (N_17389,N_16581,N_16789);
and U17390 (N_17390,N_16169,N_16622);
nor U17391 (N_17391,N_16633,N_16318);
nor U17392 (N_17392,N_16659,N_16362);
and U17393 (N_17393,N_16249,N_16695);
and U17394 (N_17394,N_16813,N_16783);
or U17395 (N_17395,N_16024,N_16029);
and U17396 (N_17396,N_16356,N_16736);
xor U17397 (N_17397,N_16969,N_16889);
nand U17398 (N_17398,N_16299,N_16893);
and U17399 (N_17399,N_16312,N_16995);
nor U17400 (N_17400,N_16676,N_16096);
nand U17401 (N_17401,N_16267,N_16781);
xnor U17402 (N_17402,N_16053,N_16624);
nor U17403 (N_17403,N_16040,N_16576);
nand U17404 (N_17404,N_16962,N_16968);
nor U17405 (N_17405,N_16434,N_16791);
or U17406 (N_17406,N_16829,N_16271);
or U17407 (N_17407,N_16847,N_16805);
nor U17408 (N_17408,N_16861,N_16894);
nand U17409 (N_17409,N_16644,N_16333);
nor U17410 (N_17410,N_16960,N_16184);
xnor U17411 (N_17411,N_16373,N_16794);
xor U17412 (N_17412,N_16170,N_16769);
nand U17413 (N_17413,N_16857,N_16399);
nand U17414 (N_17414,N_16891,N_16363);
xor U17415 (N_17415,N_16620,N_16070);
or U17416 (N_17416,N_16206,N_16936);
xnor U17417 (N_17417,N_16765,N_16725);
and U17418 (N_17418,N_16246,N_16097);
xor U17419 (N_17419,N_16415,N_16372);
or U17420 (N_17420,N_16799,N_16628);
nor U17421 (N_17421,N_16262,N_16121);
nor U17422 (N_17422,N_16639,N_16466);
nand U17423 (N_17423,N_16537,N_16099);
and U17424 (N_17424,N_16407,N_16463);
xnor U17425 (N_17425,N_16954,N_16892);
xor U17426 (N_17426,N_16837,N_16380);
nand U17427 (N_17427,N_16445,N_16853);
xnor U17428 (N_17428,N_16621,N_16851);
xor U17429 (N_17429,N_16175,N_16424);
xor U17430 (N_17430,N_16143,N_16834);
nor U17431 (N_17431,N_16844,N_16570);
or U17432 (N_17432,N_16178,N_16619);
nand U17433 (N_17433,N_16460,N_16643);
or U17434 (N_17434,N_16854,N_16066);
and U17435 (N_17435,N_16301,N_16277);
nor U17436 (N_17436,N_16368,N_16755);
or U17437 (N_17437,N_16047,N_16210);
nor U17438 (N_17438,N_16583,N_16383);
nand U17439 (N_17439,N_16094,N_16906);
xnor U17440 (N_17440,N_16293,N_16034);
nand U17441 (N_17441,N_16303,N_16715);
nor U17442 (N_17442,N_16009,N_16887);
or U17443 (N_17443,N_16929,N_16618);
xor U17444 (N_17444,N_16276,N_16830);
xor U17445 (N_17445,N_16665,N_16010);
xnor U17446 (N_17446,N_16456,N_16722);
or U17447 (N_17447,N_16898,N_16073);
and U17448 (N_17448,N_16770,N_16394);
and U17449 (N_17449,N_16104,N_16930);
nand U17450 (N_17450,N_16757,N_16447);
or U17451 (N_17451,N_16404,N_16137);
or U17452 (N_17452,N_16382,N_16554);
and U17453 (N_17453,N_16035,N_16966);
nor U17454 (N_17454,N_16069,N_16981);
nor U17455 (N_17455,N_16325,N_16219);
nand U17456 (N_17456,N_16713,N_16134);
xnor U17457 (N_17457,N_16139,N_16845);
xnor U17458 (N_17458,N_16673,N_16517);
or U17459 (N_17459,N_16150,N_16060);
nand U17460 (N_17460,N_16985,N_16119);
and U17461 (N_17461,N_16160,N_16823);
nand U17462 (N_17462,N_16653,N_16273);
xnor U17463 (N_17463,N_16149,N_16747);
and U17464 (N_17464,N_16561,N_16631);
nand U17465 (N_17465,N_16675,N_16878);
xor U17466 (N_17466,N_16020,N_16467);
or U17467 (N_17467,N_16036,N_16533);
xnor U17468 (N_17468,N_16940,N_16553);
xnor U17469 (N_17469,N_16022,N_16652);
or U17470 (N_17470,N_16412,N_16527);
or U17471 (N_17471,N_16544,N_16499);
xor U17472 (N_17472,N_16572,N_16117);
nor U17473 (N_17473,N_16566,N_16485);
xnor U17474 (N_17474,N_16552,N_16409);
nor U17475 (N_17475,N_16256,N_16288);
nand U17476 (N_17476,N_16890,N_16775);
nand U17477 (N_17477,N_16904,N_16868);
xor U17478 (N_17478,N_16147,N_16189);
nand U17479 (N_17479,N_16750,N_16284);
or U17480 (N_17480,N_16921,N_16984);
and U17481 (N_17481,N_16345,N_16386);
or U17482 (N_17482,N_16235,N_16200);
and U17483 (N_17483,N_16802,N_16961);
and U17484 (N_17484,N_16243,N_16220);
nand U17485 (N_17485,N_16339,N_16875);
and U17486 (N_17486,N_16548,N_16923);
and U17487 (N_17487,N_16075,N_16738);
nor U17488 (N_17488,N_16088,N_16818);
and U17489 (N_17489,N_16841,N_16551);
xnor U17490 (N_17490,N_16540,N_16091);
nor U17491 (N_17491,N_16127,N_16762);
xnor U17492 (N_17492,N_16827,N_16582);
nand U17493 (N_17493,N_16538,N_16471);
and U17494 (N_17494,N_16432,N_16329);
or U17495 (N_17495,N_16950,N_16716);
xor U17496 (N_17496,N_16555,N_16260);
xor U17497 (N_17497,N_16058,N_16098);
nand U17498 (N_17498,N_16971,N_16917);
xnor U17499 (N_17499,N_16610,N_16480);
or U17500 (N_17500,N_16709,N_16907);
xor U17501 (N_17501,N_16573,N_16910);
or U17502 (N_17502,N_16725,N_16538);
or U17503 (N_17503,N_16800,N_16153);
and U17504 (N_17504,N_16776,N_16971);
xor U17505 (N_17505,N_16209,N_16766);
xor U17506 (N_17506,N_16872,N_16590);
or U17507 (N_17507,N_16295,N_16532);
xnor U17508 (N_17508,N_16844,N_16767);
or U17509 (N_17509,N_16287,N_16805);
xnor U17510 (N_17510,N_16968,N_16856);
xor U17511 (N_17511,N_16053,N_16982);
or U17512 (N_17512,N_16706,N_16629);
and U17513 (N_17513,N_16766,N_16227);
nor U17514 (N_17514,N_16738,N_16031);
nand U17515 (N_17515,N_16506,N_16764);
or U17516 (N_17516,N_16253,N_16432);
nand U17517 (N_17517,N_16689,N_16516);
and U17518 (N_17518,N_16172,N_16300);
nand U17519 (N_17519,N_16704,N_16196);
nand U17520 (N_17520,N_16089,N_16075);
nor U17521 (N_17521,N_16744,N_16750);
or U17522 (N_17522,N_16146,N_16071);
nand U17523 (N_17523,N_16312,N_16152);
xor U17524 (N_17524,N_16511,N_16557);
or U17525 (N_17525,N_16978,N_16396);
and U17526 (N_17526,N_16979,N_16443);
nand U17527 (N_17527,N_16725,N_16099);
or U17528 (N_17528,N_16443,N_16880);
nand U17529 (N_17529,N_16551,N_16519);
nand U17530 (N_17530,N_16368,N_16703);
and U17531 (N_17531,N_16246,N_16858);
nor U17532 (N_17532,N_16493,N_16804);
xor U17533 (N_17533,N_16166,N_16732);
and U17534 (N_17534,N_16528,N_16752);
or U17535 (N_17535,N_16567,N_16096);
or U17536 (N_17536,N_16588,N_16254);
and U17537 (N_17537,N_16943,N_16584);
xnor U17538 (N_17538,N_16055,N_16653);
and U17539 (N_17539,N_16416,N_16434);
nor U17540 (N_17540,N_16247,N_16304);
or U17541 (N_17541,N_16524,N_16151);
xnor U17542 (N_17542,N_16471,N_16334);
and U17543 (N_17543,N_16914,N_16279);
nand U17544 (N_17544,N_16092,N_16329);
and U17545 (N_17545,N_16972,N_16303);
and U17546 (N_17546,N_16260,N_16784);
or U17547 (N_17547,N_16519,N_16812);
nor U17548 (N_17548,N_16103,N_16588);
and U17549 (N_17549,N_16739,N_16818);
nor U17550 (N_17550,N_16688,N_16242);
nor U17551 (N_17551,N_16588,N_16203);
nor U17552 (N_17552,N_16641,N_16288);
and U17553 (N_17553,N_16371,N_16945);
nand U17554 (N_17554,N_16136,N_16441);
nand U17555 (N_17555,N_16802,N_16582);
and U17556 (N_17556,N_16619,N_16432);
nor U17557 (N_17557,N_16717,N_16111);
xnor U17558 (N_17558,N_16505,N_16057);
or U17559 (N_17559,N_16910,N_16838);
and U17560 (N_17560,N_16644,N_16188);
xor U17561 (N_17561,N_16449,N_16607);
or U17562 (N_17562,N_16016,N_16652);
and U17563 (N_17563,N_16639,N_16276);
nand U17564 (N_17564,N_16401,N_16502);
xor U17565 (N_17565,N_16576,N_16911);
nor U17566 (N_17566,N_16177,N_16248);
nand U17567 (N_17567,N_16225,N_16583);
or U17568 (N_17568,N_16168,N_16497);
and U17569 (N_17569,N_16823,N_16054);
and U17570 (N_17570,N_16145,N_16144);
xor U17571 (N_17571,N_16991,N_16458);
nor U17572 (N_17572,N_16898,N_16039);
nand U17573 (N_17573,N_16534,N_16386);
and U17574 (N_17574,N_16872,N_16587);
nor U17575 (N_17575,N_16596,N_16577);
or U17576 (N_17576,N_16692,N_16025);
and U17577 (N_17577,N_16507,N_16861);
nand U17578 (N_17578,N_16996,N_16965);
nand U17579 (N_17579,N_16633,N_16908);
nor U17580 (N_17580,N_16026,N_16444);
nor U17581 (N_17581,N_16677,N_16545);
xor U17582 (N_17582,N_16932,N_16923);
nand U17583 (N_17583,N_16367,N_16945);
and U17584 (N_17584,N_16031,N_16610);
xnor U17585 (N_17585,N_16024,N_16996);
or U17586 (N_17586,N_16215,N_16655);
xnor U17587 (N_17587,N_16918,N_16488);
and U17588 (N_17588,N_16090,N_16372);
xnor U17589 (N_17589,N_16818,N_16874);
and U17590 (N_17590,N_16932,N_16642);
or U17591 (N_17591,N_16592,N_16950);
and U17592 (N_17592,N_16745,N_16915);
nor U17593 (N_17593,N_16514,N_16254);
nand U17594 (N_17594,N_16233,N_16782);
nand U17595 (N_17595,N_16786,N_16582);
or U17596 (N_17596,N_16902,N_16951);
xnor U17597 (N_17597,N_16806,N_16479);
and U17598 (N_17598,N_16418,N_16887);
nand U17599 (N_17599,N_16533,N_16310);
xor U17600 (N_17600,N_16681,N_16749);
nor U17601 (N_17601,N_16727,N_16985);
and U17602 (N_17602,N_16691,N_16551);
nand U17603 (N_17603,N_16882,N_16000);
and U17604 (N_17604,N_16555,N_16920);
nand U17605 (N_17605,N_16766,N_16211);
nand U17606 (N_17606,N_16076,N_16529);
xnor U17607 (N_17607,N_16913,N_16957);
or U17608 (N_17608,N_16779,N_16890);
nor U17609 (N_17609,N_16451,N_16902);
nor U17610 (N_17610,N_16258,N_16041);
xor U17611 (N_17611,N_16476,N_16555);
xor U17612 (N_17612,N_16186,N_16979);
xnor U17613 (N_17613,N_16010,N_16466);
xor U17614 (N_17614,N_16753,N_16693);
xnor U17615 (N_17615,N_16214,N_16381);
nand U17616 (N_17616,N_16837,N_16610);
xor U17617 (N_17617,N_16437,N_16269);
xor U17618 (N_17618,N_16397,N_16351);
xor U17619 (N_17619,N_16613,N_16269);
nor U17620 (N_17620,N_16737,N_16702);
or U17621 (N_17621,N_16699,N_16041);
and U17622 (N_17622,N_16651,N_16596);
xnor U17623 (N_17623,N_16480,N_16351);
nand U17624 (N_17624,N_16075,N_16702);
nor U17625 (N_17625,N_16253,N_16595);
nor U17626 (N_17626,N_16216,N_16173);
nand U17627 (N_17627,N_16491,N_16227);
or U17628 (N_17628,N_16451,N_16559);
nor U17629 (N_17629,N_16900,N_16285);
or U17630 (N_17630,N_16602,N_16950);
nor U17631 (N_17631,N_16617,N_16615);
xor U17632 (N_17632,N_16378,N_16793);
or U17633 (N_17633,N_16551,N_16440);
nor U17634 (N_17634,N_16571,N_16070);
xor U17635 (N_17635,N_16962,N_16627);
nand U17636 (N_17636,N_16841,N_16272);
nand U17637 (N_17637,N_16220,N_16246);
or U17638 (N_17638,N_16971,N_16210);
xor U17639 (N_17639,N_16272,N_16328);
or U17640 (N_17640,N_16803,N_16400);
nor U17641 (N_17641,N_16843,N_16577);
or U17642 (N_17642,N_16858,N_16212);
xnor U17643 (N_17643,N_16879,N_16727);
or U17644 (N_17644,N_16691,N_16018);
xnor U17645 (N_17645,N_16928,N_16529);
and U17646 (N_17646,N_16460,N_16354);
xnor U17647 (N_17647,N_16411,N_16739);
or U17648 (N_17648,N_16113,N_16006);
nor U17649 (N_17649,N_16392,N_16808);
xnor U17650 (N_17650,N_16968,N_16872);
and U17651 (N_17651,N_16866,N_16703);
or U17652 (N_17652,N_16932,N_16151);
xor U17653 (N_17653,N_16497,N_16920);
and U17654 (N_17654,N_16344,N_16932);
and U17655 (N_17655,N_16605,N_16001);
nor U17656 (N_17656,N_16237,N_16615);
xor U17657 (N_17657,N_16877,N_16455);
nand U17658 (N_17658,N_16058,N_16615);
or U17659 (N_17659,N_16440,N_16321);
xnor U17660 (N_17660,N_16877,N_16256);
xor U17661 (N_17661,N_16299,N_16986);
nor U17662 (N_17662,N_16917,N_16705);
and U17663 (N_17663,N_16412,N_16381);
or U17664 (N_17664,N_16734,N_16360);
and U17665 (N_17665,N_16074,N_16625);
nor U17666 (N_17666,N_16727,N_16694);
and U17667 (N_17667,N_16109,N_16271);
nand U17668 (N_17668,N_16081,N_16314);
nor U17669 (N_17669,N_16927,N_16606);
and U17670 (N_17670,N_16061,N_16849);
nand U17671 (N_17671,N_16922,N_16627);
nor U17672 (N_17672,N_16672,N_16106);
or U17673 (N_17673,N_16172,N_16780);
nor U17674 (N_17674,N_16422,N_16239);
or U17675 (N_17675,N_16193,N_16881);
nand U17676 (N_17676,N_16254,N_16975);
nand U17677 (N_17677,N_16274,N_16170);
and U17678 (N_17678,N_16693,N_16204);
or U17679 (N_17679,N_16154,N_16212);
nor U17680 (N_17680,N_16015,N_16173);
and U17681 (N_17681,N_16968,N_16049);
xor U17682 (N_17682,N_16169,N_16164);
or U17683 (N_17683,N_16501,N_16418);
xor U17684 (N_17684,N_16858,N_16203);
nor U17685 (N_17685,N_16568,N_16877);
and U17686 (N_17686,N_16246,N_16954);
or U17687 (N_17687,N_16266,N_16343);
xnor U17688 (N_17688,N_16469,N_16898);
and U17689 (N_17689,N_16327,N_16724);
or U17690 (N_17690,N_16069,N_16552);
nor U17691 (N_17691,N_16317,N_16635);
nor U17692 (N_17692,N_16338,N_16546);
and U17693 (N_17693,N_16969,N_16545);
xnor U17694 (N_17694,N_16694,N_16259);
nand U17695 (N_17695,N_16407,N_16918);
nand U17696 (N_17696,N_16703,N_16040);
nand U17697 (N_17697,N_16527,N_16256);
and U17698 (N_17698,N_16026,N_16732);
or U17699 (N_17699,N_16770,N_16862);
or U17700 (N_17700,N_16705,N_16307);
or U17701 (N_17701,N_16765,N_16899);
and U17702 (N_17702,N_16759,N_16919);
xor U17703 (N_17703,N_16834,N_16612);
and U17704 (N_17704,N_16010,N_16130);
xor U17705 (N_17705,N_16910,N_16228);
and U17706 (N_17706,N_16009,N_16083);
xnor U17707 (N_17707,N_16951,N_16486);
or U17708 (N_17708,N_16357,N_16231);
nand U17709 (N_17709,N_16107,N_16855);
nand U17710 (N_17710,N_16209,N_16465);
nand U17711 (N_17711,N_16744,N_16897);
xor U17712 (N_17712,N_16383,N_16102);
and U17713 (N_17713,N_16013,N_16629);
and U17714 (N_17714,N_16969,N_16861);
xnor U17715 (N_17715,N_16207,N_16106);
nor U17716 (N_17716,N_16337,N_16803);
and U17717 (N_17717,N_16896,N_16521);
or U17718 (N_17718,N_16932,N_16036);
nand U17719 (N_17719,N_16037,N_16363);
nand U17720 (N_17720,N_16971,N_16084);
or U17721 (N_17721,N_16083,N_16429);
and U17722 (N_17722,N_16099,N_16771);
nand U17723 (N_17723,N_16269,N_16747);
or U17724 (N_17724,N_16238,N_16950);
or U17725 (N_17725,N_16770,N_16957);
xor U17726 (N_17726,N_16696,N_16568);
nand U17727 (N_17727,N_16649,N_16825);
nor U17728 (N_17728,N_16984,N_16632);
nor U17729 (N_17729,N_16029,N_16559);
xnor U17730 (N_17730,N_16112,N_16544);
xor U17731 (N_17731,N_16035,N_16506);
and U17732 (N_17732,N_16665,N_16615);
or U17733 (N_17733,N_16383,N_16785);
or U17734 (N_17734,N_16525,N_16895);
and U17735 (N_17735,N_16665,N_16477);
nand U17736 (N_17736,N_16174,N_16055);
nand U17737 (N_17737,N_16009,N_16462);
nor U17738 (N_17738,N_16043,N_16766);
nand U17739 (N_17739,N_16842,N_16662);
xnor U17740 (N_17740,N_16541,N_16530);
and U17741 (N_17741,N_16459,N_16942);
nand U17742 (N_17742,N_16314,N_16309);
or U17743 (N_17743,N_16807,N_16077);
xor U17744 (N_17744,N_16011,N_16698);
xor U17745 (N_17745,N_16624,N_16949);
xor U17746 (N_17746,N_16015,N_16008);
and U17747 (N_17747,N_16612,N_16427);
and U17748 (N_17748,N_16580,N_16239);
nand U17749 (N_17749,N_16577,N_16135);
nand U17750 (N_17750,N_16180,N_16447);
xor U17751 (N_17751,N_16161,N_16412);
or U17752 (N_17752,N_16688,N_16785);
and U17753 (N_17753,N_16278,N_16310);
and U17754 (N_17754,N_16561,N_16253);
or U17755 (N_17755,N_16954,N_16161);
or U17756 (N_17756,N_16109,N_16871);
and U17757 (N_17757,N_16477,N_16457);
nand U17758 (N_17758,N_16444,N_16905);
nor U17759 (N_17759,N_16317,N_16921);
nor U17760 (N_17760,N_16296,N_16257);
nand U17761 (N_17761,N_16723,N_16796);
xor U17762 (N_17762,N_16524,N_16747);
nand U17763 (N_17763,N_16271,N_16955);
or U17764 (N_17764,N_16275,N_16781);
nand U17765 (N_17765,N_16973,N_16700);
or U17766 (N_17766,N_16767,N_16965);
or U17767 (N_17767,N_16797,N_16433);
or U17768 (N_17768,N_16499,N_16304);
nor U17769 (N_17769,N_16834,N_16869);
nand U17770 (N_17770,N_16378,N_16350);
nor U17771 (N_17771,N_16161,N_16373);
nand U17772 (N_17772,N_16185,N_16816);
xnor U17773 (N_17773,N_16288,N_16153);
and U17774 (N_17774,N_16667,N_16465);
nand U17775 (N_17775,N_16495,N_16368);
or U17776 (N_17776,N_16297,N_16301);
and U17777 (N_17777,N_16200,N_16195);
xnor U17778 (N_17778,N_16527,N_16289);
or U17779 (N_17779,N_16268,N_16301);
or U17780 (N_17780,N_16706,N_16525);
nor U17781 (N_17781,N_16048,N_16961);
or U17782 (N_17782,N_16495,N_16406);
or U17783 (N_17783,N_16409,N_16896);
nand U17784 (N_17784,N_16874,N_16956);
nand U17785 (N_17785,N_16891,N_16484);
xor U17786 (N_17786,N_16775,N_16801);
nor U17787 (N_17787,N_16091,N_16015);
xor U17788 (N_17788,N_16705,N_16924);
nand U17789 (N_17789,N_16044,N_16462);
xor U17790 (N_17790,N_16777,N_16863);
nor U17791 (N_17791,N_16056,N_16558);
or U17792 (N_17792,N_16745,N_16218);
and U17793 (N_17793,N_16954,N_16739);
or U17794 (N_17794,N_16374,N_16514);
or U17795 (N_17795,N_16607,N_16513);
and U17796 (N_17796,N_16498,N_16378);
nor U17797 (N_17797,N_16171,N_16890);
nor U17798 (N_17798,N_16069,N_16174);
nand U17799 (N_17799,N_16621,N_16242);
nor U17800 (N_17800,N_16028,N_16684);
and U17801 (N_17801,N_16542,N_16213);
nor U17802 (N_17802,N_16019,N_16378);
nor U17803 (N_17803,N_16869,N_16568);
nor U17804 (N_17804,N_16670,N_16601);
nor U17805 (N_17805,N_16129,N_16183);
xnor U17806 (N_17806,N_16222,N_16262);
nor U17807 (N_17807,N_16902,N_16424);
nand U17808 (N_17808,N_16135,N_16285);
xnor U17809 (N_17809,N_16186,N_16366);
nor U17810 (N_17810,N_16530,N_16826);
xor U17811 (N_17811,N_16912,N_16799);
nor U17812 (N_17812,N_16417,N_16038);
and U17813 (N_17813,N_16261,N_16748);
nand U17814 (N_17814,N_16247,N_16005);
xor U17815 (N_17815,N_16725,N_16424);
and U17816 (N_17816,N_16434,N_16542);
nor U17817 (N_17817,N_16582,N_16637);
or U17818 (N_17818,N_16656,N_16782);
and U17819 (N_17819,N_16130,N_16726);
xor U17820 (N_17820,N_16611,N_16912);
nand U17821 (N_17821,N_16710,N_16723);
or U17822 (N_17822,N_16641,N_16735);
or U17823 (N_17823,N_16947,N_16991);
or U17824 (N_17824,N_16054,N_16491);
nand U17825 (N_17825,N_16560,N_16765);
and U17826 (N_17826,N_16335,N_16613);
or U17827 (N_17827,N_16483,N_16520);
nor U17828 (N_17828,N_16645,N_16795);
nand U17829 (N_17829,N_16533,N_16386);
and U17830 (N_17830,N_16059,N_16202);
and U17831 (N_17831,N_16212,N_16710);
nand U17832 (N_17832,N_16635,N_16948);
and U17833 (N_17833,N_16324,N_16843);
nor U17834 (N_17834,N_16769,N_16825);
xnor U17835 (N_17835,N_16603,N_16389);
nor U17836 (N_17836,N_16785,N_16287);
nor U17837 (N_17837,N_16347,N_16637);
or U17838 (N_17838,N_16040,N_16104);
or U17839 (N_17839,N_16363,N_16709);
nor U17840 (N_17840,N_16263,N_16253);
xor U17841 (N_17841,N_16761,N_16543);
nand U17842 (N_17842,N_16664,N_16623);
or U17843 (N_17843,N_16970,N_16141);
or U17844 (N_17844,N_16026,N_16805);
or U17845 (N_17845,N_16342,N_16589);
xnor U17846 (N_17846,N_16770,N_16316);
or U17847 (N_17847,N_16944,N_16736);
xor U17848 (N_17848,N_16305,N_16827);
and U17849 (N_17849,N_16874,N_16534);
xor U17850 (N_17850,N_16752,N_16003);
or U17851 (N_17851,N_16774,N_16835);
nand U17852 (N_17852,N_16351,N_16798);
and U17853 (N_17853,N_16098,N_16017);
xnor U17854 (N_17854,N_16422,N_16750);
nand U17855 (N_17855,N_16935,N_16799);
and U17856 (N_17856,N_16983,N_16507);
nor U17857 (N_17857,N_16795,N_16979);
or U17858 (N_17858,N_16781,N_16025);
nor U17859 (N_17859,N_16420,N_16836);
and U17860 (N_17860,N_16752,N_16938);
xor U17861 (N_17861,N_16803,N_16910);
nor U17862 (N_17862,N_16913,N_16798);
and U17863 (N_17863,N_16264,N_16167);
nor U17864 (N_17864,N_16260,N_16763);
nand U17865 (N_17865,N_16230,N_16860);
and U17866 (N_17866,N_16054,N_16205);
and U17867 (N_17867,N_16035,N_16019);
xnor U17868 (N_17868,N_16828,N_16269);
xor U17869 (N_17869,N_16674,N_16788);
nand U17870 (N_17870,N_16550,N_16333);
or U17871 (N_17871,N_16708,N_16523);
nand U17872 (N_17872,N_16059,N_16230);
nor U17873 (N_17873,N_16410,N_16051);
nand U17874 (N_17874,N_16358,N_16766);
and U17875 (N_17875,N_16204,N_16668);
nor U17876 (N_17876,N_16076,N_16873);
nand U17877 (N_17877,N_16772,N_16382);
or U17878 (N_17878,N_16154,N_16365);
nor U17879 (N_17879,N_16695,N_16439);
nand U17880 (N_17880,N_16610,N_16671);
nor U17881 (N_17881,N_16549,N_16225);
nor U17882 (N_17882,N_16087,N_16395);
xnor U17883 (N_17883,N_16809,N_16911);
xor U17884 (N_17884,N_16130,N_16802);
nand U17885 (N_17885,N_16124,N_16202);
and U17886 (N_17886,N_16970,N_16343);
xnor U17887 (N_17887,N_16848,N_16339);
and U17888 (N_17888,N_16931,N_16910);
nor U17889 (N_17889,N_16884,N_16877);
or U17890 (N_17890,N_16903,N_16396);
and U17891 (N_17891,N_16081,N_16862);
and U17892 (N_17892,N_16389,N_16116);
nor U17893 (N_17893,N_16669,N_16737);
nand U17894 (N_17894,N_16139,N_16091);
xnor U17895 (N_17895,N_16912,N_16233);
or U17896 (N_17896,N_16698,N_16898);
nand U17897 (N_17897,N_16441,N_16755);
nor U17898 (N_17898,N_16978,N_16317);
or U17899 (N_17899,N_16440,N_16418);
xnor U17900 (N_17900,N_16984,N_16854);
nor U17901 (N_17901,N_16643,N_16288);
xnor U17902 (N_17902,N_16342,N_16480);
and U17903 (N_17903,N_16484,N_16527);
nand U17904 (N_17904,N_16389,N_16054);
nand U17905 (N_17905,N_16018,N_16511);
nand U17906 (N_17906,N_16303,N_16636);
nor U17907 (N_17907,N_16380,N_16841);
and U17908 (N_17908,N_16686,N_16835);
or U17909 (N_17909,N_16770,N_16114);
or U17910 (N_17910,N_16712,N_16213);
nand U17911 (N_17911,N_16922,N_16496);
nor U17912 (N_17912,N_16524,N_16754);
or U17913 (N_17913,N_16593,N_16535);
nand U17914 (N_17914,N_16298,N_16512);
xnor U17915 (N_17915,N_16012,N_16633);
and U17916 (N_17916,N_16111,N_16402);
nand U17917 (N_17917,N_16705,N_16608);
nand U17918 (N_17918,N_16577,N_16299);
xor U17919 (N_17919,N_16774,N_16863);
nor U17920 (N_17920,N_16411,N_16470);
or U17921 (N_17921,N_16890,N_16475);
nand U17922 (N_17922,N_16541,N_16402);
xnor U17923 (N_17923,N_16736,N_16475);
xor U17924 (N_17924,N_16923,N_16326);
and U17925 (N_17925,N_16902,N_16721);
xnor U17926 (N_17926,N_16077,N_16983);
and U17927 (N_17927,N_16749,N_16145);
nor U17928 (N_17928,N_16464,N_16338);
and U17929 (N_17929,N_16304,N_16561);
nor U17930 (N_17930,N_16587,N_16659);
and U17931 (N_17931,N_16863,N_16386);
or U17932 (N_17932,N_16735,N_16747);
and U17933 (N_17933,N_16705,N_16565);
or U17934 (N_17934,N_16482,N_16126);
nor U17935 (N_17935,N_16317,N_16180);
nor U17936 (N_17936,N_16401,N_16725);
nand U17937 (N_17937,N_16850,N_16183);
nand U17938 (N_17938,N_16481,N_16288);
or U17939 (N_17939,N_16479,N_16492);
xor U17940 (N_17940,N_16048,N_16173);
nand U17941 (N_17941,N_16284,N_16573);
nor U17942 (N_17942,N_16771,N_16468);
and U17943 (N_17943,N_16588,N_16698);
nor U17944 (N_17944,N_16498,N_16223);
and U17945 (N_17945,N_16076,N_16670);
and U17946 (N_17946,N_16125,N_16900);
nor U17947 (N_17947,N_16997,N_16501);
xor U17948 (N_17948,N_16901,N_16876);
nor U17949 (N_17949,N_16328,N_16746);
and U17950 (N_17950,N_16792,N_16419);
nand U17951 (N_17951,N_16755,N_16090);
and U17952 (N_17952,N_16888,N_16162);
and U17953 (N_17953,N_16627,N_16676);
or U17954 (N_17954,N_16160,N_16873);
and U17955 (N_17955,N_16400,N_16869);
nor U17956 (N_17956,N_16181,N_16923);
nor U17957 (N_17957,N_16714,N_16363);
nor U17958 (N_17958,N_16784,N_16693);
and U17959 (N_17959,N_16894,N_16390);
xor U17960 (N_17960,N_16879,N_16048);
xnor U17961 (N_17961,N_16086,N_16874);
and U17962 (N_17962,N_16230,N_16122);
or U17963 (N_17963,N_16108,N_16340);
nor U17964 (N_17964,N_16525,N_16528);
or U17965 (N_17965,N_16641,N_16764);
nand U17966 (N_17966,N_16324,N_16746);
nand U17967 (N_17967,N_16445,N_16470);
nand U17968 (N_17968,N_16249,N_16372);
or U17969 (N_17969,N_16517,N_16523);
nor U17970 (N_17970,N_16306,N_16427);
nor U17971 (N_17971,N_16997,N_16540);
nor U17972 (N_17972,N_16886,N_16037);
nor U17973 (N_17973,N_16734,N_16488);
nor U17974 (N_17974,N_16978,N_16651);
nor U17975 (N_17975,N_16440,N_16332);
or U17976 (N_17976,N_16228,N_16924);
nor U17977 (N_17977,N_16712,N_16902);
or U17978 (N_17978,N_16741,N_16496);
or U17979 (N_17979,N_16149,N_16429);
and U17980 (N_17980,N_16761,N_16507);
xnor U17981 (N_17981,N_16607,N_16279);
nor U17982 (N_17982,N_16996,N_16763);
and U17983 (N_17983,N_16463,N_16820);
xor U17984 (N_17984,N_16502,N_16427);
nand U17985 (N_17985,N_16968,N_16721);
and U17986 (N_17986,N_16852,N_16650);
nor U17987 (N_17987,N_16806,N_16978);
xor U17988 (N_17988,N_16289,N_16990);
nor U17989 (N_17989,N_16693,N_16715);
or U17990 (N_17990,N_16944,N_16227);
xnor U17991 (N_17991,N_16142,N_16368);
nor U17992 (N_17992,N_16579,N_16866);
nor U17993 (N_17993,N_16580,N_16495);
nor U17994 (N_17994,N_16215,N_16870);
or U17995 (N_17995,N_16497,N_16368);
and U17996 (N_17996,N_16190,N_16452);
nand U17997 (N_17997,N_16507,N_16956);
and U17998 (N_17998,N_16207,N_16950);
xor U17999 (N_17999,N_16264,N_16080);
nor U18000 (N_18000,N_17536,N_17485);
or U18001 (N_18001,N_17756,N_17892);
nand U18002 (N_18002,N_17941,N_17068);
nor U18003 (N_18003,N_17552,N_17030);
or U18004 (N_18004,N_17126,N_17138);
xor U18005 (N_18005,N_17064,N_17752);
and U18006 (N_18006,N_17954,N_17712);
nor U18007 (N_18007,N_17533,N_17759);
nand U18008 (N_18008,N_17402,N_17390);
nand U18009 (N_18009,N_17385,N_17491);
nand U18010 (N_18010,N_17884,N_17793);
nand U18011 (N_18011,N_17420,N_17803);
nand U18012 (N_18012,N_17155,N_17936);
or U18013 (N_18013,N_17798,N_17612);
nand U18014 (N_18014,N_17487,N_17576);
xor U18015 (N_18015,N_17422,N_17180);
or U18016 (N_18016,N_17249,N_17719);
or U18017 (N_18017,N_17111,N_17261);
nand U18018 (N_18018,N_17382,N_17010);
xor U18019 (N_18019,N_17538,N_17474);
nor U18020 (N_18020,N_17739,N_17226);
and U18021 (N_18021,N_17670,N_17925);
nand U18022 (N_18022,N_17074,N_17646);
xor U18023 (N_18023,N_17514,N_17541);
nor U18024 (N_18024,N_17366,N_17315);
nand U18025 (N_18025,N_17036,N_17707);
or U18026 (N_18026,N_17225,N_17563);
or U18027 (N_18027,N_17475,N_17592);
nand U18028 (N_18028,N_17253,N_17968);
or U18029 (N_18029,N_17800,N_17201);
nand U18030 (N_18030,N_17312,N_17205);
nand U18031 (N_18031,N_17910,N_17100);
or U18032 (N_18032,N_17096,N_17145);
nand U18033 (N_18033,N_17935,N_17280);
nor U18034 (N_18034,N_17808,N_17579);
or U18035 (N_18035,N_17848,N_17518);
xnor U18036 (N_18036,N_17499,N_17250);
nor U18037 (N_18037,N_17822,N_17147);
nand U18038 (N_18038,N_17025,N_17221);
nand U18039 (N_18039,N_17635,N_17015);
nand U18040 (N_18040,N_17160,N_17995);
nor U18041 (N_18041,N_17729,N_17715);
or U18042 (N_18042,N_17951,N_17292);
and U18043 (N_18043,N_17718,N_17634);
and U18044 (N_18044,N_17726,N_17501);
xnor U18045 (N_18045,N_17802,N_17773);
nand U18046 (N_18046,N_17983,N_17703);
xnor U18047 (N_18047,N_17710,N_17686);
and U18048 (N_18048,N_17734,N_17982);
xnor U18049 (N_18049,N_17887,N_17853);
nor U18050 (N_18050,N_17188,N_17206);
or U18051 (N_18051,N_17128,N_17316);
and U18052 (N_18052,N_17764,N_17048);
and U18053 (N_18053,N_17016,N_17108);
xnor U18054 (N_18054,N_17072,N_17319);
nand U18055 (N_18055,N_17920,N_17489);
or U18056 (N_18056,N_17886,N_17173);
nand U18057 (N_18057,N_17717,N_17926);
nand U18058 (N_18058,N_17133,N_17243);
or U18059 (N_18059,N_17512,N_17031);
xor U18060 (N_18060,N_17595,N_17400);
nor U18061 (N_18061,N_17568,N_17027);
nand U18062 (N_18062,N_17999,N_17948);
xor U18063 (N_18063,N_17905,N_17247);
nand U18064 (N_18064,N_17771,N_17866);
nor U18065 (N_18065,N_17114,N_17236);
nand U18066 (N_18066,N_17471,N_17680);
and U18067 (N_18067,N_17085,N_17813);
nor U18068 (N_18068,N_17414,N_17241);
nor U18069 (N_18069,N_17812,N_17616);
nand U18070 (N_18070,N_17934,N_17855);
nor U18071 (N_18071,N_17311,N_17796);
nand U18072 (N_18072,N_17020,N_17258);
nand U18073 (N_18073,N_17341,N_17346);
nor U18074 (N_18074,N_17164,N_17288);
nand U18075 (N_18075,N_17989,N_17478);
nor U18076 (N_18076,N_17377,N_17486);
nand U18077 (N_18077,N_17678,N_17338);
or U18078 (N_18078,N_17484,N_17349);
nor U18079 (N_18079,N_17271,N_17156);
xor U18080 (N_18080,N_17012,N_17996);
and U18081 (N_18081,N_17219,N_17668);
and U18082 (N_18082,N_17305,N_17640);
xnor U18083 (N_18083,N_17482,N_17456);
xnor U18084 (N_18084,N_17467,N_17135);
nand U18085 (N_18085,N_17902,N_17529);
xnor U18086 (N_18086,N_17861,N_17659);
nor U18087 (N_18087,N_17702,N_17768);
and U18088 (N_18088,N_17785,N_17916);
nand U18089 (N_18089,N_17539,N_17758);
and U18090 (N_18090,N_17464,N_17460);
and U18091 (N_18091,N_17748,N_17371);
or U18092 (N_18092,N_17961,N_17617);
or U18093 (N_18093,N_17110,N_17823);
and U18094 (N_18094,N_17361,N_17667);
or U18095 (N_18095,N_17778,N_17384);
xor U18096 (N_18096,N_17379,N_17921);
nor U18097 (N_18097,N_17652,N_17988);
nand U18098 (N_18098,N_17090,N_17714);
or U18099 (N_18099,N_17870,N_17880);
nor U18100 (N_18100,N_17570,N_17820);
or U18101 (N_18101,N_17291,N_17614);
xnor U18102 (N_18102,N_17666,N_17063);
nand U18103 (N_18103,N_17567,N_17875);
nor U18104 (N_18104,N_17166,N_17987);
nor U18105 (N_18105,N_17720,N_17928);
xor U18106 (N_18106,N_17628,N_17244);
or U18107 (N_18107,N_17194,N_17270);
nor U18108 (N_18108,N_17192,N_17904);
and U18109 (N_18109,N_17537,N_17300);
or U18110 (N_18110,N_17560,N_17781);
or U18111 (N_18111,N_17858,N_17769);
and U18112 (N_18112,N_17894,N_17842);
and U18113 (N_18113,N_17295,N_17237);
nand U18114 (N_18114,N_17348,N_17106);
and U18115 (N_18115,N_17607,N_17397);
nand U18116 (N_18116,N_17336,N_17028);
nand U18117 (N_18117,N_17682,N_17184);
and U18118 (N_18118,N_17801,N_17101);
or U18119 (N_18119,N_17623,N_17446);
and U18120 (N_18120,N_17962,N_17056);
nor U18121 (N_18121,N_17024,N_17955);
nand U18122 (N_18122,N_17387,N_17555);
or U18123 (N_18123,N_17774,N_17865);
nor U18124 (N_18124,N_17179,N_17692);
or U18125 (N_18125,N_17044,N_17091);
nor U18126 (N_18126,N_17797,N_17805);
or U18127 (N_18127,N_17468,N_17094);
nand U18128 (N_18128,N_17506,N_17893);
nand U18129 (N_18129,N_17980,N_17510);
nor U18130 (N_18130,N_17549,N_17564);
and U18131 (N_18131,N_17099,N_17701);
or U18132 (N_18132,N_17017,N_17942);
xnor U18133 (N_18133,N_17647,N_17411);
nand U18134 (N_18134,N_17738,N_17621);
nor U18135 (N_18135,N_17391,N_17907);
nor U18136 (N_18136,N_17151,N_17203);
or U18137 (N_18137,N_17172,N_17519);
nor U18138 (N_18138,N_17439,N_17586);
or U18139 (N_18139,N_17727,N_17424);
xor U18140 (N_18140,N_17359,N_17144);
and U18141 (N_18141,N_17867,N_17588);
and U18142 (N_18142,N_17208,N_17606);
or U18143 (N_18143,N_17814,N_17122);
xnor U18144 (N_18144,N_17932,N_17331);
nand U18145 (N_18145,N_17252,N_17087);
nor U18146 (N_18146,N_17075,N_17648);
nand U18147 (N_18147,N_17490,N_17146);
and U18148 (N_18148,N_17083,N_17217);
or U18149 (N_18149,N_17945,N_17081);
nand U18150 (N_18150,N_17076,N_17078);
nor U18151 (N_18151,N_17406,N_17055);
and U18152 (N_18152,N_17084,N_17140);
and U18153 (N_18153,N_17214,N_17791);
or U18154 (N_18154,N_17129,N_17077);
and U18155 (N_18155,N_17511,N_17381);
xnor U18156 (N_18156,N_17283,N_17974);
nor U18157 (N_18157,N_17985,N_17461);
and U18158 (N_18158,N_17417,N_17368);
nand U18159 (N_18159,N_17660,N_17161);
or U18160 (N_18160,N_17545,N_17838);
and U18161 (N_18161,N_17662,N_17515);
xnor U18162 (N_18162,N_17131,N_17363);
nor U18163 (N_18163,N_17428,N_17939);
xor U18164 (N_18164,N_17504,N_17540);
nor U18165 (N_18165,N_17594,N_17896);
xor U18166 (N_18166,N_17001,N_17903);
or U18167 (N_18167,N_17767,N_17038);
and U18168 (N_18168,N_17405,N_17704);
nor U18169 (N_18169,N_17553,N_17685);
or U18170 (N_18170,N_17223,N_17550);
and U18171 (N_18171,N_17824,N_17644);
nor U18172 (N_18172,N_17324,N_17218);
xnor U18173 (N_18173,N_17911,N_17565);
nor U18174 (N_18174,N_17760,N_17380);
nor U18175 (N_18175,N_17437,N_17859);
or U18176 (N_18176,N_17679,N_17232);
or U18177 (N_18177,N_17216,N_17517);
nand U18178 (N_18178,N_17465,N_17889);
nor U18179 (N_18179,N_17357,N_17998);
nand U18180 (N_18180,N_17345,N_17624);
xnor U18181 (N_18181,N_17642,N_17375);
nor U18182 (N_18182,N_17260,N_17722);
and U18183 (N_18183,N_17953,N_17878);
nor U18184 (N_18184,N_17693,N_17210);
nor U18185 (N_18185,N_17593,N_17011);
nor U18186 (N_18186,N_17370,N_17060);
xor U18187 (N_18187,N_17403,N_17732);
and U18188 (N_18188,N_17883,N_17170);
xnor U18189 (N_18189,N_17965,N_17435);
or U18190 (N_18190,N_17153,N_17119);
nor U18191 (N_18191,N_17211,N_17065);
and U18192 (N_18192,N_17229,N_17636);
nand U18193 (N_18193,N_17190,N_17285);
xnor U18194 (N_18194,N_17154,N_17275);
xnor U18195 (N_18195,N_17625,N_17829);
and U18196 (N_18196,N_17248,N_17834);
and U18197 (N_18197,N_17228,N_17638);
and U18198 (N_18198,N_17240,N_17990);
or U18199 (N_18199,N_17958,N_17466);
and U18200 (N_18200,N_17924,N_17169);
nor U18201 (N_18201,N_17964,N_17828);
xor U18202 (N_18202,N_17806,N_17852);
xor U18203 (N_18203,N_17535,N_17480);
and U18204 (N_18204,N_17373,N_17502);
nand U18205 (N_18205,N_17079,N_17994);
xor U18206 (N_18206,N_17868,N_17067);
nand U18207 (N_18207,N_17239,N_17672);
nor U18208 (N_18208,N_17608,N_17789);
xor U18209 (N_18209,N_17765,N_17815);
and U18210 (N_18210,N_17290,N_17917);
xnor U18211 (N_18211,N_17575,N_17620);
and U18212 (N_18212,N_17613,N_17675);
or U18213 (N_18213,N_17843,N_17627);
xnor U18214 (N_18214,N_17120,N_17849);
and U18215 (N_18215,N_17691,N_17835);
nand U18216 (N_18216,N_17947,N_17254);
and U18217 (N_18217,N_17062,N_17113);
or U18218 (N_18218,N_17654,N_17037);
nand U18219 (N_18219,N_17582,N_17195);
or U18220 (N_18220,N_17080,N_17429);
nand U18221 (N_18221,N_17209,N_17603);
nand U18222 (N_18222,N_17202,N_17699);
nand U18223 (N_18223,N_17455,N_17657);
xor U18224 (N_18224,N_17115,N_17421);
and U18225 (N_18225,N_17394,N_17423);
nor U18226 (N_18226,N_17124,N_17107);
nand U18227 (N_18227,N_17294,N_17335);
nand U18228 (N_18228,N_17671,N_17943);
xor U18229 (N_18229,N_17522,N_17329);
nand U18230 (N_18230,N_17753,N_17505);
or U18231 (N_18231,N_17137,N_17032);
nand U18232 (N_18232,N_17189,N_17493);
or U18233 (N_18233,N_17775,N_17591);
or U18234 (N_18234,N_17963,N_17061);
nand U18235 (N_18235,N_17543,N_17658);
nand U18236 (N_18236,N_17374,N_17754);
nor U18237 (N_18237,N_17117,N_17021);
nand U18238 (N_18238,N_17321,N_17503);
xnor U18239 (N_18239,N_17134,N_17182);
and U18240 (N_18240,N_17677,N_17578);
nor U18241 (N_18241,N_17314,N_17246);
nor U18242 (N_18242,N_17255,N_17600);
nand U18243 (N_18243,N_17708,N_17794);
xor U18244 (N_18244,N_17105,N_17003);
nand U18245 (N_18245,N_17334,N_17562);
or U18246 (N_18246,N_17150,N_17112);
or U18247 (N_18247,N_17799,N_17419);
or U18248 (N_18248,N_17496,N_17966);
nand U18249 (N_18249,N_17757,N_17330);
and U18250 (N_18250,N_17123,N_17443);
nor U18251 (N_18251,N_17408,N_17130);
nand U18252 (N_18252,N_17877,N_17508);
and U18253 (N_18253,N_17697,N_17973);
xor U18254 (N_18254,N_17267,N_17946);
nor U18255 (N_18255,N_17933,N_17299);
nor U18256 (N_18256,N_17454,N_17959);
xor U18257 (N_18257,N_17895,N_17093);
or U18258 (N_18258,N_17053,N_17665);
xnor U18259 (N_18259,N_17035,N_17615);
and U18260 (N_18260,N_17873,N_17470);
and U18261 (N_18261,N_17930,N_17833);
or U18262 (N_18262,N_17526,N_17304);
xor U18263 (N_18263,N_17876,N_17103);
xnor U18264 (N_18264,N_17302,N_17281);
nor U18265 (N_18265,N_17971,N_17050);
or U18266 (N_18266,N_17908,N_17817);
xor U18267 (N_18267,N_17554,N_17527);
nor U18268 (N_18268,N_17580,N_17557);
nor U18269 (N_18269,N_17197,N_17238);
or U18270 (N_18270,N_17874,N_17899);
nor U18271 (N_18271,N_17872,N_17328);
nand U18272 (N_18272,N_17006,N_17749);
and U18273 (N_18273,N_17818,N_17353);
nand U18274 (N_18274,N_17495,N_17365);
or U18275 (N_18275,N_17674,N_17610);
or U18276 (N_18276,N_17694,N_17497);
xnor U18277 (N_18277,N_17181,N_17332);
xnor U18278 (N_18278,N_17307,N_17376);
xnor U18279 (N_18279,N_17171,N_17234);
xor U18280 (N_18280,N_17746,N_17698);
nand U18281 (N_18281,N_17597,N_17297);
and U18282 (N_18282,N_17967,N_17457);
xor U18283 (N_18283,N_17816,N_17528);
or U18284 (N_18284,N_17645,N_17839);
and U18285 (N_18285,N_17742,N_17043);
or U18286 (N_18286,N_17755,N_17569);
nand U18287 (N_18287,N_17132,N_17860);
and U18288 (N_18288,N_17212,N_17199);
nand U18289 (N_18289,N_17744,N_17684);
nor U18290 (N_18290,N_17780,N_17287);
xor U18291 (N_18291,N_17441,N_17676);
and U18292 (N_18292,N_17819,N_17434);
or U18293 (N_18293,N_17398,N_17279);
xor U18294 (N_18294,N_17416,N_17022);
nand U18295 (N_18295,N_17176,N_17159);
nor U18296 (N_18296,N_17596,N_17289);
nor U18297 (N_18297,N_17763,N_17054);
nor U18298 (N_18298,N_17264,N_17811);
nor U18299 (N_18299,N_17364,N_17262);
nand U18300 (N_18300,N_17804,N_17433);
and U18301 (N_18301,N_17844,N_17949);
or U18302 (N_18302,N_17548,N_17034);
nand U18303 (N_18303,N_17918,N_17268);
or U18304 (N_18304,N_17303,N_17871);
xnor U18305 (N_18305,N_17831,N_17750);
nor U18306 (N_18306,N_17097,N_17242);
xor U18307 (N_18307,N_17204,N_17761);
nor U18308 (N_18308,N_17383,N_17730);
nand U18309 (N_18309,N_17590,N_17661);
nor U18310 (N_18310,N_17784,N_17323);
or U18311 (N_18311,N_17498,N_17599);
and U18312 (N_18312,N_17970,N_17890);
nor U18313 (N_18313,N_17779,N_17018);
nor U18314 (N_18314,N_17681,N_17436);
and U18315 (N_18315,N_17787,N_17230);
or U18316 (N_18316,N_17325,N_17040);
nor U18317 (N_18317,N_17556,N_17696);
xnor U18318 (N_18318,N_17656,N_17409);
nor U18319 (N_18319,N_17066,N_17004);
or U18320 (N_18320,N_17847,N_17278);
and U18321 (N_18321,N_17972,N_17426);
nand U18322 (N_18322,N_17125,N_17388);
nor U18323 (N_18323,N_17007,N_17837);
or U18324 (N_18324,N_17566,N_17558);
nand U18325 (N_18325,N_17919,N_17604);
nand U18326 (N_18326,N_17431,N_17534);
and U18327 (N_18327,N_17492,N_17396);
nand U18328 (N_18328,N_17452,N_17187);
xnor U18329 (N_18329,N_17263,N_17783);
nand U18330 (N_18330,N_17418,N_17574);
nor U18331 (N_18331,N_17786,N_17960);
or U18332 (N_18332,N_17997,N_17149);
or U18333 (N_18333,N_17807,N_17168);
xor U18334 (N_18334,N_17737,N_17047);
nand U18335 (N_18335,N_17864,N_17157);
xnor U18336 (N_18336,N_17898,N_17273);
nand U18337 (N_18337,N_17944,N_17045);
and U18338 (N_18338,N_17274,N_17337);
nor U18339 (N_18339,N_17602,N_17977);
nand U18340 (N_18340,N_17389,N_17673);
or U18341 (N_18341,N_17683,N_17809);
nor U18342 (N_18342,N_17913,N_17082);
xnor U18343 (N_18343,N_17029,N_17795);
and U18344 (N_18344,N_17826,N_17836);
or U18345 (N_18345,N_17631,N_17220);
nor U18346 (N_18346,N_17448,N_17709);
or U18347 (N_18347,N_17000,N_17630);
and U18348 (N_18348,N_17222,N_17412);
and U18349 (N_18349,N_17937,N_17019);
nor U18350 (N_18350,N_17444,N_17378);
and U18351 (N_18351,N_17013,N_17770);
nand U18352 (N_18352,N_17976,N_17888);
nor U18353 (N_18353,N_17601,N_17581);
nor U18354 (N_18354,N_17728,N_17162);
xor U18355 (N_18355,N_17102,N_17923);
nand U18356 (N_18356,N_17059,N_17619);
nor U18357 (N_18357,N_17788,N_17821);
or U18358 (N_18358,N_17462,N_17143);
nor U18359 (N_18359,N_17598,N_17520);
nand U18360 (N_18360,N_17825,N_17632);
nand U18361 (N_18361,N_17846,N_17320);
nor U18362 (N_18362,N_17716,N_17049);
nand U18363 (N_18363,N_17469,N_17415);
nand U18364 (N_18364,N_17731,N_17360);
nand U18365 (N_18365,N_17915,N_17741);
and U18366 (N_18366,N_17583,N_17979);
and U18367 (N_18367,N_17559,N_17463);
nand U18368 (N_18368,N_17762,N_17473);
nand U18369 (N_18369,N_17148,N_17978);
or U18370 (N_18370,N_17142,N_17981);
or U18371 (N_18371,N_17276,N_17885);
nor U18372 (N_18372,N_17909,N_17751);
or U18373 (N_18373,N_17723,N_17882);
nand U18374 (N_18374,N_17639,N_17339);
or U18375 (N_18375,N_17914,N_17792);
and U18376 (N_18376,N_17458,N_17386);
and U18377 (N_18377,N_17931,N_17929);
xnor U18378 (N_18378,N_17459,N_17743);
or U18379 (N_18379,N_17840,N_17956);
and U18380 (N_18380,N_17425,N_17185);
xor U18381 (N_18381,N_17641,N_17392);
and U18382 (N_18382,N_17183,N_17367);
xnor U18383 (N_18383,N_17139,N_17827);
and U18384 (N_18384,N_17706,N_17587);
or U18385 (N_18385,N_17927,N_17705);
nand U18386 (N_18386,N_17700,N_17663);
nand U18387 (N_18387,N_17362,N_17445);
and U18388 (N_18388,N_17098,N_17207);
and U18389 (N_18389,N_17863,N_17571);
nand U18390 (N_18390,N_17174,N_17584);
nor U18391 (N_18391,N_17393,N_17313);
xnor U18392 (N_18392,N_17284,N_17688);
or U18393 (N_18393,N_17310,N_17326);
or U18394 (N_18394,N_17224,N_17629);
and U18395 (N_18395,N_17404,N_17104);
nand U18396 (N_18396,N_17637,N_17922);
nand U18397 (N_18397,N_17879,N_17272);
and U18398 (N_18398,N_17650,N_17235);
or U18399 (N_18399,N_17810,N_17191);
nor U18400 (N_18400,N_17413,N_17088);
xor U18401 (N_18401,N_17513,N_17857);
and U18402 (N_18402,N_17440,N_17186);
or U18403 (N_18403,N_17095,N_17309);
or U18404 (N_18404,N_17561,N_17293);
and U18405 (N_18405,N_17109,N_17344);
nand U18406 (N_18406,N_17449,N_17069);
nor U18407 (N_18407,N_17286,N_17790);
or U18408 (N_18408,N_17906,N_17343);
nor U18409 (N_18409,N_17116,N_17546);
or U18410 (N_18410,N_17127,N_17735);
nand U18411 (N_18411,N_17163,N_17993);
xnor U18412 (N_18412,N_17507,N_17736);
and U18413 (N_18413,N_17488,N_17351);
nor U18414 (N_18414,N_17633,N_17724);
and U18415 (N_18415,N_17845,N_17891);
and U18416 (N_18416,N_17442,N_17118);
nor U18417 (N_18417,N_17900,N_17301);
nor U18418 (N_18418,N_17782,N_17251);
and U18419 (N_18419,N_17141,N_17327);
nand U18420 (N_18420,N_17342,N_17643);
and U18421 (N_18421,N_17296,N_17052);
or U18422 (N_18422,N_17352,N_17523);
nand U18423 (N_18423,N_17766,N_17058);
xor U18424 (N_18424,N_17957,N_17841);
xor U18425 (N_18425,N_17450,N_17950);
or U18426 (N_18426,N_17984,N_17086);
or U18427 (N_18427,N_17269,N_17651);
xor U18428 (N_18428,N_17399,N_17711);
or U18429 (N_18429,N_17009,N_17432);
and U18430 (N_18430,N_17026,N_17542);
nor U18431 (N_18431,N_17525,N_17605);
or U18432 (N_18432,N_17777,N_17483);
and U18433 (N_18433,N_17041,N_17481);
nand U18434 (N_18434,N_17227,N_17472);
nand U18435 (N_18435,N_17573,N_17215);
or U18436 (N_18436,N_17023,N_17832);
nor U18437 (N_18437,N_17350,N_17664);
nor U18438 (N_18438,N_17854,N_17008);
or U18439 (N_18439,N_17577,N_17477);
nand U18440 (N_18440,N_17725,N_17516);
and U18441 (N_18441,N_17175,N_17585);
nand U18442 (N_18442,N_17524,N_17358);
nor U18443 (N_18443,N_17282,N_17317);
nor U18444 (N_18444,N_17039,N_17695);
or U18445 (N_18445,N_17500,N_17051);
xor U18446 (N_18446,N_17057,N_17940);
and U18447 (N_18447,N_17745,N_17121);
nor U18448 (N_18448,N_17356,N_17213);
and U18449 (N_18449,N_17177,N_17669);
or U18450 (N_18450,N_17862,N_17551);
and U18451 (N_18451,N_17509,N_17046);
xor U18452 (N_18452,N_17198,N_17622);
nor U18453 (N_18453,N_17740,N_17430);
xnor U18454 (N_18454,N_17298,N_17869);
or U18455 (N_18455,N_17347,N_17609);
xor U18456 (N_18456,N_17354,N_17649);
nand U18457 (N_18457,N_17265,N_17196);
nor U18458 (N_18458,N_17395,N_17333);
xnor U18459 (N_18459,N_17689,N_17901);
nor U18460 (N_18460,N_17969,N_17033);
xnor U18461 (N_18461,N_17136,N_17521);
nor U18462 (N_18462,N_17407,N_17447);
nor U18463 (N_18463,N_17547,N_17850);
or U18464 (N_18464,N_17451,N_17092);
nand U18465 (N_18465,N_17002,N_17626);
nor U18466 (N_18466,N_17611,N_17257);
xor U18467 (N_18467,N_17733,N_17005);
and U18468 (N_18468,N_17200,N_17992);
nand U18469 (N_18469,N_17572,N_17193);
xor U18470 (N_18470,N_17231,N_17152);
nor U18471 (N_18471,N_17479,N_17308);
xor U18472 (N_18472,N_17991,N_17256);
nand U18473 (N_18473,N_17975,N_17912);
and U18474 (N_18474,N_17476,N_17372);
nand U18475 (N_18475,N_17938,N_17544);
nor U18476 (N_18476,N_17532,N_17881);
xor U18477 (N_18477,N_17687,N_17772);
or U18478 (N_18478,N_17165,N_17277);
nor U18479 (N_18479,N_17318,N_17952);
nand U18480 (N_18480,N_17158,N_17340);
nor U18481 (N_18481,N_17856,N_17071);
or U18482 (N_18482,N_17830,N_17986);
xor U18483 (N_18483,N_17245,N_17178);
and U18484 (N_18484,N_17369,N_17530);
nand U18485 (N_18485,N_17655,N_17259);
nor U18486 (N_18486,N_17427,N_17851);
or U18487 (N_18487,N_17453,N_17618);
xor U18488 (N_18488,N_17014,N_17167);
nor U18489 (N_18489,N_17721,N_17306);
nand U18490 (N_18490,N_17690,N_17531);
and U18491 (N_18491,N_17355,N_17073);
nor U18492 (N_18492,N_17747,N_17589);
or U18493 (N_18493,N_17653,N_17322);
or U18494 (N_18494,N_17776,N_17401);
nor U18495 (N_18495,N_17070,N_17042);
nand U18496 (N_18496,N_17233,N_17494);
nand U18497 (N_18497,N_17089,N_17266);
xnor U18498 (N_18498,N_17897,N_17410);
nor U18499 (N_18499,N_17438,N_17713);
nor U18500 (N_18500,N_17553,N_17062);
or U18501 (N_18501,N_17920,N_17845);
nor U18502 (N_18502,N_17548,N_17552);
or U18503 (N_18503,N_17195,N_17834);
or U18504 (N_18504,N_17165,N_17265);
nand U18505 (N_18505,N_17726,N_17815);
or U18506 (N_18506,N_17136,N_17144);
nor U18507 (N_18507,N_17400,N_17425);
or U18508 (N_18508,N_17921,N_17994);
nor U18509 (N_18509,N_17996,N_17229);
nand U18510 (N_18510,N_17847,N_17146);
xor U18511 (N_18511,N_17137,N_17335);
and U18512 (N_18512,N_17867,N_17509);
xnor U18513 (N_18513,N_17549,N_17095);
nor U18514 (N_18514,N_17927,N_17898);
nand U18515 (N_18515,N_17544,N_17832);
and U18516 (N_18516,N_17099,N_17742);
xnor U18517 (N_18517,N_17501,N_17608);
xor U18518 (N_18518,N_17352,N_17895);
and U18519 (N_18519,N_17774,N_17132);
nand U18520 (N_18520,N_17280,N_17237);
nor U18521 (N_18521,N_17610,N_17570);
or U18522 (N_18522,N_17109,N_17081);
and U18523 (N_18523,N_17109,N_17718);
or U18524 (N_18524,N_17172,N_17420);
or U18525 (N_18525,N_17111,N_17898);
nand U18526 (N_18526,N_17238,N_17868);
xnor U18527 (N_18527,N_17216,N_17433);
or U18528 (N_18528,N_17755,N_17438);
or U18529 (N_18529,N_17408,N_17106);
and U18530 (N_18530,N_17968,N_17590);
nand U18531 (N_18531,N_17754,N_17840);
xnor U18532 (N_18532,N_17076,N_17037);
xnor U18533 (N_18533,N_17064,N_17036);
nand U18534 (N_18534,N_17123,N_17477);
or U18535 (N_18535,N_17404,N_17726);
and U18536 (N_18536,N_17500,N_17827);
nor U18537 (N_18537,N_17614,N_17706);
and U18538 (N_18538,N_17908,N_17825);
xor U18539 (N_18539,N_17979,N_17121);
and U18540 (N_18540,N_17640,N_17996);
nor U18541 (N_18541,N_17982,N_17301);
xnor U18542 (N_18542,N_17924,N_17469);
xor U18543 (N_18543,N_17496,N_17004);
nor U18544 (N_18544,N_17489,N_17837);
xor U18545 (N_18545,N_17173,N_17719);
nand U18546 (N_18546,N_17956,N_17554);
nor U18547 (N_18547,N_17528,N_17027);
or U18548 (N_18548,N_17723,N_17011);
or U18549 (N_18549,N_17692,N_17698);
and U18550 (N_18550,N_17431,N_17512);
nor U18551 (N_18551,N_17245,N_17725);
and U18552 (N_18552,N_17253,N_17873);
nor U18553 (N_18553,N_17945,N_17231);
nor U18554 (N_18554,N_17977,N_17393);
nand U18555 (N_18555,N_17326,N_17906);
and U18556 (N_18556,N_17731,N_17750);
and U18557 (N_18557,N_17946,N_17807);
xor U18558 (N_18558,N_17733,N_17851);
nor U18559 (N_18559,N_17972,N_17797);
or U18560 (N_18560,N_17178,N_17053);
nand U18561 (N_18561,N_17648,N_17979);
and U18562 (N_18562,N_17367,N_17860);
xnor U18563 (N_18563,N_17781,N_17860);
nor U18564 (N_18564,N_17036,N_17832);
or U18565 (N_18565,N_17396,N_17547);
or U18566 (N_18566,N_17358,N_17834);
and U18567 (N_18567,N_17989,N_17855);
nor U18568 (N_18568,N_17413,N_17895);
xor U18569 (N_18569,N_17247,N_17498);
xnor U18570 (N_18570,N_17755,N_17002);
nor U18571 (N_18571,N_17376,N_17980);
or U18572 (N_18572,N_17691,N_17794);
nor U18573 (N_18573,N_17096,N_17702);
xnor U18574 (N_18574,N_17304,N_17357);
or U18575 (N_18575,N_17121,N_17417);
xnor U18576 (N_18576,N_17741,N_17712);
nand U18577 (N_18577,N_17557,N_17141);
xnor U18578 (N_18578,N_17921,N_17746);
nor U18579 (N_18579,N_17441,N_17419);
or U18580 (N_18580,N_17584,N_17238);
nor U18581 (N_18581,N_17557,N_17657);
or U18582 (N_18582,N_17814,N_17612);
nand U18583 (N_18583,N_17250,N_17057);
nor U18584 (N_18584,N_17489,N_17654);
or U18585 (N_18585,N_17482,N_17296);
nand U18586 (N_18586,N_17865,N_17100);
nor U18587 (N_18587,N_17269,N_17705);
or U18588 (N_18588,N_17755,N_17178);
and U18589 (N_18589,N_17903,N_17764);
nand U18590 (N_18590,N_17942,N_17285);
xnor U18591 (N_18591,N_17332,N_17338);
nand U18592 (N_18592,N_17713,N_17450);
nor U18593 (N_18593,N_17133,N_17160);
nand U18594 (N_18594,N_17351,N_17296);
nor U18595 (N_18595,N_17295,N_17017);
nand U18596 (N_18596,N_17776,N_17199);
xor U18597 (N_18597,N_17841,N_17411);
nand U18598 (N_18598,N_17627,N_17491);
xnor U18599 (N_18599,N_17606,N_17736);
nor U18600 (N_18600,N_17158,N_17751);
nor U18601 (N_18601,N_17841,N_17401);
xnor U18602 (N_18602,N_17203,N_17572);
or U18603 (N_18603,N_17217,N_17855);
and U18604 (N_18604,N_17258,N_17738);
nand U18605 (N_18605,N_17803,N_17790);
nand U18606 (N_18606,N_17297,N_17113);
xnor U18607 (N_18607,N_17841,N_17149);
and U18608 (N_18608,N_17326,N_17313);
and U18609 (N_18609,N_17414,N_17387);
xor U18610 (N_18610,N_17456,N_17448);
nor U18611 (N_18611,N_17404,N_17874);
nor U18612 (N_18612,N_17444,N_17666);
nand U18613 (N_18613,N_17615,N_17879);
or U18614 (N_18614,N_17569,N_17124);
xor U18615 (N_18615,N_17247,N_17547);
nand U18616 (N_18616,N_17970,N_17816);
nor U18617 (N_18617,N_17277,N_17712);
nand U18618 (N_18618,N_17374,N_17921);
nand U18619 (N_18619,N_17560,N_17512);
xor U18620 (N_18620,N_17701,N_17477);
nor U18621 (N_18621,N_17629,N_17312);
nor U18622 (N_18622,N_17864,N_17755);
or U18623 (N_18623,N_17872,N_17025);
and U18624 (N_18624,N_17385,N_17870);
or U18625 (N_18625,N_17590,N_17276);
and U18626 (N_18626,N_17255,N_17461);
or U18627 (N_18627,N_17092,N_17388);
or U18628 (N_18628,N_17950,N_17994);
and U18629 (N_18629,N_17413,N_17098);
and U18630 (N_18630,N_17468,N_17353);
nand U18631 (N_18631,N_17512,N_17425);
and U18632 (N_18632,N_17967,N_17807);
nor U18633 (N_18633,N_17968,N_17641);
nand U18634 (N_18634,N_17692,N_17932);
nand U18635 (N_18635,N_17786,N_17738);
xor U18636 (N_18636,N_17447,N_17101);
and U18637 (N_18637,N_17364,N_17819);
and U18638 (N_18638,N_17556,N_17477);
nor U18639 (N_18639,N_17231,N_17877);
or U18640 (N_18640,N_17535,N_17187);
nor U18641 (N_18641,N_17733,N_17483);
and U18642 (N_18642,N_17522,N_17431);
nor U18643 (N_18643,N_17479,N_17054);
or U18644 (N_18644,N_17531,N_17583);
xnor U18645 (N_18645,N_17749,N_17798);
xor U18646 (N_18646,N_17366,N_17748);
xor U18647 (N_18647,N_17495,N_17927);
and U18648 (N_18648,N_17981,N_17692);
or U18649 (N_18649,N_17186,N_17078);
or U18650 (N_18650,N_17926,N_17887);
xor U18651 (N_18651,N_17285,N_17223);
xnor U18652 (N_18652,N_17901,N_17138);
or U18653 (N_18653,N_17897,N_17920);
xor U18654 (N_18654,N_17005,N_17667);
nand U18655 (N_18655,N_17802,N_17676);
or U18656 (N_18656,N_17920,N_17604);
or U18657 (N_18657,N_17142,N_17848);
nor U18658 (N_18658,N_17133,N_17083);
or U18659 (N_18659,N_17907,N_17318);
and U18660 (N_18660,N_17777,N_17551);
nand U18661 (N_18661,N_17163,N_17193);
and U18662 (N_18662,N_17498,N_17928);
and U18663 (N_18663,N_17566,N_17370);
or U18664 (N_18664,N_17304,N_17493);
nand U18665 (N_18665,N_17190,N_17318);
nand U18666 (N_18666,N_17269,N_17696);
nand U18667 (N_18667,N_17149,N_17809);
and U18668 (N_18668,N_17675,N_17853);
nor U18669 (N_18669,N_17462,N_17781);
xnor U18670 (N_18670,N_17118,N_17961);
nand U18671 (N_18671,N_17933,N_17241);
xnor U18672 (N_18672,N_17290,N_17988);
nand U18673 (N_18673,N_17618,N_17694);
nand U18674 (N_18674,N_17420,N_17152);
xor U18675 (N_18675,N_17478,N_17456);
xor U18676 (N_18676,N_17578,N_17047);
nand U18677 (N_18677,N_17826,N_17431);
nor U18678 (N_18678,N_17992,N_17635);
nor U18679 (N_18679,N_17747,N_17607);
and U18680 (N_18680,N_17740,N_17817);
nor U18681 (N_18681,N_17672,N_17439);
or U18682 (N_18682,N_17795,N_17858);
or U18683 (N_18683,N_17800,N_17825);
xnor U18684 (N_18684,N_17564,N_17263);
xor U18685 (N_18685,N_17608,N_17744);
nand U18686 (N_18686,N_17002,N_17416);
or U18687 (N_18687,N_17270,N_17159);
or U18688 (N_18688,N_17981,N_17882);
or U18689 (N_18689,N_17202,N_17679);
nand U18690 (N_18690,N_17520,N_17997);
and U18691 (N_18691,N_17134,N_17820);
nor U18692 (N_18692,N_17061,N_17120);
xor U18693 (N_18693,N_17133,N_17903);
nor U18694 (N_18694,N_17308,N_17128);
nor U18695 (N_18695,N_17292,N_17337);
xor U18696 (N_18696,N_17838,N_17520);
or U18697 (N_18697,N_17885,N_17063);
xnor U18698 (N_18698,N_17857,N_17548);
and U18699 (N_18699,N_17615,N_17188);
xnor U18700 (N_18700,N_17250,N_17976);
or U18701 (N_18701,N_17001,N_17334);
nor U18702 (N_18702,N_17599,N_17441);
xnor U18703 (N_18703,N_17135,N_17503);
and U18704 (N_18704,N_17870,N_17111);
xor U18705 (N_18705,N_17216,N_17719);
and U18706 (N_18706,N_17456,N_17730);
or U18707 (N_18707,N_17816,N_17776);
nand U18708 (N_18708,N_17650,N_17544);
xnor U18709 (N_18709,N_17821,N_17845);
nor U18710 (N_18710,N_17569,N_17159);
xor U18711 (N_18711,N_17982,N_17581);
xor U18712 (N_18712,N_17288,N_17537);
xor U18713 (N_18713,N_17677,N_17259);
xnor U18714 (N_18714,N_17676,N_17813);
xor U18715 (N_18715,N_17583,N_17243);
nor U18716 (N_18716,N_17822,N_17847);
xor U18717 (N_18717,N_17223,N_17778);
nand U18718 (N_18718,N_17042,N_17674);
and U18719 (N_18719,N_17191,N_17959);
nand U18720 (N_18720,N_17542,N_17083);
or U18721 (N_18721,N_17240,N_17764);
or U18722 (N_18722,N_17072,N_17203);
nor U18723 (N_18723,N_17453,N_17473);
nor U18724 (N_18724,N_17904,N_17184);
nor U18725 (N_18725,N_17640,N_17325);
nor U18726 (N_18726,N_17151,N_17925);
nor U18727 (N_18727,N_17247,N_17710);
and U18728 (N_18728,N_17563,N_17714);
nand U18729 (N_18729,N_17862,N_17328);
nor U18730 (N_18730,N_17838,N_17213);
xnor U18731 (N_18731,N_17417,N_17631);
xor U18732 (N_18732,N_17517,N_17657);
or U18733 (N_18733,N_17481,N_17030);
nand U18734 (N_18734,N_17441,N_17880);
or U18735 (N_18735,N_17845,N_17003);
xnor U18736 (N_18736,N_17946,N_17610);
nand U18737 (N_18737,N_17408,N_17820);
nand U18738 (N_18738,N_17870,N_17499);
xnor U18739 (N_18739,N_17583,N_17917);
xor U18740 (N_18740,N_17462,N_17025);
and U18741 (N_18741,N_17007,N_17296);
nor U18742 (N_18742,N_17301,N_17834);
and U18743 (N_18743,N_17362,N_17536);
nand U18744 (N_18744,N_17307,N_17704);
nor U18745 (N_18745,N_17264,N_17671);
xnor U18746 (N_18746,N_17445,N_17603);
or U18747 (N_18747,N_17153,N_17083);
nor U18748 (N_18748,N_17705,N_17711);
nand U18749 (N_18749,N_17112,N_17095);
xnor U18750 (N_18750,N_17443,N_17303);
and U18751 (N_18751,N_17701,N_17394);
and U18752 (N_18752,N_17414,N_17727);
nor U18753 (N_18753,N_17682,N_17860);
nand U18754 (N_18754,N_17871,N_17076);
and U18755 (N_18755,N_17940,N_17534);
and U18756 (N_18756,N_17727,N_17515);
nand U18757 (N_18757,N_17405,N_17356);
nand U18758 (N_18758,N_17020,N_17976);
or U18759 (N_18759,N_17708,N_17913);
nor U18760 (N_18760,N_17750,N_17985);
or U18761 (N_18761,N_17817,N_17179);
xor U18762 (N_18762,N_17046,N_17404);
nor U18763 (N_18763,N_17485,N_17149);
nand U18764 (N_18764,N_17616,N_17153);
or U18765 (N_18765,N_17448,N_17724);
nand U18766 (N_18766,N_17668,N_17397);
nand U18767 (N_18767,N_17722,N_17855);
and U18768 (N_18768,N_17856,N_17678);
and U18769 (N_18769,N_17388,N_17669);
nor U18770 (N_18770,N_17464,N_17073);
xor U18771 (N_18771,N_17625,N_17031);
nand U18772 (N_18772,N_17646,N_17254);
nor U18773 (N_18773,N_17407,N_17455);
nor U18774 (N_18774,N_17538,N_17101);
or U18775 (N_18775,N_17009,N_17977);
and U18776 (N_18776,N_17466,N_17139);
nor U18777 (N_18777,N_17142,N_17763);
and U18778 (N_18778,N_17203,N_17787);
xor U18779 (N_18779,N_17548,N_17230);
or U18780 (N_18780,N_17185,N_17844);
nor U18781 (N_18781,N_17370,N_17518);
xor U18782 (N_18782,N_17288,N_17354);
xor U18783 (N_18783,N_17865,N_17146);
nor U18784 (N_18784,N_17859,N_17252);
nand U18785 (N_18785,N_17797,N_17871);
nor U18786 (N_18786,N_17546,N_17311);
or U18787 (N_18787,N_17459,N_17803);
or U18788 (N_18788,N_17403,N_17659);
xor U18789 (N_18789,N_17362,N_17541);
or U18790 (N_18790,N_17262,N_17914);
and U18791 (N_18791,N_17699,N_17295);
nand U18792 (N_18792,N_17393,N_17605);
or U18793 (N_18793,N_17054,N_17152);
nand U18794 (N_18794,N_17306,N_17073);
nor U18795 (N_18795,N_17180,N_17987);
nand U18796 (N_18796,N_17066,N_17549);
nand U18797 (N_18797,N_17959,N_17543);
nor U18798 (N_18798,N_17290,N_17407);
or U18799 (N_18799,N_17752,N_17597);
nand U18800 (N_18800,N_17417,N_17324);
and U18801 (N_18801,N_17103,N_17879);
nand U18802 (N_18802,N_17178,N_17064);
xnor U18803 (N_18803,N_17143,N_17089);
and U18804 (N_18804,N_17843,N_17948);
nand U18805 (N_18805,N_17744,N_17181);
and U18806 (N_18806,N_17187,N_17683);
nor U18807 (N_18807,N_17218,N_17067);
nor U18808 (N_18808,N_17052,N_17781);
or U18809 (N_18809,N_17027,N_17306);
nor U18810 (N_18810,N_17847,N_17292);
nor U18811 (N_18811,N_17158,N_17120);
or U18812 (N_18812,N_17666,N_17782);
xnor U18813 (N_18813,N_17937,N_17733);
xnor U18814 (N_18814,N_17024,N_17105);
and U18815 (N_18815,N_17592,N_17658);
xor U18816 (N_18816,N_17287,N_17477);
nor U18817 (N_18817,N_17691,N_17004);
nand U18818 (N_18818,N_17052,N_17099);
or U18819 (N_18819,N_17119,N_17519);
and U18820 (N_18820,N_17349,N_17457);
nand U18821 (N_18821,N_17112,N_17514);
nor U18822 (N_18822,N_17836,N_17200);
or U18823 (N_18823,N_17361,N_17325);
nand U18824 (N_18824,N_17728,N_17147);
nor U18825 (N_18825,N_17436,N_17071);
nand U18826 (N_18826,N_17126,N_17573);
nand U18827 (N_18827,N_17460,N_17166);
nand U18828 (N_18828,N_17160,N_17729);
or U18829 (N_18829,N_17969,N_17990);
nor U18830 (N_18830,N_17993,N_17572);
nand U18831 (N_18831,N_17211,N_17429);
xnor U18832 (N_18832,N_17898,N_17778);
nor U18833 (N_18833,N_17514,N_17666);
nor U18834 (N_18834,N_17675,N_17576);
nor U18835 (N_18835,N_17019,N_17644);
and U18836 (N_18836,N_17677,N_17749);
or U18837 (N_18837,N_17449,N_17053);
and U18838 (N_18838,N_17253,N_17186);
and U18839 (N_18839,N_17967,N_17335);
and U18840 (N_18840,N_17349,N_17488);
or U18841 (N_18841,N_17212,N_17975);
and U18842 (N_18842,N_17184,N_17655);
xnor U18843 (N_18843,N_17263,N_17305);
and U18844 (N_18844,N_17235,N_17416);
nand U18845 (N_18845,N_17740,N_17487);
and U18846 (N_18846,N_17977,N_17757);
and U18847 (N_18847,N_17267,N_17740);
nand U18848 (N_18848,N_17826,N_17251);
xor U18849 (N_18849,N_17676,N_17750);
and U18850 (N_18850,N_17984,N_17197);
nand U18851 (N_18851,N_17381,N_17776);
and U18852 (N_18852,N_17516,N_17661);
nor U18853 (N_18853,N_17026,N_17083);
and U18854 (N_18854,N_17688,N_17875);
xnor U18855 (N_18855,N_17429,N_17964);
or U18856 (N_18856,N_17981,N_17526);
and U18857 (N_18857,N_17585,N_17404);
or U18858 (N_18858,N_17690,N_17991);
nand U18859 (N_18859,N_17288,N_17252);
and U18860 (N_18860,N_17115,N_17167);
nor U18861 (N_18861,N_17613,N_17654);
or U18862 (N_18862,N_17830,N_17113);
nand U18863 (N_18863,N_17915,N_17854);
and U18864 (N_18864,N_17843,N_17645);
or U18865 (N_18865,N_17423,N_17861);
or U18866 (N_18866,N_17456,N_17995);
or U18867 (N_18867,N_17729,N_17462);
xnor U18868 (N_18868,N_17022,N_17173);
and U18869 (N_18869,N_17859,N_17742);
xnor U18870 (N_18870,N_17439,N_17779);
and U18871 (N_18871,N_17580,N_17841);
nand U18872 (N_18872,N_17285,N_17161);
nor U18873 (N_18873,N_17639,N_17873);
and U18874 (N_18874,N_17032,N_17404);
and U18875 (N_18875,N_17126,N_17691);
and U18876 (N_18876,N_17914,N_17955);
or U18877 (N_18877,N_17260,N_17726);
or U18878 (N_18878,N_17511,N_17548);
nor U18879 (N_18879,N_17157,N_17299);
or U18880 (N_18880,N_17468,N_17316);
or U18881 (N_18881,N_17345,N_17142);
or U18882 (N_18882,N_17064,N_17660);
xor U18883 (N_18883,N_17687,N_17754);
xor U18884 (N_18884,N_17707,N_17453);
or U18885 (N_18885,N_17885,N_17210);
or U18886 (N_18886,N_17973,N_17691);
nand U18887 (N_18887,N_17305,N_17389);
nor U18888 (N_18888,N_17047,N_17412);
nand U18889 (N_18889,N_17557,N_17177);
nand U18890 (N_18890,N_17519,N_17771);
xnor U18891 (N_18891,N_17958,N_17528);
xor U18892 (N_18892,N_17634,N_17891);
nand U18893 (N_18893,N_17869,N_17073);
and U18894 (N_18894,N_17472,N_17572);
nand U18895 (N_18895,N_17623,N_17940);
and U18896 (N_18896,N_17812,N_17973);
or U18897 (N_18897,N_17332,N_17148);
nor U18898 (N_18898,N_17661,N_17730);
nor U18899 (N_18899,N_17983,N_17287);
or U18900 (N_18900,N_17202,N_17135);
or U18901 (N_18901,N_17188,N_17192);
or U18902 (N_18902,N_17884,N_17168);
and U18903 (N_18903,N_17281,N_17919);
and U18904 (N_18904,N_17128,N_17844);
nand U18905 (N_18905,N_17430,N_17656);
and U18906 (N_18906,N_17296,N_17698);
xnor U18907 (N_18907,N_17237,N_17557);
nor U18908 (N_18908,N_17304,N_17098);
nand U18909 (N_18909,N_17193,N_17258);
nand U18910 (N_18910,N_17174,N_17323);
or U18911 (N_18911,N_17611,N_17992);
xnor U18912 (N_18912,N_17502,N_17538);
or U18913 (N_18913,N_17770,N_17460);
nor U18914 (N_18914,N_17507,N_17557);
xor U18915 (N_18915,N_17834,N_17786);
nand U18916 (N_18916,N_17253,N_17555);
nand U18917 (N_18917,N_17989,N_17976);
nor U18918 (N_18918,N_17387,N_17096);
xnor U18919 (N_18919,N_17317,N_17422);
and U18920 (N_18920,N_17141,N_17291);
or U18921 (N_18921,N_17865,N_17166);
xor U18922 (N_18922,N_17537,N_17507);
xnor U18923 (N_18923,N_17942,N_17040);
or U18924 (N_18924,N_17907,N_17532);
or U18925 (N_18925,N_17011,N_17267);
nand U18926 (N_18926,N_17562,N_17490);
nand U18927 (N_18927,N_17557,N_17199);
or U18928 (N_18928,N_17830,N_17242);
nand U18929 (N_18929,N_17526,N_17022);
and U18930 (N_18930,N_17137,N_17034);
xnor U18931 (N_18931,N_17205,N_17433);
nor U18932 (N_18932,N_17412,N_17480);
nor U18933 (N_18933,N_17055,N_17509);
and U18934 (N_18934,N_17785,N_17360);
nor U18935 (N_18935,N_17463,N_17225);
nor U18936 (N_18936,N_17601,N_17668);
and U18937 (N_18937,N_17143,N_17011);
xor U18938 (N_18938,N_17476,N_17251);
nor U18939 (N_18939,N_17270,N_17320);
nor U18940 (N_18940,N_17466,N_17570);
xnor U18941 (N_18941,N_17268,N_17966);
xor U18942 (N_18942,N_17061,N_17664);
and U18943 (N_18943,N_17469,N_17596);
or U18944 (N_18944,N_17260,N_17887);
and U18945 (N_18945,N_17185,N_17521);
nand U18946 (N_18946,N_17519,N_17931);
xor U18947 (N_18947,N_17042,N_17030);
xor U18948 (N_18948,N_17524,N_17930);
xnor U18949 (N_18949,N_17514,N_17886);
or U18950 (N_18950,N_17415,N_17988);
and U18951 (N_18951,N_17724,N_17001);
nand U18952 (N_18952,N_17443,N_17630);
or U18953 (N_18953,N_17274,N_17521);
or U18954 (N_18954,N_17257,N_17112);
xor U18955 (N_18955,N_17369,N_17597);
nand U18956 (N_18956,N_17323,N_17114);
nand U18957 (N_18957,N_17933,N_17174);
xnor U18958 (N_18958,N_17386,N_17482);
nand U18959 (N_18959,N_17277,N_17507);
nand U18960 (N_18960,N_17572,N_17890);
or U18961 (N_18961,N_17984,N_17388);
or U18962 (N_18962,N_17785,N_17324);
and U18963 (N_18963,N_17283,N_17797);
or U18964 (N_18964,N_17680,N_17549);
or U18965 (N_18965,N_17179,N_17474);
and U18966 (N_18966,N_17001,N_17983);
xnor U18967 (N_18967,N_17406,N_17433);
and U18968 (N_18968,N_17765,N_17784);
nor U18969 (N_18969,N_17039,N_17466);
or U18970 (N_18970,N_17393,N_17367);
or U18971 (N_18971,N_17934,N_17908);
or U18972 (N_18972,N_17126,N_17815);
xnor U18973 (N_18973,N_17344,N_17454);
and U18974 (N_18974,N_17583,N_17043);
or U18975 (N_18975,N_17960,N_17682);
and U18976 (N_18976,N_17266,N_17950);
or U18977 (N_18977,N_17947,N_17173);
xnor U18978 (N_18978,N_17260,N_17010);
or U18979 (N_18979,N_17879,N_17412);
xnor U18980 (N_18980,N_17983,N_17043);
nand U18981 (N_18981,N_17822,N_17807);
nand U18982 (N_18982,N_17144,N_17677);
or U18983 (N_18983,N_17641,N_17853);
and U18984 (N_18984,N_17700,N_17371);
xnor U18985 (N_18985,N_17820,N_17383);
xnor U18986 (N_18986,N_17627,N_17236);
xor U18987 (N_18987,N_17501,N_17677);
nor U18988 (N_18988,N_17444,N_17847);
and U18989 (N_18989,N_17083,N_17759);
nor U18990 (N_18990,N_17613,N_17932);
xor U18991 (N_18991,N_17777,N_17681);
and U18992 (N_18992,N_17928,N_17707);
nand U18993 (N_18993,N_17983,N_17675);
nor U18994 (N_18994,N_17395,N_17171);
nand U18995 (N_18995,N_17464,N_17743);
nand U18996 (N_18996,N_17581,N_17478);
nand U18997 (N_18997,N_17047,N_17647);
xnor U18998 (N_18998,N_17239,N_17426);
nor U18999 (N_18999,N_17029,N_17014);
nand U19000 (N_19000,N_18371,N_18928);
nand U19001 (N_19001,N_18091,N_18430);
and U19002 (N_19002,N_18609,N_18744);
nand U19003 (N_19003,N_18625,N_18965);
xnor U19004 (N_19004,N_18844,N_18575);
nand U19005 (N_19005,N_18900,N_18251);
nor U19006 (N_19006,N_18315,N_18276);
nor U19007 (N_19007,N_18878,N_18895);
nor U19008 (N_19008,N_18010,N_18016);
xnor U19009 (N_19009,N_18760,N_18946);
and U19010 (N_19010,N_18616,N_18492);
nor U19011 (N_19011,N_18327,N_18559);
nand U19012 (N_19012,N_18057,N_18097);
nor U19013 (N_19013,N_18979,N_18051);
and U19014 (N_19014,N_18291,N_18821);
nand U19015 (N_19015,N_18996,N_18148);
and U19016 (N_19016,N_18254,N_18817);
or U19017 (N_19017,N_18932,N_18083);
nor U19018 (N_19018,N_18574,N_18494);
and U19019 (N_19019,N_18506,N_18324);
or U19020 (N_19020,N_18295,N_18673);
nor U19021 (N_19021,N_18423,N_18269);
nor U19022 (N_19022,N_18508,N_18600);
nor U19023 (N_19023,N_18582,N_18432);
nor U19024 (N_19024,N_18724,N_18725);
or U19025 (N_19025,N_18563,N_18047);
nand U19026 (N_19026,N_18300,N_18845);
or U19027 (N_19027,N_18059,N_18759);
or U19028 (N_19028,N_18524,N_18119);
and U19029 (N_19029,N_18617,N_18546);
xor U19030 (N_19030,N_18282,N_18386);
nor U19031 (N_19031,N_18527,N_18024);
and U19032 (N_19032,N_18342,N_18606);
or U19033 (N_19033,N_18970,N_18983);
and U19034 (N_19034,N_18861,N_18081);
nand U19035 (N_19035,N_18767,N_18816);
or U19036 (N_19036,N_18168,N_18299);
nand U19037 (N_19037,N_18104,N_18581);
nor U19038 (N_19038,N_18444,N_18095);
nand U19039 (N_19039,N_18381,N_18441);
xnor U19040 (N_19040,N_18783,N_18820);
nand U19041 (N_19041,N_18473,N_18482);
or U19042 (N_19042,N_18337,N_18653);
nand U19043 (N_19043,N_18287,N_18583);
or U19044 (N_19044,N_18485,N_18311);
nor U19045 (N_19045,N_18697,N_18252);
or U19046 (N_19046,N_18171,N_18328);
or U19047 (N_19047,N_18781,N_18864);
nor U19048 (N_19048,N_18383,N_18340);
or U19049 (N_19049,N_18294,N_18636);
nor U19050 (N_19050,N_18692,N_18859);
xnor U19051 (N_19051,N_18448,N_18666);
and U19052 (N_19052,N_18174,N_18776);
nand U19053 (N_19053,N_18756,N_18854);
and U19054 (N_19054,N_18825,N_18812);
nor U19055 (N_19055,N_18314,N_18105);
and U19056 (N_19056,N_18195,N_18493);
nand U19057 (N_19057,N_18215,N_18253);
nand U19058 (N_19058,N_18380,N_18985);
nand U19059 (N_19059,N_18769,N_18296);
and U19060 (N_19060,N_18480,N_18657);
nand U19061 (N_19061,N_18784,N_18586);
nor U19062 (N_19062,N_18398,N_18664);
nand U19063 (N_19063,N_18579,N_18084);
or U19064 (N_19064,N_18947,N_18554);
or U19065 (N_19065,N_18108,N_18391);
nand U19066 (N_19066,N_18570,N_18860);
and U19067 (N_19067,N_18793,N_18916);
nand U19068 (N_19068,N_18421,N_18800);
xnor U19069 (N_19069,N_18213,N_18457);
and U19070 (N_19070,N_18612,N_18778);
nand U19071 (N_19071,N_18555,N_18607);
nand U19072 (N_19072,N_18735,N_18824);
nor U19073 (N_19073,N_18250,N_18741);
nor U19074 (N_19074,N_18367,N_18331);
or U19075 (N_19075,N_18856,N_18663);
or U19076 (N_19076,N_18443,N_18445);
nor U19077 (N_19077,N_18087,N_18733);
xor U19078 (N_19078,N_18220,N_18597);
nand U19079 (N_19079,N_18159,N_18308);
and U19080 (N_19080,N_18541,N_18561);
nand U19081 (N_19081,N_18855,N_18833);
or U19082 (N_19082,N_18207,N_18941);
or U19083 (N_19083,N_18446,N_18001);
nor U19084 (N_19084,N_18536,N_18644);
or U19085 (N_19085,N_18066,N_18124);
or U19086 (N_19086,N_18523,N_18713);
nand U19087 (N_19087,N_18894,N_18232);
and U19088 (N_19088,N_18418,N_18803);
xor U19089 (N_19089,N_18992,N_18533);
and U19090 (N_19090,N_18486,N_18734);
nor U19091 (N_19091,N_18588,N_18209);
or U19092 (N_19092,N_18530,N_18834);
and U19093 (N_19093,N_18263,N_18632);
and U19094 (N_19094,N_18202,N_18236);
xor U19095 (N_19095,N_18819,N_18779);
and U19096 (N_19096,N_18519,N_18490);
nor U19097 (N_19097,N_18013,N_18801);
and U19098 (N_19098,N_18589,N_18477);
nor U19099 (N_19099,N_18931,N_18434);
and U19100 (N_19100,N_18545,N_18711);
or U19101 (N_19101,N_18788,N_18547);
and U19102 (N_19102,N_18284,N_18974);
or U19103 (N_19103,N_18576,N_18611);
and U19104 (N_19104,N_18699,N_18595);
nand U19105 (N_19105,N_18658,N_18136);
xor U19106 (N_19106,N_18361,N_18170);
nor U19107 (N_19107,N_18395,N_18447);
nand U19108 (N_19108,N_18599,N_18198);
xor U19109 (N_19109,N_18873,N_18815);
nand U19110 (N_19110,N_18412,N_18107);
nand U19111 (N_19111,N_18832,N_18027);
xnor U19112 (N_19112,N_18351,N_18223);
or U19113 (N_19113,N_18507,N_18939);
xor U19114 (N_19114,N_18046,N_18467);
xor U19115 (N_19115,N_18921,N_18101);
nor U19116 (N_19116,N_18392,N_18364);
and U19117 (N_19117,N_18610,N_18571);
or U19118 (N_19118,N_18596,N_18230);
nand U19119 (N_19119,N_18323,N_18375);
nor U19120 (N_19120,N_18354,N_18106);
nor U19121 (N_19121,N_18012,N_18238);
and U19122 (N_19122,N_18768,N_18488);
or U19123 (N_19123,N_18811,N_18481);
nor U19124 (N_19124,N_18189,N_18092);
nand U19125 (N_19125,N_18660,N_18665);
and U19126 (N_19126,N_18671,N_18905);
nor U19127 (N_19127,N_18316,N_18293);
or U19128 (N_19128,N_18693,N_18133);
nor U19129 (N_19129,N_18054,N_18401);
nor U19130 (N_19130,N_18828,N_18872);
nand U19131 (N_19131,N_18281,N_18991);
and U19132 (N_19132,N_18157,N_18764);
xor U19133 (N_19133,N_18370,N_18649);
xor U19134 (N_19134,N_18417,N_18021);
and U19135 (N_19135,N_18100,N_18397);
nor U19136 (N_19136,N_18036,N_18917);
nor U19137 (N_19137,N_18376,N_18030);
nand U19138 (N_19138,N_18339,N_18898);
and U19139 (N_19139,N_18466,N_18901);
or U19140 (N_19140,N_18479,N_18216);
or U19141 (N_19141,N_18273,N_18149);
or U19142 (N_19142,N_18063,N_18453);
and U19143 (N_19143,N_18078,N_18516);
xnor U19144 (N_19144,N_18848,N_18651);
or U19145 (N_19145,N_18422,N_18019);
and U19146 (N_19146,N_18736,N_18972);
or U19147 (N_19147,N_18987,N_18163);
xnor U19148 (N_19148,N_18256,N_18279);
or U19149 (N_19149,N_18079,N_18224);
xor U19150 (N_19150,N_18850,N_18710);
nor U19151 (N_19151,N_18259,N_18694);
and U19152 (N_19152,N_18652,N_18961);
nand U19153 (N_19153,N_18714,N_18838);
xnor U19154 (N_19154,N_18945,N_18166);
xnor U19155 (N_19155,N_18025,N_18359);
nor U19156 (N_19156,N_18302,N_18085);
xnor U19157 (N_19157,N_18716,N_18912);
nand U19158 (N_19158,N_18454,N_18957);
nand U19159 (N_19159,N_18967,N_18204);
nor U19160 (N_19160,N_18067,N_18627);
or U19161 (N_19161,N_18678,N_18491);
or U19162 (N_19162,N_18497,N_18004);
xnor U19163 (N_19163,N_18145,N_18071);
xor U19164 (N_19164,N_18086,N_18818);
nor U19165 (N_19165,N_18601,N_18379);
nor U19166 (N_19166,N_18060,N_18357);
xnor U19167 (N_19167,N_18283,N_18667);
or U19168 (N_19168,N_18053,N_18048);
nand U19169 (N_19169,N_18999,N_18470);
xnor U19170 (N_19170,N_18109,N_18326);
nor U19171 (N_19171,N_18280,N_18366);
and U19172 (N_19172,N_18984,N_18998);
xnor U19173 (N_19173,N_18867,N_18404);
or U19174 (N_19174,N_18312,N_18355);
nor U19175 (N_19175,N_18330,N_18676);
nor U19176 (N_19176,N_18722,N_18709);
nand U19177 (N_19177,N_18126,N_18313);
nand U19178 (N_19178,N_18303,N_18245);
nand U19179 (N_19179,N_18499,N_18566);
or U19180 (N_19180,N_18933,N_18420);
xor U19181 (N_19181,N_18790,N_18520);
nand U19182 (N_19182,N_18304,N_18691);
nor U19183 (N_19183,N_18502,N_18843);
nor U19184 (N_19184,N_18997,N_18640);
and U19185 (N_19185,N_18911,N_18161);
nand U19186 (N_19186,N_18510,N_18680);
xor U19187 (N_19187,N_18322,N_18737);
and U19188 (N_19188,N_18474,N_18750);
nand U19189 (N_19189,N_18023,N_18943);
and U19190 (N_19190,N_18222,N_18246);
xor U19191 (N_19191,N_18462,N_18436);
nor U19192 (N_19192,N_18270,N_18573);
and U19193 (N_19193,N_18630,N_18118);
nor U19194 (N_19194,N_18853,N_18289);
xor U19195 (N_19195,N_18730,N_18435);
and U19196 (N_19196,N_18405,N_18968);
nand U19197 (N_19197,N_18647,N_18064);
xnor U19198 (N_19198,N_18568,N_18746);
xor U19199 (N_19199,N_18829,N_18178);
nor U19200 (N_19200,N_18385,N_18011);
nor U19201 (N_19201,N_18870,N_18602);
and U19202 (N_19202,N_18277,N_18766);
or U19203 (N_19203,N_18525,N_18152);
xor U19204 (N_19204,N_18134,N_18633);
xnor U19205 (N_19205,N_18000,N_18243);
xor U19206 (N_19206,N_18360,N_18188);
xnor U19207 (N_19207,N_18747,N_18622);
xor U19208 (N_19208,N_18840,N_18415);
nand U19209 (N_19209,N_18262,N_18061);
nor U19210 (N_19210,N_18585,N_18129);
xor U19211 (N_19211,N_18455,N_18286);
or U19212 (N_19212,N_18037,N_18431);
nand U19213 (N_19213,N_18637,N_18792);
and U19214 (N_19214,N_18478,N_18169);
nor U19215 (N_19215,N_18414,N_18836);
xor U19216 (N_19216,N_18908,N_18887);
xnor U19217 (N_19217,N_18701,N_18620);
and U19218 (N_19218,N_18955,N_18642);
or U19219 (N_19219,N_18549,N_18208);
or U19220 (N_19220,N_18973,N_18646);
nor U19221 (N_19221,N_18754,N_18924);
nand U19222 (N_19222,N_18785,N_18810);
and U19223 (N_19223,N_18706,N_18879);
and U19224 (N_19224,N_18338,N_18346);
xnor U19225 (N_19225,N_18677,N_18857);
nor U19226 (N_19226,N_18098,N_18876);
or U19227 (N_19227,N_18029,N_18411);
nand U19228 (N_19228,N_18298,N_18749);
xnor U19229 (N_19229,N_18951,N_18922);
or U19230 (N_19230,N_18413,N_18147);
nand U19231 (N_19231,N_18387,N_18088);
and U19232 (N_19232,N_18966,N_18685);
nor U19233 (N_19233,N_18969,N_18531);
and U19234 (N_19234,N_18073,N_18634);
or U19235 (N_19235,N_18669,N_18962);
xnor U19236 (N_19236,N_18892,N_18560);
nor U19237 (N_19237,N_18335,N_18442);
and U19238 (N_19238,N_18542,N_18723);
and U19239 (N_19239,N_18674,N_18696);
xnor U19240 (N_19240,N_18897,N_18039);
or U19241 (N_19241,N_18977,N_18613);
nor U19242 (N_19242,N_18799,N_18116);
nor U19243 (N_19243,N_18348,N_18052);
or U19244 (N_19244,N_18851,N_18180);
and U19245 (N_19245,N_18643,N_18082);
or U19246 (N_19246,N_18130,N_18437);
or U19247 (N_19247,N_18231,N_18007);
and U19248 (N_19248,N_18902,N_18650);
xor U19249 (N_19249,N_18191,N_18715);
nand U19250 (N_19250,N_18080,N_18858);
or U19251 (N_19251,N_18719,N_18952);
and U19252 (N_19252,N_18740,N_18654);
nor U19253 (N_19253,N_18459,N_18003);
nor U19254 (N_19254,N_18014,N_18112);
xor U19255 (N_19255,N_18700,N_18830);
and U19256 (N_19256,N_18707,N_18210);
nand U19257 (N_19257,N_18795,N_18672);
xor U19258 (N_19258,N_18518,N_18717);
and U19259 (N_19259,N_18475,N_18668);
xor U19260 (N_19260,N_18835,N_18074);
and U19261 (N_19261,N_18255,N_18242);
nand U19262 (N_19262,N_18628,N_18661);
nor U19263 (N_19263,N_18564,N_18089);
xnor U19264 (N_19264,N_18802,N_18374);
nand U19265 (N_19265,N_18009,N_18248);
and U19266 (N_19266,N_18639,N_18155);
or U19267 (N_19267,N_18028,N_18761);
nor U19268 (N_19268,N_18217,N_18350);
and U19269 (N_19269,N_18978,N_18496);
nand U19270 (N_19270,N_18131,N_18450);
and U19271 (N_19271,N_18020,N_18406);
or U19272 (N_19272,N_18621,N_18264);
or U19273 (N_19273,N_18940,N_18513);
or U19274 (N_19274,N_18509,N_18687);
xor U19275 (N_19275,N_18227,N_18988);
or U19276 (N_19276,N_18077,N_18923);
nor U19277 (N_19277,N_18142,N_18682);
nand U19278 (N_19278,N_18980,N_18150);
nor U19279 (N_19279,N_18846,N_18504);
nand U19280 (N_19280,N_18501,N_18199);
nand U19281 (N_19281,N_18827,N_18758);
xor U19282 (N_19282,N_18200,N_18537);
and U19283 (N_19283,N_18989,N_18805);
or U19284 (N_19284,N_18728,N_18698);
nand U19285 (N_19285,N_18772,N_18592);
and U19286 (N_19286,N_18102,N_18544);
and U19287 (N_19287,N_18393,N_18675);
or U19288 (N_19288,N_18317,N_18837);
nor U19289 (N_19289,N_18958,N_18512);
xor U19290 (N_19290,N_18813,N_18192);
nor U19291 (N_19291,N_18096,N_18689);
or U19292 (N_19292,N_18738,N_18156);
and U19293 (N_19293,N_18234,N_18786);
nor U19294 (N_19294,N_18241,N_18233);
nand U19295 (N_19295,N_18703,N_18852);
or U19296 (N_19296,N_18429,N_18938);
xnor U19297 (N_19297,N_18656,N_18890);
nand U19298 (N_19298,N_18343,N_18770);
xor U19299 (N_19299,N_18321,N_18110);
and U19300 (N_19300,N_18388,N_18272);
xnor U19301 (N_19301,N_18704,N_18796);
nand U19302 (N_19302,N_18594,N_18720);
or U19303 (N_19303,N_18789,N_18143);
or U19304 (N_19304,N_18742,N_18913);
and U19305 (N_19305,N_18993,N_18823);
xor U19306 (N_19306,N_18038,N_18033);
or U19307 (N_19307,N_18866,N_18569);
xor U19308 (N_19308,N_18261,N_18065);
and U19309 (N_19309,N_18167,N_18798);
and U19310 (N_19310,N_18604,N_18956);
and U19311 (N_19311,N_18521,N_18608);
xor U19312 (N_19312,N_18179,N_18505);
or U19313 (N_19313,N_18138,N_18954);
nor U19314 (N_19314,N_18886,N_18930);
xor U19315 (N_19315,N_18469,N_18182);
xor U19316 (N_19316,N_18146,N_18960);
nand U19317 (N_19317,N_18196,N_18266);
and U19318 (N_19318,N_18975,N_18184);
or U19319 (N_19319,N_18408,N_18572);
nor U19320 (N_19320,N_18718,N_18598);
nor U19321 (N_19321,N_18274,N_18584);
nand U19322 (N_19322,N_18807,N_18791);
xnor U19323 (N_19323,N_18702,N_18249);
nor U19324 (N_19324,N_18990,N_18229);
xnor U19325 (N_19325,N_18394,N_18183);
xor U19326 (N_19326,N_18528,N_18214);
and U19327 (N_19327,N_18212,N_18181);
nand U19328 (N_19328,N_18026,N_18522);
nor U19329 (N_19329,N_18449,N_18743);
and U19330 (N_19330,N_18885,N_18641);
or U19331 (N_19331,N_18031,N_18762);
xor U19332 (N_19332,N_18881,N_18319);
and U19333 (N_19333,N_18565,N_18332);
or U19334 (N_19334,N_18218,N_18944);
or U19335 (N_19335,N_18123,N_18333);
or U19336 (N_19336,N_18128,N_18305);
xnor U19337 (N_19337,N_18526,N_18219);
or U19338 (N_19338,N_18205,N_18550);
and U19339 (N_19339,N_18018,N_18440);
xor U19340 (N_19340,N_18139,N_18935);
or U19341 (N_19341,N_18919,N_18267);
nand U19342 (N_19342,N_18535,N_18041);
xor U19343 (N_19343,N_18164,N_18389);
and U19344 (N_19344,N_18648,N_18235);
and U19345 (N_19345,N_18534,N_18976);
nand U19346 (N_19346,N_18495,N_18301);
nand U19347 (N_19347,N_18655,N_18372);
and U19348 (N_19348,N_18880,N_18185);
xor U19349 (N_19349,N_18782,N_18117);
or U19350 (N_19350,N_18132,N_18377);
or U19351 (N_19351,N_18727,N_18726);
xnor U19352 (N_19352,N_18407,N_18175);
or U19353 (N_19353,N_18679,N_18538);
and U19354 (N_19354,N_18797,N_18099);
nor U19355 (N_19355,N_18552,N_18187);
nor U19356 (N_19356,N_18804,N_18578);
nand U19357 (N_19357,N_18461,N_18752);
nor U19358 (N_19358,N_18221,N_18907);
xor U19359 (N_19359,N_18847,N_18396);
nor U19360 (N_19360,N_18260,N_18426);
nand U19361 (N_19361,N_18684,N_18135);
nand U19362 (N_19362,N_18920,N_18540);
xnor U19363 (N_19363,N_18144,N_18986);
nor U19364 (N_19364,N_18058,N_18465);
nor U19365 (N_19365,N_18165,N_18695);
xnor U19366 (N_19366,N_18948,N_18731);
xnor U19367 (N_19367,N_18729,N_18751);
and U19368 (N_19368,N_18721,N_18732);
nand U19369 (N_19369,N_18822,N_18937);
nor U19370 (N_19370,N_18225,N_18439);
xnor U19371 (N_19371,N_18705,N_18265);
nor U19372 (N_19372,N_18580,N_18043);
xor U19373 (N_19373,N_18763,N_18556);
nand U19374 (N_19374,N_18925,N_18032);
or U19375 (N_19375,N_18121,N_18888);
or U19376 (N_19376,N_18472,N_18193);
or U19377 (N_19377,N_18757,N_18045);
xor U19378 (N_19378,N_18358,N_18874);
nor U19379 (N_19379,N_18329,N_18893);
or U19380 (N_19380,N_18949,N_18072);
nor U19381 (N_19381,N_18056,N_18950);
or U19382 (N_19382,N_18831,N_18275);
nor U19383 (N_19383,N_18120,N_18349);
or U19384 (N_19384,N_18140,N_18173);
or U19385 (N_19385,N_18906,N_18865);
xnor U19386 (N_19386,N_18748,N_18614);
nand U19387 (N_19387,N_18883,N_18197);
nand U19388 (N_19388,N_18511,N_18141);
xor U19389 (N_19389,N_18069,N_18529);
xnor U19390 (N_19390,N_18483,N_18049);
nor U19391 (N_19391,N_18869,N_18927);
nor U19392 (N_19392,N_18942,N_18390);
and U19393 (N_19393,N_18211,N_18591);
nand U19394 (N_19394,N_18982,N_18994);
xnor U19395 (N_19395,N_18427,N_18826);
xnor U19396 (N_19396,N_18618,N_18456);
and U19397 (N_19397,N_18176,N_18154);
nand U19398 (N_19398,N_18320,N_18688);
xor U19399 (N_19399,N_18484,N_18352);
nand U19400 (N_19400,N_18115,N_18288);
or U19401 (N_19401,N_18619,N_18368);
or U19402 (N_19402,N_18378,N_18093);
and U19403 (N_19403,N_18017,N_18995);
and U19404 (N_19404,N_18297,N_18503);
nor U19405 (N_19405,N_18194,N_18002);
or U19406 (N_19406,N_18042,N_18755);
or U19407 (N_19407,N_18402,N_18903);
xor U19408 (N_19408,N_18172,N_18400);
and U19409 (N_19409,N_18285,N_18015);
nand U19410 (N_19410,N_18239,N_18670);
xnor U19411 (N_19411,N_18035,N_18122);
nor U19412 (N_19412,N_18425,N_18558);
nand U19413 (N_19413,N_18050,N_18247);
or U19414 (N_19414,N_18433,N_18896);
xor U19415 (N_19415,N_18055,N_18557);
nand U19416 (N_19416,N_18226,N_18334);
nand U19417 (N_19417,N_18605,N_18373);
xor U19418 (N_19418,N_18344,N_18022);
xnor U19419 (N_19419,N_18201,N_18631);
nor U19420 (N_19420,N_18040,N_18203);
and U19421 (N_19421,N_18257,N_18623);
and U19422 (N_19422,N_18186,N_18629);
nand U19423 (N_19423,N_18626,N_18891);
nor U19424 (N_19424,N_18177,N_18292);
nand U19425 (N_19425,N_18399,N_18489);
nand U19426 (N_19426,N_18953,N_18068);
or U19427 (N_19427,N_18341,N_18753);
xor U19428 (N_19428,N_18862,N_18638);
and U19429 (N_19429,N_18787,N_18438);
or U19430 (N_19430,N_18403,N_18517);
or U19431 (N_19431,N_18452,N_18615);
xor U19432 (N_19432,N_18842,N_18271);
nor U19433 (N_19433,N_18362,N_18160);
and U19434 (N_19434,N_18353,N_18345);
or U19435 (N_19435,N_18915,N_18114);
nand U19436 (N_19436,N_18964,N_18075);
or U19437 (N_19437,N_18686,N_18662);
nor U19438 (N_19438,N_18773,N_18363);
or U19439 (N_19439,N_18683,N_18158);
xor U19440 (N_19440,N_18290,N_18356);
or U19441 (N_19441,N_18005,N_18318);
xnor U19442 (N_19442,N_18659,N_18794);
nor U19443 (N_19443,N_18877,N_18094);
nor U19444 (N_19444,N_18562,N_18471);
nor U19445 (N_19445,N_18981,N_18347);
nand U19446 (N_19446,N_18468,N_18228);
nand U19447 (N_19447,N_18382,N_18258);
nor U19448 (N_19448,N_18548,N_18237);
nand U19449 (N_19449,N_18936,N_18959);
or U19450 (N_19450,N_18111,N_18090);
and U19451 (N_19451,N_18809,N_18409);
and U19452 (N_19452,N_18635,N_18577);
nor U19453 (N_19453,N_18153,N_18365);
or U19454 (N_19454,N_18690,N_18871);
nand U19455 (N_19455,N_18076,N_18745);
xnor U19456 (N_19456,N_18553,N_18909);
xnor U19457 (N_19457,N_18151,N_18034);
nand U19458 (N_19458,N_18926,N_18567);
nand U19459 (N_19459,N_18127,N_18904);
xor U19460 (N_19460,N_18487,N_18868);
nand U19461 (N_19461,N_18808,N_18384);
or U19462 (N_19462,N_18410,N_18240);
nand U19463 (N_19463,N_18062,N_18307);
nor U19464 (N_19464,N_18587,N_18739);
nand U19465 (N_19465,N_18863,N_18884);
or U19466 (N_19466,N_18681,N_18336);
nor U19467 (N_19467,N_18306,N_18590);
nand U19468 (N_19468,N_18918,N_18889);
xnor U19469 (N_19469,N_18774,N_18424);
nor U19470 (N_19470,N_18515,N_18899);
and U19471 (N_19471,N_18103,N_18070);
and U19472 (N_19472,N_18539,N_18914);
and U19473 (N_19473,N_18244,N_18708);
or U19474 (N_19474,N_18806,N_18044);
or U19475 (N_19475,N_18551,N_18206);
xor U19476 (N_19476,N_18839,N_18369);
nand U19477 (N_19477,N_18543,N_18451);
nor U19478 (N_19478,N_18476,N_18125);
nand U19479 (N_19479,N_18771,N_18971);
or U19480 (N_19480,N_18458,N_18190);
or U19481 (N_19481,N_18325,N_18416);
or U19482 (N_19482,N_18006,N_18532);
or U19483 (N_19483,N_18841,N_18780);
nor U19484 (N_19484,N_18310,N_18500);
nor U19485 (N_19485,N_18593,N_18309);
xnor U19486 (N_19486,N_18929,N_18428);
and U19487 (N_19487,N_18814,N_18514);
xor U19488 (N_19488,N_18498,N_18460);
or U19489 (N_19489,N_18645,N_18137);
xor U19490 (N_19490,N_18934,N_18777);
nand U19491 (N_19491,N_18624,N_18775);
nor U19492 (N_19492,N_18849,N_18464);
nand U19493 (N_19493,N_18910,N_18278);
nand U19494 (N_19494,N_18268,N_18882);
nor U19495 (N_19495,N_18008,N_18113);
nand U19496 (N_19496,N_18963,N_18162);
nand U19497 (N_19497,N_18765,N_18875);
and U19498 (N_19498,N_18419,N_18463);
nand U19499 (N_19499,N_18603,N_18712);
and U19500 (N_19500,N_18348,N_18557);
nand U19501 (N_19501,N_18675,N_18756);
and U19502 (N_19502,N_18954,N_18981);
nor U19503 (N_19503,N_18262,N_18535);
and U19504 (N_19504,N_18846,N_18499);
and U19505 (N_19505,N_18196,N_18101);
and U19506 (N_19506,N_18111,N_18984);
nand U19507 (N_19507,N_18442,N_18387);
or U19508 (N_19508,N_18731,N_18846);
nand U19509 (N_19509,N_18640,N_18443);
and U19510 (N_19510,N_18060,N_18286);
nand U19511 (N_19511,N_18706,N_18857);
nand U19512 (N_19512,N_18712,N_18410);
nor U19513 (N_19513,N_18102,N_18146);
and U19514 (N_19514,N_18803,N_18737);
nor U19515 (N_19515,N_18647,N_18547);
xnor U19516 (N_19516,N_18406,N_18355);
and U19517 (N_19517,N_18199,N_18414);
or U19518 (N_19518,N_18659,N_18535);
xnor U19519 (N_19519,N_18922,N_18009);
nand U19520 (N_19520,N_18962,N_18991);
nand U19521 (N_19521,N_18276,N_18568);
xor U19522 (N_19522,N_18934,N_18852);
xor U19523 (N_19523,N_18713,N_18380);
nand U19524 (N_19524,N_18604,N_18676);
nand U19525 (N_19525,N_18526,N_18079);
nor U19526 (N_19526,N_18270,N_18102);
nand U19527 (N_19527,N_18959,N_18935);
nand U19528 (N_19528,N_18680,N_18723);
nor U19529 (N_19529,N_18194,N_18609);
nand U19530 (N_19530,N_18271,N_18941);
or U19531 (N_19531,N_18978,N_18730);
xor U19532 (N_19532,N_18297,N_18021);
nor U19533 (N_19533,N_18319,N_18772);
nand U19534 (N_19534,N_18799,N_18925);
xor U19535 (N_19535,N_18835,N_18144);
nand U19536 (N_19536,N_18775,N_18879);
and U19537 (N_19537,N_18402,N_18428);
nor U19538 (N_19538,N_18365,N_18807);
or U19539 (N_19539,N_18162,N_18102);
nand U19540 (N_19540,N_18004,N_18670);
xor U19541 (N_19541,N_18635,N_18542);
or U19542 (N_19542,N_18519,N_18937);
or U19543 (N_19543,N_18511,N_18187);
nand U19544 (N_19544,N_18068,N_18771);
nand U19545 (N_19545,N_18848,N_18673);
nor U19546 (N_19546,N_18945,N_18496);
nor U19547 (N_19547,N_18570,N_18026);
or U19548 (N_19548,N_18764,N_18662);
nand U19549 (N_19549,N_18376,N_18184);
nor U19550 (N_19550,N_18151,N_18941);
and U19551 (N_19551,N_18593,N_18338);
xor U19552 (N_19552,N_18576,N_18314);
nand U19553 (N_19553,N_18772,N_18387);
xnor U19554 (N_19554,N_18851,N_18969);
or U19555 (N_19555,N_18204,N_18856);
or U19556 (N_19556,N_18037,N_18552);
or U19557 (N_19557,N_18483,N_18081);
nor U19558 (N_19558,N_18470,N_18188);
nor U19559 (N_19559,N_18707,N_18169);
xnor U19560 (N_19560,N_18586,N_18961);
nor U19561 (N_19561,N_18262,N_18301);
nand U19562 (N_19562,N_18769,N_18041);
nand U19563 (N_19563,N_18233,N_18689);
and U19564 (N_19564,N_18404,N_18590);
or U19565 (N_19565,N_18907,N_18023);
nor U19566 (N_19566,N_18746,N_18563);
and U19567 (N_19567,N_18158,N_18014);
nor U19568 (N_19568,N_18224,N_18333);
xnor U19569 (N_19569,N_18073,N_18460);
xor U19570 (N_19570,N_18738,N_18989);
nor U19571 (N_19571,N_18060,N_18764);
or U19572 (N_19572,N_18025,N_18849);
and U19573 (N_19573,N_18773,N_18997);
and U19574 (N_19574,N_18612,N_18774);
and U19575 (N_19575,N_18094,N_18827);
and U19576 (N_19576,N_18061,N_18177);
nand U19577 (N_19577,N_18320,N_18863);
or U19578 (N_19578,N_18603,N_18457);
nand U19579 (N_19579,N_18239,N_18827);
xnor U19580 (N_19580,N_18083,N_18108);
nand U19581 (N_19581,N_18419,N_18511);
or U19582 (N_19582,N_18012,N_18945);
nand U19583 (N_19583,N_18882,N_18078);
nand U19584 (N_19584,N_18698,N_18497);
or U19585 (N_19585,N_18123,N_18361);
nand U19586 (N_19586,N_18724,N_18081);
nand U19587 (N_19587,N_18615,N_18501);
and U19588 (N_19588,N_18692,N_18955);
nor U19589 (N_19589,N_18661,N_18391);
nor U19590 (N_19590,N_18129,N_18017);
and U19591 (N_19591,N_18916,N_18341);
nor U19592 (N_19592,N_18688,N_18501);
nand U19593 (N_19593,N_18328,N_18188);
or U19594 (N_19594,N_18279,N_18851);
nand U19595 (N_19595,N_18532,N_18690);
or U19596 (N_19596,N_18426,N_18027);
and U19597 (N_19597,N_18320,N_18831);
and U19598 (N_19598,N_18487,N_18145);
nand U19599 (N_19599,N_18954,N_18627);
nand U19600 (N_19600,N_18225,N_18578);
nand U19601 (N_19601,N_18706,N_18524);
nand U19602 (N_19602,N_18220,N_18071);
xor U19603 (N_19603,N_18222,N_18121);
nor U19604 (N_19604,N_18801,N_18688);
nor U19605 (N_19605,N_18601,N_18265);
xnor U19606 (N_19606,N_18496,N_18806);
nand U19607 (N_19607,N_18934,N_18668);
or U19608 (N_19608,N_18563,N_18858);
xnor U19609 (N_19609,N_18232,N_18645);
and U19610 (N_19610,N_18302,N_18758);
nor U19611 (N_19611,N_18588,N_18275);
nand U19612 (N_19612,N_18095,N_18160);
nor U19613 (N_19613,N_18128,N_18340);
and U19614 (N_19614,N_18146,N_18007);
nor U19615 (N_19615,N_18257,N_18325);
nand U19616 (N_19616,N_18677,N_18455);
nand U19617 (N_19617,N_18836,N_18839);
and U19618 (N_19618,N_18826,N_18583);
nor U19619 (N_19619,N_18436,N_18549);
nand U19620 (N_19620,N_18445,N_18640);
nor U19621 (N_19621,N_18277,N_18947);
nor U19622 (N_19622,N_18150,N_18698);
nor U19623 (N_19623,N_18508,N_18482);
nor U19624 (N_19624,N_18386,N_18064);
nand U19625 (N_19625,N_18100,N_18459);
or U19626 (N_19626,N_18563,N_18943);
nand U19627 (N_19627,N_18608,N_18091);
and U19628 (N_19628,N_18411,N_18019);
nand U19629 (N_19629,N_18881,N_18786);
nor U19630 (N_19630,N_18600,N_18578);
or U19631 (N_19631,N_18450,N_18860);
or U19632 (N_19632,N_18298,N_18005);
nor U19633 (N_19633,N_18616,N_18768);
nor U19634 (N_19634,N_18709,N_18864);
and U19635 (N_19635,N_18608,N_18583);
xnor U19636 (N_19636,N_18605,N_18885);
and U19637 (N_19637,N_18966,N_18162);
and U19638 (N_19638,N_18824,N_18700);
nor U19639 (N_19639,N_18303,N_18330);
xor U19640 (N_19640,N_18960,N_18886);
nand U19641 (N_19641,N_18396,N_18039);
and U19642 (N_19642,N_18517,N_18979);
nor U19643 (N_19643,N_18894,N_18378);
or U19644 (N_19644,N_18007,N_18481);
xor U19645 (N_19645,N_18663,N_18819);
or U19646 (N_19646,N_18596,N_18638);
xor U19647 (N_19647,N_18554,N_18428);
or U19648 (N_19648,N_18612,N_18756);
or U19649 (N_19649,N_18929,N_18808);
nand U19650 (N_19650,N_18474,N_18499);
and U19651 (N_19651,N_18474,N_18537);
nand U19652 (N_19652,N_18752,N_18856);
nor U19653 (N_19653,N_18459,N_18354);
nor U19654 (N_19654,N_18863,N_18324);
and U19655 (N_19655,N_18511,N_18047);
and U19656 (N_19656,N_18984,N_18898);
nand U19657 (N_19657,N_18732,N_18954);
and U19658 (N_19658,N_18226,N_18266);
or U19659 (N_19659,N_18223,N_18304);
xnor U19660 (N_19660,N_18392,N_18255);
nand U19661 (N_19661,N_18179,N_18427);
nand U19662 (N_19662,N_18577,N_18585);
or U19663 (N_19663,N_18591,N_18413);
and U19664 (N_19664,N_18342,N_18578);
xnor U19665 (N_19665,N_18419,N_18922);
or U19666 (N_19666,N_18046,N_18980);
and U19667 (N_19667,N_18252,N_18182);
nor U19668 (N_19668,N_18196,N_18119);
or U19669 (N_19669,N_18128,N_18218);
nand U19670 (N_19670,N_18857,N_18397);
and U19671 (N_19671,N_18260,N_18891);
and U19672 (N_19672,N_18907,N_18982);
xnor U19673 (N_19673,N_18128,N_18653);
or U19674 (N_19674,N_18798,N_18780);
xnor U19675 (N_19675,N_18885,N_18282);
nand U19676 (N_19676,N_18819,N_18764);
or U19677 (N_19677,N_18106,N_18676);
and U19678 (N_19678,N_18578,N_18786);
nor U19679 (N_19679,N_18280,N_18333);
or U19680 (N_19680,N_18433,N_18609);
xnor U19681 (N_19681,N_18351,N_18478);
nor U19682 (N_19682,N_18679,N_18347);
or U19683 (N_19683,N_18405,N_18588);
nand U19684 (N_19684,N_18187,N_18620);
and U19685 (N_19685,N_18876,N_18631);
and U19686 (N_19686,N_18459,N_18994);
or U19687 (N_19687,N_18501,N_18012);
or U19688 (N_19688,N_18869,N_18947);
nor U19689 (N_19689,N_18460,N_18103);
xor U19690 (N_19690,N_18499,N_18658);
nor U19691 (N_19691,N_18872,N_18949);
xnor U19692 (N_19692,N_18526,N_18360);
nand U19693 (N_19693,N_18164,N_18055);
and U19694 (N_19694,N_18841,N_18914);
nor U19695 (N_19695,N_18388,N_18902);
and U19696 (N_19696,N_18244,N_18887);
nor U19697 (N_19697,N_18161,N_18538);
and U19698 (N_19698,N_18908,N_18994);
nand U19699 (N_19699,N_18524,N_18274);
nor U19700 (N_19700,N_18805,N_18153);
nor U19701 (N_19701,N_18510,N_18433);
and U19702 (N_19702,N_18204,N_18572);
nor U19703 (N_19703,N_18000,N_18164);
xnor U19704 (N_19704,N_18396,N_18876);
or U19705 (N_19705,N_18915,N_18909);
or U19706 (N_19706,N_18380,N_18147);
or U19707 (N_19707,N_18372,N_18065);
and U19708 (N_19708,N_18796,N_18087);
nand U19709 (N_19709,N_18188,N_18093);
or U19710 (N_19710,N_18965,N_18901);
nand U19711 (N_19711,N_18365,N_18244);
nor U19712 (N_19712,N_18555,N_18182);
nand U19713 (N_19713,N_18522,N_18386);
xnor U19714 (N_19714,N_18284,N_18202);
xor U19715 (N_19715,N_18256,N_18904);
and U19716 (N_19716,N_18549,N_18905);
nor U19717 (N_19717,N_18621,N_18232);
or U19718 (N_19718,N_18846,N_18177);
xor U19719 (N_19719,N_18191,N_18734);
nor U19720 (N_19720,N_18596,N_18236);
and U19721 (N_19721,N_18616,N_18751);
nor U19722 (N_19722,N_18350,N_18846);
xor U19723 (N_19723,N_18281,N_18997);
and U19724 (N_19724,N_18139,N_18898);
xor U19725 (N_19725,N_18364,N_18167);
xor U19726 (N_19726,N_18463,N_18795);
and U19727 (N_19727,N_18407,N_18047);
nand U19728 (N_19728,N_18485,N_18210);
nand U19729 (N_19729,N_18176,N_18461);
xor U19730 (N_19730,N_18258,N_18942);
or U19731 (N_19731,N_18842,N_18759);
nand U19732 (N_19732,N_18752,N_18595);
nand U19733 (N_19733,N_18541,N_18972);
nor U19734 (N_19734,N_18241,N_18069);
or U19735 (N_19735,N_18785,N_18858);
or U19736 (N_19736,N_18735,N_18617);
nor U19737 (N_19737,N_18751,N_18014);
nor U19738 (N_19738,N_18011,N_18016);
or U19739 (N_19739,N_18454,N_18431);
nand U19740 (N_19740,N_18456,N_18428);
nor U19741 (N_19741,N_18897,N_18663);
nor U19742 (N_19742,N_18245,N_18163);
xnor U19743 (N_19743,N_18900,N_18716);
nor U19744 (N_19744,N_18787,N_18744);
nand U19745 (N_19745,N_18072,N_18834);
and U19746 (N_19746,N_18300,N_18227);
and U19747 (N_19747,N_18945,N_18943);
or U19748 (N_19748,N_18389,N_18826);
or U19749 (N_19749,N_18551,N_18461);
xnor U19750 (N_19750,N_18483,N_18959);
or U19751 (N_19751,N_18328,N_18292);
nand U19752 (N_19752,N_18179,N_18827);
nand U19753 (N_19753,N_18627,N_18691);
nand U19754 (N_19754,N_18057,N_18756);
and U19755 (N_19755,N_18642,N_18880);
nor U19756 (N_19756,N_18332,N_18438);
and U19757 (N_19757,N_18843,N_18130);
and U19758 (N_19758,N_18872,N_18847);
xor U19759 (N_19759,N_18147,N_18487);
nor U19760 (N_19760,N_18754,N_18254);
xnor U19761 (N_19761,N_18700,N_18698);
or U19762 (N_19762,N_18676,N_18838);
nand U19763 (N_19763,N_18190,N_18942);
xnor U19764 (N_19764,N_18980,N_18463);
and U19765 (N_19765,N_18739,N_18107);
xnor U19766 (N_19766,N_18067,N_18077);
nand U19767 (N_19767,N_18594,N_18210);
nor U19768 (N_19768,N_18713,N_18735);
nand U19769 (N_19769,N_18595,N_18069);
and U19770 (N_19770,N_18287,N_18187);
and U19771 (N_19771,N_18288,N_18883);
and U19772 (N_19772,N_18777,N_18583);
and U19773 (N_19773,N_18847,N_18153);
xnor U19774 (N_19774,N_18539,N_18015);
or U19775 (N_19775,N_18343,N_18651);
xnor U19776 (N_19776,N_18848,N_18918);
and U19777 (N_19777,N_18064,N_18246);
xnor U19778 (N_19778,N_18183,N_18538);
nor U19779 (N_19779,N_18595,N_18516);
nor U19780 (N_19780,N_18589,N_18861);
and U19781 (N_19781,N_18499,N_18203);
nand U19782 (N_19782,N_18531,N_18073);
xnor U19783 (N_19783,N_18697,N_18285);
or U19784 (N_19784,N_18842,N_18184);
and U19785 (N_19785,N_18577,N_18610);
nand U19786 (N_19786,N_18877,N_18403);
and U19787 (N_19787,N_18284,N_18634);
or U19788 (N_19788,N_18187,N_18637);
and U19789 (N_19789,N_18693,N_18528);
xor U19790 (N_19790,N_18294,N_18942);
nand U19791 (N_19791,N_18499,N_18131);
xnor U19792 (N_19792,N_18231,N_18550);
nand U19793 (N_19793,N_18222,N_18794);
xor U19794 (N_19794,N_18039,N_18787);
or U19795 (N_19795,N_18875,N_18248);
and U19796 (N_19796,N_18525,N_18653);
nor U19797 (N_19797,N_18986,N_18885);
nor U19798 (N_19798,N_18627,N_18629);
nor U19799 (N_19799,N_18521,N_18728);
nand U19800 (N_19800,N_18843,N_18517);
and U19801 (N_19801,N_18727,N_18285);
nand U19802 (N_19802,N_18963,N_18412);
xor U19803 (N_19803,N_18119,N_18657);
nand U19804 (N_19804,N_18317,N_18351);
nand U19805 (N_19805,N_18025,N_18522);
xor U19806 (N_19806,N_18236,N_18658);
xnor U19807 (N_19807,N_18936,N_18739);
or U19808 (N_19808,N_18705,N_18609);
or U19809 (N_19809,N_18564,N_18148);
and U19810 (N_19810,N_18709,N_18786);
nor U19811 (N_19811,N_18341,N_18093);
nand U19812 (N_19812,N_18092,N_18757);
nand U19813 (N_19813,N_18074,N_18579);
xnor U19814 (N_19814,N_18010,N_18746);
nor U19815 (N_19815,N_18504,N_18268);
nor U19816 (N_19816,N_18912,N_18990);
nand U19817 (N_19817,N_18657,N_18851);
and U19818 (N_19818,N_18500,N_18570);
and U19819 (N_19819,N_18335,N_18077);
xor U19820 (N_19820,N_18154,N_18874);
and U19821 (N_19821,N_18671,N_18649);
nand U19822 (N_19822,N_18048,N_18378);
nor U19823 (N_19823,N_18604,N_18040);
and U19824 (N_19824,N_18100,N_18107);
or U19825 (N_19825,N_18564,N_18926);
or U19826 (N_19826,N_18065,N_18413);
nand U19827 (N_19827,N_18355,N_18032);
and U19828 (N_19828,N_18249,N_18113);
or U19829 (N_19829,N_18756,N_18071);
nand U19830 (N_19830,N_18445,N_18926);
nor U19831 (N_19831,N_18548,N_18987);
or U19832 (N_19832,N_18819,N_18511);
and U19833 (N_19833,N_18993,N_18577);
xnor U19834 (N_19834,N_18724,N_18875);
and U19835 (N_19835,N_18004,N_18693);
xnor U19836 (N_19836,N_18460,N_18229);
or U19837 (N_19837,N_18849,N_18613);
xnor U19838 (N_19838,N_18115,N_18940);
and U19839 (N_19839,N_18129,N_18681);
nor U19840 (N_19840,N_18245,N_18643);
or U19841 (N_19841,N_18000,N_18146);
and U19842 (N_19842,N_18669,N_18095);
and U19843 (N_19843,N_18306,N_18495);
xor U19844 (N_19844,N_18079,N_18806);
nand U19845 (N_19845,N_18065,N_18981);
and U19846 (N_19846,N_18540,N_18010);
and U19847 (N_19847,N_18573,N_18560);
and U19848 (N_19848,N_18882,N_18234);
and U19849 (N_19849,N_18838,N_18717);
nor U19850 (N_19850,N_18467,N_18621);
and U19851 (N_19851,N_18020,N_18546);
nand U19852 (N_19852,N_18943,N_18240);
or U19853 (N_19853,N_18181,N_18484);
and U19854 (N_19854,N_18733,N_18065);
xor U19855 (N_19855,N_18609,N_18644);
nor U19856 (N_19856,N_18728,N_18154);
xor U19857 (N_19857,N_18208,N_18267);
nor U19858 (N_19858,N_18432,N_18152);
nor U19859 (N_19859,N_18001,N_18861);
nor U19860 (N_19860,N_18725,N_18929);
xor U19861 (N_19861,N_18695,N_18174);
nand U19862 (N_19862,N_18843,N_18487);
or U19863 (N_19863,N_18631,N_18634);
or U19864 (N_19864,N_18229,N_18049);
xor U19865 (N_19865,N_18297,N_18461);
nor U19866 (N_19866,N_18838,N_18965);
nor U19867 (N_19867,N_18925,N_18334);
and U19868 (N_19868,N_18810,N_18424);
xnor U19869 (N_19869,N_18067,N_18525);
or U19870 (N_19870,N_18844,N_18577);
xnor U19871 (N_19871,N_18689,N_18122);
or U19872 (N_19872,N_18442,N_18500);
and U19873 (N_19873,N_18552,N_18893);
or U19874 (N_19874,N_18942,N_18768);
nand U19875 (N_19875,N_18527,N_18238);
and U19876 (N_19876,N_18834,N_18541);
nand U19877 (N_19877,N_18020,N_18705);
xnor U19878 (N_19878,N_18551,N_18757);
or U19879 (N_19879,N_18382,N_18081);
or U19880 (N_19880,N_18420,N_18449);
or U19881 (N_19881,N_18239,N_18114);
nor U19882 (N_19882,N_18234,N_18006);
or U19883 (N_19883,N_18893,N_18096);
or U19884 (N_19884,N_18006,N_18640);
or U19885 (N_19885,N_18264,N_18888);
or U19886 (N_19886,N_18597,N_18306);
xnor U19887 (N_19887,N_18526,N_18129);
and U19888 (N_19888,N_18159,N_18091);
or U19889 (N_19889,N_18943,N_18534);
nand U19890 (N_19890,N_18257,N_18377);
or U19891 (N_19891,N_18793,N_18599);
and U19892 (N_19892,N_18511,N_18423);
and U19893 (N_19893,N_18398,N_18959);
and U19894 (N_19894,N_18305,N_18158);
and U19895 (N_19895,N_18134,N_18987);
nor U19896 (N_19896,N_18724,N_18487);
or U19897 (N_19897,N_18270,N_18297);
xnor U19898 (N_19898,N_18580,N_18096);
or U19899 (N_19899,N_18571,N_18501);
nand U19900 (N_19900,N_18565,N_18314);
xor U19901 (N_19901,N_18652,N_18882);
or U19902 (N_19902,N_18889,N_18728);
or U19903 (N_19903,N_18355,N_18770);
and U19904 (N_19904,N_18108,N_18227);
xnor U19905 (N_19905,N_18897,N_18291);
nor U19906 (N_19906,N_18015,N_18002);
nor U19907 (N_19907,N_18047,N_18288);
xnor U19908 (N_19908,N_18751,N_18967);
nand U19909 (N_19909,N_18416,N_18374);
nor U19910 (N_19910,N_18754,N_18502);
xor U19911 (N_19911,N_18286,N_18567);
or U19912 (N_19912,N_18208,N_18381);
and U19913 (N_19913,N_18783,N_18829);
and U19914 (N_19914,N_18637,N_18267);
or U19915 (N_19915,N_18445,N_18789);
xnor U19916 (N_19916,N_18625,N_18258);
and U19917 (N_19917,N_18956,N_18686);
or U19918 (N_19918,N_18798,N_18568);
nor U19919 (N_19919,N_18314,N_18092);
and U19920 (N_19920,N_18769,N_18224);
xor U19921 (N_19921,N_18394,N_18416);
and U19922 (N_19922,N_18869,N_18408);
xor U19923 (N_19923,N_18597,N_18257);
xnor U19924 (N_19924,N_18700,N_18831);
or U19925 (N_19925,N_18908,N_18492);
and U19926 (N_19926,N_18643,N_18065);
or U19927 (N_19927,N_18856,N_18578);
nor U19928 (N_19928,N_18581,N_18216);
nor U19929 (N_19929,N_18924,N_18152);
nand U19930 (N_19930,N_18170,N_18077);
xor U19931 (N_19931,N_18297,N_18974);
or U19932 (N_19932,N_18665,N_18893);
or U19933 (N_19933,N_18702,N_18826);
and U19934 (N_19934,N_18581,N_18503);
nand U19935 (N_19935,N_18203,N_18445);
or U19936 (N_19936,N_18822,N_18158);
xor U19937 (N_19937,N_18608,N_18461);
and U19938 (N_19938,N_18122,N_18702);
xor U19939 (N_19939,N_18336,N_18137);
or U19940 (N_19940,N_18069,N_18308);
nor U19941 (N_19941,N_18701,N_18850);
nand U19942 (N_19942,N_18572,N_18590);
and U19943 (N_19943,N_18935,N_18990);
or U19944 (N_19944,N_18000,N_18721);
nor U19945 (N_19945,N_18801,N_18967);
nand U19946 (N_19946,N_18862,N_18099);
xor U19947 (N_19947,N_18634,N_18667);
nand U19948 (N_19948,N_18406,N_18557);
xnor U19949 (N_19949,N_18200,N_18432);
nor U19950 (N_19950,N_18574,N_18778);
or U19951 (N_19951,N_18897,N_18011);
and U19952 (N_19952,N_18329,N_18623);
xnor U19953 (N_19953,N_18525,N_18284);
xor U19954 (N_19954,N_18842,N_18523);
nor U19955 (N_19955,N_18542,N_18888);
or U19956 (N_19956,N_18847,N_18713);
or U19957 (N_19957,N_18244,N_18435);
xnor U19958 (N_19958,N_18680,N_18576);
nor U19959 (N_19959,N_18691,N_18041);
or U19960 (N_19960,N_18229,N_18784);
nand U19961 (N_19961,N_18312,N_18287);
or U19962 (N_19962,N_18189,N_18041);
nor U19963 (N_19963,N_18661,N_18878);
or U19964 (N_19964,N_18961,N_18397);
and U19965 (N_19965,N_18605,N_18830);
nor U19966 (N_19966,N_18658,N_18947);
nand U19967 (N_19967,N_18527,N_18237);
nor U19968 (N_19968,N_18616,N_18662);
or U19969 (N_19969,N_18588,N_18655);
or U19970 (N_19970,N_18919,N_18257);
nor U19971 (N_19971,N_18223,N_18774);
nand U19972 (N_19972,N_18045,N_18855);
and U19973 (N_19973,N_18062,N_18249);
or U19974 (N_19974,N_18415,N_18730);
nor U19975 (N_19975,N_18930,N_18802);
nor U19976 (N_19976,N_18601,N_18677);
nand U19977 (N_19977,N_18119,N_18942);
xor U19978 (N_19978,N_18137,N_18768);
and U19979 (N_19979,N_18154,N_18138);
nand U19980 (N_19980,N_18943,N_18758);
nor U19981 (N_19981,N_18844,N_18493);
xnor U19982 (N_19982,N_18940,N_18366);
and U19983 (N_19983,N_18565,N_18271);
and U19984 (N_19984,N_18858,N_18398);
xor U19985 (N_19985,N_18449,N_18940);
and U19986 (N_19986,N_18121,N_18580);
nand U19987 (N_19987,N_18941,N_18842);
xnor U19988 (N_19988,N_18298,N_18514);
or U19989 (N_19989,N_18396,N_18133);
or U19990 (N_19990,N_18593,N_18355);
or U19991 (N_19991,N_18668,N_18927);
nand U19992 (N_19992,N_18602,N_18366);
or U19993 (N_19993,N_18899,N_18656);
nand U19994 (N_19994,N_18486,N_18759);
nor U19995 (N_19995,N_18347,N_18898);
and U19996 (N_19996,N_18809,N_18696);
and U19997 (N_19997,N_18655,N_18553);
nand U19998 (N_19998,N_18028,N_18712);
or U19999 (N_19999,N_18904,N_18475);
or UO_0 (O_0,N_19312,N_19757);
nor UO_1 (O_1,N_19730,N_19678);
xnor UO_2 (O_2,N_19548,N_19028);
xnor UO_3 (O_3,N_19444,N_19474);
or UO_4 (O_4,N_19295,N_19531);
xor UO_5 (O_5,N_19577,N_19668);
and UO_6 (O_6,N_19773,N_19641);
or UO_7 (O_7,N_19570,N_19006);
or UO_8 (O_8,N_19137,N_19638);
or UO_9 (O_9,N_19852,N_19590);
xnor UO_10 (O_10,N_19250,N_19311);
or UO_11 (O_11,N_19973,N_19310);
or UO_12 (O_12,N_19176,N_19236);
xor UO_13 (O_13,N_19080,N_19864);
nand UO_14 (O_14,N_19631,N_19658);
nand UO_15 (O_15,N_19924,N_19732);
nor UO_16 (O_16,N_19575,N_19983);
and UO_17 (O_17,N_19323,N_19663);
or UO_18 (O_18,N_19190,N_19179);
nor UO_19 (O_19,N_19533,N_19246);
xnor UO_20 (O_20,N_19680,N_19736);
nand UO_21 (O_21,N_19065,N_19442);
xnor UO_22 (O_22,N_19596,N_19626);
and UO_23 (O_23,N_19709,N_19696);
and UO_24 (O_24,N_19768,N_19814);
or UO_25 (O_25,N_19978,N_19016);
and UO_26 (O_26,N_19748,N_19922);
xnor UO_27 (O_27,N_19933,N_19127);
xor UO_28 (O_28,N_19778,N_19745);
nand UO_29 (O_29,N_19298,N_19119);
or UO_30 (O_30,N_19530,N_19159);
nor UO_31 (O_31,N_19327,N_19164);
or UO_32 (O_32,N_19997,N_19856);
or UO_33 (O_33,N_19683,N_19829);
and UO_34 (O_34,N_19358,N_19499);
and UO_35 (O_35,N_19979,N_19661);
nor UO_36 (O_36,N_19846,N_19282);
nor UO_37 (O_37,N_19850,N_19288);
or UO_38 (O_38,N_19194,N_19656);
and UO_39 (O_39,N_19320,N_19884);
and UO_40 (O_40,N_19669,N_19302);
and UO_41 (O_41,N_19636,N_19868);
or UO_42 (O_42,N_19992,N_19999);
or UO_43 (O_43,N_19986,N_19168);
nor UO_44 (O_44,N_19875,N_19453);
xor UO_45 (O_45,N_19277,N_19685);
nand UO_46 (O_46,N_19247,N_19618);
xor UO_47 (O_47,N_19508,N_19809);
or UO_48 (O_48,N_19838,N_19177);
nor UO_49 (O_49,N_19617,N_19439);
or UO_50 (O_50,N_19431,N_19480);
or UO_51 (O_51,N_19975,N_19869);
nand UO_52 (O_52,N_19064,N_19728);
xor UO_53 (O_53,N_19202,N_19811);
nor UO_54 (O_54,N_19184,N_19557);
or UO_55 (O_55,N_19085,N_19567);
xor UO_56 (O_56,N_19723,N_19029);
xor UO_57 (O_57,N_19402,N_19645);
or UO_58 (O_58,N_19984,N_19412);
nand UO_59 (O_59,N_19138,N_19981);
or UO_60 (O_60,N_19055,N_19753);
or UO_61 (O_61,N_19970,N_19013);
nor UO_62 (O_62,N_19482,N_19813);
or UO_63 (O_63,N_19147,N_19498);
and UO_64 (O_64,N_19403,N_19964);
nand UO_65 (O_65,N_19091,N_19241);
nand UO_66 (O_66,N_19428,N_19271);
nor UO_67 (O_67,N_19654,N_19974);
xor UO_68 (O_68,N_19234,N_19321);
xor UO_69 (O_69,N_19695,N_19054);
and UO_70 (O_70,N_19361,N_19270);
or UO_71 (O_71,N_19795,N_19810);
and UO_72 (O_72,N_19681,N_19275);
and UO_73 (O_73,N_19162,N_19643);
nor UO_74 (O_74,N_19971,N_19634);
nand UO_75 (O_75,N_19892,N_19279);
nand UO_76 (O_76,N_19665,N_19576);
nor UO_77 (O_77,N_19538,N_19142);
nand UO_78 (O_78,N_19819,N_19655);
or UO_79 (O_79,N_19861,N_19827);
and UO_80 (O_80,N_19969,N_19233);
nor UO_81 (O_81,N_19607,N_19105);
nor UO_82 (O_82,N_19715,N_19502);
and UO_83 (O_83,N_19163,N_19269);
and UO_84 (O_84,N_19472,N_19896);
and UO_85 (O_85,N_19662,N_19051);
nand UO_86 (O_86,N_19747,N_19490);
xnor UO_87 (O_87,N_19647,N_19157);
nor UO_88 (O_88,N_19961,N_19552);
xnor UO_89 (O_89,N_19289,N_19468);
or UO_90 (O_90,N_19450,N_19957);
or UO_91 (O_91,N_19416,N_19521);
xnor UO_92 (O_92,N_19409,N_19877);
nor UO_93 (O_93,N_19200,N_19996);
or UO_94 (O_94,N_19382,N_19007);
or UO_95 (O_95,N_19990,N_19441);
xnor UO_96 (O_96,N_19927,N_19017);
nor UO_97 (O_97,N_19187,N_19429);
nand UO_98 (O_98,N_19229,N_19938);
and UO_99 (O_99,N_19433,N_19751);
xnor UO_100 (O_100,N_19908,N_19684);
xnor UO_101 (O_101,N_19338,N_19847);
nand UO_102 (O_102,N_19265,N_19760);
xnor UO_103 (O_103,N_19686,N_19580);
nor UO_104 (O_104,N_19722,N_19405);
nand UO_105 (O_105,N_19632,N_19204);
xor UO_106 (O_106,N_19329,N_19100);
and UO_107 (O_107,N_19769,N_19153);
and UO_108 (O_108,N_19335,N_19534);
or UO_109 (O_109,N_19789,N_19627);
nor UO_110 (O_110,N_19285,N_19144);
nor UO_111 (O_111,N_19072,N_19779);
and UO_112 (O_112,N_19860,N_19161);
and UO_113 (O_113,N_19261,N_19802);
or UO_114 (O_114,N_19232,N_19040);
nand UO_115 (O_115,N_19340,N_19420);
and UO_116 (O_116,N_19758,N_19737);
nor UO_117 (O_117,N_19267,N_19437);
nor UO_118 (O_118,N_19305,N_19995);
xnor UO_119 (O_119,N_19713,N_19793);
nor UO_120 (O_120,N_19422,N_19724);
and UO_121 (O_121,N_19824,N_19560);
and UO_122 (O_122,N_19023,N_19301);
and UO_123 (O_123,N_19395,N_19092);
nand UO_124 (O_124,N_19166,N_19484);
nand UO_125 (O_125,N_19749,N_19317);
nor UO_126 (O_126,N_19185,N_19449);
xnor UO_127 (O_127,N_19503,N_19063);
and UO_128 (O_128,N_19718,N_19421);
xnor UO_129 (O_129,N_19389,N_19701);
nand UO_130 (O_130,N_19839,N_19799);
nand UO_131 (O_131,N_19803,N_19589);
or UO_132 (O_132,N_19507,N_19294);
and UO_133 (O_133,N_19352,N_19364);
and UO_134 (O_134,N_19336,N_19096);
and UO_135 (O_135,N_19622,N_19264);
and UO_136 (O_136,N_19033,N_19511);
nand UO_137 (O_137,N_19783,N_19396);
xor UO_138 (O_138,N_19553,N_19401);
or UO_139 (O_139,N_19906,N_19619);
nor UO_140 (O_140,N_19256,N_19370);
xor UO_141 (O_141,N_19942,N_19390);
nand UO_142 (O_142,N_19316,N_19192);
and UO_143 (O_143,N_19967,N_19744);
and UO_144 (O_144,N_19280,N_19326);
nand UO_145 (O_145,N_19674,N_19909);
and UO_146 (O_146,N_19989,N_19644);
xnor UO_147 (O_147,N_19058,N_19516);
or UO_148 (O_148,N_19452,N_19203);
nor UO_149 (O_149,N_19591,N_19427);
or UO_150 (O_150,N_19487,N_19688);
nand UO_151 (O_151,N_19462,N_19633);
xnor UO_152 (O_152,N_19785,N_19331);
or UO_153 (O_153,N_19107,N_19729);
or UO_154 (O_154,N_19876,N_19239);
xor UO_155 (O_155,N_19344,N_19608);
or UO_156 (O_156,N_19337,N_19068);
or UO_157 (O_157,N_19037,N_19515);
and UO_158 (O_158,N_19777,N_19010);
nand UO_159 (O_159,N_19259,N_19598);
xor UO_160 (O_160,N_19451,N_19693);
xor UO_161 (O_161,N_19886,N_19287);
and UO_162 (O_162,N_19980,N_19394);
or UO_163 (O_163,N_19169,N_19549);
and UO_164 (O_164,N_19299,N_19489);
or UO_165 (O_165,N_19196,N_19283);
and UO_166 (O_166,N_19483,N_19035);
nand UO_167 (O_167,N_19798,N_19488);
nor UO_168 (O_168,N_19960,N_19500);
nand UO_169 (O_169,N_19457,N_19497);
and UO_170 (O_170,N_19066,N_19062);
xor UO_171 (O_171,N_19670,N_19787);
or UO_172 (O_172,N_19893,N_19284);
xor UO_173 (O_173,N_19290,N_19935);
or UO_174 (O_174,N_19805,N_19952);
xor UO_175 (O_175,N_19081,N_19426);
nor UO_176 (O_176,N_19214,N_19806);
nand UO_177 (O_177,N_19341,N_19308);
nor UO_178 (O_178,N_19380,N_19966);
or UO_179 (O_179,N_19826,N_19849);
nor UO_180 (O_180,N_19940,N_19123);
and UO_181 (O_181,N_19346,N_19817);
and UO_182 (O_182,N_19815,N_19476);
nor UO_183 (O_183,N_19821,N_19599);
nand UO_184 (O_184,N_19293,N_19628);
and UO_185 (O_185,N_19660,N_19883);
and UO_186 (O_186,N_19145,N_19198);
nand UO_187 (O_187,N_19378,N_19559);
nor UO_188 (O_188,N_19953,N_19330);
xnor UO_189 (O_189,N_19460,N_19188);
and UO_190 (O_190,N_19690,N_19889);
and UO_191 (O_191,N_19148,N_19513);
nand UO_192 (O_192,N_19637,N_19720);
or UO_193 (O_193,N_19251,N_19478);
nor UO_194 (O_194,N_19900,N_19359);
nand UO_195 (O_195,N_19630,N_19215);
or UO_196 (O_196,N_19220,N_19274);
and UO_197 (O_197,N_19003,N_19888);
nor UO_198 (O_198,N_19083,N_19620);
nor UO_199 (O_199,N_19116,N_19770);
nand UO_200 (O_200,N_19930,N_19398);
or UO_201 (O_201,N_19131,N_19871);
or UO_202 (O_202,N_19180,N_19755);
and UO_203 (O_203,N_19175,N_19550);
nand UO_204 (O_204,N_19465,N_19774);
nand UO_205 (O_205,N_19463,N_19252);
xnor UO_206 (O_206,N_19303,N_19543);
and UO_207 (O_207,N_19985,N_19300);
or UO_208 (O_208,N_19088,N_19762);
nand UO_209 (O_209,N_19791,N_19114);
nor UO_210 (O_210,N_19929,N_19958);
or UO_211 (O_211,N_19928,N_19193);
and UO_212 (O_212,N_19977,N_19613);
xnor UO_213 (O_213,N_19902,N_19309);
and UO_214 (O_214,N_19879,N_19207);
and UO_215 (O_215,N_19031,N_19495);
and UO_216 (O_216,N_19609,N_19135);
or UO_217 (O_217,N_19171,N_19725);
xor UO_218 (O_218,N_19566,N_19705);
nand UO_219 (O_219,N_19424,N_19432);
nand UO_220 (O_220,N_19243,N_19049);
xnor UO_221 (O_221,N_19694,N_19227);
nand UO_222 (O_222,N_19112,N_19077);
and UO_223 (O_223,N_19213,N_19629);
nor UO_224 (O_224,N_19959,N_19245);
xor UO_225 (O_225,N_19110,N_19368);
and UO_226 (O_226,N_19717,N_19923);
or UO_227 (O_227,N_19039,N_19520);
nor UO_228 (O_228,N_19208,N_19564);
nand UO_229 (O_229,N_19651,N_19692);
or UO_230 (O_230,N_19226,N_19012);
and UO_231 (O_231,N_19640,N_19014);
xor UO_232 (O_232,N_19915,N_19529);
xnor UO_233 (O_233,N_19845,N_19143);
xnor UO_234 (O_234,N_19676,N_19128);
and UO_235 (O_235,N_19324,N_19504);
nand UO_236 (O_236,N_19721,N_19800);
and UO_237 (O_237,N_19238,N_19649);
and UO_238 (O_238,N_19882,N_19071);
nor UO_239 (O_239,N_19963,N_19291);
xnor UO_240 (O_240,N_19895,N_19764);
nor UO_241 (O_241,N_19372,N_19501);
nand UO_242 (O_242,N_19825,N_19939);
nor UO_243 (O_243,N_19859,N_19904);
nand UO_244 (O_244,N_19339,N_19257);
nor UO_245 (O_245,N_19833,N_19170);
nand UO_246 (O_246,N_19060,N_19743);
nor UO_247 (O_247,N_19367,N_19230);
and UO_248 (O_248,N_19258,N_19746);
and UO_249 (O_249,N_19122,N_19413);
nand UO_250 (O_250,N_19820,N_19182);
nand UO_251 (O_251,N_19946,N_19244);
or UO_252 (O_252,N_19089,N_19752);
nand UO_253 (O_253,N_19255,N_19905);
nand UO_254 (O_254,N_19260,N_19881);
and UO_255 (O_255,N_19894,N_19443);
nor UO_256 (O_256,N_19509,N_19286);
nor UO_257 (O_257,N_19387,N_19150);
nor UO_258 (O_258,N_19322,N_19816);
xnor UO_259 (O_259,N_19742,N_19253);
and UO_260 (O_260,N_19120,N_19121);
xnor UO_261 (O_261,N_19854,N_19796);
xor UO_262 (O_262,N_19801,N_19750);
or UO_263 (O_263,N_19041,N_19178);
or UO_264 (O_264,N_19702,N_19972);
or UO_265 (O_265,N_19537,N_19790);
nor UO_266 (O_266,N_19624,N_19672);
nand UO_267 (O_267,N_19183,N_19991);
nand UO_268 (O_268,N_19165,N_19197);
or UO_269 (O_269,N_19414,N_19926);
xor UO_270 (O_270,N_19887,N_19399);
and UO_271 (O_271,N_19018,N_19831);
nor UO_272 (O_272,N_19406,N_19767);
xor UO_273 (O_273,N_19224,N_19872);
or UO_274 (O_274,N_19955,N_19001);
and UO_275 (O_275,N_19333,N_19074);
or UO_276 (O_276,N_19739,N_19130);
xor UO_277 (O_277,N_19385,N_19221);
xnor UO_278 (O_278,N_19351,N_19154);
nor UO_279 (O_279,N_19075,N_19571);
and UO_280 (O_280,N_19700,N_19673);
nand UO_281 (O_281,N_19697,N_19588);
and UO_282 (O_282,N_19106,N_19440);
and UO_283 (O_283,N_19532,N_19965);
xor UO_284 (O_284,N_19699,N_19400);
or UO_285 (O_285,N_19536,N_19857);
xor UO_286 (O_286,N_19334,N_19297);
nor UO_287 (O_287,N_19493,N_19461);
and UO_288 (O_288,N_19343,N_19191);
nor UO_289 (O_289,N_19830,N_19237);
or UO_290 (O_290,N_19993,N_19047);
nand UO_291 (O_291,N_19407,N_19086);
and UO_292 (O_292,N_19834,N_19002);
nand UO_293 (O_293,N_19158,N_19698);
or UO_294 (O_294,N_19318,N_19099);
nor UO_295 (O_295,N_19522,N_19761);
or UO_296 (O_296,N_19563,N_19019);
and UO_297 (O_297,N_19574,N_19411);
xnor UO_298 (O_298,N_19916,N_19603);
nand UO_299 (O_299,N_19004,N_19473);
nand UO_300 (O_300,N_19865,N_19219);
or UO_301 (O_301,N_19561,N_19082);
nor UO_302 (O_302,N_19842,N_19210);
xor UO_303 (O_303,N_19108,N_19149);
and UO_304 (O_304,N_19496,N_19353);
and UO_305 (O_305,N_19306,N_19911);
or UO_306 (O_306,N_19342,N_19103);
nor UO_307 (O_307,N_19379,N_19365);
xor UO_308 (O_308,N_19090,N_19703);
or UO_309 (O_309,N_19392,N_19542);
or UO_310 (O_310,N_19934,N_19262);
nor UO_311 (O_311,N_19126,N_19189);
and UO_312 (O_312,N_19600,N_19222);
or UO_313 (O_313,N_19155,N_19726);
nor UO_314 (O_314,N_19639,N_19217);
and UO_315 (O_315,N_19976,N_19776);
nor UO_316 (O_316,N_19467,N_19605);
nand UO_317 (O_317,N_19315,N_19383);
nor UO_318 (O_318,N_19945,N_19804);
xnor UO_319 (O_319,N_19913,N_19870);
and UO_320 (O_320,N_19034,N_19470);
nor UO_321 (O_321,N_19206,N_19592);
and UO_322 (O_322,N_19417,N_19505);
and UO_323 (O_323,N_19486,N_19418);
and UO_324 (O_324,N_19573,N_19456);
and UO_325 (O_325,N_19026,N_19038);
or UO_326 (O_326,N_19714,N_19348);
xnor UO_327 (O_327,N_19113,N_19195);
xnor UO_328 (O_328,N_19623,N_19218);
and UO_329 (O_329,N_19841,N_19679);
and UO_330 (O_330,N_19373,N_19491);
nand UO_331 (O_331,N_19863,N_19652);
and UO_332 (O_332,N_19766,N_19272);
xnor UO_333 (O_333,N_19139,N_19587);
and UO_334 (O_334,N_19936,N_19067);
xor UO_335 (O_335,N_19044,N_19707);
nand UO_336 (O_336,N_19347,N_19818);
nor UO_337 (O_337,N_19837,N_19242);
and UO_338 (O_338,N_19635,N_19786);
or UO_339 (O_339,N_19606,N_19941);
nand UO_340 (O_340,N_19097,N_19156);
and UO_341 (O_341,N_19932,N_19078);
nor UO_342 (O_342,N_19307,N_19281);
xnor UO_343 (O_343,N_19912,N_19181);
xor UO_344 (O_344,N_19050,N_19363);
and UO_345 (O_345,N_19209,N_19172);
nand UO_346 (O_346,N_19951,N_19510);
nor UO_347 (O_347,N_19921,N_19731);
xor UO_348 (O_348,N_19225,N_19759);
nor UO_349 (O_349,N_19585,N_19073);
or UO_350 (O_350,N_19249,N_19551);
nand UO_351 (O_351,N_19201,N_19374);
or UO_352 (O_352,N_19582,N_19046);
nand UO_353 (O_353,N_19677,N_19059);
or UO_354 (O_354,N_19949,N_19266);
nand UO_355 (O_355,N_19350,N_19797);
nor UO_356 (O_356,N_19292,N_19093);
and UO_357 (O_357,N_19371,N_19891);
or UO_358 (O_358,N_19835,N_19944);
nor UO_359 (O_359,N_19998,N_19782);
xor UO_360 (O_360,N_19741,N_19558);
nand UO_361 (O_361,N_19586,N_19430);
nand UO_362 (O_362,N_19011,N_19987);
nor UO_363 (O_363,N_19937,N_19212);
nor UO_364 (O_364,N_19360,N_19578);
nand UO_365 (O_365,N_19812,N_19962);
and UO_366 (O_366,N_19319,N_19765);
nand UO_367 (O_367,N_19711,N_19314);
nand UO_368 (O_368,N_19866,N_19056);
or UO_369 (O_369,N_19512,N_19556);
nor UO_370 (O_370,N_19328,N_19492);
xor UO_371 (O_371,N_19988,N_19691);
and UO_372 (O_372,N_19410,N_19612);
and UO_373 (O_373,N_19118,N_19419);
nor UO_374 (O_374,N_19648,N_19706);
nor UO_375 (O_375,N_19712,N_19393);
or UO_376 (O_376,N_19057,N_19445);
xnor UO_377 (O_377,N_19061,N_19527);
nor UO_378 (O_378,N_19015,N_19653);
or UO_379 (O_379,N_19048,N_19828);
nand UO_380 (O_380,N_19541,N_19356);
and UO_381 (O_381,N_19231,N_19756);
nor UO_382 (O_382,N_19920,N_19994);
nand UO_383 (O_383,N_19919,N_19601);
nor UO_384 (O_384,N_19141,N_19027);
nand UO_385 (O_385,N_19880,N_19947);
or UO_386 (O_386,N_19727,N_19174);
and UO_387 (O_387,N_19458,N_19982);
and UO_388 (O_388,N_19447,N_19901);
or UO_389 (O_389,N_19384,N_19167);
nor UO_390 (O_390,N_19925,N_19362);
or UO_391 (O_391,N_19772,N_19084);
or UO_392 (O_392,N_19784,N_19771);
xnor UO_393 (O_393,N_19117,N_19124);
nor UO_394 (O_394,N_19376,N_19740);
nor UO_395 (O_395,N_19518,N_19710);
nor UO_396 (O_396,N_19349,N_19228);
or UO_397 (O_397,N_19565,N_19528);
xnor UO_398 (O_398,N_19425,N_19675);
and UO_399 (O_399,N_19140,N_19519);
xnor UO_400 (O_400,N_19102,N_19211);
and UO_401 (O_401,N_19775,N_19525);
and UO_402 (O_402,N_19547,N_19614);
nor UO_403 (O_403,N_19898,N_19115);
nor UO_404 (O_404,N_19263,N_19545);
nand UO_405 (O_405,N_19597,N_19369);
or UO_406 (O_406,N_19716,N_19325);
and UO_407 (O_407,N_19205,N_19604);
nor UO_408 (O_408,N_19708,N_19794);
or UO_409 (O_409,N_19240,N_19781);
xor UO_410 (O_410,N_19754,N_19595);
xor UO_411 (O_411,N_19646,N_19602);
xor UO_412 (O_412,N_19079,N_19583);
nand UO_413 (O_413,N_19151,N_19862);
and UO_414 (O_414,N_19822,N_19304);
nand UO_415 (O_415,N_19523,N_19069);
nor UO_416 (O_416,N_19524,N_19009);
nand UO_417 (O_417,N_19111,N_19948);
nand UO_418 (O_418,N_19455,N_19903);
or UO_419 (O_419,N_19036,N_19873);
nor UO_420 (O_420,N_19485,N_19733);
nand UO_421 (O_421,N_19667,N_19555);
and UO_422 (O_422,N_19173,N_19133);
nor UO_423 (O_423,N_19332,N_19836);
nand UO_424 (O_424,N_19832,N_19354);
nor UO_425 (O_425,N_19621,N_19687);
xor UO_426 (O_426,N_19569,N_19950);
xnor UO_427 (O_427,N_19546,N_19366);
or UO_428 (O_428,N_19535,N_19625);
xor UO_429 (O_429,N_19907,N_19780);
xnor UO_430 (O_430,N_19464,N_19436);
nor UO_431 (O_431,N_19021,N_19568);
xor UO_432 (O_432,N_19268,N_19851);
and UO_433 (O_433,N_19823,N_19381);
xor UO_434 (O_434,N_19642,N_19448);
nor UO_435 (O_435,N_19276,N_19664);
or UO_436 (O_436,N_19734,N_19719);
and UO_437 (O_437,N_19296,N_19514);
nand UO_438 (O_438,N_19554,N_19788);
or UO_439 (O_439,N_19098,N_19005);
xor UO_440 (O_440,N_19704,N_19022);
and UO_441 (O_441,N_19132,N_19235);
or UO_442 (O_442,N_19375,N_19763);
nor UO_443 (O_443,N_19539,N_19404);
xnor UO_444 (O_444,N_19045,N_19377);
nor UO_445 (O_445,N_19397,N_19109);
nand UO_446 (O_446,N_19659,N_19223);
nand UO_447 (O_447,N_19562,N_19471);
nand UO_448 (O_448,N_19844,N_19899);
nor UO_449 (O_449,N_19840,N_19584);
or UO_450 (O_450,N_19479,N_19160);
xnor UO_451 (O_451,N_19650,N_19738);
nand UO_452 (O_452,N_19572,N_19735);
nor UO_453 (O_453,N_19689,N_19943);
nand UO_454 (O_454,N_19855,N_19087);
or UO_455 (O_455,N_19469,N_19910);
xor UO_456 (O_456,N_19129,N_19477);
nand UO_457 (O_457,N_19248,N_19101);
nand UO_458 (O_458,N_19459,N_19792);
and UO_459 (O_459,N_19053,N_19125);
nand UO_460 (O_460,N_19391,N_19918);
or UO_461 (O_461,N_19666,N_19579);
nor UO_462 (O_462,N_19858,N_19446);
xor UO_463 (O_463,N_19423,N_19136);
xnor UO_464 (O_464,N_19024,N_19076);
nand UO_465 (O_465,N_19070,N_19517);
nor UO_466 (O_466,N_19956,N_19494);
nor UO_467 (O_467,N_19671,N_19475);
nand UO_468 (O_468,N_19273,N_19917);
xor UO_469 (O_469,N_19874,N_19438);
or UO_470 (O_470,N_19186,N_19615);
nor UO_471 (O_471,N_19526,N_19807);
or UO_472 (O_472,N_19914,N_19931);
and UO_473 (O_473,N_19025,N_19853);
and UO_474 (O_474,N_19415,N_19435);
xnor UO_475 (O_475,N_19885,N_19216);
nand UO_476 (O_476,N_19408,N_19094);
nor UO_477 (O_477,N_19146,N_19355);
nor UO_478 (O_478,N_19345,N_19042);
or UO_479 (O_479,N_19540,N_19000);
or UO_480 (O_480,N_19386,N_19454);
or UO_481 (O_481,N_19032,N_19506);
or UO_482 (O_482,N_19254,N_19052);
or UO_483 (O_483,N_19030,N_19657);
xor UO_484 (O_484,N_19388,N_19848);
nor UO_485 (O_485,N_19008,N_19095);
nor UO_486 (O_486,N_19313,N_19968);
xnor UO_487 (O_487,N_19611,N_19890);
and UO_488 (O_488,N_19043,N_19954);
or UO_489 (O_489,N_19481,N_19434);
xor UO_490 (O_490,N_19544,N_19593);
or UO_491 (O_491,N_19897,N_19152);
or UO_492 (O_492,N_19682,N_19466);
nor UO_493 (O_493,N_19808,N_19199);
nand UO_494 (O_494,N_19878,N_19134);
nor UO_495 (O_495,N_19594,N_19616);
xor UO_496 (O_496,N_19020,N_19843);
and UO_497 (O_497,N_19610,N_19867);
xnor UO_498 (O_498,N_19357,N_19278);
nor UO_499 (O_499,N_19581,N_19104);
xor UO_500 (O_500,N_19134,N_19101);
xnor UO_501 (O_501,N_19666,N_19939);
nor UO_502 (O_502,N_19526,N_19236);
or UO_503 (O_503,N_19984,N_19454);
xor UO_504 (O_504,N_19888,N_19871);
nand UO_505 (O_505,N_19669,N_19800);
nand UO_506 (O_506,N_19867,N_19882);
nor UO_507 (O_507,N_19053,N_19055);
nor UO_508 (O_508,N_19835,N_19167);
and UO_509 (O_509,N_19918,N_19304);
xnor UO_510 (O_510,N_19648,N_19757);
or UO_511 (O_511,N_19193,N_19251);
nand UO_512 (O_512,N_19423,N_19168);
or UO_513 (O_513,N_19627,N_19646);
nor UO_514 (O_514,N_19595,N_19381);
and UO_515 (O_515,N_19812,N_19820);
xnor UO_516 (O_516,N_19981,N_19034);
and UO_517 (O_517,N_19174,N_19102);
and UO_518 (O_518,N_19663,N_19751);
and UO_519 (O_519,N_19364,N_19001);
and UO_520 (O_520,N_19716,N_19746);
xnor UO_521 (O_521,N_19625,N_19154);
nand UO_522 (O_522,N_19959,N_19429);
nor UO_523 (O_523,N_19511,N_19081);
and UO_524 (O_524,N_19874,N_19635);
and UO_525 (O_525,N_19631,N_19486);
xor UO_526 (O_526,N_19478,N_19267);
and UO_527 (O_527,N_19054,N_19916);
nor UO_528 (O_528,N_19656,N_19751);
nor UO_529 (O_529,N_19013,N_19791);
nand UO_530 (O_530,N_19232,N_19540);
nand UO_531 (O_531,N_19032,N_19156);
and UO_532 (O_532,N_19627,N_19271);
xor UO_533 (O_533,N_19511,N_19499);
nand UO_534 (O_534,N_19880,N_19410);
nor UO_535 (O_535,N_19809,N_19605);
and UO_536 (O_536,N_19171,N_19188);
xor UO_537 (O_537,N_19322,N_19613);
xor UO_538 (O_538,N_19635,N_19784);
nor UO_539 (O_539,N_19217,N_19926);
xor UO_540 (O_540,N_19445,N_19038);
and UO_541 (O_541,N_19130,N_19222);
or UO_542 (O_542,N_19874,N_19757);
and UO_543 (O_543,N_19583,N_19314);
and UO_544 (O_544,N_19960,N_19715);
nor UO_545 (O_545,N_19091,N_19605);
xor UO_546 (O_546,N_19726,N_19572);
nor UO_547 (O_547,N_19728,N_19255);
nor UO_548 (O_548,N_19407,N_19739);
and UO_549 (O_549,N_19475,N_19139);
nor UO_550 (O_550,N_19051,N_19438);
or UO_551 (O_551,N_19079,N_19848);
nor UO_552 (O_552,N_19792,N_19508);
or UO_553 (O_553,N_19957,N_19685);
nor UO_554 (O_554,N_19981,N_19350);
nor UO_555 (O_555,N_19838,N_19249);
xnor UO_556 (O_556,N_19832,N_19851);
nand UO_557 (O_557,N_19292,N_19127);
nand UO_558 (O_558,N_19567,N_19306);
or UO_559 (O_559,N_19700,N_19514);
nor UO_560 (O_560,N_19194,N_19963);
nand UO_561 (O_561,N_19655,N_19625);
or UO_562 (O_562,N_19642,N_19991);
or UO_563 (O_563,N_19083,N_19753);
nor UO_564 (O_564,N_19225,N_19160);
nand UO_565 (O_565,N_19056,N_19280);
nand UO_566 (O_566,N_19694,N_19209);
nand UO_567 (O_567,N_19028,N_19332);
and UO_568 (O_568,N_19977,N_19878);
xnor UO_569 (O_569,N_19510,N_19531);
nor UO_570 (O_570,N_19382,N_19250);
or UO_571 (O_571,N_19500,N_19120);
xnor UO_572 (O_572,N_19760,N_19594);
nand UO_573 (O_573,N_19885,N_19766);
or UO_574 (O_574,N_19458,N_19193);
nand UO_575 (O_575,N_19815,N_19836);
nand UO_576 (O_576,N_19870,N_19344);
and UO_577 (O_577,N_19452,N_19451);
xor UO_578 (O_578,N_19211,N_19721);
xnor UO_579 (O_579,N_19804,N_19308);
nand UO_580 (O_580,N_19687,N_19445);
or UO_581 (O_581,N_19927,N_19284);
nand UO_582 (O_582,N_19898,N_19182);
nor UO_583 (O_583,N_19570,N_19562);
xor UO_584 (O_584,N_19264,N_19573);
xnor UO_585 (O_585,N_19536,N_19558);
and UO_586 (O_586,N_19499,N_19633);
nand UO_587 (O_587,N_19355,N_19751);
xnor UO_588 (O_588,N_19973,N_19071);
xor UO_589 (O_589,N_19836,N_19561);
or UO_590 (O_590,N_19156,N_19056);
xnor UO_591 (O_591,N_19458,N_19159);
nor UO_592 (O_592,N_19982,N_19776);
nor UO_593 (O_593,N_19721,N_19542);
nand UO_594 (O_594,N_19559,N_19688);
and UO_595 (O_595,N_19830,N_19398);
and UO_596 (O_596,N_19715,N_19653);
nor UO_597 (O_597,N_19360,N_19678);
and UO_598 (O_598,N_19564,N_19996);
nor UO_599 (O_599,N_19459,N_19547);
nand UO_600 (O_600,N_19142,N_19555);
or UO_601 (O_601,N_19099,N_19526);
nor UO_602 (O_602,N_19627,N_19041);
xor UO_603 (O_603,N_19689,N_19089);
or UO_604 (O_604,N_19580,N_19953);
and UO_605 (O_605,N_19413,N_19978);
xnor UO_606 (O_606,N_19510,N_19746);
nand UO_607 (O_607,N_19461,N_19679);
or UO_608 (O_608,N_19888,N_19874);
and UO_609 (O_609,N_19503,N_19955);
or UO_610 (O_610,N_19816,N_19091);
nor UO_611 (O_611,N_19447,N_19526);
xor UO_612 (O_612,N_19073,N_19113);
nand UO_613 (O_613,N_19551,N_19485);
and UO_614 (O_614,N_19913,N_19030);
nand UO_615 (O_615,N_19286,N_19667);
xnor UO_616 (O_616,N_19770,N_19293);
nand UO_617 (O_617,N_19811,N_19477);
or UO_618 (O_618,N_19821,N_19336);
xor UO_619 (O_619,N_19934,N_19349);
and UO_620 (O_620,N_19503,N_19751);
and UO_621 (O_621,N_19198,N_19679);
nand UO_622 (O_622,N_19332,N_19574);
xnor UO_623 (O_623,N_19608,N_19669);
xnor UO_624 (O_624,N_19014,N_19179);
xor UO_625 (O_625,N_19440,N_19567);
xor UO_626 (O_626,N_19019,N_19071);
xor UO_627 (O_627,N_19504,N_19124);
nand UO_628 (O_628,N_19998,N_19382);
or UO_629 (O_629,N_19903,N_19579);
nor UO_630 (O_630,N_19924,N_19884);
nor UO_631 (O_631,N_19562,N_19192);
or UO_632 (O_632,N_19177,N_19295);
xnor UO_633 (O_633,N_19031,N_19509);
nand UO_634 (O_634,N_19378,N_19568);
nor UO_635 (O_635,N_19666,N_19176);
nor UO_636 (O_636,N_19496,N_19224);
or UO_637 (O_637,N_19567,N_19258);
nand UO_638 (O_638,N_19784,N_19400);
xnor UO_639 (O_639,N_19986,N_19587);
and UO_640 (O_640,N_19215,N_19405);
nor UO_641 (O_641,N_19191,N_19371);
xor UO_642 (O_642,N_19421,N_19686);
and UO_643 (O_643,N_19971,N_19579);
xnor UO_644 (O_644,N_19042,N_19417);
nor UO_645 (O_645,N_19518,N_19171);
xor UO_646 (O_646,N_19081,N_19688);
nor UO_647 (O_647,N_19237,N_19986);
nand UO_648 (O_648,N_19897,N_19061);
and UO_649 (O_649,N_19176,N_19968);
and UO_650 (O_650,N_19499,N_19732);
xor UO_651 (O_651,N_19819,N_19414);
or UO_652 (O_652,N_19639,N_19136);
nor UO_653 (O_653,N_19303,N_19045);
nor UO_654 (O_654,N_19665,N_19938);
nor UO_655 (O_655,N_19127,N_19330);
or UO_656 (O_656,N_19212,N_19175);
nand UO_657 (O_657,N_19891,N_19619);
or UO_658 (O_658,N_19557,N_19852);
xnor UO_659 (O_659,N_19038,N_19056);
and UO_660 (O_660,N_19198,N_19401);
or UO_661 (O_661,N_19656,N_19163);
or UO_662 (O_662,N_19354,N_19415);
nor UO_663 (O_663,N_19164,N_19734);
nand UO_664 (O_664,N_19821,N_19089);
or UO_665 (O_665,N_19246,N_19194);
and UO_666 (O_666,N_19100,N_19307);
and UO_667 (O_667,N_19130,N_19984);
xor UO_668 (O_668,N_19310,N_19171);
nor UO_669 (O_669,N_19262,N_19045);
nor UO_670 (O_670,N_19341,N_19199);
nand UO_671 (O_671,N_19127,N_19771);
nand UO_672 (O_672,N_19993,N_19709);
and UO_673 (O_673,N_19122,N_19123);
nor UO_674 (O_674,N_19558,N_19977);
and UO_675 (O_675,N_19100,N_19695);
nor UO_676 (O_676,N_19061,N_19080);
or UO_677 (O_677,N_19231,N_19921);
xor UO_678 (O_678,N_19561,N_19390);
and UO_679 (O_679,N_19165,N_19724);
xor UO_680 (O_680,N_19354,N_19448);
xnor UO_681 (O_681,N_19250,N_19830);
nand UO_682 (O_682,N_19867,N_19447);
and UO_683 (O_683,N_19615,N_19049);
or UO_684 (O_684,N_19602,N_19506);
and UO_685 (O_685,N_19843,N_19826);
or UO_686 (O_686,N_19081,N_19092);
xor UO_687 (O_687,N_19015,N_19409);
xnor UO_688 (O_688,N_19399,N_19276);
nand UO_689 (O_689,N_19049,N_19352);
nand UO_690 (O_690,N_19409,N_19328);
nand UO_691 (O_691,N_19954,N_19497);
xor UO_692 (O_692,N_19555,N_19519);
nand UO_693 (O_693,N_19411,N_19694);
or UO_694 (O_694,N_19043,N_19484);
xor UO_695 (O_695,N_19043,N_19105);
or UO_696 (O_696,N_19353,N_19498);
and UO_697 (O_697,N_19408,N_19537);
nor UO_698 (O_698,N_19557,N_19820);
and UO_699 (O_699,N_19291,N_19808);
or UO_700 (O_700,N_19455,N_19117);
and UO_701 (O_701,N_19089,N_19503);
nor UO_702 (O_702,N_19217,N_19885);
and UO_703 (O_703,N_19682,N_19722);
nor UO_704 (O_704,N_19304,N_19764);
nor UO_705 (O_705,N_19019,N_19652);
nor UO_706 (O_706,N_19825,N_19520);
nand UO_707 (O_707,N_19755,N_19814);
xor UO_708 (O_708,N_19685,N_19021);
or UO_709 (O_709,N_19964,N_19413);
nor UO_710 (O_710,N_19300,N_19128);
nand UO_711 (O_711,N_19966,N_19806);
or UO_712 (O_712,N_19680,N_19765);
nand UO_713 (O_713,N_19415,N_19787);
nand UO_714 (O_714,N_19861,N_19828);
or UO_715 (O_715,N_19334,N_19181);
nand UO_716 (O_716,N_19014,N_19499);
nand UO_717 (O_717,N_19428,N_19334);
xor UO_718 (O_718,N_19326,N_19459);
nand UO_719 (O_719,N_19325,N_19718);
nand UO_720 (O_720,N_19172,N_19316);
nand UO_721 (O_721,N_19646,N_19194);
nand UO_722 (O_722,N_19305,N_19958);
nand UO_723 (O_723,N_19355,N_19053);
and UO_724 (O_724,N_19089,N_19964);
or UO_725 (O_725,N_19646,N_19226);
xor UO_726 (O_726,N_19057,N_19023);
nor UO_727 (O_727,N_19453,N_19379);
and UO_728 (O_728,N_19984,N_19109);
nand UO_729 (O_729,N_19718,N_19884);
or UO_730 (O_730,N_19947,N_19308);
nand UO_731 (O_731,N_19180,N_19971);
or UO_732 (O_732,N_19694,N_19006);
and UO_733 (O_733,N_19950,N_19406);
nor UO_734 (O_734,N_19340,N_19253);
nand UO_735 (O_735,N_19015,N_19524);
nand UO_736 (O_736,N_19580,N_19126);
xor UO_737 (O_737,N_19567,N_19529);
or UO_738 (O_738,N_19155,N_19079);
and UO_739 (O_739,N_19404,N_19750);
or UO_740 (O_740,N_19570,N_19596);
nor UO_741 (O_741,N_19026,N_19889);
nor UO_742 (O_742,N_19601,N_19825);
nand UO_743 (O_743,N_19542,N_19152);
nand UO_744 (O_744,N_19893,N_19619);
nor UO_745 (O_745,N_19177,N_19947);
nand UO_746 (O_746,N_19092,N_19937);
or UO_747 (O_747,N_19376,N_19350);
or UO_748 (O_748,N_19275,N_19219);
nand UO_749 (O_749,N_19883,N_19849);
and UO_750 (O_750,N_19231,N_19827);
xnor UO_751 (O_751,N_19572,N_19791);
nor UO_752 (O_752,N_19932,N_19826);
and UO_753 (O_753,N_19228,N_19922);
nand UO_754 (O_754,N_19770,N_19964);
or UO_755 (O_755,N_19101,N_19703);
and UO_756 (O_756,N_19373,N_19134);
xor UO_757 (O_757,N_19385,N_19845);
xnor UO_758 (O_758,N_19678,N_19382);
xnor UO_759 (O_759,N_19564,N_19609);
nand UO_760 (O_760,N_19759,N_19486);
and UO_761 (O_761,N_19871,N_19215);
or UO_762 (O_762,N_19778,N_19288);
and UO_763 (O_763,N_19517,N_19398);
xnor UO_764 (O_764,N_19958,N_19026);
xor UO_765 (O_765,N_19547,N_19738);
and UO_766 (O_766,N_19667,N_19481);
xnor UO_767 (O_767,N_19685,N_19439);
xnor UO_768 (O_768,N_19986,N_19105);
xnor UO_769 (O_769,N_19401,N_19006);
xor UO_770 (O_770,N_19693,N_19270);
xnor UO_771 (O_771,N_19832,N_19615);
xnor UO_772 (O_772,N_19604,N_19899);
and UO_773 (O_773,N_19078,N_19253);
and UO_774 (O_774,N_19432,N_19290);
nor UO_775 (O_775,N_19856,N_19989);
or UO_776 (O_776,N_19121,N_19831);
nor UO_777 (O_777,N_19234,N_19151);
and UO_778 (O_778,N_19333,N_19371);
xnor UO_779 (O_779,N_19107,N_19069);
xor UO_780 (O_780,N_19853,N_19785);
or UO_781 (O_781,N_19463,N_19953);
nand UO_782 (O_782,N_19449,N_19190);
xor UO_783 (O_783,N_19637,N_19476);
and UO_784 (O_784,N_19247,N_19644);
and UO_785 (O_785,N_19723,N_19300);
or UO_786 (O_786,N_19024,N_19514);
and UO_787 (O_787,N_19927,N_19388);
and UO_788 (O_788,N_19941,N_19449);
or UO_789 (O_789,N_19795,N_19713);
nand UO_790 (O_790,N_19248,N_19738);
xor UO_791 (O_791,N_19656,N_19568);
xnor UO_792 (O_792,N_19544,N_19053);
nand UO_793 (O_793,N_19056,N_19000);
or UO_794 (O_794,N_19774,N_19652);
or UO_795 (O_795,N_19164,N_19063);
xor UO_796 (O_796,N_19547,N_19418);
xor UO_797 (O_797,N_19545,N_19133);
nor UO_798 (O_798,N_19713,N_19929);
nor UO_799 (O_799,N_19213,N_19831);
or UO_800 (O_800,N_19982,N_19435);
nor UO_801 (O_801,N_19134,N_19144);
and UO_802 (O_802,N_19661,N_19414);
nor UO_803 (O_803,N_19344,N_19696);
nor UO_804 (O_804,N_19284,N_19577);
xnor UO_805 (O_805,N_19847,N_19952);
xnor UO_806 (O_806,N_19822,N_19383);
nor UO_807 (O_807,N_19655,N_19177);
or UO_808 (O_808,N_19763,N_19146);
and UO_809 (O_809,N_19848,N_19277);
nand UO_810 (O_810,N_19230,N_19220);
nand UO_811 (O_811,N_19122,N_19033);
and UO_812 (O_812,N_19200,N_19717);
nor UO_813 (O_813,N_19167,N_19799);
xnor UO_814 (O_814,N_19703,N_19375);
xor UO_815 (O_815,N_19101,N_19129);
nor UO_816 (O_816,N_19351,N_19590);
or UO_817 (O_817,N_19971,N_19001);
or UO_818 (O_818,N_19254,N_19363);
xor UO_819 (O_819,N_19244,N_19167);
xor UO_820 (O_820,N_19368,N_19819);
nor UO_821 (O_821,N_19912,N_19620);
nand UO_822 (O_822,N_19824,N_19126);
or UO_823 (O_823,N_19438,N_19314);
nor UO_824 (O_824,N_19501,N_19069);
or UO_825 (O_825,N_19254,N_19290);
or UO_826 (O_826,N_19455,N_19244);
and UO_827 (O_827,N_19136,N_19743);
nor UO_828 (O_828,N_19020,N_19961);
nor UO_829 (O_829,N_19463,N_19837);
nand UO_830 (O_830,N_19018,N_19336);
and UO_831 (O_831,N_19980,N_19812);
or UO_832 (O_832,N_19416,N_19230);
xnor UO_833 (O_833,N_19358,N_19349);
nand UO_834 (O_834,N_19089,N_19487);
and UO_835 (O_835,N_19231,N_19165);
nor UO_836 (O_836,N_19648,N_19068);
nor UO_837 (O_837,N_19969,N_19376);
and UO_838 (O_838,N_19661,N_19276);
nand UO_839 (O_839,N_19990,N_19802);
nand UO_840 (O_840,N_19888,N_19451);
nor UO_841 (O_841,N_19652,N_19139);
and UO_842 (O_842,N_19841,N_19604);
or UO_843 (O_843,N_19983,N_19388);
nor UO_844 (O_844,N_19247,N_19624);
xor UO_845 (O_845,N_19461,N_19277);
and UO_846 (O_846,N_19729,N_19869);
nand UO_847 (O_847,N_19123,N_19915);
nand UO_848 (O_848,N_19248,N_19001);
or UO_849 (O_849,N_19281,N_19595);
and UO_850 (O_850,N_19078,N_19929);
or UO_851 (O_851,N_19912,N_19238);
and UO_852 (O_852,N_19254,N_19732);
nand UO_853 (O_853,N_19483,N_19358);
nor UO_854 (O_854,N_19173,N_19294);
xor UO_855 (O_855,N_19432,N_19043);
nor UO_856 (O_856,N_19553,N_19867);
or UO_857 (O_857,N_19067,N_19780);
or UO_858 (O_858,N_19585,N_19379);
nand UO_859 (O_859,N_19308,N_19530);
xnor UO_860 (O_860,N_19854,N_19457);
xnor UO_861 (O_861,N_19485,N_19373);
and UO_862 (O_862,N_19089,N_19003);
xor UO_863 (O_863,N_19817,N_19135);
xor UO_864 (O_864,N_19342,N_19499);
and UO_865 (O_865,N_19270,N_19026);
and UO_866 (O_866,N_19739,N_19016);
nand UO_867 (O_867,N_19256,N_19588);
nand UO_868 (O_868,N_19604,N_19916);
nand UO_869 (O_869,N_19825,N_19853);
or UO_870 (O_870,N_19203,N_19829);
or UO_871 (O_871,N_19114,N_19661);
nand UO_872 (O_872,N_19215,N_19043);
xnor UO_873 (O_873,N_19493,N_19483);
nand UO_874 (O_874,N_19824,N_19878);
or UO_875 (O_875,N_19174,N_19982);
or UO_876 (O_876,N_19311,N_19251);
xor UO_877 (O_877,N_19712,N_19798);
xor UO_878 (O_878,N_19581,N_19506);
nor UO_879 (O_879,N_19523,N_19482);
nand UO_880 (O_880,N_19675,N_19165);
nor UO_881 (O_881,N_19131,N_19238);
nand UO_882 (O_882,N_19520,N_19035);
xor UO_883 (O_883,N_19289,N_19422);
or UO_884 (O_884,N_19304,N_19317);
or UO_885 (O_885,N_19645,N_19114);
xor UO_886 (O_886,N_19554,N_19861);
nor UO_887 (O_887,N_19491,N_19006);
xor UO_888 (O_888,N_19684,N_19609);
xor UO_889 (O_889,N_19385,N_19694);
or UO_890 (O_890,N_19507,N_19913);
xor UO_891 (O_891,N_19064,N_19918);
nor UO_892 (O_892,N_19758,N_19170);
xnor UO_893 (O_893,N_19007,N_19909);
or UO_894 (O_894,N_19398,N_19202);
or UO_895 (O_895,N_19375,N_19808);
nor UO_896 (O_896,N_19120,N_19070);
xnor UO_897 (O_897,N_19053,N_19452);
and UO_898 (O_898,N_19342,N_19060);
or UO_899 (O_899,N_19403,N_19841);
nand UO_900 (O_900,N_19222,N_19335);
or UO_901 (O_901,N_19505,N_19454);
or UO_902 (O_902,N_19320,N_19809);
nand UO_903 (O_903,N_19145,N_19270);
or UO_904 (O_904,N_19818,N_19844);
nand UO_905 (O_905,N_19620,N_19543);
xor UO_906 (O_906,N_19640,N_19463);
and UO_907 (O_907,N_19629,N_19154);
nor UO_908 (O_908,N_19323,N_19636);
nand UO_909 (O_909,N_19908,N_19107);
nand UO_910 (O_910,N_19136,N_19850);
nand UO_911 (O_911,N_19157,N_19707);
or UO_912 (O_912,N_19150,N_19134);
nor UO_913 (O_913,N_19184,N_19502);
xor UO_914 (O_914,N_19510,N_19774);
nor UO_915 (O_915,N_19669,N_19712);
nand UO_916 (O_916,N_19478,N_19586);
and UO_917 (O_917,N_19267,N_19510);
nor UO_918 (O_918,N_19013,N_19533);
nor UO_919 (O_919,N_19142,N_19995);
nor UO_920 (O_920,N_19223,N_19140);
or UO_921 (O_921,N_19731,N_19716);
nand UO_922 (O_922,N_19702,N_19587);
xnor UO_923 (O_923,N_19922,N_19711);
xor UO_924 (O_924,N_19319,N_19687);
or UO_925 (O_925,N_19493,N_19691);
or UO_926 (O_926,N_19280,N_19953);
nor UO_927 (O_927,N_19938,N_19622);
nand UO_928 (O_928,N_19532,N_19609);
xnor UO_929 (O_929,N_19702,N_19520);
and UO_930 (O_930,N_19678,N_19818);
nor UO_931 (O_931,N_19691,N_19008);
and UO_932 (O_932,N_19438,N_19349);
nor UO_933 (O_933,N_19924,N_19361);
nor UO_934 (O_934,N_19721,N_19706);
or UO_935 (O_935,N_19427,N_19724);
nand UO_936 (O_936,N_19319,N_19961);
xnor UO_937 (O_937,N_19177,N_19468);
or UO_938 (O_938,N_19774,N_19313);
or UO_939 (O_939,N_19993,N_19156);
nor UO_940 (O_940,N_19739,N_19772);
nand UO_941 (O_941,N_19752,N_19712);
and UO_942 (O_942,N_19466,N_19434);
nand UO_943 (O_943,N_19772,N_19948);
nand UO_944 (O_944,N_19288,N_19491);
or UO_945 (O_945,N_19378,N_19779);
nor UO_946 (O_946,N_19454,N_19258);
and UO_947 (O_947,N_19606,N_19617);
nor UO_948 (O_948,N_19233,N_19461);
or UO_949 (O_949,N_19707,N_19488);
nor UO_950 (O_950,N_19972,N_19550);
nand UO_951 (O_951,N_19176,N_19761);
xor UO_952 (O_952,N_19539,N_19204);
xnor UO_953 (O_953,N_19472,N_19526);
or UO_954 (O_954,N_19616,N_19158);
nand UO_955 (O_955,N_19636,N_19717);
or UO_956 (O_956,N_19420,N_19442);
or UO_957 (O_957,N_19660,N_19763);
or UO_958 (O_958,N_19219,N_19963);
and UO_959 (O_959,N_19109,N_19167);
xnor UO_960 (O_960,N_19238,N_19237);
xor UO_961 (O_961,N_19655,N_19386);
nor UO_962 (O_962,N_19109,N_19836);
or UO_963 (O_963,N_19646,N_19536);
nor UO_964 (O_964,N_19833,N_19189);
xnor UO_965 (O_965,N_19498,N_19231);
and UO_966 (O_966,N_19845,N_19796);
xor UO_967 (O_967,N_19927,N_19646);
and UO_968 (O_968,N_19922,N_19058);
xor UO_969 (O_969,N_19760,N_19403);
nand UO_970 (O_970,N_19749,N_19240);
or UO_971 (O_971,N_19518,N_19324);
xor UO_972 (O_972,N_19584,N_19858);
nand UO_973 (O_973,N_19162,N_19355);
nor UO_974 (O_974,N_19502,N_19354);
or UO_975 (O_975,N_19560,N_19471);
nand UO_976 (O_976,N_19767,N_19506);
or UO_977 (O_977,N_19697,N_19867);
xnor UO_978 (O_978,N_19274,N_19393);
nand UO_979 (O_979,N_19189,N_19789);
nand UO_980 (O_980,N_19912,N_19417);
nor UO_981 (O_981,N_19792,N_19253);
nor UO_982 (O_982,N_19541,N_19401);
or UO_983 (O_983,N_19181,N_19484);
and UO_984 (O_984,N_19067,N_19297);
or UO_985 (O_985,N_19850,N_19338);
nand UO_986 (O_986,N_19271,N_19632);
and UO_987 (O_987,N_19362,N_19160);
nor UO_988 (O_988,N_19648,N_19299);
or UO_989 (O_989,N_19168,N_19666);
nor UO_990 (O_990,N_19415,N_19322);
nor UO_991 (O_991,N_19324,N_19770);
and UO_992 (O_992,N_19863,N_19903);
or UO_993 (O_993,N_19713,N_19142);
or UO_994 (O_994,N_19819,N_19723);
xnor UO_995 (O_995,N_19194,N_19597);
or UO_996 (O_996,N_19124,N_19456);
or UO_997 (O_997,N_19824,N_19283);
nand UO_998 (O_998,N_19467,N_19004);
nor UO_999 (O_999,N_19544,N_19888);
nand UO_1000 (O_1000,N_19197,N_19182);
nand UO_1001 (O_1001,N_19790,N_19675);
xor UO_1002 (O_1002,N_19365,N_19928);
nor UO_1003 (O_1003,N_19829,N_19331);
nor UO_1004 (O_1004,N_19555,N_19997);
or UO_1005 (O_1005,N_19055,N_19616);
xor UO_1006 (O_1006,N_19150,N_19870);
nor UO_1007 (O_1007,N_19354,N_19074);
nand UO_1008 (O_1008,N_19801,N_19738);
or UO_1009 (O_1009,N_19939,N_19556);
xor UO_1010 (O_1010,N_19799,N_19318);
and UO_1011 (O_1011,N_19782,N_19326);
and UO_1012 (O_1012,N_19158,N_19579);
and UO_1013 (O_1013,N_19179,N_19465);
xnor UO_1014 (O_1014,N_19678,N_19050);
and UO_1015 (O_1015,N_19635,N_19946);
and UO_1016 (O_1016,N_19362,N_19316);
nand UO_1017 (O_1017,N_19285,N_19158);
or UO_1018 (O_1018,N_19732,N_19392);
and UO_1019 (O_1019,N_19545,N_19141);
or UO_1020 (O_1020,N_19121,N_19647);
nor UO_1021 (O_1021,N_19914,N_19050);
or UO_1022 (O_1022,N_19392,N_19606);
and UO_1023 (O_1023,N_19792,N_19368);
nor UO_1024 (O_1024,N_19403,N_19204);
xor UO_1025 (O_1025,N_19838,N_19382);
nand UO_1026 (O_1026,N_19230,N_19222);
nor UO_1027 (O_1027,N_19582,N_19187);
nand UO_1028 (O_1028,N_19047,N_19116);
nand UO_1029 (O_1029,N_19810,N_19945);
and UO_1030 (O_1030,N_19880,N_19665);
or UO_1031 (O_1031,N_19566,N_19795);
xor UO_1032 (O_1032,N_19528,N_19024);
nand UO_1033 (O_1033,N_19627,N_19412);
or UO_1034 (O_1034,N_19457,N_19106);
xor UO_1035 (O_1035,N_19917,N_19020);
or UO_1036 (O_1036,N_19665,N_19998);
nor UO_1037 (O_1037,N_19954,N_19767);
nor UO_1038 (O_1038,N_19948,N_19221);
nand UO_1039 (O_1039,N_19220,N_19450);
xnor UO_1040 (O_1040,N_19410,N_19196);
nor UO_1041 (O_1041,N_19680,N_19204);
nand UO_1042 (O_1042,N_19209,N_19083);
nor UO_1043 (O_1043,N_19569,N_19123);
nand UO_1044 (O_1044,N_19261,N_19775);
xnor UO_1045 (O_1045,N_19454,N_19638);
nor UO_1046 (O_1046,N_19732,N_19561);
nand UO_1047 (O_1047,N_19899,N_19337);
nor UO_1048 (O_1048,N_19838,N_19348);
or UO_1049 (O_1049,N_19984,N_19463);
xor UO_1050 (O_1050,N_19977,N_19825);
nand UO_1051 (O_1051,N_19611,N_19964);
xnor UO_1052 (O_1052,N_19607,N_19366);
or UO_1053 (O_1053,N_19380,N_19739);
nand UO_1054 (O_1054,N_19843,N_19145);
nor UO_1055 (O_1055,N_19836,N_19249);
nor UO_1056 (O_1056,N_19741,N_19135);
nand UO_1057 (O_1057,N_19287,N_19588);
xnor UO_1058 (O_1058,N_19114,N_19025);
xor UO_1059 (O_1059,N_19259,N_19951);
or UO_1060 (O_1060,N_19537,N_19414);
or UO_1061 (O_1061,N_19206,N_19409);
nor UO_1062 (O_1062,N_19176,N_19533);
nor UO_1063 (O_1063,N_19136,N_19903);
xor UO_1064 (O_1064,N_19714,N_19587);
nand UO_1065 (O_1065,N_19050,N_19948);
and UO_1066 (O_1066,N_19581,N_19424);
nand UO_1067 (O_1067,N_19340,N_19373);
nand UO_1068 (O_1068,N_19336,N_19048);
nor UO_1069 (O_1069,N_19953,N_19059);
nand UO_1070 (O_1070,N_19024,N_19121);
nand UO_1071 (O_1071,N_19574,N_19441);
xnor UO_1072 (O_1072,N_19150,N_19033);
nand UO_1073 (O_1073,N_19335,N_19036);
nand UO_1074 (O_1074,N_19791,N_19787);
or UO_1075 (O_1075,N_19274,N_19203);
or UO_1076 (O_1076,N_19979,N_19429);
and UO_1077 (O_1077,N_19329,N_19009);
or UO_1078 (O_1078,N_19297,N_19750);
or UO_1079 (O_1079,N_19470,N_19919);
nor UO_1080 (O_1080,N_19118,N_19675);
nor UO_1081 (O_1081,N_19345,N_19769);
or UO_1082 (O_1082,N_19825,N_19639);
nand UO_1083 (O_1083,N_19893,N_19029);
nor UO_1084 (O_1084,N_19443,N_19709);
xnor UO_1085 (O_1085,N_19780,N_19339);
and UO_1086 (O_1086,N_19593,N_19691);
nand UO_1087 (O_1087,N_19331,N_19768);
and UO_1088 (O_1088,N_19310,N_19875);
or UO_1089 (O_1089,N_19944,N_19264);
nand UO_1090 (O_1090,N_19381,N_19826);
xnor UO_1091 (O_1091,N_19281,N_19620);
nand UO_1092 (O_1092,N_19313,N_19727);
or UO_1093 (O_1093,N_19332,N_19390);
xnor UO_1094 (O_1094,N_19145,N_19242);
xnor UO_1095 (O_1095,N_19968,N_19850);
and UO_1096 (O_1096,N_19827,N_19185);
or UO_1097 (O_1097,N_19550,N_19735);
and UO_1098 (O_1098,N_19673,N_19490);
or UO_1099 (O_1099,N_19910,N_19567);
or UO_1100 (O_1100,N_19327,N_19346);
and UO_1101 (O_1101,N_19099,N_19167);
xor UO_1102 (O_1102,N_19594,N_19740);
nor UO_1103 (O_1103,N_19639,N_19874);
xor UO_1104 (O_1104,N_19038,N_19110);
nor UO_1105 (O_1105,N_19679,N_19572);
nand UO_1106 (O_1106,N_19143,N_19534);
nor UO_1107 (O_1107,N_19445,N_19272);
or UO_1108 (O_1108,N_19895,N_19802);
nand UO_1109 (O_1109,N_19184,N_19495);
or UO_1110 (O_1110,N_19678,N_19085);
nor UO_1111 (O_1111,N_19817,N_19794);
xnor UO_1112 (O_1112,N_19180,N_19856);
and UO_1113 (O_1113,N_19813,N_19682);
or UO_1114 (O_1114,N_19093,N_19811);
or UO_1115 (O_1115,N_19065,N_19063);
xor UO_1116 (O_1116,N_19279,N_19310);
nor UO_1117 (O_1117,N_19838,N_19022);
or UO_1118 (O_1118,N_19307,N_19881);
and UO_1119 (O_1119,N_19065,N_19351);
nand UO_1120 (O_1120,N_19188,N_19693);
nor UO_1121 (O_1121,N_19882,N_19551);
xnor UO_1122 (O_1122,N_19649,N_19243);
nand UO_1123 (O_1123,N_19880,N_19208);
nor UO_1124 (O_1124,N_19403,N_19568);
or UO_1125 (O_1125,N_19602,N_19727);
nand UO_1126 (O_1126,N_19308,N_19912);
nor UO_1127 (O_1127,N_19154,N_19787);
and UO_1128 (O_1128,N_19868,N_19284);
and UO_1129 (O_1129,N_19965,N_19008);
xor UO_1130 (O_1130,N_19351,N_19195);
or UO_1131 (O_1131,N_19845,N_19480);
and UO_1132 (O_1132,N_19468,N_19759);
or UO_1133 (O_1133,N_19767,N_19066);
or UO_1134 (O_1134,N_19718,N_19867);
xnor UO_1135 (O_1135,N_19765,N_19766);
xnor UO_1136 (O_1136,N_19254,N_19566);
xor UO_1137 (O_1137,N_19718,N_19638);
nand UO_1138 (O_1138,N_19014,N_19529);
or UO_1139 (O_1139,N_19759,N_19921);
nand UO_1140 (O_1140,N_19285,N_19738);
or UO_1141 (O_1141,N_19428,N_19338);
and UO_1142 (O_1142,N_19436,N_19710);
nand UO_1143 (O_1143,N_19478,N_19853);
or UO_1144 (O_1144,N_19141,N_19348);
or UO_1145 (O_1145,N_19181,N_19299);
and UO_1146 (O_1146,N_19206,N_19270);
and UO_1147 (O_1147,N_19578,N_19100);
nor UO_1148 (O_1148,N_19505,N_19999);
nor UO_1149 (O_1149,N_19406,N_19627);
or UO_1150 (O_1150,N_19777,N_19089);
or UO_1151 (O_1151,N_19511,N_19708);
and UO_1152 (O_1152,N_19168,N_19798);
and UO_1153 (O_1153,N_19394,N_19091);
nand UO_1154 (O_1154,N_19903,N_19645);
nor UO_1155 (O_1155,N_19969,N_19862);
and UO_1156 (O_1156,N_19562,N_19126);
and UO_1157 (O_1157,N_19454,N_19113);
and UO_1158 (O_1158,N_19529,N_19908);
xnor UO_1159 (O_1159,N_19370,N_19584);
xor UO_1160 (O_1160,N_19871,N_19732);
xnor UO_1161 (O_1161,N_19408,N_19582);
and UO_1162 (O_1162,N_19395,N_19640);
nor UO_1163 (O_1163,N_19353,N_19692);
nor UO_1164 (O_1164,N_19780,N_19928);
or UO_1165 (O_1165,N_19734,N_19272);
nand UO_1166 (O_1166,N_19701,N_19143);
xor UO_1167 (O_1167,N_19883,N_19381);
xnor UO_1168 (O_1168,N_19706,N_19562);
nand UO_1169 (O_1169,N_19564,N_19230);
nor UO_1170 (O_1170,N_19543,N_19964);
nor UO_1171 (O_1171,N_19229,N_19904);
nor UO_1172 (O_1172,N_19991,N_19593);
and UO_1173 (O_1173,N_19968,N_19721);
xnor UO_1174 (O_1174,N_19601,N_19990);
nand UO_1175 (O_1175,N_19805,N_19834);
or UO_1176 (O_1176,N_19528,N_19144);
nand UO_1177 (O_1177,N_19462,N_19646);
or UO_1178 (O_1178,N_19333,N_19117);
or UO_1179 (O_1179,N_19933,N_19669);
or UO_1180 (O_1180,N_19394,N_19096);
nand UO_1181 (O_1181,N_19431,N_19707);
xor UO_1182 (O_1182,N_19181,N_19888);
or UO_1183 (O_1183,N_19668,N_19131);
nor UO_1184 (O_1184,N_19851,N_19541);
and UO_1185 (O_1185,N_19493,N_19586);
nand UO_1186 (O_1186,N_19348,N_19126);
xor UO_1187 (O_1187,N_19674,N_19765);
xor UO_1188 (O_1188,N_19872,N_19515);
and UO_1189 (O_1189,N_19814,N_19306);
or UO_1190 (O_1190,N_19843,N_19298);
and UO_1191 (O_1191,N_19278,N_19955);
nor UO_1192 (O_1192,N_19173,N_19274);
or UO_1193 (O_1193,N_19634,N_19474);
nor UO_1194 (O_1194,N_19558,N_19309);
xnor UO_1195 (O_1195,N_19010,N_19992);
and UO_1196 (O_1196,N_19445,N_19337);
nand UO_1197 (O_1197,N_19193,N_19159);
and UO_1198 (O_1198,N_19472,N_19047);
xor UO_1199 (O_1199,N_19209,N_19748);
xor UO_1200 (O_1200,N_19104,N_19329);
and UO_1201 (O_1201,N_19315,N_19809);
nand UO_1202 (O_1202,N_19051,N_19157);
nor UO_1203 (O_1203,N_19194,N_19753);
or UO_1204 (O_1204,N_19337,N_19878);
and UO_1205 (O_1205,N_19147,N_19837);
nand UO_1206 (O_1206,N_19534,N_19506);
nor UO_1207 (O_1207,N_19682,N_19867);
and UO_1208 (O_1208,N_19726,N_19404);
xnor UO_1209 (O_1209,N_19161,N_19993);
xnor UO_1210 (O_1210,N_19974,N_19266);
or UO_1211 (O_1211,N_19502,N_19086);
nand UO_1212 (O_1212,N_19262,N_19057);
xnor UO_1213 (O_1213,N_19237,N_19399);
or UO_1214 (O_1214,N_19380,N_19144);
nand UO_1215 (O_1215,N_19774,N_19099);
nor UO_1216 (O_1216,N_19098,N_19579);
nor UO_1217 (O_1217,N_19061,N_19282);
or UO_1218 (O_1218,N_19493,N_19947);
nor UO_1219 (O_1219,N_19403,N_19090);
xor UO_1220 (O_1220,N_19014,N_19773);
or UO_1221 (O_1221,N_19004,N_19448);
and UO_1222 (O_1222,N_19618,N_19110);
nand UO_1223 (O_1223,N_19849,N_19390);
or UO_1224 (O_1224,N_19626,N_19365);
nor UO_1225 (O_1225,N_19692,N_19348);
xnor UO_1226 (O_1226,N_19647,N_19412);
xor UO_1227 (O_1227,N_19239,N_19570);
or UO_1228 (O_1228,N_19989,N_19307);
nor UO_1229 (O_1229,N_19102,N_19656);
xor UO_1230 (O_1230,N_19403,N_19938);
and UO_1231 (O_1231,N_19794,N_19434);
nor UO_1232 (O_1232,N_19101,N_19554);
nand UO_1233 (O_1233,N_19502,N_19926);
nor UO_1234 (O_1234,N_19443,N_19872);
and UO_1235 (O_1235,N_19943,N_19754);
or UO_1236 (O_1236,N_19390,N_19290);
nand UO_1237 (O_1237,N_19107,N_19253);
xor UO_1238 (O_1238,N_19490,N_19449);
xnor UO_1239 (O_1239,N_19814,N_19392);
nor UO_1240 (O_1240,N_19995,N_19006);
or UO_1241 (O_1241,N_19483,N_19190);
nand UO_1242 (O_1242,N_19839,N_19430);
nand UO_1243 (O_1243,N_19514,N_19857);
nand UO_1244 (O_1244,N_19099,N_19235);
nor UO_1245 (O_1245,N_19766,N_19472);
xnor UO_1246 (O_1246,N_19687,N_19461);
nor UO_1247 (O_1247,N_19097,N_19972);
or UO_1248 (O_1248,N_19122,N_19603);
nor UO_1249 (O_1249,N_19831,N_19968);
xor UO_1250 (O_1250,N_19905,N_19535);
nand UO_1251 (O_1251,N_19050,N_19953);
and UO_1252 (O_1252,N_19161,N_19501);
and UO_1253 (O_1253,N_19981,N_19645);
and UO_1254 (O_1254,N_19004,N_19898);
nor UO_1255 (O_1255,N_19538,N_19977);
nor UO_1256 (O_1256,N_19179,N_19627);
nor UO_1257 (O_1257,N_19131,N_19886);
nor UO_1258 (O_1258,N_19870,N_19396);
xor UO_1259 (O_1259,N_19854,N_19618);
or UO_1260 (O_1260,N_19149,N_19428);
nand UO_1261 (O_1261,N_19371,N_19292);
and UO_1262 (O_1262,N_19361,N_19671);
and UO_1263 (O_1263,N_19767,N_19194);
nor UO_1264 (O_1264,N_19864,N_19107);
and UO_1265 (O_1265,N_19688,N_19671);
nor UO_1266 (O_1266,N_19998,N_19557);
or UO_1267 (O_1267,N_19479,N_19254);
or UO_1268 (O_1268,N_19590,N_19317);
nor UO_1269 (O_1269,N_19109,N_19022);
nand UO_1270 (O_1270,N_19696,N_19777);
nor UO_1271 (O_1271,N_19418,N_19166);
and UO_1272 (O_1272,N_19648,N_19179);
nor UO_1273 (O_1273,N_19340,N_19085);
xnor UO_1274 (O_1274,N_19411,N_19506);
and UO_1275 (O_1275,N_19856,N_19298);
xor UO_1276 (O_1276,N_19029,N_19382);
and UO_1277 (O_1277,N_19112,N_19938);
and UO_1278 (O_1278,N_19894,N_19856);
nor UO_1279 (O_1279,N_19480,N_19379);
or UO_1280 (O_1280,N_19377,N_19102);
xor UO_1281 (O_1281,N_19096,N_19698);
nor UO_1282 (O_1282,N_19049,N_19018);
nor UO_1283 (O_1283,N_19788,N_19854);
or UO_1284 (O_1284,N_19146,N_19063);
or UO_1285 (O_1285,N_19412,N_19925);
or UO_1286 (O_1286,N_19130,N_19945);
or UO_1287 (O_1287,N_19181,N_19453);
and UO_1288 (O_1288,N_19007,N_19870);
and UO_1289 (O_1289,N_19978,N_19600);
or UO_1290 (O_1290,N_19911,N_19964);
or UO_1291 (O_1291,N_19851,N_19406);
or UO_1292 (O_1292,N_19381,N_19391);
or UO_1293 (O_1293,N_19733,N_19189);
and UO_1294 (O_1294,N_19430,N_19299);
and UO_1295 (O_1295,N_19543,N_19725);
nand UO_1296 (O_1296,N_19716,N_19604);
or UO_1297 (O_1297,N_19727,N_19592);
xor UO_1298 (O_1298,N_19877,N_19261);
nor UO_1299 (O_1299,N_19845,N_19280);
and UO_1300 (O_1300,N_19391,N_19596);
xor UO_1301 (O_1301,N_19134,N_19183);
nand UO_1302 (O_1302,N_19368,N_19928);
or UO_1303 (O_1303,N_19673,N_19893);
or UO_1304 (O_1304,N_19196,N_19096);
nand UO_1305 (O_1305,N_19008,N_19671);
or UO_1306 (O_1306,N_19185,N_19783);
nor UO_1307 (O_1307,N_19555,N_19610);
or UO_1308 (O_1308,N_19814,N_19023);
xor UO_1309 (O_1309,N_19988,N_19428);
xor UO_1310 (O_1310,N_19078,N_19641);
nor UO_1311 (O_1311,N_19946,N_19486);
or UO_1312 (O_1312,N_19893,N_19954);
or UO_1313 (O_1313,N_19656,N_19171);
nor UO_1314 (O_1314,N_19908,N_19833);
xor UO_1315 (O_1315,N_19578,N_19656);
xnor UO_1316 (O_1316,N_19817,N_19920);
and UO_1317 (O_1317,N_19571,N_19909);
or UO_1318 (O_1318,N_19551,N_19364);
and UO_1319 (O_1319,N_19475,N_19632);
nor UO_1320 (O_1320,N_19215,N_19106);
nor UO_1321 (O_1321,N_19484,N_19836);
nand UO_1322 (O_1322,N_19164,N_19714);
nand UO_1323 (O_1323,N_19837,N_19535);
xnor UO_1324 (O_1324,N_19303,N_19808);
xor UO_1325 (O_1325,N_19630,N_19527);
and UO_1326 (O_1326,N_19673,N_19258);
and UO_1327 (O_1327,N_19492,N_19011);
nor UO_1328 (O_1328,N_19692,N_19118);
nor UO_1329 (O_1329,N_19663,N_19343);
nand UO_1330 (O_1330,N_19888,N_19066);
or UO_1331 (O_1331,N_19033,N_19360);
nor UO_1332 (O_1332,N_19268,N_19563);
and UO_1333 (O_1333,N_19738,N_19410);
and UO_1334 (O_1334,N_19562,N_19611);
and UO_1335 (O_1335,N_19142,N_19571);
and UO_1336 (O_1336,N_19972,N_19917);
nand UO_1337 (O_1337,N_19578,N_19071);
nand UO_1338 (O_1338,N_19325,N_19383);
nor UO_1339 (O_1339,N_19510,N_19915);
and UO_1340 (O_1340,N_19367,N_19848);
nor UO_1341 (O_1341,N_19835,N_19318);
xnor UO_1342 (O_1342,N_19902,N_19054);
and UO_1343 (O_1343,N_19053,N_19824);
nand UO_1344 (O_1344,N_19937,N_19910);
or UO_1345 (O_1345,N_19396,N_19456);
nor UO_1346 (O_1346,N_19704,N_19221);
and UO_1347 (O_1347,N_19001,N_19253);
nor UO_1348 (O_1348,N_19937,N_19334);
or UO_1349 (O_1349,N_19981,N_19383);
nand UO_1350 (O_1350,N_19602,N_19673);
or UO_1351 (O_1351,N_19918,N_19057);
nor UO_1352 (O_1352,N_19322,N_19451);
nor UO_1353 (O_1353,N_19249,N_19630);
xor UO_1354 (O_1354,N_19813,N_19651);
nor UO_1355 (O_1355,N_19236,N_19968);
xor UO_1356 (O_1356,N_19833,N_19858);
xnor UO_1357 (O_1357,N_19238,N_19250);
xnor UO_1358 (O_1358,N_19420,N_19772);
and UO_1359 (O_1359,N_19572,N_19747);
nor UO_1360 (O_1360,N_19948,N_19475);
nor UO_1361 (O_1361,N_19373,N_19801);
or UO_1362 (O_1362,N_19842,N_19527);
or UO_1363 (O_1363,N_19635,N_19795);
nand UO_1364 (O_1364,N_19422,N_19225);
nand UO_1365 (O_1365,N_19981,N_19453);
and UO_1366 (O_1366,N_19908,N_19052);
xor UO_1367 (O_1367,N_19986,N_19995);
nor UO_1368 (O_1368,N_19361,N_19400);
nor UO_1369 (O_1369,N_19956,N_19172);
nand UO_1370 (O_1370,N_19982,N_19850);
and UO_1371 (O_1371,N_19292,N_19728);
or UO_1372 (O_1372,N_19241,N_19102);
and UO_1373 (O_1373,N_19046,N_19540);
nor UO_1374 (O_1374,N_19193,N_19887);
nand UO_1375 (O_1375,N_19766,N_19188);
or UO_1376 (O_1376,N_19563,N_19764);
xor UO_1377 (O_1377,N_19841,N_19299);
and UO_1378 (O_1378,N_19226,N_19037);
or UO_1379 (O_1379,N_19257,N_19104);
xor UO_1380 (O_1380,N_19454,N_19978);
or UO_1381 (O_1381,N_19705,N_19798);
xor UO_1382 (O_1382,N_19469,N_19384);
nor UO_1383 (O_1383,N_19114,N_19540);
and UO_1384 (O_1384,N_19876,N_19997);
nor UO_1385 (O_1385,N_19665,N_19248);
or UO_1386 (O_1386,N_19106,N_19248);
nand UO_1387 (O_1387,N_19142,N_19327);
nor UO_1388 (O_1388,N_19626,N_19535);
and UO_1389 (O_1389,N_19250,N_19470);
nand UO_1390 (O_1390,N_19771,N_19227);
nor UO_1391 (O_1391,N_19010,N_19653);
or UO_1392 (O_1392,N_19130,N_19113);
nor UO_1393 (O_1393,N_19354,N_19984);
xnor UO_1394 (O_1394,N_19150,N_19558);
xnor UO_1395 (O_1395,N_19110,N_19995);
and UO_1396 (O_1396,N_19657,N_19833);
nand UO_1397 (O_1397,N_19180,N_19774);
nand UO_1398 (O_1398,N_19879,N_19334);
and UO_1399 (O_1399,N_19068,N_19537);
and UO_1400 (O_1400,N_19428,N_19327);
or UO_1401 (O_1401,N_19229,N_19165);
or UO_1402 (O_1402,N_19889,N_19656);
and UO_1403 (O_1403,N_19753,N_19390);
nor UO_1404 (O_1404,N_19081,N_19698);
or UO_1405 (O_1405,N_19633,N_19921);
nor UO_1406 (O_1406,N_19965,N_19382);
xnor UO_1407 (O_1407,N_19124,N_19283);
or UO_1408 (O_1408,N_19803,N_19837);
xor UO_1409 (O_1409,N_19510,N_19542);
xor UO_1410 (O_1410,N_19563,N_19929);
nor UO_1411 (O_1411,N_19873,N_19822);
or UO_1412 (O_1412,N_19467,N_19448);
xor UO_1413 (O_1413,N_19311,N_19159);
nor UO_1414 (O_1414,N_19402,N_19456);
nor UO_1415 (O_1415,N_19336,N_19796);
nor UO_1416 (O_1416,N_19105,N_19324);
nand UO_1417 (O_1417,N_19699,N_19381);
or UO_1418 (O_1418,N_19234,N_19466);
and UO_1419 (O_1419,N_19289,N_19070);
or UO_1420 (O_1420,N_19201,N_19717);
xor UO_1421 (O_1421,N_19183,N_19565);
xnor UO_1422 (O_1422,N_19493,N_19352);
nor UO_1423 (O_1423,N_19705,N_19847);
nand UO_1424 (O_1424,N_19007,N_19838);
nand UO_1425 (O_1425,N_19484,N_19029);
and UO_1426 (O_1426,N_19696,N_19713);
nand UO_1427 (O_1427,N_19457,N_19534);
or UO_1428 (O_1428,N_19363,N_19234);
xnor UO_1429 (O_1429,N_19703,N_19097);
xnor UO_1430 (O_1430,N_19451,N_19839);
nor UO_1431 (O_1431,N_19615,N_19163);
and UO_1432 (O_1432,N_19352,N_19596);
or UO_1433 (O_1433,N_19249,N_19288);
xor UO_1434 (O_1434,N_19011,N_19699);
xor UO_1435 (O_1435,N_19750,N_19855);
and UO_1436 (O_1436,N_19992,N_19302);
nor UO_1437 (O_1437,N_19810,N_19755);
and UO_1438 (O_1438,N_19699,N_19646);
xor UO_1439 (O_1439,N_19893,N_19603);
xnor UO_1440 (O_1440,N_19521,N_19300);
and UO_1441 (O_1441,N_19771,N_19732);
nor UO_1442 (O_1442,N_19229,N_19372);
or UO_1443 (O_1443,N_19101,N_19385);
and UO_1444 (O_1444,N_19569,N_19305);
xor UO_1445 (O_1445,N_19801,N_19938);
nor UO_1446 (O_1446,N_19198,N_19457);
nor UO_1447 (O_1447,N_19680,N_19907);
and UO_1448 (O_1448,N_19745,N_19267);
or UO_1449 (O_1449,N_19868,N_19241);
nand UO_1450 (O_1450,N_19811,N_19070);
xor UO_1451 (O_1451,N_19757,N_19741);
or UO_1452 (O_1452,N_19838,N_19576);
and UO_1453 (O_1453,N_19532,N_19163);
and UO_1454 (O_1454,N_19966,N_19967);
nor UO_1455 (O_1455,N_19210,N_19183);
xnor UO_1456 (O_1456,N_19473,N_19903);
and UO_1457 (O_1457,N_19673,N_19263);
nand UO_1458 (O_1458,N_19752,N_19754);
or UO_1459 (O_1459,N_19601,N_19109);
nor UO_1460 (O_1460,N_19444,N_19864);
or UO_1461 (O_1461,N_19372,N_19140);
and UO_1462 (O_1462,N_19062,N_19512);
nand UO_1463 (O_1463,N_19966,N_19113);
nor UO_1464 (O_1464,N_19171,N_19352);
or UO_1465 (O_1465,N_19092,N_19500);
or UO_1466 (O_1466,N_19811,N_19010);
or UO_1467 (O_1467,N_19337,N_19212);
nand UO_1468 (O_1468,N_19401,N_19518);
or UO_1469 (O_1469,N_19581,N_19342);
nand UO_1470 (O_1470,N_19999,N_19638);
and UO_1471 (O_1471,N_19268,N_19428);
or UO_1472 (O_1472,N_19218,N_19261);
nand UO_1473 (O_1473,N_19746,N_19440);
and UO_1474 (O_1474,N_19434,N_19220);
nand UO_1475 (O_1475,N_19069,N_19556);
nand UO_1476 (O_1476,N_19259,N_19829);
or UO_1477 (O_1477,N_19611,N_19862);
nor UO_1478 (O_1478,N_19207,N_19183);
nand UO_1479 (O_1479,N_19426,N_19876);
xor UO_1480 (O_1480,N_19967,N_19302);
and UO_1481 (O_1481,N_19776,N_19253);
xor UO_1482 (O_1482,N_19771,N_19345);
or UO_1483 (O_1483,N_19991,N_19073);
and UO_1484 (O_1484,N_19631,N_19540);
nand UO_1485 (O_1485,N_19344,N_19680);
nor UO_1486 (O_1486,N_19415,N_19021);
xnor UO_1487 (O_1487,N_19362,N_19059);
or UO_1488 (O_1488,N_19881,N_19589);
nor UO_1489 (O_1489,N_19990,N_19740);
and UO_1490 (O_1490,N_19626,N_19152);
nor UO_1491 (O_1491,N_19950,N_19891);
xor UO_1492 (O_1492,N_19478,N_19769);
or UO_1493 (O_1493,N_19770,N_19637);
xnor UO_1494 (O_1494,N_19967,N_19543);
nor UO_1495 (O_1495,N_19195,N_19581);
or UO_1496 (O_1496,N_19933,N_19174);
and UO_1497 (O_1497,N_19749,N_19721);
nor UO_1498 (O_1498,N_19834,N_19400);
xor UO_1499 (O_1499,N_19112,N_19600);
nand UO_1500 (O_1500,N_19977,N_19192);
nor UO_1501 (O_1501,N_19199,N_19937);
nor UO_1502 (O_1502,N_19880,N_19747);
and UO_1503 (O_1503,N_19065,N_19808);
or UO_1504 (O_1504,N_19683,N_19465);
nand UO_1505 (O_1505,N_19887,N_19101);
xnor UO_1506 (O_1506,N_19272,N_19303);
and UO_1507 (O_1507,N_19053,N_19825);
nand UO_1508 (O_1508,N_19650,N_19461);
nor UO_1509 (O_1509,N_19270,N_19914);
xnor UO_1510 (O_1510,N_19851,N_19021);
xor UO_1511 (O_1511,N_19356,N_19245);
and UO_1512 (O_1512,N_19891,N_19993);
or UO_1513 (O_1513,N_19424,N_19003);
or UO_1514 (O_1514,N_19307,N_19413);
xnor UO_1515 (O_1515,N_19786,N_19839);
and UO_1516 (O_1516,N_19954,N_19867);
nand UO_1517 (O_1517,N_19636,N_19850);
xnor UO_1518 (O_1518,N_19052,N_19195);
nand UO_1519 (O_1519,N_19331,N_19558);
and UO_1520 (O_1520,N_19308,N_19622);
xor UO_1521 (O_1521,N_19875,N_19520);
or UO_1522 (O_1522,N_19842,N_19053);
or UO_1523 (O_1523,N_19998,N_19321);
nor UO_1524 (O_1524,N_19056,N_19934);
or UO_1525 (O_1525,N_19911,N_19550);
nor UO_1526 (O_1526,N_19326,N_19454);
xor UO_1527 (O_1527,N_19735,N_19933);
or UO_1528 (O_1528,N_19230,N_19911);
or UO_1529 (O_1529,N_19281,N_19849);
nand UO_1530 (O_1530,N_19493,N_19678);
nor UO_1531 (O_1531,N_19012,N_19995);
or UO_1532 (O_1532,N_19166,N_19458);
xnor UO_1533 (O_1533,N_19419,N_19841);
and UO_1534 (O_1534,N_19116,N_19217);
and UO_1535 (O_1535,N_19640,N_19916);
nor UO_1536 (O_1536,N_19988,N_19525);
nor UO_1537 (O_1537,N_19402,N_19989);
or UO_1538 (O_1538,N_19957,N_19771);
nand UO_1539 (O_1539,N_19935,N_19624);
xnor UO_1540 (O_1540,N_19119,N_19855);
or UO_1541 (O_1541,N_19163,N_19485);
xnor UO_1542 (O_1542,N_19358,N_19162);
xnor UO_1543 (O_1543,N_19199,N_19394);
and UO_1544 (O_1544,N_19343,N_19839);
nor UO_1545 (O_1545,N_19842,N_19909);
or UO_1546 (O_1546,N_19633,N_19968);
nor UO_1547 (O_1547,N_19431,N_19023);
or UO_1548 (O_1548,N_19284,N_19154);
nand UO_1549 (O_1549,N_19954,N_19308);
nor UO_1550 (O_1550,N_19417,N_19841);
nand UO_1551 (O_1551,N_19788,N_19577);
or UO_1552 (O_1552,N_19836,N_19739);
and UO_1553 (O_1553,N_19214,N_19469);
xnor UO_1554 (O_1554,N_19970,N_19522);
xor UO_1555 (O_1555,N_19481,N_19245);
nor UO_1556 (O_1556,N_19342,N_19578);
or UO_1557 (O_1557,N_19234,N_19573);
nor UO_1558 (O_1558,N_19608,N_19577);
and UO_1559 (O_1559,N_19990,N_19437);
and UO_1560 (O_1560,N_19044,N_19255);
and UO_1561 (O_1561,N_19020,N_19597);
and UO_1562 (O_1562,N_19327,N_19838);
and UO_1563 (O_1563,N_19162,N_19506);
nand UO_1564 (O_1564,N_19653,N_19935);
or UO_1565 (O_1565,N_19832,N_19138);
nor UO_1566 (O_1566,N_19624,N_19437);
or UO_1567 (O_1567,N_19231,N_19594);
and UO_1568 (O_1568,N_19431,N_19681);
nand UO_1569 (O_1569,N_19051,N_19495);
xor UO_1570 (O_1570,N_19052,N_19796);
and UO_1571 (O_1571,N_19086,N_19038);
or UO_1572 (O_1572,N_19995,N_19164);
xnor UO_1573 (O_1573,N_19050,N_19215);
nand UO_1574 (O_1574,N_19837,N_19152);
nor UO_1575 (O_1575,N_19179,N_19896);
or UO_1576 (O_1576,N_19075,N_19861);
and UO_1577 (O_1577,N_19958,N_19813);
or UO_1578 (O_1578,N_19173,N_19610);
xnor UO_1579 (O_1579,N_19581,N_19164);
xor UO_1580 (O_1580,N_19073,N_19735);
nor UO_1581 (O_1581,N_19899,N_19134);
nand UO_1582 (O_1582,N_19108,N_19244);
nor UO_1583 (O_1583,N_19869,N_19333);
nand UO_1584 (O_1584,N_19758,N_19843);
and UO_1585 (O_1585,N_19505,N_19748);
or UO_1586 (O_1586,N_19759,N_19421);
nand UO_1587 (O_1587,N_19811,N_19549);
and UO_1588 (O_1588,N_19430,N_19163);
or UO_1589 (O_1589,N_19241,N_19563);
and UO_1590 (O_1590,N_19416,N_19772);
and UO_1591 (O_1591,N_19570,N_19183);
nor UO_1592 (O_1592,N_19590,N_19927);
nor UO_1593 (O_1593,N_19006,N_19202);
and UO_1594 (O_1594,N_19695,N_19115);
or UO_1595 (O_1595,N_19381,N_19128);
xnor UO_1596 (O_1596,N_19532,N_19075);
nand UO_1597 (O_1597,N_19865,N_19593);
or UO_1598 (O_1598,N_19357,N_19290);
or UO_1599 (O_1599,N_19959,N_19438);
nand UO_1600 (O_1600,N_19274,N_19661);
xnor UO_1601 (O_1601,N_19600,N_19291);
and UO_1602 (O_1602,N_19428,N_19461);
or UO_1603 (O_1603,N_19525,N_19140);
or UO_1604 (O_1604,N_19314,N_19921);
nor UO_1605 (O_1605,N_19344,N_19949);
nor UO_1606 (O_1606,N_19598,N_19370);
nand UO_1607 (O_1607,N_19409,N_19768);
and UO_1608 (O_1608,N_19508,N_19538);
xnor UO_1609 (O_1609,N_19163,N_19497);
or UO_1610 (O_1610,N_19912,N_19434);
nand UO_1611 (O_1611,N_19002,N_19754);
nor UO_1612 (O_1612,N_19506,N_19531);
nor UO_1613 (O_1613,N_19322,N_19234);
nand UO_1614 (O_1614,N_19659,N_19773);
nand UO_1615 (O_1615,N_19757,N_19870);
nor UO_1616 (O_1616,N_19212,N_19548);
or UO_1617 (O_1617,N_19555,N_19179);
xnor UO_1618 (O_1618,N_19528,N_19415);
nand UO_1619 (O_1619,N_19760,N_19264);
and UO_1620 (O_1620,N_19608,N_19858);
nand UO_1621 (O_1621,N_19713,N_19662);
and UO_1622 (O_1622,N_19890,N_19246);
and UO_1623 (O_1623,N_19332,N_19411);
xor UO_1624 (O_1624,N_19236,N_19762);
nor UO_1625 (O_1625,N_19242,N_19053);
nand UO_1626 (O_1626,N_19983,N_19940);
xor UO_1627 (O_1627,N_19576,N_19890);
or UO_1628 (O_1628,N_19455,N_19573);
nor UO_1629 (O_1629,N_19040,N_19437);
nor UO_1630 (O_1630,N_19036,N_19193);
xnor UO_1631 (O_1631,N_19433,N_19375);
or UO_1632 (O_1632,N_19177,N_19321);
xor UO_1633 (O_1633,N_19616,N_19181);
nand UO_1634 (O_1634,N_19205,N_19440);
xor UO_1635 (O_1635,N_19993,N_19536);
xnor UO_1636 (O_1636,N_19197,N_19316);
xnor UO_1637 (O_1637,N_19156,N_19755);
and UO_1638 (O_1638,N_19405,N_19345);
and UO_1639 (O_1639,N_19388,N_19625);
nor UO_1640 (O_1640,N_19216,N_19151);
xor UO_1641 (O_1641,N_19329,N_19339);
nor UO_1642 (O_1642,N_19576,N_19012);
nand UO_1643 (O_1643,N_19460,N_19846);
nand UO_1644 (O_1644,N_19848,N_19172);
nor UO_1645 (O_1645,N_19017,N_19460);
xor UO_1646 (O_1646,N_19429,N_19255);
nor UO_1647 (O_1647,N_19596,N_19532);
xor UO_1648 (O_1648,N_19496,N_19129);
and UO_1649 (O_1649,N_19092,N_19572);
nor UO_1650 (O_1650,N_19966,N_19297);
and UO_1651 (O_1651,N_19983,N_19903);
or UO_1652 (O_1652,N_19238,N_19265);
or UO_1653 (O_1653,N_19790,N_19771);
or UO_1654 (O_1654,N_19162,N_19056);
nor UO_1655 (O_1655,N_19389,N_19665);
nand UO_1656 (O_1656,N_19459,N_19087);
nor UO_1657 (O_1657,N_19109,N_19268);
xnor UO_1658 (O_1658,N_19985,N_19606);
nor UO_1659 (O_1659,N_19825,N_19522);
nand UO_1660 (O_1660,N_19602,N_19963);
nor UO_1661 (O_1661,N_19586,N_19301);
xor UO_1662 (O_1662,N_19287,N_19320);
nand UO_1663 (O_1663,N_19595,N_19085);
nor UO_1664 (O_1664,N_19305,N_19637);
xnor UO_1665 (O_1665,N_19781,N_19981);
nand UO_1666 (O_1666,N_19001,N_19333);
nand UO_1667 (O_1667,N_19195,N_19569);
or UO_1668 (O_1668,N_19965,N_19416);
nand UO_1669 (O_1669,N_19646,N_19778);
xnor UO_1670 (O_1670,N_19456,N_19539);
nor UO_1671 (O_1671,N_19520,N_19164);
nor UO_1672 (O_1672,N_19566,N_19043);
and UO_1673 (O_1673,N_19230,N_19146);
or UO_1674 (O_1674,N_19196,N_19584);
or UO_1675 (O_1675,N_19824,N_19357);
or UO_1676 (O_1676,N_19566,N_19429);
nand UO_1677 (O_1677,N_19662,N_19614);
and UO_1678 (O_1678,N_19802,N_19040);
nand UO_1679 (O_1679,N_19646,N_19342);
nand UO_1680 (O_1680,N_19260,N_19059);
and UO_1681 (O_1681,N_19904,N_19771);
xor UO_1682 (O_1682,N_19885,N_19010);
and UO_1683 (O_1683,N_19364,N_19969);
or UO_1684 (O_1684,N_19116,N_19754);
nor UO_1685 (O_1685,N_19964,N_19110);
and UO_1686 (O_1686,N_19973,N_19031);
or UO_1687 (O_1687,N_19421,N_19398);
nor UO_1688 (O_1688,N_19125,N_19086);
xnor UO_1689 (O_1689,N_19144,N_19762);
nand UO_1690 (O_1690,N_19487,N_19271);
or UO_1691 (O_1691,N_19650,N_19670);
xor UO_1692 (O_1692,N_19382,N_19508);
and UO_1693 (O_1693,N_19885,N_19546);
nor UO_1694 (O_1694,N_19726,N_19558);
or UO_1695 (O_1695,N_19769,N_19839);
nand UO_1696 (O_1696,N_19980,N_19350);
nor UO_1697 (O_1697,N_19341,N_19946);
or UO_1698 (O_1698,N_19400,N_19552);
and UO_1699 (O_1699,N_19586,N_19878);
nand UO_1700 (O_1700,N_19688,N_19771);
nand UO_1701 (O_1701,N_19105,N_19074);
xnor UO_1702 (O_1702,N_19095,N_19707);
and UO_1703 (O_1703,N_19344,N_19186);
nand UO_1704 (O_1704,N_19098,N_19676);
and UO_1705 (O_1705,N_19003,N_19729);
or UO_1706 (O_1706,N_19782,N_19253);
and UO_1707 (O_1707,N_19053,N_19580);
xor UO_1708 (O_1708,N_19485,N_19962);
xor UO_1709 (O_1709,N_19210,N_19360);
xor UO_1710 (O_1710,N_19412,N_19175);
nand UO_1711 (O_1711,N_19903,N_19701);
nand UO_1712 (O_1712,N_19714,N_19877);
nor UO_1713 (O_1713,N_19411,N_19376);
nor UO_1714 (O_1714,N_19221,N_19875);
nand UO_1715 (O_1715,N_19482,N_19776);
and UO_1716 (O_1716,N_19461,N_19528);
nor UO_1717 (O_1717,N_19519,N_19863);
or UO_1718 (O_1718,N_19087,N_19238);
nor UO_1719 (O_1719,N_19447,N_19699);
xor UO_1720 (O_1720,N_19763,N_19215);
and UO_1721 (O_1721,N_19701,N_19519);
nand UO_1722 (O_1722,N_19941,N_19882);
and UO_1723 (O_1723,N_19097,N_19189);
nor UO_1724 (O_1724,N_19427,N_19865);
and UO_1725 (O_1725,N_19969,N_19636);
nand UO_1726 (O_1726,N_19688,N_19872);
nor UO_1727 (O_1727,N_19518,N_19629);
nor UO_1728 (O_1728,N_19154,N_19780);
and UO_1729 (O_1729,N_19386,N_19078);
or UO_1730 (O_1730,N_19427,N_19548);
nor UO_1731 (O_1731,N_19791,N_19239);
and UO_1732 (O_1732,N_19471,N_19113);
and UO_1733 (O_1733,N_19330,N_19696);
nor UO_1734 (O_1734,N_19085,N_19243);
and UO_1735 (O_1735,N_19797,N_19027);
nor UO_1736 (O_1736,N_19430,N_19992);
nand UO_1737 (O_1737,N_19151,N_19664);
and UO_1738 (O_1738,N_19177,N_19200);
and UO_1739 (O_1739,N_19142,N_19286);
nor UO_1740 (O_1740,N_19907,N_19087);
or UO_1741 (O_1741,N_19528,N_19843);
xnor UO_1742 (O_1742,N_19002,N_19054);
nor UO_1743 (O_1743,N_19404,N_19363);
or UO_1744 (O_1744,N_19161,N_19470);
or UO_1745 (O_1745,N_19080,N_19772);
nand UO_1746 (O_1746,N_19196,N_19408);
or UO_1747 (O_1747,N_19740,N_19014);
nand UO_1748 (O_1748,N_19576,N_19254);
nand UO_1749 (O_1749,N_19472,N_19711);
or UO_1750 (O_1750,N_19290,N_19271);
nand UO_1751 (O_1751,N_19682,N_19006);
xnor UO_1752 (O_1752,N_19683,N_19561);
nor UO_1753 (O_1753,N_19726,N_19732);
nor UO_1754 (O_1754,N_19275,N_19725);
nand UO_1755 (O_1755,N_19346,N_19247);
nand UO_1756 (O_1756,N_19616,N_19528);
nor UO_1757 (O_1757,N_19678,N_19993);
xnor UO_1758 (O_1758,N_19207,N_19899);
or UO_1759 (O_1759,N_19774,N_19711);
and UO_1760 (O_1760,N_19808,N_19304);
or UO_1761 (O_1761,N_19175,N_19304);
nor UO_1762 (O_1762,N_19570,N_19313);
xnor UO_1763 (O_1763,N_19812,N_19031);
and UO_1764 (O_1764,N_19607,N_19286);
nor UO_1765 (O_1765,N_19113,N_19729);
nor UO_1766 (O_1766,N_19930,N_19784);
and UO_1767 (O_1767,N_19298,N_19668);
nor UO_1768 (O_1768,N_19302,N_19424);
nand UO_1769 (O_1769,N_19544,N_19170);
and UO_1770 (O_1770,N_19429,N_19595);
or UO_1771 (O_1771,N_19974,N_19175);
xor UO_1772 (O_1772,N_19051,N_19855);
nand UO_1773 (O_1773,N_19891,N_19474);
nand UO_1774 (O_1774,N_19488,N_19402);
or UO_1775 (O_1775,N_19793,N_19661);
xor UO_1776 (O_1776,N_19090,N_19233);
and UO_1777 (O_1777,N_19959,N_19444);
or UO_1778 (O_1778,N_19181,N_19084);
xor UO_1779 (O_1779,N_19604,N_19315);
nand UO_1780 (O_1780,N_19138,N_19583);
xnor UO_1781 (O_1781,N_19096,N_19801);
xnor UO_1782 (O_1782,N_19884,N_19252);
nand UO_1783 (O_1783,N_19212,N_19470);
nor UO_1784 (O_1784,N_19753,N_19250);
or UO_1785 (O_1785,N_19012,N_19723);
or UO_1786 (O_1786,N_19786,N_19248);
xor UO_1787 (O_1787,N_19207,N_19060);
nor UO_1788 (O_1788,N_19240,N_19821);
and UO_1789 (O_1789,N_19796,N_19048);
nor UO_1790 (O_1790,N_19308,N_19370);
xor UO_1791 (O_1791,N_19473,N_19053);
and UO_1792 (O_1792,N_19033,N_19436);
nand UO_1793 (O_1793,N_19919,N_19782);
and UO_1794 (O_1794,N_19005,N_19828);
xnor UO_1795 (O_1795,N_19691,N_19394);
nand UO_1796 (O_1796,N_19499,N_19179);
or UO_1797 (O_1797,N_19894,N_19828);
and UO_1798 (O_1798,N_19867,N_19173);
or UO_1799 (O_1799,N_19184,N_19468);
or UO_1800 (O_1800,N_19755,N_19571);
nor UO_1801 (O_1801,N_19739,N_19043);
nand UO_1802 (O_1802,N_19879,N_19305);
nor UO_1803 (O_1803,N_19709,N_19228);
nand UO_1804 (O_1804,N_19844,N_19399);
and UO_1805 (O_1805,N_19967,N_19056);
xor UO_1806 (O_1806,N_19834,N_19983);
nand UO_1807 (O_1807,N_19415,N_19731);
and UO_1808 (O_1808,N_19585,N_19958);
nor UO_1809 (O_1809,N_19159,N_19687);
xor UO_1810 (O_1810,N_19182,N_19151);
and UO_1811 (O_1811,N_19809,N_19567);
xnor UO_1812 (O_1812,N_19529,N_19768);
xor UO_1813 (O_1813,N_19747,N_19766);
or UO_1814 (O_1814,N_19871,N_19578);
nand UO_1815 (O_1815,N_19144,N_19406);
nand UO_1816 (O_1816,N_19009,N_19845);
nand UO_1817 (O_1817,N_19816,N_19102);
or UO_1818 (O_1818,N_19355,N_19509);
or UO_1819 (O_1819,N_19095,N_19469);
or UO_1820 (O_1820,N_19705,N_19593);
or UO_1821 (O_1821,N_19749,N_19707);
nand UO_1822 (O_1822,N_19947,N_19423);
or UO_1823 (O_1823,N_19594,N_19612);
and UO_1824 (O_1824,N_19633,N_19037);
nand UO_1825 (O_1825,N_19064,N_19885);
nor UO_1826 (O_1826,N_19667,N_19402);
and UO_1827 (O_1827,N_19293,N_19176);
and UO_1828 (O_1828,N_19315,N_19919);
and UO_1829 (O_1829,N_19889,N_19308);
xor UO_1830 (O_1830,N_19740,N_19540);
nand UO_1831 (O_1831,N_19710,N_19019);
or UO_1832 (O_1832,N_19191,N_19743);
nor UO_1833 (O_1833,N_19748,N_19550);
nor UO_1834 (O_1834,N_19214,N_19920);
xnor UO_1835 (O_1835,N_19446,N_19570);
xnor UO_1836 (O_1836,N_19925,N_19951);
xor UO_1837 (O_1837,N_19526,N_19365);
and UO_1838 (O_1838,N_19461,N_19129);
nor UO_1839 (O_1839,N_19597,N_19129);
and UO_1840 (O_1840,N_19310,N_19454);
xor UO_1841 (O_1841,N_19104,N_19665);
and UO_1842 (O_1842,N_19723,N_19023);
xnor UO_1843 (O_1843,N_19072,N_19760);
or UO_1844 (O_1844,N_19546,N_19339);
and UO_1845 (O_1845,N_19151,N_19418);
nand UO_1846 (O_1846,N_19184,N_19615);
nor UO_1847 (O_1847,N_19433,N_19681);
nand UO_1848 (O_1848,N_19583,N_19373);
nor UO_1849 (O_1849,N_19316,N_19334);
nand UO_1850 (O_1850,N_19469,N_19926);
nor UO_1851 (O_1851,N_19533,N_19111);
nand UO_1852 (O_1852,N_19067,N_19823);
or UO_1853 (O_1853,N_19031,N_19524);
and UO_1854 (O_1854,N_19954,N_19734);
and UO_1855 (O_1855,N_19628,N_19701);
nor UO_1856 (O_1856,N_19555,N_19938);
nand UO_1857 (O_1857,N_19908,N_19955);
nor UO_1858 (O_1858,N_19299,N_19882);
and UO_1859 (O_1859,N_19207,N_19007);
and UO_1860 (O_1860,N_19762,N_19783);
xnor UO_1861 (O_1861,N_19761,N_19859);
or UO_1862 (O_1862,N_19647,N_19983);
xnor UO_1863 (O_1863,N_19335,N_19114);
and UO_1864 (O_1864,N_19946,N_19304);
xor UO_1865 (O_1865,N_19123,N_19616);
or UO_1866 (O_1866,N_19660,N_19852);
nand UO_1867 (O_1867,N_19187,N_19337);
xor UO_1868 (O_1868,N_19059,N_19110);
nor UO_1869 (O_1869,N_19567,N_19387);
and UO_1870 (O_1870,N_19833,N_19853);
xor UO_1871 (O_1871,N_19234,N_19257);
nor UO_1872 (O_1872,N_19879,N_19934);
and UO_1873 (O_1873,N_19992,N_19721);
or UO_1874 (O_1874,N_19934,N_19891);
xor UO_1875 (O_1875,N_19004,N_19211);
or UO_1876 (O_1876,N_19652,N_19171);
and UO_1877 (O_1877,N_19362,N_19738);
or UO_1878 (O_1878,N_19832,N_19323);
or UO_1879 (O_1879,N_19100,N_19076);
xor UO_1880 (O_1880,N_19354,N_19238);
nor UO_1881 (O_1881,N_19716,N_19960);
or UO_1882 (O_1882,N_19241,N_19652);
and UO_1883 (O_1883,N_19390,N_19638);
and UO_1884 (O_1884,N_19627,N_19899);
nor UO_1885 (O_1885,N_19508,N_19681);
nor UO_1886 (O_1886,N_19396,N_19439);
nand UO_1887 (O_1887,N_19210,N_19642);
nor UO_1888 (O_1888,N_19069,N_19384);
nand UO_1889 (O_1889,N_19796,N_19058);
and UO_1890 (O_1890,N_19972,N_19388);
nor UO_1891 (O_1891,N_19978,N_19237);
or UO_1892 (O_1892,N_19881,N_19093);
and UO_1893 (O_1893,N_19871,N_19038);
and UO_1894 (O_1894,N_19318,N_19726);
nor UO_1895 (O_1895,N_19799,N_19674);
nand UO_1896 (O_1896,N_19776,N_19739);
xor UO_1897 (O_1897,N_19058,N_19630);
xor UO_1898 (O_1898,N_19575,N_19553);
and UO_1899 (O_1899,N_19664,N_19093);
nor UO_1900 (O_1900,N_19925,N_19439);
nor UO_1901 (O_1901,N_19700,N_19696);
nor UO_1902 (O_1902,N_19789,N_19000);
nand UO_1903 (O_1903,N_19050,N_19018);
nand UO_1904 (O_1904,N_19937,N_19764);
xor UO_1905 (O_1905,N_19460,N_19330);
or UO_1906 (O_1906,N_19590,N_19383);
xnor UO_1907 (O_1907,N_19864,N_19267);
or UO_1908 (O_1908,N_19592,N_19548);
and UO_1909 (O_1909,N_19746,N_19206);
or UO_1910 (O_1910,N_19281,N_19479);
and UO_1911 (O_1911,N_19253,N_19007);
and UO_1912 (O_1912,N_19314,N_19128);
and UO_1913 (O_1913,N_19310,N_19910);
or UO_1914 (O_1914,N_19562,N_19482);
or UO_1915 (O_1915,N_19039,N_19004);
nand UO_1916 (O_1916,N_19617,N_19414);
or UO_1917 (O_1917,N_19125,N_19919);
and UO_1918 (O_1918,N_19411,N_19791);
and UO_1919 (O_1919,N_19828,N_19530);
nor UO_1920 (O_1920,N_19281,N_19246);
nor UO_1921 (O_1921,N_19091,N_19454);
nor UO_1922 (O_1922,N_19672,N_19862);
xor UO_1923 (O_1923,N_19098,N_19565);
or UO_1924 (O_1924,N_19964,N_19548);
xor UO_1925 (O_1925,N_19223,N_19523);
nor UO_1926 (O_1926,N_19413,N_19314);
or UO_1927 (O_1927,N_19430,N_19461);
or UO_1928 (O_1928,N_19432,N_19743);
nor UO_1929 (O_1929,N_19633,N_19795);
xor UO_1930 (O_1930,N_19105,N_19659);
nand UO_1931 (O_1931,N_19960,N_19045);
or UO_1932 (O_1932,N_19368,N_19594);
xnor UO_1933 (O_1933,N_19119,N_19808);
or UO_1934 (O_1934,N_19724,N_19805);
or UO_1935 (O_1935,N_19676,N_19968);
or UO_1936 (O_1936,N_19317,N_19843);
or UO_1937 (O_1937,N_19735,N_19291);
nand UO_1938 (O_1938,N_19587,N_19471);
and UO_1939 (O_1939,N_19355,N_19787);
nand UO_1940 (O_1940,N_19402,N_19151);
xor UO_1941 (O_1941,N_19525,N_19560);
xor UO_1942 (O_1942,N_19660,N_19489);
xnor UO_1943 (O_1943,N_19699,N_19082);
or UO_1944 (O_1944,N_19245,N_19175);
and UO_1945 (O_1945,N_19102,N_19886);
and UO_1946 (O_1946,N_19908,N_19244);
nand UO_1947 (O_1947,N_19351,N_19189);
or UO_1948 (O_1948,N_19942,N_19726);
xnor UO_1949 (O_1949,N_19997,N_19867);
nand UO_1950 (O_1950,N_19691,N_19731);
xnor UO_1951 (O_1951,N_19265,N_19500);
or UO_1952 (O_1952,N_19500,N_19597);
xor UO_1953 (O_1953,N_19467,N_19002);
nand UO_1954 (O_1954,N_19773,N_19646);
or UO_1955 (O_1955,N_19329,N_19122);
or UO_1956 (O_1956,N_19624,N_19909);
or UO_1957 (O_1957,N_19108,N_19594);
and UO_1958 (O_1958,N_19172,N_19804);
and UO_1959 (O_1959,N_19416,N_19727);
nand UO_1960 (O_1960,N_19471,N_19114);
xnor UO_1961 (O_1961,N_19732,N_19585);
and UO_1962 (O_1962,N_19683,N_19806);
nand UO_1963 (O_1963,N_19040,N_19063);
nor UO_1964 (O_1964,N_19620,N_19910);
or UO_1965 (O_1965,N_19469,N_19603);
nor UO_1966 (O_1966,N_19756,N_19959);
nor UO_1967 (O_1967,N_19336,N_19260);
nor UO_1968 (O_1968,N_19594,N_19391);
nor UO_1969 (O_1969,N_19355,N_19917);
or UO_1970 (O_1970,N_19545,N_19772);
nand UO_1971 (O_1971,N_19706,N_19270);
or UO_1972 (O_1972,N_19025,N_19860);
xor UO_1973 (O_1973,N_19506,N_19171);
xor UO_1974 (O_1974,N_19398,N_19007);
nor UO_1975 (O_1975,N_19044,N_19840);
nor UO_1976 (O_1976,N_19034,N_19740);
nor UO_1977 (O_1977,N_19069,N_19472);
nand UO_1978 (O_1978,N_19785,N_19074);
or UO_1979 (O_1979,N_19774,N_19299);
and UO_1980 (O_1980,N_19129,N_19514);
nand UO_1981 (O_1981,N_19854,N_19375);
and UO_1982 (O_1982,N_19777,N_19824);
xnor UO_1983 (O_1983,N_19449,N_19055);
and UO_1984 (O_1984,N_19650,N_19794);
and UO_1985 (O_1985,N_19266,N_19138);
and UO_1986 (O_1986,N_19981,N_19279);
nor UO_1987 (O_1987,N_19514,N_19494);
or UO_1988 (O_1988,N_19909,N_19954);
nor UO_1989 (O_1989,N_19149,N_19150);
and UO_1990 (O_1990,N_19478,N_19000);
xnor UO_1991 (O_1991,N_19213,N_19957);
xor UO_1992 (O_1992,N_19466,N_19008);
nor UO_1993 (O_1993,N_19935,N_19144);
or UO_1994 (O_1994,N_19969,N_19038);
nor UO_1995 (O_1995,N_19099,N_19647);
nor UO_1996 (O_1996,N_19615,N_19663);
or UO_1997 (O_1997,N_19200,N_19169);
nor UO_1998 (O_1998,N_19784,N_19821);
xnor UO_1999 (O_1999,N_19334,N_19170);
nand UO_2000 (O_2000,N_19848,N_19769);
nand UO_2001 (O_2001,N_19692,N_19747);
and UO_2002 (O_2002,N_19212,N_19575);
xnor UO_2003 (O_2003,N_19789,N_19785);
and UO_2004 (O_2004,N_19345,N_19729);
or UO_2005 (O_2005,N_19034,N_19080);
and UO_2006 (O_2006,N_19581,N_19418);
nor UO_2007 (O_2007,N_19715,N_19149);
nor UO_2008 (O_2008,N_19296,N_19692);
or UO_2009 (O_2009,N_19078,N_19611);
nor UO_2010 (O_2010,N_19681,N_19109);
and UO_2011 (O_2011,N_19481,N_19742);
or UO_2012 (O_2012,N_19482,N_19979);
and UO_2013 (O_2013,N_19306,N_19443);
and UO_2014 (O_2014,N_19933,N_19570);
or UO_2015 (O_2015,N_19298,N_19798);
xor UO_2016 (O_2016,N_19468,N_19902);
or UO_2017 (O_2017,N_19924,N_19330);
and UO_2018 (O_2018,N_19473,N_19275);
nor UO_2019 (O_2019,N_19014,N_19004);
nor UO_2020 (O_2020,N_19805,N_19058);
or UO_2021 (O_2021,N_19497,N_19948);
nand UO_2022 (O_2022,N_19795,N_19346);
nor UO_2023 (O_2023,N_19190,N_19649);
nand UO_2024 (O_2024,N_19209,N_19419);
xnor UO_2025 (O_2025,N_19472,N_19305);
and UO_2026 (O_2026,N_19087,N_19562);
and UO_2027 (O_2027,N_19345,N_19287);
xnor UO_2028 (O_2028,N_19770,N_19507);
and UO_2029 (O_2029,N_19379,N_19895);
and UO_2030 (O_2030,N_19900,N_19759);
nor UO_2031 (O_2031,N_19985,N_19134);
or UO_2032 (O_2032,N_19555,N_19374);
or UO_2033 (O_2033,N_19098,N_19547);
xor UO_2034 (O_2034,N_19204,N_19796);
nand UO_2035 (O_2035,N_19029,N_19770);
or UO_2036 (O_2036,N_19012,N_19138);
or UO_2037 (O_2037,N_19053,N_19827);
nand UO_2038 (O_2038,N_19817,N_19507);
and UO_2039 (O_2039,N_19785,N_19226);
nor UO_2040 (O_2040,N_19376,N_19763);
or UO_2041 (O_2041,N_19822,N_19428);
nand UO_2042 (O_2042,N_19893,N_19881);
nand UO_2043 (O_2043,N_19884,N_19125);
or UO_2044 (O_2044,N_19298,N_19322);
xnor UO_2045 (O_2045,N_19056,N_19121);
and UO_2046 (O_2046,N_19083,N_19496);
and UO_2047 (O_2047,N_19790,N_19928);
nand UO_2048 (O_2048,N_19218,N_19050);
nand UO_2049 (O_2049,N_19075,N_19249);
nor UO_2050 (O_2050,N_19793,N_19393);
and UO_2051 (O_2051,N_19841,N_19205);
nand UO_2052 (O_2052,N_19726,N_19087);
xor UO_2053 (O_2053,N_19742,N_19043);
or UO_2054 (O_2054,N_19215,N_19629);
and UO_2055 (O_2055,N_19356,N_19655);
nor UO_2056 (O_2056,N_19325,N_19095);
and UO_2057 (O_2057,N_19970,N_19656);
nor UO_2058 (O_2058,N_19223,N_19550);
nor UO_2059 (O_2059,N_19761,N_19569);
or UO_2060 (O_2060,N_19173,N_19495);
nand UO_2061 (O_2061,N_19524,N_19516);
or UO_2062 (O_2062,N_19003,N_19749);
or UO_2063 (O_2063,N_19558,N_19519);
xor UO_2064 (O_2064,N_19284,N_19482);
and UO_2065 (O_2065,N_19951,N_19463);
nand UO_2066 (O_2066,N_19675,N_19007);
nor UO_2067 (O_2067,N_19079,N_19900);
or UO_2068 (O_2068,N_19457,N_19603);
nor UO_2069 (O_2069,N_19700,N_19808);
nor UO_2070 (O_2070,N_19414,N_19846);
nand UO_2071 (O_2071,N_19802,N_19382);
nand UO_2072 (O_2072,N_19167,N_19666);
nor UO_2073 (O_2073,N_19565,N_19890);
xnor UO_2074 (O_2074,N_19438,N_19919);
nand UO_2075 (O_2075,N_19405,N_19326);
and UO_2076 (O_2076,N_19274,N_19278);
and UO_2077 (O_2077,N_19096,N_19178);
nand UO_2078 (O_2078,N_19837,N_19276);
nand UO_2079 (O_2079,N_19354,N_19416);
nor UO_2080 (O_2080,N_19513,N_19670);
or UO_2081 (O_2081,N_19388,N_19736);
or UO_2082 (O_2082,N_19271,N_19425);
xor UO_2083 (O_2083,N_19761,N_19562);
xnor UO_2084 (O_2084,N_19756,N_19463);
or UO_2085 (O_2085,N_19262,N_19781);
or UO_2086 (O_2086,N_19531,N_19949);
or UO_2087 (O_2087,N_19773,N_19269);
xor UO_2088 (O_2088,N_19688,N_19847);
nand UO_2089 (O_2089,N_19638,N_19125);
nand UO_2090 (O_2090,N_19839,N_19561);
nand UO_2091 (O_2091,N_19989,N_19367);
xor UO_2092 (O_2092,N_19025,N_19631);
or UO_2093 (O_2093,N_19597,N_19611);
nor UO_2094 (O_2094,N_19068,N_19442);
nor UO_2095 (O_2095,N_19382,N_19955);
and UO_2096 (O_2096,N_19394,N_19920);
nor UO_2097 (O_2097,N_19954,N_19931);
xnor UO_2098 (O_2098,N_19256,N_19780);
and UO_2099 (O_2099,N_19438,N_19665);
or UO_2100 (O_2100,N_19989,N_19976);
or UO_2101 (O_2101,N_19295,N_19759);
nand UO_2102 (O_2102,N_19360,N_19074);
xnor UO_2103 (O_2103,N_19869,N_19256);
and UO_2104 (O_2104,N_19318,N_19495);
and UO_2105 (O_2105,N_19105,N_19217);
nand UO_2106 (O_2106,N_19297,N_19212);
nand UO_2107 (O_2107,N_19372,N_19190);
and UO_2108 (O_2108,N_19880,N_19023);
nor UO_2109 (O_2109,N_19063,N_19052);
nand UO_2110 (O_2110,N_19949,N_19352);
xnor UO_2111 (O_2111,N_19575,N_19029);
xor UO_2112 (O_2112,N_19457,N_19191);
nor UO_2113 (O_2113,N_19603,N_19960);
and UO_2114 (O_2114,N_19903,N_19566);
or UO_2115 (O_2115,N_19400,N_19049);
or UO_2116 (O_2116,N_19762,N_19473);
nor UO_2117 (O_2117,N_19315,N_19085);
xnor UO_2118 (O_2118,N_19694,N_19083);
nand UO_2119 (O_2119,N_19551,N_19235);
and UO_2120 (O_2120,N_19935,N_19809);
or UO_2121 (O_2121,N_19698,N_19658);
xnor UO_2122 (O_2122,N_19884,N_19744);
or UO_2123 (O_2123,N_19185,N_19363);
xor UO_2124 (O_2124,N_19750,N_19235);
and UO_2125 (O_2125,N_19772,N_19840);
and UO_2126 (O_2126,N_19791,N_19450);
xor UO_2127 (O_2127,N_19626,N_19900);
xnor UO_2128 (O_2128,N_19797,N_19965);
and UO_2129 (O_2129,N_19219,N_19082);
nand UO_2130 (O_2130,N_19681,N_19461);
xor UO_2131 (O_2131,N_19543,N_19627);
and UO_2132 (O_2132,N_19629,N_19119);
nand UO_2133 (O_2133,N_19117,N_19184);
and UO_2134 (O_2134,N_19462,N_19786);
and UO_2135 (O_2135,N_19565,N_19018);
nor UO_2136 (O_2136,N_19435,N_19529);
or UO_2137 (O_2137,N_19334,N_19320);
xor UO_2138 (O_2138,N_19585,N_19829);
nand UO_2139 (O_2139,N_19028,N_19290);
xor UO_2140 (O_2140,N_19532,N_19062);
xnor UO_2141 (O_2141,N_19090,N_19557);
nor UO_2142 (O_2142,N_19993,N_19576);
nand UO_2143 (O_2143,N_19137,N_19727);
nand UO_2144 (O_2144,N_19053,N_19835);
and UO_2145 (O_2145,N_19839,N_19759);
and UO_2146 (O_2146,N_19378,N_19328);
xnor UO_2147 (O_2147,N_19235,N_19611);
nor UO_2148 (O_2148,N_19339,N_19937);
nor UO_2149 (O_2149,N_19153,N_19145);
or UO_2150 (O_2150,N_19283,N_19022);
nand UO_2151 (O_2151,N_19095,N_19006);
or UO_2152 (O_2152,N_19208,N_19134);
xor UO_2153 (O_2153,N_19583,N_19602);
and UO_2154 (O_2154,N_19519,N_19525);
xor UO_2155 (O_2155,N_19841,N_19491);
xor UO_2156 (O_2156,N_19912,N_19798);
or UO_2157 (O_2157,N_19757,N_19556);
nand UO_2158 (O_2158,N_19505,N_19344);
xnor UO_2159 (O_2159,N_19564,N_19249);
nand UO_2160 (O_2160,N_19219,N_19264);
or UO_2161 (O_2161,N_19891,N_19445);
xor UO_2162 (O_2162,N_19371,N_19518);
nand UO_2163 (O_2163,N_19207,N_19714);
nor UO_2164 (O_2164,N_19118,N_19574);
and UO_2165 (O_2165,N_19673,N_19530);
xnor UO_2166 (O_2166,N_19452,N_19531);
and UO_2167 (O_2167,N_19277,N_19287);
nor UO_2168 (O_2168,N_19657,N_19962);
and UO_2169 (O_2169,N_19582,N_19725);
xor UO_2170 (O_2170,N_19151,N_19625);
nor UO_2171 (O_2171,N_19393,N_19692);
xor UO_2172 (O_2172,N_19723,N_19789);
nand UO_2173 (O_2173,N_19559,N_19610);
and UO_2174 (O_2174,N_19805,N_19853);
or UO_2175 (O_2175,N_19264,N_19667);
xnor UO_2176 (O_2176,N_19050,N_19043);
nor UO_2177 (O_2177,N_19188,N_19410);
nor UO_2178 (O_2178,N_19643,N_19060);
or UO_2179 (O_2179,N_19293,N_19869);
xor UO_2180 (O_2180,N_19455,N_19208);
xor UO_2181 (O_2181,N_19664,N_19886);
nand UO_2182 (O_2182,N_19579,N_19004);
nand UO_2183 (O_2183,N_19537,N_19608);
nand UO_2184 (O_2184,N_19279,N_19860);
or UO_2185 (O_2185,N_19457,N_19169);
xor UO_2186 (O_2186,N_19705,N_19695);
or UO_2187 (O_2187,N_19137,N_19519);
nand UO_2188 (O_2188,N_19658,N_19970);
and UO_2189 (O_2189,N_19235,N_19174);
xor UO_2190 (O_2190,N_19484,N_19335);
nor UO_2191 (O_2191,N_19000,N_19277);
nor UO_2192 (O_2192,N_19356,N_19433);
nor UO_2193 (O_2193,N_19432,N_19533);
and UO_2194 (O_2194,N_19916,N_19790);
and UO_2195 (O_2195,N_19476,N_19006);
or UO_2196 (O_2196,N_19725,N_19577);
nand UO_2197 (O_2197,N_19573,N_19791);
and UO_2198 (O_2198,N_19877,N_19980);
xnor UO_2199 (O_2199,N_19263,N_19758);
xor UO_2200 (O_2200,N_19805,N_19209);
xnor UO_2201 (O_2201,N_19768,N_19255);
nand UO_2202 (O_2202,N_19963,N_19052);
or UO_2203 (O_2203,N_19264,N_19657);
nor UO_2204 (O_2204,N_19007,N_19860);
nand UO_2205 (O_2205,N_19602,N_19961);
and UO_2206 (O_2206,N_19901,N_19818);
nand UO_2207 (O_2207,N_19300,N_19941);
and UO_2208 (O_2208,N_19668,N_19371);
nand UO_2209 (O_2209,N_19346,N_19363);
nand UO_2210 (O_2210,N_19540,N_19274);
nor UO_2211 (O_2211,N_19133,N_19594);
nand UO_2212 (O_2212,N_19690,N_19514);
xnor UO_2213 (O_2213,N_19116,N_19063);
xnor UO_2214 (O_2214,N_19218,N_19336);
xnor UO_2215 (O_2215,N_19389,N_19589);
and UO_2216 (O_2216,N_19072,N_19433);
xnor UO_2217 (O_2217,N_19469,N_19010);
or UO_2218 (O_2218,N_19030,N_19993);
nor UO_2219 (O_2219,N_19703,N_19546);
nor UO_2220 (O_2220,N_19644,N_19160);
nor UO_2221 (O_2221,N_19097,N_19245);
nand UO_2222 (O_2222,N_19722,N_19721);
xnor UO_2223 (O_2223,N_19159,N_19421);
nand UO_2224 (O_2224,N_19937,N_19035);
nand UO_2225 (O_2225,N_19434,N_19411);
xnor UO_2226 (O_2226,N_19738,N_19689);
nand UO_2227 (O_2227,N_19831,N_19146);
and UO_2228 (O_2228,N_19302,N_19713);
nand UO_2229 (O_2229,N_19832,N_19119);
or UO_2230 (O_2230,N_19471,N_19061);
nand UO_2231 (O_2231,N_19055,N_19781);
nor UO_2232 (O_2232,N_19469,N_19434);
nor UO_2233 (O_2233,N_19919,N_19100);
xnor UO_2234 (O_2234,N_19028,N_19964);
nand UO_2235 (O_2235,N_19505,N_19533);
or UO_2236 (O_2236,N_19113,N_19537);
or UO_2237 (O_2237,N_19494,N_19943);
xor UO_2238 (O_2238,N_19292,N_19286);
and UO_2239 (O_2239,N_19507,N_19253);
and UO_2240 (O_2240,N_19126,N_19777);
nor UO_2241 (O_2241,N_19779,N_19388);
xnor UO_2242 (O_2242,N_19298,N_19710);
xor UO_2243 (O_2243,N_19933,N_19306);
and UO_2244 (O_2244,N_19033,N_19205);
nor UO_2245 (O_2245,N_19001,N_19107);
nand UO_2246 (O_2246,N_19510,N_19757);
xor UO_2247 (O_2247,N_19840,N_19876);
and UO_2248 (O_2248,N_19266,N_19993);
and UO_2249 (O_2249,N_19741,N_19245);
or UO_2250 (O_2250,N_19418,N_19163);
xor UO_2251 (O_2251,N_19792,N_19656);
or UO_2252 (O_2252,N_19386,N_19559);
xor UO_2253 (O_2253,N_19289,N_19778);
nand UO_2254 (O_2254,N_19737,N_19242);
xnor UO_2255 (O_2255,N_19267,N_19147);
nor UO_2256 (O_2256,N_19700,N_19290);
nand UO_2257 (O_2257,N_19592,N_19119);
nor UO_2258 (O_2258,N_19670,N_19451);
or UO_2259 (O_2259,N_19803,N_19870);
or UO_2260 (O_2260,N_19996,N_19657);
nand UO_2261 (O_2261,N_19592,N_19656);
xnor UO_2262 (O_2262,N_19795,N_19565);
or UO_2263 (O_2263,N_19919,N_19905);
nor UO_2264 (O_2264,N_19686,N_19498);
nand UO_2265 (O_2265,N_19505,N_19253);
or UO_2266 (O_2266,N_19757,N_19334);
or UO_2267 (O_2267,N_19674,N_19166);
and UO_2268 (O_2268,N_19888,N_19920);
or UO_2269 (O_2269,N_19476,N_19817);
or UO_2270 (O_2270,N_19491,N_19254);
or UO_2271 (O_2271,N_19250,N_19321);
or UO_2272 (O_2272,N_19011,N_19638);
and UO_2273 (O_2273,N_19208,N_19595);
or UO_2274 (O_2274,N_19853,N_19975);
or UO_2275 (O_2275,N_19479,N_19267);
xnor UO_2276 (O_2276,N_19626,N_19176);
nor UO_2277 (O_2277,N_19182,N_19555);
nand UO_2278 (O_2278,N_19622,N_19949);
nor UO_2279 (O_2279,N_19327,N_19866);
and UO_2280 (O_2280,N_19565,N_19536);
xnor UO_2281 (O_2281,N_19964,N_19290);
or UO_2282 (O_2282,N_19769,N_19809);
nor UO_2283 (O_2283,N_19421,N_19492);
nand UO_2284 (O_2284,N_19165,N_19785);
or UO_2285 (O_2285,N_19807,N_19550);
nor UO_2286 (O_2286,N_19429,N_19329);
or UO_2287 (O_2287,N_19618,N_19499);
nand UO_2288 (O_2288,N_19774,N_19572);
nor UO_2289 (O_2289,N_19597,N_19935);
or UO_2290 (O_2290,N_19620,N_19204);
xnor UO_2291 (O_2291,N_19365,N_19753);
xor UO_2292 (O_2292,N_19139,N_19597);
xor UO_2293 (O_2293,N_19052,N_19295);
xor UO_2294 (O_2294,N_19568,N_19718);
or UO_2295 (O_2295,N_19453,N_19856);
or UO_2296 (O_2296,N_19665,N_19556);
nand UO_2297 (O_2297,N_19224,N_19660);
nor UO_2298 (O_2298,N_19636,N_19779);
xor UO_2299 (O_2299,N_19097,N_19885);
nor UO_2300 (O_2300,N_19742,N_19868);
xor UO_2301 (O_2301,N_19837,N_19234);
nand UO_2302 (O_2302,N_19320,N_19680);
and UO_2303 (O_2303,N_19701,N_19420);
nand UO_2304 (O_2304,N_19020,N_19103);
or UO_2305 (O_2305,N_19620,N_19527);
or UO_2306 (O_2306,N_19822,N_19407);
nand UO_2307 (O_2307,N_19961,N_19355);
xor UO_2308 (O_2308,N_19498,N_19416);
nand UO_2309 (O_2309,N_19076,N_19658);
or UO_2310 (O_2310,N_19753,N_19737);
and UO_2311 (O_2311,N_19552,N_19265);
nand UO_2312 (O_2312,N_19890,N_19603);
and UO_2313 (O_2313,N_19756,N_19118);
nand UO_2314 (O_2314,N_19773,N_19619);
nor UO_2315 (O_2315,N_19563,N_19427);
and UO_2316 (O_2316,N_19866,N_19232);
nor UO_2317 (O_2317,N_19951,N_19544);
nand UO_2318 (O_2318,N_19026,N_19870);
xor UO_2319 (O_2319,N_19974,N_19680);
and UO_2320 (O_2320,N_19567,N_19807);
nand UO_2321 (O_2321,N_19416,N_19767);
nand UO_2322 (O_2322,N_19237,N_19585);
xnor UO_2323 (O_2323,N_19252,N_19389);
and UO_2324 (O_2324,N_19420,N_19891);
nand UO_2325 (O_2325,N_19977,N_19339);
or UO_2326 (O_2326,N_19394,N_19694);
xor UO_2327 (O_2327,N_19742,N_19263);
nand UO_2328 (O_2328,N_19991,N_19646);
xnor UO_2329 (O_2329,N_19254,N_19400);
xor UO_2330 (O_2330,N_19293,N_19025);
or UO_2331 (O_2331,N_19490,N_19425);
and UO_2332 (O_2332,N_19746,N_19636);
nor UO_2333 (O_2333,N_19366,N_19759);
xnor UO_2334 (O_2334,N_19845,N_19256);
or UO_2335 (O_2335,N_19689,N_19493);
nand UO_2336 (O_2336,N_19669,N_19497);
or UO_2337 (O_2337,N_19313,N_19492);
or UO_2338 (O_2338,N_19482,N_19334);
and UO_2339 (O_2339,N_19283,N_19926);
nor UO_2340 (O_2340,N_19410,N_19222);
and UO_2341 (O_2341,N_19602,N_19863);
and UO_2342 (O_2342,N_19864,N_19214);
xnor UO_2343 (O_2343,N_19206,N_19307);
nor UO_2344 (O_2344,N_19658,N_19894);
or UO_2345 (O_2345,N_19142,N_19373);
or UO_2346 (O_2346,N_19486,N_19499);
nand UO_2347 (O_2347,N_19825,N_19593);
nor UO_2348 (O_2348,N_19348,N_19857);
xor UO_2349 (O_2349,N_19838,N_19707);
nor UO_2350 (O_2350,N_19667,N_19503);
nand UO_2351 (O_2351,N_19196,N_19136);
nand UO_2352 (O_2352,N_19512,N_19439);
nor UO_2353 (O_2353,N_19308,N_19185);
nand UO_2354 (O_2354,N_19979,N_19194);
or UO_2355 (O_2355,N_19100,N_19451);
nand UO_2356 (O_2356,N_19648,N_19823);
nor UO_2357 (O_2357,N_19319,N_19541);
xnor UO_2358 (O_2358,N_19792,N_19698);
xor UO_2359 (O_2359,N_19102,N_19985);
nor UO_2360 (O_2360,N_19592,N_19911);
nor UO_2361 (O_2361,N_19288,N_19827);
nand UO_2362 (O_2362,N_19842,N_19047);
or UO_2363 (O_2363,N_19808,N_19053);
or UO_2364 (O_2364,N_19702,N_19089);
xnor UO_2365 (O_2365,N_19218,N_19823);
xnor UO_2366 (O_2366,N_19014,N_19497);
nor UO_2367 (O_2367,N_19692,N_19014);
nand UO_2368 (O_2368,N_19124,N_19776);
xor UO_2369 (O_2369,N_19259,N_19936);
and UO_2370 (O_2370,N_19870,N_19076);
xnor UO_2371 (O_2371,N_19977,N_19547);
xor UO_2372 (O_2372,N_19469,N_19716);
or UO_2373 (O_2373,N_19833,N_19568);
or UO_2374 (O_2374,N_19456,N_19278);
nor UO_2375 (O_2375,N_19881,N_19823);
or UO_2376 (O_2376,N_19738,N_19300);
and UO_2377 (O_2377,N_19559,N_19323);
and UO_2378 (O_2378,N_19838,N_19500);
xnor UO_2379 (O_2379,N_19956,N_19009);
nor UO_2380 (O_2380,N_19962,N_19636);
nor UO_2381 (O_2381,N_19496,N_19261);
or UO_2382 (O_2382,N_19822,N_19887);
or UO_2383 (O_2383,N_19403,N_19748);
xor UO_2384 (O_2384,N_19318,N_19515);
nand UO_2385 (O_2385,N_19879,N_19383);
xor UO_2386 (O_2386,N_19351,N_19962);
nand UO_2387 (O_2387,N_19964,N_19116);
xnor UO_2388 (O_2388,N_19232,N_19257);
or UO_2389 (O_2389,N_19404,N_19323);
xnor UO_2390 (O_2390,N_19509,N_19011);
and UO_2391 (O_2391,N_19566,N_19399);
nand UO_2392 (O_2392,N_19620,N_19807);
and UO_2393 (O_2393,N_19364,N_19218);
and UO_2394 (O_2394,N_19573,N_19784);
nor UO_2395 (O_2395,N_19508,N_19951);
nor UO_2396 (O_2396,N_19182,N_19863);
nand UO_2397 (O_2397,N_19038,N_19752);
and UO_2398 (O_2398,N_19947,N_19496);
nand UO_2399 (O_2399,N_19598,N_19318);
or UO_2400 (O_2400,N_19831,N_19793);
nand UO_2401 (O_2401,N_19875,N_19424);
and UO_2402 (O_2402,N_19107,N_19123);
nand UO_2403 (O_2403,N_19837,N_19481);
nand UO_2404 (O_2404,N_19607,N_19636);
or UO_2405 (O_2405,N_19769,N_19510);
or UO_2406 (O_2406,N_19763,N_19405);
nor UO_2407 (O_2407,N_19367,N_19556);
nand UO_2408 (O_2408,N_19579,N_19377);
and UO_2409 (O_2409,N_19179,N_19924);
nor UO_2410 (O_2410,N_19022,N_19405);
or UO_2411 (O_2411,N_19985,N_19485);
xnor UO_2412 (O_2412,N_19237,N_19354);
or UO_2413 (O_2413,N_19073,N_19393);
and UO_2414 (O_2414,N_19825,N_19434);
and UO_2415 (O_2415,N_19593,N_19566);
or UO_2416 (O_2416,N_19005,N_19725);
and UO_2417 (O_2417,N_19746,N_19379);
xor UO_2418 (O_2418,N_19701,N_19918);
and UO_2419 (O_2419,N_19479,N_19622);
xnor UO_2420 (O_2420,N_19225,N_19000);
and UO_2421 (O_2421,N_19651,N_19591);
and UO_2422 (O_2422,N_19146,N_19309);
or UO_2423 (O_2423,N_19602,N_19238);
and UO_2424 (O_2424,N_19317,N_19167);
and UO_2425 (O_2425,N_19405,N_19683);
nand UO_2426 (O_2426,N_19384,N_19558);
nor UO_2427 (O_2427,N_19498,N_19243);
nor UO_2428 (O_2428,N_19268,N_19536);
xnor UO_2429 (O_2429,N_19664,N_19550);
nand UO_2430 (O_2430,N_19343,N_19766);
xor UO_2431 (O_2431,N_19437,N_19953);
nor UO_2432 (O_2432,N_19400,N_19939);
or UO_2433 (O_2433,N_19244,N_19413);
nand UO_2434 (O_2434,N_19673,N_19888);
or UO_2435 (O_2435,N_19402,N_19459);
nor UO_2436 (O_2436,N_19449,N_19781);
xor UO_2437 (O_2437,N_19702,N_19177);
nand UO_2438 (O_2438,N_19824,N_19906);
nor UO_2439 (O_2439,N_19541,N_19575);
or UO_2440 (O_2440,N_19836,N_19010);
and UO_2441 (O_2441,N_19729,N_19412);
xor UO_2442 (O_2442,N_19907,N_19838);
and UO_2443 (O_2443,N_19992,N_19887);
and UO_2444 (O_2444,N_19548,N_19073);
nor UO_2445 (O_2445,N_19512,N_19077);
and UO_2446 (O_2446,N_19117,N_19843);
xor UO_2447 (O_2447,N_19253,N_19594);
nor UO_2448 (O_2448,N_19639,N_19206);
nand UO_2449 (O_2449,N_19075,N_19782);
and UO_2450 (O_2450,N_19927,N_19215);
or UO_2451 (O_2451,N_19113,N_19689);
nor UO_2452 (O_2452,N_19638,N_19012);
nor UO_2453 (O_2453,N_19662,N_19642);
and UO_2454 (O_2454,N_19643,N_19447);
nand UO_2455 (O_2455,N_19242,N_19401);
or UO_2456 (O_2456,N_19498,N_19476);
or UO_2457 (O_2457,N_19768,N_19840);
xor UO_2458 (O_2458,N_19050,N_19227);
or UO_2459 (O_2459,N_19926,N_19426);
nor UO_2460 (O_2460,N_19978,N_19488);
nor UO_2461 (O_2461,N_19998,N_19708);
nand UO_2462 (O_2462,N_19739,N_19271);
or UO_2463 (O_2463,N_19626,N_19497);
or UO_2464 (O_2464,N_19593,N_19258);
xor UO_2465 (O_2465,N_19110,N_19822);
and UO_2466 (O_2466,N_19737,N_19650);
nor UO_2467 (O_2467,N_19417,N_19553);
xnor UO_2468 (O_2468,N_19452,N_19694);
and UO_2469 (O_2469,N_19096,N_19666);
nor UO_2470 (O_2470,N_19048,N_19584);
and UO_2471 (O_2471,N_19529,N_19526);
nand UO_2472 (O_2472,N_19414,N_19040);
and UO_2473 (O_2473,N_19881,N_19134);
and UO_2474 (O_2474,N_19703,N_19749);
nand UO_2475 (O_2475,N_19006,N_19874);
nor UO_2476 (O_2476,N_19999,N_19497);
or UO_2477 (O_2477,N_19166,N_19245);
nor UO_2478 (O_2478,N_19505,N_19823);
nor UO_2479 (O_2479,N_19316,N_19002);
and UO_2480 (O_2480,N_19279,N_19754);
nand UO_2481 (O_2481,N_19650,N_19847);
or UO_2482 (O_2482,N_19678,N_19142);
xor UO_2483 (O_2483,N_19717,N_19818);
nand UO_2484 (O_2484,N_19269,N_19064);
nor UO_2485 (O_2485,N_19552,N_19612);
nand UO_2486 (O_2486,N_19123,N_19697);
or UO_2487 (O_2487,N_19440,N_19658);
nand UO_2488 (O_2488,N_19399,N_19489);
and UO_2489 (O_2489,N_19089,N_19045);
or UO_2490 (O_2490,N_19076,N_19860);
or UO_2491 (O_2491,N_19323,N_19561);
nand UO_2492 (O_2492,N_19188,N_19548);
and UO_2493 (O_2493,N_19986,N_19390);
and UO_2494 (O_2494,N_19892,N_19273);
nand UO_2495 (O_2495,N_19979,N_19716);
or UO_2496 (O_2496,N_19791,N_19859);
or UO_2497 (O_2497,N_19120,N_19544);
and UO_2498 (O_2498,N_19340,N_19488);
or UO_2499 (O_2499,N_19789,N_19522);
endmodule