module basic_1000_10000_1500_50_levels_2xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nand U0 (N_0,In_248,In_71);
nand U1 (N_1,In_466,In_717);
nor U2 (N_2,In_526,In_806);
or U3 (N_3,In_225,In_97);
nand U4 (N_4,In_131,In_651);
nor U5 (N_5,In_317,In_306);
and U6 (N_6,In_856,In_340);
nor U7 (N_7,In_375,In_871);
nor U8 (N_8,In_984,In_289);
and U9 (N_9,In_274,In_851);
or U10 (N_10,In_218,In_534);
or U11 (N_11,In_140,In_293);
and U12 (N_12,In_518,In_144);
or U13 (N_13,In_133,In_76);
nor U14 (N_14,In_88,In_100);
and U15 (N_15,In_496,In_124);
or U16 (N_16,In_908,In_26);
nor U17 (N_17,In_882,In_721);
nand U18 (N_18,In_497,In_290);
nor U19 (N_19,In_404,In_962);
nor U20 (N_20,In_96,In_555);
nand U21 (N_21,In_792,In_7);
and U22 (N_22,In_85,In_460);
and U23 (N_23,In_125,In_59);
nor U24 (N_24,In_780,In_535);
nand U25 (N_25,In_401,In_513);
nor U26 (N_26,In_938,In_132);
or U27 (N_27,In_318,In_590);
and U28 (N_28,In_729,In_628);
nand U29 (N_29,In_32,In_454);
or U30 (N_30,In_839,In_393);
or U31 (N_31,In_808,In_752);
nand U32 (N_32,In_79,In_834);
nor U33 (N_33,In_202,In_431);
or U34 (N_34,In_942,In_127);
or U35 (N_35,In_996,In_877);
or U36 (N_36,In_870,In_146);
nor U37 (N_37,In_945,In_700);
xor U38 (N_38,In_272,In_970);
nor U39 (N_39,In_120,In_621);
nor U40 (N_40,In_482,In_686);
nor U41 (N_41,In_241,In_119);
nand U42 (N_42,In_911,In_972);
and U43 (N_43,In_81,In_958);
or U44 (N_44,In_749,In_742);
and U45 (N_45,In_315,In_593);
nand U46 (N_46,In_776,In_400);
nand U47 (N_47,In_398,In_874);
and U48 (N_48,In_585,In_34);
or U49 (N_49,In_50,In_502);
and U50 (N_50,In_109,In_656);
or U51 (N_51,In_521,In_715);
nand U52 (N_52,In_793,In_909);
or U53 (N_53,In_764,In_149);
and U54 (N_54,In_688,In_990);
xnor U55 (N_55,In_444,In_250);
nor U56 (N_56,In_410,In_150);
or U57 (N_57,In_963,In_260);
nor U58 (N_58,In_452,In_761);
or U59 (N_59,In_872,In_505);
and U60 (N_60,In_292,In_989);
and U61 (N_61,In_592,In_731);
or U62 (N_62,In_933,In_33);
or U63 (N_63,In_435,In_671);
nor U64 (N_64,In_470,In_756);
nand U65 (N_65,In_895,In_240);
and U66 (N_66,In_38,In_524);
xnor U67 (N_67,In_489,In_301);
or U68 (N_68,In_845,In_203);
nand U69 (N_69,In_354,In_840);
nand U70 (N_70,In_860,In_921);
nor U71 (N_71,In_214,In_771);
and U72 (N_72,In_216,In_447);
or U73 (N_73,In_672,In_319);
and U74 (N_74,In_416,In_605);
or U75 (N_75,In_819,In_625);
nand U76 (N_76,In_620,In_221);
nor U77 (N_77,In_881,In_779);
nor U78 (N_78,In_713,In_186);
and U79 (N_79,In_817,In_423);
or U80 (N_80,In_812,In_153);
or U81 (N_81,In_259,In_428);
or U82 (N_82,In_980,In_956);
and U83 (N_83,In_481,In_598);
nand U84 (N_84,In_782,In_645);
nand U85 (N_85,In_987,In_352);
or U86 (N_86,In_491,In_701);
nand U87 (N_87,In_44,In_693);
and U88 (N_88,In_334,In_1);
nor U89 (N_89,In_560,In_857);
nand U90 (N_90,In_276,In_99);
or U91 (N_91,In_210,In_308);
or U92 (N_92,In_784,In_356);
or U93 (N_93,In_608,In_46);
nor U94 (N_94,In_130,In_953);
nand U95 (N_95,In_951,In_583);
or U96 (N_96,In_16,In_166);
nand U97 (N_97,In_121,In_287);
or U98 (N_98,In_422,In_712);
nand U99 (N_99,In_878,In_284);
nand U100 (N_100,In_6,In_624);
nor U101 (N_101,In_200,In_324);
and U102 (N_102,In_519,In_763);
nand U103 (N_103,In_825,In_328);
nand U104 (N_104,In_329,In_440);
or U105 (N_105,In_969,In_873);
or U106 (N_106,In_949,In_421);
and U107 (N_107,In_189,In_243);
or U108 (N_108,In_134,In_252);
or U109 (N_109,In_233,In_662);
and U110 (N_110,In_735,In_90);
and U111 (N_111,In_683,In_687);
nand U112 (N_112,In_843,In_802);
and U113 (N_113,In_930,In_443);
nand U114 (N_114,In_530,In_462);
nor U115 (N_115,In_589,In_868);
and U116 (N_116,In_697,In_42);
and U117 (N_117,In_775,In_668);
or U118 (N_118,In_762,In_361);
nor U119 (N_119,In_72,In_93);
nor U120 (N_120,In_685,In_795);
nor U121 (N_121,In_343,In_254);
nor U122 (N_122,In_737,In_888);
nor U123 (N_123,In_377,In_809);
or U124 (N_124,In_271,In_704);
nand U125 (N_125,In_168,In_514);
or U126 (N_126,In_915,In_420);
nor U127 (N_127,In_245,In_234);
nor U128 (N_128,In_719,In_477);
nand U129 (N_129,In_709,In_769);
nor U130 (N_130,In_280,In_267);
nand U131 (N_131,In_531,In_927);
nand U132 (N_132,In_858,In_372);
nand U133 (N_133,In_249,In_547);
or U134 (N_134,In_17,In_407);
nand U135 (N_135,In_296,In_611);
nor U136 (N_136,In_786,In_538);
or U137 (N_137,In_931,In_914);
or U138 (N_138,In_902,In_955);
and U139 (N_139,In_4,In_787);
or U140 (N_140,In_223,In_607);
and U141 (N_141,In_18,In_741);
and U142 (N_142,In_13,In_618);
and U143 (N_143,In_275,In_307);
or U144 (N_144,In_601,In_371);
or U145 (N_145,In_395,In_488);
or U146 (N_146,In_926,In_396);
nor U147 (N_147,In_60,In_244);
or U148 (N_148,In_177,In_800);
or U149 (N_149,In_586,In_434);
or U150 (N_150,In_879,In_635);
or U151 (N_151,In_652,In_378);
nor U152 (N_152,In_865,In_569);
or U153 (N_153,In_773,In_610);
and U154 (N_154,In_449,In_522);
nand U155 (N_155,In_368,In_894);
or U156 (N_156,In_478,In_627);
nand U157 (N_157,In_884,In_486);
nand U158 (N_158,In_327,In_426);
and U159 (N_159,In_432,In_384);
nand U160 (N_160,In_630,In_537);
nand U161 (N_161,In_886,In_745);
nand U162 (N_162,In_600,In_78);
and U163 (N_163,In_405,In_357);
nor U164 (N_164,In_442,In_476);
and U165 (N_165,In_509,In_382);
or U166 (N_166,In_944,In_451);
and U167 (N_167,In_748,In_103);
or U168 (N_168,In_348,In_917);
nand U169 (N_169,In_999,In_781);
nor U170 (N_170,In_774,In_70);
nand U171 (N_171,In_811,In_545);
nor U172 (N_172,In_438,In_559);
and U173 (N_173,In_386,In_550);
nand U174 (N_174,In_302,In_880);
nor U175 (N_175,In_828,In_388);
nor U176 (N_176,In_824,In_362);
or U177 (N_177,In_936,In_413);
nor U178 (N_178,In_597,In_571);
nor U179 (N_179,In_41,In_567);
and U180 (N_180,In_394,In_54);
nand U181 (N_181,In_788,In_141);
nor U182 (N_182,In_409,In_30);
and U183 (N_183,In_558,In_772);
nand U184 (N_184,In_708,In_660);
or U185 (N_185,In_212,In_655);
nand U186 (N_186,In_118,In_650);
nor U187 (N_187,In_644,In_759);
nand U188 (N_188,In_543,In_137);
or U189 (N_189,In_445,In_948);
and U190 (N_190,In_8,In_667);
nor U191 (N_191,In_932,In_485);
nand U192 (N_192,In_151,In_504);
nand U193 (N_193,In_968,In_746);
nand U194 (N_194,In_457,In_602);
nor U195 (N_195,In_459,In_575);
or U196 (N_196,In_353,In_734);
nor U197 (N_197,In_580,In_235);
or U198 (N_198,In_916,In_294);
nand U199 (N_199,In_229,In_957);
and U200 (N_200,In_975,In_901);
and U201 (N_201,In_480,In_805);
and U202 (N_202,In_810,In_722);
and U203 (N_203,N_158,N_177);
and U204 (N_204,In_563,In_747);
nand U205 (N_205,N_185,In_39);
and U206 (N_206,In_653,In_501);
or U207 (N_207,In_510,In_833);
or U208 (N_208,In_247,In_947);
and U209 (N_209,N_127,In_172);
nor U210 (N_210,In_347,In_157);
nor U211 (N_211,N_77,In_219);
or U212 (N_212,In_689,In_129);
nor U213 (N_213,In_154,In_974);
and U214 (N_214,In_814,In_281);
or U215 (N_215,In_922,N_27);
and U216 (N_216,In_669,In_791);
nor U217 (N_217,In_866,In_570);
nor U218 (N_218,In_728,In_852);
and U219 (N_219,In_291,In_204);
or U220 (N_220,In_339,In_226);
xnor U221 (N_221,N_20,In_152);
or U222 (N_222,In_336,N_73);
xnor U223 (N_223,N_170,In_114);
nand U224 (N_224,In_441,In_475);
nor U225 (N_225,In_487,In_716);
or U226 (N_226,In_646,N_135);
and U227 (N_227,In_220,In_883);
or U228 (N_228,In_896,In_25);
xor U229 (N_229,In_211,In_63);
xor U230 (N_230,N_19,In_251);
nor U231 (N_231,N_119,N_65);
and U232 (N_232,In_572,N_124);
nand U233 (N_233,N_96,N_105);
and U234 (N_234,N_168,In_842);
and U235 (N_235,N_192,N_163);
and U236 (N_236,N_70,In_228);
and U237 (N_237,In_295,In_677);
or U238 (N_238,In_298,In_108);
or U239 (N_239,In_900,In_167);
or U240 (N_240,In_62,In_184);
nor U241 (N_241,In_193,In_66);
and U242 (N_242,In_511,N_150);
or U243 (N_243,N_58,In_224);
and U244 (N_244,N_33,In_123);
or U245 (N_245,In_821,In_503);
and U246 (N_246,In_217,In_924);
or U247 (N_247,N_118,In_699);
nor U248 (N_248,In_278,In_730);
and U249 (N_249,In_359,In_160);
or U250 (N_250,N_3,N_160);
nand U251 (N_251,In_606,In_588);
xnor U252 (N_252,In_379,In_29);
or U253 (N_253,In_813,In_40);
nor U254 (N_254,In_467,N_50);
and U255 (N_255,In_778,N_52);
nand U256 (N_256,In_982,N_172);
nor U257 (N_257,In_322,N_111);
nand U258 (N_258,In_913,In_777);
nor U259 (N_259,In_403,In_187);
and U260 (N_260,In_615,N_74);
and U261 (N_261,N_4,In_997);
nor U262 (N_262,N_23,In_979);
and U263 (N_263,In_27,In_562);
or U264 (N_264,In_316,In_208);
nand U265 (N_265,In_28,In_331);
and U266 (N_266,In_506,In_299);
and U267 (N_267,N_63,N_36);
or U268 (N_268,In_841,In_818);
nor U269 (N_269,N_162,In_68);
nor U270 (N_270,N_112,In_499);
and U271 (N_271,In_861,N_132);
or U272 (N_272,N_175,N_62);
and U273 (N_273,In_961,In_58);
nor U274 (N_274,N_95,In_549);
or U275 (N_275,In_55,N_47);
nand U276 (N_276,In_330,In_995);
nor U277 (N_277,In_564,In_849);
or U278 (N_278,In_684,In_711);
or U279 (N_279,N_171,In_623);
or U280 (N_280,In_707,In_231);
nand U281 (N_281,In_53,In_128);
and U282 (N_282,In_139,N_117);
nor U283 (N_283,N_102,In_390);
nand U284 (N_284,N_28,In_920);
or U285 (N_285,In_724,In_57);
nor U286 (N_286,In_262,N_98);
nand U287 (N_287,N_167,In_626);
or U288 (N_288,In_760,In_750);
nor U289 (N_289,N_179,In_227);
nand U290 (N_290,N_121,N_146);
and U291 (N_291,In_928,In_789);
nor U292 (N_292,In_551,In_389);
or U293 (N_293,N_152,In_138);
and U294 (N_294,N_141,In_631);
nor U295 (N_295,N_174,In_163);
nand U296 (N_296,N_71,In_529);
nand U297 (N_297,In_935,In_837);
nand U298 (N_298,In_471,In_110);
and U299 (N_299,In_65,In_617);
nand U300 (N_300,In_269,N_189);
nand U301 (N_301,N_21,In_536);
nand U302 (N_302,In_893,In_381);
nor U303 (N_303,N_44,In_702);
nand U304 (N_304,In_889,N_104);
or U305 (N_305,In_898,In_94);
nor U306 (N_306,N_144,In_494);
nand U307 (N_307,N_101,In_367);
or U308 (N_308,In_369,In_946);
nand U309 (N_309,In_766,In_213);
or U310 (N_310,In_215,N_8);
nand U311 (N_311,In_807,In_516);
nand U312 (N_312,In_176,In_582);
or U313 (N_313,In_179,In_885);
and U314 (N_314,In_767,In_678);
nand U315 (N_315,In_2,In_288);
nor U316 (N_316,In_320,N_34);
nand U317 (N_317,In_539,In_964);
or U318 (N_318,N_191,In_576);
or U319 (N_319,In_829,N_76);
nor U320 (N_320,N_7,In_691);
and U321 (N_321,In_540,N_106);
nand U322 (N_322,In_397,In_270);
and U323 (N_323,In_726,In_136);
or U324 (N_324,N_6,N_110);
nor U325 (N_325,N_136,N_198);
or U326 (N_326,In_976,In_84);
and U327 (N_327,In_816,In_392);
nor U328 (N_328,In_994,In_581);
and U329 (N_329,In_483,N_45);
nor U330 (N_330,N_108,In_145);
nand U331 (N_331,In_661,N_100);
or U332 (N_332,In_544,N_90);
or U333 (N_333,In_616,N_149);
or U334 (N_334,In_937,In_333);
nand U335 (N_335,N_46,In_863);
or U336 (N_336,In_998,In_798);
or U337 (N_337,In_207,N_22);
and U338 (N_338,In_910,N_182);
or U339 (N_339,In_692,In_633);
nand U340 (N_340,In_574,In_736);
or U341 (N_341,In_345,N_147);
nor U342 (N_342,In_753,N_68);
or U343 (N_343,In_342,In_614);
nor U344 (N_344,N_125,In_399);
or U345 (N_345,In_991,In_0);
nand U346 (N_346,In_351,In_439);
nand U347 (N_347,N_5,N_31);
nand U348 (N_348,In_847,In_246);
nand U349 (N_349,In_364,In_934);
nor U350 (N_350,In_642,N_24);
or U351 (N_351,N_13,In_433);
or U352 (N_352,In_674,In_566);
nand U353 (N_353,In_321,N_48);
nor U354 (N_354,In_402,N_196);
nor U355 (N_355,In_568,In_197);
or U356 (N_356,N_107,In_694);
nand U357 (N_357,In_658,In_238);
nand U358 (N_358,In_11,In_376);
and U359 (N_359,In_173,N_14);
or U360 (N_360,In_876,In_854);
nor U361 (N_361,In_523,In_20);
nor U362 (N_362,In_323,N_180);
or U363 (N_363,In_905,In_609);
and U364 (N_364,In_822,In_178);
nand U365 (N_365,In_733,In_458);
nor U366 (N_366,N_159,N_25);
nor U367 (N_367,In_21,In_770);
nand U368 (N_368,In_232,In_890);
nor U369 (N_369,In_51,In_67);
nor U370 (N_370,N_38,In_966);
nor U371 (N_371,In_195,In_565);
or U372 (N_372,N_148,In_468);
and U373 (N_373,In_106,In_801);
or U374 (N_374,In_257,In_417);
nor U375 (N_375,N_173,In_629);
or U376 (N_376,In_744,In_940);
nand U377 (N_377,In_256,In_727);
xor U378 (N_378,In_436,In_573);
nand U379 (N_379,In_527,In_10);
and U380 (N_380,In_309,In_619);
xnor U381 (N_381,In_579,In_169);
nor U382 (N_382,In_429,In_350);
and U383 (N_383,In_198,In_637);
nor U384 (N_384,In_22,In_277);
nand U385 (N_385,In_222,N_69);
and U386 (N_386,In_182,In_846);
nand U387 (N_387,In_622,In_310);
and U388 (N_388,In_666,In_665);
or U389 (N_389,In_48,In_263);
and U390 (N_390,In_595,In_332);
nor U391 (N_391,In_490,N_88);
nand U392 (N_392,N_181,In_188);
nor U393 (N_393,In_92,In_279);
nor U394 (N_394,In_255,N_113);
or U395 (N_395,In_64,N_164);
nor U396 (N_396,In_862,In_799);
nor U397 (N_397,In_335,N_129);
and U398 (N_398,In_365,N_12);
and U399 (N_399,In_236,In_919);
nor U400 (N_400,In_584,In_556);
nor U401 (N_401,In_408,In_918);
xor U402 (N_402,In_500,In_532);
nand U403 (N_403,N_134,N_184);
and U404 (N_404,In_493,In_815);
nand U405 (N_405,N_166,N_120);
xnor U406 (N_406,N_363,In_875);
nor U407 (N_407,N_1,In_768);
xnor U408 (N_408,N_351,In_366);
or U409 (N_409,In_869,N_392);
and U410 (N_410,N_257,In_9);
and U411 (N_411,N_264,In_698);
nand U412 (N_412,In_113,In_983);
nand U413 (N_413,In_673,In_180);
nand U414 (N_414,N_332,N_366);
nand U415 (N_415,N_85,In_69);
and U416 (N_416,In_725,N_313);
or U417 (N_417,N_138,N_330);
or U418 (N_418,N_390,N_320);
and U419 (N_419,N_251,N_268);
nor U420 (N_420,In_758,N_399);
nand U421 (N_421,N_388,N_261);
nand U422 (N_422,In_192,In_418);
and U423 (N_423,In_950,In_242);
nor U424 (N_424,N_140,In_446);
and U425 (N_425,In_751,N_317);
or U426 (N_426,N_37,In_196);
nand U427 (N_427,N_262,N_40);
nor U428 (N_428,In_971,In_52);
and U429 (N_429,In_385,N_126);
and U430 (N_430,N_256,N_333);
or U431 (N_431,N_271,In_143);
nor U432 (N_432,In_835,In_554);
and U433 (N_433,N_302,N_308);
and U434 (N_434,N_291,In_230);
nor U435 (N_435,N_373,N_339);
nor U436 (N_436,In_887,N_10);
nand U437 (N_437,N_2,In_533);
or U438 (N_438,N_263,N_224);
nand U439 (N_439,N_282,In_785);
or U440 (N_440,In_943,N_356);
xnor U441 (N_441,In_162,In_156);
and U442 (N_442,In_341,N_344);
nand U443 (N_443,N_115,N_331);
nor U444 (N_444,In_664,In_803);
or U445 (N_445,N_116,N_369);
nand U446 (N_446,In_670,In_304);
or U447 (N_447,N_240,In_300);
nand U448 (N_448,N_190,In_891);
nand U449 (N_449,In_206,N_329);
nor U450 (N_450,In_978,In_338);
nor U451 (N_451,N_87,In_515);
and U452 (N_452,In_325,In_850);
or U453 (N_453,In_406,In_696);
nand U454 (N_454,N_187,In_453);
and U455 (N_455,In_743,In_939);
nor U456 (N_456,N_368,In_237);
or U457 (N_457,N_137,N_321);
or U458 (N_458,N_336,N_139);
nand U459 (N_459,N_9,N_323);
nor U460 (N_460,In_101,N_169);
or U461 (N_461,In_718,N_337);
nand U462 (N_462,N_327,In_107);
or U463 (N_463,In_548,In_122);
nor U464 (N_464,N_383,N_156);
or U465 (N_465,N_215,N_371);
and U466 (N_466,N_377,In_591);
or U467 (N_467,In_844,In_720);
and U468 (N_468,N_280,In_639);
nor U469 (N_469,N_145,In_23);
nor U470 (N_470,N_188,N_209);
nand U471 (N_471,N_86,In_577);
nor U472 (N_472,N_393,N_355);
nor U473 (N_473,In_906,N_0);
or U474 (N_474,N_202,In_498);
nor U475 (N_475,N_53,N_229);
nand U476 (N_476,In_363,N_306);
and U477 (N_477,N_266,In_732);
nor U478 (N_478,In_820,N_296);
nand U479 (N_479,In_380,In_552);
or U480 (N_480,In_632,N_376);
nand U481 (N_481,N_303,N_238);
nor U482 (N_482,In_557,In_738);
nor U483 (N_483,N_287,In_604);
nand U484 (N_484,N_217,In_425);
nand U485 (N_485,In_448,In_190);
nor U486 (N_486,N_316,In_147);
or U487 (N_487,In_424,N_32);
nand U488 (N_488,In_19,In_261);
nor U489 (N_489,In_520,N_334);
nor U490 (N_490,N_60,In_517);
nand U491 (N_491,N_258,In_831);
or U492 (N_492,In_286,N_310);
and U493 (N_493,In_358,N_309);
or U494 (N_494,In_804,In_98);
nor U495 (N_495,In_492,N_360);
nor U496 (N_496,N_380,In_757);
nand U497 (N_497,N_353,N_91);
and U498 (N_498,In_484,N_59);
nor U499 (N_499,N_49,In_525);
and U500 (N_500,N_265,In_461);
nor U501 (N_501,N_197,N_250);
nand U502 (N_502,N_109,N_365);
nand U503 (N_503,In_427,N_276);
nand U504 (N_504,In_102,N_300);
or U505 (N_505,In_859,In_643);
and U506 (N_506,N_204,In_636);
nand U507 (N_507,N_157,In_903);
nor U508 (N_508,N_18,N_312);
or U509 (N_509,In_383,N_315);
nand U510 (N_510,In_148,N_212);
nand U511 (N_511,N_286,N_89);
and U512 (N_512,N_122,In_14);
or U513 (N_513,N_226,In_313);
or U514 (N_514,N_133,In_473);
nor U515 (N_515,In_191,In_283);
nand U516 (N_516,In_112,N_237);
and U517 (N_517,In_973,N_361);
nor U518 (N_518,In_508,N_247);
nand U519 (N_519,In_312,In_61);
and U520 (N_520,N_239,N_78);
nor U521 (N_521,N_200,In_897);
nand U522 (N_522,In_853,N_338);
or U523 (N_523,In_415,In_981);
nor U524 (N_524,N_26,In_649);
xor U525 (N_525,N_193,In_528);
and U526 (N_526,In_73,In_360);
and U527 (N_527,In_456,N_165);
and U528 (N_528,In_638,In_663);
and U529 (N_529,N_207,In_205);
or U530 (N_530,N_176,In_159);
nand U531 (N_531,N_80,N_72);
or U532 (N_532,In_104,In_3);
nand U533 (N_533,In_414,N_275);
xor U534 (N_534,In_464,N_252);
and U535 (N_535,N_272,In_373);
nand U536 (N_536,N_142,In_47);
nor U537 (N_537,N_382,In_797);
xor U538 (N_538,N_11,In_239);
nor U539 (N_539,In_171,N_210);
nor U540 (N_540,N_340,N_347);
and U541 (N_541,In_135,In_867);
nand U542 (N_542,In_297,N_227);
nor U543 (N_543,In_174,In_266);
and U544 (N_544,In_268,In_794);
nand U545 (N_545,N_213,N_66);
or U546 (N_546,In_126,N_241);
or U547 (N_547,In_561,In_370);
or U548 (N_548,In_864,N_178);
or U549 (N_549,In_594,N_29);
nor U550 (N_550,In_12,N_346);
nor U551 (N_551,In_115,In_155);
nand U552 (N_552,N_294,In_765);
nor U553 (N_553,N_364,In_929);
nor U554 (N_554,N_231,N_211);
and U555 (N_555,N_82,In_848);
nand U556 (N_556,N_260,N_234);
and U557 (N_557,N_290,In_105);
or U558 (N_558,In_314,In_941);
nand U559 (N_559,N_97,N_154);
xor U560 (N_560,In_706,In_391);
and U561 (N_561,N_161,In_679);
or U562 (N_562,In_904,In_892);
nor U563 (N_563,In_282,N_205);
or U564 (N_564,N_301,N_288);
nand U565 (N_565,N_379,N_389);
or U566 (N_566,N_341,In_832);
and U567 (N_567,N_79,In_739);
nand U568 (N_568,In_985,N_203);
or U569 (N_569,In_265,N_57);
nor U570 (N_570,N_143,N_386);
or U571 (N_571,In_986,In_654);
or U572 (N_572,N_367,In_754);
nand U573 (N_573,In_952,N_304);
nand U574 (N_574,N_41,N_285);
and U575 (N_575,In_412,N_269);
or U576 (N_576,N_99,N_318);
nand U577 (N_577,N_328,N_219);
and U578 (N_578,N_299,N_345);
nand U579 (N_579,In_648,N_378);
nand U580 (N_580,In_36,In_116);
nand U581 (N_581,N_155,In_553);
or U582 (N_582,In_31,In_634);
xnor U583 (N_583,N_206,In_142);
nor U584 (N_584,N_289,N_314);
and U585 (N_585,In_542,N_283);
or U586 (N_586,In_91,In_258);
and U587 (N_587,In_690,N_208);
nand U588 (N_588,In_49,N_103);
xnor U589 (N_589,N_246,N_222);
or U590 (N_590,In_960,N_279);
nand U591 (N_591,N_30,In_411);
and U592 (N_592,In_827,N_297);
nor U593 (N_593,N_395,In_185);
nand U594 (N_594,N_42,N_243);
or U595 (N_595,In_305,N_292);
or U596 (N_596,N_228,In_472);
and U597 (N_597,N_61,N_43);
nand U598 (N_598,In_912,In_437);
nor U599 (N_599,N_64,N_259);
and U600 (N_600,In_675,N_92);
and U601 (N_601,N_419,N_548);
nand U602 (N_602,N_556,N_358);
and U603 (N_603,N_568,N_199);
nor U604 (N_604,In_181,In_796);
nand U605 (N_605,In_15,In_45);
and U606 (N_606,N_153,N_434);
or U607 (N_607,In_273,N_16);
and U608 (N_608,N_426,In_264);
nor U609 (N_609,N_335,In_495);
nand U610 (N_610,In_790,In_680);
nor U611 (N_611,N_519,N_591);
nand U612 (N_612,In_855,N_558);
and U613 (N_613,N_580,N_39);
nand U614 (N_614,N_487,In_344);
nor U615 (N_615,N_83,In_965);
nand U616 (N_616,N_15,N_555);
nand U617 (N_617,N_539,N_438);
or U618 (N_618,N_236,N_582);
nor U619 (N_619,N_502,N_566);
or U620 (N_620,In_165,N_599);
nand U621 (N_621,N_455,N_131);
and U622 (N_622,N_93,N_510);
nor U623 (N_623,In_199,N_151);
nand U624 (N_624,In_988,N_547);
xnor U625 (N_625,N_518,N_472);
and U626 (N_626,In_612,In_285);
and U627 (N_627,N_442,In_326);
and U628 (N_628,N_417,N_587);
and U629 (N_629,N_403,N_576);
or U630 (N_630,N_521,N_281);
nand U631 (N_631,In_603,N_412);
and U632 (N_632,N_589,In_77);
nor U633 (N_633,N_374,N_407);
or U634 (N_634,N_75,N_427);
or U635 (N_635,In_647,In_682);
nand U636 (N_636,In_755,N_186);
and U637 (N_637,N_443,N_456);
and U638 (N_638,N_435,N_216);
and U639 (N_639,N_492,N_319);
and U640 (N_640,N_594,In_253);
nor U641 (N_641,In_907,In_899);
and U642 (N_642,N_420,N_491);
or U643 (N_643,N_509,N_496);
or U644 (N_644,N_531,N_586);
nand U645 (N_645,N_248,N_391);
and U646 (N_646,In_512,N_503);
and U647 (N_647,N_354,N_352);
or U648 (N_648,In_783,N_428);
and U649 (N_649,N_486,In_463);
nand U650 (N_650,N_569,In_455);
and U651 (N_651,N_35,In_923);
and U652 (N_652,N_463,N_592);
and U653 (N_653,N_574,N_221);
or U654 (N_654,N_422,N_423);
nand U655 (N_655,N_84,N_530);
and U656 (N_656,N_230,N_67);
nor U657 (N_657,N_563,N_557);
nor U658 (N_658,N_253,N_54);
or U659 (N_659,N_526,N_220);
nor U660 (N_660,N_481,In_450);
and U661 (N_661,In_35,In_161);
and U662 (N_662,N_56,N_450);
nand U663 (N_663,In_710,N_324);
nand U664 (N_664,N_498,N_490);
or U665 (N_665,N_577,In_681);
nor U666 (N_666,N_440,N_225);
xnor U667 (N_667,In_714,N_493);
nand U668 (N_668,N_402,In_387);
nand U669 (N_669,In_587,N_544);
nand U670 (N_670,N_512,In_74);
nor U671 (N_671,N_536,N_433);
or U672 (N_672,In_82,N_397);
nor U673 (N_673,N_342,N_460);
or U674 (N_674,N_533,N_552);
nand U675 (N_675,In_993,N_593);
or U676 (N_676,N_464,N_270);
or U677 (N_677,N_583,N_254);
nor U678 (N_678,In_346,N_578);
and U679 (N_679,N_410,N_545);
or U680 (N_680,In_37,In_703);
nor U681 (N_681,In_80,In_823);
nor U682 (N_682,In_640,N_218);
nor U683 (N_683,N_501,In_954);
or U684 (N_684,N_527,N_244);
nor U685 (N_685,N_404,In_546);
nand U686 (N_686,N_401,N_396);
nor U687 (N_687,N_384,N_232);
xor U688 (N_688,N_429,In_641);
nor U689 (N_689,N_362,In_303);
and U690 (N_690,N_284,N_416);
nor U691 (N_691,N_554,N_551);
and U692 (N_692,N_17,N_81);
nor U693 (N_693,In_474,In_925);
and U694 (N_694,N_476,N_541);
nand U695 (N_695,N_553,N_457);
or U696 (N_696,N_477,In_695);
nand U697 (N_697,N_559,N_567);
nand U698 (N_698,N_528,N_445);
nor U699 (N_699,N_585,In_507);
nor U700 (N_700,In_311,In_723);
nand U701 (N_701,In_89,N_408);
and U702 (N_702,In_337,In_967);
nor U703 (N_703,N_513,N_597);
or U704 (N_704,N_520,N_451);
and U705 (N_705,N_350,N_183);
or U706 (N_706,N_223,N_542);
and U707 (N_707,N_305,N_488);
nor U708 (N_708,N_277,In_164);
nand U709 (N_709,In_175,In_111);
and U710 (N_710,N_415,N_55);
nor U711 (N_711,In_705,N_595);
nor U712 (N_712,N_590,N_381);
nor U713 (N_713,N_130,N_575);
or U714 (N_714,N_94,In_613);
nand U715 (N_715,In_183,N_598);
nand U716 (N_716,N_499,N_515);
nor U717 (N_717,N_500,In_836);
and U718 (N_718,N_394,In_75);
nor U719 (N_719,N_516,In_977);
nor U720 (N_720,N_465,N_581);
nor U721 (N_721,N_448,N_255);
nor U722 (N_722,In_469,N_444);
or U723 (N_723,N_550,N_293);
nor U724 (N_724,N_128,N_267);
and U725 (N_725,In_374,N_480);
and U726 (N_726,N_495,In_95);
or U727 (N_727,N_572,N_461);
or U728 (N_728,In_86,N_298);
nor U729 (N_729,In_201,N_194);
nand U730 (N_730,N_579,N_370);
and U731 (N_731,N_233,N_508);
and U732 (N_732,N_538,In_158);
nand U733 (N_733,In_992,N_385);
nor U734 (N_734,N_245,In_541);
and U735 (N_735,N_505,N_561);
or U736 (N_736,In_87,N_235);
or U737 (N_737,In_5,N_406);
nor U738 (N_738,In_578,N_483);
and U739 (N_739,N_506,N_523);
nand U740 (N_740,N_549,N_504);
or U741 (N_741,N_471,N_537);
nand U742 (N_742,N_560,N_123);
xor U743 (N_743,N_398,In_479);
and U744 (N_744,In_430,N_357);
xor U745 (N_745,N_375,In_170);
xnor U746 (N_746,In_826,N_447);
nor U747 (N_747,N_458,N_485);
nand U748 (N_748,In_596,In_209);
nand U749 (N_749,N_469,N_430);
and U750 (N_750,In_117,N_425);
nor U751 (N_751,In_419,N_565);
xnor U752 (N_752,In_355,N_242);
nor U753 (N_753,N_475,N_359);
or U754 (N_754,N_372,N_274);
nand U755 (N_755,In_740,N_439);
or U756 (N_756,N_525,N_584);
and U757 (N_757,N_534,N_479);
nor U758 (N_758,N_466,N_311);
and U759 (N_759,N_441,N_201);
nand U760 (N_760,In_676,N_511);
nor U761 (N_761,N_343,In_83);
nor U762 (N_762,N_322,In_56);
nand U763 (N_763,N_529,N_562);
nor U764 (N_764,N_413,N_411);
nand U765 (N_765,N_452,N_418);
or U766 (N_766,N_409,N_387);
or U767 (N_767,N_524,N_195);
and U768 (N_768,N_414,N_514);
and U769 (N_769,N_295,N_467);
or U770 (N_770,N_424,N_573);
nand U771 (N_771,N_326,In_43);
or U772 (N_772,N_532,N_51);
and U773 (N_773,N_517,In_830);
nor U774 (N_774,N_474,N_405);
nand U775 (N_775,In_657,N_484);
or U776 (N_776,N_273,N_570);
or U777 (N_777,N_348,N_596);
nor U778 (N_778,N_432,N_468);
nand U779 (N_779,N_307,N_497);
or U780 (N_780,N_437,In_838);
and U781 (N_781,N_588,N_446);
nor U782 (N_782,In_349,In_194);
and U783 (N_783,N_543,N_494);
nor U784 (N_784,In_599,N_470);
nor U785 (N_785,N_473,N_507);
nand U786 (N_786,N_214,In_465);
nand U787 (N_787,N_546,N_449);
and U788 (N_788,N_400,N_114);
xor U789 (N_789,N_459,N_278);
or U790 (N_790,N_421,N_482);
nand U791 (N_791,N_454,In_959);
nor U792 (N_792,N_489,N_349);
nor U793 (N_793,N_249,N_431);
and U794 (N_794,N_571,N_462);
nand U795 (N_795,In_24,N_522);
and U796 (N_796,N_325,N_535);
and U797 (N_797,N_436,N_564);
nor U798 (N_798,N_478,N_540);
nand U799 (N_799,N_453,In_659);
and U800 (N_800,N_762,N_646);
nand U801 (N_801,N_702,N_700);
nand U802 (N_802,N_763,N_604);
nand U803 (N_803,N_798,N_660);
or U804 (N_804,N_701,N_754);
or U805 (N_805,N_687,N_792);
nand U806 (N_806,N_621,N_765);
or U807 (N_807,N_784,N_623);
and U808 (N_808,N_773,N_601);
nand U809 (N_809,N_723,N_799);
nor U810 (N_810,N_732,N_661);
or U811 (N_811,N_636,N_710);
nand U812 (N_812,N_649,N_603);
or U813 (N_813,N_709,N_635);
or U814 (N_814,N_731,N_712);
or U815 (N_815,N_776,N_714);
nand U816 (N_816,N_713,N_741);
nand U817 (N_817,N_655,N_629);
and U818 (N_818,N_653,N_654);
or U819 (N_819,N_766,N_613);
and U820 (N_820,N_694,N_727);
nor U821 (N_821,N_724,N_738);
nand U822 (N_822,N_602,N_683);
or U823 (N_823,N_698,N_674);
nand U824 (N_824,N_615,N_715);
xnor U825 (N_825,N_606,N_767);
or U826 (N_826,N_616,N_663);
nor U827 (N_827,N_600,N_786);
nand U828 (N_828,N_778,N_685);
nor U829 (N_829,N_764,N_611);
and U830 (N_830,N_617,N_774);
or U831 (N_831,N_612,N_691);
nand U832 (N_832,N_783,N_703);
nor U833 (N_833,N_684,N_642);
nor U834 (N_834,N_772,N_650);
or U835 (N_835,N_729,N_697);
and U836 (N_836,N_639,N_682);
nand U837 (N_837,N_777,N_749);
nand U838 (N_838,N_782,N_696);
or U839 (N_839,N_757,N_633);
and U840 (N_840,N_736,N_716);
nand U841 (N_841,N_705,N_728);
and U842 (N_842,N_672,N_662);
or U843 (N_843,N_718,N_659);
nand U844 (N_844,N_620,N_740);
nor U845 (N_845,N_630,N_758);
nand U846 (N_846,N_619,N_751);
nand U847 (N_847,N_607,N_711);
nand U848 (N_848,N_677,N_768);
and U849 (N_849,N_695,N_790);
or U850 (N_850,N_609,N_706);
or U851 (N_851,N_648,N_614);
nor U852 (N_852,N_761,N_622);
and U853 (N_853,N_708,N_690);
nand U854 (N_854,N_610,N_780);
nand U855 (N_855,N_689,N_647);
nor U856 (N_856,N_605,N_725);
nor U857 (N_857,N_669,N_671);
and U858 (N_858,N_771,N_752);
nand U859 (N_859,N_734,N_651);
nor U860 (N_860,N_722,N_668);
nor U861 (N_861,N_760,N_785);
or U862 (N_862,N_657,N_796);
nor U863 (N_863,N_769,N_618);
nand U864 (N_864,N_750,N_634);
nor U865 (N_865,N_656,N_681);
and U866 (N_866,N_626,N_673);
or U867 (N_867,N_733,N_746);
xor U868 (N_868,N_735,N_631);
xor U869 (N_869,N_688,N_666);
or U870 (N_870,N_781,N_795);
nor U871 (N_871,N_627,N_788);
or U872 (N_872,N_719,N_667);
nand U873 (N_873,N_624,N_787);
or U874 (N_874,N_726,N_756);
and U875 (N_875,N_789,N_676);
or U876 (N_876,N_720,N_608);
nand U877 (N_877,N_753,N_641);
nand U878 (N_878,N_704,N_721);
and U879 (N_879,N_678,N_730);
and U880 (N_880,N_686,N_744);
and U881 (N_881,N_759,N_675);
xor U882 (N_882,N_707,N_743);
nor U883 (N_883,N_644,N_739);
and U884 (N_884,N_679,N_794);
or U885 (N_885,N_747,N_791);
or U886 (N_886,N_652,N_638);
and U887 (N_887,N_755,N_770);
and U888 (N_888,N_665,N_717);
and U889 (N_889,N_670,N_640);
nor U890 (N_890,N_779,N_692);
nand U891 (N_891,N_693,N_775);
and U892 (N_892,N_645,N_628);
and U893 (N_893,N_793,N_699);
nand U894 (N_894,N_643,N_680);
nand U895 (N_895,N_745,N_625);
or U896 (N_896,N_664,N_637);
nand U897 (N_897,N_737,N_748);
nor U898 (N_898,N_632,N_742);
nand U899 (N_899,N_658,N_797);
xor U900 (N_900,N_687,N_686);
or U901 (N_901,N_745,N_670);
or U902 (N_902,N_626,N_760);
nand U903 (N_903,N_603,N_735);
xor U904 (N_904,N_679,N_657);
or U905 (N_905,N_707,N_694);
nor U906 (N_906,N_632,N_784);
nor U907 (N_907,N_666,N_656);
nor U908 (N_908,N_742,N_728);
nand U909 (N_909,N_617,N_733);
nand U910 (N_910,N_669,N_738);
nor U911 (N_911,N_603,N_698);
and U912 (N_912,N_628,N_746);
and U913 (N_913,N_697,N_645);
nor U914 (N_914,N_724,N_621);
nor U915 (N_915,N_751,N_779);
nor U916 (N_916,N_632,N_799);
nor U917 (N_917,N_758,N_605);
or U918 (N_918,N_766,N_614);
nor U919 (N_919,N_737,N_604);
and U920 (N_920,N_749,N_731);
nor U921 (N_921,N_780,N_738);
or U922 (N_922,N_773,N_750);
or U923 (N_923,N_677,N_617);
or U924 (N_924,N_662,N_780);
nor U925 (N_925,N_606,N_610);
or U926 (N_926,N_728,N_657);
xnor U927 (N_927,N_670,N_739);
and U928 (N_928,N_724,N_687);
and U929 (N_929,N_630,N_688);
and U930 (N_930,N_715,N_606);
and U931 (N_931,N_794,N_710);
and U932 (N_932,N_631,N_699);
or U933 (N_933,N_741,N_738);
or U934 (N_934,N_704,N_645);
nand U935 (N_935,N_627,N_684);
nand U936 (N_936,N_787,N_618);
xor U937 (N_937,N_756,N_745);
nand U938 (N_938,N_757,N_622);
nor U939 (N_939,N_789,N_775);
and U940 (N_940,N_718,N_664);
nor U941 (N_941,N_644,N_610);
nor U942 (N_942,N_687,N_769);
or U943 (N_943,N_796,N_702);
nand U944 (N_944,N_677,N_745);
and U945 (N_945,N_734,N_653);
nor U946 (N_946,N_768,N_775);
and U947 (N_947,N_672,N_610);
nand U948 (N_948,N_695,N_742);
and U949 (N_949,N_624,N_644);
nand U950 (N_950,N_767,N_754);
nor U951 (N_951,N_694,N_640);
nor U952 (N_952,N_797,N_633);
and U953 (N_953,N_710,N_632);
or U954 (N_954,N_781,N_724);
or U955 (N_955,N_630,N_729);
nand U956 (N_956,N_795,N_662);
and U957 (N_957,N_702,N_738);
and U958 (N_958,N_605,N_700);
nand U959 (N_959,N_772,N_761);
nand U960 (N_960,N_620,N_693);
or U961 (N_961,N_709,N_737);
and U962 (N_962,N_693,N_719);
and U963 (N_963,N_773,N_783);
nand U964 (N_964,N_609,N_611);
or U965 (N_965,N_780,N_778);
nand U966 (N_966,N_600,N_780);
nor U967 (N_967,N_721,N_648);
nand U968 (N_968,N_787,N_793);
nor U969 (N_969,N_652,N_626);
and U970 (N_970,N_721,N_660);
nor U971 (N_971,N_671,N_633);
and U972 (N_972,N_689,N_665);
and U973 (N_973,N_712,N_684);
and U974 (N_974,N_647,N_679);
nor U975 (N_975,N_776,N_788);
nand U976 (N_976,N_785,N_693);
xor U977 (N_977,N_750,N_644);
nor U978 (N_978,N_683,N_784);
nand U979 (N_979,N_775,N_750);
nand U980 (N_980,N_743,N_612);
nor U981 (N_981,N_706,N_723);
nand U982 (N_982,N_794,N_754);
and U983 (N_983,N_700,N_651);
nand U984 (N_984,N_793,N_681);
nand U985 (N_985,N_644,N_765);
nor U986 (N_986,N_799,N_654);
nor U987 (N_987,N_674,N_742);
or U988 (N_988,N_712,N_773);
or U989 (N_989,N_765,N_709);
and U990 (N_990,N_611,N_608);
and U991 (N_991,N_734,N_632);
nor U992 (N_992,N_643,N_755);
or U993 (N_993,N_777,N_735);
nor U994 (N_994,N_643,N_660);
nor U995 (N_995,N_646,N_739);
or U996 (N_996,N_625,N_731);
nand U997 (N_997,N_649,N_612);
and U998 (N_998,N_772,N_627);
or U999 (N_999,N_699,N_720);
nor U1000 (N_1000,N_909,N_807);
or U1001 (N_1001,N_998,N_981);
or U1002 (N_1002,N_929,N_954);
or U1003 (N_1003,N_991,N_983);
nand U1004 (N_1004,N_876,N_971);
and U1005 (N_1005,N_955,N_915);
nor U1006 (N_1006,N_801,N_838);
or U1007 (N_1007,N_905,N_943);
nor U1008 (N_1008,N_860,N_854);
and U1009 (N_1009,N_881,N_990);
and U1010 (N_1010,N_936,N_968);
nand U1011 (N_1011,N_977,N_864);
xnor U1012 (N_1012,N_960,N_997);
and U1013 (N_1013,N_853,N_809);
nand U1014 (N_1014,N_986,N_872);
nor U1015 (N_1015,N_850,N_966);
or U1016 (N_1016,N_994,N_873);
nor U1017 (N_1017,N_825,N_822);
nor U1018 (N_1018,N_871,N_842);
nor U1019 (N_1019,N_824,N_874);
nor U1020 (N_1020,N_805,N_914);
and U1021 (N_1021,N_878,N_973);
or U1022 (N_1022,N_826,N_904);
nor U1023 (N_1023,N_880,N_916);
nor U1024 (N_1024,N_887,N_867);
nand U1025 (N_1025,N_821,N_804);
and U1026 (N_1026,N_931,N_948);
and U1027 (N_1027,N_933,N_894);
nor U1028 (N_1028,N_843,N_819);
nand U1029 (N_1029,N_999,N_829);
or U1030 (N_1030,N_859,N_988);
nor U1031 (N_1031,N_925,N_811);
and U1032 (N_1032,N_951,N_861);
or U1033 (N_1033,N_852,N_942);
nand U1034 (N_1034,N_939,N_893);
and U1035 (N_1035,N_820,N_908);
nand U1036 (N_1036,N_906,N_803);
or U1037 (N_1037,N_984,N_982);
nand U1038 (N_1038,N_972,N_932);
and U1039 (N_1039,N_985,N_888);
xnor U1040 (N_1040,N_978,N_810);
nand U1041 (N_1041,N_800,N_993);
nor U1042 (N_1042,N_814,N_926);
or U1043 (N_1043,N_958,N_910);
nor U1044 (N_1044,N_987,N_827);
nor U1045 (N_1045,N_848,N_913);
nand U1046 (N_1046,N_862,N_815);
nand U1047 (N_1047,N_969,N_844);
nand U1048 (N_1048,N_901,N_956);
or U1049 (N_1049,N_828,N_980);
or U1050 (N_1050,N_947,N_961);
or U1051 (N_1051,N_866,N_930);
nand U1052 (N_1052,N_865,N_953);
nor U1053 (N_1053,N_989,N_875);
or U1054 (N_1054,N_856,N_938);
and U1055 (N_1055,N_917,N_802);
and U1056 (N_1056,N_835,N_941);
nor U1057 (N_1057,N_899,N_884);
or U1058 (N_1058,N_920,N_857);
or U1059 (N_1059,N_952,N_895);
nand U1060 (N_1060,N_911,N_992);
nand U1061 (N_1061,N_863,N_849);
nor U1062 (N_1062,N_927,N_995);
and U1063 (N_1063,N_922,N_975);
nor U1064 (N_1064,N_890,N_806);
nand U1065 (N_1065,N_879,N_897);
nor U1066 (N_1066,N_841,N_847);
or U1067 (N_1067,N_834,N_869);
or U1068 (N_1068,N_817,N_945);
and U1069 (N_1069,N_846,N_957);
or U1070 (N_1070,N_912,N_858);
and U1071 (N_1071,N_963,N_831);
or U1072 (N_1072,N_979,N_974);
and U1073 (N_1073,N_959,N_891);
and U1074 (N_1074,N_902,N_845);
nor U1075 (N_1075,N_921,N_907);
nand U1076 (N_1076,N_883,N_935);
nor U1077 (N_1077,N_976,N_839);
nor U1078 (N_1078,N_900,N_924);
nand U1079 (N_1079,N_896,N_812);
nand U1080 (N_1080,N_944,N_950);
nor U1081 (N_1081,N_882,N_816);
nand U1082 (N_1082,N_885,N_836);
nor U1083 (N_1083,N_937,N_918);
or U1084 (N_1084,N_877,N_919);
nor U1085 (N_1085,N_830,N_928);
and U1086 (N_1086,N_889,N_832);
or U1087 (N_1087,N_965,N_833);
or U1088 (N_1088,N_949,N_996);
and U1089 (N_1089,N_837,N_923);
nand U1090 (N_1090,N_818,N_940);
nand U1091 (N_1091,N_892,N_962);
and U1092 (N_1092,N_808,N_870);
nand U1093 (N_1093,N_886,N_855);
nor U1094 (N_1094,N_970,N_903);
nor U1095 (N_1095,N_851,N_934);
xor U1096 (N_1096,N_840,N_823);
or U1097 (N_1097,N_967,N_898);
or U1098 (N_1098,N_964,N_946);
xor U1099 (N_1099,N_868,N_813);
and U1100 (N_1100,N_829,N_985);
or U1101 (N_1101,N_873,N_849);
and U1102 (N_1102,N_942,N_883);
nor U1103 (N_1103,N_965,N_801);
nand U1104 (N_1104,N_872,N_978);
or U1105 (N_1105,N_943,N_915);
nand U1106 (N_1106,N_905,N_808);
or U1107 (N_1107,N_920,N_978);
nor U1108 (N_1108,N_954,N_979);
nor U1109 (N_1109,N_840,N_842);
nor U1110 (N_1110,N_989,N_980);
and U1111 (N_1111,N_848,N_967);
nand U1112 (N_1112,N_904,N_853);
nand U1113 (N_1113,N_822,N_943);
nand U1114 (N_1114,N_996,N_906);
nand U1115 (N_1115,N_838,N_802);
or U1116 (N_1116,N_907,N_946);
nor U1117 (N_1117,N_983,N_924);
or U1118 (N_1118,N_940,N_947);
nand U1119 (N_1119,N_804,N_897);
and U1120 (N_1120,N_806,N_901);
nor U1121 (N_1121,N_802,N_989);
nand U1122 (N_1122,N_854,N_849);
nor U1123 (N_1123,N_933,N_912);
and U1124 (N_1124,N_866,N_933);
and U1125 (N_1125,N_836,N_958);
nor U1126 (N_1126,N_955,N_916);
and U1127 (N_1127,N_936,N_975);
nand U1128 (N_1128,N_963,N_919);
nor U1129 (N_1129,N_972,N_897);
or U1130 (N_1130,N_806,N_976);
and U1131 (N_1131,N_818,N_903);
nor U1132 (N_1132,N_835,N_826);
nand U1133 (N_1133,N_911,N_917);
or U1134 (N_1134,N_914,N_970);
or U1135 (N_1135,N_958,N_846);
and U1136 (N_1136,N_981,N_880);
and U1137 (N_1137,N_949,N_840);
and U1138 (N_1138,N_857,N_840);
nor U1139 (N_1139,N_965,N_982);
nor U1140 (N_1140,N_953,N_912);
and U1141 (N_1141,N_879,N_918);
and U1142 (N_1142,N_807,N_875);
xor U1143 (N_1143,N_975,N_812);
nand U1144 (N_1144,N_839,N_966);
nand U1145 (N_1145,N_841,N_951);
nor U1146 (N_1146,N_887,N_990);
nor U1147 (N_1147,N_900,N_912);
and U1148 (N_1148,N_935,N_955);
nand U1149 (N_1149,N_944,N_832);
nand U1150 (N_1150,N_834,N_802);
or U1151 (N_1151,N_885,N_823);
nand U1152 (N_1152,N_858,N_915);
nor U1153 (N_1153,N_958,N_808);
and U1154 (N_1154,N_880,N_833);
nor U1155 (N_1155,N_951,N_849);
and U1156 (N_1156,N_891,N_841);
xnor U1157 (N_1157,N_997,N_975);
nor U1158 (N_1158,N_961,N_941);
and U1159 (N_1159,N_816,N_965);
and U1160 (N_1160,N_830,N_828);
nand U1161 (N_1161,N_898,N_910);
or U1162 (N_1162,N_958,N_999);
nor U1163 (N_1163,N_932,N_800);
xnor U1164 (N_1164,N_988,N_847);
and U1165 (N_1165,N_865,N_825);
and U1166 (N_1166,N_975,N_974);
nor U1167 (N_1167,N_994,N_849);
and U1168 (N_1168,N_859,N_972);
or U1169 (N_1169,N_819,N_987);
nor U1170 (N_1170,N_835,N_958);
nor U1171 (N_1171,N_954,N_915);
xor U1172 (N_1172,N_911,N_932);
or U1173 (N_1173,N_833,N_919);
nand U1174 (N_1174,N_931,N_923);
nor U1175 (N_1175,N_829,N_804);
nand U1176 (N_1176,N_989,N_884);
or U1177 (N_1177,N_992,N_972);
nand U1178 (N_1178,N_954,N_862);
nand U1179 (N_1179,N_843,N_955);
or U1180 (N_1180,N_836,N_893);
and U1181 (N_1181,N_834,N_997);
nand U1182 (N_1182,N_878,N_898);
nor U1183 (N_1183,N_882,N_961);
and U1184 (N_1184,N_847,N_800);
nor U1185 (N_1185,N_925,N_977);
or U1186 (N_1186,N_846,N_888);
and U1187 (N_1187,N_822,N_866);
and U1188 (N_1188,N_986,N_870);
nand U1189 (N_1189,N_953,N_922);
nor U1190 (N_1190,N_906,N_882);
and U1191 (N_1191,N_876,N_986);
nor U1192 (N_1192,N_996,N_839);
and U1193 (N_1193,N_896,N_875);
or U1194 (N_1194,N_877,N_939);
and U1195 (N_1195,N_836,N_832);
and U1196 (N_1196,N_999,N_869);
and U1197 (N_1197,N_952,N_914);
nor U1198 (N_1198,N_958,N_843);
nand U1199 (N_1199,N_892,N_882);
nor U1200 (N_1200,N_1056,N_1058);
xnor U1201 (N_1201,N_1031,N_1080);
nand U1202 (N_1202,N_1059,N_1015);
or U1203 (N_1203,N_1071,N_1074);
or U1204 (N_1204,N_1036,N_1060);
nand U1205 (N_1205,N_1155,N_1077);
or U1206 (N_1206,N_1005,N_1083);
and U1207 (N_1207,N_1079,N_1021);
nand U1208 (N_1208,N_1085,N_1142);
nand U1209 (N_1209,N_1160,N_1014);
nor U1210 (N_1210,N_1184,N_1019);
nor U1211 (N_1211,N_1001,N_1131);
nor U1212 (N_1212,N_1157,N_1076);
nor U1213 (N_1213,N_1165,N_1175);
or U1214 (N_1214,N_1087,N_1182);
and U1215 (N_1215,N_1010,N_1018);
nand U1216 (N_1216,N_1053,N_1129);
nor U1217 (N_1217,N_1061,N_1012);
nand U1218 (N_1218,N_1191,N_1063);
and U1219 (N_1219,N_1180,N_1123);
nand U1220 (N_1220,N_1064,N_1047);
nor U1221 (N_1221,N_1177,N_1172);
and U1222 (N_1222,N_1179,N_1150);
nor U1223 (N_1223,N_1037,N_1054);
or U1224 (N_1224,N_1032,N_1065);
nand U1225 (N_1225,N_1039,N_1190);
nand U1226 (N_1226,N_1072,N_1116);
nor U1227 (N_1227,N_1088,N_1057);
and U1228 (N_1228,N_1062,N_1133);
nand U1229 (N_1229,N_1183,N_1089);
nand U1230 (N_1230,N_1169,N_1096);
or U1231 (N_1231,N_1049,N_1055);
and U1232 (N_1232,N_1176,N_1112);
nor U1233 (N_1233,N_1187,N_1097);
or U1234 (N_1234,N_1107,N_1066);
nand U1235 (N_1235,N_1038,N_1126);
and U1236 (N_1236,N_1178,N_1025);
or U1237 (N_1237,N_1004,N_1051);
nor U1238 (N_1238,N_1167,N_1152);
nand U1239 (N_1239,N_1048,N_1104);
nand U1240 (N_1240,N_1171,N_1111);
and U1241 (N_1241,N_1106,N_1029);
or U1242 (N_1242,N_1134,N_1026);
nand U1243 (N_1243,N_1086,N_1017);
nor U1244 (N_1244,N_1198,N_1090);
or U1245 (N_1245,N_1052,N_1113);
nand U1246 (N_1246,N_1078,N_1141);
nand U1247 (N_1247,N_1185,N_1007);
nor U1248 (N_1248,N_1144,N_1151);
nor U1249 (N_1249,N_1117,N_1122);
or U1250 (N_1250,N_1114,N_1003);
nand U1251 (N_1251,N_1110,N_1188);
nand U1252 (N_1252,N_1093,N_1068);
nand U1253 (N_1253,N_1154,N_1130);
nor U1254 (N_1254,N_1069,N_1011);
xor U1255 (N_1255,N_1162,N_1043);
and U1256 (N_1256,N_1098,N_1164);
nand U1257 (N_1257,N_1101,N_1070);
and U1258 (N_1258,N_1092,N_1199);
nand U1259 (N_1259,N_1121,N_1000);
and U1260 (N_1260,N_1148,N_1149);
nand U1261 (N_1261,N_1020,N_1163);
and U1262 (N_1262,N_1067,N_1091);
or U1263 (N_1263,N_1196,N_1094);
and U1264 (N_1264,N_1103,N_1042);
nor U1265 (N_1265,N_1136,N_1009);
or U1266 (N_1266,N_1181,N_1194);
nand U1267 (N_1267,N_1034,N_1033);
nand U1268 (N_1268,N_1044,N_1195);
nand U1269 (N_1269,N_1041,N_1138);
nand U1270 (N_1270,N_1016,N_1105);
or U1271 (N_1271,N_1146,N_1173);
nor U1272 (N_1272,N_1099,N_1013);
nor U1273 (N_1273,N_1045,N_1166);
nand U1274 (N_1274,N_1028,N_1027);
and U1275 (N_1275,N_1161,N_1158);
nor U1276 (N_1276,N_1073,N_1137);
nor U1277 (N_1277,N_1170,N_1002);
nand U1278 (N_1278,N_1125,N_1118);
or U1279 (N_1279,N_1168,N_1006);
or U1280 (N_1280,N_1147,N_1082);
nand U1281 (N_1281,N_1174,N_1145);
or U1282 (N_1282,N_1030,N_1102);
nand U1283 (N_1283,N_1139,N_1120);
nand U1284 (N_1284,N_1075,N_1197);
nor U1285 (N_1285,N_1100,N_1008);
and U1286 (N_1286,N_1040,N_1193);
and U1287 (N_1287,N_1192,N_1095);
nor U1288 (N_1288,N_1108,N_1084);
nand U1289 (N_1289,N_1132,N_1128);
nand U1290 (N_1290,N_1081,N_1022);
nor U1291 (N_1291,N_1035,N_1050);
or U1292 (N_1292,N_1140,N_1156);
or U1293 (N_1293,N_1124,N_1046);
nand U1294 (N_1294,N_1024,N_1153);
nand U1295 (N_1295,N_1159,N_1119);
or U1296 (N_1296,N_1109,N_1186);
or U1297 (N_1297,N_1023,N_1143);
nor U1298 (N_1298,N_1127,N_1115);
nand U1299 (N_1299,N_1135,N_1189);
nand U1300 (N_1300,N_1085,N_1021);
or U1301 (N_1301,N_1133,N_1188);
xor U1302 (N_1302,N_1086,N_1194);
or U1303 (N_1303,N_1170,N_1024);
or U1304 (N_1304,N_1032,N_1176);
and U1305 (N_1305,N_1065,N_1117);
nor U1306 (N_1306,N_1194,N_1134);
and U1307 (N_1307,N_1114,N_1130);
nor U1308 (N_1308,N_1035,N_1048);
or U1309 (N_1309,N_1056,N_1136);
nor U1310 (N_1310,N_1048,N_1011);
nor U1311 (N_1311,N_1120,N_1100);
or U1312 (N_1312,N_1004,N_1049);
nand U1313 (N_1313,N_1192,N_1005);
nor U1314 (N_1314,N_1160,N_1172);
nand U1315 (N_1315,N_1092,N_1046);
nand U1316 (N_1316,N_1141,N_1003);
nor U1317 (N_1317,N_1087,N_1077);
xor U1318 (N_1318,N_1012,N_1022);
and U1319 (N_1319,N_1113,N_1015);
nand U1320 (N_1320,N_1089,N_1068);
nor U1321 (N_1321,N_1135,N_1127);
or U1322 (N_1322,N_1139,N_1104);
or U1323 (N_1323,N_1026,N_1087);
nand U1324 (N_1324,N_1049,N_1148);
nor U1325 (N_1325,N_1069,N_1020);
nand U1326 (N_1326,N_1044,N_1087);
or U1327 (N_1327,N_1001,N_1082);
or U1328 (N_1328,N_1107,N_1135);
nor U1329 (N_1329,N_1147,N_1189);
or U1330 (N_1330,N_1014,N_1021);
nand U1331 (N_1331,N_1175,N_1094);
and U1332 (N_1332,N_1117,N_1093);
and U1333 (N_1333,N_1150,N_1151);
or U1334 (N_1334,N_1116,N_1097);
nor U1335 (N_1335,N_1069,N_1063);
nand U1336 (N_1336,N_1140,N_1193);
nand U1337 (N_1337,N_1070,N_1000);
or U1338 (N_1338,N_1177,N_1051);
nor U1339 (N_1339,N_1043,N_1064);
nor U1340 (N_1340,N_1121,N_1012);
nand U1341 (N_1341,N_1013,N_1088);
nand U1342 (N_1342,N_1058,N_1068);
nand U1343 (N_1343,N_1048,N_1056);
nand U1344 (N_1344,N_1084,N_1058);
nand U1345 (N_1345,N_1072,N_1085);
nor U1346 (N_1346,N_1057,N_1059);
and U1347 (N_1347,N_1140,N_1104);
nand U1348 (N_1348,N_1176,N_1169);
or U1349 (N_1349,N_1084,N_1099);
or U1350 (N_1350,N_1135,N_1059);
nand U1351 (N_1351,N_1070,N_1088);
and U1352 (N_1352,N_1011,N_1087);
or U1353 (N_1353,N_1022,N_1052);
xnor U1354 (N_1354,N_1027,N_1038);
nor U1355 (N_1355,N_1028,N_1142);
nand U1356 (N_1356,N_1069,N_1031);
nor U1357 (N_1357,N_1144,N_1089);
or U1358 (N_1358,N_1078,N_1119);
and U1359 (N_1359,N_1154,N_1095);
or U1360 (N_1360,N_1057,N_1022);
nand U1361 (N_1361,N_1028,N_1191);
nor U1362 (N_1362,N_1042,N_1078);
nand U1363 (N_1363,N_1025,N_1003);
and U1364 (N_1364,N_1158,N_1132);
and U1365 (N_1365,N_1127,N_1092);
and U1366 (N_1366,N_1104,N_1022);
and U1367 (N_1367,N_1118,N_1183);
and U1368 (N_1368,N_1153,N_1165);
nor U1369 (N_1369,N_1056,N_1000);
and U1370 (N_1370,N_1152,N_1017);
or U1371 (N_1371,N_1105,N_1140);
nand U1372 (N_1372,N_1184,N_1160);
and U1373 (N_1373,N_1096,N_1165);
nand U1374 (N_1374,N_1157,N_1162);
nand U1375 (N_1375,N_1165,N_1058);
nand U1376 (N_1376,N_1056,N_1123);
and U1377 (N_1377,N_1130,N_1004);
or U1378 (N_1378,N_1173,N_1137);
and U1379 (N_1379,N_1037,N_1140);
nand U1380 (N_1380,N_1076,N_1119);
and U1381 (N_1381,N_1128,N_1068);
or U1382 (N_1382,N_1122,N_1076);
nand U1383 (N_1383,N_1084,N_1090);
or U1384 (N_1384,N_1107,N_1100);
and U1385 (N_1385,N_1081,N_1056);
nand U1386 (N_1386,N_1154,N_1034);
or U1387 (N_1387,N_1036,N_1015);
xnor U1388 (N_1388,N_1014,N_1072);
nor U1389 (N_1389,N_1006,N_1046);
or U1390 (N_1390,N_1142,N_1011);
or U1391 (N_1391,N_1060,N_1173);
or U1392 (N_1392,N_1058,N_1149);
or U1393 (N_1393,N_1045,N_1176);
nor U1394 (N_1394,N_1012,N_1078);
nor U1395 (N_1395,N_1029,N_1105);
nor U1396 (N_1396,N_1045,N_1123);
and U1397 (N_1397,N_1045,N_1162);
nand U1398 (N_1398,N_1159,N_1046);
xnor U1399 (N_1399,N_1198,N_1142);
nor U1400 (N_1400,N_1330,N_1353);
or U1401 (N_1401,N_1216,N_1282);
and U1402 (N_1402,N_1385,N_1305);
nand U1403 (N_1403,N_1272,N_1296);
and U1404 (N_1404,N_1284,N_1292);
and U1405 (N_1405,N_1271,N_1313);
nand U1406 (N_1406,N_1234,N_1246);
nand U1407 (N_1407,N_1396,N_1325);
nand U1408 (N_1408,N_1295,N_1302);
nor U1409 (N_1409,N_1386,N_1338);
nand U1410 (N_1410,N_1254,N_1274);
nor U1411 (N_1411,N_1339,N_1291);
nor U1412 (N_1412,N_1280,N_1281);
nand U1413 (N_1413,N_1245,N_1208);
nand U1414 (N_1414,N_1279,N_1275);
or U1415 (N_1415,N_1345,N_1357);
nand U1416 (N_1416,N_1373,N_1365);
and U1417 (N_1417,N_1362,N_1389);
nand U1418 (N_1418,N_1321,N_1209);
and U1419 (N_1419,N_1372,N_1287);
nand U1420 (N_1420,N_1260,N_1202);
xnor U1421 (N_1421,N_1348,N_1257);
nand U1422 (N_1422,N_1381,N_1203);
nand U1423 (N_1423,N_1212,N_1352);
or U1424 (N_1424,N_1300,N_1326);
nor U1425 (N_1425,N_1363,N_1374);
or U1426 (N_1426,N_1344,N_1200);
nor U1427 (N_1427,N_1244,N_1359);
nor U1428 (N_1428,N_1239,N_1355);
or U1429 (N_1429,N_1301,N_1205);
and U1430 (N_1430,N_1343,N_1368);
nor U1431 (N_1431,N_1380,N_1384);
nand U1432 (N_1432,N_1224,N_1327);
nor U1433 (N_1433,N_1371,N_1306);
or U1434 (N_1434,N_1298,N_1351);
nand U1435 (N_1435,N_1304,N_1247);
or U1436 (N_1436,N_1370,N_1337);
nand U1437 (N_1437,N_1248,N_1236);
and U1438 (N_1438,N_1349,N_1207);
and U1439 (N_1439,N_1297,N_1223);
nand U1440 (N_1440,N_1261,N_1204);
or U1441 (N_1441,N_1273,N_1394);
nand U1442 (N_1442,N_1294,N_1311);
nand U1443 (N_1443,N_1342,N_1308);
nor U1444 (N_1444,N_1331,N_1328);
nand U1445 (N_1445,N_1390,N_1232);
or U1446 (N_1446,N_1219,N_1316);
and U1447 (N_1447,N_1268,N_1379);
and U1448 (N_1448,N_1387,N_1354);
and U1449 (N_1449,N_1356,N_1332);
or U1450 (N_1450,N_1392,N_1315);
and U1451 (N_1451,N_1270,N_1231);
nand U1452 (N_1452,N_1206,N_1350);
nand U1453 (N_1453,N_1347,N_1312);
and U1454 (N_1454,N_1201,N_1217);
or U1455 (N_1455,N_1259,N_1210);
nor U1456 (N_1456,N_1240,N_1366);
or U1457 (N_1457,N_1263,N_1251);
nand U1458 (N_1458,N_1375,N_1382);
nor U1459 (N_1459,N_1220,N_1269);
nand U1460 (N_1460,N_1388,N_1237);
or U1461 (N_1461,N_1230,N_1293);
nand U1462 (N_1462,N_1395,N_1225);
and U1463 (N_1463,N_1299,N_1360);
nor U1464 (N_1464,N_1277,N_1253);
or U1465 (N_1465,N_1314,N_1285);
or U1466 (N_1466,N_1226,N_1391);
nand U1467 (N_1467,N_1318,N_1229);
nand U1468 (N_1468,N_1341,N_1399);
and U1469 (N_1469,N_1317,N_1358);
or U1470 (N_1470,N_1369,N_1264);
nor U1471 (N_1471,N_1323,N_1278);
nand U1472 (N_1472,N_1265,N_1276);
nand U1473 (N_1473,N_1227,N_1290);
and U1474 (N_1474,N_1233,N_1393);
and U1475 (N_1475,N_1242,N_1250);
nand U1476 (N_1476,N_1333,N_1266);
and U1477 (N_1477,N_1286,N_1340);
or U1478 (N_1478,N_1252,N_1310);
or U1479 (N_1479,N_1364,N_1221);
or U1480 (N_1480,N_1256,N_1213);
or U1481 (N_1481,N_1329,N_1335);
nand U1482 (N_1482,N_1255,N_1322);
and U1483 (N_1483,N_1235,N_1309);
or U1484 (N_1484,N_1378,N_1267);
and U1485 (N_1485,N_1346,N_1218);
nor U1486 (N_1486,N_1319,N_1303);
nand U1487 (N_1487,N_1249,N_1361);
and U1488 (N_1488,N_1367,N_1289);
nor U1489 (N_1489,N_1238,N_1336);
nand U1490 (N_1490,N_1241,N_1397);
nand U1491 (N_1491,N_1243,N_1215);
and U1492 (N_1492,N_1283,N_1258);
or U1493 (N_1493,N_1398,N_1228);
nor U1494 (N_1494,N_1262,N_1334);
nor U1495 (N_1495,N_1307,N_1288);
or U1496 (N_1496,N_1214,N_1320);
or U1497 (N_1497,N_1376,N_1211);
or U1498 (N_1498,N_1222,N_1383);
nand U1499 (N_1499,N_1377,N_1324);
or U1500 (N_1500,N_1358,N_1279);
nor U1501 (N_1501,N_1356,N_1350);
nor U1502 (N_1502,N_1321,N_1330);
nand U1503 (N_1503,N_1249,N_1325);
nor U1504 (N_1504,N_1235,N_1306);
nor U1505 (N_1505,N_1329,N_1241);
and U1506 (N_1506,N_1210,N_1241);
nand U1507 (N_1507,N_1354,N_1218);
nor U1508 (N_1508,N_1238,N_1319);
or U1509 (N_1509,N_1218,N_1361);
or U1510 (N_1510,N_1290,N_1278);
nand U1511 (N_1511,N_1336,N_1235);
xor U1512 (N_1512,N_1399,N_1212);
nand U1513 (N_1513,N_1345,N_1298);
nor U1514 (N_1514,N_1265,N_1211);
or U1515 (N_1515,N_1306,N_1355);
nand U1516 (N_1516,N_1204,N_1377);
and U1517 (N_1517,N_1333,N_1397);
and U1518 (N_1518,N_1256,N_1350);
nor U1519 (N_1519,N_1319,N_1217);
nand U1520 (N_1520,N_1363,N_1351);
nor U1521 (N_1521,N_1378,N_1335);
nand U1522 (N_1522,N_1346,N_1294);
or U1523 (N_1523,N_1228,N_1347);
nor U1524 (N_1524,N_1274,N_1219);
xor U1525 (N_1525,N_1279,N_1219);
or U1526 (N_1526,N_1216,N_1327);
xnor U1527 (N_1527,N_1306,N_1263);
nor U1528 (N_1528,N_1359,N_1376);
nor U1529 (N_1529,N_1260,N_1327);
nor U1530 (N_1530,N_1377,N_1323);
nand U1531 (N_1531,N_1301,N_1231);
nor U1532 (N_1532,N_1382,N_1388);
nor U1533 (N_1533,N_1203,N_1262);
or U1534 (N_1534,N_1238,N_1327);
and U1535 (N_1535,N_1260,N_1287);
nand U1536 (N_1536,N_1248,N_1330);
or U1537 (N_1537,N_1317,N_1335);
or U1538 (N_1538,N_1369,N_1383);
or U1539 (N_1539,N_1348,N_1223);
nor U1540 (N_1540,N_1302,N_1373);
or U1541 (N_1541,N_1336,N_1399);
nand U1542 (N_1542,N_1319,N_1317);
or U1543 (N_1543,N_1368,N_1208);
or U1544 (N_1544,N_1389,N_1275);
or U1545 (N_1545,N_1274,N_1351);
or U1546 (N_1546,N_1374,N_1269);
nor U1547 (N_1547,N_1271,N_1212);
nand U1548 (N_1548,N_1346,N_1245);
nand U1549 (N_1549,N_1219,N_1363);
nand U1550 (N_1550,N_1206,N_1393);
nor U1551 (N_1551,N_1332,N_1359);
nor U1552 (N_1552,N_1210,N_1224);
and U1553 (N_1553,N_1292,N_1235);
nand U1554 (N_1554,N_1376,N_1321);
nor U1555 (N_1555,N_1360,N_1241);
and U1556 (N_1556,N_1391,N_1279);
nor U1557 (N_1557,N_1383,N_1396);
and U1558 (N_1558,N_1344,N_1370);
nor U1559 (N_1559,N_1307,N_1215);
nor U1560 (N_1560,N_1275,N_1218);
nand U1561 (N_1561,N_1293,N_1326);
or U1562 (N_1562,N_1316,N_1237);
or U1563 (N_1563,N_1265,N_1305);
nor U1564 (N_1564,N_1399,N_1218);
xnor U1565 (N_1565,N_1292,N_1206);
nand U1566 (N_1566,N_1344,N_1254);
and U1567 (N_1567,N_1376,N_1365);
nand U1568 (N_1568,N_1322,N_1315);
nand U1569 (N_1569,N_1322,N_1264);
or U1570 (N_1570,N_1392,N_1384);
and U1571 (N_1571,N_1350,N_1359);
nand U1572 (N_1572,N_1386,N_1251);
nand U1573 (N_1573,N_1385,N_1356);
nor U1574 (N_1574,N_1370,N_1207);
nor U1575 (N_1575,N_1365,N_1338);
or U1576 (N_1576,N_1328,N_1325);
and U1577 (N_1577,N_1335,N_1214);
and U1578 (N_1578,N_1318,N_1203);
nor U1579 (N_1579,N_1267,N_1242);
nand U1580 (N_1580,N_1274,N_1347);
nor U1581 (N_1581,N_1357,N_1389);
or U1582 (N_1582,N_1242,N_1362);
or U1583 (N_1583,N_1301,N_1381);
and U1584 (N_1584,N_1294,N_1239);
and U1585 (N_1585,N_1390,N_1316);
and U1586 (N_1586,N_1240,N_1309);
nor U1587 (N_1587,N_1297,N_1259);
or U1588 (N_1588,N_1239,N_1226);
nand U1589 (N_1589,N_1217,N_1374);
or U1590 (N_1590,N_1234,N_1274);
or U1591 (N_1591,N_1325,N_1296);
nor U1592 (N_1592,N_1347,N_1208);
nand U1593 (N_1593,N_1316,N_1322);
or U1594 (N_1594,N_1284,N_1364);
nand U1595 (N_1595,N_1313,N_1312);
and U1596 (N_1596,N_1251,N_1378);
xor U1597 (N_1597,N_1335,N_1392);
xor U1598 (N_1598,N_1320,N_1366);
or U1599 (N_1599,N_1283,N_1371);
and U1600 (N_1600,N_1594,N_1422);
nor U1601 (N_1601,N_1468,N_1406);
nand U1602 (N_1602,N_1407,N_1556);
nand U1603 (N_1603,N_1444,N_1587);
or U1604 (N_1604,N_1501,N_1533);
nand U1605 (N_1605,N_1483,N_1534);
or U1606 (N_1606,N_1452,N_1549);
nand U1607 (N_1607,N_1548,N_1436);
and U1608 (N_1608,N_1428,N_1405);
or U1609 (N_1609,N_1460,N_1409);
nand U1610 (N_1610,N_1448,N_1511);
and U1611 (N_1611,N_1562,N_1583);
and U1612 (N_1612,N_1521,N_1536);
nor U1613 (N_1613,N_1506,N_1507);
or U1614 (N_1614,N_1478,N_1596);
nor U1615 (N_1615,N_1535,N_1429);
nand U1616 (N_1616,N_1426,N_1504);
or U1617 (N_1617,N_1545,N_1408);
nand U1618 (N_1618,N_1414,N_1411);
and U1619 (N_1619,N_1563,N_1427);
and U1620 (N_1620,N_1580,N_1463);
or U1621 (N_1621,N_1592,N_1480);
nor U1622 (N_1622,N_1418,N_1443);
nor U1623 (N_1623,N_1514,N_1567);
nand U1624 (N_1624,N_1569,N_1518);
and U1625 (N_1625,N_1470,N_1430);
nor U1626 (N_1626,N_1477,N_1599);
nand U1627 (N_1627,N_1525,N_1502);
xnor U1628 (N_1628,N_1522,N_1449);
and U1629 (N_1629,N_1447,N_1571);
nand U1630 (N_1630,N_1403,N_1459);
and U1631 (N_1631,N_1494,N_1446);
nand U1632 (N_1632,N_1473,N_1462);
nand U1633 (N_1633,N_1584,N_1552);
nor U1634 (N_1634,N_1519,N_1465);
and U1635 (N_1635,N_1503,N_1538);
nand U1636 (N_1636,N_1526,N_1438);
nor U1637 (N_1637,N_1581,N_1445);
nand U1638 (N_1638,N_1486,N_1410);
nand U1639 (N_1639,N_1566,N_1516);
or U1640 (N_1640,N_1453,N_1475);
nor U1641 (N_1641,N_1543,N_1528);
nor U1642 (N_1642,N_1439,N_1493);
nand U1643 (N_1643,N_1597,N_1554);
or U1644 (N_1644,N_1472,N_1544);
or U1645 (N_1645,N_1487,N_1496);
nand U1646 (N_1646,N_1455,N_1454);
nand U1647 (N_1647,N_1512,N_1450);
or U1648 (N_1648,N_1495,N_1404);
and U1649 (N_1649,N_1458,N_1591);
nor U1650 (N_1650,N_1442,N_1529);
and U1651 (N_1651,N_1433,N_1542);
nor U1652 (N_1652,N_1489,N_1540);
and U1653 (N_1653,N_1457,N_1451);
nor U1654 (N_1654,N_1421,N_1479);
nor U1655 (N_1655,N_1456,N_1579);
or U1656 (N_1656,N_1417,N_1537);
and U1657 (N_1657,N_1508,N_1467);
or U1658 (N_1658,N_1550,N_1440);
nor U1659 (N_1659,N_1432,N_1485);
or U1660 (N_1660,N_1484,N_1531);
nand U1661 (N_1661,N_1585,N_1499);
nor U1662 (N_1662,N_1578,N_1574);
and U1663 (N_1663,N_1568,N_1573);
nand U1664 (N_1664,N_1488,N_1590);
and U1665 (N_1665,N_1497,N_1572);
or U1666 (N_1666,N_1476,N_1505);
or U1667 (N_1667,N_1500,N_1523);
nor U1668 (N_1668,N_1415,N_1491);
or U1669 (N_1669,N_1586,N_1598);
nand U1670 (N_1670,N_1419,N_1510);
nor U1671 (N_1671,N_1423,N_1588);
or U1672 (N_1672,N_1595,N_1547);
and U1673 (N_1673,N_1435,N_1541);
and U1674 (N_1674,N_1520,N_1461);
nor U1675 (N_1675,N_1492,N_1402);
and U1676 (N_1676,N_1471,N_1559);
or U1677 (N_1677,N_1431,N_1555);
or U1678 (N_1678,N_1413,N_1582);
and U1679 (N_1679,N_1441,N_1412);
xnor U1680 (N_1680,N_1551,N_1524);
and U1681 (N_1681,N_1560,N_1424);
nand U1682 (N_1682,N_1437,N_1401);
nand U1683 (N_1683,N_1490,N_1466);
or U1684 (N_1684,N_1515,N_1530);
nand U1685 (N_1685,N_1575,N_1589);
nor U1686 (N_1686,N_1481,N_1558);
nand U1687 (N_1687,N_1416,N_1420);
nand U1688 (N_1688,N_1577,N_1464);
nor U1689 (N_1689,N_1469,N_1517);
and U1690 (N_1690,N_1498,N_1434);
and U1691 (N_1691,N_1576,N_1593);
nand U1692 (N_1692,N_1527,N_1482);
or U1693 (N_1693,N_1565,N_1539);
or U1694 (N_1694,N_1553,N_1400);
or U1695 (N_1695,N_1532,N_1425);
nor U1696 (N_1696,N_1513,N_1564);
nand U1697 (N_1697,N_1474,N_1509);
nor U1698 (N_1698,N_1570,N_1561);
nor U1699 (N_1699,N_1546,N_1557);
and U1700 (N_1700,N_1568,N_1496);
nor U1701 (N_1701,N_1500,N_1504);
and U1702 (N_1702,N_1574,N_1409);
nor U1703 (N_1703,N_1590,N_1581);
nor U1704 (N_1704,N_1594,N_1513);
nand U1705 (N_1705,N_1437,N_1531);
nor U1706 (N_1706,N_1409,N_1454);
nor U1707 (N_1707,N_1491,N_1414);
or U1708 (N_1708,N_1425,N_1534);
nand U1709 (N_1709,N_1437,N_1509);
nor U1710 (N_1710,N_1542,N_1506);
and U1711 (N_1711,N_1577,N_1499);
or U1712 (N_1712,N_1436,N_1537);
nand U1713 (N_1713,N_1479,N_1457);
nand U1714 (N_1714,N_1473,N_1584);
and U1715 (N_1715,N_1448,N_1431);
nand U1716 (N_1716,N_1427,N_1532);
or U1717 (N_1717,N_1572,N_1527);
nand U1718 (N_1718,N_1586,N_1454);
nor U1719 (N_1719,N_1564,N_1549);
and U1720 (N_1720,N_1465,N_1406);
nor U1721 (N_1721,N_1590,N_1532);
nand U1722 (N_1722,N_1514,N_1495);
or U1723 (N_1723,N_1462,N_1438);
or U1724 (N_1724,N_1486,N_1542);
nor U1725 (N_1725,N_1454,N_1482);
xnor U1726 (N_1726,N_1442,N_1451);
nand U1727 (N_1727,N_1401,N_1571);
and U1728 (N_1728,N_1464,N_1465);
nor U1729 (N_1729,N_1419,N_1516);
nor U1730 (N_1730,N_1435,N_1462);
nor U1731 (N_1731,N_1402,N_1406);
nand U1732 (N_1732,N_1422,N_1553);
and U1733 (N_1733,N_1409,N_1513);
nand U1734 (N_1734,N_1475,N_1482);
nand U1735 (N_1735,N_1510,N_1407);
and U1736 (N_1736,N_1567,N_1507);
nand U1737 (N_1737,N_1530,N_1580);
nor U1738 (N_1738,N_1545,N_1504);
and U1739 (N_1739,N_1486,N_1557);
and U1740 (N_1740,N_1413,N_1471);
and U1741 (N_1741,N_1477,N_1592);
nor U1742 (N_1742,N_1524,N_1560);
nand U1743 (N_1743,N_1473,N_1528);
or U1744 (N_1744,N_1549,N_1463);
nor U1745 (N_1745,N_1419,N_1426);
and U1746 (N_1746,N_1556,N_1421);
or U1747 (N_1747,N_1458,N_1432);
nand U1748 (N_1748,N_1535,N_1469);
nand U1749 (N_1749,N_1490,N_1444);
nand U1750 (N_1750,N_1436,N_1577);
nor U1751 (N_1751,N_1537,N_1420);
and U1752 (N_1752,N_1551,N_1437);
or U1753 (N_1753,N_1551,N_1536);
nand U1754 (N_1754,N_1521,N_1484);
nor U1755 (N_1755,N_1467,N_1547);
nor U1756 (N_1756,N_1466,N_1421);
or U1757 (N_1757,N_1597,N_1489);
nor U1758 (N_1758,N_1457,N_1493);
or U1759 (N_1759,N_1478,N_1502);
or U1760 (N_1760,N_1430,N_1551);
and U1761 (N_1761,N_1544,N_1447);
and U1762 (N_1762,N_1442,N_1432);
xor U1763 (N_1763,N_1411,N_1409);
nand U1764 (N_1764,N_1492,N_1585);
or U1765 (N_1765,N_1415,N_1439);
or U1766 (N_1766,N_1516,N_1486);
and U1767 (N_1767,N_1498,N_1505);
nor U1768 (N_1768,N_1430,N_1563);
nand U1769 (N_1769,N_1550,N_1549);
or U1770 (N_1770,N_1483,N_1406);
nand U1771 (N_1771,N_1466,N_1474);
or U1772 (N_1772,N_1582,N_1487);
nand U1773 (N_1773,N_1411,N_1487);
xnor U1774 (N_1774,N_1510,N_1526);
or U1775 (N_1775,N_1497,N_1415);
nand U1776 (N_1776,N_1534,N_1504);
or U1777 (N_1777,N_1592,N_1530);
or U1778 (N_1778,N_1453,N_1432);
nor U1779 (N_1779,N_1434,N_1499);
nor U1780 (N_1780,N_1410,N_1472);
and U1781 (N_1781,N_1567,N_1456);
and U1782 (N_1782,N_1525,N_1413);
nand U1783 (N_1783,N_1449,N_1466);
nor U1784 (N_1784,N_1444,N_1424);
or U1785 (N_1785,N_1514,N_1560);
nand U1786 (N_1786,N_1570,N_1494);
nor U1787 (N_1787,N_1407,N_1557);
or U1788 (N_1788,N_1518,N_1536);
nor U1789 (N_1789,N_1468,N_1478);
nand U1790 (N_1790,N_1508,N_1591);
or U1791 (N_1791,N_1504,N_1419);
nand U1792 (N_1792,N_1406,N_1446);
nor U1793 (N_1793,N_1547,N_1445);
nor U1794 (N_1794,N_1594,N_1434);
and U1795 (N_1795,N_1517,N_1443);
or U1796 (N_1796,N_1496,N_1411);
or U1797 (N_1797,N_1498,N_1534);
nor U1798 (N_1798,N_1432,N_1477);
nand U1799 (N_1799,N_1451,N_1454);
and U1800 (N_1800,N_1648,N_1735);
nand U1801 (N_1801,N_1782,N_1651);
and U1802 (N_1802,N_1681,N_1606);
nor U1803 (N_1803,N_1750,N_1660);
nor U1804 (N_1804,N_1783,N_1751);
or U1805 (N_1805,N_1694,N_1717);
and U1806 (N_1806,N_1766,N_1642);
nand U1807 (N_1807,N_1776,N_1673);
or U1808 (N_1808,N_1640,N_1778);
nand U1809 (N_1809,N_1798,N_1628);
and U1810 (N_1810,N_1637,N_1763);
and U1811 (N_1811,N_1720,N_1710);
nor U1812 (N_1812,N_1629,N_1609);
and U1813 (N_1813,N_1711,N_1746);
or U1814 (N_1814,N_1713,N_1686);
nand U1815 (N_1815,N_1755,N_1659);
and U1816 (N_1816,N_1761,N_1610);
nand U1817 (N_1817,N_1754,N_1608);
or U1818 (N_1818,N_1740,N_1669);
nor U1819 (N_1819,N_1601,N_1605);
or U1820 (N_1820,N_1718,N_1616);
or U1821 (N_1821,N_1725,N_1726);
or U1822 (N_1822,N_1768,N_1736);
and U1823 (N_1823,N_1715,N_1724);
nand U1824 (N_1824,N_1636,N_1621);
nand U1825 (N_1825,N_1787,N_1773);
nand U1826 (N_1826,N_1602,N_1742);
and U1827 (N_1827,N_1641,N_1622);
and U1828 (N_1828,N_1721,N_1714);
nor U1829 (N_1829,N_1771,N_1646);
nand U1830 (N_1830,N_1632,N_1655);
nand U1831 (N_1831,N_1770,N_1623);
and U1832 (N_1832,N_1685,N_1625);
nor U1833 (N_1833,N_1614,N_1767);
nand U1834 (N_1834,N_1745,N_1676);
nand U1835 (N_1835,N_1774,N_1775);
nor U1836 (N_1836,N_1760,N_1657);
and U1837 (N_1837,N_1696,N_1674);
nor U1838 (N_1838,N_1688,N_1730);
and U1839 (N_1839,N_1789,N_1650);
or U1840 (N_1840,N_1667,N_1679);
nor U1841 (N_1841,N_1607,N_1683);
or U1842 (N_1842,N_1678,N_1691);
and U1843 (N_1843,N_1693,N_1633);
and U1844 (N_1844,N_1635,N_1727);
and U1845 (N_1845,N_1743,N_1682);
nand U1846 (N_1846,N_1748,N_1744);
and U1847 (N_1847,N_1604,N_1627);
or U1848 (N_1848,N_1747,N_1695);
nand U1849 (N_1849,N_1684,N_1731);
nor U1850 (N_1850,N_1662,N_1664);
nand U1851 (N_1851,N_1799,N_1618);
and U1852 (N_1852,N_1764,N_1779);
nor U1853 (N_1853,N_1709,N_1665);
and U1854 (N_1854,N_1677,N_1753);
nor U1855 (N_1855,N_1707,N_1643);
and U1856 (N_1856,N_1708,N_1663);
nor U1857 (N_1857,N_1781,N_1794);
or U1858 (N_1858,N_1670,N_1791);
and U1859 (N_1859,N_1716,N_1759);
nand U1860 (N_1860,N_1793,N_1697);
or U1861 (N_1861,N_1666,N_1672);
or U1862 (N_1862,N_1668,N_1790);
nand U1863 (N_1863,N_1706,N_1723);
nor U1864 (N_1864,N_1712,N_1784);
nor U1865 (N_1865,N_1700,N_1728);
nand U1866 (N_1866,N_1741,N_1644);
nor U1867 (N_1867,N_1719,N_1645);
nor U1868 (N_1868,N_1757,N_1613);
nor U1869 (N_1869,N_1603,N_1653);
and U1870 (N_1870,N_1654,N_1630);
or U1871 (N_1871,N_1611,N_1617);
and U1872 (N_1872,N_1756,N_1738);
xnor U1873 (N_1873,N_1704,N_1658);
nand U1874 (N_1874,N_1649,N_1739);
or U1875 (N_1875,N_1634,N_1772);
or U1876 (N_1876,N_1675,N_1661);
xnor U1877 (N_1877,N_1796,N_1626);
and U1878 (N_1878,N_1687,N_1758);
and U1879 (N_1879,N_1702,N_1689);
nor U1880 (N_1880,N_1647,N_1797);
and U1881 (N_1881,N_1734,N_1752);
and U1882 (N_1882,N_1698,N_1732);
nand U1883 (N_1883,N_1786,N_1788);
nand U1884 (N_1884,N_1639,N_1624);
and U1885 (N_1885,N_1703,N_1722);
or U1886 (N_1886,N_1705,N_1762);
nor U1887 (N_1887,N_1690,N_1612);
or U1888 (N_1888,N_1769,N_1600);
nand U1889 (N_1889,N_1671,N_1729);
nand U1890 (N_1890,N_1699,N_1638);
nor U1891 (N_1891,N_1785,N_1692);
nor U1892 (N_1892,N_1620,N_1701);
and U1893 (N_1893,N_1652,N_1656);
nand U1894 (N_1894,N_1777,N_1749);
or U1895 (N_1895,N_1765,N_1615);
nand U1896 (N_1896,N_1680,N_1792);
nand U1897 (N_1897,N_1795,N_1619);
nand U1898 (N_1898,N_1631,N_1780);
and U1899 (N_1899,N_1737,N_1733);
and U1900 (N_1900,N_1705,N_1607);
or U1901 (N_1901,N_1621,N_1788);
nand U1902 (N_1902,N_1677,N_1652);
or U1903 (N_1903,N_1747,N_1604);
nor U1904 (N_1904,N_1781,N_1640);
xor U1905 (N_1905,N_1656,N_1645);
xor U1906 (N_1906,N_1714,N_1733);
nand U1907 (N_1907,N_1612,N_1609);
nand U1908 (N_1908,N_1722,N_1756);
nor U1909 (N_1909,N_1797,N_1747);
and U1910 (N_1910,N_1740,N_1750);
nor U1911 (N_1911,N_1747,N_1726);
or U1912 (N_1912,N_1754,N_1669);
nor U1913 (N_1913,N_1716,N_1681);
nand U1914 (N_1914,N_1635,N_1726);
or U1915 (N_1915,N_1794,N_1633);
nor U1916 (N_1916,N_1619,N_1623);
or U1917 (N_1917,N_1619,N_1732);
and U1918 (N_1918,N_1631,N_1758);
or U1919 (N_1919,N_1779,N_1725);
nand U1920 (N_1920,N_1710,N_1775);
nand U1921 (N_1921,N_1600,N_1603);
or U1922 (N_1922,N_1724,N_1654);
or U1923 (N_1923,N_1634,N_1684);
and U1924 (N_1924,N_1740,N_1736);
and U1925 (N_1925,N_1676,N_1689);
and U1926 (N_1926,N_1726,N_1698);
nor U1927 (N_1927,N_1708,N_1729);
nor U1928 (N_1928,N_1745,N_1605);
or U1929 (N_1929,N_1724,N_1748);
and U1930 (N_1930,N_1767,N_1737);
nand U1931 (N_1931,N_1673,N_1625);
nor U1932 (N_1932,N_1789,N_1710);
nand U1933 (N_1933,N_1652,N_1660);
or U1934 (N_1934,N_1771,N_1724);
and U1935 (N_1935,N_1617,N_1781);
nor U1936 (N_1936,N_1745,N_1751);
nand U1937 (N_1937,N_1665,N_1755);
nand U1938 (N_1938,N_1653,N_1722);
or U1939 (N_1939,N_1782,N_1757);
and U1940 (N_1940,N_1746,N_1766);
nor U1941 (N_1941,N_1646,N_1679);
and U1942 (N_1942,N_1627,N_1798);
and U1943 (N_1943,N_1751,N_1688);
or U1944 (N_1944,N_1718,N_1609);
and U1945 (N_1945,N_1683,N_1796);
nor U1946 (N_1946,N_1602,N_1753);
or U1947 (N_1947,N_1658,N_1612);
nand U1948 (N_1948,N_1759,N_1664);
nor U1949 (N_1949,N_1718,N_1682);
nor U1950 (N_1950,N_1762,N_1649);
nor U1951 (N_1951,N_1711,N_1602);
and U1952 (N_1952,N_1603,N_1658);
nor U1953 (N_1953,N_1709,N_1671);
or U1954 (N_1954,N_1621,N_1782);
nand U1955 (N_1955,N_1646,N_1610);
nor U1956 (N_1956,N_1684,N_1686);
nand U1957 (N_1957,N_1787,N_1757);
and U1958 (N_1958,N_1744,N_1630);
or U1959 (N_1959,N_1688,N_1655);
nand U1960 (N_1960,N_1699,N_1631);
and U1961 (N_1961,N_1653,N_1627);
and U1962 (N_1962,N_1618,N_1623);
nor U1963 (N_1963,N_1704,N_1743);
nand U1964 (N_1964,N_1702,N_1725);
nor U1965 (N_1965,N_1606,N_1617);
and U1966 (N_1966,N_1777,N_1770);
and U1967 (N_1967,N_1617,N_1753);
nor U1968 (N_1968,N_1625,N_1732);
nand U1969 (N_1969,N_1667,N_1643);
and U1970 (N_1970,N_1759,N_1739);
nand U1971 (N_1971,N_1743,N_1702);
or U1972 (N_1972,N_1792,N_1645);
and U1973 (N_1973,N_1619,N_1798);
or U1974 (N_1974,N_1648,N_1740);
or U1975 (N_1975,N_1692,N_1666);
nand U1976 (N_1976,N_1738,N_1783);
nand U1977 (N_1977,N_1707,N_1717);
nand U1978 (N_1978,N_1740,N_1726);
and U1979 (N_1979,N_1678,N_1685);
and U1980 (N_1980,N_1695,N_1657);
nand U1981 (N_1981,N_1762,N_1621);
and U1982 (N_1982,N_1602,N_1601);
nand U1983 (N_1983,N_1754,N_1739);
or U1984 (N_1984,N_1600,N_1637);
and U1985 (N_1985,N_1663,N_1773);
xnor U1986 (N_1986,N_1791,N_1752);
nand U1987 (N_1987,N_1651,N_1622);
nor U1988 (N_1988,N_1782,N_1670);
and U1989 (N_1989,N_1710,N_1666);
and U1990 (N_1990,N_1643,N_1618);
and U1991 (N_1991,N_1732,N_1649);
and U1992 (N_1992,N_1660,N_1638);
nor U1993 (N_1993,N_1781,N_1765);
nand U1994 (N_1994,N_1624,N_1629);
nand U1995 (N_1995,N_1605,N_1775);
or U1996 (N_1996,N_1676,N_1713);
and U1997 (N_1997,N_1788,N_1791);
nor U1998 (N_1998,N_1649,N_1770);
xnor U1999 (N_1999,N_1766,N_1605);
nor U2000 (N_2000,N_1964,N_1945);
and U2001 (N_2001,N_1831,N_1887);
nor U2002 (N_2002,N_1873,N_1820);
nand U2003 (N_2003,N_1882,N_1978);
and U2004 (N_2004,N_1929,N_1846);
or U2005 (N_2005,N_1817,N_1934);
nor U2006 (N_2006,N_1813,N_1862);
and U2007 (N_2007,N_1879,N_1843);
nand U2008 (N_2008,N_1811,N_1832);
xor U2009 (N_2009,N_1953,N_1958);
nand U2010 (N_2010,N_1916,N_1860);
and U2011 (N_2011,N_1976,N_1957);
nand U2012 (N_2012,N_1968,N_1907);
nor U2013 (N_2013,N_1854,N_1823);
and U2014 (N_2014,N_1876,N_1858);
or U2015 (N_2015,N_1810,N_1919);
nand U2016 (N_2016,N_1963,N_1905);
xor U2017 (N_2017,N_1999,N_1926);
nor U2018 (N_2018,N_1954,N_1833);
nor U2019 (N_2019,N_1848,N_1972);
nor U2020 (N_2020,N_1912,N_1807);
nand U2021 (N_2021,N_1901,N_1900);
xnor U2022 (N_2022,N_1840,N_1949);
nand U2023 (N_2023,N_1917,N_1885);
nand U2024 (N_2024,N_1996,N_1986);
nor U2025 (N_2025,N_1921,N_1928);
nor U2026 (N_2026,N_1889,N_1877);
nand U2027 (N_2027,N_1801,N_1839);
xor U2028 (N_2028,N_1822,N_1899);
nor U2029 (N_2029,N_1850,N_1891);
and U2030 (N_2030,N_1966,N_1909);
or U2031 (N_2031,N_1974,N_1925);
or U2032 (N_2032,N_1849,N_1967);
and U2033 (N_2033,N_1874,N_1821);
nor U2034 (N_2034,N_1951,N_1910);
nor U2035 (N_2035,N_1878,N_1948);
nand U2036 (N_2036,N_1844,N_1800);
nand U2037 (N_2037,N_1973,N_1838);
nand U2038 (N_2038,N_1947,N_1959);
and U2039 (N_2039,N_1895,N_1955);
or U2040 (N_2040,N_1856,N_1865);
or U2041 (N_2041,N_1825,N_1875);
or U2042 (N_2042,N_1881,N_1994);
nand U2043 (N_2043,N_1880,N_1990);
nor U2044 (N_2044,N_1939,N_1961);
or U2045 (N_2045,N_1851,N_1952);
and U2046 (N_2046,N_1868,N_1806);
nor U2047 (N_2047,N_1903,N_1893);
nor U2048 (N_2048,N_1960,N_1979);
nor U2049 (N_2049,N_1970,N_1935);
nor U2050 (N_2050,N_1812,N_1908);
nor U2051 (N_2051,N_1834,N_1892);
nand U2052 (N_2052,N_1842,N_1956);
nor U2053 (N_2053,N_1824,N_1869);
or U2054 (N_2054,N_1931,N_1932);
and U2055 (N_2055,N_1888,N_1837);
and U2056 (N_2056,N_1923,N_1965);
or U2057 (N_2057,N_1918,N_1870);
and U2058 (N_2058,N_1897,N_1827);
and U2059 (N_2059,N_1997,N_1989);
or U2060 (N_2060,N_1896,N_1941);
nand U2061 (N_2061,N_1867,N_1803);
nand U2062 (N_2062,N_1922,N_1815);
nor U2063 (N_2063,N_1982,N_1991);
nor U2064 (N_2064,N_1835,N_1980);
or U2065 (N_2065,N_1969,N_1809);
nand U2066 (N_2066,N_1985,N_1914);
nand U2067 (N_2067,N_1940,N_1902);
and U2068 (N_2068,N_1971,N_1836);
nand U2069 (N_2069,N_1829,N_1927);
and U2070 (N_2070,N_1861,N_1894);
or U2071 (N_2071,N_1871,N_1818);
nand U2072 (N_2072,N_1946,N_1906);
nand U2073 (N_2073,N_1855,N_1944);
or U2074 (N_2074,N_1816,N_1830);
nor U2075 (N_2075,N_1814,N_1938);
and U2076 (N_2076,N_1962,N_1890);
nor U2077 (N_2077,N_1853,N_1904);
or U2078 (N_2078,N_1984,N_1992);
nor U2079 (N_2079,N_1863,N_1988);
nor U2080 (N_2080,N_1998,N_1936);
nor U2081 (N_2081,N_1913,N_1924);
nor U2082 (N_2082,N_1864,N_1826);
or U2083 (N_2083,N_1943,N_1866);
nor U2084 (N_2084,N_1805,N_1915);
or U2085 (N_2085,N_1828,N_1911);
nor U2086 (N_2086,N_1886,N_1884);
nand U2087 (N_2087,N_1847,N_1977);
nand U2088 (N_2088,N_1987,N_1819);
or U2089 (N_2089,N_1872,N_1950);
nand U2090 (N_2090,N_1975,N_1920);
nor U2091 (N_2091,N_1883,N_1808);
or U2092 (N_2092,N_1898,N_1993);
nor U2093 (N_2093,N_1930,N_1983);
and U2094 (N_2094,N_1981,N_1937);
and U2095 (N_2095,N_1804,N_1995);
nand U2096 (N_2096,N_1859,N_1852);
and U2097 (N_2097,N_1933,N_1857);
nor U2098 (N_2098,N_1845,N_1942);
and U2099 (N_2099,N_1841,N_1802);
and U2100 (N_2100,N_1861,N_1974);
nand U2101 (N_2101,N_1904,N_1967);
and U2102 (N_2102,N_1892,N_1819);
or U2103 (N_2103,N_1941,N_1918);
or U2104 (N_2104,N_1827,N_1855);
or U2105 (N_2105,N_1886,N_1819);
or U2106 (N_2106,N_1905,N_1969);
nor U2107 (N_2107,N_1995,N_1931);
and U2108 (N_2108,N_1987,N_1820);
nor U2109 (N_2109,N_1958,N_1932);
xnor U2110 (N_2110,N_1830,N_1808);
or U2111 (N_2111,N_1824,N_1969);
and U2112 (N_2112,N_1854,N_1819);
nor U2113 (N_2113,N_1935,N_1808);
and U2114 (N_2114,N_1980,N_1972);
nand U2115 (N_2115,N_1947,N_1802);
nor U2116 (N_2116,N_1959,N_1992);
nor U2117 (N_2117,N_1941,N_1805);
or U2118 (N_2118,N_1825,N_1936);
nand U2119 (N_2119,N_1879,N_1929);
nand U2120 (N_2120,N_1984,N_1900);
nand U2121 (N_2121,N_1815,N_1860);
nand U2122 (N_2122,N_1876,N_1820);
or U2123 (N_2123,N_1901,N_1881);
or U2124 (N_2124,N_1845,N_1813);
nand U2125 (N_2125,N_1887,N_1994);
nor U2126 (N_2126,N_1860,N_1825);
nand U2127 (N_2127,N_1955,N_1981);
or U2128 (N_2128,N_1890,N_1964);
nor U2129 (N_2129,N_1854,N_1810);
nor U2130 (N_2130,N_1971,N_1959);
xnor U2131 (N_2131,N_1832,N_1965);
or U2132 (N_2132,N_1900,N_1828);
nand U2133 (N_2133,N_1817,N_1807);
nor U2134 (N_2134,N_1814,N_1906);
or U2135 (N_2135,N_1937,N_1916);
and U2136 (N_2136,N_1893,N_1945);
nor U2137 (N_2137,N_1889,N_1891);
and U2138 (N_2138,N_1809,N_1975);
xnor U2139 (N_2139,N_1980,N_1993);
and U2140 (N_2140,N_1973,N_1925);
or U2141 (N_2141,N_1984,N_1971);
nor U2142 (N_2142,N_1873,N_1810);
nand U2143 (N_2143,N_1813,N_1851);
nand U2144 (N_2144,N_1946,N_1992);
or U2145 (N_2145,N_1909,N_1815);
nand U2146 (N_2146,N_1803,N_1995);
and U2147 (N_2147,N_1927,N_1920);
nor U2148 (N_2148,N_1805,N_1991);
or U2149 (N_2149,N_1898,N_1873);
or U2150 (N_2150,N_1826,N_1801);
and U2151 (N_2151,N_1873,N_1839);
or U2152 (N_2152,N_1845,N_1850);
or U2153 (N_2153,N_1822,N_1958);
or U2154 (N_2154,N_1931,N_1817);
and U2155 (N_2155,N_1976,N_1852);
nand U2156 (N_2156,N_1845,N_1848);
or U2157 (N_2157,N_1943,N_1958);
nor U2158 (N_2158,N_1856,N_1826);
or U2159 (N_2159,N_1863,N_1832);
and U2160 (N_2160,N_1905,N_1961);
xnor U2161 (N_2161,N_1902,N_1999);
nor U2162 (N_2162,N_1820,N_1916);
nor U2163 (N_2163,N_1924,N_1819);
nor U2164 (N_2164,N_1928,N_1821);
nand U2165 (N_2165,N_1874,N_1944);
and U2166 (N_2166,N_1928,N_1936);
or U2167 (N_2167,N_1838,N_1974);
or U2168 (N_2168,N_1869,N_1989);
or U2169 (N_2169,N_1877,N_1928);
or U2170 (N_2170,N_1999,N_1857);
or U2171 (N_2171,N_1898,N_1872);
and U2172 (N_2172,N_1992,N_1958);
nor U2173 (N_2173,N_1903,N_1845);
nand U2174 (N_2174,N_1886,N_1833);
or U2175 (N_2175,N_1830,N_1975);
or U2176 (N_2176,N_1990,N_1806);
or U2177 (N_2177,N_1921,N_1847);
or U2178 (N_2178,N_1960,N_1859);
nor U2179 (N_2179,N_1889,N_1830);
and U2180 (N_2180,N_1920,N_1847);
nor U2181 (N_2181,N_1904,N_1969);
nor U2182 (N_2182,N_1981,N_1916);
and U2183 (N_2183,N_1975,N_1804);
nor U2184 (N_2184,N_1966,N_1961);
nor U2185 (N_2185,N_1963,N_1830);
or U2186 (N_2186,N_1801,N_1924);
and U2187 (N_2187,N_1997,N_1806);
and U2188 (N_2188,N_1952,N_1926);
nand U2189 (N_2189,N_1987,N_1941);
nor U2190 (N_2190,N_1831,N_1835);
or U2191 (N_2191,N_1856,N_1858);
and U2192 (N_2192,N_1872,N_1845);
nor U2193 (N_2193,N_1950,N_1873);
and U2194 (N_2194,N_1915,N_1833);
nand U2195 (N_2195,N_1851,N_1956);
nand U2196 (N_2196,N_1925,N_1982);
nor U2197 (N_2197,N_1912,N_1947);
nand U2198 (N_2198,N_1974,N_1834);
or U2199 (N_2199,N_1882,N_1936);
and U2200 (N_2200,N_2178,N_2006);
nand U2201 (N_2201,N_2000,N_2074);
and U2202 (N_2202,N_2156,N_2059);
nand U2203 (N_2203,N_2139,N_2123);
nand U2204 (N_2204,N_2021,N_2100);
and U2205 (N_2205,N_2192,N_2096);
or U2206 (N_2206,N_2141,N_2130);
nor U2207 (N_2207,N_2002,N_2189);
and U2208 (N_2208,N_2035,N_2152);
nand U2209 (N_2209,N_2098,N_2064);
and U2210 (N_2210,N_2171,N_2039);
nor U2211 (N_2211,N_2012,N_2165);
nand U2212 (N_2212,N_2174,N_2062);
nand U2213 (N_2213,N_2122,N_2125);
and U2214 (N_2214,N_2083,N_2082);
or U2215 (N_2215,N_2115,N_2131);
nor U2216 (N_2216,N_2190,N_2113);
or U2217 (N_2217,N_2187,N_2117);
nand U2218 (N_2218,N_2175,N_2066);
and U2219 (N_2219,N_2011,N_2069);
or U2220 (N_2220,N_2079,N_2181);
or U2221 (N_2221,N_2157,N_2055);
or U2222 (N_2222,N_2153,N_2183);
nor U2223 (N_2223,N_2060,N_2080);
xor U2224 (N_2224,N_2101,N_2112);
nor U2225 (N_2225,N_2032,N_2145);
nand U2226 (N_2226,N_2163,N_2196);
or U2227 (N_2227,N_2084,N_2065);
nor U2228 (N_2228,N_2159,N_2017);
and U2229 (N_2229,N_2118,N_2048);
nor U2230 (N_2230,N_2133,N_2132);
xor U2231 (N_2231,N_2013,N_2151);
and U2232 (N_2232,N_2168,N_2107);
or U2233 (N_2233,N_2007,N_2023);
and U2234 (N_2234,N_2193,N_2028);
nand U2235 (N_2235,N_2050,N_2126);
nor U2236 (N_2236,N_2137,N_2049);
nand U2237 (N_2237,N_2018,N_2036);
and U2238 (N_2238,N_2169,N_2073);
and U2239 (N_2239,N_2185,N_2092);
nor U2240 (N_2240,N_2146,N_2086);
or U2241 (N_2241,N_2182,N_2162);
nor U2242 (N_2242,N_2143,N_2186);
nor U2243 (N_2243,N_2005,N_2078);
or U2244 (N_2244,N_2054,N_2158);
nand U2245 (N_2245,N_2010,N_2105);
or U2246 (N_2246,N_2097,N_2024);
or U2247 (N_2247,N_2135,N_2104);
or U2248 (N_2248,N_2176,N_2184);
nand U2249 (N_2249,N_2191,N_2003);
nand U2250 (N_2250,N_2087,N_2094);
and U2251 (N_2251,N_2026,N_2119);
or U2252 (N_2252,N_2091,N_2045);
or U2253 (N_2253,N_2063,N_2128);
or U2254 (N_2254,N_2161,N_2172);
xor U2255 (N_2255,N_2046,N_2016);
and U2256 (N_2256,N_2194,N_2030);
nand U2257 (N_2257,N_2150,N_2170);
or U2258 (N_2258,N_2103,N_2042);
nor U2259 (N_2259,N_2188,N_2110);
or U2260 (N_2260,N_2077,N_2124);
or U2261 (N_2261,N_2076,N_2154);
nor U2262 (N_2262,N_2052,N_2136);
or U2263 (N_2263,N_2167,N_2095);
or U2264 (N_2264,N_2040,N_2106);
or U2265 (N_2265,N_2058,N_2198);
nor U2266 (N_2266,N_2047,N_2071);
or U2267 (N_2267,N_2027,N_2015);
nor U2268 (N_2268,N_2034,N_2138);
and U2269 (N_2269,N_2085,N_2142);
nand U2270 (N_2270,N_2037,N_2116);
or U2271 (N_2271,N_2075,N_2056);
nand U2272 (N_2272,N_2164,N_2111);
and U2273 (N_2273,N_2108,N_2009);
and U2274 (N_2274,N_2089,N_2144);
xor U2275 (N_2275,N_2041,N_2070);
nor U2276 (N_2276,N_2134,N_2127);
and U2277 (N_2277,N_2114,N_2102);
and U2278 (N_2278,N_2180,N_2090);
nor U2279 (N_2279,N_2025,N_2099);
and U2280 (N_2280,N_2001,N_2197);
or U2281 (N_2281,N_2109,N_2014);
and U2282 (N_2282,N_2053,N_2072);
nor U2283 (N_2283,N_2179,N_2044);
and U2284 (N_2284,N_2155,N_2008);
nor U2285 (N_2285,N_2020,N_2068);
nor U2286 (N_2286,N_2088,N_2022);
or U2287 (N_2287,N_2140,N_2067);
nor U2288 (N_2288,N_2129,N_2081);
nand U2289 (N_2289,N_2160,N_2004);
and U2290 (N_2290,N_2120,N_2121);
nor U2291 (N_2291,N_2033,N_2199);
or U2292 (N_2292,N_2148,N_2166);
nor U2293 (N_2293,N_2093,N_2029);
and U2294 (N_2294,N_2051,N_2038);
or U2295 (N_2295,N_2031,N_2177);
nand U2296 (N_2296,N_2057,N_2061);
nand U2297 (N_2297,N_2173,N_2149);
nand U2298 (N_2298,N_2043,N_2147);
or U2299 (N_2299,N_2195,N_2019);
or U2300 (N_2300,N_2160,N_2136);
or U2301 (N_2301,N_2018,N_2199);
or U2302 (N_2302,N_2083,N_2191);
nor U2303 (N_2303,N_2185,N_2123);
and U2304 (N_2304,N_2176,N_2005);
and U2305 (N_2305,N_2005,N_2011);
nor U2306 (N_2306,N_2034,N_2045);
or U2307 (N_2307,N_2065,N_2003);
or U2308 (N_2308,N_2175,N_2103);
xor U2309 (N_2309,N_2082,N_2107);
nand U2310 (N_2310,N_2187,N_2119);
or U2311 (N_2311,N_2084,N_2057);
and U2312 (N_2312,N_2083,N_2016);
nand U2313 (N_2313,N_2093,N_2036);
nor U2314 (N_2314,N_2028,N_2110);
and U2315 (N_2315,N_2035,N_2029);
nand U2316 (N_2316,N_2178,N_2130);
and U2317 (N_2317,N_2120,N_2166);
nand U2318 (N_2318,N_2138,N_2195);
nor U2319 (N_2319,N_2154,N_2020);
or U2320 (N_2320,N_2190,N_2049);
and U2321 (N_2321,N_2133,N_2154);
nand U2322 (N_2322,N_2124,N_2176);
nor U2323 (N_2323,N_2018,N_2043);
nand U2324 (N_2324,N_2049,N_2066);
nor U2325 (N_2325,N_2038,N_2023);
and U2326 (N_2326,N_2183,N_2186);
nor U2327 (N_2327,N_2014,N_2107);
nand U2328 (N_2328,N_2069,N_2112);
nand U2329 (N_2329,N_2066,N_2051);
or U2330 (N_2330,N_2061,N_2048);
or U2331 (N_2331,N_2131,N_2068);
or U2332 (N_2332,N_2065,N_2122);
and U2333 (N_2333,N_2129,N_2196);
and U2334 (N_2334,N_2170,N_2061);
or U2335 (N_2335,N_2124,N_2173);
or U2336 (N_2336,N_2123,N_2075);
nand U2337 (N_2337,N_2125,N_2077);
nand U2338 (N_2338,N_2039,N_2159);
and U2339 (N_2339,N_2125,N_2142);
and U2340 (N_2340,N_2159,N_2077);
nor U2341 (N_2341,N_2143,N_2010);
or U2342 (N_2342,N_2138,N_2054);
or U2343 (N_2343,N_2084,N_2005);
nor U2344 (N_2344,N_2059,N_2092);
or U2345 (N_2345,N_2072,N_2027);
or U2346 (N_2346,N_2066,N_2102);
and U2347 (N_2347,N_2112,N_2184);
or U2348 (N_2348,N_2026,N_2182);
or U2349 (N_2349,N_2195,N_2086);
nand U2350 (N_2350,N_2080,N_2031);
or U2351 (N_2351,N_2189,N_2059);
nand U2352 (N_2352,N_2174,N_2112);
or U2353 (N_2353,N_2146,N_2142);
or U2354 (N_2354,N_2066,N_2129);
or U2355 (N_2355,N_2058,N_2196);
and U2356 (N_2356,N_2178,N_2020);
or U2357 (N_2357,N_2128,N_2145);
or U2358 (N_2358,N_2040,N_2160);
nor U2359 (N_2359,N_2040,N_2042);
nand U2360 (N_2360,N_2189,N_2060);
nand U2361 (N_2361,N_2031,N_2060);
or U2362 (N_2362,N_2112,N_2178);
and U2363 (N_2363,N_2028,N_2109);
nor U2364 (N_2364,N_2109,N_2146);
and U2365 (N_2365,N_2086,N_2194);
or U2366 (N_2366,N_2156,N_2140);
nand U2367 (N_2367,N_2008,N_2100);
and U2368 (N_2368,N_2095,N_2064);
nor U2369 (N_2369,N_2053,N_2184);
nor U2370 (N_2370,N_2163,N_2168);
and U2371 (N_2371,N_2130,N_2134);
nand U2372 (N_2372,N_2138,N_2167);
nor U2373 (N_2373,N_2034,N_2026);
or U2374 (N_2374,N_2034,N_2178);
or U2375 (N_2375,N_2015,N_2139);
nand U2376 (N_2376,N_2159,N_2199);
nor U2377 (N_2377,N_2132,N_2082);
or U2378 (N_2378,N_2093,N_2081);
nand U2379 (N_2379,N_2055,N_2148);
xor U2380 (N_2380,N_2152,N_2043);
or U2381 (N_2381,N_2101,N_2026);
and U2382 (N_2382,N_2107,N_2109);
and U2383 (N_2383,N_2143,N_2062);
and U2384 (N_2384,N_2093,N_2020);
nor U2385 (N_2385,N_2102,N_2087);
and U2386 (N_2386,N_2161,N_2116);
and U2387 (N_2387,N_2040,N_2038);
nand U2388 (N_2388,N_2042,N_2060);
or U2389 (N_2389,N_2173,N_2100);
nand U2390 (N_2390,N_2162,N_2066);
xor U2391 (N_2391,N_2020,N_2038);
nand U2392 (N_2392,N_2190,N_2059);
or U2393 (N_2393,N_2004,N_2185);
or U2394 (N_2394,N_2120,N_2182);
xnor U2395 (N_2395,N_2006,N_2032);
or U2396 (N_2396,N_2041,N_2149);
and U2397 (N_2397,N_2146,N_2116);
and U2398 (N_2398,N_2186,N_2064);
or U2399 (N_2399,N_2011,N_2193);
and U2400 (N_2400,N_2346,N_2308);
and U2401 (N_2401,N_2256,N_2222);
nor U2402 (N_2402,N_2329,N_2315);
or U2403 (N_2403,N_2372,N_2267);
xor U2404 (N_2404,N_2352,N_2397);
nor U2405 (N_2405,N_2236,N_2269);
or U2406 (N_2406,N_2284,N_2369);
and U2407 (N_2407,N_2215,N_2338);
and U2408 (N_2408,N_2304,N_2335);
and U2409 (N_2409,N_2207,N_2341);
xor U2410 (N_2410,N_2312,N_2272);
or U2411 (N_2411,N_2374,N_2219);
nand U2412 (N_2412,N_2317,N_2293);
or U2413 (N_2413,N_2208,N_2362);
nor U2414 (N_2414,N_2251,N_2387);
nor U2415 (N_2415,N_2376,N_2339);
xnor U2416 (N_2416,N_2309,N_2370);
nor U2417 (N_2417,N_2203,N_2368);
nor U2418 (N_2418,N_2386,N_2231);
xor U2419 (N_2419,N_2205,N_2380);
nor U2420 (N_2420,N_2201,N_2384);
or U2421 (N_2421,N_2225,N_2307);
or U2422 (N_2422,N_2233,N_2393);
or U2423 (N_2423,N_2381,N_2286);
nand U2424 (N_2424,N_2212,N_2248);
nand U2425 (N_2425,N_2318,N_2295);
nand U2426 (N_2426,N_2358,N_2282);
or U2427 (N_2427,N_2323,N_2273);
and U2428 (N_2428,N_2213,N_2328);
nor U2429 (N_2429,N_2396,N_2357);
nand U2430 (N_2430,N_2363,N_2230);
and U2431 (N_2431,N_2217,N_2302);
nor U2432 (N_2432,N_2324,N_2390);
and U2433 (N_2433,N_2259,N_2237);
and U2434 (N_2434,N_2264,N_2361);
and U2435 (N_2435,N_2223,N_2200);
and U2436 (N_2436,N_2377,N_2257);
nor U2437 (N_2437,N_2221,N_2331);
nand U2438 (N_2438,N_2296,N_2306);
nand U2439 (N_2439,N_2316,N_2245);
or U2440 (N_2440,N_2399,N_2266);
or U2441 (N_2441,N_2395,N_2210);
and U2442 (N_2442,N_2303,N_2322);
xor U2443 (N_2443,N_2206,N_2263);
or U2444 (N_2444,N_2297,N_2244);
nand U2445 (N_2445,N_2355,N_2277);
nor U2446 (N_2446,N_2239,N_2270);
or U2447 (N_2447,N_2343,N_2228);
and U2448 (N_2448,N_2226,N_2385);
nand U2449 (N_2449,N_2276,N_2294);
and U2450 (N_2450,N_2271,N_2325);
nand U2451 (N_2451,N_2389,N_2373);
nor U2452 (N_2452,N_2242,N_2275);
nand U2453 (N_2453,N_2319,N_2224);
nor U2454 (N_2454,N_2383,N_2349);
or U2455 (N_2455,N_2249,N_2285);
nor U2456 (N_2456,N_2364,N_2252);
nor U2457 (N_2457,N_2337,N_2262);
or U2458 (N_2458,N_2209,N_2365);
nor U2459 (N_2459,N_2243,N_2246);
or U2460 (N_2460,N_2391,N_2238);
nor U2461 (N_2461,N_2340,N_2394);
nor U2462 (N_2462,N_2332,N_2378);
or U2463 (N_2463,N_2289,N_2311);
nand U2464 (N_2464,N_2356,N_2298);
and U2465 (N_2465,N_2392,N_2281);
nor U2466 (N_2466,N_2287,N_2371);
nand U2467 (N_2467,N_2204,N_2314);
or U2468 (N_2468,N_2300,N_2348);
nand U2469 (N_2469,N_2260,N_2388);
nor U2470 (N_2470,N_2274,N_2354);
nand U2471 (N_2471,N_2327,N_2218);
or U2472 (N_2472,N_2216,N_2220);
nor U2473 (N_2473,N_2214,N_2350);
xor U2474 (N_2474,N_2344,N_2268);
and U2475 (N_2475,N_2310,N_2250);
and U2476 (N_2476,N_2288,N_2353);
nor U2477 (N_2477,N_2254,N_2336);
and U2478 (N_2478,N_2235,N_2326);
or U2479 (N_2479,N_2313,N_2279);
and U2480 (N_2480,N_2299,N_2247);
nor U2481 (N_2481,N_2292,N_2241);
nand U2482 (N_2482,N_2320,N_2301);
nor U2483 (N_2483,N_2345,N_2382);
or U2484 (N_2484,N_2280,N_2334);
nor U2485 (N_2485,N_2366,N_2232);
or U2486 (N_2486,N_2229,N_2255);
nand U2487 (N_2487,N_2261,N_2321);
or U2488 (N_2488,N_2305,N_2290);
and U2489 (N_2489,N_2330,N_2398);
nor U2490 (N_2490,N_2211,N_2202);
or U2491 (N_2491,N_2265,N_2234);
nand U2492 (N_2492,N_2367,N_2351);
xnor U2493 (N_2493,N_2278,N_2347);
and U2494 (N_2494,N_2359,N_2360);
nor U2495 (N_2495,N_2253,N_2258);
nor U2496 (N_2496,N_2379,N_2240);
nor U2497 (N_2497,N_2227,N_2291);
nor U2498 (N_2498,N_2333,N_2283);
nor U2499 (N_2499,N_2375,N_2342);
nor U2500 (N_2500,N_2351,N_2373);
nand U2501 (N_2501,N_2216,N_2201);
nor U2502 (N_2502,N_2294,N_2392);
nand U2503 (N_2503,N_2323,N_2249);
nand U2504 (N_2504,N_2355,N_2208);
and U2505 (N_2505,N_2211,N_2389);
and U2506 (N_2506,N_2307,N_2233);
xnor U2507 (N_2507,N_2307,N_2379);
or U2508 (N_2508,N_2286,N_2386);
nor U2509 (N_2509,N_2309,N_2320);
and U2510 (N_2510,N_2223,N_2306);
or U2511 (N_2511,N_2256,N_2341);
nand U2512 (N_2512,N_2322,N_2352);
nand U2513 (N_2513,N_2366,N_2230);
nand U2514 (N_2514,N_2371,N_2261);
nand U2515 (N_2515,N_2234,N_2286);
and U2516 (N_2516,N_2245,N_2330);
nand U2517 (N_2517,N_2338,N_2331);
nand U2518 (N_2518,N_2209,N_2244);
nand U2519 (N_2519,N_2357,N_2213);
nor U2520 (N_2520,N_2316,N_2261);
or U2521 (N_2521,N_2362,N_2356);
or U2522 (N_2522,N_2311,N_2200);
nand U2523 (N_2523,N_2322,N_2258);
nor U2524 (N_2524,N_2208,N_2376);
and U2525 (N_2525,N_2289,N_2357);
or U2526 (N_2526,N_2256,N_2381);
nor U2527 (N_2527,N_2267,N_2390);
nand U2528 (N_2528,N_2333,N_2287);
or U2529 (N_2529,N_2359,N_2240);
and U2530 (N_2530,N_2360,N_2324);
and U2531 (N_2531,N_2327,N_2329);
nor U2532 (N_2532,N_2227,N_2269);
nand U2533 (N_2533,N_2233,N_2264);
or U2534 (N_2534,N_2274,N_2326);
or U2535 (N_2535,N_2247,N_2337);
nor U2536 (N_2536,N_2342,N_2206);
nor U2537 (N_2537,N_2234,N_2211);
and U2538 (N_2538,N_2226,N_2293);
and U2539 (N_2539,N_2209,N_2343);
or U2540 (N_2540,N_2354,N_2356);
or U2541 (N_2541,N_2206,N_2253);
and U2542 (N_2542,N_2285,N_2219);
nand U2543 (N_2543,N_2363,N_2240);
or U2544 (N_2544,N_2322,N_2366);
nand U2545 (N_2545,N_2214,N_2380);
and U2546 (N_2546,N_2298,N_2309);
or U2547 (N_2547,N_2245,N_2309);
nand U2548 (N_2548,N_2206,N_2314);
and U2549 (N_2549,N_2332,N_2245);
nor U2550 (N_2550,N_2363,N_2398);
nor U2551 (N_2551,N_2248,N_2334);
nor U2552 (N_2552,N_2277,N_2301);
and U2553 (N_2553,N_2253,N_2280);
nor U2554 (N_2554,N_2219,N_2232);
nor U2555 (N_2555,N_2243,N_2291);
and U2556 (N_2556,N_2379,N_2237);
nor U2557 (N_2557,N_2219,N_2323);
or U2558 (N_2558,N_2395,N_2258);
or U2559 (N_2559,N_2206,N_2327);
and U2560 (N_2560,N_2228,N_2217);
or U2561 (N_2561,N_2224,N_2361);
nor U2562 (N_2562,N_2246,N_2305);
nor U2563 (N_2563,N_2397,N_2363);
and U2564 (N_2564,N_2263,N_2363);
nor U2565 (N_2565,N_2200,N_2221);
and U2566 (N_2566,N_2391,N_2235);
nand U2567 (N_2567,N_2277,N_2386);
or U2568 (N_2568,N_2212,N_2228);
nand U2569 (N_2569,N_2215,N_2376);
nor U2570 (N_2570,N_2308,N_2340);
nor U2571 (N_2571,N_2387,N_2260);
or U2572 (N_2572,N_2247,N_2365);
nand U2573 (N_2573,N_2289,N_2281);
or U2574 (N_2574,N_2272,N_2307);
nand U2575 (N_2575,N_2390,N_2278);
nand U2576 (N_2576,N_2369,N_2373);
and U2577 (N_2577,N_2383,N_2241);
and U2578 (N_2578,N_2218,N_2281);
nand U2579 (N_2579,N_2237,N_2229);
nor U2580 (N_2580,N_2309,N_2284);
nand U2581 (N_2581,N_2313,N_2360);
nor U2582 (N_2582,N_2344,N_2345);
nor U2583 (N_2583,N_2305,N_2273);
or U2584 (N_2584,N_2391,N_2228);
or U2585 (N_2585,N_2276,N_2267);
nor U2586 (N_2586,N_2250,N_2391);
nand U2587 (N_2587,N_2255,N_2385);
nand U2588 (N_2588,N_2262,N_2388);
or U2589 (N_2589,N_2283,N_2256);
nand U2590 (N_2590,N_2308,N_2330);
and U2591 (N_2591,N_2278,N_2320);
nand U2592 (N_2592,N_2285,N_2289);
nor U2593 (N_2593,N_2325,N_2331);
xnor U2594 (N_2594,N_2313,N_2382);
xnor U2595 (N_2595,N_2352,N_2206);
nand U2596 (N_2596,N_2302,N_2269);
nor U2597 (N_2597,N_2279,N_2229);
nor U2598 (N_2598,N_2273,N_2345);
nor U2599 (N_2599,N_2288,N_2210);
and U2600 (N_2600,N_2400,N_2551);
and U2601 (N_2601,N_2485,N_2525);
nand U2602 (N_2602,N_2481,N_2435);
and U2603 (N_2603,N_2473,N_2430);
nand U2604 (N_2604,N_2476,N_2433);
and U2605 (N_2605,N_2445,N_2508);
and U2606 (N_2606,N_2513,N_2571);
nor U2607 (N_2607,N_2480,N_2450);
or U2608 (N_2608,N_2470,N_2500);
nor U2609 (N_2609,N_2415,N_2514);
nor U2610 (N_2610,N_2575,N_2568);
or U2611 (N_2611,N_2589,N_2558);
or U2612 (N_2612,N_2465,N_2419);
nand U2613 (N_2613,N_2520,N_2518);
nand U2614 (N_2614,N_2507,N_2454);
nand U2615 (N_2615,N_2488,N_2572);
and U2616 (N_2616,N_2417,N_2538);
nor U2617 (N_2617,N_2505,N_2545);
nor U2618 (N_2618,N_2526,N_2477);
nand U2619 (N_2619,N_2464,N_2584);
nand U2620 (N_2620,N_2401,N_2421);
or U2621 (N_2621,N_2418,N_2493);
nand U2622 (N_2622,N_2489,N_2527);
nand U2623 (N_2623,N_2595,N_2528);
nor U2624 (N_2624,N_2586,N_2449);
nand U2625 (N_2625,N_2497,N_2591);
or U2626 (N_2626,N_2599,N_2482);
or U2627 (N_2627,N_2455,N_2533);
nor U2628 (N_2628,N_2561,N_2451);
and U2629 (N_2629,N_2587,N_2524);
nand U2630 (N_2630,N_2531,N_2462);
and U2631 (N_2631,N_2427,N_2407);
nand U2632 (N_2632,N_2429,N_2544);
or U2633 (N_2633,N_2490,N_2475);
and U2634 (N_2634,N_2425,N_2569);
nor U2635 (N_2635,N_2557,N_2576);
or U2636 (N_2636,N_2516,N_2431);
nor U2637 (N_2637,N_2532,N_2484);
or U2638 (N_2638,N_2494,N_2550);
or U2639 (N_2639,N_2438,N_2502);
and U2640 (N_2640,N_2441,N_2487);
xor U2641 (N_2641,N_2456,N_2578);
xor U2642 (N_2642,N_2521,N_2588);
nand U2643 (N_2643,N_2432,N_2553);
nor U2644 (N_2644,N_2512,N_2519);
xnor U2645 (N_2645,N_2463,N_2406);
and U2646 (N_2646,N_2403,N_2556);
nor U2647 (N_2647,N_2579,N_2597);
nand U2648 (N_2648,N_2469,N_2426);
nor U2649 (N_2649,N_2436,N_2453);
nand U2650 (N_2650,N_2444,N_2496);
nand U2651 (N_2651,N_2548,N_2536);
or U2652 (N_2652,N_2459,N_2420);
or U2653 (N_2653,N_2468,N_2580);
and U2654 (N_2654,N_2478,N_2534);
nor U2655 (N_2655,N_2539,N_2428);
or U2656 (N_2656,N_2509,N_2565);
nand U2657 (N_2657,N_2461,N_2592);
or U2658 (N_2658,N_2416,N_2452);
or U2659 (N_2659,N_2559,N_2535);
or U2660 (N_2660,N_2479,N_2474);
nand U2661 (N_2661,N_2555,N_2540);
nand U2662 (N_2662,N_2404,N_2408);
nor U2663 (N_2663,N_2501,N_2537);
nand U2664 (N_2664,N_2590,N_2447);
nor U2665 (N_2665,N_2495,N_2547);
or U2666 (N_2666,N_2446,N_2577);
nand U2667 (N_2667,N_2504,N_2522);
and U2668 (N_2668,N_2457,N_2471);
or U2669 (N_2669,N_2424,N_2409);
nor U2670 (N_2670,N_2552,N_2411);
nor U2671 (N_2671,N_2412,N_2563);
and U2672 (N_2672,N_2510,N_2570);
nor U2673 (N_2673,N_2582,N_2499);
and U2674 (N_2674,N_2439,N_2574);
or U2675 (N_2675,N_2546,N_2414);
and U2676 (N_2676,N_2562,N_2529);
xor U2677 (N_2677,N_2581,N_2492);
nand U2678 (N_2678,N_2434,N_2498);
and U2679 (N_2679,N_2560,N_2573);
and U2680 (N_2680,N_2402,N_2437);
nor U2681 (N_2681,N_2472,N_2467);
nand U2682 (N_2682,N_2486,N_2413);
nor U2683 (N_2683,N_2460,N_2466);
xnor U2684 (N_2684,N_2440,N_2598);
or U2685 (N_2685,N_2506,N_2530);
nand U2686 (N_2686,N_2549,N_2442);
nor U2687 (N_2687,N_2443,N_2423);
and U2688 (N_2688,N_2517,N_2554);
nor U2689 (N_2689,N_2594,N_2543);
or U2690 (N_2690,N_2491,N_2458);
and U2691 (N_2691,N_2422,N_2483);
nand U2692 (N_2692,N_2542,N_2596);
nand U2693 (N_2693,N_2585,N_2448);
nand U2694 (N_2694,N_2567,N_2511);
and U2695 (N_2695,N_2515,N_2523);
or U2696 (N_2696,N_2410,N_2541);
nand U2697 (N_2697,N_2564,N_2405);
or U2698 (N_2698,N_2503,N_2566);
or U2699 (N_2699,N_2583,N_2593);
and U2700 (N_2700,N_2506,N_2591);
or U2701 (N_2701,N_2453,N_2496);
or U2702 (N_2702,N_2563,N_2479);
nand U2703 (N_2703,N_2583,N_2422);
or U2704 (N_2704,N_2461,N_2536);
nand U2705 (N_2705,N_2402,N_2514);
and U2706 (N_2706,N_2509,N_2539);
nand U2707 (N_2707,N_2542,N_2563);
nor U2708 (N_2708,N_2520,N_2424);
or U2709 (N_2709,N_2515,N_2561);
or U2710 (N_2710,N_2450,N_2580);
nor U2711 (N_2711,N_2417,N_2585);
nand U2712 (N_2712,N_2587,N_2506);
nand U2713 (N_2713,N_2506,N_2444);
nand U2714 (N_2714,N_2591,N_2527);
nor U2715 (N_2715,N_2542,N_2571);
xor U2716 (N_2716,N_2424,N_2554);
nand U2717 (N_2717,N_2598,N_2457);
or U2718 (N_2718,N_2499,N_2458);
and U2719 (N_2719,N_2593,N_2502);
nor U2720 (N_2720,N_2430,N_2515);
and U2721 (N_2721,N_2490,N_2504);
nor U2722 (N_2722,N_2499,N_2459);
and U2723 (N_2723,N_2457,N_2497);
nor U2724 (N_2724,N_2572,N_2592);
nor U2725 (N_2725,N_2455,N_2400);
xnor U2726 (N_2726,N_2480,N_2494);
nand U2727 (N_2727,N_2517,N_2448);
and U2728 (N_2728,N_2432,N_2482);
or U2729 (N_2729,N_2588,N_2410);
nand U2730 (N_2730,N_2415,N_2492);
or U2731 (N_2731,N_2481,N_2434);
nand U2732 (N_2732,N_2554,N_2418);
nor U2733 (N_2733,N_2483,N_2429);
or U2734 (N_2734,N_2534,N_2559);
and U2735 (N_2735,N_2451,N_2404);
and U2736 (N_2736,N_2577,N_2425);
nor U2737 (N_2737,N_2493,N_2590);
or U2738 (N_2738,N_2591,N_2405);
or U2739 (N_2739,N_2523,N_2545);
nor U2740 (N_2740,N_2593,N_2530);
xnor U2741 (N_2741,N_2492,N_2419);
or U2742 (N_2742,N_2453,N_2462);
and U2743 (N_2743,N_2438,N_2554);
nor U2744 (N_2744,N_2599,N_2553);
and U2745 (N_2745,N_2426,N_2558);
or U2746 (N_2746,N_2417,N_2527);
or U2747 (N_2747,N_2431,N_2560);
nor U2748 (N_2748,N_2563,N_2428);
xnor U2749 (N_2749,N_2441,N_2554);
and U2750 (N_2750,N_2411,N_2529);
nand U2751 (N_2751,N_2594,N_2504);
nor U2752 (N_2752,N_2595,N_2555);
or U2753 (N_2753,N_2484,N_2488);
nand U2754 (N_2754,N_2458,N_2571);
and U2755 (N_2755,N_2402,N_2448);
nor U2756 (N_2756,N_2596,N_2591);
nor U2757 (N_2757,N_2598,N_2406);
or U2758 (N_2758,N_2562,N_2502);
and U2759 (N_2759,N_2504,N_2552);
nand U2760 (N_2760,N_2488,N_2506);
nand U2761 (N_2761,N_2589,N_2525);
nand U2762 (N_2762,N_2402,N_2508);
and U2763 (N_2763,N_2445,N_2580);
nor U2764 (N_2764,N_2536,N_2552);
and U2765 (N_2765,N_2433,N_2412);
nor U2766 (N_2766,N_2429,N_2490);
or U2767 (N_2767,N_2526,N_2470);
and U2768 (N_2768,N_2404,N_2589);
nor U2769 (N_2769,N_2535,N_2446);
and U2770 (N_2770,N_2536,N_2544);
or U2771 (N_2771,N_2445,N_2496);
nand U2772 (N_2772,N_2439,N_2545);
nand U2773 (N_2773,N_2494,N_2457);
nand U2774 (N_2774,N_2430,N_2518);
or U2775 (N_2775,N_2519,N_2545);
or U2776 (N_2776,N_2540,N_2576);
or U2777 (N_2777,N_2416,N_2406);
nor U2778 (N_2778,N_2441,N_2523);
or U2779 (N_2779,N_2498,N_2482);
nand U2780 (N_2780,N_2573,N_2593);
or U2781 (N_2781,N_2509,N_2469);
or U2782 (N_2782,N_2548,N_2422);
or U2783 (N_2783,N_2485,N_2535);
xnor U2784 (N_2784,N_2541,N_2403);
nand U2785 (N_2785,N_2498,N_2510);
and U2786 (N_2786,N_2542,N_2541);
nor U2787 (N_2787,N_2593,N_2469);
or U2788 (N_2788,N_2566,N_2454);
or U2789 (N_2789,N_2427,N_2481);
and U2790 (N_2790,N_2550,N_2520);
or U2791 (N_2791,N_2460,N_2437);
and U2792 (N_2792,N_2423,N_2495);
nand U2793 (N_2793,N_2553,N_2426);
and U2794 (N_2794,N_2592,N_2563);
or U2795 (N_2795,N_2467,N_2497);
nand U2796 (N_2796,N_2502,N_2557);
and U2797 (N_2797,N_2517,N_2475);
nand U2798 (N_2798,N_2526,N_2428);
and U2799 (N_2799,N_2485,N_2472);
or U2800 (N_2800,N_2785,N_2710);
and U2801 (N_2801,N_2743,N_2773);
nor U2802 (N_2802,N_2675,N_2715);
and U2803 (N_2803,N_2667,N_2765);
or U2804 (N_2804,N_2629,N_2700);
nand U2805 (N_2805,N_2607,N_2644);
or U2806 (N_2806,N_2712,N_2732);
nor U2807 (N_2807,N_2796,N_2620);
or U2808 (N_2808,N_2774,N_2779);
nand U2809 (N_2809,N_2631,N_2693);
nand U2810 (N_2810,N_2786,N_2672);
and U2811 (N_2811,N_2709,N_2737);
nand U2812 (N_2812,N_2604,N_2782);
and U2813 (N_2813,N_2600,N_2744);
nor U2814 (N_2814,N_2689,N_2741);
nor U2815 (N_2815,N_2777,N_2795);
nand U2816 (N_2816,N_2764,N_2756);
nor U2817 (N_2817,N_2701,N_2725);
nand U2818 (N_2818,N_2688,N_2770);
nand U2819 (N_2819,N_2625,N_2703);
nor U2820 (N_2820,N_2720,N_2788);
and U2821 (N_2821,N_2601,N_2747);
or U2822 (N_2822,N_2781,N_2727);
and U2823 (N_2823,N_2618,N_2642);
nor U2824 (N_2824,N_2608,N_2664);
or U2825 (N_2825,N_2706,N_2739);
nand U2826 (N_2826,N_2661,N_2750);
or U2827 (N_2827,N_2665,N_2656);
or U2828 (N_2828,N_2673,N_2617);
nand U2829 (N_2829,N_2746,N_2717);
nor U2830 (N_2830,N_2679,N_2798);
nand U2831 (N_2831,N_2775,N_2692);
xnor U2832 (N_2832,N_2682,N_2632);
nor U2833 (N_2833,N_2799,N_2695);
and U2834 (N_2834,N_2767,N_2610);
nor U2835 (N_2835,N_2748,N_2615);
and U2836 (N_2836,N_2776,N_2755);
or U2837 (N_2837,N_2702,N_2762);
and U2838 (N_2838,N_2766,N_2694);
and U2839 (N_2839,N_2760,N_2622);
or U2840 (N_2840,N_2678,N_2635);
nand U2841 (N_2841,N_2787,N_2687);
nor U2842 (N_2842,N_2613,N_2722);
nand U2843 (N_2843,N_2714,N_2657);
nor U2844 (N_2844,N_2794,N_2772);
nand U2845 (N_2845,N_2699,N_2628);
nand U2846 (N_2846,N_2789,N_2690);
and U2847 (N_2847,N_2677,N_2757);
or U2848 (N_2848,N_2745,N_2684);
nor U2849 (N_2849,N_2650,N_2666);
or U2850 (N_2850,N_2645,N_2705);
or U2851 (N_2851,N_2680,N_2659);
nand U2852 (N_2852,N_2754,N_2738);
nand U2853 (N_2853,N_2609,N_2627);
or U2854 (N_2854,N_2728,N_2637);
nor U2855 (N_2855,N_2638,N_2771);
nor U2856 (N_2856,N_2780,N_2749);
nand U2857 (N_2857,N_2752,N_2653);
or U2858 (N_2858,N_2730,N_2648);
and U2859 (N_2859,N_2669,N_2671);
nor U2860 (N_2860,N_2654,N_2704);
nor U2861 (N_2861,N_2621,N_2668);
nand U2862 (N_2862,N_2792,N_2655);
xor U2863 (N_2863,N_2611,N_2734);
or U2864 (N_2864,N_2753,N_2691);
or U2865 (N_2865,N_2751,N_2683);
and U2866 (N_2866,N_2778,N_2769);
or U2867 (N_2867,N_2763,N_2793);
nor U2868 (N_2868,N_2652,N_2731);
nor U2869 (N_2869,N_2640,N_2686);
nand U2870 (N_2870,N_2797,N_2740);
nor U2871 (N_2871,N_2658,N_2681);
nand U2872 (N_2872,N_2724,N_2616);
and U2873 (N_2873,N_2729,N_2707);
nand U2874 (N_2874,N_2761,N_2643);
or U2875 (N_2875,N_2735,N_2624);
and U2876 (N_2876,N_2719,N_2612);
and U2877 (N_2877,N_2649,N_2718);
nor U2878 (N_2878,N_2606,N_2742);
or U2879 (N_2879,N_2721,N_2783);
or U2880 (N_2880,N_2713,N_2736);
or U2881 (N_2881,N_2790,N_2660);
nand U2882 (N_2882,N_2662,N_2676);
nor U2883 (N_2883,N_2634,N_2758);
nand U2884 (N_2884,N_2602,N_2711);
nand U2885 (N_2885,N_2674,N_2716);
nand U2886 (N_2886,N_2685,N_2733);
nand U2887 (N_2887,N_2623,N_2614);
or U2888 (N_2888,N_2670,N_2641);
nor U2889 (N_2889,N_2605,N_2708);
or U2890 (N_2890,N_2726,N_2636);
nor U2891 (N_2891,N_2647,N_2626);
and U2892 (N_2892,N_2723,N_2630);
and U2893 (N_2893,N_2651,N_2663);
nand U2894 (N_2894,N_2603,N_2791);
and U2895 (N_2895,N_2696,N_2697);
nor U2896 (N_2896,N_2759,N_2633);
nand U2897 (N_2897,N_2619,N_2768);
nand U2898 (N_2898,N_2784,N_2639);
nand U2899 (N_2899,N_2698,N_2646);
or U2900 (N_2900,N_2745,N_2664);
nor U2901 (N_2901,N_2668,N_2660);
nand U2902 (N_2902,N_2745,N_2754);
nand U2903 (N_2903,N_2629,N_2616);
and U2904 (N_2904,N_2726,N_2785);
and U2905 (N_2905,N_2775,N_2766);
and U2906 (N_2906,N_2718,N_2617);
and U2907 (N_2907,N_2640,N_2770);
and U2908 (N_2908,N_2637,N_2737);
nor U2909 (N_2909,N_2701,N_2628);
nand U2910 (N_2910,N_2695,N_2757);
and U2911 (N_2911,N_2634,N_2754);
and U2912 (N_2912,N_2682,N_2652);
and U2913 (N_2913,N_2690,N_2666);
or U2914 (N_2914,N_2627,N_2771);
xnor U2915 (N_2915,N_2707,N_2789);
nand U2916 (N_2916,N_2607,N_2672);
nor U2917 (N_2917,N_2737,N_2749);
nand U2918 (N_2918,N_2699,N_2721);
nor U2919 (N_2919,N_2725,N_2610);
nand U2920 (N_2920,N_2782,N_2629);
or U2921 (N_2921,N_2718,N_2687);
nor U2922 (N_2922,N_2725,N_2664);
nand U2923 (N_2923,N_2673,N_2706);
and U2924 (N_2924,N_2635,N_2755);
and U2925 (N_2925,N_2627,N_2622);
nor U2926 (N_2926,N_2765,N_2716);
nor U2927 (N_2927,N_2733,N_2785);
and U2928 (N_2928,N_2760,N_2709);
and U2929 (N_2929,N_2745,N_2708);
or U2930 (N_2930,N_2654,N_2732);
xor U2931 (N_2931,N_2756,N_2606);
and U2932 (N_2932,N_2632,N_2679);
nand U2933 (N_2933,N_2623,N_2626);
and U2934 (N_2934,N_2645,N_2661);
and U2935 (N_2935,N_2710,N_2709);
and U2936 (N_2936,N_2691,N_2656);
or U2937 (N_2937,N_2619,N_2753);
nand U2938 (N_2938,N_2639,N_2706);
and U2939 (N_2939,N_2666,N_2673);
or U2940 (N_2940,N_2606,N_2769);
or U2941 (N_2941,N_2729,N_2739);
and U2942 (N_2942,N_2611,N_2711);
or U2943 (N_2943,N_2799,N_2684);
xor U2944 (N_2944,N_2712,N_2665);
or U2945 (N_2945,N_2793,N_2709);
or U2946 (N_2946,N_2608,N_2615);
or U2947 (N_2947,N_2763,N_2626);
and U2948 (N_2948,N_2732,N_2634);
or U2949 (N_2949,N_2764,N_2795);
or U2950 (N_2950,N_2602,N_2651);
and U2951 (N_2951,N_2617,N_2628);
nand U2952 (N_2952,N_2750,N_2666);
or U2953 (N_2953,N_2713,N_2732);
nor U2954 (N_2954,N_2604,N_2738);
or U2955 (N_2955,N_2661,N_2655);
nand U2956 (N_2956,N_2638,N_2731);
or U2957 (N_2957,N_2684,N_2705);
nand U2958 (N_2958,N_2715,N_2620);
and U2959 (N_2959,N_2621,N_2680);
nor U2960 (N_2960,N_2644,N_2716);
nand U2961 (N_2961,N_2602,N_2731);
nand U2962 (N_2962,N_2712,N_2760);
nor U2963 (N_2963,N_2717,N_2698);
and U2964 (N_2964,N_2706,N_2672);
or U2965 (N_2965,N_2797,N_2669);
nor U2966 (N_2966,N_2718,N_2629);
nor U2967 (N_2967,N_2664,N_2774);
nand U2968 (N_2968,N_2752,N_2672);
nor U2969 (N_2969,N_2690,N_2732);
and U2970 (N_2970,N_2793,N_2688);
and U2971 (N_2971,N_2799,N_2716);
or U2972 (N_2972,N_2776,N_2618);
nor U2973 (N_2973,N_2784,N_2673);
and U2974 (N_2974,N_2639,N_2698);
nand U2975 (N_2975,N_2759,N_2640);
nand U2976 (N_2976,N_2670,N_2642);
nand U2977 (N_2977,N_2704,N_2619);
nand U2978 (N_2978,N_2611,N_2799);
or U2979 (N_2979,N_2727,N_2695);
nor U2980 (N_2980,N_2761,N_2658);
and U2981 (N_2981,N_2793,N_2762);
or U2982 (N_2982,N_2660,N_2688);
or U2983 (N_2983,N_2684,N_2633);
nand U2984 (N_2984,N_2765,N_2618);
or U2985 (N_2985,N_2693,N_2740);
nand U2986 (N_2986,N_2688,N_2725);
or U2987 (N_2987,N_2704,N_2680);
or U2988 (N_2988,N_2716,N_2608);
and U2989 (N_2989,N_2717,N_2793);
or U2990 (N_2990,N_2686,N_2786);
or U2991 (N_2991,N_2670,N_2688);
nand U2992 (N_2992,N_2722,N_2730);
and U2993 (N_2993,N_2674,N_2638);
xnor U2994 (N_2994,N_2674,N_2745);
or U2995 (N_2995,N_2686,N_2773);
nor U2996 (N_2996,N_2658,N_2660);
or U2997 (N_2997,N_2783,N_2715);
nand U2998 (N_2998,N_2646,N_2757);
nor U2999 (N_2999,N_2749,N_2605);
nand U3000 (N_3000,N_2929,N_2949);
nand U3001 (N_3001,N_2977,N_2881);
and U3002 (N_3002,N_2850,N_2854);
nand U3003 (N_3003,N_2955,N_2825);
and U3004 (N_3004,N_2951,N_2991);
and U3005 (N_3005,N_2865,N_2911);
and U3006 (N_3006,N_2832,N_2873);
and U3007 (N_3007,N_2844,N_2984);
or U3008 (N_3008,N_2979,N_2805);
or U3009 (N_3009,N_2941,N_2950);
nand U3010 (N_3010,N_2961,N_2834);
nand U3011 (N_3011,N_2824,N_2947);
nor U3012 (N_3012,N_2988,N_2922);
nand U3013 (N_3013,N_2811,N_2924);
nor U3014 (N_3014,N_2931,N_2934);
nand U3015 (N_3015,N_2875,N_2972);
nand U3016 (N_3016,N_2957,N_2859);
nand U3017 (N_3017,N_2887,N_2855);
or U3018 (N_3018,N_2997,N_2851);
and U3019 (N_3019,N_2915,N_2971);
or U3020 (N_3020,N_2866,N_2815);
nand U3021 (N_3021,N_2898,N_2963);
or U3022 (N_3022,N_2993,N_2920);
nor U3023 (N_3023,N_2877,N_2980);
or U3024 (N_3024,N_2831,N_2982);
and U3025 (N_3025,N_2871,N_2852);
nand U3026 (N_3026,N_2846,N_2917);
nand U3027 (N_3027,N_2822,N_2912);
or U3028 (N_3028,N_2879,N_2999);
and U3029 (N_3029,N_2944,N_2989);
nand U3030 (N_3030,N_2974,N_2816);
nor U3031 (N_3031,N_2807,N_2861);
or U3032 (N_3032,N_2841,N_2857);
nor U3033 (N_3033,N_2826,N_2833);
or U3034 (N_3034,N_2975,N_2820);
or U3035 (N_3035,N_2876,N_2998);
xor U3036 (N_3036,N_2830,N_2872);
or U3037 (N_3037,N_2995,N_2933);
xnor U3038 (N_3038,N_2870,N_2883);
or U3039 (N_3039,N_2835,N_2894);
nand U3040 (N_3040,N_2829,N_2899);
and U3041 (N_3041,N_2992,N_2897);
nor U3042 (N_3042,N_2886,N_2940);
and U3043 (N_3043,N_2891,N_2839);
or U3044 (N_3044,N_2869,N_2828);
or U3045 (N_3045,N_2808,N_2803);
nor U3046 (N_3046,N_2942,N_2985);
and U3047 (N_3047,N_2962,N_2878);
nor U3048 (N_3048,N_2904,N_2823);
nor U3049 (N_3049,N_2845,N_2827);
nor U3050 (N_3050,N_2862,N_2976);
or U3051 (N_3051,N_2867,N_2840);
or U3052 (N_3052,N_2914,N_2892);
or U3053 (N_3053,N_2900,N_2801);
nor U3054 (N_3054,N_2952,N_2968);
nand U3055 (N_3055,N_2916,N_2885);
nand U3056 (N_3056,N_2946,N_2960);
nand U3057 (N_3057,N_2923,N_2802);
nor U3058 (N_3058,N_2893,N_2842);
or U3059 (N_3059,N_2965,N_2927);
or U3060 (N_3060,N_2838,N_2938);
and U3061 (N_3061,N_2928,N_2956);
or U3062 (N_3062,N_2905,N_2800);
xor U3063 (N_3063,N_2804,N_2856);
nor U3064 (N_3064,N_2909,N_2868);
or U3065 (N_3065,N_2945,N_2814);
and U3066 (N_3066,N_2990,N_2902);
and U3067 (N_3067,N_2994,N_2849);
nor U3068 (N_3068,N_2864,N_2903);
and U3069 (N_3069,N_2848,N_2809);
nand U3070 (N_3070,N_2843,N_2847);
and U3071 (N_3071,N_2821,N_2926);
or U3072 (N_3072,N_2853,N_2958);
nand U3073 (N_3073,N_2987,N_2930);
nand U3074 (N_3074,N_2889,N_2863);
or U3075 (N_3075,N_2880,N_2817);
or U3076 (N_3076,N_2978,N_2890);
or U3077 (N_3077,N_2981,N_2818);
nand U3078 (N_3078,N_2937,N_2964);
nand U3079 (N_3079,N_2954,N_2939);
and U3080 (N_3080,N_2906,N_2959);
nor U3081 (N_3081,N_2925,N_2948);
and U3082 (N_3082,N_2969,N_2935);
or U3083 (N_3083,N_2943,N_2812);
and U3084 (N_3084,N_2874,N_2966);
nand U3085 (N_3085,N_2836,N_2996);
nor U3086 (N_3086,N_2936,N_2970);
nand U3087 (N_3087,N_2813,N_2913);
nor U3088 (N_3088,N_2810,N_2806);
nand U3089 (N_3089,N_2858,N_2901);
and U3090 (N_3090,N_2918,N_2908);
nand U3091 (N_3091,N_2837,N_2860);
and U3092 (N_3092,N_2921,N_2983);
nand U3093 (N_3093,N_2973,N_2888);
or U3094 (N_3094,N_2819,N_2932);
or U3095 (N_3095,N_2895,N_2882);
and U3096 (N_3096,N_2884,N_2919);
or U3097 (N_3097,N_2896,N_2967);
nand U3098 (N_3098,N_2910,N_2986);
nand U3099 (N_3099,N_2907,N_2953);
nor U3100 (N_3100,N_2874,N_2928);
and U3101 (N_3101,N_2810,N_2908);
or U3102 (N_3102,N_2876,N_2971);
or U3103 (N_3103,N_2940,N_2972);
nand U3104 (N_3104,N_2859,N_2856);
nor U3105 (N_3105,N_2907,N_2898);
or U3106 (N_3106,N_2859,N_2912);
nand U3107 (N_3107,N_2995,N_2872);
nor U3108 (N_3108,N_2991,N_2843);
nand U3109 (N_3109,N_2980,N_2947);
nor U3110 (N_3110,N_2876,N_2822);
and U3111 (N_3111,N_2833,N_2976);
and U3112 (N_3112,N_2991,N_2846);
and U3113 (N_3113,N_2922,N_2843);
nand U3114 (N_3114,N_2924,N_2846);
nand U3115 (N_3115,N_2950,N_2951);
nand U3116 (N_3116,N_2974,N_2882);
nand U3117 (N_3117,N_2928,N_2826);
or U3118 (N_3118,N_2885,N_2878);
nor U3119 (N_3119,N_2912,N_2845);
nand U3120 (N_3120,N_2869,N_2977);
nor U3121 (N_3121,N_2886,N_2859);
and U3122 (N_3122,N_2861,N_2867);
and U3123 (N_3123,N_2813,N_2914);
nand U3124 (N_3124,N_2887,N_2924);
or U3125 (N_3125,N_2840,N_2983);
and U3126 (N_3126,N_2985,N_2965);
or U3127 (N_3127,N_2835,N_2833);
and U3128 (N_3128,N_2820,N_2894);
nand U3129 (N_3129,N_2878,N_2863);
and U3130 (N_3130,N_2954,N_2876);
nand U3131 (N_3131,N_2928,N_2922);
nand U3132 (N_3132,N_2863,N_2979);
and U3133 (N_3133,N_2817,N_2906);
nor U3134 (N_3134,N_2904,N_2865);
nor U3135 (N_3135,N_2861,N_2827);
or U3136 (N_3136,N_2926,N_2913);
nand U3137 (N_3137,N_2982,N_2946);
nand U3138 (N_3138,N_2807,N_2958);
nand U3139 (N_3139,N_2833,N_2988);
nand U3140 (N_3140,N_2979,N_2896);
nand U3141 (N_3141,N_2998,N_2809);
or U3142 (N_3142,N_2802,N_2822);
and U3143 (N_3143,N_2980,N_2862);
nor U3144 (N_3144,N_2807,N_2801);
nor U3145 (N_3145,N_2870,N_2897);
and U3146 (N_3146,N_2999,N_2906);
nor U3147 (N_3147,N_2997,N_2875);
and U3148 (N_3148,N_2899,N_2813);
nor U3149 (N_3149,N_2869,N_2987);
nor U3150 (N_3150,N_2848,N_2841);
nor U3151 (N_3151,N_2945,N_2861);
or U3152 (N_3152,N_2912,N_2820);
or U3153 (N_3153,N_2970,N_2980);
and U3154 (N_3154,N_2932,N_2999);
or U3155 (N_3155,N_2958,N_2912);
and U3156 (N_3156,N_2874,N_2896);
and U3157 (N_3157,N_2898,N_2919);
nor U3158 (N_3158,N_2830,N_2865);
and U3159 (N_3159,N_2911,N_2986);
nor U3160 (N_3160,N_2896,N_2921);
and U3161 (N_3161,N_2866,N_2975);
and U3162 (N_3162,N_2953,N_2809);
and U3163 (N_3163,N_2888,N_2994);
nor U3164 (N_3164,N_2953,N_2861);
nor U3165 (N_3165,N_2923,N_2846);
and U3166 (N_3166,N_2834,N_2836);
nor U3167 (N_3167,N_2872,N_2999);
nand U3168 (N_3168,N_2884,N_2883);
and U3169 (N_3169,N_2813,N_2891);
nand U3170 (N_3170,N_2907,N_2860);
or U3171 (N_3171,N_2874,N_2981);
and U3172 (N_3172,N_2908,N_2813);
and U3173 (N_3173,N_2846,N_2942);
nor U3174 (N_3174,N_2951,N_2870);
and U3175 (N_3175,N_2885,N_2970);
and U3176 (N_3176,N_2915,N_2972);
or U3177 (N_3177,N_2888,N_2826);
or U3178 (N_3178,N_2967,N_2976);
nand U3179 (N_3179,N_2946,N_2834);
nand U3180 (N_3180,N_2993,N_2858);
nand U3181 (N_3181,N_2967,N_2999);
and U3182 (N_3182,N_2888,N_2975);
nor U3183 (N_3183,N_2868,N_2930);
nor U3184 (N_3184,N_2974,N_2963);
and U3185 (N_3185,N_2932,N_2938);
nor U3186 (N_3186,N_2913,N_2968);
or U3187 (N_3187,N_2956,N_2870);
and U3188 (N_3188,N_2800,N_2864);
and U3189 (N_3189,N_2993,N_2811);
nor U3190 (N_3190,N_2877,N_2905);
and U3191 (N_3191,N_2828,N_2946);
nand U3192 (N_3192,N_2942,N_2844);
or U3193 (N_3193,N_2992,N_2987);
nor U3194 (N_3194,N_2831,N_2932);
or U3195 (N_3195,N_2856,N_2972);
or U3196 (N_3196,N_2950,N_2952);
nor U3197 (N_3197,N_2920,N_2815);
nand U3198 (N_3198,N_2946,N_2818);
or U3199 (N_3199,N_2945,N_2862);
or U3200 (N_3200,N_3068,N_3014);
nor U3201 (N_3201,N_3029,N_3084);
nand U3202 (N_3202,N_3158,N_3108);
and U3203 (N_3203,N_3182,N_3153);
and U3204 (N_3204,N_3168,N_3189);
nand U3205 (N_3205,N_3069,N_3046);
nor U3206 (N_3206,N_3144,N_3131);
nor U3207 (N_3207,N_3083,N_3129);
and U3208 (N_3208,N_3071,N_3113);
xor U3209 (N_3209,N_3097,N_3141);
and U3210 (N_3210,N_3171,N_3162);
and U3211 (N_3211,N_3061,N_3054);
and U3212 (N_3212,N_3124,N_3198);
nand U3213 (N_3213,N_3098,N_3107);
nand U3214 (N_3214,N_3056,N_3018);
nor U3215 (N_3215,N_3127,N_3121);
nand U3216 (N_3216,N_3125,N_3183);
or U3217 (N_3217,N_3042,N_3188);
and U3218 (N_3218,N_3157,N_3166);
and U3219 (N_3219,N_3092,N_3004);
or U3220 (N_3220,N_3185,N_3101);
or U3221 (N_3221,N_3077,N_3074);
and U3222 (N_3222,N_3050,N_3000);
nor U3223 (N_3223,N_3133,N_3102);
or U3224 (N_3224,N_3019,N_3040);
or U3225 (N_3225,N_3152,N_3106);
nor U3226 (N_3226,N_3167,N_3063);
or U3227 (N_3227,N_3088,N_3138);
or U3228 (N_3228,N_3184,N_3159);
or U3229 (N_3229,N_3066,N_3165);
nor U3230 (N_3230,N_3080,N_3156);
nand U3231 (N_3231,N_3003,N_3137);
nand U3232 (N_3232,N_3006,N_3044);
or U3233 (N_3233,N_3199,N_3030);
and U3234 (N_3234,N_3049,N_3053);
nor U3235 (N_3235,N_3142,N_3007);
and U3236 (N_3236,N_3015,N_3169);
nor U3237 (N_3237,N_3145,N_3178);
and U3238 (N_3238,N_3120,N_3076);
and U3239 (N_3239,N_3024,N_3073);
xor U3240 (N_3240,N_3013,N_3005);
or U3241 (N_3241,N_3174,N_3010);
nand U3242 (N_3242,N_3051,N_3105);
nor U3243 (N_3243,N_3196,N_3177);
and U3244 (N_3244,N_3002,N_3012);
and U3245 (N_3245,N_3147,N_3082);
nand U3246 (N_3246,N_3136,N_3031);
nand U3247 (N_3247,N_3059,N_3095);
and U3248 (N_3248,N_3170,N_3028);
nor U3249 (N_3249,N_3027,N_3067);
nor U3250 (N_3250,N_3037,N_3026);
nand U3251 (N_3251,N_3187,N_3192);
or U3252 (N_3252,N_3060,N_3111);
nand U3253 (N_3253,N_3135,N_3081);
or U3254 (N_3254,N_3052,N_3043);
or U3255 (N_3255,N_3047,N_3191);
nand U3256 (N_3256,N_3070,N_3093);
nor U3257 (N_3257,N_3173,N_3181);
or U3258 (N_3258,N_3079,N_3020);
or U3259 (N_3259,N_3130,N_3195);
and U3260 (N_3260,N_3033,N_3115);
nor U3261 (N_3261,N_3087,N_3036);
or U3262 (N_3262,N_3186,N_3001);
nand U3263 (N_3263,N_3175,N_3025);
nor U3264 (N_3264,N_3114,N_3140);
nand U3265 (N_3265,N_3134,N_3104);
nor U3266 (N_3266,N_3062,N_3151);
and U3267 (N_3267,N_3154,N_3039);
or U3268 (N_3268,N_3176,N_3022);
or U3269 (N_3269,N_3055,N_3109);
and U3270 (N_3270,N_3096,N_3072);
nand U3271 (N_3271,N_3180,N_3090);
nand U3272 (N_3272,N_3146,N_3112);
nor U3273 (N_3273,N_3190,N_3058);
nor U3274 (N_3274,N_3032,N_3078);
nor U3275 (N_3275,N_3038,N_3197);
and U3276 (N_3276,N_3122,N_3123);
nand U3277 (N_3277,N_3160,N_3132);
nand U3278 (N_3278,N_3091,N_3110);
and U3279 (N_3279,N_3094,N_3041);
or U3280 (N_3280,N_3065,N_3048);
and U3281 (N_3281,N_3089,N_3117);
or U3282 (N_3282,N_3021,N_3099);
and U3283 (N_3283,N_3100,N_3057);
nand U3284 (N_3284,N_3034,N_3148);
nand U3285 (N_3285,N_3119,N_3116);
and U3286 (N_3286,N_3164,N_3193);
and U3287 (N_3287,N_3008,N_3128);
nand U3288 (N_3288,N_3179,N_3126);
nor U3289 (N_3289,N_3161,N_3118);
nand U3290 (N_3290,N_3139,N_3163);
nand U3291 (N_3291,N_3064,N_3172);
or U3292 (N_3292,N_3016,N_3035);
nor U3293 (N_3293,N_3143,N_3150);
nand U3294 (N_3294,N_3086,N_3085);
and U3295 (N_3295,N_3155,N_3023);
or U3296 (N_3296,N_3194,N_3103);
nand U3297 (N_3297,N_3009,N_3075);
nand U3298 (N_3298,N_3045,N_3149);
nand U3299 (N_3299,N_3017,N_3011);
or U3300 (N_3300,N_3195,N_3156);
or U3301 (N_3301,N_3189,N_3084);
or U3302 (N_3302,N_3028,N_3057);
and U3303 (N_3303,N_3164,N_3066);
and U3304 (N_3304,N_3099,N_3058);
or U3305 (N_3305,N_3178,N_3139);
nand U3306 (N_3306,N_3144,N_3023);
nor U3307 (N_3307,N_3126,N_3040);
nor U3308 (N_3308,N_3090,N_3118);
and U3309 (N_3309,N_3157,N_3173);
nor U3310 (N_3310,N_3080,N_3133);
nor U3311 (N_3311,N_3102,N_3197);
nor U3312 (N_3312,N_3016,N_3077);
nor U3313 (N_3313,N_3061,N_3123);
nand U3314 (N_3314,N_3026,N_3077);
nand U3315 (N_3315,N_3136,N_3143);
or U3316 (N_3316,N_3017,N_3039);
nor U3317 (N_3317,N_3108,N_3022);
nand U3318 (N_3318,N_3138,N_3141);
nor U3319 (N_3319,N_3027,N_3009);
nand U3320 (N_3320,N_3097,N_3134);
and U3321 (N_3321,N_3014,N_3001);
and U3322 (N_3322,N_3093,N_3103);
nor U3323 (N_3323,N_3094,N_3172);
and U3324 (N_3324,N_3010,N_3138);
and U3325 (N_3325,N_3156,N_3108);
or U3326 (N_3326,N_3085,N_3040);
or U3327 (N_3327,N_3002,N_3166);
and U3328 (N_3328,N_3046,N_3113);
or U3329 (N_3329,N_3079,N_3025);
and U3330 (N_3330,N_3062,N_3073);
nand U3331 (N_3331,N_3153,N_3150);
and U3332 (N_3332,N_3055,N_3127);
nor U3333 (N_3333,N_3191,N_3046);
and U3334 (N_3334,N_3005,N_3116);
nand U3335 (N_3335,N_3153,N_3009);
and U3336 (N_3336,N_3035,N_3181);
and U3337 (N_3337,N_3162,N_3049);
nand U3338 (N_3338,N_3093,N_3173);
and U3339 (N_3339,N_3176,N_3159);
nor U3340 (N_3340,N_3036,N_3060);
nor U3341 (N_3341,N_3144,N_3124);
and U3342 (N_3342,N_3072,N_3053);
nor U3343 (N_3343,N_3171,N_3038);
nand U3344 (N_3344,N_3008,N_3169);
nand U3345 (N_3345,N_3116,N_3014);
nor U3346 (N_3346,N_3173,N_3074);
or U3347 (N_3347,N_3154,N_3147);
nand U3348 (N_3348,N_3154,N_3094);
or U3349 (N_3349,N_3035,N_3161);
or U3350 (N_3350,N_3128,N_3119);
xor U3351 (N_3351,N_3132,N_3061);
nand U3352 (N_3352,N_3132,N_3075);
nand U3353 (N_3353,N_3087,N_3124);
and U3354 (N_3354,N_3170,N_3179);
and U3355 (N_3355,N_3022,N_3185);
nor U3356 (N_3356,N_3150,N_3047);
nand U3357 (N_3357,N_3102,N_3155);
and U3358 (N_3358,N_3169,N_3002);
nor U3359 (N_3359,N_3130,N_3165);
xor U3360 (N_3360,N_3036,N_3169);
and U3361 (N_3361,N_3116,N_3101);
nor U3362 (N_3362,N_3180,N_3094);
nor U3363 (N_3363,N_3016,N_3083);
nand U3364 (N_3364,N_3079,N_3159);
nor U3365 (N_3365,N_3144,N_3044);
and U3366 (N_3366,N_3184,N_3048);
and U3367 (N_3367,N_3075,N_3015);
nand U3368 (N_3368,N_3057,N_3195);
and U3369 (N_3369,N_3157,N_3190);
nand U3370 (N_3370,N_3144,N_3086);
or U3371 (N_3371,N_3112,N_3080);
or U3372 (N_3372,N_3028,N_3105);
or U3373 (N_3373,N_3105,N_3073);
nand U3374 (N_3374,N_3003,N_3126);
nor U3375 (N_3375,N_3165,N_3047);
and U3376 (N_3376,N_3187,N_3035);
and U3377 (N_3377,N_3115,N_3031);
nor U3378 (N_3378,N_3065,N_3075);
nor U3379 (N_3379,N_3162,N_3113);
nor U3380 (N_3380,N_3194,N_3156);
and U3381 (N_3381,N_3127,N_3182);
nand U3382 (N_3382,N_3002,N_3172);
nand U3383 (N_3383,N_3195,N_3121);
and U3384 (N_3384,N_3018,N_3078);
nand U3385 (N_3385,N_3180,N_3196);
and U3386 (N_3386,N_3161,N_3081);
and U3387 (N_3387,N_3196,N_3116);
and U3388 (N_3388,N_3088,N_3108);
and U3389 (N_3389,N_3174,N_3052);
or U3390 (N_3390,N_3029,N_3142);
nor U3391 (N_3391,N_3092,N_3019);
xnor U3392 (N_3392,N_3144,N_3039);
nand U3393 (N_3393,N_3170,N_3120);
nand U3394 (N_3394,N_3126,N_3014);
nand U3395 (N_3395,N_3116,N_3175);
nand U3396 (N_3396,N_3124,N_3030);
nand U3397 (N_3397,N_3050,N_3176);
nand U3398 (N_3398,N_3186,N_3160);
nand U3399 (N_3399,N_3126,N_3198);
and U3400 (N_3400,N_3311,N_3392);
or U3401 (N_3401,N_3396,N_3322);
nand U3402 (N_3402,N_3289,N_3275);
or U3403 (N_3403,N_3266,N_3298);
xor U3404 (N_3404,N_3252,N_3319);
or U3405 (N_3405,N_3350,N_3251);
and U3406 (N_3406,N_3358,N_3265);
and U3407 (N_3407,N_3215,N_3260);
or U3408 (N_3408,N_3329,N_3205);
or U3409 (N_3409,N_3206,N_3390);
nand U3410 (N_3410,N_3303,N_3352);
nor U3411 (N_3411,N_3310,N_3236);
nand U3412 (N_3412,N_3344,N_3321);
nand U3413 (N_3413,N_3226,N_3261);
nand U3414 (N_3414,N_3225,N_3375);
nand U3415 (N_3415,N_3294,N_3351);
nand U3416 (N_3416,N_3354,N_3302);
nand U3417 (N_3417,N_3247,N_3280);
and U3418 (N_3418,N_3283,N_3397);
nor U3419 (N_3419,N_3307,N_3301);
nor U3420 (N_3420,N_3245,N_3361);
and U3421 (N_3421,N_3279,N_3372);
and U3422 (N_3422,N_3254,N_3389);
nand U3423 (N_3423,N_3258,N_3315);
nand U3424 (N_3424,N_3250,N_3272);
nor U3425 (N_3425,N_3367,N_3211);
nor U3426 (N_3426,N_3316,N_3263);
and U3427 (N_3427,N_3274,N_3218);
or U3428 (N_3428,N_3239,N_3388);
or U3429 (N_3429,N_3207,N_3234);
nand U3430 (N_3430,N_3297,N_3393);
nand U3431 (N_3431,N_3328,N_3314);
nand U3432 (N_3432,N_3231,N_3355);
nand U3433 (N_3433,N_3313,N_3208);
nor U3434 (N_3434,N_3334,N_3256);
nand U3435 (N_3435,N_3369,N_3336);
nand U3436 (N_3436,N_3229,N_3366);
or U3437 (N_3437,N_3235,N_3217);
nor U3438 (N_3438,N_3306,N_3379);
or U3439 (N_3439,N_3339,N_3230);
or U3440 (N_3440,N_3359,N_3320);
or U3441 (N_3441,N_3202,N_3399);
nor U3442 (N_3442,N_3387,N_3305);
or U3443 (N_3443,N_3349,N_3284);
nor U3444 (N_3444,N_3377,N_3323);
and U3445 (N_3445,N_3296,N_3395);
and U3446 (N_3446,N_3286,N_3368);
and U3447 (N_3447,N_3227,N_3295);
nand U3448 (N_3448,N_3278,N_3391);
nor U3449 (N_3449,N_3385,N_3337);
or U3450 (N_3450,N_3262,N_3242);
and U3451 (N_3451,N_3243,N_3380);
or U3452 (N_3452,N_3304,N_3222);
nand U3453 (N_3453,N_3267,N_3273);
and U3454 (N_3454,N_3212,N_3219);
or U3455 (N_3455,N_3257,N_3290);
nor U3456 (N_3456,N_3288,N_3210);
and U3457 (N_3457,N_3353,N_3214);
nor U3458 (N_3458,N_3382,N_3381);
and U3459 (N_3459,N_3348,N_3287);
nand U3460 (N_3460,N_3386,N_3356);
or U3461 (N_3461,N_3271,N_3233);
nor U3462 (N_3462,N_3221,N_3241);
or U3463 (N_3463,N_3340,N_3276);
and U3464 (N_3464,N_3220,N_3371);
or U3465 (N_3465,N_3364,N_3270);
and U3466 (N_3466,N_3333,N_3335);
or U3467 (N_3467,N_3378,N_3324);
and U3468 (N_3468,N_3384,N_3345);
nor U3469 (N_3469,N_3223,N_3255);
and U3470 (N_3470,N_3291,N_3376);
nor U3471 (N_3471,N_3201,N_3300);
nor U3472 (N_3472,N_3394,N_3332);
nor U3473 (N_3473,N_3268,N_3360);
nand U3474 (N_3474,N_3216,N_3326);
nand U3475 (N_3475,N_3281,N_3325);
and U3476 (N_3476,N_3338,N_3240);
or U3477 (N_3477,N_3347,N_3373);
or U3478 (N_3478,N_3285,N_3357);
and U3479 (N_3479,N_3249,N_3228);
nand U3480 (N_3480,N_3312,N_3200);
nand U3481 (N_3481,N_3213,N_3398);
nor U3482 (N_3482,N_3330,N_3342);
nand U3483 (N_3483,N_3374,N_3264);
and U3484 (N_3484,N_3253,N_3317);
nor U3485 (N_3485,N_3269,N_3308);
nand U3486 (N_3486,N_3259,N_3299);
nand U3487 (N_3487,N_3232,N_3346);
nor U3488 (N_3488,N_3209,N_3246);
and U3489 (N_3489,N_3203,N_3383);
and U3490 (N_3490,N_3237,N_3309);
nor U3491 (N_3491,N_3248,N_3204);
xnor U3492 (N_3492,N_3327,N_3224);
and U3493 (N_3493,N_3293,N_3370);
or U3494 (N_3494,N_3362,N_3365);
and U3495 (N_3495,N_3331,N_3363);
nand U3496 (N_3496,N_3244,N_3282);
and U3497 (N_3497,N_3292,N_3238);
nand U3498 (N_3498,N_3318,N_3277);
or U3499 (N_3499,N_3343,N_3341);
xor U3500 (N_3500,N_3267,N_3240);
or U3501 (N_3501,N_3357,N_3284);
or U3502 (N_3502,N_3382,N_3347);
and U3503 (N_3503,N_3260,N_3349);
or U3504 (N_3504,N_3345,N_3365);
and U3505 (N_3505,N_3254,N_3335);
or U3506 (N_3506,N_3352,N_3237);
and U3507 (N_3507,N_3226,N_3309);
xnor U3508 (N_3508,N_3244,N_3225);
and U3509 (N_3509,N_3218,N_3244);
xor U3510 (N_3510,N_3279,N_3355);
nor U3511 (N_3511,N_3348,N_3394);
nand U3512 (N_3512,N_3389,N_3242);
nor U3513 (N_3513,N_3237,N_3261);
nand U3514 (N_3514,N_3358,N_3259);
or U3515 (N_3515,N_3232,N_3337);
and U3516 (N_3516,N_3371,N_3281);
and U3517 (N_3517,N_3286,N_3328);
nor U3518 (N_3518,N_3307,N_3272);
and U3519 (N_3519,N_3204,N_3202);
nand U3520 (N_3520,N_3217,N_3269);
or U3521 (N_3521,N_3316,N_3313);
nand U3522 (N_3522,N_3345,N_3219);
nor U3523 (N_3523,N_3364,N_3294);
xor U3524 (N_3524,N_3243,N_3350);
nor U3525 (N_3525,N_3373,N_3377);
or U3526 (N_3526,N_3275,N_3262);
nor U3527 (N_3527,N_3201,N_3314);
or U3528 (N_3528,N_3203,N_3221);
or U3529 (N_3529,N_3243,N_3229);
or U3530 (N_3530,N_3334,N_3329);
nor U3531 (N_3531,N_3358,N_3291);
nor U3532 (N_3532,N_3313,N_3205);
nor U3533 (N_3533,N_3275,N_3369);
or U3534 (N_3534,N_3292,N_3390);
nor U3535 (N_3535,N_3242,N_3292);
or U3536 (N_3536,N_3375,N_3377);
or U3537 (N_3537,N_3218,N_3380);
nor U3538 (N_3538,N_3398,N_3375);
nand U3539 (N_3539,N_3250,N_3352);
nor U3540 (N_3540,N_3244,N_3332);
nor U3541 (N_3541,N_3275,N_3366);
nand U3542 (N_3542,N_3397,N_3358);
or U3543 (N_3543,N_3268,N_3208);
nor U3544 (N_3544,N_3244,N_3280);
nand U3545 (N_3545,N_3337,N_3230);
or U3546 (N_3546,N_3274,N_3336);
nor U3547 (N_3547,N_3312,N_3276);
nand U3548 (N_3548,N_3318,N_3307);
or U3549 (N_3549,N_3252,N_3285);
nor U3550 (N_3550,N_3251,N_3288);
nand U3551 (N_3551,N_3347,N_3264);
or U3552 (N_3552,N_3364,N_3303);
nor U3553 (N_3553,N_3291,N_3211);
nand U3554 (N_3554,N_3304,N_3289);
nor U3555 (N_3555,N_3278,N_3248);
and U3556 (N_3556,N_3369,N_3223);
or U3557 (N_3557,N_3316,N_3264);
nor U3558 (N_3558,N_3246,N_3211);
or U3559 (N_3559,N_3375,N_3378);
or U3560 (N_3560,N_3321,N_3288);
nand U3561 (N_3561,N_3377,N_3211);
or U3562 (N_3562,N_3253,N_3346);
nor U3563 (N_3563,N_3250,N_3234);
and U3564 (N_3564,N_3230,N_3225);
nand U3565 (N_3565,N_3288,N_3325);
and U3566 (N_3566,N_3377,N_3210);
nand U3567 (N_3567,N_3287,N_3247);
and U3568 (N_3568,N_3354,N_3256);
or U3569 (N_3569,N_3342,N_3264);
and U3570 (N_3570,N_3340,N_3214);
or U3571 (N_3571,N_3334,N_3399);
nor U3572 (N_3572,N_3283,N_3311);
xnor U3573 (N_3573,N_3214,N_3267);
nand U3574 (N_3574,N_3333,N_3363);
and U3575 (N_3575,N_3284,N_3258);
nand U3576 (N_3576,N_3365,N_3335);
nand U3577 (N_3577,N_3385,N_3390);
xor U3578 (N_3578,N_3343,N_3226);
nand U3579 (N_3579,N_3266,N_3230);
nor U3580 (N_3580,N_3313,N_3203);
and U3581 (N_3581,N_3291,N_3250);
nor U3582 (N_3582,N_3272,N_3213);
nand U3583 (N_3583,N_3328,N_3355);
nand U3584 (N_3584,N_3257,N_3262);
or U3585 (N_3585,N_3304,N_3399);
and U3586 (N_3586,N_3268,N_3381);
and U3587 (N_3587,N_3215,N_3236);
and U3588 (N_3588,N_3321,N_3307);
and U3589 (N_3589,N_3305,N_3254);
nor U3590 (N_3590,N_3278,N_3265);
or U3591 (N_3591,N_3263,N_3304);
nor U3592 (N_3592,N_3338,N_3391);
and U3593 (N_3593,N_3265,N_3370);
or U3594 (N_3594,N_3237,N_3225);
nor U3595 (N_3595,N_3291,N_3229);
and U3596 (N_3596,N_3319,N_3363);
nand U3597 (N_3597,N_3343,N_3213);
nand U3598 (N_3598,N_3346,N_3231);
and U3599 (N_3599,N_3230,N_3250);
nand U3600 (N_3600,N_3535,N_3515);
and U3601 (N_3601,N_3520,N_3476);
or U3602 (N_3602,N_3447,N_3564);
nand U3603 (N_3603,N_3433,N_3531);
nand U3604 (N_3604,N_3415,N_3582);
nand U3605 (N_3605,N_3548,N_3420);
xnor U3606 (N_3606,N_3454,N_3424);
and U3607 (N_3607,N_3426,N_3563);
nand U3608 (N_3608,N_3503,N_3525);
nand U3609 (N_3609,N_3423,N_3498);
nand U3610 (N_3610,N_3436,N_3590);
or U3611 (N_3611,N_3522,N_3524);
and U3612 (N_3612,N_3443,N_3510);
or U3613 (N_3613,N_3560,N_3591);
xnor U3614 (N_3614,N_3541,N_3592);
nor U3615 (N_3615,N_3407,N_3465);
nor U3616 (N_3616,N_3400,N_3562);
or U3617 (N_3617,N_3506,N_3568);
or U3618 (N_3618,N_3473,N_3482);
nand U3619 (N_3619,N_3526,N_3406);
nand U3620 (N_3620,N_3478,N_3460);
nor U3621 (N_3621,N_3561,N_3480);
and U3622 (N_3622,N_3446,N_3431);
nand U3623 (N_3623,N_3428,N_3581);
nand U3624 (N_3624,N_3502,N_3444);
and U3625 (N_3625,N_3457,N_3501);
nand U3626 (N_3626,N_3536,N_3599);
or U3627 (N_3627,N_3507,N_3516);
or U3628 (N_3628,N_3519,N_3416);
nor U3629 (N_3629,N_3418,N_3573);
or U3630 (N_3630,N_3453,N_3570);
and U3631 (N_3631,N_3499,N_3435);
nand U3632 (N_3632,N_3569,N_3451);
and U3633 (N_3633,N_3505,N_3471);
nor U3634 (N_3634,N_3412,N_3544);
or U3635 (N_3635,N_3538,N_3421);
nor U3636 (N_3636,N_3487,N_3546);
and U3637 (N_3637,N_3558,N_3474);
xor U3638 (N_3638,N_3529,N_3575);
and U3639 (N_3639,N_3540,N_3484);
nor U3640 (N_3640,N_3442,N_3477);
nor U3641 (N_3641,N_3517,N_3437);
nor U3642 (N_3642,N_3513,N_3528);
nand U3643 (N_3643,N_3448,N_3411);
and U3644 (N_3644,N_3410,N_3583);
and U3645 (N_3645,N_3547,N_3508);
nor U3646 (N_3646,N_3588,N_3597);
and U3647 (N_3647,N_3596,N_3533);
nor U3648 (N_3648,N_3552,N_3488);
nor U3649 (N_3649,N_3574,N_3557);
nand U3650 (N_3650,N_3509,N_3419);
nand U3651 (N_3651,N_3464,N_3537);
nor U3652 (N_3652,N_3438,N_3593);
nor U3653 (N_3653,N_3427,N_3475);
nor U3654 (N_3654,N_3550,N_3572);
nand U3655 (N_3655,N_3408,N_3527);
or U3656 (N_3656,N_3492,N_3585);
or U3657 (N_3657,N_3579,N_3430);
nor U3658 (N_3658,N_3532,N_3469);
nor U3659 (N_3659,N_3461,N_3425);
nor U3660 (N_3660,N_3402,N_3576);
nor U3661 (N_3661,N_3458,N_3584);
and U3662 (N_3662,N_3518,N_3405);
nand U3663 (N_3663,N_3455,N_3472);
nand U3664 (N_3664,N_3459,N_3449);
or U3665 (N_3665,N_3463,N_3494);
nand U3666 (N_3666,N_3422,N_3439);
or U3667 (N_3667,N_3468,N_3456);
and U3668 (N_3668,N_3489,N_3594);
and U3669 (N_3669,N_3504,N_3493);
nand U3670 (N_3670,N_3496,N_3445);
and U3671 (N_3671,N_3555,N_3495);
nand U3672 (N_3672,N_3556,N_3434);
xor U3673 (N_3673,N_3466,N_3490);
nor U3674 (N_3674,N_3414,N_3497);
nand U3675 (N_3675,N_3566,N_3491);
nor U3676 (N_3676,N_3589,N_3598);
nor U3677 (N_3677,N_3565,N_3543);
and U3678 (N_3678,N_3530,N_3432);
xor U3679 (N_3679,N_3417,N_3441);
and U3680 (N_3680,N_3413,N_3559);
and U3681 (N_3681,N_3580,N_3523);
nor U3682 (N_3682,N_3554,N_3539);
nand U3683 (N_3683,N_3545,N_3440);
nand U3684 (N_3684,N_3595,N_3462);
nor U3685 (N_3685,N_3470,N_3534);
nand U3686 (N_3686,N_3514,N_3500);
and U3687 (N_3687,N_3429,N_3404);
nand U3688 (N_3688,N_3450,N_3549);
or U3689 (N_3689,N_3401,N_3542);
and U3690 (N_3690,N_3578,N_3553);
nand U3691 (N_3691,N_3567,N_3577);
nand U3692 (N_3692,N_3486,N_3571);
or U3693 (N_3693,N_3479,N_3481);
nor U3694 (N_3694,N_3485,N_3586);
nand U3695 (N_3695,N_3551,N_3587);
or U3696 (N_3696,N_3521,N_3452);
and U3697 (N_3697,N_3409,N_3483);
nand U3698 (N_3698,N_3512,N_3511);
and U3699 (N_3699,N_3467,N_3403);
xnor U3700 (N_3700,N_3400,N_3481);
nand U3701 (N_3701,N_3489,N_3524);
nand U3702 (N_3702,N_3533,N_3431);
and U3703 (N_3703,N_3569,N_3435);
and U3704 (N_3704,N_3516,N_3473);
nor U3705 (N_3705,N_3576,N_3410);
nor U3706 (N_3706,N_3441,N_3574);
nor U3707 (N_3707,N_3457,N_3537);
nor U3708 (N_3708,N_3523,N_3551);
nor U3709 (N_3709,N_3430,N_3427);
nand U3710 (N_3710,N_3559,N_3480);
nand U3711 (N_3711,N_3439,N_3414);
nand U3712 (N_3712,N_3489,N_3550);
nor U3713 (N_3713,N_3411,N_3513);
or U3714 (N_3714,N_3489,N_3436);
or U3715 (N_3715,N_3407,N_3477);
nand U3716 (N_3716,N_3422,N_3483);
nand U3717 (N_3717,N_3528,N_3408);
nand U3718 (N_3718,N_3445,N_3577);
nand U3719 (N_3719,N_3593,N_3524);
nor U3720 (N_3720,N_3457,N_3498);
and U3721 (N_3721,N_3453,N_3403);
or U3722 (N_3722,N_3537,N_3519);
and U3723 (N_3723,N_3456,N_3478);
and U3724 (N_3724,N_3569,N_3488);
or U3725 (N_3725,N_3587,N_3516);
nand U3726 (N_3726,N_3519,N_3485);
or U3727 (N_3727,N_3409,N_3422);
nor U3728 (N_3728,N_3512,N_3403);
and U3729 (N_3729,N_3558,N_3593);
or U3730 (N_3730,N_3555,N_3404);
and U3731 (N_3731,N_3476,N_3532);
xnor U3732 (N_3732,N_3461,N_3432);
nor U3733 (N_3733,N_3450,N_3465);
nor U3734 (N_3734,N_3503,N_3488);
and U3735 (N_3735,N_3530,N_3566);
nand U3736 (N_3736,N_3584,N_3404);
nor U3737 (N_3737,N_3426,N_3570);
nand U3738 (N_3738,N_3438,N_3451);
nor U3739 (N_3739,N_3449,N_3487);
nand U3740 (N_3740,N_3425,N_3482);
or U3741 (N_3741,N_3466,N_3556);
or U3742 (N_3742,N_3547,N_3534);
nor U3743 (N_3743,N_3473,N_3565);
or U3744 (N_3744,N_3517,N_3577);
nor U3745 (N_3745,N_3443,N_3547);
nor U3746 (N_3746,N_3491,N_3506);
nor U3747 (N_3747,N_3545,N_3508);
and U3748 (N_3748,N_3474,N_3559);
and U3749 (N_3749,N_3555,N_3417);
nor U3750 (N_3750,N_3402,N_3419);
nor U3751 (N_3751,N_3560,N_3470);
or U3752 (N_3752,N_3429,N_3538);
nor U3753 (N_3753,N_3592,N_3572);
nor U3754 (N_3754,N_3582,N_3572);
or U3755 (N_3755,N_3443,N_3586);
nor U3756 (N_3756,N_3457,N_3504);
nor U3757 (N_3757,N_3577,N_3490);
and U3758 (N_3758,N_3560,N_3515);
and U3759 (N_3759,N_3547,N_3452);
or U3760 (N_3760,N_3567,N_3484);
and U3761 (N_3761,N_3512,N_3518);
or U3762 (N_3762,N_3430,N_3485);
nor U3763 (N_3763,N_3577,N_3524);
and U3764 (N_3764,N_3428,N_3534);
and U3765 (N_3765,N_3590,N_3431);
or U3766 (N_3766,N_3567,N_3433);
or U3767 (N_3767,N_3548,N_3456);
nand U3768 (N_3768,N_3476,N_3418);
nand U3769 (N_3769,N_3576,N_3473);
and U3770 (N_3770,N_3505,N_3410);
and U3771 (N_3771,N_3510,N_3502);
and U3772 (N_3772,N_3437,N_3451);
nor U3773 (N_3773,N_3515,N_3522);
nand U3774 (N_3774,N_3588,N_3432);
and U3775 (N_3775,N_3466,N_3521);
nand U3776 (N_3776,N_3579,N_3474);
nand U3777 (N_3777,N_3431,N_3555);
nand U3778 (N_3778,N_3586,N_3596);
or U3779 (N_3779,N_3481,N_3535);
nor U3780 (N_3780,N_3449,N_3411);
xnor U3781 (N_3781,N_3501,N_3435);
or U3782 (N_3782,N_3404,N_3483);
and U3783 (N_3783,N_3404,N_3537);
or U3784 (N_3784,N_3501,N_3477);
nor U3785 (N_3785,N_3506,N_3452);
and U3786 (N_3786,N_3520,N_3458);
nor U3787 (N_3787,N_3454,N_3506);
nor U3788 (N_3788,N_3479,N_3409);
or U3789 (N_3789,N_3522,N_3469);
and U3790 (N_3790,N_3403,N_3588);
and U3791 (N_3791,N_3534,N_3519);
nand U3792 (N_3792,N_3475,N_3593);
or U3793 (N_3793,N_3450,N_3551);
nor U3794 (N_3794,N_3461,N_3565);
nor U3795 (N_3795,N_3533,N_3552);
nor U3796 (N_3796,N_3409,N_3567);
or U3797 (N_3797,N_3487,N_3446);
nand U3798 (N_3798,N_3555,N_3457);
nand U3799 (N_3799,N_3525,N_3449);
or U3800 (N_3800,N_3742,N_3740);
nand U3801 (N_3801,N_3769,N_3646);
nand U3802 (N_3802,N_3739,N_3621);
nor U3803 (N_3803,N_3689,N_3765);
and U3804 (N_3804,N_3793,N_3788);
nor U3805 (N_3805,N_3760,N_3732);
or U3806 (N_3806,N_3761,N_3659);
and U3807 (N_3807,N_3703,N_3613);
or U3808 (N_3808,N_3705,N_3609);
or U3809 (N_3809,N_3662,N_3757);
nand U3810 (N_3810,N_3784,N_3714);
nand U3811 (N_3811,N_3605,N_3617);
and U3812 (N_3812,N_3794,N_3730);
and U3813 (N_3813,N_3622,N_3669);
nand U3814 (N_3814,N_3683,N_3666);
nand U3815 (N_3815,N_3670,N_3686);
nor U3816 (N_3816,N_3789,N_3672);
nor U3817 (N_3817,N_3638,N_3653);
nor U3818 (N_3818,N_3762,N_3658);
and U3819 (N_3819,N_3787,N_3717);
or U3820 (N_3820,N_3756,N_3770);
nor U3821 (N_3821,N_3719,N_3636);
nor U3822 (N_3822,N_3779,N_3624);
or U3823 (N_3823,N_3615,N_3734);
or U3824 (N_3824,N_3688,N_3652);
and U3825 (N_3825,N_3750,N_3764);
or U3826 (N_3826,N_3713,N_3712);
nor U3827 (N_3827,N_3641,N_3720);
and U3828 (N_3828,N_3664,N_3618);
or U3829 (N_3829,N_3637,N_3663);
nor U3830 (N_3830,N_3655,N_3731);
and U3831 (N_3831,N_3639,N_3702);
and U3832 (N_3832,N_3772,N_3709);
and U3833 (N_3833,N_3644,N_3774);
nand U3834 (N_3834,N_3735,N_3758);
nand U3835 (N_3835,N_3642,N_3674);
or U3836 (N_3836,N_3629,N_3648);
nor U3837 (N_3837,N_3773,N_3699);
nand U3838 (N_3838,N_3775,N_3738);
or U3839 (N_3839,N_3797,N_3700);
nor U3840 (N_3840,N_3679,N_3616);
or U3841 (N_3841,N_3791,N_3799);
nor U3842 (N_3842,N_3675,N_3634);
or U3843 (N_3843,N_3657,N_3623);
or U3844 (N_3844,N_3747,N_3630);
or U3845 (N_3845,N_3710,N_3614);
nor U3846 (N_3846,N_3628,N_3635);
nor U3847 (N_3847,N_3681,N_3723);
nand U3848 (N_3848,N_3647,N_3729);
or U3849 (N_3849,N_3656,N_3610);
nor U3850 (N_3850,N_3776,N_3667);
or U3851 (N_3851,N_3744,N_3694);
and U3852 (N_3852,N_3786,N_3736);
nand U3853 (N_3853,N_3654,N_3781);
nand U3854 (N_3854,N_3661,N_3725);
nor U3855 (N_3855,N_3745,N_3727);
nand U3856 (N_3856,N_3753,N_3754);
nor U3857 (N_3857,N_3778,N_3695);
nor U3858 (N_3858,N_3706,N_3696);
or U3859 (N_3859,N_3708,N_3766);
nand U3860 (N_3860,N_3677,N_3668);
and U3861 (N_3861,N_3768,N_3697);
xor U3862 (N_3862,N_3606,N_3660);
nand U3863 (N_3863,N_3746,N_3604);
or U3864 (N_3864,N_3627,N_3782);
nand U3865 (N_3865,N_3741,N_3625);
nand U3866 (N_3866,N_3722,N_3608);
or U3867 (N_3867,N_3690,N_3759);
nand U3868 (N_3868,N_3733,N_3743);
and U3869 (N_3869,N_3633,N_3798);
or U3870 (N_3870,N_3611,N_3749);
nand U3871 (N_3871,N_3698,N_3620);
nand U3872 (N_3872,N_3691,N_3716);
or U3873 (N_3873,N_3796,N_3651);
nor U3874 (N_3874,N_3626,N_3783);
or U3875 (N_3875,N_3721,N_3685);
nor U3876 (N_3876,N_3780,N_3715);
nand U3877 (N_3877,N_3678,N_3792);
nor U3878 (N_3878,N_3619,N_3649);
nand U3879 (N_3879,N_3640,N_3600);
nand U3880 (N_3880,N_3601,N_3671);
or U3881 (N_3881,N_3701,N_3777);
nor U3882 (N_3882,N_3763,N_3643);
nand U3883 (N_3883,N_3650,N_3707);
or U3884 (N_3884,N_3632,N_3751);
nand U3885 (N_3885,N_3676,N_3704);
nor U3886 (N_3886,N_3752,N_3767);
or U3887 (N_3887,N_3755,N_3790);
or U3888 (N_3888,N_3687,N_3726);
nor U3889 (N_3889,N_3631,N_3673);
or U3890 (N_3890,N_3684,N_3682);
or U3891 (N_3891,N_3771,N_3602);
or U3892 (N_3892,N_3785,N_3603);
nand U3893 (N_3893,N_3665,N_3728);
nand U3894 (N_3894,N_3718,N_3737);
nand U3895 (N_3895,N_3795,N_3693);
nor U3896 (N_3896,N_3692,N_3711);
nand U3897 (N_3897,N_3607,N_3724);
nand U3898 (N_3898,N_3748,N_3612);
nor U3899 (N_3899,N_3680,N_3645);
and U3900 (N_3900,N_3693,N_3611);
nor U3901 (N_3901,N_3764,N_3641);
and U3902 (N_3902,N_3764,N_3667);
nand U3903 (N_3903,N_3756,N_3741);
or U3904 (N_3904,N_3734,N_3664);
nand U3905 (N_3905,N_3700,N_3768);
nand U3906 (N_3906,N_3731,N_3609);
nor U3907 (N_3907,N_3680,N_3737);
nand U3908 (N_3908,N_3707,N_3796);
or U3909 (N_3909,N_3719,N_3704);
and U3910 (N_3910,N_3687,N_3783);
or U3911 (N_3911,N_3663,N_3602);
nand U3912 (N_3912,N_3747,N_3709);
or U3913 (N_3913,N_3765,N_3750);
xor U3914 (N_3914,N_3647,N_3735);
or U3915 (N_3915,N_3690,N_3791);
and U3916 (N_3916,N_3723,N_3695);
nor U3917 (N_3917,N_3736,N_3777);
nor U3918 (N_3918,N_3727,N_3668);
and U3919 (N_3919,N_3633,N_3750);
or U3920 (N_3920,N_3685,N_3652);
or U3921 (N_3921,N_3707,N_3613);
or U3922 (N_3922,N_3695,N_3600);
nor U3923 (N_3923,N_3629,N_3680);
nor U3924 (N_3924,N_3738,N_3608);
nand U3925 (N_3925,N_3703,N_3640);
nand U3926 (N_3926,N_3642,N_3776);
xnor U3927 (N_3927,N_3629,N_3604);
or U3928 (N_3928,N_3794,N_3796);
or U3929 (N_3929,N_3721,N_3620);
and U3930 (N_3930,N_3782,N_3686);
and U3931 (N_3931,N_3730,N_3623);
and U3932 (N_3932,N_3620,N_3653);
nor U3933 (N_3933,N_3702,N_3790);
nor U3934 (N_3934,N_3702,N_3651);
or U3935 (N_3935,N_3645,N_3623);
and U3936 (N_3936,N_3794,N_3707);
or U3937 (N_3937,N_3775,N_3751);
nor U3938 (N_3938,N_3617,N_3743);
or U3939 (N_3939,N_3617,N_3635);
and U3940 (N_3940,N_3684,N_3701);
and U3941 (N_3941,N_3722,N_3783);
or U3942 (N_3942,N_3603,N_3697);
or U3943 (N_3943,N_3793,N_3645);
or U3944 (N_3944,N_3746,N_3744);
or U3945 (N_3945,N_3752,N_3747);
or U3946 (N_3946,N_3737,N_3751);
nor U3947 (N_3947,N_3607,N_3733);
nand U3948 (N_3948,N_3724,N_3649);
xnor U3949 (N_3949,N_3632,N_3695);
and U3950 (N_3950,N_3650,N_3701);
and U3951 (N_3951,N_3607,N_3663);
and U3952 (N_3952,N_3626,N_3645);
and U3953 (N_3953,N_3667,N_3737);
nor U3954 (N_3954,N_3615,N_3682);
nor U3955 (N_3955,N_3706,N_3665);
nand U3956 (N_3956,N_3751,N_3690);
and U3957 (N_3957,N_3690,N_3634);
and U3958 (N_3958,N_3693,N_3745);
nor U3959 (N_3959,N_3670,N_3614);
and U3960 (N_3960,N_3757,N_3673);
or U3961 (N_3961,N_3694,N_3779);
or U3962 (N_3962,N_3677,N_3755);
nor U3963 (N_3963,N_3612,N_3736);
and U3964 (N_3964,N_3622,N_3647);
and U3965 (N_3965,N_3758,N_3721);
nand U3966 (N_3966,N_3616,N_3647);
and U3967 (N_3967,N_3742,N_3791);
nor U3968 (N_3968,N_3789,N_3703);
nor U3969 (N_3969,N_3763,N_3681);
or U3970 (N_3970,N_3669,N_3601);
or U3971 (N_3971,N_3745,N_3651);
nor U3972 (N_3972,N_3725,N_3775);
nor U3973 (N_3973,N_3738,N_3659);
or U3974 (N_3974,N_3770,N_3713);
or U3975 (N_3975,N_3708,N_3655);
and U3976 (N_3976,N_3789,N_3613);
nor U3977 (N_3977,N_3736,N_3785);
or U3978 (N_3978,N_3603,N_3676);
nand U3979 (N_3979,N_3613,N_3604);
nand U3980 (N_3980,N_3611,N_3797);
and U3981 (N_3981,N_3607,N_3687);
and U3982 (N_3982,N_3768,N_3776);
nand U3983 (N_3983,N_3696,N_3639);
nand U3984 (N_3984,N_3672,N_3776);
nor U3985 (N_3985,N_3689,N_3611);
and U3986 (N_3986,N_3696,N_3750);
or U3987 (N_3987,N_3639,N_3667);
or U3988 (N_3988,N_3717,N_3606);
nand U3989 (N_3989,N_3627,N_3636);
nor U3990 (N_3990,N_3614,N_3798);
and U3991 (N_3991,N_3695,N_3698);
nor U3992 (N_3992,N_3623,N_3610);
and U3993 (N_3993,N_3708,N_3745);
or U3994 (N_3994,N_3755,N_3628);
nand U3995 (N_3995,N_3736,N_3763);
or U3996 (N_3996,N_3779,N_3603);
and U3997 (N_3997,N_3744,N_3785);
nand U3998 (N_3998,N_3718,N_3637);
nor U3999 (N_3999,N_3604,N_3761);
nand U4000 (N_4000,N_3948,N_3937);
nand U4001 (N_4001,N_3836,N_3926);
nor U4002 (N_4002,N_3882,N_3806);
and U4003 (N_4003,N_3914,N_3827);
and U4004 (N_4004,N_3972,N_3936);
nor U4005 (N_4005,N_3977,N_3952);
or U4006 (N_4006,N_3903,N_3930);
and U4007 (N_4007,N_3838,N_3970);
nand U4008 (N_4008,N_3818,N_3996);
and U4009 (N_4009,N_3848,N_3857);
nand U4010 (N_4010,N_3992,N_3958);
or U4011 (N_4011,N_3912,N_3802);
or U4012 (N_4012,N_3891,N_3847);
and U4013 (N_4013,N_3815,N_3889);
or U4014 (N_4014,N_3879,N_3834);
or U4015 (N_4015,N_3976,N_3951);
nand U4016 (N_4016,N_3820,N_3925);
nor U4017 (N_4017,N_3991,N_3869);
nor U4018 (N_4018,N_3899,N_3931);
xnor U4019 (N_4019,N_3949,N_3844);
and U4020 (N_4020,N_3947,N_3933);
and U4021 (N_4021,N_3942,N_3893);
nor U4022 (N_4022,N_3957,N_3805);
nand U4023 (N_4023,N_3884,N_3814);
nor U4024 (N_4024,N_3812,N_3974);
or U4025 (N_4025,N_3966,N_3975);
nand U4026 (N_4026,N_3953,N_3856);
nand U4027 (N_4027,N_3923,N_3973);
or U4028 (N_4028,N_3829,N_3868);
nand U4029 (N_4029,N_3900,N_3995);
and U4030 (N_4030,N_3855,N_3983);
and U4031 (N_4031,N_3984,N_3934);
nor U4032 (N_4032,N_3885,N_3831);
nor U4033 (N_4033,N_3928,N_3842);
nand U4034 (N_4034,N_3998,N_3927);
nor U4035 (N_4035,N_3908,N_3811);
and U4036 (N_4036,N_3898,N_3870);
and U4037 (N_4037,N_3804,N_3968);
xnor U4038 (N_4038,N_3994,N_3935);
nor U4039 (N_4039,N_3852,N_3999);
nor U4040 (N_4040,N_3807,N_3924);
nand U4041 (N_4041,N_3997,N_3978);
and U4042 (N_4042,N_3967,N_3918);
and U4043 (N_4043,N_3840,N_3828);
nand U4044 (N_4044,N_3866,N_3982);
nand U4045 (N_4045,N_3830,N_3904);
nand U4046 (N_4046,N_3886,N_3905);
or U4047 (N_4047,N_3919,N_3946);
or U4048 (N_4048,N_3878,N_3888);
or U4049 (N_4049,N_3841,N_3892);
nor U4050 (N_4050,N_3846,N_3960);
nand U4051 (N_4051,N_3965,N_3833);
and U4052 (N_4052,N_3859,N_3932);
and U4053 (N_4053,N_3961,N_3962);
nor U4054 (N_4054,N_3909,N_3823);
or U4055 (N_4055,N_3938,N_3963);
and U4056 (N_4056,N_3813,N_3971);
and U4057 (N_4057,N_3808,N_3993);
nor U4058 (N_4058,N_3837,N_3944);
nand U4059 (N_4059,N_3987,N_3801);
nor U4060 (N_4060,N_3862,N_3890);
or U4061 (N_4061,N_3921,N_3881);
or U4062 (N_4062,N_3876,N_3985);
and U4063 (N_4063,N_3810,N_3850);
or U4064 (N_4064,N_3959,N_3920);
and U4065 (N_4065,N_3988,N_3849);
or U4066 (N_4066,N_3824,N_3956);
nand U4067 (N_4067,N_3863,N_3939);
nor U4068 (N_4068,N_3954,N_3981);
nand U4069 (N_4069,N_3800,N_3887);
nor U4070 (N_4070,N_3864,N_3803);
and U4071 (N_4071,N_3832,N_3872);
nor U4072 (N_4072,N_3941,N_3874);
and U4073 (N_4073,N_3894,N_3858);
or U4074 (N_4074,N_3986,N_3943);
or U4075 (N_4075,N_3860,N_3969);
nor U4076 (N_4076,N_3826,N_3913);
or U4077 (N_4077,N_3851,N_3945);
or U4078 (N_4078,N_3854,N_3809);
nor U4079 (N_4079,N_3839,N_3867);
or U4080 (N_4080,N_3990,N_3955);
nand U4081 (N_4081,N_3817,N_3922);
nand U4082 (N_4082,N_3915,N_3911);
nand U4083 (N_4083,N_3822,N_3875);
and U4084 (N_4084,N_3835,N_3979);
nor U4085 (N_4085,N_3843,N_3895);
nor U4086 (N_4086,N_3902,N_3916);
and U4087 (N_4087,N_3816,N_3873);
or U4088 (N_4088,N_3825,N_3910);
nand U4089 (N_4089,N_3865,N_3877);
nand U4090 (N_4090,N_3883,N_3845);
and U4091 (N_4091,N_3871,N_3980);
nand U4092 (N_4092,N_3964,N_3907);
nor U4093 (N_4093,N_3989,N_3861);
or U4094 (N_4094,N_3929,N_3950);
and U4095 (N_4095,N_3901,N_3940);
xor U4096 (N_4096,N_3821,N_3880);
nor U4097 (N_4097,N_3906,N_3853);
or U4098 (N_4098,N_3896,N_3917);
nand U4099 (N_4099,N_3819,N_3897);
nand U4100 (N_4100,N_3863,N_3862);
nor U4101 (N_4101,N_3916,N_3804);
nor U4102 (N_4102,N_3873,N_3982);
nand U4103 (N_4103,N_3981,N_3859);
and U4104 (N_4104,N_3871,N_3947);
nor U4105 (N_4105,N_3843,N_3862);
or U4106 (N_4106,N_3847,N_3851);
nand U4107 (N_4107,N_3801,N_3803);
nor U4108 (N_4108,N_3850,N_3833);
and U4109 (N_4109,N_3871,N_3887);
nor U4110 (N_4110,N_3886,N_3865);
or U4111 (N_4111,N_3813,N_3948);
nand U4112 (N_4112,N_3832,N_3969);
nand U4113 (N_4113,N_3976,N_3897);
or U4114 (N_4114,N_3813,N_3832);
nand U4115 (N_4115,N_3890,N_3879);
nor U4116 (N_4116,N_3909,N_3963);
nor U4117 (N_4117,N_3935,N_3907);
nor U4118 (N_4118,N_3970,N_3877);
and U4119 (N_4119,N_3962,N_3949);
nor U4120 (N_4120,N_3920,N_3999);
nand U4121 (N_4121,N_3965,N_3983);
or U4122 (N_4122,N_3864,N_3969);
nor U4123 (N_4123,N_3996,N_3943);
and U4124 (N_4124,N_3859,N_3940);
nand U4125 (N_4125,N_3808,N_3826);
nor U4126 (N_4126,N_3967,N_3962);
or U4127 (N_4127,N_3963,N_3890);
nor U4128 (N_4128,N_3988,N_3853);
or U4129 (N_4129,N_3957,N_3920);
or U4130 (N_4130,N_3942,N_3904);
or U4131 (N_4131,N_3921,N_3876);
or U4132 (N_4132,N_3879,N_3831);
nor U4133 (N_4133,N_3940,N_3887);
nand U4134 (N_4134,N_3912,N_3920);
or U4135 (N_4135,N_3825,N_3981);
and U4136 (N_4136,N_3840,N_3920);
and U4137 (N_4137,N_3914,N_3905);
or U4138 (N_4138,N_3983,N_3917);
and U4139 (N_4139,N_3851,N_3969);
or U4140 (N_4140,N_3954,N_3805);
nand U4141 (N_4141,N_3996,N_3966);
and U4142 (N_4142,N_3891,N_3819);
xnor U4143 (N_4143,N_3857,N_3927);
or U4144 (N_4144,N_3992,N_3932);
nor U4145 (N_4145,N_3900,N_3827);
or U4146 (N_4146,N_3975,N_3999);
xnor U4147 (N_4147,N_3834,N_3877);
nor U4148 (N_4148,N_3999,N_3972);
or U4149 (N_4149,N_3930,N_3851);
nand U4150 (N_4150,N_3868,N_3927);
nand U4151 (N_4151,N_3905,N_3997);
nand U4152 (N_4152,N_3914,N_3986);
and U4153 (N_4153,N_3983,N_3884);
or U4154 (N_4154,N_3839,N_3963);
nand U4155 (N_4155,N_3978,N_3867);
nand U4156 (N_4156,N_3865,N_3891);
and U4157 (N_4157,N_3918,N_3965);
and U4158 (N_4158,N_3827,N_3958);
nand U4159 (N_4159,N_3892,N_3830);
or U4160 (N_4160,N_3885,N_3988);
nand U4161 (N_4161,N_3913,N_3841);
nor U4162 (N_4162,N_3970,N_3848);
or U4163 (N_4163,N_3964,N_3854);
nor U4164 (N_4164,N_3926,N_3891);
and U4165 (N_4165,N_3992,N_3994);
xor U4166 (N_4166,N_3984,N_3876);
and U4167 (N_4167,N_3912,N_3926);
and U4168 (N_4168,N_3804,N_3887);
or U4169 (N_4169,N_3994,N_3955);
nand U4170 (N_4170,N_3907,N_3980);
and U4171 (N_4171,N_3816,N_3832);
or U4172 (N_4172,N_3947,N_3968);
and U4173 (N_4173,N_3966,N_3988);
nor U4174 (N_4174,N_3867,N_3855);
and U4175 (N_4175,N_3981,N_3839);
nand U4176 (N_4176,N_3837,N_3809);
nor U4177 (N_4177,N_3813,N_3872);
or U4178 (N_4178,N_3814,N_3867);
and U4179 (N_4179,N_3929,N_3803);
or U4180 (N_4180,N_3810,N_3911);
nor U4181 (N_4181,N_3827,N_3975);
and U4182 (N_4182,N_3898,N_3981);
nand U4183 (N_4183,N_3979,N_3987);
nor U4184 (N_4184,N_3954,N_3986);
nor U4185 (N_4185,N_3886,N_3825);
nor U4186 (N_4186,N_3965,N_3886);
nor U4187 (N_4187,N_3998,N_3847);
nor U4188 (N_4188,N_3877,N_3955);
or U4189 (N_4189,N_3820,N_3804);
or U4190 (N_4190,N_3914,N_3982);
and U4191 (N_4191,N_3939,N_3897);
xnor U4192 (N_4192,N_3933,N_3823);
nand U4193 (N_4193,N_3835,N_3963);
nand U4194 (N_4194,N_3872,N_3919);
nor U4195 (N_4195,N_3879,N_3923);
and U4196 (N_4196,N_3884,N_3826);
or U4197 (N_4197,N_3965,N_3843);
nand U4198 (N_4198,N_3870,N_3857);
nand U4199 (N_4199,N_3822,N_3883);
and U4200 (N_4200,N_4151,N_4167);
nand U4201 (N_4201,N_4129,N_4139);
or U4202 (N_4202,N_4075,N_4035);
and U4203 (N_4203,N_4156,N_4168);
xor U4204 (N_4204,N_4196,N_4111);
nor U4205 (N_4205,N_4098,N_4056);
and U4206 (N_4206,N_4149,N_4161);
nand U4207 (N_4207,N_4188,N_4070);
nor U4208 (N_4208,N_4079,N_4185);
nand U4209 (N_4209,N_4158,N_4050);
xor U4210 (N_4210,N_4010,N_4174);
nand U4211 (N_4211,N_4060,N_4181);
nand U4212 (N_4212,N_4143,N_4085);
nand U4213 (N_4213,N_4072,N_4178);
nand U4214 (N_4214,N_4117,N_4131);
or U4215 (N_4215,N_4091,N_4033);
nand U4216 (N_4216,N_4121,N_4045);
or U4217 (N_4217,N_4047,N_4146);
nand U4218 (N_4218,N_4113,N_4136);
or U4219 (N_4219,N_4027,N_4066);
nor U4220 (N_4220,N_4059,N_4042);
and U4221 (N_4221,N_4133,N_4134);
nand U4222 (N_4222,N_4030,N_4002);
and U4223 (N_4223,N_4171,N_4165);
nand U4224 (N_4224,N_4062,N_4106);
nor U4225 (N_4225,N_4065,N_4150);
or U4226 (N_4226,N_4198,N_4071);
or U4227 (N_4227,N_4140,N_4166);
nand U4228 (N_4228,N_4063,N_4018);
nor U4229 (N_4229,N_4105,N_4123);
and U4230 (N_4230,N_4017,N_4159);
or U4231 (N_4231,N_4080,N_4088);
and U4232 (N_4232,N_4046,N_4005);
nand U4233 (N_4233,N_4144,N_4154);
or U4234 (N_4234,N_4054,N_4038);
and U4235 (N_4235,N_4122,N_4162);
or U4236 (N_4236,N_4084,N_4192);
or U4237 (N_4237,N_4053,N_4128);
or U4238 (N_4238,N_4015,N_4100);
nand U4239 (N_4239,N_4004,N_4182);
and U4240 (N_4240,N_4157,N_4126);
nand U4241 (N_4241,N_4094,N_4041);
nor U4242 (N_4242,N_4049,N_4120);
nand U4243 (N_4243,N_4077,N_4110);
nor U4244 (N_4244,N_4081,N_4177);
nand U4245 (N_4245,N_4189,N_4170);
xor U4246 (N_4246,N_4073,N_4012);
and U4247 (N_4247,N_4020,N_4114);
nor U4248 (N_4248,N_4039,N_4090);
or U4249 (N_4249,N_4104,N_4031);
and U4250 (N_4250,N_4026,N_4093);
and U4251 (N_4251,N_4097,N_4029);
and U4252 (N_4252,N_4019,N_4006);
nor U4253 (N_4253,N_4199,N_4078);
and U4254 (N_4254,N_4180,N_4191);
nand U4255 (N_4255,N_4096,N_4024);
and U4256 (N_4256,N_4124,N_4175);
nor U4257 (N_4257,N_4083,N_4130);
and U4258 (N_4258,N_4099,N_4116);
or U4259 (N_4259,N_4197,N_4001);
nor U4260 (N_4260,N_4135,N_4118);
and U4261 (N_4261,N_4064,N_4068);
nor U4262 (N_4262,N_4142,N_4176);
or U4263 (N_4263,N_4016,N_4119);
nor U4264 (N_4264,N_4011,N_4164);
or U4265 (N_4265,N_4132,N_4115);
nand U4266 (N_4266,N_4037,N_4013);
nor U4267 (N_4267,N_4007,N_4160);
and U4268 (N_4268,N_4187,N_4112);
or U4269 (N_4269,N_4108,N_4125);
and U4270 (N_4270,N_4152,N_4101);
and U4271 (N_4271,N_4194,N_4055);
nand U4272 (N_4272,N_4032,N_4076);
nand U4273 (N_4273,N_4000,N_4195);
and U4274 (N_4274,N_4008,N_4009);
and U4275 (N_4275,N_4023,N_4040);
or U4276 (N_4276,N_4014,N_4043);
and U4277 (N_4277,N_4082,N_4057);
or U4278 (N_4278,N_4193,N_4021);
nor U4279 (N_4279,N_4022,N_4061);
or U4280 (N_4280,N_4169,N_4069);
or U4281 (N_4281,N_4052,N_4051);
nand U4282 (N_4282,N_4138,N_4058);
nor U4283 (N_4283,N_4127,N_4089);
nor U4284 (N_4284,N_4028,N_4103);
and U4285 (N_4285,N_4147,N_4036);
nand U4286 (N_4286,N_4092,N_4086);
and U4287 (N_4287,N_4155,N_4025);
nor U4288 (N_4288,N_4107,N_4163);
nor U4289 (N_4289,N_4034,N_4044);
nand U4290 (N_4290,N_4067,N_4183);
and U4291 (N_4291,N_4074,N_4003);
or U4292 (N_4292,N_4141,N_4190);
or U4293 (N_4293,N_4186,N_4179);
or U4294 (N_4294,N_4137,N_4148);
and U4295 (N_4295,N_4153,N_4145);
and U4296 (N_4296,N_4109,N_4173);
nand U4297 (N_4297,N_4087,N_4102);
or U4298 (N_4298,N_4095,N_4048);
nor U4299 (N_4299,N_4184,N_4172);
or U4300 (N_4300,N_4164,N_4121);
and U4301 (N_4301,N_4154,N_4153);
nor U4302 (N_4302,N_4046,N_4145);
or U4303 (N_4303,N_4081,N_4128);
nor U4304 (N_4304,N_4079,N_4085);
or U4305 (N_4305,N_4054,N_4089);
nor U4306 (N_4306,N_4079,N_4161);
nor U4307 (N_4307,N_4009,N_4001);
or U4308 (N_4308,N_4137,N_4183);
and U4309 (N_4309,N_4154,N_4131);
nor U4310 (N_4310,N_4028,N_4066);
nand U4311 (N_4311,N_4132,N_4009);
nand U4312 (N_4312,N_4056,N_4091);
or U4313 (N_4313,N_4149,N_4106);
or U4314 (N_4314,N_4079,N_4107);
and U4315 (N_4315,N_4111,N_4190);
or U4316 (N_4316,N_4003,N_4028);
nor U4317 (N_4317,N_4088,N_4160);
nand U4318 (N_4318,N_4042,N_4031);
nor U4319 (N_4319,N_4026,N_4010);
nor U4320 (N_4320,N_4129,N_4025);
or U4321 (N_4321,N_4009,N_4119);
nand U4322 (N_4322,N_4085,N_4033);
nand U4323 (N_4323,N_4157,N_4079);
xor U4324 (N_4324,N_4186,N_4106);
or U4325 (N_4325,N_4173,N_4137);
and U4326 (N_4326,N_4077,N_4045);
or U4327 (N_4327,N_4141,N_4089);
or U4328 (N_4328,N_4054,N_4035);
and U4329 (N_4329,N_4168,N_4123);
nor U4330 (N_4330,N_4170,N_4068);
or U4331 (N_4331,N_4152,N_4035);
nor U4332 (N_4332,N_4062,N_4065);
or U4333 (N_4333,N_4144,N_4173);
nand U4334 (N_4334,N_4168,N_4089);
and U4335 (N_4335,N_4045,N_4159);
nand U4336 (N_4336,N_4177,N_4142);
or U4337 (N_4337,N_4073,N_4151);
or U4338 (N_4338,N_4101,N_4073);
nand U4339 (N_4339,N_4178,N_4081);
nor U4340 (N_4340,N_4066,N_4055);
nand U4341 (N_4341,N_4108,N_4008);
or U4342 (N_4342,N_4055,N_4082);
or U4343 (N_4343,N_4142,N_4188);
nand U4344 (N_4344,N_4167,N_4196);
or U4345 (N_4345,N_4189,N_4076);
nor U4346 (N_4346,N_4159,N_4062);
nand U4347 (N_4347,N_4168,N_4125);
and U4348 (N_4348,N_4128,N_4162);
or U4349 (N_4349,N_4019,N_4037);
nand U4350 (N_4350,N_4193,N_4159);
nor U4351 (N_4351,N_4003,N_4186);
and U4352 (N_4352,N_4194,N_4012);
xor U4353 (N_4353,N_4181,N_4109);
and U4354 (N_4354,N_4135,N_4033);
and U4355 (N_4355,N_4186,N_4084);
and U4356 (N_4356,N_4117,N_4076);
and U4357 (N_4357,N_4003,N_4173);
nand U4358 (N_4358,N_4101,N_4193);
or U4359 (N_4359,N_4164,N_4088);
or U4360 (N_4360,N_4087,N_4099);
nand U4361 (N_4361,N_4104,N_4147);
nand U4362 (N_4362,N_4020,N_4069);
nor U4363 (N_4363,N_4112,N_4096);
nand U4364 (N_4364,N_4135,N_4038);
nand U4365 (N_4365,N_4068,N_4057);
or U4366 (N_4366,N_4011,N_4079);
or U4367 (N_4367,N_4191,N_4159);
nand U4368 (N_4368,N_4018,N_4009);
and U4369 (N_4369,N_4027,N_4154);
or U4370 (N_4370,N_4121,N_4199);
or U4371 (N_4371,N_4157,N_4192);
or U4372 (N_4372,N_4106,N_4173);
and U4373 (N_4373,N_4171,N_4189);
and U4374 (N_4374,N_4113,N_4005);
and U4375 (N_4375,N_4132,N_4080);
or U4376 (N_4376,N_4138,N_4192);
and U4377 (N_4377,N_4067,N_4070);
or U4378 (N_4378,N_4122,N_4022);
or U4379 (N_4379,N_4029,N_4173);
or U4380 (N_4380,N_4174,N_4061);
or U4381 (N_4381,N_4069,N_4027);
and U4382 (N_4382,N_4031,N_4162);
or U4383 (N_4383,N_4052,N_4018);
and U4384 (N_4384,N_4085,N_4119);
nor U4385 (N_4385,N_4117,N_4192);
or U4386 (N_4386,N_4042,N_4161);
and U4387 (N_4387,N_4056,N_4157);
and U4388 (N_4388,N_4108,N_4172);
or U4389 (N_4389,N_4188,N_4046);
nand U4390 (N_4390,N_4142,N_4152);
or U4391 (N_4391,N_4029,N_4047);
or U4392 (N_4392,N_4165,N_4183);
nor U4393 (N_4393,N_4108,N_4120);
nor U4394 (N_4394,N_4066,N_4098);
nand U4395 (N_4395,N_4031,N_4028);
nor U4396 (N_4396,N_4113,N_4104);
nor U4397 (N_4397,N_4148,N_4114);
and U4398 (N_4398,N_4062,N_4031);
and U4399 (N_4399,N_4104,N_4106);
nor U4400 (N_4400,N_4371,N_4364);
nor U4401 (N_4401,N_4387,N_4217);
and U4402 (N_4402,N_4268,N_4326);
nand U4403 (N_4403,N_4212,N_4298);
and U4404 (N_4404,N_4274,N_4249);
or U4405 (N_4405,N_4359,N_4270);
or U4406 (N_4406,N_4372,N_4292);
nor U4407 (N_4407,N_4368,N_4236);
or U4408 (N_4408,N_4202,N_4308);
nand U4409 (N_4409,N_4351,N_4214);
and U4410 (N_4410,N_4201,N_4231);
or U4411 (N_4411,N_4340,N_4337);
nor U4412 (N_4412,N_4238,N_4376);
nor U4413 (N_4413,N_4240,N_4253);
nor U4414 (N_4414,N_4304,N_4234);
and U4415 (N_4415,N_4206,N_4283);
xor U4416 (N_4416,N_4235,N_4317);
and U4417 (N_4417,N_4209,N_4345);
nand U4418 (N_4418,N_4336,N_4357);
or U4419 (N_4419,N_4284,N_4385);
nor U4420 (N_4420,N_4393,N_4362);
nor U4421 (N_4421,N_4379,N_4369);
nor U4422 (N_4422,N_4287,N_4245);
and U4423 (N_4423,N_4386,N_4289);
nand U4424 (N_4424,N_4338,N_4220);
or U4425 (N_4425,N_4248,N_4224);
nand U4426 (N_4426,N_4313,N_4394);
nand U4427 (N_4427,N_4255,N_4204);
nor U4428 (N_4428,N_4203,N_4205);
xnor U4429 (N_4429,N_4280,N_4318);
nor U4430 (N_4430,N_4276,N_4353);
and U4431 (N_4431,N_4391,N_4327);
or U4432 (N_4432,N_4277,N_4389);
xnor U4433 (N_4433,N_4228,N_4380);
nor U4434 (N_4434,N_4230,N_4264);
or U4435 (N_4435,N_4267,N_4324);
or U4436 (N_4436,N_4250,N_4223);
nor U4437 (N_4437,N_4349,N_4307);
or U4438 (N_4438,N_4365,N_4272);
and U4439 (N_4439,N_4260,N_4208);
nor U4440 (N_4440,N_4328,N_4286);
nand U4441 (N_4441,N_4261,N_4269);
nor U4442 (N_4442,N_4233,N_4388);
nand U4443 (N_4443,N_4232,N_4335);
nor U4444 (N_4444,N_4291,N_4303);
nand U4445 (N_4445,N_4399,N_4305);
nor U4446 (N_4446,N_4299,N_4354);
nor U4447 (N_4447,N_4211,N_4381);
or U4448 (N_4448,N_4251,N_4219);
nor U4449 (N_4449,N_4358,N_4315);
or U4450 (N_4450,N_4221,N_4302);
nor U4451 (N_4451,N_4310,N_4239);
nor U4452 (N_4452,N_4259,N_4363);
or U4453 (N_4453,N_4216,N_4344);
nor U4454 (N_4454,N_4382,N_4256);
and U4455 (N_4455,N_4397,N_4306);
nand U4456 (N_4456,N_4330,N_4398);
and U4457 (N_4457,N_4229,N_4275);
and U4458 (N_4458,N_4300,N_4237);
nor U4459 (N_4459,N_4366,N_4384);
xnor U4460 (N_4460,N_4314,N_4347);
nand U4461 (N_4461,N_4244,N_4271);
nand U4462 (N_4462,N_4341,N_4282);
nor U4463 (N_4463,N_4373,N_4222);
and U4464 (N_4464,N_4301,N_4375);
and U4465 (N_4465,N_4218,N_4348);
nor U4466 (N_4466,N_4213,N_4396);
nand U4467 (N_4467,N_4273,N_4395);
and U4468 (N_4468,N_4254,N_4200);
and U4469 (N_4469,N_4262,N_4295);
xor U4470 (N_4470,N_4339,N_4311);
nor U4471 (N_4471,N_4322,N_4383);
or U4472 (N_4472,N_4266,N_4207);
or U4473 (N_4473,N_4243,N_4390);
nor U4474 (N_4474,N_4252,N_4279);
nor U4475 (N_4475,N_4331,N_4225);
nand U4476 (N_4476,N_4377,N_4293);
nor U4477 (N_4477,N_4352,N_4265);
nand U4478 (N_4478,N_4285,N_4332);
and U4479 (N_4479,N_4333,N_4281);
nand U4480 (N_4480,N_4361,N_4309);
or U4481 (N_4481,N_4246,N_4320);
or U4482 (N_4482,N_4296,N_4258);
nand U4483 (N_4483,N_4257,N_4319);
and U4484 (N_4484,N_4392,N_4343);
or U4485 (N_4485,N_4210,N_4215);
or U4486 (N_4486,N_4355,N_4278);
xor U4487 (N_4487,N_4242,N_4288);
or U4488 (N_4488,N_4329,N_4294);
or U4489 (N_4489,N_4360,N_4312);
and U4490 (N_4490,N_4263,N_4321);
nand U4491 (N_4491,N_4297,N_4325);
and U4492 (N_4492,N_4346,N_4367);
nor U4493 (N_4493,N_4247,N_4378);
and U4494 (N_4494,N_4316,N_4350);
nand U4495 (N_4495,N_4226,N_4342);
nor U4496 (N_4496,N_4334,N_4323);
and U4497 (N_4497,N_4241,N_4374);
nor U4498 (N_4498,N_4356,N_4370);
and U4499 (N_4499,N_4227,N_4290);
nand U4500 (N_4500,N_4318,N_4333);
nor U4501 (N_4501,N_4295,N_4225);
nand U4502 (N_4502,N_4259,N_4361);
nor U4503 (N_4503,N_4358,N_4200);
nand U4504 (N_4504,N_4388,N_4243);
and U4505 (N_4505,N_4371,N_4300);
nand U4506 (N_4506,N_4218,N_4206);
nor U4507 (N_4507,N_4371,N_4275);
nand U4508 (N_4508,N_4356,N_4275);
and U4509 (N_4509,N_4343,N_4326);
xor U4510 (N_4510,N_4216,N_4232);
nand U4511 (N_4511,N_4356,N_4224);
xnor U4512 (N_4512,N_4240,N_4232);
or U4513 (N_4513,N_4311,N_4220);
or U4514 (N_4514,N_4203,N_4289);
nor U4515 (N_4515,N_4396,N_4280);
and U4516 (N_4516,N_4355,N_4328);
xnor U4517 (N_4517,N_4309,N_4380);
or U4518 (N_4518,N_4396,N_4228);
and U4519 (N_4519,N_4392,N_4279);
or U4520 (N_4520,N_4366,N_4263);
nand U4521 (N_4521,N_4256,N_4273);
and U4522 (N_4522,N_4333,N_4370);
and U4523 (N_4523,N_4235,N_4359);
and U4524 (N_4524,N_4375,N_4200);
nor U4525 (N_4525,N_4309,N_4228);
xor U4526 (N_4526,N_4271,N_4305);
nor U4527 (N_4527,N_4328,N_4296);
xor U4528 (N_4528,N_4242,N_4271);
xnor U4529 (N_4529,N_4206,N_4228);
and U4530 (N_4530,N_4339,N_4372);
or U4531 (N_4531,N_4271,N_4211);
or U4532 (N_4532,N_4267,N_4348);
or U4533 (N_4533,N_4261,N_4302);
and U4534 (N_4534,N_4203,N_4396);
or U4535 (N_4535,N_4355,N_4280);
and U4536 (N_4536,N_4380,N_4367);
or U4537 (N_4537,N_4281,N_4371);
nand U4538 (N_4538,N_4309,N_4331);
or U4539 (N_4539,N_4369,N_4377);
or U4540 (N_4540,N_4366,N_4207);
or U4541 (N_4541,N_4206,N_4234);
nand U4542 (N_4542,N_4244,N_4263);
nor U4543 (N_4543,N_4291,N_4289);
nor U4544 (N_4544,N_4263,N_4383);
and U4545 (N_4545,N_4334,N_4277);
nand U4546 (N_4546,N_4269,N_4365);
or U4547 (N_4547,N_4275,N_4242);
and U4548 (N_4548,N_4338,N_4368);
nor U4549 (N_4549,N_4367,N_4394);
and U4550 (N_4550,N_4275,N_4225);
nand U4551 (N_4551,N_4309,N_4327);
nor U4552 (N_4552,N_4353,N_4255);
or U4553 (N_4553,N_4337,N_4327);
nor U4554 (N_4554,N_4380,N_4348);
or U4555 (N_4555,N_4331,N_4339);
or U4556 (N_4556,N_4269,N_4354);
and U4557 (N_4557,N_4292,N_4324);
nand U4558 (N_4558,N_4216,N_4371);
and U4559 (N_4559,N_4254,N_4312);
nor U4560 (N_4560,N_4240,N_4244);
or U4561 (N_4561,N_4293,N_4314);
and U4562 (N_4562,N_4213,N_4303);
nand U4563 (N_4563,N_4268,N_4212);
and U4564 (N_4564,N_4238,N_4311);
nand U4565 (N_4565,N_4374,N_4214);
and U4566 (N_4566,N_4275,N_4274);
or U4567 (N_4567,N_4354,N_4223);
nor U4568 (N_4568,N_4353,N_4278);
nand U4569 (N_4569,N_4395,N_4317);
and U4570 (N_4570,N_4265,N_4377);
or U4571 (N_4571,N_4268,N_4366);
nor U4572 (N_4572,N_4202,N_4365);
or U4573 (N_4573,N_4241,N_4311);
and U4574 (N_4574,N_4209,N_4288);
nand U4575 (N_4575,N_4382,N_4311);
and U4576 (N_4576,N_4203,N_4224);
nand U4577 (N_4577,N_4218,N_4330);
nor U4578 (N_4578,N_4261,N_4210);
and U4579 (N_4579,N_4233,N_4348);
or U4580 (N_4580,N_4344,N_4279);
and U4581 (N_4581,N_4257,N_4276);
nor U4582 (N_4582,N_4204,N_4222);
nor U4583 (N_4583,N_4261,N_4218);
or U4584 (N_4584,N_4389,N_4385);
nor U4585 (N_4585,N_4359,N_4222);
and U4586 (N_4586,N_4389,N_4213);
or U4587 (N_4587,N_4386,N_4393);
nor U4588 (N_4588,N_4208,N_4396);
or U4589 (N_4589,N_4263,N_4331);
nor U4590 (N_4590,N_4386,N_4276);
or U4591 (N_4591,N_4325,N_4333);
or U4592 (N_4592,N_4213,N_4298);
nand U4593 (N_4593,N_4200,N_4261);
nor U4594 (N_4594,N_4338,N_4209);
nand U4595 (N_4595,N_4246,N_4364);
nand U4596 (N_4596,N_4377,N_4264);
and U4597 (N_4597,N_4257,N_4240);
nor U4598 (N_4598,N_4270,N_4372);
and U4599 (N_4599,N_4273,N_4356);
nor U4600 (N_4600,N_4453,N_4579);
nor U4601 (N_4601,N_4533,N_4534);
nor U4602 (N_4602,N_4486,N_4563);
and U4603 (N_4603,N_4530,N_4473);
nand U4604 (N_4604,N_4487,N_4446);
and U4605 (N_4605,N_4516,N_4430);
nand U4606 (N_4606,N_4440,N_4583);
and U4607 (N_4607,N_4434,N_4466);
nand U4608 (N_4608,N_4403,N_4523);
nand U4609 (N_4609,N_4452,N_4432);
or U4610 (N_4610,N_4577,N_4515);
nand U4611 (N_4611,N_4413,N_4506);
nand U4612 (N_4612,N_4475,N_4522);
nor U4613 (N_4613,N_4401,N_4484);
nand U4614 (N_4614,N_4570,N_4468);
and U4615 (N_4615,N_4404,N_4444);
nor U4616 (N_4616,N_4548,N_4589);
or U4617 (N_4617,N_4472,N_4525);
and U4618 (N_4618,N_4580,N_4594);
nor U4619 (N_4619,N_4595,N_4598);
and U4620 (N_4620,N_4471,N_4553);
nor U4621 (N_4621,N_4584,N_4459);
nand U4622 (N_4622,N_4517,N_4443);
nor U4623 (N_4623,N_4496,N_4441);
xor U4624 (N_4624,N_4429,N_4596);
and U4625 (N_4625,N_4442,N_4504);
and U4626 (N_4626,N_4480,N_4560);
and U4627 (N_4627,N_4508,N_4541);
and U4628 (N_4628,N_4435,N_4501);
or U4629 (N_4629,N_4479,N_4426);
and U4630 (N_4630,N_4410,N_4477);
nor U4631 (N_4631,N_4546,N_4561);
nor U4632 (N_4632,N_4428,N_4512);
or U4633 (N_4633,N_4437,N_4542);
or U4634 (N_4634,N_4538,N_4456);
nor U4635 (N_4635,N_4491,N_4599);
nor U4636 (N_4636,N_4463,N_4550);
nand U4637 (N_4637,N_4511,N_4592);
nand U4638 (N_4638,N_4489,N_4564);
nor U4639 (N_4639,N_4558,N_4520);
and U4640 (N_4640,N_4573,N_4519);
or U4641 (N_4641,N_4562,N_4539);
nor U4642 (N_4642,N_4421,N_4445);
or U4643 (N_4643,N_4524,N_4518);
nand U4644 (N_4644,N_4503,N_4510);
and U4645 (N_4645,N_4572,N_4587);
nand U4646 (N_4646,N_4449,N_4494);
or U4647 (N_4647,N_4591,N_4526);
xor U4648 (N_4648,N_4566,N_4425);
nor U4649 (N_4649,N_4551,N_4419);
or U4650 (N_4650,N_4492,N_4549);
or U4651 (N_4651,N_4568,N_4438);
and U4652 (N_4652,N_4439,N_4557);
or U4653 (N_4653,N_4531,N_4588);
nor U4654 (N_4654,N_4405,N_4532);
and U4655 (N_4655,N_4590,N_4482);
or U4656 (N_4656,N_4597,N_4470);
nand U4657 (N_4657,N_4574,N_4460);
nand U4658 (N_4658,N_4567,N_4455);
or U4659 (N_4659,N_4544,N_4556);
nand U4660 (N_4660,N_4528,N_4581);
nor U4661 (N_4661,N_4424,N_4414);
nor U4662 (N_4662,N_4535,N_4474);
nor U4663 (N_4663,N_4409,N_4586);
and U4664 (N_4664,N_4521,N_4420);
or U4665 (N_4665,N_4485,N_4465);
or U4666 (N_4666,N_4529,N_4527);
or U4667 (N_4667,N_4407,N_4476);
nor U4668 (N_4668,N_4411,N_4402);
and U4669 (N_4669,N_4457,N_4450);
nor U4670 (N_4670,N_4447,N_4540);
and U4671 (N_4671,N_4509,N_4507);
nor U4672 (N_4672,N_4493,N_4481);
nor U4673 (N_4673,N_4469,N_4461);
or U4674 (N_4674,N_4433,N_4488);
or U4675 (N_4675,N_4408,N_4406);
or U4676 (N_4676,N_4412,N_4545);
nand U4677 (N_4677,N_4448,N_4547);
or U4678 (N_4678,N_4400,N_4513);
nor U4679 (N_4679,N_4576,N_4483);
or U4680 (N_4680,N_4418,N_4514);
and U4681 (N_4681,N_4415,N_4490);
or U4682 (N_4682,N_4552,N_4575);
or U4683 (N_4683,N_4569,N_4495);
nor U4684 (N_4684,N_4505,N_4582);
and U4685 (N_4685,N_4464,N_4571);
nand U4686 (N_4686,N_4417,N_4431);
nor U4687 (N_4687,N_4537,N_4462);
and U4688 (N_4688,N_4436,N_4543);
or U4689 (N_4689,N_4478,N_4593);
nand U4690 (N_4690,N_4422,N_4498);
and U4691 (N_4691,N_4585,N_4536);
or U4692 (N_4692,N_4578,N_4467);
or U4693 (N_4693,N_4451,N_4454);
and U4694 (N_4694,N_4423,N_4565);
nor U4695 (N_4695,N_4458,N_4502);
nor U4696 (N_4696,N_4416,N_4497);
and U4697 (N_4697,N_4499,N_4555);
and U4698 (N_4698,N_4427,N_4554);
nand U4699 (N_4699,N_4500,N_4559);
and U4700 (N_4700,N_4405,N_4555);
or U4701 (N_4701,N_4439,N_4520);
or U4702 (N_4702,N_4466,N_4520);
nand U4703 (N_4703,N_4475,N_4582);
or U4704 (N_4704,N_4503,N_4509);
and U4705 (N_4705,N_4461,N_4446);
and U4706 (N_4706,N_4532,N_4587);
and U4707 (N_4707,N_4422,N_4476);
nor U4708 (N_4708,N_4598,N_4539);
xor U4709 (N_4709,N_4539,N_4514);
nand U4710 (N_4710,N_4500,N_4413);
nor U4711 (N_4711,N_4554,N_4406);
nor U4712 (N_4712,N_4401,N_4516);
nor U4713 (N_4713,N_4576,N_4451);
nor U4714 (N_4714,N_4480,N_4444);
nor U4715 (N_4715,N_4492,N_4587);
and U4716 (N_4716,N_4554,N_4553);
or U4717 (N_4717,N_4471,N_4522);
or U4718 (N_4718,N_4569,N_4511);
xnor U4719 (N_4719,N_4591,N_4582);
nand U4720 (N_4720,N_4549,N_4506);
nand U4721 (N_4721,N_4417,N_4512);
and U4722 (N_4722,N_4435,N_4541);
nand U4723 (N_4723,N_4482,N_4533);
nor U4724 (N_4724,N_4572,N_4569);
nand U4725 (N_4725,N_4498,N_4540);
and U4726 (N_4726,N_4523,N_4471);
and U4727 (N_4727,N_4577,N_4410);
nor U4728 (N_4728,N_4522,N_4525);
or U4729 (N_4729,N_4587,N_4515);
and U4730 (N_4730,N_4470,N_4515);
nor U4731 (N_4731,N_4405,N_4484);
nand U4732 (N_4732,N_4482,N_4450);
nor U4733 (N_4733,N_4448,N_4437);
nand U4734 (N_4734,N_4517,N_4457);
and U4735 (N_4735,N_4452,N_4436);
nor U4736 (N_4736,N_4539,N_4497);
nand U4737 (N_4737,N_4461,N_4466);
nand U4738 (N_4738,N_4416,N_4586);
nand U4739 (N_4739,N_4588,N_4565);
nor U4740 (N_4740,N_4482,N_4580);
and U4741 (N_4741,N_4502,N_4448);
and U4742 (N_4742,N_4414,N_4453);
nand U4743 (N_4743,N_4406,N_4462);
nor U4744 (N_4744,N_4502,N_4479);
nor U4745 (N_4745,N_4487,N_4517);
or U4746 (N_4746,N_4501,N_4550);
nand U4747 (N_4747,N_4439,N_4410);
nor U4748 (N_4748,N_4590,N_4435);
and U4749 (N_4749,N_4440,N_4420);
nor U4750 (N_4750,N_4556,N_4584);
or U4751 (N_4751,N_4456,N_4415);
or U4752 (N_4752,N_4556,N_4579);
nor U4753 (N_4753,N_4425,N_4564);
and U4754 (N_4754,N_4533,N_4513);
and U4755 (N_4755,N_4442,N_4433);
or U4756 (N_4756,N_4505,N_4423);
and U4757 (N_4757,N_4485,N_4471);
nor U4758 (N_4758,N_4507,N_4587);
and U4759 (N_4759,N_4520,N_4440);
or U4760 (N_4760,N_4421,N_4502);
or U4761 (N_4761,N_4472,N_4432);
or U4762 (N_4762,N_4563,N_4401);
and U4763 (N_4763,N_4443,N_4433);
and U4764 (N_4764,N_4559,N_4583);
nor U4765 (N_4765,N_4547,N_4555);
nand U4766 (N_4766,N_4569,N_4429);
nor U4767 (N_4767,N_4549,N_4575);
and U4768 (N_4768,N_4528,N_4471);
nand U4769 (N_4769,N_4551,N_4426);
or U4770 (N_4770,N_4487,N_4495);
and U4771 (N_4771,N_4537,N_4554);
or U4772 (N_4772,N_4531,N_4545);
nor U4773 (N_4773,N_4467,N_4496);
nor U4774 (N_4774,N_4512,N_4477);
nor U4775 (N_4775,N_4462,N_4440);
nand U4776 (N_4776,N_4598,N_4474);
or U4777 (N_4777,N_4546,N_4445);
or U4778 (N_4778,N_4413,N_4549);
and U4779 (N_4779,N_4482,N_4571);
nand U4780 (N_4780,N_4584,N_4539);
or U4781 (N_4781,N_4455,N_4537);
or U4782 (N_4782,N_4581,N_4477);
and U4783 (N_4783,N_4466,N_4413);
and U4784 (N_4784,N_4503,N_4493);
or U4785 (N_4785,N_4489,N_4459);
nor U4786 (N_4786,N_4464,N_4554);
nor U4787 (N_4787,N_4444,N_4494);
or U4788 (N_4788,N_4596,N_4545);
nor U4789 (N_4789,N_4595,N_4589);
or U4790 (N_4790,N_4524,N_4539);
nor U4791 (N_4791,N_4588,N_4415);
nand U4792 (N_4792,N_4461,N_4511);
and U4793 (N_4793,N_4499,N_4463);
nor U4794 (N_4794,N_4473,N_4490);
nor U4795 (N_4795,N_4555,N_4400);
or U4796 (N_4796,N_4456,N_4483);
or U4797 (N_4797,N_4452,N_4553);
nor U4798 (N_4798,N_4565,N_4494);
and U4799 (N_4799,N_4497,N_4412);
nand U4800 (N_4800,N_4674,N_4611);
or U4801 (N_4801,N_4658,N_4715);
nand U4802 (N_4802,N_4765,N_4751);
and U4803 (N_4803,N_4693,N_4666);
nand U4804 (N_4804,N_4682,N_4767);
or U4805 (N_4805,N_4793,N_4761);
xor U4806 (N_4806,N_4607,N_4694);
xnor U4807 (N_4807,N_4796,N_4713);
or U4808 (N_4808,N_4687,N_4643);
nor U4809 (N_4809,N_4732,N_4706);
xnor U4810 (N_4810,N_4613,N_4781);
and U4811 (N_4811,N_4776,N_4712);
nand U4812 (N_4812,N_4791,N_4616);
or U4813 (N_4813,N_4700,N_4645);
and U4814 (N_4814,N_4782,N_4688);
or U4815 (N_4815,N_4759,N_4755);
nand U4816 (N_4816,N_4698,N_4632);
nand U4817 (N_4817,N_4655,N_4737);
or U4818 (N_4818,N_4663,N_4654);
nor U4819 (N_4819,N_4702,N_4790);
nand U4820 (N_4820,N_4725,N_4748);
nand U4821 (N_4821,N_4710,N_4617);
nand U4822 (N_4822,N_4707,N_4756);
and U4823 (N_4823,N_4699,N_4639);
and U4824 (N_4824,N_4640,N_4681);
or U4825 (N_4825,N_4745,N_4768);
and U4826 (N_4826,N_4680,N_4672);
nand U4827 (N_4827,N_4614,N_4685);
or U4828 (N_4828,N_4665,N_4622);
nand U4829 (N_4829,N_4637,N_4692);
nor U4830 (N_4830,N_4734,N_4775);
nor U4831 (N_4831,N_4600,N_4621);
and U4832 (N_4832,N_4628,N_4608);
and U4833 (N_4833,N_4615,N_4642);
and U4834 (N_4834,N_4619,N_4729);
nand U4835 (N_4835,N_4757,N_4684);
or U4836 (N_4836,N_4605,N_4606);
or U4837 (N_4837,N_4722,N_4749);
nor U4838 (N_4838,N_4669,N_4733);
or U4839 (N_4839,N_4763,N_4742);
nor U4840 (N_4840,N_4668,N_4770);
and U4841 (N_4841,N_4653,N_4670);
nand U4842 (N_4842,N_4696,N_4744);
nand U4843 (N_4843,N_4726,N_4704);
nor U4844 (N_4844,N_4738,N_4774);
and U4845 (N_4845,N_4769,N_4676);
or U4846 (N_4846,N_4758,N_4739);
and U4847 (N_4847,N_4648,N_4603);
or U4848 (N_4848,N_4679,N_4634);
or U4849 (N_4849,N_4691,N_4703);
and U4850 (N_4850,N_4728,N_4612);
nand U4851 (N_4851,N_4683,N_4766);
nand U4852 (N_4852,N_4778,N_4623);
nand U4853 (N_4853,N_4720,N_4656);
and U4854 (N_4854,N_4794,N_4743);
and U4855 (N_4855,N_4650,N_4786);
or U4856 (N_4856,N_4711,N_4741);
nand U4857 (N_4857,N_4626,N_4785);
and U4858 (N_4858,N_4718,N_4671);
nor U4859 (N_4859,N_4708,N_4661);
xnor U4860 (N_4860,N_4610,N_4636);
nand U4861 (N_4861,N_4660,N_4797);
nand U4862 (N_4862,N_4675,N_4752);
nand U4863 (N_4863,N_4602,N_4719);
and U4864 (N_4864,N_4717,N_4764);
nand U4865 (N_4865,N_4601,N_4667);
and U4866 (N_4866,N_4627,N_4659);
nand U4867 (N_4867,N_4705,N_4618);
nand U4868 (N_4868,N_4754,N_4772);
or U4869 (N_4869,N_4686,N_4746);
nand U4870 (N_4870,N_4795,N_4792);
and U4871 (N_4871,N_4678,N_4721);
and U4872 (N_4872,N_4780,N_4773);
nand U4873 (N_4873,N_4625,N_4662);
and U4874 (N_4874,N_4633,N_4677);
nand U4875 (N_4875,N_4753,N_4760);
and U4876 (N_4876,N_4624,N_4664);
and U4877 (N_4877,N_4727,N_4673);
and U4878 (N_4878,N_4697,N_4604);
and U4879 (N_4879,N_4620,N_4788);
or U4880 (N_4880,N_4714,N_4798);
nor U4881 (N_4881,N_4701,N_4735);
nand U4882 (N_4882,N_4747,N_4724);
or U4883 (N_4883,N_4631,N_4635);
nand U4884 (N_4884,N_4789,N_4771);
nand U4885 (N_4885,N_4736,N_4731);
nand U4886 (N_4886,N_4689,N_4730);
and U4887 (N_4887,N_4783,N_4644);
and U4888 (N_4888,N_4762,N_4750);
or U4889 (N_4889,N_4740,N_4652);
nor U4890 (N_4890,N_4695,N_4651);
nand U4891 (N_4891,N_4647,N_4646);
or U4892 (N_4892,N_4690,N_4709);
and U4893 (N_4893,N_4630,N_4716);
and U4894 (N_4894,N_4777,N_4638);
nand U4895 (N_4895,N_4784,N_4641);
nand U4896 (N_4896,N_4649,N_4629);
or U4897 (N_4897,N_4723,N_4779);
nor U4898 (N_4898,N_4799,N_4787);
nor U4899 (N_4899,N_4657,N_4609);
or U4900 (N_4900,N_4725,N_4784);
nand U4901 (N_4901,N_4727,N_4650);
nor U4902 (N_4902,N_4679,N_4788);
or U4903 (N_4903,N_4764,N_4772);
nor U4904 (N_4904,N_4680,N_4762);
and U4905 (N_4905,N_4637,N_4670);
nor U4906 (N_4906,N_4645,N_4698);
and U4907 (N_4907,N_4756,N_4694);
and U4908 (N_4908,N_4623,N_4609);
or U4909 (N_4909,N_4729,N_4639);
nor U4910 (N_4910,N_4609,N_4659);
or U4911 (N_4911,N_4661,N_4677);
nor U4912 (N_4912,N_4696,N_4694);
or U4913 (N_4913,N_4736,N_4782);
and U4914 (N_4914,N_4615,N_4614);
nor U4915 (N_4915,N_4707,N_4600);
or U4916 (N_4916,N_4718,N_4682);
and U4917 (N_4917,N_4710,N_4664);
or U4918 (N_4918,N_4781,N_4607);
nand U4919 (N_4919,N_4641,N_4702);
nor U4920 (N_4920,N_4768,N_4673);
nand U4921 (N_4921,N_4687,N_4724);
nand U4922 (N_4922,N_4654,N_4607);
nor U4923 (N_4923,N_4677,N_4683);
nand U4924 (N_4924,N_4798,N_4638);
nor U4925 (N_4925,N_4607,N_4658);
and U4926 (N_4926,N_4642,N_4626);
nand U4927 (N_4927,N_4640,N_4642);
nor U4928 (N_4928,N_4651,N_4738);
xnor U4929 (N_4929,N_4720,N_4776);
nand U4930 (N_4930,N_4755,N_4639);
and U4931 (N_4931,N_4688,N_4633);
and U4932 (N_4932,N_4653,N_4721);
or U4933 (N_4933,N_4758,N_4717);
and U4934 (N_4934,N_4782,N_4695);
or U4935 (N_4935,N_4760,N_4656);
nand U4936 (N_4936,N_4700,N_4621);
nor U4937 (N_4937,N_4747,N_4641);
nor U4938 (N_4938,N_4607,N_4693);
or U4939 (N_4939,N_4644,N_4700);
nand U4940 (N_4940,N_4703,N_4602);
or U4941 (N_4941,N_4718,N_4660);
nand U4942 (N_4942,N_4755,N_4750);
nand U4943 (N_4943,N_4722,N_4658);
nand U4944 (N_4944,N_4705,N_4684);
nor U4945 (N_4945,N_4736,N_4646);
and U4946 (N_4946,N_4723,N_4764);
or U4947 (N_4947,N_4656,N_4717);
nor U4948 (N_4948,N_4775,N_4641);
and U4949 (N_4949,N_4688,N_4737);
and U4950 (N_4950,N_4733,N_4642);
and U4951 (N_4951,N_4735,N_4643);
nor U4952 (N_4952,N_4739,N_4782);
nor U4953 (N_4953,N_4702,N_4723);
nor U4954 (N_4954,N_4711,N_4787);
and U4955 (N_4955,N_4737,N_4670);
nor U4956 (N_4956,N_4793,N_4788);
and U4957 (N_4957,N_4743,N_4779);
nand U4958 (N_4958,N_4645,N_4663);
or U4959 (N_4959,N_4689,N_4724);
or U4960 (N_4960,N_4635,N_4623);
nand U4961 (N_4961,N_4670,N_4770);
nand U4962 (N_4962,N_4736,N_4665);
and U4963 (N_4963,N_4762,N_4613);
nor U4964 (N_4964,N_4735,N_4777);
and U4965 (N_4965,N_4732,N_4716);
or U4966 (N_4966,N_4695,N_4622);
and U4967 (N_4967,N_4600,N_4765);
and U4968 (N_4968,N_4635,N_4784);
and U4969 (N_4969,N_4766,N_4608);
nor U4970 (N_4970,N_4602,N_4785);
nor U4971 (N_4971,N_4632,N_4620);
xor U4972 (N_4972,N_4757,N_4615);
and U4973 (N_4973,N_4611,N_4771);
or U4974 (N_4974,N_4648,N_4672);
nor U4975 (N_4975,N_4779,N_4679);
or U4976 (N_4976,N_4781,N_4775);
or U4977 (N_4977,N_4708,N_4705);
or U4978 (N_4978,N_4687,N_4720);
nor U4979 (N_4979,N_4643,N_4716);
and U4980 (N_4980,N_4779,N_4787);
nand U4981 (N_4981,N_4641,N_4692);
and U4982 (N_4982,N_4707,N_4773);
nand U4983 (N_4983,N_4768,N_4662);
and U4984 (N_4984,N_4755,N_4733);
or U4985 (N_4985,N_4658,N_4754);
nor U4986 (N_4986,N_4728,N_4727);
or U4987 (N_4987,N_4739,N_4605);
nor U4988 (N_4988,N_4774,N_4694);
nor U4989 (N_4989,N_4631,N_4623);
nor U4990 (N_4990,N_4632,N_4773);
nor U4991 (N_4991,N_4759,N_4774);
nand U4992 (N_4992,N_4673,N_4648);
or U4993 (N_4993,N_4794,N_4754);
or U4994 (N_4994,N_4760,N_4624);
nand U4995 (N_4995,N_4797,N_4671);
nand U4996 (N_4996,N_4790,N_4794);
nand U4997 (N_4997,N_4646,N_4607);
and U4998 (N_4998,N_4726,N_4636);
and U4999 (N_4999,N_4712,N_4695);
or U5000 (N_5000,N_4915,N_4988);
nand U5001 (N_5001,N_4943,N_4999);
nand U5002 (N_5002,N_4948,N_4854);
nor U5003 (N_5003,N_4875,N_4892);
nor U5004 (N_5004,N_4924,N_4886);
or U5005 (N_5005,N_4807,N_4871);
and U5006 (N_5006,N_4974,N_4955);
and U5007 (N_5007,N_4976,N_4899);
or U5008 (N_5008,N_4856,N_4897);
nor U5009 (N_5009,N_4929,N_4824);
nor U5010 (N_5010,N_4970,N_4939);
nand U5011 (N_5011,N_4872,N_4967);
nand U5012 (N_5012,N_4983,N_4878);
or U5013 (N_5013,N_4885,N_4819);
and U5014 (N_5014,N_4850,N_4989);
or U5015 (N_5015,N_4947,N_4866);
nor U5016 (N_5016,N_4858,N_4873);
or U5017 (N_5017,N_4839,N_4860);
nand U5018 (N_5018,N_4831,N_4890);
nor U5019 (N_5019,N_4905,N_4908);
or U5020 (N_5020,N_4887,N_4870);
and U5021 (N_5021,N_4906,N_4916);
or U5022 (N_5022,N_4863,N_4889);
xor U5023 (N_5023,N_4972,N_4898);
and U5024 (N_5024,N_4997,N_4953);
and U5025 (N_5025,N_4882,N_4944);
or U5026 (N_5026,N_4998,N_4954);
nand U5027 (N_5027,N_4923,N_4951);
nand U5028 (N_5028,N_4904,N_4816);
nor U5029 (N_5029,N_4865,N_4836);
nor U5030 (N_5030,N_4849,N_4909);
or U5031 (N_5031,N_4981,N_4968);
nor U5032 (N_5032,N_4920,N_4965);
nor U5033 (N_5033,N_4935,N_4940);
and U5034 (N_5034,N_4930,N_4803);
nor U5035 (N_5035,N_4817,N_4913);
or U5036 (N_5036,N_4814,N_4962);
nand U5037 (N_5037,N_4966,N_4928);
and U5038 (N_5038,N_4808,N_4977);
nor U5039 (N_5039,N_4861,N_4901);
nand U5040 (N_5040,N_4903,N_4868);
nor U5041 (N_5041,N_4827,N_4978);
and U5042 (N_5042,N_4867,N_4821);
nand U5043 (N_5043,N_4888,N_4949);
nor U5044 (N_5044,N_4937,N_4829);
or U5045 (N_5045,N_4809,N_4986);
nor U5046 (N_5046,N_4830,N_4879);
or U5047 (N_5047,N_4884,N_4802);
or U5048 (N_5048,N_4969,N_4975);
or U5049 (N_5049,N_4812,N_4843);
nor U5050 (N_5050,N_4841,N_4927);
and U5051 (N_5051,N_4848,N_4941);
and U5052 (N_5052,N_4893,N_4926);
nor U5053 (N_5053,N_4945,N_4996);
or U5054 (N_5054,N_4925,N_4917);
or U5055 (N_5055,N_4933,N_4846);
or U5056 (N_5056,N_4958,N_4956);
nand U5057 (N_5057,N_4826,N_4957);
or U5058 (N_5058,N_4993,N_4995);
xor U5059 (N_5059,N_4832,N_4852);
nand U5060 (N_5060,N_4874,N_4833);
and U5061 (N_5061,N_4869,N_4961);
nor U5062 (N_5062,N_4918,N_4804);
or U5063 (N_5063,N_4902,N_4971);
nand U5064 (N_5064,N_4881,N_4921);
and U5065 (N_5065,N_4805,N_4840);
nor U5066 (N_5066,N_4979,N_4952);
and U5067 (N_5067,N_4823,N_4876);
nor U5068 (N_5068,N_4801,N_4859);
xor U5069 (N_5069,N_4825,N_4991);
nand U5070 (N_5070,N_4914,N_4855);
or U5071 (N_5071,N_4851,N_4895);
nor U5072 (N_5072,N_4847,N_4837);
nor U5073 (N_5073,N_4835,N_4946);
or U5074 (N_5074,N_4992,N_4984);
nor U5075 (N_5075,N_4844,N_4896);
and U5076 (N_5076,N_4842,N_4942);
nor U5077 (N_5077,N_4964,N_4813);
xor U5078 (N_5078,N_4938,N_4911);
and U5079 (N_5079,N_4822,N_4838);
and U5080 (N_5080,N_4891,N_4932);
or U5081 (N_5081,N_4845,N_4880);
nand U5082 (N_5082,N_4985,N_4907);
or U5083 (N_5083,N_4811,N_4877);
or U5084 (N_5084,N_4818,N_4936);
nand U5085 (N_5085,N_4973,N_4862);
and U5086 (N_5086,N_4934,N_4806);
and U5087 (N_5087,N_4853,N_4820);
or U5088 (N_5088,N_4960,N_4959);
nand U5089 (N_5089,N_4800,N_4864);
nor U5090 (N_5090,N_4931,N_4987);
or U5091 (N_5091,N_4894,N_4910);
nand U5092 (N_5092,N_4919,N_4994);
or U5093 (N_5093,N_4834,N_4810);
nand U5094 (N_5094,N_4980,N_4900);
nor U5095 (N_5095,N_4912,N_4815);
nor U5096 (N_5096,N_4950,N_4990);
or U5097 (N_5097,N_4883,N_4963);
nand U5098 (N_5098,N_4922,N_4982);
or U5099 (N_5099,N_4828,N_4857);
or U5100 (N_5100,N_4980,N_4983);
or U5101 (N_5101,N_4942,N_4929);
or U5102 (N_5102,N_4891,N_4897);
nor U5103 (N_5103,N_4839,N_4974);
nand U5104 (N_5104,N_4803,N_4820);
nor U5105 (N_5105,N_4936,N_4850);
xor U5106 (N_5106,N_4999,N_4937);
and U5107 (N_5107,N_4892,N_4942);
or U5108 (N_5108,N_4801,N_4964);
and U5109 (N_5109,N_4822,N_4846);
nor U5110 (N_5110,N_4957,N_4880);
and U5111 (N_5111,N_4836,N_4803);
nand U5112 (N_5112,N_4961,N_4936);
and U5113 (N_5113,N_4982,N_4854);
nor U5114 (N_5114,N_4879,N_4974);
nand U5115 (N_5115,N_4876,N_4921);
and U5116 (N_5116,N_4889,N_4897);
nor U5117 (N_5117,N_4994,N_4881);
nand U5118 (N_5118,N_4827,N_4822);
and U5119 (N_5119,N_4990,N_4862);
nor U5120 (N_5120,N_4968,N_4974);
xnor U5121 (N_5121,N_4984,N_4835);
nor U5122 (N_5122,N_4863,N_4955);
nand U5123 (N_5123,N_4990,N_4995);
nor U5124 (N_5124,N_4967,N_4924);
nor U5125 (N_5125,N_4963,N_4972);
nor U5126 (N_5126,N_4894,N_4898);
or U5127 (N_5127,N_4946,N_4985);
and U5128 (N_5128,N_4894,N_4983);
nand U5129 (N_5129,N_4806,N_4979);
or U5130 (N_5130,N_4998,N_4938);
nor U5131 (N_5131,N_4994,N_4862);
nor U5132 (N_5132,N_4803,N_4872);
and U5133 (N_5133,N_4956,N_4918);
nor U5134 (N_5134,N_4892,N_4953);
nor U5135 (N_5135,N_4827,N_4810);
or U5136 (N_5136,N_4828,N_4928);
nor U5137 (N_5137,N_4859,N_4892);
or U5138 (N_5138,N_4825,N_4924);
nor U5139 (N_5139,N_4991,N_4987);
nor U5140 (N_5140,N_4924,N_4900);
nand U5141 (N_5141,N_4873,N_4808);
and U5142 (N_5142,N_4888,N_4821);
or U5143 (N_5143,N_4931,N_4806);
nor U5144 (N_5144,N_4948,N_4974);
nand U5145 (N_5145,N_4991,N_4942);
nand U5146 (N_5146,N_4956,N_4802);
nor U5147 (N_5147,N_4957,N_4966);
or U5148 (N_5148,N_4872,N_4858);
and U5149 (N_5149,N_4893,N_4896);
or U5150 (N_5150,N_4887,N_4956);
and U5151 (N_5151,N_4973,N_4807);
nand U5152 (N_5152,N_4915,N_4851);
or U5153 (N_5153,N_4989,N_4861);
and U5154 (N_5154,N_4874,N_4954);
and U5155 (N_5155,N_4970,N_4825);
nor U5156 (N_5156,N_4967,N_4895);
or U5157 (N_5157,N_4888,N_4950);
nand U5158 (N_5158,N_4864,N_4935);
nand U5159 (N_5159,N_4858,N_4930);
or U5160 (N_5160,N_4895,N_4972);
nand U5161 (N_5161,N_4807,N_4910);
nor U5162 (N_5162,N_4858,N_4993);
nand U5163 (N_5163,N_4922,N_4816);
or U5164 (N_5164,N_4944,N_4865);
nand U5165 (N_5165,N_4882,N_4959);
or U5166 (N_5166,N_4851,N_4884);
or U5167 (N_5167,N_4994,N_4930);
nor U5168 (N_5168,N_4896,N_4888);
nor U5169 (N_5169,N_4806,N_4964);
nor U5170 (N_5170,N_4850,N_4824);
or U5171 (N_5171,N_4853,N_4917);
nand U5172 (N_5172,N_4961,N_4892);
and U5173 (N_5173,N_4979,N_4893);
or U5174 (N_5174,N_4977,N_4968);
or U5175 (N_5175,N_4909,N_4898);
nand U5176 (N_5176,N_4954,N_4860);
nand U5177 (N_5177,N_4991,N_4984);
and U5178 (N_5178,N_4915,N_4844);
or U5179 (N_5179,N_4802,N_4980);
or U5180 (N_5180,N_4849,N_4801);
nor U5181 (N_5181,N_4803,N_4906);
nor U5182 (N_5182,N_4933,N_4960);
nor U5183 (N_5183,N_4909,N_4838);
nand U5184 (N_5184,N_4945,N_4843);
or U5185 (N_5185,N_4850,N_4839);
nor U5186 (N_5186,N_4890,N_4982);
or U5187 (N_5187,N_4935,N_4866);
nor U5188 (N_5188,N_4958,N_4928);
nand U5189 (N_5189,N_4831,N_4820);
nand U5190 (N_5190,N_4936,N_4949);
and U5191 (N_5191,N_4895,N_4912);
nand U5192 (N_5192,N_4881,N_4915);
xnor U5193 (N_5193,N_4993,N_4845);
nand U5194 (N_5194,N_4967,N_4857);
or U5195 (N_5195,N_4825,N_4927);
nor U5196 (N_5196,N_4920,N_4984);
and U5197 (N_5197,N_4861,N_4999);
nand U5198 (N_5198,N_4988,N_4883);
or U5199 (N_5199,N_4907,N_4867);
and U5200 (N_5200,N_5119,N_5060);
nor U5201 (N_5201,N_5098,N_5195);
nor U5202 (N_5202,N_5124,N_5061);
xor U5203 (N_5203,N_5084,N_5174);
and U5204 (N_5204,N_5029,N_5130);
nand U5205 (N_5205,N_5015,N_5095);
and U5206 (N_5206,N_5148,N_5050);
and U5207 (N_5207,N_5137,N_5134);
or U5208 (N_5208,N_5080,N_5022);
and U5209 (N_5209,N_5139,N_5069);
or U5210 (N_5210,N_5155,N_5018);
or U5211 (N_5211,N_5164,N_5064);
and U5212 (N_5212,N_5034,N_5036);
and U5213 (N_5213,N_5016,N_5070);
nor U5214 (N_5214,N_5120,N_5152);
nor U5215 (N_5215,N_5051,N_5063);
nand U5216 (N_5216,N_5025,N_5185);
and U5217 (N_5217,N_5177,N_5001);
nand U5218 (N_5218,N_5062,N_5048);
nor U5219 (N_5219,N_5165,N_5189);
or U5220 (N_5220,N_5076,N_5187);
and U5221 (N_5221,N_5154,N_5083);
or U5222 (N_5222,N_5169,N_5089);
or U5223 (N_5223,N_5026,N_5009);
nand U5224 (N_5224,N_5047,N_5088);
nand U5225 (N_5225,N_5106,N_5144);
nand U5226 (N_5226,N_5162,N_5086);
nor U5227 (N_5227,N_5149,N_5003);
nor U5228 (N_5228,N_5030,N_5156);
or U5229 (N_5229,N_5056,N_5143);
nor U5230 (N_5230,N_5075,N_5138);
nand U5231 (N_5231,N_5127,N_5002);
or U5232 (N_5232,N_5140,N_5142);
nor U5233 (N_5233,N_5090,N_5104);
or U5234 (N_5234,N_5053,N_5163);
and U5235 (N_5235,N_5128,N_5096);
nand U5236 (N_5236,N_5122,N_5173);
or U5237 (N_5237,N_5091,N_5166);
or U5238 (N_5238,N_5093,N_5188);
or U5239 (N_5239,N_5125,N_5150);
or U5240 (N_5240,N_5109,N_5017);
nor U5241 (N_5241,N_5181,N_5014);
and U5242 (N_5242,N_5141,N_5057);
or U5243 (N_5243,N_5184,N_5147);
nor U5244 (N_5244,N_5191,N_5146);
and U5245 (N_5245,N_5035,N_5028);
nand U5246 (N_5246,N_5092,N_5197);
nor U5247 (N_5247,N_5082,N_5079);
or U5248 (N_5248,N_5081,N_5037);
nand U5249 (N_5249,N_5193,N_5186);
nand U5250 (N_5250,N_5054,N_5033);
and U5251 (N_5251,N_5123,N_5020);
or U5252 (N_5252,N_5021,N_5041);
nand U5253 (N_5253,N_5110,N_5010);
nor U5254 (N_5254,N_5102,N_5097);
and U5255 (N_5255,N_5077,N_5115);
nor U5256 (N_5256,N_5179,N_5004);
xnor U5257 (N_5257,N_5199,N_5032);
nand U5258 (N_5258,N_5170,N_5135);
or U5259 (N_5259,N_5019,N_5118);
or U5260 (N_5260,N_5111,N_5176);
and U5261 (N_5261,N_5129,N_5011);
and U5262 (N_5262,N_5024,N_5145);
nand U5263 (N_5263,N_5023,N_5121);
and U5264 (N_5264,N_5159,N_5132);
or U5265 (N_5265,N_5108,N_5105);
nand U5266 (N_5266,N_5043,N_5113);
or U5267 (N_5267,N_5192,N_5087);
nor U5268 (N_5268,N_5196,N_5073);
and U5269 (N_5269,N_5008,N_5042);
nand U5270 (N_5270,N_5099,N_5044);
nand U5271 (N_5271,N_5068,N_5103);
nand U5272 (N_5272,N_5085,N_5178);
nand U5273 (N_5273,N_5151,N_5074);
nor U5274 (N_5274,N_5067,N_5031);
or U5275 (N_5275,N_5027,N_5136);
nand U5276 (N_5276,N_5052,N_5059);
or U5277 (N_5277,N_5194,N_5126);
nor U5278 (N_5278,N_5078,N_5157);
nand U5279 (N_5279,N_5040,N_5112);
and U5280 (N_5280,N_5171,N_5116);
and U5281 (N_5281,N_5158,N_5172);
nor U5282 (N_5282,N_5100,N_5045);
nor U5283 (N_5283,N_5005,N_5055);
and U5284 (N_5284,N_5058,N_5101);
and U5285 (N_5285,N_5049,N_5038);
or U5286 (N_5286,N_5007,N_5168);
and U5287 (N_5287,N_5190,N_5167);
or U5288 (N_5288,N_5039,N_5071);
or U5289 (N_5289,N_5094,N_5000);
nand U5290 (N_5290,N_5065,N_5182);
and U5291 (N_5291,N_5006,N_5114);
nand U5292 (N_5292,N_5161,N_5153);
nand U5293 (N_5293,N_5072,N_5133);
or U5294 (N_5294,N_5117,N_5012);
or U5295 (N_5295,N_5046,N_5180);
xnor U5296 (N_5296,N_5198,N_5183);
nand U5297 (N_5297,N_5175,N_5107);
and U5298 (N_5298,N_5066,N_5013);
and U5299 (N_5299,N_5131,N_5160);
nand U5300 (N_5300,N_5014,N_5037);
and U5301 (N_5301,N_5103,N_5076);
and U5302 (N_5302,N_5180,N_5056);
nand U5303 (N_5303,N_5101,N_5005);
and U5304 (N_5304,N_5189,N_5085);
nand U5305 (N_5305,N_5004,N_5076);
and U5306 (N_5306,N_5161,N_5063);
nand U5307 (N_5307,N_5101,N_5085);
and U5308 (N_5308,N_5108,N_5000);
or U5309 (N_5309,N_5118,N_5140);
and U5310 (N_5310,N_5157,N_5015);
or U5311 (N_5311,N_5019,N_5028);
or U5312 (N_5312,N_5086,N_5041);
and U5313 (N_5313,N_5144,N_5063);
nor U5314 (N_5314,N_5080,N_5072);
nor U5315 (N_5315,N_5176,N_5033);
nor U5316 (N_5316,N_5173,N_5090);
or U5317 (N_5317,N_5079,N_5097);
nand U5318 (N_5318,N_5039,N_5017);
and U5319 (N_5319,N_5145,N_5176);
nand U5320 (N_5320,N_5139,N_5173);
and U5321 (N_5321,N_5071,N_5014);
nor U5322 (N_5322,N_5067,N_5128);
nand U5323 (N_5323,N_5060,N_5093);
and U5324 (N_5324,N_5181,N_5115);
or U5325 (N_5325,N_5143,N_5177);
nand U5326 (N_5326,N_5145,N_5149);
or U5327 (N_5327,N_5057,N_5131);
and U5328 (N_5328,N_5053,N_5173);
nand U5329 (N_5329,N_5084,N_5141);
nand U5330 (N_5330,N_5149,N_5161);
or U5331 (N_5331,N_5135,N_5166);
xor U5332 (N_5332,N_5162,N_5163);
nand U5333 (N_5333,N_5092,N_5040);
and U5334 (N_5334,N_5135,N_5079);
xor U5335 (N_5335,N_5016,N_5184);
and U5336 (N_5336,N_5125,N_5080);
or U5337 (N_5337,N_5090,N_5159);
and U5338 (N_5338,N_5066,N_5153);
or U5339 (N_5339,N_5030,N_5099);
or U5340 (N_5340,N_5187,N_5158);
and U5341 (N_5341,N_5071,N_5157);
nand U5342 (N_5342,N_5183,N_5188);
or U5343 (N_5343,N_5098,N_5055);
and U5344 (N_5344,N_5178,N_5173);
nand U5345 (N_5345,N_5144,N_5119);
nand U5346 (N_5346,N_5117,N_5078);
and U5347 (N_5347,N_5190,N_5044);
xnor U5348 (N_5348,N_5000,N_5059);
nor U5349 (N_5349,N_5197,N_5115);
or U5350 (N_5350,N_5144,N_5070);
nand U5351 (N_5351,N_5074,N_5119);
nor U5352 (N_5352,N_5041,N_5045);
or U5353 (N_5353,N_5078,N_5143);
or U5354 (N_5354,N_5163,N_5164);
nand U5355 (N_5355,N_5001,N_5114);
and U5356 (N_5356,N_5136,N_5041);
nor U5357 (N_5357,N_5065,N_5104);
or U5358 (N_5358,N_5139,N_5042);
nor U5359 (N_5359,N_5161,N_5016);
and U5360 (N_5360,N_5048,N_5119);
nand U5361 (N_5361,N_5044,N_5100);
and U5362 (N_5362,N_5065,N_5143);
or U5363 (N_5363,N_5191,N_5151);
xor U5364 (N_5364,N_5148,N_5103);
or U5365 (N_5365,N_5129,N_5034);
or U5366 (N_5366,N_5135,N_5143);
and U5367 (N_5367,N_5144,N_5073);
and U5368 (N_5368,N_5130,N_5033);
xnor U5369 (N_5369,N_5153,N_5076);
nor U5370 (N_5370,N_5025,N_5101);
nand U5371 (N_5371,N_5186,N_5102);
nor U5372 (N_5372,N_5011,N_5015);
nor U5373 (N_5373,N_5154,N_5189);
and U5374 (N_5374,N_5062,N_5003);
nor U5375 (N_5375,N_5119,N_5094);
nand U5376 (N_5376,N_5147,N_5156);
nand U5377 (N_5377,N_5088,N_5074);
and U5378 (N_5378,N_5051,N_5020);
nand U5379 (N_5379,N_5045,N_5122);
and U5380 (N_5380,N_5149,N_5195);
nor U5381 (N_5381,N_5124,N_5135);
or U5382 (N_5382,N_5143,N_5137);
nor U5383 (N_5383,N_5045,N_5081);
nand U5384 (N_5384,N_5011,N_5097);
nand U5385 (N_5385,N_5016,N_5169);
and U5386 (N_5386,N_5198,N_5182);
and U5387 (N_5387,N_5067,N_5057);
nor U5388 (N_5388,N_5199,N_5197);
xnor U5389 (N_5389,N_5100,N_5024);
nor U5390 (N_5390,N_5197,N_5102);
and U5391 (N_5391,N_5030,N_5054);
nand U5392 (N_5392,N_5152,N_5042);
and U5393 (N_5393,N_5054,N_5060);
nand U5394 (N_5394,N_5041,N_5176);
and U5395 (N_5395,N_5135,N_5188);
and U5396 (N_5396,N_5126,N_5002);
nor U5397 (N_5397,N_5065,N_5049);
nor U5398 (N_5398,N_5118,N_5198);
and U5399 (N_5399,N_5173,N_5126);
and U5400 (N_5400,N_5359,N_5345);
and U5401 (N_5401,N_5370,N_5323);
or U5402 (N_5402,N_5290,N_5303);
or U5403 (N_5403,N_5230,N_5333);
nand U5404 (N_5404,N_5352,N_5377);
nand U5405 (N_5405,N_5311,N_5291);
and U5406 (N_5406,N_5374,N_5305);
xnor U5407 (N_5407,N_5320,N_5245);
or U5408 (N_5408,N_5331,N_5243);
nor U5409 (N_5409,N_5354,N_5286);
nand U5410 (N_5410,N_5375,N_5228);
nor U5411 (N_5411,N_5205,N_5337);
or U5412 (N_5412,N_5244,N_5292);
nand U5413 (N_5413,N_5268,N_5317);
nand U5414 (N_5414,N_5269,N_5262);
and U5415 (N_5415,N_5253,N_5260);
or U5416 (N_5416,N_5240,N_5294);
or U5417 (N_5417,N_5275,N_5288);
nand U5418 (N_5418,N_5383,N_5273);
or U5419 (N_5419,N_5369,N_5381);
and U5420 (N_5420,N_5327,N_5256);
or U5421 (N_5421,N_5324,N_5224);
and U5422 (N_5422,N_5254,N_5242);
nor U5423 (N_5423,N_5271,N_5364);
nor U5424 (N_5424,N_5239,N_5236);
xnor U5425 (N_5425,N_5265,N_5299);
nor U5426 (N_5426,N_5241,N_5343);
xnor U5427 (N_5427,N_5201,N_5363);
nor U5428 (N_5428,N_5223,N_5225);
and U5429 (N_5429,N_5306,N_5391);
nor U5430 (N_5430,N_5274,N_5332);
and U5431 (N_5431,N_5379,N_5367);
or U5432 (N_5432,N_5221,N_5395);
nor U5433 (N_5433,N_5272,N_5348);
nor U5434 (N_5434,N_5368,N_5214);
nor U5435 (N_5435,N_5233,N_5284);
and U5436 (N_5436,N_5362,N_5296);
or U5437 (N_5437,N_5219,N_5285);
nor U5438 (N_5438,N_5289,N_5335);
nor U5439 (N_5439,N_5339,N_5315);
or U5440 (N_5440,N_5338,N_5279);
nand U5441 (N_5441,N_5227,N_5267);
nor U5442 (N_5442,N_5329,N_5378);
and U5443 (N_5443,N_5394,N_5220);
or U5444 (N_5444,N_5257,N_5204);
nand U5445 (N_5445,N_5390,N_5347);
and U5446 (N_5446,N_5229,N_5341);
nor U5447 (N_5447,N_5218,N_5388);
nand U5448 (N_5448,N_5266,N_5358);
nand U5449 (N_5449,N_5261,N_5360);
nand U5450 (N_5450,N_5319,N_5237);
nand U5451 (N_5451,N_5309,N_5313);
and U5452 (N_5452,N_5246,N_5396);
and U5453 (N_5453,N_5316,N_5304);
and U5454 (N_5454,N_5353,N_5312);
nand U5455 (N_5455,N_5384,N_5344);
nor U5456 (N_5456,N_5307,N_5398);
nand U5457 (N_5457,N_5356,N_5278);
nor U5458 (N_5458,N_5361,N_5212);
nor U5459 (N_5459,N_5231,N_5297);
or U5460 (N_5460,N_5302,N_5216);
and U5461 (N_5461,N_5211,N_5397);
nor U5462 (N_5462,N_5217,N_5203);
or U5463 (N_5463,N_5258,N_5282);
and U5464 (N_5464,N_5200,N_5264);
or U5465 (N_5465,N_5371,N_5365);
nand U5466 (N_5466,N_5399,N_5330);
nor U5467 (N_5467,N_5259,N_5300);
nor U5468 (N_5468,N_5222,N_5340);
or U5469 (N_5469,N_5393,N_5382);
and U5470 (N_5470,N_5342,N_5366);
nand U5471 (N_5471,N_5336,N_5208);
and U5472 (N_5472,N_5326,N_5255);
and U5473 (N_5473,N_5349,N_5318);
or U5474 (N_5474,N_5380,N_5252);
xor U5475 (N_5475,N_5346,N_5276);
nand U5476 (N_5476,N_5357,N_5226);
and U5477 (N_5477,N_5283,N_5351);
nand U5478 (N_5478,N_5301,N_5373);
and U5479 (N_5479,N_5251,N_5250);
or U5480 (N_5480,N_5281,N_5389);
nand U5481 (N_5481,N_5248,N_5328);
or U5482 (N_5482,N_5280,N_5207);
nor U5483 (N_5483,N_5209,N_5322);
nand U5484 (N_5484,N_5295,N_5263);
and U5485 (N_5485,N_5235,N_5385);
or U5486 (N_5486,N_5376,N_5215);
and U5487 (N_5487,N_5325,N_5386);
or U5488 (N_5488,N_5249,N_5206);
or U5489 (N_5489,N_5202,N_5321);
nand U5490 (N_5490,N_5355,N_5213);
or U5491 (N_5491,N_5298,N_5234);
and U5492 (N_5492,N_5232,N_5238);
or U5493 (N_5493,N_5287,N_5277);
nand U5494 (N_5494,N_5270,N_5293);
nand U5495 (N_5495,N_5334,N_5350);
nand U5496 (N_5496,N_5308,N_5247);
nand U5497 (N_5497,N_5392,N_5310);
or U5498 (N_5498,N_5372,N_5210);
nand U5499 (N_5499,N_5387,N_5314);
and U5500 (N_5500,N_5352,N_5234);
xor U5501 (N_5501,N_5256,N_5245);
nand U5502 (N_5502,N_5282,N_5243);
nor U5503 (N_5503,N_5362,N_5221);
nor U5504 (N_5504,N_5285,N_5381);
xor U5505 (N_5505,N_5231,N_5292);
nor U5506 (N_5506,N_5377,N_5297);
nor U5507 (N_5507,N_5297,N_5371);
nor U5508 (N_5508,N_5347,N_5290);
xor U5509 (N_5509,N_5384,N_5379);
and U5510 (N_5510,N_5378,N_5252);
nor U5511 (N_5511,N_5363,N_5300);
and U5512 (N_5512,N_5271,N_5395);
and U5513 (N_5513,N_5395,N_5241);
or U5514 (N_5514,N_5334,N_5211);
xor U5515 (N_5515,N_5206,N_5350);
nand U5516 (N_5516,N_5295,N_5392);
nor U5517 (N_5517,N_5200,N_5210);
nor U5518 (N_5518,N_5202,N_5326);
and U5519 (N_5519,N_5288,N_5351);
and U5520 (N_5520,N_5271,N_5326);
or U5521 (N_5521,N_5207,N_5219);
nand U5522 (N_5522,N_5214,N_5247);
or U5523 (N_5523,N_5242,N_5255);
nand U5524 (N_5524,N_5325,N_5290);
nand U5525 (N_5525,N_5294,N_5378);
nand U5526 (N_5526,N_5280,N_5388);
nand U5527 (N_5527,N_5316,N_5352);
or U5528 (N_5528,N_5265,N_5319);
nor U5529 (N_5529,N_5236,N_5381);
nor U5530 (N_5530,N_5340,N_5276);
nand U5531 (N_5531,N_5314,N_5247);
and U5532 (N_5532,N_5292,N_5366);
or U5533 (N_5533,N_5308,N_5342);
or U5534 (N_5534,N_5373,N_5350);
or U5535 (N_5535,N_5221,N_5291);
nand U5536 (N_5536,N_5371,N_5201);
nand U5537 (N_5537,N_5229,N_5230);
and U5538 (N_5538,N_5285,N_5335);
nand U5539 (N_5539,N_5328,N_5272);
and U5540 (N_5540,N_5268,N_5289);
or U5541 (N_5541,N_5281,N_5283);
or U5542 (N_5542,N_5333,N_5335);
nor U5543 (N_5543,N_5271,N_5301);
nand U5544 (N_5544,N_5394,N_5333);
nor U5545 (N_5545,N_5314,N_5257);
xnor U5546 (N_5546,N_5326,N_5346);
nor U5547 (N_5547,N_5343,N_5276);
or U5548 (N_5548,N_5396,N_5368);
and U5549 (N_5549,N_5219,N_5235);
nor U5550 (N_5550,N_5271,N_5249);
nor U5551 (N_5551,N_5325,N_5313);
and U5552 (N_5552,N_5210,N_5396);
and U5553 (N_5553,N_5212,N_5364);
and U5554 (N_5554,N_5388,N_5380);
nand U5555 (N_5555,N_5284,N_5315);
nand U5556 (N_5556,N_5398,N_5291);
nand U5557 (N_5557,N_5243,N_5338);
or U5558 (N_5558,N_5384,N_5371);
or U5559 (N_5559,N_5299,N_5388);
or U5560 (N_5560,N_5351,N_5379);
and U5561 (N_5561,N_5370,N_5379);
nor U5562 (N_5562,N_5299,N_5253);
nor U5563 (N_5563,N_5299,N_5383);
and U5564 (N_5564,N_5222,N_5369);
or U5565 (N_5565,N_5202,N_5380);
and U5566 (N_5566,N_5235,N_5239);
or U5567 (N_5567,N_5395,N_5240);
nor U5568 (N_5568,N_5208,N_5376);
nand U5569 (N_5569,N_5392,N_5249);
and U5570 (N_5570,N_5379,N_5203);
and U5571 (N_5571,N_5266,N_5316);
nand U5572 (N_5572,N_5306,N_5264);
xor U5573 (N_5573,N_5220,N_5314);
nor U5574 (N_5574,N_5218,N_5264);
nor U5575 (N_5575,N_5342,N_5254);
or U5576 (N_5576,N_5335,N_5252);
nand U5577 (N_5577,N_5258,N_5204);
or U5578 (N_5578,N_5285,N_5365);
or U5579 (N_5579,N_5379,N_5386);
and U5580 (N_5580,N_5289,N_5269);
or U5581 (N_5581,N_5213,N_5245);
or U5582 (N_5582,N_5237,N_5368);
nor U5583 (N_5583,N_5320,N_5224);
or U5584 (N_5584,N_5283,N_5234);
nand U5585 (N_5585,N_5379,N_5378);
or U5586 (N_5586,N_5230,N_5311);
nor U5587 (N_5587,N_5354,N_5313);
or U5588 (N_5588,N_5348,N_5291);
nand U5589 (N_5589,N_5260,N_5344);
nor U5590 (N_5590,N_5388,N_5335);
and U5591 (N_5591,N_5335,N_5321);
and U5592 (N_5592,N_5319,N_5235);
nor U5593 (N_5593,N_5202,N_5398);
nand U5594 (N_5594,N_5247,N_5334);
and U5595 (N_5595,N_5274,N_5252);
nor U5596 (N_5596,N_5248,N_5393);
nor U5597 (N_5597,N_5200,N_5369);
and U5598 (N_5598,N_5380,N_5382);
nor U5599 (N_5599,N_5328,N_5354);
xor U5600 (N_5600,N_5509,N_5495);
and U5601 (N_5601,N_5457,N_5466);
nand U5602 (N_5602,N_5502,N_5482);
or U5603 (N_5603,N_5467,N_5551);
and U5604 (N_5604,N_5591,N_5487);
nor U5605 (N_5605,N_5492,N_5571);
or U5606 (N_5606,N_5557,N_5471);
nand U5607 (N_5607,N_5519,N_5576);
and U5608 (N_5608,N_5419,N_5527);
nor U5609 (N_5609,N_5564,N_5444);
or U5610 (N_5610,N_5511,N_5448);
or U5611 (N_5611,N_5453,N_5418);
nand U5612 (N_5612,N_5479,N_5537);
nor U5613 (N_5613,N_5447,N_5497);
or U5614 (N_5614,N_5589,N_5553);
or U5615 (N_5615,N_5508,N_5540);
and U5616 (N_5616,N_5555,N_5427);
or U5617 (N_5617,N_5547,N_5524);
nor U5618 (N_5618,N_5568,N_5562);
or U5619 (N_5619,N_5599,N_5405);
nand U5620 (N_5620,N_5433,N_5480);
nand U5621 (N_5621,N_5516,N_5408);
xnor U5622 (N_5622,N_5422,N_5426);
nor U5623 (N_5623,N_5460,N_5545);
nand U5624 (N_5624,N_5563,N_5401);
nand U5625 (N_5625,N_5507,N_5512);
and U5626 (N_5626,N_5446,N_5424);
nand U5627 (N_5627,N_5420,N_5456);
nand U5628 (N_5628,N_5543,N_5485);
nor U5629 (N_5629,N_5423,N_5577);
or U5630 (N_5630,N_5435,N_5454);
or U5631 (N_5631,N_5569,N_5469);
nand U5632 (N_5632,N_5414,N_5526);
or U5633 (N_5633,N_5538,N_5406);
nand U5634 (N_5634,N_5499,N_5478);
and U5635 (N_5635,N_5410,N_5597);
or U5636 (N_5636,N_5494,N_5461);
nand U5637 (N_5637,N_5596,N_5458);
and U5638 (N_5638,N_5522,N_5473);
nand U5639 (N_5639,N_5443,N_5504);
nor U5640 (N_5640,N_5415,N_5536);
or U5641 (N_5641,N_5412,N_5585);
nor U5642 (N_5642,N_5486,N_5490);
and U5643 (N_5643,N_5430,N_5594);
or U5644 (N_5644,N_5409,N_5592);
nor U5645 (N_5645,N_5438,N_5500);
or U5646 (N_5646,N_5575,N_5570);
and U5647 (N_5647,N_5400,N_5528);
or U5648 (N_5648,N_5450,N_5407);
and U5649 (N_5649,N_5417,N_5581);
and U5650 (N_5650,N_5558,N_5488);
and U5651 (N_5651,N_5404,N_5539);
or U5652 (N_5652,N_5574,N_5525);
nand U5653 (N_5653,N_5403,N_5477);
or U5654 (N_5654,N_5475,N_5428);
nor U5655 (N_5655,N_5464,N_5421);
nor U5656 (N_5656,N_5465,N_5436);
nand U5657 (N_5657,N_5529,N_5449);
xor U5658 (N_5658,N_5532,N_5561);
nor U5659 (N_5659,N_5432,N_5484);
and U5660 (N_5660,N_5565,N_5552);
and U5661 (N_5661,N_5546,N_5442);
nor U5662 (N_5662,N_5550,N_5413);
nor U5663 (N_5663,N_5411,N_5593);
nor U5664 (N_5664,N_5518,N_5513);
or U5665 (N_5665,N_5584,N_5566);
nor U5666 (N_5666,N_5425,N_5580);
nor U5667 (N_5667,N_5431,N_5481);
nand U5668 (N_5668,N_5541,N_5533);
and U5669 (N_5669,N_5556,N_5587);
or U5670 (N_5670,N_5462,N_5554);
nor U5671 (N_5671,N_5586,N_5489);
nand U5672 (N_5672,N_5437,N_5514);
nand U5673 (N_5673,N_5416,N_5493);
or U5674 (N_5674,N_5451,N_5501);
or U5675 (N_5675,N_5463,N_5583);
nand U5676 (N_5676,N_5441,N_5523);
nand U5677 (N_5677,N_5595,N_5440);
nand U5678 (N_5678,N_5505,N_5483);
or U5679 (N_5679,N_5498,N_5503);
nand U5680 (N_5680,N_5567,N_5506);
nand U5681 (N_5681,N_5582,N_5470);
or U5682 (N_5682,N_5572,N_5531);
and U5683 (N_5683,N_5517,N_5530);
and U5684 (N_5684,N_5445,N_5559);
nor U5685 (N_5685,N_5542,N_5474);
nor U5686 (N_5686,N_5472,N_5452);
nand U5687 (N_5687,N_5496,N_5434);
nand U5688 (N_5688,N_5429,N_5590);
nand U5689 (N_5689,N_5515,N_5491);
or U5690 (N_5690,N_5459,N_5534);
nand U5691 (N_5691,N_5579,N_5468);
nor U5692 (N_5692,N_5598,N_5578);
nor U5693 (N_5693,N_5535,N_5455);
nor U5694 (N_5694,N_5520,N_5521);
nand U5695 (N_5695,N_5560,N_5510);
nor U5696 (N_5696,N_5439,N_5402);
and U5697 (N_5697,N_5544,N_5548);
nand U5698 (N_5698,N_5588,N_5549);
nor U5699 (N_5699,N_5573,N_5476);
nor U5700 (N_5700,N_5534,N_5506);
nand U5701 (N_5701,N_5581,N_5462);
or U5702 (N_5702,N_5488,N_5552);
and U5703 (N_5703,N_5587,N_5585);
and U5704 (N_5704,N_5552,N_5582);
nand U5705 (N_5705,N_5562,N_5494);
or U5706 (N_5706,N_5507,N_5572);
nor U5707 (N_5707,N_5490,N_5529);
nand U5708 (N_5708,N_5459,N_5498);
and U5709 (N_5709,N_5466,N_5580);
nand U5710 (N_5710,N_5525,N_5537);
nand U5711 (N_5711,N_5421,N_5433);
nand U5712 (N_5712,N_5422,N_5535);
nor U5713 (N_5713,N_5458,N_5587);
nor U5714 (N_5714,N_5471,N_5571);
and U5715 (N_5715,N_5407,N_5547);
and U5716 (N_5716,N_5401,N_5466);
nand U5717 (N_5717,N_5479,N_5534);
and U5718 (N_5718,N_5404,N_5457);
and U5719 (N_5719,N_5501,N_5552);
and U5720 (N_5720,N_5560,N_5495);
nor U5721 (N_5721,N_5520,N_5580);
and U5722 (N_5722,N_5544,N_5435);
nor U5723 (N_5723,N_5423,N_5521);
nor U5724 (N_5724,N_5507,N_5458);
nor U5725 (N_5725,N_5441,N_5599);
nand U5726 (N_5726,N_5490,N_5493);
nand U5727 (N_5727,N_5424,N_5410);
nand U5728 (N_5728,N_5427,N_5418);
xnor U5729 (N_5729,N_5400,N_5462);
or U5730 (N_5730,N_5437,N_5575);
or U5731 (N_5731,N_5563,N_5517);
nor U5732 (N_5732,N_5421,N_5582);
and U5733 (N_5733,N_5525,N_5425);
and U5734 (N_5734,N_5479,N_5473);
nand U5735 (N_5735,N_5486,N_5485);
or U5736 (N_5736,N_5533,N_5540);
and U5737 (N_5737,N_5427,N_5521);
nor U5738 (N_5738,N_5455,N_5400);
and U5739 (N_5739,N_5472,N_5564);
nor U5740 (N_5740,N_5506,N_5473);
or U5741 (N_5741,N_5533,N_5473);
nor U5742 (N_5742,N_5444,N_5434);
and U5743 (N_5743,N_5404,N_5591);
or U5744 (N_5744,N_5499,N_5583);
or U5745 (N_5745,N_5526,N_5476);
xnor U5746 (N_5746,N_5590,N_5460);
or U5747 (N_5747,N_5422,N_5587);
or U5748 (N_5748,N_5593,N_5433);
and U5749 (N_5749,N_5419,N_5475);
nand U5750 (N_5750,N_5480,N_5500);
and U5751 (N_5751,N_5545,N_5576);
nand U5752 (N_5752,N_5555,N_5473);
nand U5753 (N_5753,N_5460,N_5499);
nor U5754 (N_5754,N_5577,N_5552);
nand U5755 (N_5755,N_5443,N_5580);
and U5756 (N_5756,N_5565,N_5446);
xor U5757 (N_5757,N_5402,N_5518);
nand U5758 (N_5758,N_5430,N_5540);
or U5759 (N_5759,N_5503,N_5517);
and U5760 (N_5760,N_5550,N_5470);
nand U5761 (N_5761,N_5536,N_5562);
and U5762 (N_5762,N_5560,N_5547);
xor U5763 (N_5763,N_5410,N_5461);
or U5764 (N_5764,N_5555,N_5546);
nand U5765 (N_5765,N_5479,N_5471);
or U5766 (N_5766,N_5554,N_5406);
or U5767 (N_5767,N_5555,N_5586);
or U5768 (N_5768,N_5580,N_5444);
and U5769 (N_5769,N_5593,N_5426);
or U5770 (N_5770,N_5488,N_5480);
nand U5771 (N_5771,N_5485,N_5420);
and U5772 (N_5772,N_5547,N_5433);
nor U5773 (N_5773,N_5430,N_5543);
nor U5774 (N_5774,N_5442,N_5410);
or U5775 (N_5775,N_5451,N_5464);
nor U5776 (N_5776,N_5519,N_5516);
and U5777 (N_5777,N_5565,N_5413);
nor U5778 (N_5778,N_5556,N_5478);
nand U5779 (N_5779,N_5527,N_5522);
and U5780 (N_5780,N_5477,N_5511);
or U5781 (N_5781,N_5493,N_5567);
or U5782 (N_5782,N_5516,N_5581);
and U5783 (N_5783,N_5568,N_5534);
nand U5784 (N_5784,N_5534,N_5424);
or U5785 (N_5785,N_5427,N_5454);
nand U5786 (N_5786,N_5525,N_5420);
xnor U5787 (N_5787,N_5552,N_5525);
nand U5788 (N_5788,N_5563,N_5504);
nor U5789 (N_5789,N_5574,N_5485);
and U5790 (N_5790,N_5544,N_5502);
nor U5791 (N_5791,N_5452,N_5568);
and U5792 (N_5792,N_5411,N_5557);
nand U5793 (N_5793,N_5510,N_5432);
nor U5794 (N_5794,N_5492,N_5572);
nand U5795 (N_5795,N_5556,N_5574);
or U5796 (N_5796,N_5503,N_5594);
nand U5797 (N_5797,N_5521,N_5443);
and U5798 (N_5798,N_5533,N_5552);
or U5799 (N_5799,N_5540,N_5442);
nand U5800 (N_5800,N_5708,N_5648);
nand U5801 (N_5801,N_5659,N_5600);
or U5802 (N_5802,N_5639,N_5742);
nor U5803 (N_5803,N_5628,N_5612);
and U5804 (N_5804,N_5795,N_5718);
and U5805 (N_5805,N_5661,N_5652);
nor U5806 (N_5806,N_5698,N_5691);
or U5807 (N_5807,N_5699,N_5697);
or U5808 (N_5808,N_5721,N_5704);
and U5809 (N_5809,N_5679,N_5650);
nand U5810 (N_5810,N_5616,N_5717);
nand U5811 (N_5811,N_5642,N_5644);
and U5812 (N_5812,N_5687,N_5752);
and U5813 (N_5813,N_5634,N_5711);
nand U5814 (N_5814,N_5636,N_5759);
nor U5815 (N_5815,N_5793,N_5774);
nand U5816 (N_5816,N_5707,N_5604);
nand U5817 (N_5817,N_5620,N_5790);
or U5818 (N_5818,N_5710,N_5619);
nor U5819 (N_5819,N_5608,N_5673);
nor U5820 (N_5820,N_5631,N_5734);
and U5821 (N_5821,N_5794,N_5702);
or U5822 (N_5822,N_5762,N_5743);
and U5823 (N_5823,N_5739,N_5658);
and U5824 (N_5824,N_5719,N_5725);
and U5825 (N_5825,N_5680,N_5667);
nand U5826 (N_5826,N_5764,N_5615);
nand U5827 (N_5827,N_5611,N_5748);
or U5828 (N_5828,N_5773,N_5741);
and U5829 (N_5829,N_5695,N_5617);
or U5830 (N_5830,N_5689,N_5723);
xnor U5831 (N_5831,N_5760,N_5668);
and U5832 (N_5832,N_5749,N_5675);
nand U5833 (N_5833,N_5692,N_5602);
and U5834 (N_5834,N_5745,N_5789);
xnor U5835 (N_5835,N_5685,N_5714);
nand U5836 (N_5836,N_5610,N_5732);
and U5837 (N_5837,N_5798,N_5603);
nor U5838 (N_5838,N_5766,N_5788);
or U5839 (N_5839,N_5783,N_5666);
or U5840 (N_5840,N_5606,N_5753);
nor U5841 (N_5841,N_5756,N_5646);
or U5842 (N_5842,N_5637,N_5633);
and U5843 (N_5843,N_5657,N_5638);
nand U5844 (N_5844,N_5799,N_5792);
nand U5845 (N_5845,N_5765,N_5772);
nand U5846 (N_5846,N_5676,N_5700);
nor U5847 (N_5847,N_5640,N_5750);
or U5848 (N_5848,N_5733,N_5609);
nand U5849 (N_5849,N_5709,N_5769);
or U5850 (N_5850,N_5715,N_5728);
or U5851 (N_5851,N_5746,N_5713);
nor U5852 (N_5852,N_5730,N_5607);
and U5853 (N_5853,N_5625,N_5643);
xnor U5854 (N_5854,N_5731,N_5621);
or U5855 (N_5855,N_5786,N_5776);
nor U5856 (N_5856,N_5779,N_5662);
or U5857 (N_5857,N_5672,N_5651);
or U5858 (N_5858,N_5744,N_5647);
and U5859 (N_5859,N_5797,N_5684);
nand U5860 (N_5860,N_5751,N_5635);
and U5861 (N_5861,N_5771,N_5665);
nor U5862 (N_5862,N_5706,N_5624);
and U5863 (N_5863,N_5686,N_5670);
or U5864 (N_5864,N_5682,N_5683);
nor U5865 (N_5865,N_5664,N_5701);
or U5866 (N_5866,N_5653,N_5694);
or U5867 (N_5867,N_5618,N_5770);
nor U5868 (N_5868,N_5735,N_5712);
nand U5869 (N_5869,N_5720,N_5740);
or U5870 (N_5870,N_5654,N_5663);
and U5871 (N_5871,N_5768,N_5784);
or U5872 (N_5872,N_5613,N_5645);
or U5873 (N_5873,N_5722,N_5641);
nand U5874 (N_5874,N_5605,N_5655);
or U5875 (N_5875,N_5778,N_5690);
nand U5876 (N_5876,N_5796,N_5622);
and U5877 (N_5877,N_5787,N_5660);
nand U5878 (N_5878,N_5671,N_5780);
nor U5879 (N_5879,N_5649,N_5629);
nand U5880 (N_5880,N_5705,N_5761);
nand U5881 (N_5881,N_5677,N_5696);
nor U5882 (N_5882,N_5757,N_5703);
nor U5883 (N_5883,N_5777,N_5781);
and U5884 (N_5884,N_5747,N_5791);
nor U5885 (N_5885,N_5736,N_5681);
nor U5886 (N_5886,N_5688,N_5754);
nand U5887 (N_5887,N_5623,N_5716);
nand U5888 (N_5888,N_5678,N_5626);
or U5889 (N_5889,N_5767,N_5726);
and U5890 (N_5890,N_5724,N_5601);
or U5891 (N_5891,N_5785,N_5627);
and U5892 (N_5892,N_5674,N_5630);
or U5893 (N_5893,N_5727,N_5729);
nor U5894 (N_5894,N_5758,N_5669);
and U5895 (N_5895,N_5782,N_5693);
nor U5896 (N_5896,N_5632,N_5738);
nand U5897 (N_5897,N_5737,N_5755);
and U5898 (N_5898,N_5656,N_5763);
nand U5899 (N_5899,N_5775,N_5614);
and U5900 (N_5900,N_5613,N_5790);
or U5901 (N_5901,N_5652,N_5605);
nor U5902 (N_5902,N_5732,N_5723);
nor U5903 (N_5903,N_5660,N_5704);
nand U5904 (N_5904,N_5610,N_5600);
and U5905 (N_5905,N_5629,N_5642);
nand U5906 (N_5906,N_5649,N_5656);
nand U5907 (N_5907,N_5637,N_5789);
and U5908 (N_5908,N_5784,N_5625);
nand U5909 (N_5909,N_5775,N_5609);
nor U5910 (N_5910,N_5699,N_5689);
and U5911 (N_5911,N_5612,N_5734);
or U5912 (N_5912,N_5797,N_5658);
or U5913 (N_5913,N_5625,N_5616);
nand U5914 (N_5914,N_5742,N_5673);
nand U5915 (N_5915,N_5659,N_5692);
or U5916 (N_5916,N_5732,N_5611);
nand U5917 (N_5917,N_5785,N_5692);
or U5918 (N_5918,N_5605,N_5694);
nand U5919 (N_5919,N_5787,N_5711);
and U5920 (N_5920,N_5708,N_5684);
and U5921 (N_5921,N_5706,N_5781);
xnor U5922 (N_5922,N_5696,N_5730);
or U5923 (N_5923,N_5644,N_5699);
nor U5924 (N_5924,N_5791,N_5671);
and U5925 (N_5925,N_5696,N_5687);
and U5926 (N_5926,N_5743,N_5731);
nand U5927 (N_5927,N_5721,N_5638);
nand U5928 (N_5928,N_5758,N_5637);
or U5929 (N_5929,N_5708,N_5614);
and U5930 (N_5930,N_5793,N_5735);
nand U5931 (N_5931,N_5688,N_5702);
or U5932 (N_5932,N_5718,N_5661);
or U5933 (N_5933,N_5758,N_5615);
nor U5934 (N_5934,N_5773,N_5614);
or U5935 (N_5935,N_5664,N_5728);
or U5936 (N_5936,N_5705,N_5758);
nand U5937 (N_5937,N_5700,N_5784);
and U5938 (N_5938,N_5774,N_5771);
or U5939 (N_5939,N_5603,N_5734);
and U5940 (N_5940,N_5696,N_5663);
nor U5941 (N_5941,N_5769,N_5745);
or U5942 (N_5942,N_5698,N_5747);
xor U5943 (N_5943,N_5733,N_5771);
nand U5944 (N_5944,N_5649,N_5721);
nor U5945 (N_5945,N_5760,N_5737);
and U5946 (N_5946,N_5701,N_5614);
nand U5947 (N_5947,N_5768,N_5696);
or U5948 (N_5948,N_5657,N_5673);
and U5949 (N_5949,N_5601,N_5707);
nand U5950 (N_5950,N_5689,N_5614);
or U5951 (N_5951,N_5726,N_5700);
nand U5952 (N_5952,N_5600,N_5728);
or U5953 (N_5953,N_5758,N_5775);
or U5954 (N_5954,N_5753,N_5614);
or U5955 (N_5955,N_5759,N_5647);
nand U5956 (N_5956,N_5601,N_5607);
nand U5957 (N_5957,N_5773,N_5665);
or U5958 (N_5958,N_5621,N_5641);
and U5959 (N_5959,N_5630,N_5738);
nor U5960 (N_5960,N_5683,N_5751);
and U5961 (N_5961,N_5692,N_5675);
nor U5962 (N_5962,N_5784,N_5750);
or U5963 (N_5963,N_5736,N_5684);
nand U5964 (N_5964,N_5707,N_5652);
nor U5965 (N_5965,N_5767,N_5657);
nand U5966 (N_5966,N_5790,N_5665);
nor U5967 (N_5967,N_5681,N_5620);
and U5968 (N_5968,N_5648,N_5662);
nand U5969 (N_5969,N_5775,N_5719);
or U5970 (N_5970,N_5725,N_5776);
or U5971 (N_5971,N_5674,N_5627);
or U5972 (N_5972,N_5686,N_5605);
nor U5973 (N_5973,N_5778,N_5610);
nor U5974 (N_5974,N_5607,N_5722);
nand U5975 (N_5975,N_5737,N_5744);
or U5976 (N_5976,N_5646,N_5731);
or U5977 (N_5977,N_5648,N_5786);
nand U5978 (N_5978,N_5686,N_5638);
and U5979 (N_5979,N_5683,N_5702);
nor U5980 (N_5980,N_5672,N_5668);
nor U5981 (N_5981,N_5750,N_5612);
or U5982 (N_5982,N_5611,N_5721);
and U5983 (N_5983,N_5659,N_5685);
nand U5984 (N_5984,N_5640,N_5654);
or U5985 (N_5985,N_5602,N_5744);
nor U5986 (N_5986,N_5704,N_5624);
or U5987 (N_5987,N_5615,N_5752);
nand U5988 (N_5988,N_5649,N_5641);
or U5989 (N_5989,N_5600,N_5651);
or U5990 (N_5990,N_5642,N_5640);
nor U5991 (N_5991,N_5657,N_5635);
or U5992 (N_5992,N_5614,N_5726);
and U5993 (N_5993,N_5741,N_5724);
nand U5994 (N_5994,N_5793,N_5755);
and U5995 (N_5995,N_5748,N_5743);
or U5996 (N_5996,N_5753,N_5689);
nor U5997 (N_5997,N_5761,N_5653);
and U5998 (N_5998,N_5625,N_5730);
or U5999 (N_5999,N_5664,N_5758);
nor U6000 (N_6000,N_5944,N_5983);
or U6001 (N_6001,N_5996,N_5964);
nor U6002 (N_6002,N_5999,N_5873);
xnor U6003 (N_6003,N_5853,N_5975);
or U6004 (N_6004,N_5997,N_5821);
and U6005 (N_6005,N_5800,N_5921);
and U6006 (N_6006,N_5813,N_5959);
or U6007 (N_6007,N_5859,N_5801);
and U6008 (N_6008,N_5877,N_5829);
nand U6009 (N_6009,N_5994,N_5846);
nor U6010 (N_6010,N_5989,N_5832);
nor U6011 (N_6011,N_5828,N_5909);
nand U6012 (N_6012,N_5984,N_5874);
nand U6013 (N_6013,N_5971,N_5955);
nand U6014 (N_6014,N_5865,N_5844);
nor U6015 (N_6015,N_5904,N_5917);
or U6016 (N_6016,N_5988,N_5812);
nand U6017 (N_6017,N_5835,N_5869);
nor U6018 (N_6018,N_5903,N_5913);
nor U6019 (N_6019,N_5926,N_5930);
nor U6020 (N_6020,N_5923,N_5876);
nor U6021 (N_6021,N_5942,N_5939);
nand U6022 (N_6022,N_5890,N_5976);
and U6023 (N_6023,N_5875,N_5855);
nand U6024 (N_6024,N_5900,N_5948);
nor U6025 (N_6025,N_5963,N_5852);
and U6026 (N_6026,N_5811,N_5820);
and U6027 (N_6027,N_5928,N_5891);
nand U6028 (N_6028,N_5974,N_5929);
nor U6029 (N_6029,N_5961,N_5927);
or U6030 (N_6030,N_5956,N_5945);
xor U6031 (N_6031,N_5907,N_5987);
nand U6032 (N_6032,N_5953,N_5985);
and U6033 (N_6033,N_5847,N_5836);
nor U6034 (N_6034,N_5868,N_5886);
nor U6035 (N_6035,N_5978,N_5951);
nand U6036 (N_6036,N_5823,N_5901);
nor U6037 (N_6037,N_5937,N_5915);
nand U6038 (N_6038,N_5882,N_5981);
nand U6039 (N_6039,N_5980,N_5833);
or U6040 (N_6040,N_5932,N_5841);
and U6041 (N_6041,N_5973,N_5962);
and U6042 (N_6042,N_5970,N_5965);
nand U6043 (N_6043,N_5908,N_5938);
nor U6044 (N_6044,N_5840,N_5850);
and U6045 (N_6045,N_5918,N_5831);
or U6046 (N_6046,N_5960,N_5816);
or U6047 (N_6047,N_5910,N_5922);
and U6048 (N_6048,N_5858,N_5920);
nand U6049 (N_6049,N_5954,N_5993);
nand U6050 (N_6050,N_5824,N_5940);
and U6051 (N_6051,N_5883,N_5884);
nand U6052 (N_6052,N_5856,N_5935);
or U6053 (N_6053,N_5992,N_5849);
or U6054 (N_6054,N_5854,N_5827);
and U6055 (N_6055,N_5815,N_5843);
nand U6056 (N_6056,N_5864,N_5845);
or U6057 (N_6057,N_5952,N_5969);
nor U6058 (N_6058,N_5897,N_5943);
nand U6059 (N_6059,N_5804,N_5894);
nor U6060 (N_6060,N_5861,N_5839);
and U6061 (N_6061,N_5879,N_5977);
nand U6062 (N_6062,N_5896,N_5991);
nor U6063 (N_6063,N_5880,N_5887);
nor U6064 (N_6064,N_5912,N_5979);
and U6065 (N_6065,N_5914,N_5802);
nor U6066 (N_6066,N_5822,N_5866);
nand U6067 (N_6067,N_5872,N_5924);
nor U6068 (N_6068,N_5867,N_5941);
and U6069 (N_6069,N_5911,N_5986);
or U6070 (N_6070,N_5817,N_5819);
nand U6071 (N_6071,N_5809,N_5826);
nand U6072 (N_6072,N_5947,N_5889);
and U6073 (N_6073,N_5878,N_5934);
and U6074 (N_6074,N_5807,N_5803);
or U6075 (N_6075,N_5881,N_5950);
or U6076 (N_6076,N_5967,N_5936);
and U6077 (N_6077,N_5830,N_5860);
nand U6078 (N_6078,N_5902,N_5946);
nor U6079 (N_6079,N_5933,N_5893);
or U6080 (N_6080,N_5808,N_5905);
or U6081 (N_6081,N_5895,N_5863);
or U6082 (N_6082,N_5919,N_5998);
nand U6083 (N_6083,N_5848,N_5958);
nor U6084 (N_6084,N_5931,N_5972);
or U6085 (N_6085,N_5857,N_5885);
nor U6086 (N_6086,N_5806,N_5837);
or U6087 (N_6087,N_5825,N_5906);
and U6088 (N_6088,N_5838,N_5898);
nor U6089 (N_6089,N_5949,N_5834);
nor U6090 (N_6090,N_5916,N_5870);
nand U6091 (N_6091,N_5966,N_5925);
or U6092 (N_6092,N_5810,N_5871);
nand U6093 (N_6093,N_5968,N_5842);
or U6094 (N_6094,N_5982,N_5899);
xnor U6095 (N_6095,N_5995,N_5990);
nand U6096 (N_6096,N_5892,N_5814);
and U6097 (N_6097,N_5957,N_5818);
and U6098 (N_6098,N_5851,N_5862);
nor U6099 (N_6099,N_5805,N_5888);
and U6100 (N_6100,N_5859,N_5986);
or U6101 (N_6101,N_5851,N_5839);
nand U6102 (N_6102,N_5930,N_5894);
and U6103 (N_6103,N_5914,N_5992);
and U6104 (N_6104,N_5908,N_5851);
or U6105 (N_6105,N_5914,N_5959);
nor U6106 (N_6106,N_5945,N_5998);
nand U6107 (N_6107,N_5871,N_5999);
or U6108 (N_6108,N_5889,N_5967);
or U6109 (N_6109,N_5872,N_5967);
or U6110 (N_6110,N_5890,N_5961);
nor U6111 (N_6111,N_5809,N_5856);
or U6112 (N_6112,N_5817,N_5832);
nand U6113 (N_6113,N_5912,N_5957);
and U6114 (N_6114,N_5820,N_5997);
or U6115 (N_6115,N_5842,N_5857);
nor U6116 (N_6116,N_5916,N_5915);
or U6117 (N_6117,N_5835,N_5966);
nand U6118 (N_6118,N_5939,N_5891);
nor U6119 (N_6119,N_5975,N_5984);
nand U6120 (N_6120,N_5896,N_5827);
nor U6121 (N_6121,N_5942,N_5871);
and U6122 (N_6122,N_5940,N_5836);
nor U6123 (N_6123,N_5839,N_5977);
or U6124 (N_6124,N_5992,N_5802);
or U6125 (N_6125,N_5922,N_5958);
and U6126 (N_6126,N_5920,N_5836);
nand U6127 (N_6127,N_5889,N_5982);
nand U6128 (N_6128,N_5829,N_5945);
and U6129 (N_6129,N_5964,N_5906);
nand U6130 (N_6130,N_5809,N_5878);
xnor U6131 (N_6131,N_5822,N_5856);
nand U6132 (N_6132,N_5845,N_5909);
and U6133 (N_6133,N_5895,N_5902);
nor U6134 (N_6134,N_5897,N_5902);
nor U6135 (N_6135,N_5999,N_5984);
nor U6136 (N_6136,N_5980,N_5916);
and U6137 (N_6137,N_5922,N_5997);
nor U6138 (N_6138,N_5960,N_5857);
or U6139 (N_6139,N_5962,N_5989);
or U6140 (N_6140,N_5848,N_5955);
nor U6141 (N_6141,N_5908,N_5895);
and U6142 (N_6142,N_5845,N_5986);
xor U6143 (N_6143,N_5857,N_5887);
nand U6144 (N_6144,N_5922,N_5890);
nand U6145 (N_6145,N_5957,N_5801);
nor U6146 (N_6146,N_5934,N_5984);
and U6147 (N_6147,N_5947,N_5836);
or U6148 (N_6148,N_5981,N_5969);
and U6149 (N_6149,N_5963,N_5971);
or U6150 (N_6150,N_5835,N_5870);
or U6151 (N_6151,N_5899,N_5855);
and U6152 (N_6152,N_5817,N_5954);
and U6153 (N_6153,N_5974,N_5822);
nor U6154 (N_6154,N_5891,N_5905);
nand U6155 (N_6155,N_5945,N_5920);
and U6156 (N_6156,N_5917,N_5856);
or U6157 (N_6157,N_5903,N_5907);
nand U6158 (N_6158,N_5849,N_5834);
and U6159 (N_6159,N_5847,N_5912);
nor U6160 (N_6160,N_5803,N_5877);
nand U6161 (N_6161,N_5999,N_5857);
and U6162 (N_6162,N_5949,N_5900);
nand U6163 (N_6163,N_5893,N_5815);
and U6164 (N_6164,N_5897,N_5817);
nand U6165 (N_6165,N_5973,N_5993);
or U6166 (N_6166,N_5941,N_5891);
or U6167 (N_6167,N_5851,N_5959);
nand U6168 (N_6168,N_5938,N_5976);
nand U6169 (N_6169,N_5975,N_5897);
and U6170 (N_6170,N_5943,N_5945);
and U6171 (N_6171,N_5970,N_5911);
or U6172 (N_6172,N_5974,N_5911);
nor U6173 (N_6173,N_5801,N_5987);
nor U6174 (N_6174,N_5935,N_5812);
and U6175 (N_6175,N_5878,N_5928);
or U6176 (N_6176,N_5926,N_5992);
nand U6177 (N_6177,N_5979,N_5908);
or U6178 (N_6178,N_5802,N_5866);
xnor U6179 (N_6179,N_5874,N_5980);
nand U6180 (N_6180,N_5916,N_5812);
and U6181 (N_6181,N_5923,N_5900);
and U6182 (N_6182,N_5833,N_5906);
xor U6183 (N_6183,N_5802,N_5969);
nand U6184 (N_6184,N_5961,N_5985);
nand U6185 (N_6185,N_5918,N_5965);
and U6186 (N_6186,N_5895,N_5937);
nor U6187 (N_6187,N_5811,N_5844);
and U6188 (N_6188,N_5958,N_5992);
or U6189 (N_6189,N_5830,N_5926);
or U6190 (N_6190,N_5888,N_5868);
and U6191 (N_6191,N_5865,N_5882);
and U6192 (N_6192,N_5895,N_5995);
nor U6193 (N_6193,N_5829,N_5895);
nor U6194 (N_6194,N_5828,N_5918);
and U6195 (N_6195,N_5985,N_5921);
nand U6196 (N_6196,N_5882,N_5923);
and U6197 (N_6197,N_5862,N_5838);
nor U6198 (N_6198,N_5942,N_5829);
or U6199 (N_6199,N_5981,N_5873);
nor U6200 (N_6200,N_6182,N_6001);
and U6201 (N_6201,N_6154,N_6124);
nor U6202 (N_6202,N_6050,N_6085);
nand U6203 (N_6203,N_6089,N_6105);
and U6204 (N_6204,N_6044,N_6103);
nand U6205 (N_6205,N_6034,N_6101);
nand U6206 (N_6206,N_6068,N_6125);
and U6207 (N_6207,N_6057,N_6082);
and U6208 (N_6208,N_6111,N_6183);
nand U6209 (N_6209,N_6168,N_6115);
nor U6210 (N_6210,N_6065,N_6176);
xnor U6211 (N_6211,N_6175,N_6131);
or U6212 (N_6212,N_6196,N_6126);
or U6213 (N_6213,N_6099,N_6002);
and U6214 (N_6214,N_6136,N_6010);
nor U6215 (N_6215,N_6157,N_6108);
and U6216 (N_6216,N_6166,N_6112);
or U6217 (N_6217,N_6162,N_6056);
and U6218 (N_6218,N_6193,N_6097);
and U6219 (N_6219,N_6077,N_6106);
nand U6220 (N_6220,N_6164,N_6022);
nand U6221 (N_6221,N_6011,N_6070);
nand U6222 (N_6222,N_6110,N_6086);
xnor U6223 (N_6223,N_6170,N_6051);
nand U6224 (N_6224,N_6169,N_6003);
nor U6225 (N_6225,N_6081,N_6100);
nand U6226 (N_6226,N_6198,N_6141);
nand U6227 (N_6227,N_6120,N_6040);
and U6228 (N_6228,N_6107,N_6046);
and U6229 (N_6229,N_6018,N_6083);
nand U6230 (N_6230,N_6015,N_6054);
xor U6231 (N_6231,N_6167,N_6029);
nor U6232 (N_6232,N_6045,N_6043);
or U6233 (N_6233,N_6074,N_6178);
nor U6234 (N_6234,N_6037,N_6071);
nand U6235 (N_6235,N_6041,N_6104);
and U6236 (N_6236,N_6118,N_6152);
and U6237 (N_6237,N_6060,N_6028);
nor U6238 (N_6238,N_6165,N_6181);
and U6239 (N_6239,N_6121,N_6146);
or U6240 (N_6240,N_6113,N_6163);
nor U6241 (N_6241,N_6032,N_6147);
or U6242 (N_6242,N_6109,N_6135);
and U6243 (N_6243,N_6139,N_6186);
nor U6244 (N_6244,N_6004,N_6021);
and U6245 (N_6245,N_6066,N_6067);
or U6246 (N_6246,N_6160,N_6013);
or U6247 (N_6247,N_6150,N_6014);
or U6248 (N_6248,N_6171,N_6038);
nand U6249 (N_6249,N_6127,N_6130);
or U6250 (N_6250,N_6094,N_6187);
nand U6251 (N_6251,N_6129,N_6161);
xor U6252 (N_6252,N_6078,N_6143);
nor U6253 (N_6253,N_6008,N_6095);
nand U6254 (N_6254,N_6027,N_6059);
nand U6255 (N_6255,N_6180,N_6090);
nor U6256 (N_6256,N_6184,N_6075);
and U6257 (N_6257,N_6158,N_6092);
nand U6258 (N_6258,N_6138,N_6000);
nand U6259 (N_6259,N_6128,N_6006);
and U6260 (N_6260,N_6192,N_6199);
nor U6261 (N_6261,N_6102,N_6123);
or U6262 (N_6262,N_6019,N_6079);
and U6263 (N_6263,N_6088,N_6191);
nor U6264 (N_6264,N_6172,N_6073);
or U6265 (N_6265,N_6185,N_6119);
and U6266 (N_6266,N_6096,N_6132);
or U6267 (N_6267,N_6047,N_6133);
and U6268 (N_6268,N_6093,N_6144);
nor U6269 (N_6269,N_6061,N_6025);
or U6270 (N_6270,N_6055,N_6179);
or U6271 (N_6271,N_6155,N_6145);
or U6272 (N_6272,N_6030,N_6149);
nand U6273 (N_6273,N_6194,N_6053);
nand U6274 (N_6274,N_6049,N_6173);
xor U6275 (N_6275,N_6159,N_6042);
and U6276 (N_6276,N_6035,N_6023);
nand U6277 (N_6277,N_6005,N_6137);
nand U6278 (N_6278,N_6062,N_6190);
nor U6279 (N_6279,N_6069,N_6052);
nand U6280 (N_6280,N_6177,N_6072);
and U6281 (N_6281,N_6048,N_6148);
nor U6282 (N_6282,N_6012,N_6026);
nor U6283 (N_6283,N_6117,N_6020);
or U6284 (N_6284,N_6017,N_6116);
nor U6285 (N_6285,N_6114,N_6091);
nand U6286 (N_6286,N_6156,N_6122);
or U6287 (N_6287,N_6007,N_6142);
nand U6288 (N_6288,N_6016,N_6063);
or U6289 (N_6289,N_6058,N_6033);
and U6290 (N_6290,N_6080,N_6009);
or U6291 (N_6291,N_6064,N_6195);
nor U6292 (N_6292,N_6087,N_6153);
or U6293 (N_6293,N_6024,N_6134);
nor U6294 (N_6294,N_6084,N_6189);
and U6295 (N_6295,N_6076,N_6036);
nand U6296 (N_6296,N_6151,N_6174);
nor U6297 (N_6297,N_6039,N_6197);
and U6298 (N_6298,N_6098,N_6140);
and U6299 (N_6299,N_6188,N_6031);
and U6300 (N_6300,N_6118,N_6122);
nor U6301 (N_6301,N_6017,N_6029);
nand U6302 (N_6302,N_6073,N_6092);
nand U6303 (N_6303,N_6098,N_6122);
nor U6304 (N_6304,N_6111,N_6118);
or U6305 (N_6305,N_6017,N_6151);
and U6306 (N_6306,N_6067,N_6012);
nor U6307 (N_6307,N_6143,N_6100);
and U6308 (N_6308,N_6165,N_6131);
or U6309 (N_6309,N_6000,N_6139);
or U6310 (N_6310,N_6046,N_6134);
and U6311 (N_6311,N_6149,N_6114);
nand U6312 (N_6312,N_6000,N_6036);
nand U6313 (N_6313,N_6035,N_6128);
nor U6314 (N_6314,N_6127,N_6143);
and U6315 (N_6315,N_6019,N_6072);
nor U6316 (N_6316,N_6130,N_6166);
nor U6317 (N_6317,N_6014,N_6042);
nand U6318 (N_6318,N_6056,N_6087);
and U6319 (N_6319,N_6075,N_6181);
nand U6320 (N_6320,N_6077,N_6167);
or U6321 (N_6321,N_6042,N_6104);
and U6322 (N_6322,N_6063,N_6041);
or U6323 (N_6323,N_6028,N_6065);
nand U6324 (N_6324,N_6145,N_6162);
xor U6325 (N_6325,N_6058,N_6141);
and U6326 (N_6326,N_6015,N_6053);
nand U6327 (N_6327,N_6176,N_6100);
nand U6328 (N_6328,N_6136,N_6195);
or U6329 (N_6329,N_6088,N_6017);
nor U6330 (N_6330,N_6080,N_6109);
nor U6331 (N_6331,N_6162,N_6097);
or U6332 (N_6332,N_6119,N_6035);
nand U6333 (N_6333,N_6197,N_6173);
nand U6334 (N_6334,N_6049,N_6034);
nor U6335 (N_6335,N_6181,N_6188);
nand U6336 (N_6336,N_6080,N_6167);
and U6337 (N_6337,N_6122,N_6094);
nand U6338 (N_6338,N_6198,N_6087);
and U6339 (N_6339,N_6027,N_6037);
nand U6340 (N_6340,N_6123,N_6117);
nand U6341 (N_6341,N_6015,N_6137);
and U6342 (N_6342,N_6169,N_6008);
nand U6343 (N_6343,N_6043,N_6067);
and U6344 (N_6344,N_6042,N_6062);
and U6345 (N_6345,N_6050,N_6036);
nand U6346 (N_6346,N_6173,N_6030);
or U6347 (N_6347,N_6151,N_6012);
nor U6348 (N_6348,N_6035,N_6022);
nand U6349 (N_6349,N_6033,N_6049);
nor U6350 (N_6350,N_6003,N_6155);
or U6351 (N_6351,N_6103,N_6118);
and U6352 (N_6352,N_6125,N_6051);
and U6353 (N_6353,N_6103,N_6017);
xnor U6354 (N_6354,N_6106,N_6178);
and U6355 (N_6355,N_6113,N_6139);
and U6356 (N_6356,N_6105,N_6020);
or U6357 (N_6357,N_6151,N_6083);
nor U6358 (N_6358,N_6079,N_6000);
nor U6359 (N_6359,N_6077,N_6097);
or U6360 (N_6360,N_6198,N_6093);
nand U6361 (N_6361,N_6083,N_6015);
and U6362 (N_6362,N_6196,N_6078);
nor U6363 (N_6363,N_6127,N_6181);
nand U6364 (N_6364,N_6066,N_6167);
and U6365 (N_6365,N_6033,N_6012);
nand U6366 (N_6366,N_6095,N_6157);
nand U6367 (N_6367,N_6120,N_6131);
or U6368 (N_6368,N_6031,N_6077);
nand U6369 (N_6369,N_6051,N_6076);
and U6370 (N_6370,N_6038,N_6100);
nor U6371 (N_6371,N_6122,N_6007);
nor U6372 (N_6372,N_6114,N_6165);
nor U6373 (N_6373,N_6073,N_6090);
nand U6374 (N_6374,N_6048,N_6045);
or U6375 (N_6375,N_6030,N_6032);
nand U6376 (N_6376,N_6098,N_6107);
nand U6377 (N_6377,N_6172,N_6060);
and U6378 (N_6378,N_6126,N_6122);
nand U6379 (N_6379,N_6147,N_6062);
nand U6380 (N_6380,N_6015,N_6045);
and U6381 (N_6381,N_6184,N_6019);
and U6382 (N_6382,N_6026,N_6093);
and U6383 (N_6383,N_6077,N_6137);
and U6384 (N_6384,N_6026,N_6108);
nor U6385 (N_6385,N_6114,N_6030);
or U6386 (N_6386,N_6117,N_6053);
nand U6387 (N_6387,N_6064,N_6105);
and U6388 (N_6388,N_6052,N_6182);
nor U6389 (N_6389,N_6104,N_6063);
nand U6390 (N_6390,N_6037,N_6012);
or U6391 (N_6391,N_6145,N_6134);
or U6392 (N_6392,N_6001,N_6012);
and U6393 (N_6393,N_6026,N_6172);
nand U6394 (N_6394,N_6107,N_6125);
nor U6395 (N_6395,N_6066,N_6053);
nor U6396 (N_6396,N_6123,N_6099);
or U6397 (N_6397,N_6050,N_6004);
nand U6398 (N_6398,N_6181,N_6105);
or U6399 (N_6399,N_6173,N_6014);
nand U6400 (N_6400,N_6228,N_6373);
nor U6401 (N_6401,N_6287,N_6246);
xor U6402 (N_6402,N_6240,N_6219);
or U6403 (N_6403,N_6285,N_6381);
nand U6404 (N_6404,N_6380,N_6366);
or U6405 (N_6405,N_6351,N_6320);
and U6406 (N_6406,N_6398,N_6203);
nor U6407 (N_6407,N_6204,N_6334);
or U6408 (N_6408,N_6368,N_6249);
and U6409 (N_6409,N_6394,N_6215);
nor U6410 (N_6410,N_6376,N_6393);
nor U6411 (N_6411,N_6254,N_6382);
and U6412 (N_6412,N_6278,N_6311);
or U6413 (N_6413,N_6325,N_6205);
or U6414 (N_6414,N_6377,N_6383);
and U6415 (N_6415,N_6353,N_6250);
nor U6416 (N_6416,N_6297,N_6346);
and U6417 (N_6417,N_6315,N_6293);
and U6418 (N_6418,N_6303,N_6288);
nor U6419 (N_6419,N_6358,N_6357);
and U6420 (N_6420,N_6255,N_6302);
and U6421 (N_6421,N_6369,N_6291);
and U6422 (N_6422,N_6345,N_6280);
or U6423 (N_6423,N_6391,N_6387);
or U6424 (N_6424,N_6284,N_6209);
nor U6425 (N_6425,N_6313,N_6226);
nand U6426 (N_6426,N_6257,N_6251);
nor U6427 (N_6427,N_6333,N_6201);
or U6428 (N_6428,N_6244,N_6227);
nor U6429 (N_6429,N_6367,N_6339);
nand U6430 (N_6430,N_6350,N_6340);
nor U6431 (N_6431,N_6232,N_6332);
and U6432 (N_6432,N_6370,N_6281);
nor U6433 (N_6433,N_6309,N_6225);
nand U6434 (N_6434,N_6307,N_6295);
and U6435 (N_6435,N_6263,N_6396);
nand U6436 (N_6436,N_6348,N_6214);
nor U6437 (N_6437,N_6261,N_6319);
or U6438 (N_6438,N_6399,N_6359);
nor U6439 (N_6439,N_6323,N_6304);
or U6440 (N_6440,N_6222,N_6270);
and U6441 (N_6441,N_6327,N_6384);
nand U6442 (N_6442,N_6231,N_6264);
nand U6443 (N_6443,N_6216,N_6212);
or U6444 (N_6444,N_6397,N_6324);
and U6445 (N_6445,N_6385,N_6312);
and U6446 (N_6446,N_6349,N_6317);
or U6447 (N_6447,N_6289,N_6355);
or U6448 (N_6448,N_6272,N_6268);
or U6449 (N_6449,N_6229,N_6364);
nand U6450 (N_6450,N_6259,N_6378);
xnor U6451 (N_6451,N_6375,N_6300);
xnor U6452 (N_6452,N_6245,N_6274);
xor U6453 (N_6453,N_6276,N_6301);
and U6454 (N_6454,N_6386,N_6218);
or U6455 (N_6455,N_6310,N_6234);
and U6456 (N_6456,N_6262,N_6354);
nor U6457 (N_6457,N_6267,N_6256);
nor U6458 (N_6458,N_6336,N_6316);
and U6459 (N_6459,N_6248,N_6388);
or U6460 (N_6460,N_6286,N_6236);
and U6461 (N_6461,N_6243,N_6260);
nand U6462 (N_6462,N_6352,N_6202);
nand U6463 (N_6463,N_6330,N_6223);
or U6464 (N_6464,N_6269,N_6211);
or U6465 (N_6465,N_6224,N_6242);
nand U6466 (N_6466,N_6230,N_6241);
and U6467 (N_6467,N_6338,N_6342);
xor U6468 (N_6468,N_6344,N_6273);
nor U6469 (N_6469,N_6258,N_6329);
or U6470 (N_6470,N_6271,N_6322);
nor U6471 (N_6471,N_6347,N_6362);
nor U6472 (N_6472,N_6206,N_6335);
nor U6473 (N_6473,N_6207,N_6379);
nor U6474 (N_6474,N_6296,N_6314);
and U6475 (N_6475,N_6363,N_6252);
xor U6476 (N_6476,N_6371,N_6360);
nor U6477 (N_6477,N_6372,N_6290);
nor U6478 (N_6478,N_6210,N_6208);
nor U6479 (N_6479,N_6321,N_6283);
or U6480 (N_6480,N_6239,N_6305);
and U6481 (N_6481,N_6299,N_6356);
nor U6482 (N_6482,N_6266,N_6265);
or U6483 (N_6483,N_6292,N_6337);
and U6484 (N_6484,N_6217,N_6200);
xnor U6485 (N_6485,N_6361,N_6253);
or U6486 (N_6486,N_6294,N_6306);
xor U6487 (N_6487,N_6213,N_6275);
nand U6488 (N_6488,N_6237,N_6343);
nand U6489 (N_6489,N_6374,N_6235);
and U6490 (N_6490,N_6395,N_6331);
nand U6491 (N_6491,N_6279,N_6298);
or U6492 (N_6492,N_6365,N_6220);
and U6493 (N_6493,N_6328,N_6390);
and U6494 (N_6494,N_6341,N_6277);
and U6495 (N_6495,N_6221,N_6389);
nor U6496 (N_6496,N_6233,N_6318);
or U6497 (N_6497,N_6238,N_6392);
and U6498 (N_6498,N_6247,N_6282);
and U6499 (N_6499,N_6326,N_6308);
or U6500 (N_6500,N_6237,N_6250);
or U6501 (N_6501,N_6293,N_6276);
or U6502 (N_6502,N_6390,N_6200);
or U6503 (N_6503,N_6292,N_6253);
or U6504 (N_6504,N_6266,N_6330);
nand U6505 (N_6505,N_6329,N_6364);
and U6506 (N_6506,N_6314,N_6334);
or U6507 (N_6507,N_6256,N_6280);
nor U6508 (N_6508,N_6259,N_6258);
or U6509 (N_6509,N_6209,N_6238);
nand U6510 (N_6510,N_6223,N_6349);
or U6511 (N_6511,N_6373,N_6307);
or U6512 (N_6512,N_6368,N_6209);
and U6513 (N_6513,N_6330,N_6369);
and U6514 (N_6514,N_6296,N_6249);
or U6515 (N_6515,N_6271,N_6247);
and U6516 (N_6516,N_6259,N_6310);
nand U6517 (N_6517,N_6277,N_6371);
nand U6518 (N_6518,N_6386,N_6388);
or U6519 (N_6519,N_6342,N_6335);
nand U6520 (N_6520,N_6209,N_6212);
nand U6521 (N_6521,N_6200,N_6307);
nor U6522 (N_6522,N_6371,N_6298);
nand U6523 (N_6523,N_6226,N_6360);
nor U6524 (N_6524,N_6301,N_6310);
and U6525 (N_6525,N_6217,N_6308);
nand U6526 (N_6526,N_6336,N_6326);
and U6527 (N_6527,N_6383,N_6211);
nor U6528 (N_6528,N_6361,N_6254);
nor U6529 (N_6529,N_6234,N_6312);
nand U6530 (N_6530,N_6399,N_6286);
nand U6531 (N_6531,N_6286,N_6239);
nor U6532 (N_6532,N_6367,N_6290);
nor U6533 (N_6533,N_6270,N_6371);
and U6534 (N_6534,N_6318,N_6211);
nand U6535 (N_6535,N_6285,N_6276);
nand U6536 (N_6536,N_6374,N_6324);
xor U6537 (N_6537,N_6273,N_6258);
nand U6538 (N_6538,N_6343,N_6270);
and U6539 (N_6539,N_6337,N_6250);
or U6540 (N_6540,N_6233,N_6266);
and U6541 (N_6541,N_6297,N_6224);
nor U6542 (N_6542,N_6362,N_6297);
or U6543 (N_6543,N_6205,N_6220);
nand U6544 (N_6544,N_6244,N_6328);
nand U6545 (N_6545,N_6347,N_6343);
nor U6546 (N_6546,N_6264,N_6216);
or U6547 (N_6547,N_6339,N_6307);
and U6548 (N_6548,N_6222,N_6398);
nor U6549 (N_6549,N_6215,N_6227);
nor U6550 (N_6550,N_6353,N_6375);
and U6551 (N_6551,N_6321,N_6353);
nand U6552 (N_6552,N_6350,N_6240);
and U6553 (N_6553,N_6221,N_6360);
and U6554 (N_6554,N_6276,N_6286);
and U6555 (N_6555,N_6395,N_6339);
nand U6556 (N_6556,N_6271,N_6339);
or U6557 (N_6557,N_6251,N_6350);
nand U6558 (N_6558,N_6237,N_6359);
and U6559 (N_6559,N_6381,N_6271);
or U6560 (N_6560,N_6383,N_6316);
or U6561 (N_6561,N_6323,N_6238);
nand U6562 (N_6562,N_6329,N_6390);
or U6563 (N_6563,N_6258,N_6257);
or U6564 (N_6564,N_6296,N_6209);
and U6565 (N_6565,N_6338,N_6201);
nor U6566 (N_6566,N_6271,N_6396);
nor U6567 (N_6567,N_6231,N_6308);
nand U6568 (N_6568,N_6219,N_6281);
nand U6569 (N_6569,N_6235,N_6341);
nor U6570 (N_6570,N_6312,N_6356);
or U6571 (N_6571,N_6243,N_6383);
or U6572 (N_6572,N_6337,N_6236);
nand U6573 (N_6573,N_6382,N_6323);
xor U6574 (N_6574,N_6239,N_6292);
and U6575 (N_6575,N_6247,N_6366);
nor U6576 (N_6576,N_6300,N_6327);
and U6577 (N_6577,N_6347,N_6385);
and U6578 (N_6578,N_6263,N_6266);
nor U6579 (N_6579,N_6292,N_6364);
nand U6580 (N_6580,N_6210,N_6343);
nor U6581 (N_6581,N_6363,N_6357);
nor U6582 (N_6582,N_6306,N_6241);
and U6583 (N_6583,N_6352,N_6237);
nand U6584 (N_6584,N_6323,N_6273);
and U6585 (N_6585,N_6392,N_6374);
nand U6586 (N_6586,N_6203,N_6369);
nor U6587 (N_6587,N_6218,N_6371);
or U6588 (N_6588,N_6249,N_6366);
nor U6589 (N_6589,N_6295,N_6340);
or U6590 (N_6590,N_6349,N_6364);
or U6591 (N_6591,N_6215,N_6360);
or U6592 (N_6592,N_6312,N_6382);
and U6593 (N_6593,N_6223,N_6291);
nand U6594 (N_6594,N_6225,N_6371);
nand U6595 (N_6595,N_6398,N_6385);
or U6596 (N_6596,N_6366,N_6332);
nor U6597 (N_6597,N_6347,N_6211);
or U6598 (N_6598,N_6339,N_6393);
nor U6599 (N_6599,N_6335,N_6332);
or U6600 (N_6600,N_6519,N_6508);
and U6601 (N_6601,N_6461,N_6413);
nand U6602 (N_6602,N_6419,N_6432);
nor U6603 (N_6603,N_6502,N_6516);
or U6604 (N_6604,N_6415,N_6459);
xnor U6605 (N_6605,N_6423,N_6538);
nor U6606 (N_6606,N_6581,N_6456);
or U6607 (N_6607,N_6414,N_6515);
nand U6608 (N_6608,N_6514,N_6547);
nand U6609 (N_6609,N_6557,N_6481);
or U6610 (N_6610,N_6537,N_6549);
and U6611 (N_6611,N_6500,N_6512);
nor U6612 (N_6612,N_6572,N_6412);
nor U6613 (N_6613,N_6401,N_6532);
and U6614 (N_6614,N_6442,N_6513);
and U6615 (N_6615,N_6529,N_6584);
nand U6616 (N_6616,N_6530,N_6510);
or U6617 (N_6617,N_6465,N_6463);
nor U6618 (N_6618,N_6410,N_6409);
or U6619 (N_6619,N_6476,N_6418);
and U6620 (N_6620,N_6539,N_6569);
nand U6621 (N_6621,N_6488,N_6478);
or U6622 (N_6622,N_6427,N_6585);
and U6623 (N_6623,N_6449,N_6499);
nand U6624 (N_6624,N_6404,N_6573);
nand U6625 (N_6625,N_6441,N_6430);
nand U6626 (N_6626,N_6565,N_6533);
and U6627 (N_6627,N_6424,N_6405);
nand U6628 (N_6628,N_6436,N_6588);
or U6629 (N_6629,N_6462,N_6440);
nor U6630 (N_6630,N_6560,N_6439);
nand U6631 (N_6631,N_6551,N_6496);
nor U6632 (N_6632,N_6451,N_6559);
nor U6633 (N_6633,N_6417,N_6596);
nor U6634 (N_6634,N_6503,N_6536);
and U6635 (N_6635,N_6567,N_6593);
nor U6636 (N_6636,N_6470,N_6595);
or U6637 (N_6637,N_6580,N_6523);
or U6638 (N_6638,N_6446,N_6426);
nand U6639 (N_6639,N_6583,N_6467);
xor U6640 (N_6640,N_6437,N_6468);
or U6641 (N_6641,N_6522,N_6590);
nor U6642 (N_6642,N_6403,N_6587);
and U6643 (N_6643,N_6431,N_6526);
nand U6644 (N_6644,N_6542,N_6576);
and U6645 (N_6645,N_6540,N_6472);
or U6646 (N_6646,N_6517,N_6420);
nor U6647 (N_6647,N_6509,N_6479);
nand U6648 (N_6648,N_6591,N_6524);
nand U6649 (N_6649,N_6599,N_6407);
nand U6650 (N_6650,N_6555,N_6422);
or U6651 (N_6651,N_6425,N_6448);
nand U6652 (N_6652,N_6582,N_6571);
or U6653 (N_6653,N_6561,N_6406);
nor U6654 (N_6654,N_6553,N_6505);
or U6655 (N_6655,N_6563,N_6518);
nand U6656 (N_6656,N_6433,N_6445);
nand U6657 (N_6657,N_6589,N_6554);
xnor U6658 (N_6658,N_6545,N_6491);
nand U6659 (N_6659,N_6464,N_6469);
xor U6660 (N_6660,N_6490,N_6501);
nand U6661 (N_6661,N_6527,N_6552);
and U6662 (N_6662,N_6562,N_6434);
or U6663 (N_6663,N_6568,N_6447);
nand U6664 (N_6664,N_6507,N_6458);
nand U6665 (N_6665,N_6429,N_6497);
nand U6666 (N_6666,N_6483,N_6550);
nand U6667 (N_6667,N_6457,N_6485);
nand U6668 (N_6668,N_6486,N_6471);
nor U6669 (N_6669,N_6475,N_6574);
or U6670 (N_6670,N_6450,N_6438);
xor U6671 (N_6671,N_6428,N_6493);
or U6672 (N_6672,N_6531,N_6477);
nor U6673 (N_6673,N_6487,N_6544);
nand U6674 (N_6674,N_6535,N_6577);
nor U6675 (N_6675,N_6594,N_6598);
nor U6676 (N_6676,N_6400,N_6578);
and U6677 (N_6677,N_6482,N_6511);
and U6678 (N_6678,N_6474,N_6528);
or U6679 (N_6679,N_6579,N_6494);
nand U6680 (N_6680,N_6454,N_6564);
nand U6681 (N_6681,N_6570,N_6546);
or U6682 (N_6682,N_6506,N_6444);
nor U6683 (N_6683,N_6435,N_6408);
nor U6684 (N_6684,N_6575,N_6489);
xor U6685 (N_6685,N_6520,N_6492);
nand U6686 (N_6686,N_6484,N_6521);
or U6687 (N_6687,N_6473,N_6455);
nand U6688 (N_6688,N_6402,N_6421);
nor U6689 (N_6689,N_6460,N_6504);
nor U6690 (N_6690,N_6466,N_6543);
or U6691 (N_6691,N_6498,N_6452);
and U6692 (N_6692,N_6566,N_6597);
nand U6693 (N_6693,N_6416,N_6443);
nor U6694 (N_6694,N_6556,N_6534);
nand U6695 (N_6695,N_6586,N_6592);
or U6696 (N_6696,N_6525,N_6480);
nand U6697 (N_6697,N_6495,N_6411);
or U6698 (N_6698,N_6541,N_6548);
or U6699 (N_6699,N_6558,N_6453);
nor U6700 (N_6700,N_6491,N_6425);
nand U6701 (N_6701,N_6451,N_6417);
and U6702 (N_6702,N_6407,N_6476);
and U6703 (N_6703,N_6513,N_6405);
xnor U6704 (N_6704,N_6592,N_6578);
and U6705 (N_6705,N_6549,N_6419);
nand U6706 (N_6706,N_6466,N_6561);
or U6707 (N_6707,N_6572,N_6552);
nor U6708 (N_6708,N_6505,N_6525);
or U6709 (N_6709,N_6590,N_6409);
or U6710 (N_6710,N_6472,N_6587);
nand U6711 (N_6711,N_6580,N_6420);
or U6712 (N_6712,N_6512,N_6591);
nor U6713 (N_6713,N_6426,N_6598);
nor U6714 (N_6714,N_6535,N_6485);
nor U6715 (N_6715,N_6437,N_6481);
xnor U6716 (N_6716,N_6572,N_6569);
and U6717 (N_6717,N_6466,N_6579);
nor U6718 (N_6718,N_6501,N_6561);
or U6719 (N_6719,N_6505,N_6581);
nor U6720 (N_6720,N_6581,N_6508);
nor U6721 (N_6721,N_6431,N_6494);
nand U6722 (N_6722,N_6521,N_6494);
nand U6723 (N_6723,N_6518,N_6595);
nor U6724 (N_6724,N_6547,N_6565);
nor U6725 (N_6725,N_6491,N_6459);
nor U6726 (N_6726,N_6512,N_6488);
and U6727 (N_6727,N_6478,N_6503);
nand U6728 (N_6728,N_6537,N_6497);
and U6729 (N_6729,N_6508,N_6420);
or U6730 (N_6730,N_6577,N_6527);
nor U6731 (N_6731,N_6438,N_6526);
nor U6732 (N_6732,N_6549,N_6569);
nand U6733 (N_6733,N_6464,N_6408);
nand U6734 (N_6734,N_6435,N_6491);
or U6735 (N_6735,N_6461,N_6454);
or U6736 (N_6736,N_6410,N_6561);
nand U6737 (N_6737,N_6522,N_6436);
nor U6738 (N_6738,N_6473,N_6488);
or U6739 (N_6739,N_6532,N_6460);
nand U6740 (N_6740,N_6576,N_6560);
and U6741 (N_6741,N_6555,N_6476);
and U6742 (N_6742,N_6596,N_6516);
nand U6743 (N_6743,N_6569,N_6419);
or U6744 (N_6744,N_6485,N_6559);
or U6745 (N_6745,N_6594,N_6432);
or U6746 (N_6746,N_6588,N_6596);
or U6747 (N_6747,N_6581,N_6431);
and U6748 (N_6748,N_6490,N_6436);
nand U6749 (N_6749,N_6487,N_6483);
and U6750 (N_6750,N_6402,N_6461);
or U6751 (N_6751,N_6485,N_6548);
or U6752 (N_6752,N_6442,N_6441);
nand U6753 (N_6753,N_6429,N_6516);
nor U6754 (N_6754,N_6535,N_6434);
or U6755 (N_6755,N_6533,N_6535);
nor U6756 (N_6756,N_6474,N_6447);
and U6757 (N_6757,N_6452,N_6438);
or U6758 (N_6758,N_6566,N_6474);
nor U6759 (N_6759,N_6497,N_6477);
or U6760 (N_6760,N_6583,N_6570);
nor U6761 (N_6761,N_6596,N_6478);
nor U6762 (N_6762,N_6532,N_6588);
or U6763 (N_6763,N_6564,N_6593);
nand U6764 (N_6764,N_6542,N_6561);
xnor U6765 (N_6765,N_6545,N_6428);
and U6766 (N_6766,N_6507,N_6564);
nor U6767 (N_6767,N_6519,N_6404);
nand U6768 (N_6768,N_6493,N_6577);
nand U6769 (N_6769,N_6443,N_6584);
nor U6770 (N_6770,N_6543,N_6504);
and U6771 (N_6771,N_6593,N_6562);
nor U6772 (N_6772,N_6496,N_6473);
nor U6773 (N_6773,N_6589,N_6564);
and U6774 (N_6774,N_6471,N_6570);
xor U6775 (N_6775,N_6558,N_6423);
or U6776 (N_6776,N_6576,N_6519);
nand U6777 (N_6777,N_6441,N_6439);
or U6778 (N_6778,N_6407,N_6522);
or U6779 (N_6779,N_6587,N_6571);
or U6780 (N_6780,N_6506,N_6501);
and U6781 (N_6781,N_6434,N_6423);
or U6782 (N_6782,N_6401,N_6510);
nor U6783 (N_6783,N_6516,N_6430);
or U6784 (N_6784,N_6546,N_6469);
nor U6785 (N_6785,N_6478,N_6577);
and U6786 (N_6786,N_6495,N_6589);
and U6787 (N_6787,N_6521,N_6478);
nand U6788 (N_6788,N_6467,N_6591);
and U6789 (N_6789,N_6506,N_6531);
and U6790 (N_6790,N_6553,N_6417);
and U6791 (N_6791,N_6508,N_6425);
and U6792 (N_6792,N_6450,N_6549);
xor U6793 (N_6793,N_6457,N_6439);
and U6794 (N_6794,N_6453,N_6504);
and U6795 (N_6795,N_6464,N_6522);
nand U6796 (N_6796,N_6591,N_6460);
or U6797 (N_6797,N_6567,N_6512);
nand U6798 (N_6798,N_6565,N_6406);
nand U6799 (N_6799,N_6501,N_6581);
or U6800 (N_6800,N_6627,N_6659);
nor U6801 (N_6801,N_6715,N_6622);
nor U6802 (N_6802,N_6698,N_6692);
or U6803 (N_6803,N_6705,N_6759);
and U6804 (N_6804,N_6617,N_6625);
and U6805 (N_6805,N_6666,N_6675);
nand U6806 (N_6806,N_6610,N_6661);
and U6807 (N_6807,N_6785,N_6719);
and U6808 (N_6808,N_6615,N_6762);
nand U6809 (N_6809,N_6652,N_6760);
or U6810 (N_6810,N_6720,N_6729);
nand U6811 (N_6811,N_6711,N_6786);
nor U6812 (N_6812,N_6697,N_6793);
nand U6813 (N_6813,N_6624,N_6693);
or U6814 (N_6814,N_6783,N_6630);
nand U6815 (N_6815,N_6732,N_6601);
or U6816 (N_6816,N_6704,N_6678);
or U6817 (N_6817,N_6743,N_6751);
or U6818 (N_6818,N_6744,N_6618);
or U6819 (N_6819,N_6796,N_6686);
and U6820 (N_6820,N_6670,N_6741);
nand U6821 (N_6821,N_6616,N_6723);
nand U6822 (N_6822,N_6782,N_6792);
nand U6823 (N_6823,N_6763,N_6695);
nor U6824 (N_6824,N_6603,N_6673);
xor U6825 (N_6825,N_6674,N_6749);
nor U6826 (N_6826,N_6799,N_6791);
nand U6827 (N_6827,N_6689,N_6789);
and U6828 (N_6828,N_6716,N_6680);
and U6829 (N_6829,N_6734,N_6702);
nand U6830 (N_6830,N_6605,N_6638);
nand U6831 (N_6831,N_6687,N_6708);
and U6832 (N_6832,N_6777,N_6643);
or U6833 (N_6833,N_6649,N_6608);
nor U6834 (N_6834,N_6747,N_6694);
nor U6835 (N_6835,N_6776,N_6740);
xor U6836 (N_6836,N_6628,N_6737);
and U6837 (N_6837,N_6619,N_6699);
nand U6838 (N_6838,N_6707,N_6644);
and U6839 (N_6839,N_6775,N_6631);
nand U6840 (N_6840,N_6768,N_6733);
nor U6841 (N_6841,N_6611,N_6765);
or U6842 (N_6842,N_6648,N_6798);
or U6843 (N_6843,N_6646,N_6780);
or U6844 (N_6844,N_6685,N_6722);
nor U6845 (N_6845,N_6641,N_6756);
or U6846 (N_6846,N_6683,N_6753);
or U6847 (N_6847,N_6745,N_6781);
xnor U6848 (N_6848,N_6676,N_6653);
nand U6849 (N_6849,N_6614,N_6794);
and U6850 (N_6850,N_6724,N_6736);
nor U6851 (N_6851,N_6677,N_6613);
or U6852 (N_6852,N_6725,N_6769);
or U6853 (N_6853,N_6634,N_6767);
xor U6854 (N_6854,N_6787,N_6713);
and U6855 (N_6855,N_6606,N_6651);
nor U6856 (N_6856,N_6623,N_6612);
nand U6857 (N_6857,N_6773,N_6731);
or U6858 (N_6858,N_6688,N_6672);
and U6859 (N_6859,N_6779,N_6600);
or U6860 (N_6860,N_6764,N_6728);
and U6861 (N_6861,N_6658,N_6607);
and U6862 (N_6862,N_6701,N_6735);
and U6863 (N_6863,N_6621,N_6727);
and U6864 (N_6864,N_6714,N_6691);
and U6865 (N_6865,N_6640,N_6726);
nand U6866 (N_6866,N_6710,N_6750);
nor U6867 (N_6867,N_6682,N_6795);
nand U6868 (N_6868,N_6752,N_6645);
nand U6869 (N_6869,N_6706,N_6730);
nand U6870 (N_6870,N_6718,N_6626);
and U6871 (N_6871,N_6657,N_6656);
or U6872 (N_6872,N_6668,N_6742);
xor U6873 (N_6873,N_6665,N_6774);
nand U6874 (N_6874,N_6721,N_6754);
or U6875 (N_6875,N_6717,N_6669);
nand U6876 (N_6876,N_6609,N_6671);
or U6877 (N_6877,N_6772,N_6770);
and U6878 (N_6878,N_6797,N_6690);
xor U6879 (N_6879,N_6633,N_6778);
and U6880 (N_6880,N_6637,N_6681);
and U6881 (N_6881,N_6604,N_6679);
nor U6882 (N_6882,N_6655,N_6703);
nor U6883 (N_6883,N_6748,N_6790);
nor U6884 (N_6884,N_6660,N_6664);
nor U6885 (N_6885,N_6757,N_6761);
nor U6886 (N_6886,N_6602,N_6788);
or U6887 (N_6887,N_6784,N_6684);
nor U6888 (N_6888,N_6667,N_6712);
nand U6889 (N_6889,N_6663,N_6758);
nand U6890 (N_6890,N_6632,N_6636);
or U6891 (N_6891,N_6639,N_6746);
or U6892 (N_6892,N_6696,N_6738);
or U6893 (N_6893,N_6662,N_6635);
nor U6894 (N_6894,N_6620,N_6629);
or U6895 (N_6895,N_6739,N_6709);
nand U6896 (N_6896,N_6654,N_6771);
or U6897 (N_6897,N_6755,N_6642);
nand U6898 (N_6898,N_6647,N_6766);
and U6899 (N_6899,N_6650,N_6700);
or U6900 (N_6900,N_6737,N_6708);
nand U6901 (N_6901,N_6716,N_6758);
and U6902 (N_6902,N_6737,N_6773);
nand U6903 (N_6903,N_6666,N_6662);
nand U6904 (N_6904,N_6799,N_6758);
nand U6905 (N_6905,N_6666,N_6768);
and U6906 (N_6906,N_6714,N_6643);
nor U6907 (N_6907,N_6612,N_6618);
nand U6908 (N_6908,N_6674,N_6770);
and U6909 (N_6909,N_6731,N_6658);
or U6910 (N_6910,N_6788,N_6714);
or U6911 (N_6911,N_6615,N_6677);
and U6912 (N_6912,N_6791,N_6639);
nand U6913 (N_6913,N_6627,N_6737);
or U6914 (N_6914,N_6726,N_6660);
and U6915 (N_6915,N_6792,N_6639);
nand U6916 (N_6916,N_6638,N_6771);
and U6917 (N_6917,N_6623,N_6709);
nor U6918 (N_6918,N_6631,N_6749);
or U6919 (N_6919,N_6659,N_6687);
and U6920 (N_6920,N_6675,N_6722);
nor U6921 (N_6921,N_6615,N_6717);
or U6922 (N_6922,N_6630,N_6608);
or U6923 (N_6923,N_6716,N_6669);
or U6924 (N_6924,N_6769,N_6759);
nor U6925 (N_6925,N_6737,N_6743);
or U6926 (N_6926,N_6728,N_6644);
or U6927 (N_6927,N_6601,N_6683);
nor U6928 (N_6928,N_6688,N_6631);
nand U6929 (N_6929,N_6601,N_6767);
or U6930 (N_6930,N_6725,N_6660);
or U6931 (N_6931,N_6618,N_6621);
or U6932 (N_6932,N_6725,N_6662);
and U6933 (N_6933,N_6724,N_6600);
nor U6934 (N_6934,N_6697,N_6655);
or U6935 (N_6935,N_6613,N_6792);
or U6936 (N_6936,N_6604,N_6784);
or U6937 (N_6937,N_6643,N_6797);
and U6938 (N_6938,N_6686,N_6644);
nand U6939 (N_6939,N_6614,N_6692);
nor U6940 (N_6940,N_6705,N_6700);
and U6941 (N_6941,N_6625,N_6743);
nor U6942 (N_6942,N_6602,N_6701);
and U6943 (N_6943,N_6719,N_6673);
and U6944 (N_6944,N_6748,N_6708);
xor U6945 (N_6945,N_6619,N_6793);
or U6946 (N_6946,N_6616,N_6722);
and U6947 (N_6947,N_6780,N_6697);
or U6948 (N_6948,N_6763,N_6677);
nand U6949 (N_6949,N_6658,N_6625);
nor U6950 (N_6950,N_6750,N_6787);
and U6951 (N_6951,N_6752,N_6698);
or U6952 (N_6952,N_6790,N_6619);
and U6953 (N_6953,N_6761,N_6732);
or U6954 (N_6954,N_6710,N_6635);
or U6955 (N_6955,N_6727,N_6756);
and U6956 (N_6956,N_6612,N_6798);
nor U6957 (N_6957,N_6647,N_6624);
nor U6958 (N_6958,N_6782,N_6732);
or U6959 (N_6959,N_6741,N_6652);
xor U6960 (N_6960,N_6641,N_6688);
or U6961 (N_6961,N_6725,N_6659);
nor U6962 (N_6962,N_6686,N_6732);
nor U6963 (N_6963,N_6671,N_6678);
xnor U6964 (N_6964,N_6784,N_6647);
and U6965 (N_6965,N_6616,N_6752);
or U6966 (N_6966,N_6722,N_6757);
nand U6967 (N_6967,N_6659,N_6729);
or U6968 (N_6968,N_6746,N_6617);
or U6969 (N_6969,N_6605,N_6697);
and U6970 (N_6970,N_6683,N_6720);
nor U6971 (N_6971,N_6784,N_6722);
or U6972 (N_6972,N_6762,N_6721);
and U6973 (N_6973,N_6651,N_6716);
and U6974 (N_6974,N_6677,N_6606);
and U6975 (N_6975,N_6606,N_6695);
nor U6976 (N_6976,N_6707,N_6789);
or U6977 (N_6977,N_6697,N_6759);
nand U6978 (N_6978,N_6674,N_6698);
nor U6979 (N_6979,N_6753,N_6656);
nand U6980 (N_6980,N_6670,N_6786);
nand U6981 (N_6981,N_6783,N_6712);
nor U6982 (N_6982,N_6791,N_6752);
or U6983 (N_6983,N_6671,N_6665);
and U6984 (N_6984,N_6670,N_6628);
nor U6985 (N_6985,N_6679,N_6676);
nand U6986 (N_6986,N_6677,N_6706);
or U6987 (N_6987,N_6694,N_6730);
nor U6988 (N_6988,N_6777,N_6768);
nor U6989 (N_6989,N_6651,N_6771);
nor U6990 (N_6990,N_6637,N_6779);
and U6991 (N_6991,N_6656,N_6725);
nor U6992 (N_6992,N_6687,N_6726);
nor U6993 (N_6993,N_6743,N_6778);
or U6994 (N_6994,N_6670,N_6669);
nor U6995 (N_6995,N_6671,N_6706);
nor U6996 (N_6996,N_6731,N_6745);
or U6997 (N_6997,N_6644,N_6705);
nor U6998 (N_6998,N_6604,N_6694);
and U6999 (N_6999,N_6670,N_6702);
or U7000 (N_7000,N_6899,N_6846);
or U7001 (N_7001,N_6843,N_6949);
and U7002 (N_7002,N_6978,N_6951);
nor U7003 (N_7003,N_6962,N_6989);
nor U7004 (N_7004,N_6803,N_6825);
and U7005 (N_7005,N_6826,N_6896);
or U7006 (N_7006,N_6854,N_6996);
nand U7007 (N_7007,N_6878,N_6813);
nor U7008 (N_7008,N_6849,N_6927);
or U7009 (N_7009,N_6982,N_6894);
and U7010 (N_7010,N_6935,N_6980);
nor U7011 (N_7011,N_6869,N_6873);
nand U7012 (N_7012,N_6867,N_6850);
nor U7013 (N_7013,N_6955,N_6833);
nand U7014 (N_7014,N_6905,N_6808);
nand U7015 (N_7015,N_6875,N_6883);
or U7016 (N_7016,N_6964,N_6863);
nor U7017 (N_7017,N_6804,N_6811);
nor U7018 (N_7018,N_6966,N_6972);
nor U7019 (N_7019,N_6948,N_6872);
nor U7020 (N_7020,N_6889,N_6998);
and U7021 (N_7021,N_6819,N_6914);
and U7022 (N_7022,N_6834,N_6963);
and U7023 (N_7023,N_6926,N_6992);
or U7024 (N_7024,N_6801,N_6909);
nor U7025 (N_7025,N_6942,N_6810);
or U7026 (N_7026,N_6944,N_6816);
nand U7027 (N_7027,N_6911,N_6973);
xor U7028 (N_7028,N_6877,N_6910);
nand U7029 (N_7029,N_6876,N_6806);
nor U7030 (N_7030,N_6929,N_6895);
nand U7031 (N_7031,N_6925,N_6969);
and U7032 (N_7032,N_6871,N_6897);
nor U7033 (N_7033,N_6977,N_6956);
or U7034 (N_7034,N_6859,N_6979);
or U7035 (N_7035,N_6997,N_6852);
xnor U7036 (N_7036,N_6960,N_6994);
or U7037 (N_7037,N_6991,N_6839);
and U7038 (N_7038,N_6809,N_6892);
nor U7039 (N_7039,N_6965,N_6938);
nor U7040 (N_7040,N_6882,N_6886);
or U7041 (N_7041,N_6890,N_6860);
or U7042 (N_7042,N_6906,N_6968);
nand U7043 (N_7043,N_6837,N_6880);
nor U7044 (N_7044,N_6845,N_6824);
xnor U7045 (N_7045,N_6934,N_6928);
nor U7046 (N_7046,N_6903,N_6884);
nand U7047 (N_7047,N_6908,N_6821);
nor U7048 (N_7048,N_6932,N_6902);
and U7049 (N_7049,N_6836,N_6901);
or U7050 (N_7050,N_6993,N_6832);
nor U7051 (N_7051,N_6817,N_6923);
nor U7052 (N_7052,N_6995,N_6891);
or U7053 (N_7053,N_6933,N_6822);
and U7054 (N_7054,N_6990,N_6898);
or U7055 (N_7055,N_6885,N_6818);
or U7056 (N_7056,N_6842,N_6976);
nor U7057 (N_7057,N_6864,N_6917);
and U7058 (N_7058,N_6970,N_6814);
nor U7059 (N_7059,N_6975,N_6844);
nor U7060 (N_7060,N_6805,N_6987);
and U7061 (N_7061,N_6907,N_6848);
nor U7062 (N_7062,N_6800,N_6967);
nand U7063 (N_7063,N_6835,N_6831);
nand U7064 (N_7064,N_6931,N_6930);
and U7065 (N_7065,N_6865,N_6830);
xor U7066 (N_7066,N_6815,N_6900);
and U7067 (N_7067,N_6866,N_6913);
nor U7068 (N_7068,N_6957,N_6840);
xor U7069 (N_7069,N_6855,N_6904);
and U7070 (N_7070,N_6999,N_6986);
or U7071 (N_7071,N_6879,N_6971);
and U7072 (N_7072,N_6941,N_6954);
xor U7073 (N_7073,N_6838,N_6961);
and U7074 (N_7074,N_6888,N_6856);
nor U7075 (N_7075,N_6812,N_6924);
xnor U7076 (N_7076,N_6915,N_6981);
or U7077 (N_7077,N_6947,N_6823);
or U7078 (N_7078,N_6950,N_6857);
and U7079 (N_7079,N_6916,N_6939);
or U7080 (N_7080,N_6820,N_6945);
and U7081 (N_7081,N_6862,N_6868);
nand U7082 (N_7082,N_6828,N_6841);
or U7083 (N_7083,N_6940,N_6959);
nand U7084 (N_7084,N_6985,N_6988);
nand U7085 (N_7085,N_6921,N_6829);
nor U7086 (N_7086,N_6952,N_6861);
xor U7087 (N_7087,N_6936,N_6920);
or U7088 (N_7088,N_6918,N_6922);
nand U7089 (N_7089,N_6858,N_6958);
and U7090 (N_7090,N_6870,N_6887);
nand U7091 (N_7091,N_6847,N_6946);
nor U7092 (N_7092,N_6853,N_6851);
nand U7093 (N_7093,N_6919,N_6974);
or U7094 (N_7094,N_6874,N_6881);
nand U7095 (N_7095,N_6937,N_6943);
or U7096 (N_7096,N_6827,N_6983);
nand U7097 (N_7097,N_6893,N_6953);
nor U7098 (N_7098,N_6984,N_6912);
or U7099 (N_7099,N_6802,N_6807);
nor U7100 (N_7100,N_6998,N_6838);
and U7101 (N_7101,N_6898,N_6967);
nor U7102 (N_7102,N_6824,N_6803);
or U7103 (N_7103,N_6805,N_6842);
nand U7104 (N_7104,N_6892,N_6973);
nand U7105 (N_7105,N_6823,N_6800);
and U7106 (N_7106,N_6820,N_6847);
and U7107 (N_7107,N_6804,N_6877);
nand U7108 (N_7108,N_6854,N_6889);
nor U7109 (N_7109,N_6939,N_6952);
nand U7110 (N_7110,N_6969,N_6903);
or U7111 (N_7111,N_6830,N_6871);
and U7112 (N_7112,N_6914,N_6887);
and U7113 (N_7113,N_6914,N_6991);
or U7114 (N_7114,N_6822,N_6969);
or U7115 (N_7115,N_6829,N_6936);
nor U7116 (N_7116,N_6882,N_6833);
nor U7117 (N_7117,N_6805,N_6813);
nor U7118 (N_7118,N_6968,N_6861);
nand U7119 (N_7119,N_6822,N_6905);
and U7120 (N_7120,N_6959,N_6882);
nor U7121 (N_7121,N_6917,N_6936);
nand U7122 (N_7122,N_6870,N_6844);
nor U7123 (N_7123,N_6942,N_6843);
or U7124 (N_7124,N_6835,N_6923);
nor U7125 (N_7125,N_6840,N_6865);
and U7126 (N_7126,N_6976,N_6950);
or U7127 (N_7127,N_6970,N_6906);
nand U7128 (N_7128,N_6829,N_6835);
nor U7129 (N_7129,N_6882,N_6926);
nor U7130 (N_7130,N_6999,N_6969);
and U7131 (N_7131,N_6892,N_6932);
or U7132 (N_7132,N_6813,N_6855);
nor U7133 (N_7133,N_6886,N_6849);
nor U7134 (N_7134,N_6947,N_6963);
or U7135 (N_7135,N_6989,N_6992);
and U7136 (N_7136,N_6986,N_6913);
nand U7137 (N_7137,N_6965,N_6940);
or U7138 (N_7138,N_6935,N_6811);
or U7139 (N_7139,N_6989,N_6862);
nor U7140 (N_7140,N_6866,N_6823);
and U7141 (N_7141,N_6990,N_6879);
and U7142 (N_7142,N_6929,N_6897);
nor U7143 (N_7143,N_6810,N_6969);
and U7144 (N_7144,N_6960,N_6859);
nor U7145 (N_7145,N_6894,N_6853);
xor U7146 (N_7146,N_6825,N_6863);
nor U7147 (N_7147,N_6860,N_6843);
nor U7148 (N_7148,N_6997,N_6853);
or U7149 (N_7149,N_6860,N_6852);
and U7150 (N_7150,N_6896,N_6903);
nor U7151 (N_7151,N_6939,N_6943);
or U7152 (N_7152,N_6934,N_6945);
and U7153 (N_7153,N_6919,N_6830);
and U7154 (N_7154,N_6890,N_6962);
and U7155 (N_7155,N_6907,N_6867);
xor U7156 (N_7156,N_6809,N_6924);
nand U7157 (N_7157,N_6913,N_6902);
and U7158 (N_7158,N_6817,N_6836);
nand U7159 (N_7159,N_6853,N_6908);
nand U7160 (N_7160,N_6831,N_6913);
and U7161 (N_7161,N_6942,N_6914);
nand U7162 (N_7162,N_6828,N_6884);
nor U7163 (N_7163,N_6833,N_6938);
nor U7164 (N_7164,N_6994,N_6992);
and U7165 (N_7165,N_6847,N_6903);
and U7166 (N_7166,N_6907,N_6959);
xor U7167 (N_7167,N_6915,N_6849);
or U7168 (N_7168,N_6971,N_6999);
and U7169 (N_7169,N_6818,N_6812);
nor U7170 (N_7170,N_6834,N_6925);
or U7171 (N_7171,N_6831,N_6827);
xor U7172 (N_7172,N_6998,N_6980);
or U7173 (N_7173,N_6966,N_6944);
and U7174 (N_7174,N_6813,N_6918);
and U7175 (N_7175,N_6965,N_6866);
and U7176 (N_7176,N_6943,N_6906);
or U7177 (N_7177,N_6968,N_6850);
nand U7178 (N_7178,N_6887,N_6999);
or U7179 (N_7179,N_6885,N_6864);
or U7180 (N_7180,N_6971,N_6952);
nor U7181 (N_7181,N_6882,N_6943);
nand U7182 (N_7182,N_6852,N_6819);
and U7183 (N_7183,N_6844,N_6857);
nor U7184 (N_7184,N_6927,N_6826);
nor U7185 (N_7185,N_6895,N_6963);
or U7186 (N_7186,N_6949,N_6802);
and U7187 (N_7187,N_6978,N_6880);
xor U7188 (N_7188,N_6858,N_6935);
or U7189 (N_7189,N_6933,N_6969);
xor U7190 (N_7190,N_6934,N_6881);
or U7191 (N_7191,N_6975,N_6815);
or U7192 (N_7192,N_6895,N_6805);
nor U7193 (N_7193,N_6864,N_6861);
nand U7194 (N_7194,N_6942,N_6878);
nor U7195 (N_7195,N_6965,N_6966);
nand U7196 (N_7196,N_6962,N_6830);
nand U7197 (N_7197,N_6971,N_6918);
nand U7198 (N_7198,N_6934,N_6876);
nand U7199 (N_7199,N_6859,N_6834);
nor U7200 (N_7200,N_7199,N_7004);
nand U7201 (N_7201,N_7024,N_7113);
nor U7202 (N_7202,N_7077,N_7128);
or U7203 (N_7203,N_7151,N_7121);
or U7204 (N_7204,N_7053,N_7020);
nor U7205 (N_7205,N_7062,N_7019);
nor U7206 (N_7206,N_7154,N_7099);
and U7207 (N_7207,N_7040,N_7067);
nand U7208 (N_7208,N_7031,N_7102);
nand U7209 (N_7209,N_7167,N_7188);
or U7210 (N_7210,N_7098,N_7017);
or U7211 (N_7211,N_7133,N_7041);
nand U7212 (N_7212,N_7005,N_7139);
and U7213 (N_7213,N_7048,N_7076);
or U7214 (N_7214,N_7089,N_7071);
or U7215 (N_7215,N_7164,N_7138);
nor U7216 (N_7216,N_7184,N_7153);
nor U7217 (N_7217,N_7009,N_7035);
nor U7218 (N_7218,N_7185,N_7174);
or U7219 (N_7219,N_7027,N_7150);
nand U7220 (N_7220,N_7070,N_7110);
and U7221 (N_7221,N_7045,N_7096);
nand U7222 (N_7222,N_7037,N_7000);
nand U7223 (N_7223,N_7021,N_7001);
nand U7224 (N_7224,N_7180,N_7013);
nand U7225 (N_7225,N_7068,N_7125);
nand U7226 (N_7226,N_7175,N_7126);
and U7227 (N_7227,N_7016,N_7039);
nand U7228 (N_7228,N_7119,N_7115);
nand U7229 (N_7229,N_7152,N_7073);
and U7230 (N_7230,N_7131,N_7084);
nor U7231 (N_7231,N_7055,N_7038);
or U7232 (N_7232,N_7085,N_7034);
and U7233 (N_7233,N_7191,N_7108);
xor U7234 (N_7234,N_7047,N_7182);
or U7235 (N_7235,N_7087,N_7163);
nor U7236 (N_7236,N_7132,N_7170);
or U7237 (N_7237,N_7065,N_7118);
nor U7238 (N_7238,N_7074,N_7183);
nor U7239 (N_7239,N_7036,N_7060);
and U7240 (N_7240,N_7127,N_7006);
and U7241 (N_7241,N_7135,N_7157);
nor U7242 (N_7242,N_7111,N_7046);
xor U7243 (N_7243,N_7148,N_7193);
nor U7244 (N_7244,N_7072,N_7026);
and U7245 (N_7245,N_7172,N_7091);
nand U7246 (N_7246,N_7134,N_7082);
nor U7247 (N_7247,N_7018,N_7169);
nor U7248 (N_7248,N_7160,N_7064);
or U7249 (N_7249,N_7114,N_7149);
and U7250 (N_7250,N_7058,N_7141);
and U7251 (N_7251,N_7195,N_7095);
and U7252 (N_7252,N_7156,N_7106);
nand U7253 (N_7253,N_7145,N_7112);
and U7254 (N_7254,N_7173,N_7061);
or U7255 (N_7255,N_7008,N_7130);
nor U7256 (N_7256,N_7162,N_7063);
nand U7257 (N_7257,N_7007,N_7025);
or U7258 (N_7258,N_7181,N_7107);
nor U7259 (N_7259,N_7168,N_7120);
or U7260 (N_7260,N_7176,N_7092);
nor U7261 (N_7261,N_7083,N_7075);
nor U7262 (N_7262,N_7011,N_7088);
nor U7263 (N_7263,N_7050,N_7059);
or U7264 (N_7264,N_7010,N_7147);
or U7265 (N_7265,N_7196,N_7159);
nor U7266 (N_7266,N_7078,N_7144);
nand U7267 (N_7267,N_7002,N_7030);
nand U7268 (N_7268,N_7136,N_7124);
or U7269 (N_7269,N_7178,N_7081);
and U7270 (N_7270,N_7033,N_7103);
xor U7271 (N_7271,N_7043,N_7042);
or U7272 (N_7272,N_7186,N_7093);
and U7273 (N_7273,N_7123,N_7052);
nor U7274 (N_7274,N_7198,N_7094);
nand U7275 (N_7275,N_7056,N_7079);
nand U7276 (N_7276,N_7161,N_7192);
nor U7277 (N_7277,N_7122,N_7101);
nor U7278 (N_7278,N_7146,N_7116);
and U7279 (N_7279,N_7022,N_7189);
nand U7280 (N_7280,N_7032,N_7165);
nand U7281 (N_7281,N_7143,N_7028);
and U7282 (N_7282,N_7069,N_7090);
nand U7283 (N_7283,N_7100,N_7049);
and U7284 (N_7284,N_7190,N_7023);
nor U7285 (N_7285,N_7104,N_7014);
or U7286 (N_7286,N_7171,N_7080);
and U7287 (N_7287,N_7137,N_7044);
and U7288 (N_7288,N_7155,N_7105);
nor U7289 (N_7289,N_7158,N_7015);
nand U7290 (N_7290,N_7066,N_7029);
nand U7291 (N_7291,N_7179,N_7012);
nor U7292 (N_7292,N_7140,N_7177);
nand U7293 (N_7293,N_7097,N_7003);
nand U7294 (N_7294,N_7054,N_7057);
and U7295 (N_7295,N_7109,N_7129);
nand U7296 (N_7296,N_7166,N_7194);
nand U7297 (N_7297,N_7142,N_7117);
nor U7298 (N_7298,N_7197,N_7086);
xor U7299 (N_7299,N_7051,N_7187);
nand U7300 (N_7300,N_7013,N_7000);
and U7301 (N_7301,N_7065,N_7074);
nor U7302 (N_7302,N_7179,N_7024);
or U7303 (N_7303,N_7194,N_7182);
nor U7304 (N_7304,N_7100,N_7126);
and U7305 (N_7305,N_7047,N_7006);
and U7306 (N_7306,N_7051,N_7087);
and U7307 (N_7307,N_7165,N_7166);
nor U7308 (N_7308,N_7038,N_7198);
and U7309 (N_7309,N_7095,N_7104);
nand U7310 (N_7310,N_7073,N_7141);
nand U7311 (N_7311,N_7016,N_7163);
or U7312 (N_7312,N_7054,N_7150);
or U7313 (N_7313,N_7187,N_7055);
nand U7314 (N_7314,N_7053,N_7048);
or U7315 (N_7315,N_7116,N_7042);
and U7316 (N_7316,N_7005,N_7076);
or U7317 (N_7317,N_7037,N_7163);
or U7318 (N_7318,N_7174,N_7118);
nand U7319 (N_7319,N_7062,N_7156);
or U7320 (N_7320,N_7119,N_7088);
nor U7321 (N_7321,N_7120,N_7109);
and U7322 (N_7322,N_7105,N_7137);
and U7323 (N_7323,N_7193,N_7179);
nor U7324 (N_7324,N_7027,N_7031);
nand U7325 (N_7325,N_7021,N_7188);
or U7326 (N_7326,N_7098,N_7030);
xnor U7327 (N_7327,N_7099,N_7037);
nor U7328 (N_7328,N_7109,N_7068);
or U7329 (N_7329,N_7119,N_7117);
nor U7330 (N_7330,N_7022,N_7037);
nor U7331 (N_7331,N_7162,N_7003);
nand U7332 (N_7332,N_7043,N_7186);
nor U7333 (N_7333,N_7067,N_7193);
nand U7334 (N_7334,N_7133,N_7094);
nand U7335 (N_7335,N_7189,N_7063);
nor U7336 (N_7336,N_7125,N_7176);
nor U7337 (N_7337,N_7063,N_7071);
and U7338 (N_7338,N_7124,N_7038);
nand U7339 (N_7339,N_7160,N_7029);
nand U7340 (N_7340,N_7186,N_7154);
or U7341 (N_7341,N_7108,N_7124);
or U7342 (N_7342,N_7165,N_7011);
nand U7343 (N_7343,N_7068,N_7164);
nor U7344 (N_7344,N_7152,N_7028);
nor U7345 (N_7345,N_7043,N_7148);
nand U7346 (N_7346,N_7176,N_7191);
and U7347 (N_7347,N_7093,N_7187);
and U7348 (N_7348,N_7177,N_7076);
and U7349 (N_7349,N_7007,N_7039);
and U7350 (N_7350,N_7198,N_7009);
nor U7351 (N_7351,N_7029,N_7196);
nand U7352 (N_7352,N_7157,N_7103);
or U7353 (N_7353,N_7028,N_7166);
nand U7354 (N_7354,N_7091,N_7185);
or U7355 (N_7355,N_7149,N_7156);
nor U7356 (N_7356,N_7094,N_7079);
nor U7357 (N_7357,N_7148,N_7180);
and U7358 (N_7358,N_7142,N_7007);
and U7359 (N_7359,N_7151,N_7156);
or U7360 (N_7360,N_7072,N_7000);
and U7361 (N_7361,N_7085,N_7110);
nor U7362 (N_7362,N_7169,N_7092);
nor U7363 (N_7363,N_7032,N_7140);
nor U7364 (N_7364,N_7185,N_7104);
nor U7365 (N_7365,N_7198,N_7100);
nor U7366 (N_7366,N_7152,N_7174);
nor U7367 (N_7367,N_7009,N_7188);
nand U7368 (N_7368,N_7112,N_7195);
or U7369 (N_7369,N_7007,N_7009);
nor U7370 (N_7370,N_7118,N_7177);
xnor U7371 (N_7371,N_7195,N_7059);
and U7372 (N_7372,N_7124,N_7113);
nor U7373 (N_7373,N_7042,N_7047);
or U7374 (N_7374,N_7077,N_7080);
nand U7375 (N_7375,N_7047,N_7112);
or U7376 (N_7376,N_7100,N_7146);
or U7377 (N_7377,N_7061,N_7059);
and U7378 (N_7378,N_7031,N_7074);
nand U7379 (N_7379,N_7055,N_7156);
nor U7380 (N_7380,N_7055,N_7199);
and U7381 (N_7381,N_7030,N_7148);
or U7382 (N_7382,N_7002,N_7171);
nand U7383 (N_7383,N_7149,N_7135);
and U7384 (N_7384,N_7157,N_7022);
or U7385 (N_7385,N_7143,N_7005);
or U7386 (N_7386,N_7054,N_7034);
nor U7387 (N_7387,N_7157,N_7168);
nand U7388 (N_7388,N_7148,N_7192);
nor U7389 (N_7389,N_7046,N_7142);
nand U7390 (N_7390,N_7025,N_7150);
and U7391 (N_7391,N_7081,N_7154);
xor U7392 (N_7392,N_7132,N_7056);
or U7393 (N_7393,N_7118,N_7045);
or U7394 (N_7394,N_7117,N_7154);
xnor U7395 (N_7395,N_7126,N_7005);
nor U7396 (N_7396,N_7128,N_7015);
nor U7397 (N_7397,N_7178,N_7089);
and U7398 (N_7398,N_7000,N_7151);
nand U7399 (N_7399,N_7055,N_7036);
nor U7400 (N_7400,N_7324,N_7308);
nand U7401 (N_7401,N_7296,N_7282);
nand U7402 (N_7402,N_7235,N_7220);
and U7403 (N_7403,N_7207,N_7266);
nor U7404 (N_7404,N_7341,N_7323);
and U7405 (N_7405,N_7351,N_7258);
nor U7406 (N_7406,N_7352,N_7377);
and U7407 (N_7407,N_7217,N_7211);
or U7408 (N_7408,N_7290,N_7229);
nor U7409 (N_7409,N_7301,N_7239);
and U7410 (N_7410,N_7236,N_7332);
or U7411 (N_7411,N_7271,N_7264);
or U7412 (N_7412,N_7309,N_7283);
and U7413 (N_7413,N_7303,N_7261);
nor U7414 (N_7414,N_7326,N_7298);
nand U7415 (N_7415,N_7367,N_7322);
nand U7416 (N_7416,N_7294,N_7200);
or U7417 (N_7417,N_7355,N_7230);
nand U7418 (N_7418,N_7209,N_7276);
nor U7419 (N_7419,N_7291,N_7250);
nand U7420 (N_7420,N_7202,N_7218);
nor U7421 (N_7421,N_7399,N_7278);
or U7422 (N_7422,N_7379,N_7317);
nor U7423 (N_7423,N_7320,N_7274);
and U7424 (N_7424,N_7292,N_7225);
nand U7425 (N_7425,N_7255,N_7380);
xor U7426 (N_7426,N_7279,N_7381);
nand U7427 (N_7427,N_7385,N_7299);
or U7428 (N_7428,N_7372,N_7371);
and U7429 (N_7429,N_7215,N_7213);
and U7430 (N_7430,N_7289,N_7210);
nand U7431 (N_7431,N_7306,N_7263);
nor U7432 (N_7432,N_7304,N_7275);
nor U7433 (N_7433,N_7214,N_7391);
nand U7434 (N_7434,N_7302,N_7387);
nand U7435 (N_7435,N_7243,N_7343);
and U7436 (N_7436,N_7262,N_7347);
and U7437 (N_7437,N_7321,N_7319);
nand U7438 (N_7438,N_7314,N_7393);
and U7439 (N_7439,N_7237,N_7226);
or U7440 (N_7440,N_7222,N_7256);
nand U7441 (N_7441,N_7267,N_7336);
nand U7442 (N_7442,N_7313,N_7241);
nor U7443 (N_7443,N_7373,N_7221);
nor U7444 (N_7444,N_7305,N_7281);
nor U7445 (N_7445,N_7375,N_7328);
or U7446 (N_7446,N_7376,N_7334);
and U7447 (N_7447,N_7339,N_7345);
nand U7448 (N_7448,N_7231,N_7201);
and U7449 (N_7449,N_7329,N_7223);
xor U7450 (N_7450,N_7206,N_7318);
and U7451 (N_7451,N_7348,N_7245);
or U7452 (N_7452,N_7398,N_7205);
nor U7453 (N_7453,N_7280,N_7240);
or U7454 (N_7454,N_7254,N_7242);
nor U7455 (N_7455,N_7369,N_7390);
and U7456 (N_7456,N_7316,N_7232);
and U7457 (N_7457,N_7325,N_7286);
or U7458 (N_7458,N_7358,N_7384);
and U7459 (N_7459,N_7395,N_7312);
nand U7460 (N_7460,N_7233,N_7204);
or U7461 (N_7461,N_7260,N_7247);
nor U7462 (N_7462,N_7269,N_7330);
nand U7463 (N_7463,N_7353,N_7310);
nor U7464 (N_7464,N_7364,N_7361);
nor U7465 (N_7465,N_7383,N_7342);
nand U7466 (N_7466,N_7354,N_7272);
or U7467 (N_7467,N_7340,N_7365);
or U7468 (N_7468,N_7337,N_7327);
or U7469 (N_7469,N_7307,N_7259);
nand U7470 (N_7470,N_7219,N_7244);
and U7471 (N_7471,N_7356,N_7311);
nor U7472 (N_7472,N_7378,N_7388);
or U7473 (N_7473,N_7238,N_7397);
or U7474 (N_7474,N_7234,N_7394);
or U7475 (N_7475,N_7257,N_7295);
or U7476 (N_7476,N_7350,N_7300);
and U7477 (N_7477,N_7227,N_7382);
and U7478 (N_7478,N_7333,N_7203);
nand U7479 (N_7479,N_7335,N_7346);
nand U7480 (N_7480,N_7392,N_7252);
nor U7481 (N_7481,N_7228,N_7273);
or U7482 (N_7482,N_7248,N_7251);
or U7483 (N_7483,N_7331,N_7386);
nor U7484 (N_7484,N_7268,N_7370);
and U7485 (N_7485,N_7277,N_7253);
and U7486 (N_7486,N_7246,N_7368);
xor U7487 (N_7487,N_7360,N_7285);
nor U7488 (N_7488,N_7366,N_7265);
and U7489 (N_7489,N_7288,N_7362);
and U7490 (N_7490,N_7344,N_7396);
nand U7491 (N_7491,N_7212,N_7363);
or U7492 (N_7492,N_7224,N_7297);
nand U7493 (N_7493,N_7315,N_7359);
or U7494 (N_7494,N_7208,N_7374);
and U7495 (N_7495,N_7216,N_7270);
and U7496 (N_7496,N_7284,N_7357);
nor U7497 (N_7497,N_7349,N_7389);
nor U7498 (N_7498,N_7338,N_7293);
and U7499 (N_7499,N_7249,N_7287);
nor U7500 (N_7500,N_7309,N_7316);
nor U7501 (N_7501,N_7392,N_7312);
nor U7502 (N_7502,N_7322,N_7341);
and U7503 (N_7503,N_7314,N_7218);
or U7504 (N_7504,N_7343,N_7202);
and U7505 (N_7505,N_7387,N_7325);
and U7506 (N_7506,N_7379,N_7369);
or U7507 (N_7507,N_7353,N_7237);
nand U7508 (N_7508,N_7377,N_7318);
and U7509 (N_7509,N_7375,N_7269);
xnor U7510 (N_7510,N_7330,N_7259);
nand U7511 (N_7511,N_7237,N_7224);
and U7512 (N_7512,N_7326,N_7395);
and U7513 (N_7513,N_7314,N_7262);
or U7514 (N_7514,N_7319,N_7351);
nor U7515 (N_7515,N_7376,N_7287);
nor U7516 (N_7516,N_7259,N_7203);
and U7517 (N_7517,N_7210,N_7216);
or U7518 (N_7518,N_7317,N_7287);
or U7519 (N_7519,N_7225,N_7361);
and U7520 (N_7520,N_7274,N_7269);
and U7521 (N_7521,N_7338,N_7281);
xor U7522 (N_7522,N_7355,N_7357);
or U7523 (N_7523,N_7209,N_7267);
and U7524 (N_7524,N_7323,N_7257);
and U7525 (N_7525,N_7399,N_7346);
xor U7526 (N_7526,N_7258,N_7222);
or U7527 (N_7527,N_7371,N_7385);
nand U7528 (N_7528,N_7252,N_7305);
nor U7529 (N_7529,N_7313,N_7264);
nand U7530 (N_7530,N_7346,N_7289);
or U7531 (N_7531,N_7370,N_7253);
or U7532 (N_7532,N_7248,N_7234);
or U7533 (N_7533,N_7314,N_7299);
and U7534 (N_7534,N_7274,N_7360);
and U7535 (N_7535,N_7291,N_7367);
nand U7536 (N_7536,N_7368,N_7396);
nand U7537 (N_7537,N_7339,N_7373);
or U7538 (N_7538,N_7215,N_7330);
and U7539 (N_7539,N_7246,N_7392);
nor U7540 (N_7540,N_7374,N_7307);
or U7541 (N_7541,N_7234,N_7331);
nor U7542 (N_7542,N_7362,N_7263);
or U7543 (N_7543,N_7347,N_7209);
nand U7544 (N_7544,N_7381,N_7211);
and U7545 (N_7545,N_7358,N_7252);
nor U7546 (N_7546,N_7221,N_7268);
nand U7547 (N_7547,N_7279,N_7278);
and U7548 (N_7548,N_7257,N_7297);
and U7549 (N_7549,N_7396,N_7229);
nor U7550 (N_7550,N_7318,N_7302);
nor U7551 (N_7551,N_7293,N_7389);
nand U7552 (N_7552,N_7395,N_7280);
nand U7553 (N_7553,N_7254,N_7275);
nand U7554 (N_7554,N_7210,N_7247);
nand U7555 (N_7555,N_7287,N_7288);
xnor U7556 (N_7556,N_7333,N_7397);
nand U7557 (N_7557,N_7371,N_7310);
or U7558 (N_7558,N_7278,N_7313);
nor U7559 (N_7559,N_7319,N_7209);
or U7560 (N_7560,N_7252,N_7301);
and U7561 (N_7561,N_7296,N_7396);
and U7562 (N_7562,N_7236,N_7396);
nand U7563 (N_7563,N_7246,N_7312);
nor U7564 (N_7564,N_7214,N_7213);
and U7565 (N_7565,N_7370,N_7312);
nor U7566 (N_7566,N_7230,N_7279);
and U7567 (N_7567,N_7325,N_7354);
and U7568 (N_7568,N_7313,N_7237);
nor U7569 (N_7569,N_7345,N_7201);
and U7570 (N_7570,N_7226,N_7329);
and U7571 (N_7571,N_7349,N_7293);
and U7572 (N_7572,N_7285,N_7299);
nand U7573 (N_7573,N_7292,N_7329);
and U7574 (N_7574,N_7316,N_7201);
nor U7575 (N_7575,N_7234,N_7300);
nand U7576 (N_7576,N_7212,N_7322);
and U7577 (N_7577,N_7242,N_7394);
and U7578 (N_7578,N_7265,N_7284);
nor U7579 (N_7579,N_7396,N_7275);
nor U7580 (N_7580,N_7335,N_7329);
nor U7581 (N_7581,N_7363,N_7310);
nor U7582 (N_7582,N_7266,N_7208);
and U7583 (N_7583,N_7312,N_7224);
xnor U7584 (N_7584,N_7228,N_7314);
and U7585 (N_7585,N_7389,N_7350);
nand U7586 (N_7586,N_7219,N_7276);
xnor U7587 (N_7587,N_7322,N_7276);
or U7588 (N_7588,N_7367,N_7230);
nand U7589 (N_7589,N_7253,N_7331);
or U7590 (N_7590,N_7328,N_7228);
nand U7591 (N_7591,N_7362,N_7277);
nand U7592 (N_7592,N_7329,N_7350);
nor U7593 (N_7593,N_7220,N_7348);
nand U7594 (N_7594,N_7260,N_7374);
and U7595 (N_7595,N_7218,N_7376);
and U7596 (N_7596,N_7228,N_7391);
nor U7597 (N_7597,N_7349,N_7271);
xnor U7598 (N_7598,N_7360,N_7371);
and U7599 (N_7599,N_7330,N_7359);
nand U7600 (N_7600,N_7523,N_7440);
or U7601 (N_7601,N_7555,N_7585);
nand U7602 (N_7602,N_7495,N_7489);
and U7603 (N_7603,N_7561,N_7432);
and U7604 (N_7604,N_7514,N_7461);
and U7605 (N_7605,N_7579,N_7431);
nand U7606 (N_7606,N_7529,N_7481);
or U7607 (N_7607,N_7583,N_7447);
nand U7608 (N_7608,N_7449,N_7546);
and U7609 (N_7609,N_7455,N_7429);
or U7610 (N_7610,N_7571,N_7423);
nand U7611 (N_7611,N_7596,N_7493);
nand U7612 (N_7612,N_7444,N_7487);
xnor U7613 (N_7613,N_7412,N_7451);
nor U7614 (N_7614,N_7470,N_7509);
or U7615 (N_7615,N_7522,N_7434);
and U7616 (N_7616,N_7593,N_7413);
nor U7617 (N_7617,N_7468,N_7511);
nand U7618 (N_7618,N_7516,N_7492);
nand U7619 (N_7619,N_7425,N_7586);
nor U7620 (N_7620,N_7474,N_7454);
nor U7621 (N_7621,N_7537,N_7591);
and U7622 (N_7622,N_7491,N_7581);
nor U7623 (N_7623,N_7452,N_7435);
or U7624 (N_7624,N_7551,N_7521);
or U7625 (N_7625,N_7415,N_7480);
nand U7626 (N_7626,N_7402,N_7498);
or U7627 (N_7627,N_7421,N_7476);
xor U7628 (N_7628,N_7578,N_7408);
or U7629 (N_7629,N_7524,N_7506);
or U7630 (N_7630,N_7515,N_7460);
nor U7631 (N_7631,N_7549,N_7564);
and U7632 (N_7632,N_7598,N_7545);
nor U7633 (N_7633,N_7528,N_7544);
and U7634 (N_7634,N_7490,N_7443);
and U7635 (N_7635,N_7436,N_7482);
or U7636 (N_7636,N_7462,N_7448);
nand U7637 (N_7637,N_7401,N_7483);
or U7638 (N_7638,N_7477,N_7590);
and U7639 (N_7639,N_7594,N_7418);
or U7640 (N_7640,N_7450,N_7539);
or U7641 (N_7641,N_7445,N_7497);
and U7642 (N_7642,N_7428,N_7419);
or U7643 (N_7643,N_7526,N_7456);
nand U7644 (N_7644,N_7488,N_7560);
and U7645 (N_7645,N_7573,N_7486);
and U7646 (N_7646,N_7400,N_7563);
nor U7647 (N_7647,N_7508,N_7533);
and U7648 (N_7648,N_7442,N_7405);
nand U7649 (N_7649,N_7505,N_7439);
and U7650 (N_7650,N_7407,N_7404);
nand U7651 (N_7651,N_7577,N_7588);
nand U7652 (N_7652,N_7513,N_7584);
nand U7653 (N_7653,N_7536,N_7503);
xor U7654 (N_7654,N_7507,N_7430);
and U7655 (N_7655,N_7466,N_7446);
nand U7656 (N_7656,N_7441,N_7599);
nand U7657 (N_7657,N_7531,N_7475);
nor U7658 (N_7658,N_7478,N_7433);
nor U7659 (N_7659,N_7518,N_7530);
and U7660 (N_7660,N_7467,N_7542);
nand U7661 (N_7661,N_7416,N_7473);
nand U7662 (N_7662,N_7438,N_7406);
nor U7663 (N_7663,N_7472,N_7504);
or U7664 (N_7664,N_7566,N_7459);
or U7665 (N_7665,N_7540,N_7485);
or U7666 (N_7666,N_7437,N_7538);
or U7667 (N_7667,N_7567,N_7541);
and U7668 (N_7668,N_7453,N_7414);
nand U7669 (N_7669,N_7420,N_7458);
and U7670 (N_7670,N_7465,N_7422);
nand U7671 (N_7671,N_7574,N_7572);
or U7672 (N_7672,N_7424,N_7548);
or U7673 (N_7673,N_7587,N_7410);
and U7674 (N_7674,N_7427,N_7502);
xor U7675 (N_7675,N_7527,N_7576);
and U7676 (N_7676,N_7457,N_7580);
nor U7677 (N_7677,N_7550,N_7559);
nor U7678 (N_7678,N_7553,N_7525);
or U7679 (N_7679,N_7463,N_7479);
nor U7680 (N_7680,N_7535,N_7595);
nand U7681 (N_7681,N_7597,N_7517);
nand U7682 (N_7682,N_7547,N_7512);
or U7683 (N_7683,N_7501,N_7471);
and U7684 (N_7684,N_7565,N_7556);
or U7685 (N_7685,N_7519,N_7557);
nand U7686 (N_7686,N_7575,N_7589);
and U7687 (N_7687,N_7570,N_7464);
nor U7688 (N_7688,N_7500,N_7417);
and U7689 (N_7689,N_7403,N_7554);
or U7690 (N_7690,N_7534,N_7494);
nand U7691 (N_7691,N_7568,N_7532);
and U7692 (N_7692,N_7592,N_7510);
nand U7693 (N_7693,N_7496,N_7562);
and U7694 (N_7694,N_7543,N_7558);
or U7695 (N_7695,N_7484,N_7469);
xnor U7696 (N_7696,N_7569,N_7409);
and U7697 (N_7697,N_7552,N_7426);
and U7698 (N_7698,N_7499,N_7411);
or U7699 (N_7699,N_7582,N_7520);
nor U7700 (N_7700,N_7432,N_7559);
nand U7701 (N_7701,N_7583,N_7503);
nor U7702 (N_7702,N_7517,N_7465);
or U7703 (N_7703,N_7466,N_7477);
and U7704 (N_7704,N_7554,N_7525);
or U7705 (N_7705,N_7426,N_7481);
or U7706 (N_7706,N_7425,N_7563);
nand U7707 (N_7707,N_7561,N_7509);
nand U7708 (N_7708,N_7441,N_7538);
and U7709 (N_7709,N_7405,N_7558);
and U7710 (N_7710,N_7591,N_7530);
or U7711 (N_7711,N_7497,N_7549);
and U7712 (N_7712,N_7424,N_7411);
or U7713 (N_7713,N_7534,N_7489);
and U7714 (N_7714,N_7475,N_7575);
nor U7715 (N_7715,N_7473,N_7452);
nand U7716 (N_7716,N_7411,N_7500);
nor U7717 (N_7717,N_7518,N_7458);
and U7718 (N_7718,N_7514,N_7498);
nor U7719 (N_7719,N_7593,N_7596);
nand U7720 (N_7720,N_7436,N_7588);
or U7721 (N_7721,N_7549,N_7500);
or U7722 (N_7722,N_7518,N_7425);
nor U7723 (N_7723,N_7549,N_7495);
or U7724 (N_7724,N_7485,N_7575);
nor U7725 (N_7725,N_7546,N_7591);
or U7726 (N_7726,N_7588,N_7427);
and U7727 (N_7727,N_7454,N_7402);
or U7728 (N_7728,N_7490,N_7474);
or U7729 (N_7729,N_7437,N_7409);
and U7730 (N_7730,N_7467,N_7547);
and U7731 (N_7731,N_7452,N_7510);
or U7732 (N_7732,N_7550,N_7435);
nand U7733 (N_7733,N_7523,N_7498);
nor U7734 (N_7734,N_7560,N_7549);
or U7735 (N_7735,N_7485,N_7418);
and U7736 (N_7736,N_7512,N_7567);
or U7737 (N_7737,N_7480,N_7533);
or U7738 (N_7738,N_7488,N_7500);
or U7739 (N_7739,N_7589,N_7560);
and U7740 (N_7740,N_7476,N_7468);
nand U7741 (N_7741,N_7546,N_7533);
and U7742 (N_7742,N_7551,N_7525);
nand U7743 (N_7743,N_7407,N_7592);
and U7744 (N_7744,N_7419,N_7598);
nor U7745 (N_7745,N_7483,N_7506);
nor U7746 (N_7746,N_7443,N_7488);
nor U7747 (N_7747,N_7535,N_7455);
nor U7748 (N_7748,N_7594,N_7523);
or U7749 (N_7749,N_7575,N_7456);
and U7750 (N_7750,N_7406,N_7457);
nor U7751 (N_7751,N_7538,N_7462);
nor U7752 (N_7752,N_7584,N_7593);
and U7753 (N_7753,N_7407,N_7411);
nor U7754 (N_7754,N_7490,N_7453);
and U7755 (N_7755,N_7544,N_7467);
nand U7756 (N_7756,N_7479,N_7488);
nor U7757 (N_7757,N_7590,N_7539);
or U7758 (N_7758,N_7517,N_7479);
nor U7759 (N_7759,N_7462,N_7531);
xnor U7760 (N_7760,N_7526,N_7584);
or U7761 (N_7761,N_7559,N_7571);
nor U7762 (N_7762,N_7537,N_7426);
and U7763 (N_7763,N_7535,N_7466);
nor U7764 (N_7764,N_7404,N_7586);
or U7765 (N_7765,N_7548,N_7453);
or U7766 (N_7766,N_7542,N_7429);
and U7767 (N_7767,N_7474,N_7516);
nand U7768 (N_7768,N_7439,N_7409);
nor U7769 (N_7769,N_7464,N_7479);
nor U7770 (N_7770,N_7453,N_7593);
xnor U7771 (N_7771,N_7527,N_7446);
and U7772 (N_7772,N_7574,N_7567);
or U7773 (N_7773,N_7518,N_7408);
or U7774 (N_7774,N_7422,N_7545);
and U7775 (N_7775,N_7572,N_7587);
or U7776 (N_7776,N_7432,N_7470);
nand U7777 (N_7777,N_7414,N_7597);
and U7778 (N_7778,N_7479,N_7558);
or U7779 (N_7779,N_7529,N_7496);
or U7780 (N_7780,N_7444,N_7406);
nor U7781 (N_7781,N_7547,N_7401);
nand U7782 (N_7782,N_7469,N_7561);
nor U7783 (N_7783,N_7579,N_7556);
or U7784 (N_7784,N_7561,N_7555);
or U7785 (N_7785,N_7576,N_7548);
and U7786 (N_7786,N_7535,N_7597);
nand U7787 (N_7787,N_7522,N_7546);
nor U7788 (N_7788,N_7591,N_7503);
and U7789 (N_7789,N_7412,N_7568);
and U7790 (N_7790,N_7511,N_7546);
or U7791 (N_7791,N_7547,N_7409);
nand U7792 (N_7792,N_7492,N_7482);
nor U7793 (N_7793,N_7444,N_7436);
nand U7794 (N_7794,N_7418,N_7441);
nand U7795 (N_7795,N_7559,N_7426);
and U7796 (N_7796,N_7413,N_7493);
nor U7797 (N_7797,N_7430,N_7529);
and U7798 (N_7798,N_7594,N_7472);
or U7799 (N_7799,N_7526,N_7512);
nand U7800 (N_7800,N_7706,N_7799);
and U7801 (N_7801,N_7632,N_7736);
and U7802 (N_7802,N_7780,N_7631);
and U7803 (N_7803,N_7650,N_7749);
nand U7804 (N_7804,N_7619,N_7759);
or U7805 (N_7805,N_7621,N_7757);
and U7806 (N_7806,N_7689,N_7639);
or U7807 (N_7807,N_7748,N_7646);
or U7808 (N_7808,N_7755,N_7788);
and U7809 (N_7809,N_7781,N_7658);
or U7810 (N_7810,N_7662,N_7610);
nand U7811 (N_7811,N_7665,N_7681);
or U7812 (N_7812,N_7764,N_7645);
nor U7813 (N_7813,N_7737,N_7739);
nor U7814 (N_7814,N_7654,N_7611);
nand U7815 (N_7815,N_7684,N_7740);
or U7816 (N_7816,N_7769,N_7742);
nand U7817 (N_7817,N_7783,N_7734);
and U7818 (N_7818,N_7660,N_7672);
or U7819 (N_7819,N_7745,N_7655);
xor U7820 (N_7820,N_7784,N_7702);
or U7821 (N_7821,N_7765,N_7791);
and U7822 (N_7822,N_7679,N_7717);
nor U7823 (N_7823,N_7715,N_7793);
or U7824 (N_7824,N_7648,N_7713);
and U7825 (N_7825,N_7667,N_7735);
xor U7826 (N_7826,N_7721,N_7692);
nor U7827 (N_7827,N_7612,N_7618);
and U7828 (N_7828,N_7615,N_7635);
or U7829 (N_7829,N_7756,N_7698);
nand U7830 (N_7830,N_7602,N_7709);
nor U7831 (N_7831,N_7629,N_7644);
or U7832 (N_7832,N_7703,N_7763);
or U7833 (N_7833,N_7704,N_7601);
or U7834 (N_7834,N_7607,N_7640);
or U7835 (N_7835,N_7637,N_7664);
xor U7836 (N_7836,N_7643,N_7790);
nor U7837 (N_7837,N_7787,N_7733);
nand U7838 (N_7838,N_7718,N_7760);
or U7839 (N_7839,N_7731,N_7753);
and U7840 (N_7840,N_7633,N_7777);
nor U7841 (N_7841,N_7685,N_7673);
nand U7842 (N_7842,N_7636,N_7659);
nor U7843 (N_7843,N_7642,N_7649);
or U7844 (N_7844,N_7700,N_7716);
and U7845 (N_7845,N_7691,N_7729);
and U7846 (N_7846,N_7669,N_7626);
nor U7847 (N_7847,N_7786,N_7798);
or U7848 (N_7848,N_7688,N_7627);
xor U7849 (N_7849,N_7779,N_7675);
or U7850 (N_7850,N_7604,N_7705);
nand U7851 (N_7851,N_7747,N_7624);
nand U7852 (N_7852,N_7670,N_7617);
and U7853 (N_7853,N_7775,N_7778);
nand U7854 (N_7854,N_7711,N_7680);
and U7855 (N_7855,N_7647,N_7725);
nand U7856 (N_7856,N_7651,N_7652);
nand U7857 (N_7857,N_7714,N_7693);
nor U7858 (N_7858,N_7634,N_7744);
or U7859 (N_7859,N_7690,N_7794);
and U7860 (N_7860,N_7767,N_7708);
and U7861 (N_7861,N_7726,N_7656);
and U7862 (N_7862,N_7761,N_7609);
xnor U7863 (N_7863,N_7728,N_7710);
or U7864 (N_7864,N_7625,N_7653);
or U7865 (N_7865,N_7797,N_7641);
or U7866 (N_7866,N_7677,N_7789);
nor U7867 (N_7867,N_7657,N_7730);
nand U7868 (N_7868,N_7623,N_7697);
nor U7869 (N_7869,N_7683,N_7608);
nand U7870 (N_7870,N_7603,N_7613);
nand U7871 (N_7871,N_7600,N_7720);
and U7872 (N_7872,N_7614,N_7622);
and U7873 (N_7873,N_7682,N_7638);
nand U7874 (N_7874,N_7616,N_7738);
and U7875 (N_7875,N_7687,N_7671);
or U7876 (N_7876,N_7686,N_7727);
nor U7877 (N_7877,N_7782,N_7751);
or U7878 (N_7878,N_7661,N_7796);
nand U7879 (N_7879,N_7766,N_7771);
xor U7880 (N_7880,N_7754,N_7668);
or U7881 (N_7881,N_7758,N_7776);
and U7882 (N_7882,N_7723,N_7722);
and U7883 (N_7883,N_7743,N_7719);
or U7884 (N_7884,N_7774,N_7741);
and U7885 (N_7885,N_7605,N_7666);
nand U7886 (N_7886,N_7768,N_7732);
nor U7887 (N_7887,N_7694,N_7772);
nor U7888 (N_7888,N_7785,N_7630);
or U7889 (N_7889,N_7712,N_7678);
nor U7890 (N_7890,N_7701,N_7606);
and U7891 (N_7891,N_7674,N_7750);
nor U7892 (N_7892,N_7676,N_7792);
or U7893 (N_7893,N_7663,N_7770);
nor U7894 (N_7894,N_7620,N_7746);
nor U7895 (N_7895,N_7699,N_7695);
nand U7896 (N_7896,N_7752,N_7696);
xnor U7897 (N_7897,N_7707,N_7795);
or U7898 (N_7898,N_7724,N_7762);
nand U7899 (N_7899,N_7628,N_7773);
nor U7900 (N_7900,N_7770,N_7790);
and U7901 (N_7901,N_7688,N_7648);
or U7902 (N_7902,N_7751,N_7679);
nor U7903 (N_7903,N_7700,N_7686);
nor U7904 (N_7904,N_7703,N_7715);
or U7905 (N_7905,N_7675,N_7644);
or U7906 (N_7906,N_7711,N_7631);
or U7907 (N_7907,N_7652,N_7722);
nand U7908 (N_7908,N_7760,N_7746);
or U7909 (N_7909,N_7646,N_7638);
and U7910 (N_7910,N_7655,N_7639);
or U7911 (N_7911,N_7791,N_7769);
nor U7912 (N_7912,N_7745,N_7736);
or U7913 (N_7913,N_7683,N_7638);
or U7914 (N_7914,N_7712,N_7785);
or U7915 (N_7915,N_7624,N_7680);
and U7916 (N_7916,N_7651,N_7658);
nor U7917 (N_7917,N_7715,N_7601);
and U7918 (N_7918,N_7716,N_7778);
or U7919 (N_7919,N_7625,N_7680);
nand U7920 (N_7920,N_7701,N_7664);
nor U7921 (N_7921,N_7741,N_7728);
and U7922 (N_7922,N_7690,N_7610);
nand U7923 (N_7923,N_7601,N_7724);
nor U7924 (N_7924,N_7653,N_7683);
and U7925 (N_7925,N_7646,N_7754);
nand U7926 (N_7926,N_7644,N_7767);
nor U7927 (N_7927,N_7629,N_7714);
or U7928 (N_7928,N_7611,N_7766);
and U7929 (N_7929,N_7654,N_7629);
or U7930 (N_7930,N_7748,N_7754);
nor U7931 (N_7931,N_7767,N_7728);
or U7932 (N_7932,N_7623,N_7746);
nand U7933 (N_7933,N_7748,N_7747);
nand U7934 (N_7934,N_7787,N_7691);
nand U7935 (N_7935,N_7774,N_7756);
or U7936 (N_7936,N_7645,N_7739);
and U7937 (N_7937,N_7728,N_7659);
nor U7938 (N_7938,N_7757,N_7762);
nor U7939 (N_7939,N_7726,N_7629);
nor U7940 (N_7940,N_7696,N_7745);
nand U7941 (N_7941,N_7798,N_7702);
xor U7942 (N_7942,N_7691,N_7649);
nand U7943 (N_7943,N_7727,N_7698);
and U7944 (N_7944,N_7735,N_7619);
nand U7945 (N_7945,N_7759,N_7615);
and U7946 (N_7946,N_7730,N_7728);
or U7947 (N_7947,N_7698,N_7654);
or U7948 (N_7948,N_7698,N_7609);
or U7949 (N_7949,N_7746,N_7630);
and U7950 (N_7950,N_7674,N_7797);
nand U7951 (N_7951,N_7691,N_7646);
or U7952 (N_7952,N_7695,N_7609);
or U7953 (N_7953,N_7665,N_7608);
nand U7954 (N_7954,N_7773,N_7604);
nand U7955 (N_7955,N_7676,N_7789);
nor U7956 (N_7956,N_7684,N_7768);
nor U7957 (N_7957,N_7740,N_7797);
nor U7958 (N_7958,N_7732,N_7645);
or U7959 (N_7959,N_7649,N_7675);
xnor U7960 (N_7960,N_7634,N_7653);
nand U7961 (N_7961,N_7760,N_7729);
or U7962 (N_7962,N_7698,N_7613);
nand U7963 (N_7963,N_7668,N_7732);
and U7964 (N_7964,N_7633,N_7674);
and U7965 (N_7965,N_7640,N_7757);
or U7966 (N_7966,N_7724,N_7653);
or U7967 (N_7967,N_7756,N_7632);
and U7968 (N_7968,N_7745,N_7699);
and U7969 (N_7969,N_7704,N_7624);
nand U7970 (N_7970,N_7626,N_7641);
nand U7971 (N_7971,N_7716,N_7753);
and U7972 (N_7972,N_7769,N_7745);
nand U7973 (N_7973,N_7613,N_7721);
or U7974 (N_7974,N_7774,N_7696);
and U7975 (N_7975,N_7607,N_7785);
xnor U7976 (N_7976,N_7632,N_7668);
or U7977 (N_7977,N_7757,N_7710);
nor U7978 (N_7978,N_7691,N_7759);
nand U7979 (N_7979,N_7739,N_7696);
and U7980 (N_7980,N_7775,N_7714);
nand U7981 (N_7981,N_7633,N_7787);
xnor U7982 (N_7982,N_7634,N_7773);
nand U7983 (N_7983,N_7727,N_7648);
xnor U7984 (N_7984,N_7718,N_7678);
nor U7985 (N_7985,N_7768,N_7757);
and U7986 (N_7986,N_7613,N_7648);
or U7987 (N_7987,N_7620,N_7633);
nand U7988 (N_7988,N_7783,N_7658);
and U7989 (N_7989,N_7766,N_7671);
or U7990 (N_7990,N_7602,N_7727);
and U7991 (N_7991,N_7724,N_7676);
or U7992 (N_7992,N_7796,N_7612);
and U7993 (N_7993,N_7795,N_7655);
nor U7994 (N_7994,N_7628,N_7603);
or U7995 (N_7995,N_7764,N_7605);
and U7996 (N_7996,N_7610,N_7650);
nand U7997 (N_7997,N_7662,N_7667);
and U7998 (N_7998,N_7784,N_7675);
or U7999 (N_7999,N_7692,N_7718);
or U8000 (N_8000,N_7923,N_7937);
or U8001 (N_8001,N_7958,N_7864);
nor U8002 (N_8002,N_7991,N_7850);
and U8003 (N_8003,N_7944,N_7874);
nand U8004 (N_8004,N_7969,N_7911);
or U8005 (N_8005,N_7854,N_7856);
nor U8006 (N_8006,N_7838,N_7857);
nor U8007 (N_8007,N_7842,N_7921);
nor U8008 (N_8008,N_7908,N_7974);
nor U8009 (N_8009,N_7929,N_7881);
nand U8010 (N_8010,N_7887,N_7953);
or U8011 (N_8011,N_7815,N_7833);
nand U8012 (N_8012,N_7938,N_7810);
and U8013 (N_8013,N_7878,N_7860);
and U8014 (N_8014,N_7822,N_7992);
or U8015 (N_8015,N_7903,N_7951);
nand U8016 (N_8016,N_7843,N_7862);
nor U8017 (N_8017,N_7806,N_7895);
nand U8018 (N_8018,N_7970,N_7826);
xnor U8019 (N_8019,N_7845,N_7914);
xor U8020 (N_8020,N_7891,N_7859);
and U8021 (N_8021,N_7883,N_7886);
nand U8022 (N_8022,N_7959,N_7972);
nor U8023 (N_8023,N_7851,N_7831);
nor U8024 (N_8024,N_7888,N_7968);
nand U8025 (N_8025,N_7976,N_7917);
and U8026 (N_8026,N_7997,N_7824);
nand U8027 (N_8027,N_7852,N_7830);
or U8028 (N_8028,N_7947,N_7990);
or U8029 (N_8029,N_7933,N_7812);
or U8030 (N_8030,N_7880,N_7855);
nor U8031 (N_8031,N_7912,N_7834);
nor U8032 (N_8032,N_7966,N_7873);
and U8033 (N_8033,N_7853,N_7863);
nor U8034 (N_8034,N_7920,N_7896);
and U8035 (N_8035,N_7820,N_7890);
or U8036 (N_8036,N_7954,N_7889);
nor U8037 (N_8037,N_7924,N_7829);
or U8038 (N_8038,N_7870,N_7823);
and U8039 (N_8039,N_7910,N_7871);
and U8040 (N_8040,N_7978,N_7807);
and U8041 (N_8041,N_7861,N_7986);
nand U8042 (N_8042,N_7865,N_7835);
nor U8043 (N_8043,N_7902,N_7918);
and U8044 (N_8044,N_7821,N_7981);
or U8045 (N_8045,N_7872,N_7805);
or U8046 (N_8046,N_7808,N_7922);
nand U8047 (N_8047,N_7956,N_7939);
nand U8048 (N_8048,N_7876,N_7819);
nor U8049 (N_8049,N_7868,N_7905);
nand U8050 (N_8050,N_7932,N_7915);
nor U8051 (N_8051,N_7975,N_7955);
nor U8052 (N_8052,N_7841,N_7867);
and U8053 (N_8053,N_7900,N_7899);
or U8054 (N_8054,N_7893,N_7879);
nand U8055 (N_8055,N_7875,N_7935);
xor U8056 (N_8056,N_7963,N_7832);
nor U8057 (N_8057,N_7809,N_7985);
nor U8058 (N_8058,N_7919,N_7901);
or U8059 (N_8059,N_7803,N_7952);
xor U8060 (N_8060,N_7816,N_7931);
nor U8061 (N_8061,N_7877,N_7836);
nand U8062 (N_8062,N_7849,N_7847);
nand U8063 (N_8063,N_7898,N_7892);
xnor U8064 (N_8064,N_7993,N_7943);
and U8065 (N_8065,N_7999,N_7949);
or U8066 (N_8066,N_7946,N_7934);
and U8067 (N_8067,N_7804,N_7936);
and U8068 (N_8068,N_7884,N_7961);
nand U8069 (N_8069,N_7945,N_7825);
nor U8070 (N_8070,N_7828,N_7840);
nor U8071 (N_8071,N_7967,N_7817);
nand U8072 (N_8072,N_7988,N_7960);
or U8073 (N_8073,N_7925,N_7894);
or U8074 (N_8074,N_7957,N_7801);
nand U8075 (N_8075,N_7971,N_7907);
and U8076 (N_8076,N_7980,N_7998);
nand U8077 (N_8077,N_7965,N_7964);
and U8078 (N_8078,N_7909,N_7942);
and U8079 (N_8079,N_7882,N_7800);
and U8080 (N_8080,N_7897,N_7941);
nand U8081 (N_8081,N_7948,N_7928);
or U8082 (N_8082,N_7813,N_7846);
nand U8083 (N_8083,N_7987,N_7996);
or U8084 (N_8084,N_7848,N_7818);
nor U8085 (N_8085,N_7979,N_7869);
and U8086 (N_8086,N_7973,N_7913);
nand U8087 (N_8087,N_7904,N_7844);
nand U8088 (N_8088,N_7916,N_7811);
nand U8089 (N_8089,N_7989,N_7837);
or U8090 (N_8090,N_7858,N_7983);
and U8091 (N_8091,N_7885,N_7866);
and U8092 (N_8092,N_7940,N_7977);
nor U8093 (N_8093,N_7906,N_7802);
nor U8094 (N_8094,N_7814,N_7950);
or U8095 (N_8095,N_7984,N_7962);
and U8096 (N_8096,N_7927,N_7982);
nor U8097 (N_8097,N_7994,N_7926);
or U8098 (N_8098,N_7930,N_7995);
nor U8099 (N_8099,N_7839,N_7827);
nand U8100 (N_8100,N_7947,N_7928);
or U8101 (N_8101,N_7852,N_7960);
nor U8102 (N_8102,N_7863,N_7919);
and U8103 (N_8103,N_7825,N_7815);
nand U8104 (N_8104,N_7890,N_7831);
nor U8105 (N_8105,N_7836,N_7806);
nor U8106 (N_8106,N_7837,N_7816);
nor U8107 (N_8107,N_7944,N_7994);
nor U8108 (N_8108,N_7814,N_7828);
nor U8109 (N_8109,N_7856,N_7872);
and U8110 (N_8110,N_7800,N_7965);
or U8111 (N_8111,N_7818,N_7948);
and U8112 (N_8112,N_7857,N_7880);
nand U8113 (N_8113,N_7862,N_7889);
nor U8114 (N_8114,N_7900,N_7974);
and U8115 (N_8115,N_7896,N_7925);
and U8116 (N_8116,N_7901,N_7953);
nand U8117 (N_8117,N_7880,N_7997);
nor U8118 (N_8118,N_7880,N_7840);
or U8119 (N_8119,N_7826,N_7908);
nor U8120 (N_8120,N_7970,N_7959);
or U8121 (N_8121,N_7998,N_7811);
nand U8122 (N_8122,N_7889,N_7935);
nor U8123 (N_8123,N_7865,N_7850);
or U8124 (N_8124,N_7961,N_7869);
nand U8125 (N_8125,N_7960,N_7879);
nor U8126 (N_8126,N_7817,N_7902);
nor U8127 (N_8127,N_7878,N_7969);
nor U8128 (N_8128,N_7932,N_7957);
nor U8129 (N_8129,N_7937,N_7842);
and U8130 (N_8130,N_7942,N_7810);
or U8131 (N_8131,N_7964,N_7857);
and U8132 (N_8132,N_7806,N_7918);
and U8133 (N_8133,N_7848,N_7982);
or U8134 (N_8134,N_7904,N_7895);
nand U8135 (N_8135,N_7907,N_7960);
or U8136 (N_8136,N_7825,N_7959);
and U8137 (N_8137,N_7822,N_7896);
and U8138 (N_8138,N_7880,N_7828);
nor U8139 (N_8139,N_7888,N_7918);
nand U8140 (N_8140,N_7964,N_7981);
or U8141 (N_8141,N_7913,N_7990);
nand U8142 (N_8142,N_7885,N_7850);
nor U8143 (N_8143,N_7839,N_7896);
and U8144 (N_8144,N_7957,N_7919);
nor U8145 (N_8145,N_7827,N_7972);
and U8146 (N_8146,N_7844,N_7819);
and U8147 (N_8147,N_7929,N_7842);
or U8148 (N_8148,N_7895,N_7950);
nand U8149 (N_8149,N_7863,N_7910);
and U8150 (N_8150,N_7979,N_7847);
or U8151 (N_8151,N_7912,N_7955);
nor U8152 (N_8152,N_7813,N_7844);
nor U8153 (N_8153,N_7840,N_7939);
and U8154 (N_8154,N_7821,N_7833);
nand U8155 (N_8155,N_7880,N_7951);
nor U8156 (N_8156,N_7883,N_7869);
nand U8157 (N_8157,N_7859,N_7994);
nand U8158 (N_8158,N_7900,N_7926);
or U8159 (N_8159,N_7980,N_7839);
nor U8160 (N_8160,N_7888,N_7800);
nand U8161 (N_8161,N_7983,N_7882);
or U8162 (N_8162,N_7886,N_7991);
nand U8163 (N_8163,N_7967,N_7911);
or U8164 (N_8164,N_7846,N_7821);
or U8165 (N_8165,N_7904,N_7886);
nor U8166 (N_8166,N_7921,N_7841);
or U8167 (N_8167,N_7841,N_7932);
and U8168 (N_8168,N_7911,N_7974);
nand U8169 (N_8169,N_7813,N_7802);
nor U8170 (N_8170,N_7806,N_7828);
and U8171 (N_8171,N_7976,N_7835);
or U8172 (N_8172,N_7873,N_7970);
or U8173 (N_8173,N_7942,N_7990);
and U8174 (N_8174,N_7927,N_7970);
and U8175 (N_8175,N_7884,N_7887);
or U8176 (N_8176,N_7849,N_7917);
nand U8177 (N_8177,N_7976,N_7993);
or U8178 (N_8178,N_7961,N_7905);
or U8179 (N_8179,N_7849,N_7882);
or U8180 (N_8180,N_7986,N_7928);
nand U8181 (N_8181,N_7988,N_7966);
nor U8182 (N_8182,N_7922,N_7993);
nor U8183 (N_8183,N_7945,N_7965);
and U8184 (N_8184,N_7975,N_7988);
or U8185 (N_8185,N_7819,N_7920);
and U8186 (N_8186,N_7965,N_7818);
nor U8187 (N_8187,N_7997,N_7931);
and U8188 (N_8188,N_7968,N_7831);
or U8189 (N_8189,N_7858,N_7950);
and U8190 (N_8190,N_7950,N_7927);
or U8191 (N_8191,N_7984,N_7959);
nand U8192 (N_8192,N_7997,N_7832);
or U8193 (N_8193,N_7825,N_7951);
nor U8194 (N_8194,N_7938,N_7936);
and U8195 (N_8195,N_7848,N_7990);
nand U8196 (N_8196,N_7943,N_7987);
nor U8197 (N_8197,N_7940,N_7927);
and U8198 (N_8198,N_7890,N_7862);
nor U8199 (N_8199,N_7996,N_7811);
nor U8200 (N_8200,N_8169,N_8011);
or U8201 (N_8201,N_8013,N_8110);
and U8202 (N_8202,N_8053,N_8117);
and U8203 (N_8203,N_8015,N_8083);
nor U8204 (N_8204,N_8174,N_8033);
nor U8205 (N_8205,N_8163,N_8170);
nand U8206 (N_8206,N_8104,N_8161);
xnor U8207 (N_8207,N_8040,N_8115);
nor U8208 (N_8208,N_8096,N_8128);
and U8209 (N_8209,N_8063,N_8078);
and U8210 (N_8210,N_8131,N_8024);
and U8211 (N_8211,N_8003,N_8106);
nor U8212 (N_8212,N_8025,N_8031);
and U8213 (N_8213,N_8046,N_8137);
nor U8214 (N_8214,N_8178,N_8149);
nor U8215 (N_8215,N_8026,N_8043);
and U8216 (N_8216,N_8060,N_8181);
or U8217 (N_8217,N_8176,N_8114);
nor U8218 (N_8218,N_8165,N_8172);
or U8219 (N_8219,N_8134,N_8132);
xor U8220 (N_8220,N_8085,N_8167);
nand U8221 (N_8221,N_8099,N_8067);
or U8222 (N_8222,N_8111,N_8194);
and U8223 (N_8223,N_8023,N_8069);
or U8224 (N_8224,N_8092,N_8120);
nor U8225 (N_8225,N_8034,N_8183);
nor U8226 (N_8226,N_8101,N_8164);
nor U8227 (N_8227,N_8074,N_8056);
nand U8228 (N_8228,N_8080,N_8029);
and U8229 (N_8229,N_8156,N_8190);
nand U8230 (N_8230,N_8150,N_8144);
nand U8231 (N_8231,N_8135,N_8180);
nor U8232 (N_8232,N_8084,N_8058);
nand U8233 (N_8233,N_8186,N_8059);
or U8234 (N_8234,N_8103,N_8151);
or U8235 (N_8235,N_8038,N_8062);
nor U8236 (N_8236,N_8065,N_8055);
nand U8237 (N_8237,N_8197,N_8154);
and U8238 (N_8238,N_8079,N_8054);
nor U8239 (N_8239,N_8073,N_8061);
and U8240 (N_8240,N_8009,N_8173);
or U8241 (N_8241,N_8094,N_8121);
nand U8242 (N_8242,N_8095,N_8116);
nor U8243 (N_8243,N_8126,N_8051);
nor U8244 (N_8244,N_8097,N_8019);
or U8245 (N_8245,N_8123,N_8010);
and U8246 (N_8246,N_8168,N_8005);
or U8247 (N_8247,N_8159,N_8050);
and U8248 (N_8248,N_8036,N_8185);
or U8249 (N_8249,N_8157,N_8153);
or U8250 (N_8250,N_8192,N_8158);
nand U8251 (N_8251,N_8048,N_8160);
and U8252 (N_8252,N_8018,N_8027);
or U8253 (N_8253,N_8093,N_8112);
or U8254 (N_8254,N_8130,N_8166);
and U8255 (N_8255,N_8017,N_8057);
nand U8256 (N_8256,N_8066,N_8146);
and U8257 (N_8257,N_8087,N_8070);
nand U8258 (N_8258,N_8090,N_8039);
nor U8259 (N_8259,N_8102,N_8012);
nand U8260 (N_8260,N_8072,N_8196);
xor U8261 (N_8261,N_8136,N_8171);
or U8262 (N_8262,N_8047,N_8145);
and U8263 (N_8263,N_8077,N_8091);
xnor U8264 (N_8264,N_8139,N_8098);
or U8265 (N_8265,N_8022,N_8141);
or U8266 (N_8266,N_8037,N_8014);
nand U8267 (N_8267,N_8199,N_8042);
nor U8268 (N_8268,N_8032,N_8142);
nand U8269 (N_8269,N_8075,N_8089);
or U8270 (N_8270,N_8041,N_8044);
nor U8271 (N_8271,N_8081,N_8035);
nand U8272 (N_8272,N_8088,N_8086);
nand U8273 (N_8273,N_8155,N_8107);
or U8274 (N_8274,N_8184,N_8100);
or U8275 (N_8275,N_8068,N_8129);
nor U8276 (N_8276,N_8133,N_8105);
or U8277 (N_8277,N_8030,N_8076);
nor U8278 (N_8278,N_8109,N_8020);
and U8279 (N_8279,N_8001,N_8187);
nor U8280 (N_8280,N_8148,N_8140);
and U8281 (N_8281,N_8175,N_8189);
or U8282 (N_8282,N_8188,N_8045);
or U8283 (N_8283,N_8198,N_8124);
and U8284 (N_8284,N_8064,N_8119);
nor U8285 (N_8285,N_8177,N_8147);
xor U8286 (N_8286,N_8108,N_8127);
xnor U8287 (N_8287,N_8052,N_8113);
nand U8288 (N_8288,N_8162,N_8049);
nand U8289 (N_8289,N_8191,N_8000);
or U8290 (N_8290,N_8138,N_8195);
nor U8291 (N_8291,N_8021,N_8143);
or U8292 (N_8292,N_8193,N_8122);
and U8293 (N_8293,N_8004,N_8002);
or U8294 (N_8294,N_8006,N_8028);
or U8295 (N_8295,N_8125,N_8152);
nand U8296 (N_8296,N_8179,N_8008);
nor U8297 (N_8297,N_8182,N_8082);
and U8298 (N_8298,N_8007,N_8118);
or U8299 (N_8299,N_8071,N_8016);
nand U8300 (N_8300,N_8075,N_8024);
or U8301 (N_8301,N_8103,N_8058);
nor U8302 (N_8302,N_8139,N_8164);
nor U8303 (N_8303,N_8105,N_8011);
or U8304 (N_8304,N_8059,N_8090);
or U8305 (N_8305,N_8102,N_8188);
and U8306 (N_8306,N_8147,N_8143);
or U8307 (N_8307,N_8198,N_8056);
nor U8308 (N_8308,N_8148,N_8137);
nand U8309 (N_8309,N_8066,N_8121);
or U8310 (N_8310,N_8048,N_8176);
nand U8311 (N_8311,N_8013,N_8187);
nand U8312 (N_8312,N_8072,N_8089);
nor U8313 (N_8313,N_8051,N_8009);
and U8314 (N_8314,N_8028,N_8033);
or U8315 (N_8315,N_8083,N_8164);
or U8316 (N_8316,N_8148,N_8005);
or U8317 (N_8317,N_8088,N_8145);
nor U8318 (N_8318,N_8016,N_8041);
or U8319 (N_8319,N_8106,N_8127);
or U8320 (N_8320,N_8146,N_8058);
nand U8321 (N_8321,N_8031,N_8092);
or U8322 (N_8322,N_8139,N_8052);
nand U8323 (N_8323,N_8073,N_8119);
nand U8324 (N_8324,N_8149,N_8152);
nand U8325 (N_8325,N_8036,N_8075);
nand U8326 (N_8326,N_8116,N_8077);
and U8327 (N_8327,N_8026,N_8190);
nand U8328 (N_8328,N_8062,N_8171);
nor U8329 (N_8329,N_8104,N_8038);
and U8330 (N_8330,N_8009,N_8085);
and U8331 (N_8331,N_8029,N_8001);
nor U8332 (N_8332,N_8152,N_8114);
nand U8333 (N_8333,N_8023,N_8079);
nand U8334 (N_8334,N_8149,N_8062);
nor U8335 (N_8335,N_8104,N_8168);
nor U8336 (N_8336,N_8139,N_8083);
or U8337 (N_8337,N_8005,N_8093);
nand U8338 (N_8338,N_8076,N_8038);
and U8339 (N_8339,N_8143,N_8113);
nand U8340 (N_8340,N_8045,N_8011);
xor U8341 (N_8341,N_8083,N_8076);
nor U8342 (N_8342,N_8144,N_8037);
xnor U8343 (N_8343,N_8191,N_8123);
nand U8344 (N_8344,N_8063,N_8188);
or U8345 (N_8345,N_8068,N_8037);
or U8346 (N_8346,N_8164,N_8082);
or U8347 (N_8347,N_8057,N_8058);
nand U8348 (N_8348,N_8189,N_8090);
or U8349 (N_8349,N_8020,N_8130);
nand U8350 (N_8350,N_8091,N_8043);
nand U8351 (N_8351,N_8027,N_8072);
and U8352 (N_8352,N_8048,N_8047);
xnor U8353 (N_8353,N_8099,N_8068);
xnor U8354 (N_8354,N_8033,N_8133);
or U8355 (N_8355,N_8106,N_8050);
or U8356 (N_8356,N_8114,N_8135);
nand U8357 (N_8357,N_8129,N_8139);
and U8358 (N_8358,N_8108,N_8050);
nand U8359 (N_8359,N_8042,N_8140);
nor U8360 (N_8360,N_8143,N_8015);
and U8361 (N_8361,N_8103,N_8191);
nand U8362 (N_8362,N_8004,N_8053);
nand U8363 (N_8363,N_8191,N_8197);
nor U8364 (N_8364,N_8062,N_8086);
nand U8365 (N_8365,N_8050,N_8139);
and U8366 (N_8366,N_8145,N_8021);
nor U8367 (N_8367,N_8086,N_8118);
nand U8368 (N_8368,N_8105,N_8012);
nand U8369 (N_8369,N_8171,N_8074);
or U8370 (N_8370,N_8139,N_8008);
and U8371 (N_8371,N_8181,N_8139);
nand U8372 (N_8372,N_8158,N_8146);
and U8373 (N_8373,N_8157,N_8192);
nor U8374 (N_8374,N_8120,N_8186);
nor U8375 (N_8375,N_8110,N_8101);
and U8376 (N_8376,N_8174,N_8177);
nand U8377 (N_8377,N_8089,N_8179);
nor U8378 (N_8378,N_8041,N_8049);
nand U8379 (N_8379,N_8004,N_8035);
and U8380 (N_8380,N_8177,N_8089);
nor U8381 (N_8381,N_8110,N_8040);
nand U8382 (N_8382,N_8142,N_8133);
and U8383 (N_8383,N_8071,N_8089);
or U8384 (N_8384,N_8181,N_8186);
and U8385 (N_8385,N_8166,N_8052);
or U8386 (N_8386,N_8154,N_8171);
nor U8387 (N_8387,N_8116,N_8165);
nor U8388 (N_8388,N_8170,N_8126);
nand U8389 (N_8389,N_8039,N_8075);
or U8390 (N_8390,N_8061,N_8157);
nor U8391 (N_8391,N_8056,N_8153);
nand U8392 (N_8392,N_8025,N_8070);
or U8393 (N_8393,N_8148,N_8057);
nor U8394 (N_8394,N_8070,N_8113);
or U8395 (N_8395,N_8019,N_8076);
and U8396 (N_8396,N_8040,N_8011);
and U8397 (N_8397,N_8070,N_8111);
nor U8398 (N_8398,N_8122,N_8033);
or U8399 (N_8399,N_8046,N_8014);
nand U8400 (N_8400,N_8223,N_8277);
and U8401 (N_8401,N_8398,N_8320);
nand U8402 (N_8402,N_8292,N_8299);
and U8403 (N_8403,N_8388,N_8366);
and U8404 (N_8404,N_8318,N_8250);
or U8405 (N_8405,N_8236,N_8367);
nor U8406 (N_8406,N_8317,N_8343);
nor U8407 (N_8407,N_8330,N_8247);
or U8408 (N_8408,N_8363,N_8322);
and U8409 (N_8409,N_8259,N_8339);
or U8410 (N_8410,N_8238,N_8224);
nand U8411 (N_8411,N_8387,N_8204);
nand U8412 (N_8412,N_8389,N_8270);
nand U8413 (N_8413,N_8274,N_8218);
and U8414 (N_8414,N_8346,N_8258);
or U8415 (N_8415,N_8289,N_8329);
and U8416 (N_8416,N_8311,N_8231);
nand U8417 (N_8417,N_8206,N_8337);
nand U8418 (N_8418,N_8378,N_8350);
and U8419 (N_8419,N_8371,N_8243);
nand U8420 (N_8420,N_8385,N_8272);
nor U8421 (N_8421,N_8280,N_8278);
and U8422 (N_8422,N_8240,N_8351);
or U8423 (N_8423,N_8325,N_8319);
nor U8424 (N_8424,N_8365,N_8281);
or U8425 (N_8425,N_8241,N_8205);
or U8426 (N_8426,N_8390,N_8321);
nor U8427 (N_8427,N_8324,N_8380);
nor U8428 (N_8428,N_8239,N_8296);
nor U8429 (N_8429,N_8225,N_8227);
or U8430 (N_8430,N_8235,N_8370);
nand U8431 (N_8431,N_8384,N_8354);
and U8432 (N_8432,N_8298,N_8248);
and U8433 (N_8433,N_8294,N_8356);
or U8434 (N_8434,N_8251,N_8300);
nor U8435 (N_8435,N_8359,N_8266);
nand U8436 (N_8436,N_8207,N_8364);
xor U8437 (N_8437,N_8312,N_8349);
nand U8438 (N_8438,N_8373,N_8328);
or U8439 (N_8439,N_8357,N_8233);
nor U8440 (N_8440,N_8263,N_8210);
nor U8441 (N_8441,N_8301,N_8331);
or U8442 (N_8442,N_8309,N_8372);
nand U8443 (N_8443,N_8336,N_8276);
and U8444 (N_8444,N_8334,N_8392);
or U8445 (N_8445,N_8382,N_8262);
nor U8446 (N_8446,N_8313,N_8374);
or U8447 (N_8447,N_8244,N_8308);
nand U8448 (N_8448,N_8303,N_8326);
nand U8449 (N_8449,N_8215,N_8291);
or U8450 (N_8450,N_8302,N_8232);
nor U8451 (N_8451,N_8341,N_8253);
nand U8452 (N_8452,N_8310,N_8249);
nand U8453 (N_8453,N_8315,N_8216);
nor U8454 (N_8454,N_8245,N_8369);
or U8455 (N_8455,N_8344,N_8273);
nand U8456 (N_8456,N_8304,N_8201);
nand U8457 (N_8457,N_8285,N_8267);
and U8458 (N_8458,N_8255,N_8217);
or U8459 (N_8459,N_8284,N_8338);
or U8460 (N_8460,N_8348,N_8265);
or U8461 (N_8461,N_8282,N_8316);
nor U8462 (N_8462,N_8360,N_8202);
nor U8463 (N_8463,N_8230,N_8213);
nor U8464 (N_8464,N_8261,N_8226);
and U8465 (N_8465,N_8288,N_8305);
or U8466 (N_8466,N_8394,N_8333);
or U8467 (N_8467,N_8286,N_8393);
or U8468 (N_8468,N_8375,N_8347);
nand U8469 (N_8469,N_8327,N_8229);
or U8470 (N_8470,N_8295,N_8275);
or U8471 (N_8471,N_8377,N_8264);
or U8472 (N_8472,N_8256,N_8212);
or U8473 (N_8473,N_8342,N_8391);
nor U8474 (N_8474,N_8221,N_8297);
nor U8475 (N_8475,N_8345,N_8376);
or U8476 (N_8476,N_8283,N_8368);
nand U8477 (N_8477,N_8386,N_8381);
and U8478 (N_8478,N_8361,N_8332);
nor U8479 (N_8479,N_8246,N_8355);
and U8480 (N_8480,N_8234,N_8257);
nor U8481 (N_8481,N_8395,N_8252);
and U8482 (N_8482,N_8287,N_8314);
or U8483 (N_8483,N_8242,N_8379);
and U8484 (N_8484,N_8269,N_8219);
nor U8485 (N_8485,N_8323,N_8200);
nand U8486 (N_8486,N_8306,N_8220);
nor U8487 (N_8487,N_8293,N_8211);
and U8488 (N_8488,N_8397,N_8399);
or U8489 (N_8489,N_8222,N_8214);
nor U8490 (N_8490,N_8203,N_8352);
and U8491 (N_8491,N_8208,N_8362);
nor U8492 (N_8492,N_8271,N_8340);
and U8493 (N_8493,N_8268,N_8335);
nor U8494 (N_8494,N_8228,N_8358);
nor U8495 (N_8495,N_8237,N_8279);
nor U8496 (N_8496,N_8307,N_8396);
or U8497 (N_8497,N_8383,N_8260);
or U8498 (N_8498,N_8290,N_8209);
or U8499 (N_8499,N_8254,N_8353);
nand U8500 (N_8500,N_8383,N_8362);
nor U8501 (N_8501,N_8281,N_8341);
and U8502 (N_8502,N_8329,N_8239);
nor U8503 (N_8503,N_8386,N_8336);
nor U8504 (N_8504,N_8325,N_8285);
nor U8505 (N_8505,N_8239,N_8260);
or U8506 (N_8506,N_8326,N_8391);
nor U8507 (N_8507,N_8258,N_8325);
or U8508 (N_8508,N_8217,N_8395);
or U8509 (N_8509,N_8212,N_8347);
nor U8510 (N_8510,N_8338,N_8368);
or U8511 (N_8511,N_8328,N_8343);
nand U8512 (N_8512,N_8290,N_8334);
xnor U8513 (N_8513,N_8215,N_8284);
xor U8514 (N_8514,N_8277,N_8263);
nor U8515 (N_8515,N_8345,N_8358);
or U8516 (N_8516,N_8208,N_8209);
or U8517 (N_8517,N_8361,N_8255);
and U8518 (N_8518,N_8262,N_8274);
nor U8519 (N_8519,N_8320,N_8267);
nand U8520 (N_8520,N_8310,N_8303);
nand U8521 (N_8521,N_8221,N_8397);
nand U8522 (N_8522,N_8301,N_8338);
or U8523 (N_8523,N_8374,N_8272);
and U8524 (N_8524,N_8389,N_8269);
and U8525 (N_8525,N_8245,N_8283);
or U8526 (N_8526,N_8219,N_8342);
nor U8527 (N_8527,N_8241,N_8249);
nor U8528 (N_8528,N_8211,N_8202);
or U8529 (N_8529,N_8347,N_8323);
nor U8530 (N_8530,N_8257,N_8200);
or U8531 (N_8531,N_8311,N_8284);
nand U8532 (N_8532,N_8253,N_8254);
nor U8533 (N_8533,N_8300,N_8385);
or U8534 (N_8534,N_8327,N_8346);
or U8535 (N_8535,N_8387,N_8367);
or U8536 (N_8536,N_8316,N_8213);
nand U8537 (N_8537,N_8303,N_8377);
and U8538 (N_8538,N_8306,N_8334);
nor U8539 (N_8539,N_8383,N_8216);
nor U8540 (N_8540,N_8210,N_8317);
nor U8541 (N_8541,N_8369,N_8258);
nor U8542 (N_8542,N_8249,N_8205);
or U8543 (N_8543,N_8378,N_8289);
nor U8544 (N_8544,N_8321,N_8237);
or U8545 (N_8545,N_8373,N_8209);
nand U8546 (N_8546,N_8321,N_8286);
or U8547 (N_8547,N_8209,N_8232);
nor U8548 (N_8548,N_8344,N_8260);
and U8549 (N_8549,N_8371,N_8397);
nand U8550 (N_8550,N_8343,N_8371);
or U8551 (N_8551,N_8275,N_8348);
or U8552 (N_8552,N_8302,N_8333);
nor U8553 (N_8553,N_8372,N_8267);
or U8554 (N_8554,N_8356,N_8276);
xnor U8555 (N_8555,N_8259,N_8376);
xnor U8556 (N_8556,N_8341,N_8324);
nor U8557 (N_8557,N_8278,N_8200);
nand U8558 (N_8558,N_8367,N_8259);
xnor U8559 (N_8559,N_8247,N_8378);
and U8560 (N_8560,N_8369,N_8241);
nor U8561 (N_8561,N_8326,N_8213);
nor U8562 (N_8562,N_8252,N_8318);
nand U8563 (N_8563,N_8300,N_8250);
nor U8564 (N_8564,N_8376,N_8352);
and U8565 (N_8565,N_8333,N_8331);
or U8566 (N_8566,N_8201,N_8212);
nor U8567 (N_8567,N_8290,N_8202);
and U8568 (N_8568,N_8243,N_8378);
nor U8569 (N_8569,N_8204,N_8356);
nor U8570 (N_8570,N_8279,N_8317);
and U8571 (N_8571,N_8345,N_8208);
nor U8572 (N_8572,N_8235,N_8272);
nor U8573 (N_8573,N_8278,N_8396);
nand U8574 (N_8574,N_8356,N_8285);
and U8575 (N_8575,N_8215,N_8395);
or U8576 (N_8576,N_8289,N_8217);
nand U8577 (N_8577,N_8293,N_8298);
nor U8578 (N_8578,N_8266,N_8398);
and U8579 (N_8579,N_8229,N_8243);
and U8580 (N_8580,N_8274,N_8304);
and U8581 (N_8581,N_8369,N_8250);
nor U8582 (N_8582,N_8390,N_8245);
and U8583 (N_8583,N_8337,N_8372);
and U8584 (N_8584,N_8318,N_8325);
nor U8585 (N_8585,N_8250,N_8371);
or U8586 (N_8586,N_8271,N_8236);
and U8587 (N_8587,N_8224,N_8292);
or U8588 (N_8588,N_8317,N_8212);
xor U8589 (N_8589,N_8321,N_8342);
and U8590 (N_8590,N_8234,N_8264);
and U8591 (N_8591,N_8386,N_8200);
and U8592 (N_8592,N_8387,N_8229);
nor U8593 (N_8593,N_8343,N_8334);
and U8594 (N_8594,N_8241,N_8263);
and U8595 (N_8595,N_8293,N_8332);
nand U8596 (N_8596,N_8219,N_8353);
nor U8597 (N_8597,N_8260,N_8274);
nand U8598 (N_8598,N_8231,N_8366);
xor U8599 (N_8599,N_8210,N_8369);
or U8600 (N_8600,N_8556,N_8428);
or U8601 (N_8601,N_8567,N_8485);
or U8602 (N_8602,N_8580,N_8586);
or U8603 (N_8603,N_8588,N_8450);
or U8604 (N_8604,N_8599,N_8577);
nand U8605 (N_8605,N_8405,N_8597);
nand U8606 (N_8606,N_8499,N_8593);
nor U8607 (N_8607,N_8458,N_8560);
nand U8608 (N_8608,N_8594,N_8420);
or U8609 (N_8609,N_8406,N_8557);
xor U8610 (N_8610,N_8595,N_8472);
nand U8611 (N_8611,N_8473,N_8494);
and U8612 (N_8612,N_8486,N_8481);
and U8613 (N_8613,N_8585,N_8554);
and U8614 (N_8614,N_8546,N_8497);
nand U8615 (N_8615,N_8407,N_8598);
nand U8616 (N_8616,N_8455,N_8492);
or U8617 (N_8617,N_8456,N_8482);
or U8618 (N_8618,N_8442,N_8570);
or U8619 (N_8619,N_8489,N_8477);
or U8620 (N_8620,N_8464,N_8581);
and U8621 (N_8621,N_8490,N_8511);
nor U8622 (N_8622,N_8507,N_8518);
nand U8623 (N_8623,N_8596,N_8487);
and U8624 (N_8624,N_8475,N_8572);
nor U8625 (N_8625,N_8539,N_8467);
or U8626 (N_8626,N_8545,N_8509);
and U8627 (N_8627,N_8532,N_8548);
nor U8628 (N_8628,N_8402,N_8410);
nor U8629 (N_8629,N_8495,N_8404);
nor U8630 (N_8630,N_8483,N_8504);
nor U8631 (N_8631,N_8535,N_8491);
nor U8632 (N_8632,N_8441,N_8538);
or U8633 (N_8633,N_8564,N_8445);
nor U8634 (N_8634,N_8496,N_8421);
or U8635 (N_8635,N_8531,N_8503);
nand U8636 (N_8636,N_8505,N_8500);
nor U8637 (N_8637,N_8444,N_8448);
and U8638 (N_8638,N_8521,N_8573);
nor U8639 (N_8639,N_8578,N_8543);
nand U8640 (N_8640,N_8575,N_8431);
or U8641 (N_8641,N_8529,N_8547);
nor U8642 (N_8642,N_8435,N_8468);
nor U8643 (N_8643,N_8436,N_8424);
nor U8644 (N_8644,N_8540,N_8584);
nand U8645 (N_8645,N_8403,N_8466);
nand U8646 (N_8646,N_8517,N_8569);
nand U8647 (N_8647,N_8592,N_8443);
nor U8648 (N_8648,N_8488,N_8550);
nand U8649 (N_8649,N_8558,N_8457);
and U8650 (N_8650,N_8512,N_8426);
or U8651 (N_8651,N_8549,N_8544);
or U8652 (N_8652,N_8565,N_8498);
and U8653 (N_8653,N_8536,N_8527);
nand U8654 (N_8654,N_8419,N_8510);
or U8655 (N_8655,N_8479,N_8566);
nor U8656 (N_8656,N_8414,N_8542);
nand U8657 (N_8657,N_8551,N_8552);
nand U8658 (N_8658,N_8415,N_8528);
or U8659 (N_8659,N_8590,N_8462);
nor U8660 (N_8660,N_8541,N_8454);
nand U8661 (N_8661,N_8422,N_8568);
and U8662 (N_8662,N_8587,N_8471);
nand U8663 (N_8663,N_8523,N_8520);
nor U8664 (N_8664,N_8461,N_8478);
and U8665 (N_8665,N_8574,N_8537);
and U8666 (N_8666,N_8484,N_8408);
and U8667 (N_8667,N_8401,N_8591);
nor U8668 (N_8668,N_8513,N_8579);
nand U8669 (N_8669,N_8463,N_8576);
or U8670 (N_8670,N_8519,N_8525);
and U8671 (N_8671,N_8418,N_8559);
or U8672 (N_8672,N_8449,N_8508);
nand U8673 (N_8673,N_8516,N_8480);
and U8674 (N_8674,N_8476,N_8400);
nor U8675 (N_8675,N_8526,N_8515);
and U8676 (N_8676,N_8493,N_8583);
nand U8677 (N_8677,N_8553,N_8502);
nand U8678 (N_8678,N_8453,N_8474);
and U8679 (N_8679,N_8562,N_8530);
nor U8680 (N_8680,N_8465,N_8412);
or U8681 (N_8681,N_8429,N_8430);
nor U8682 (N_8682,N_8439,N_8459);
or U8683 (N_8683,N_8582,N_8411);
and U8684 (N_8684,N_8524,N_8409);
nor U8685 (N_8685,N_8423,N_8425);
and U8686 (N_8686,N_8433,N_8452);
nand U8687 (N_8687,N_8416,N_8501);
and U8688 (N_8688,N_8563,N_8534);
and U8689 (N_8689,N_8447,N_8434);
nand U8690 (N_8690,N_8470,N_8555);
or U8691 (N_8691,N_8413,N_8460);
nand U8692 (N_8692,N_8446,N_8506);
and U8693 (N_8693,N_8427,N_8561);
nor U8694 (N_8694,N_8440,N_8522);
nor U8695 (N_8695,N_8589,N_8451);
or U8696 (N_8696,N_8437,N_8514);
nand U8697 (N_8697,N_8533,N_8438);
nand U8698 (N_8698,N_8432,N_8469);
and U8699 (N_8699,N_8417,N_8571);
or U8700 (N_8700,N_8502,N_8498);
nand U8701 (N_8701,N_8527,N_8494);
nor U8702 (N_8702,N_8421,N_8536);
nor U8703 (N_8703,N_8574,N_8509);
and U8704 (N_8704,N_8451,N_8427);
and U8705 (N_8705,N_8528,N_8456);
nor U8706 (N_8706,N_8569,N_8449);
nor U8707 (N_8707,N_8418,N_8406);
nor U8708 (N_8708,N_8417,N_8548);
or U8709 (N_8709,N_8422,N_8428);
and U8710 (N_8710,N_8452,N_8549);
nor U8711 (N_8711,N_8529,N_8446);
nand U8712 (N_8712,N_8518,N_8465);
nand U8713 (N_8713,N_8532,N_8523);
and U8714 (N_8714,N_8425,N_8426);
xnor U8715 (N_8715,N_8448,N_8541);
or U8716 (N_8716,N_8407,N_8569);
and U8717 (N_8717,N_8527,N_8414);
or U8718 (N_8718,N_8524,N_8488);
or U8719 (N_8719,N_8481,N_8571);
nand U8720 (N_8720,N_8512,N_8427);
or U8721 (N_8721,N_8400,N_8404);
or U8722 (N_8722,N_8490,N_8575);
nor U8723 (N_8723,N_8461,N_8422);
nand U8724 (N_8724,N_8454,N_8536);
and U8725 (N_8725,N_8431,N_8428);
nand U8726 (N_8726,N_8462,N_8419);
nor U8727 (N_8727,N_8514,N_8423);
and U8728 (N_8728,N_8497,N_8430);
and U8729 (N_8729,N_8580,N_8566);
or U8730 (N_8730,N_8596,N_8411);
nor U8731 (N_8731,N_8494,N_8479);
nor U8732 (N_8732,N_8423,N_8557);
or U8733 (N_8733,N_8508,N_8477);
nand U8734 (N_8734,N_8536,N_8444);
nor U8735 (N_8735,N_8542,N_8503);
or U8736 (N_8736,N_8518,N_8407);
nor U8737 (N_8737,N_8592,N_8426);
or U8738 (N_8738,N_8566,N_8405);
or U8739 (N_8739,N_8584,N_8585);
nand U8740 (N_8740,N_8581,N_8473);
and U8741 (N_8741,N_8463,N_8560);
nor U8742 (N_8742,N_8510,N_8453);
nor U8743 (N_8743,N_8483,N_8573);
and U8744 (N_8744,N_8500,N_8462);
and U8745 (N_8745,N_8520,N_8403);
and U8746 (N_8746,N_8419,N_8585);
or U8747 (N_8747,N_8490,N_8438);
or U8748 (N_8748,N_8424,N_8465);
nand U8749 (N_8749,N_8587,N_8449);
or U8750 (N_8750,N_8489,N_8555);
nor U8751 (N_8751,N_8511,N_8485);
and U8752 (N_8752,N_8410,N_8443);
nor U8753 (N_8753,N_8539,N_8466);
nor U8754 (N_8754,N_8511,N_8595);
nor U8755 (N_8755,N_8497,N_8515);
nand U8756 (N_8756,N_8522,N_8447);
nor U8757 (N_8757,N_8493,N_8507);
nor U8758 (N_8758,N_8560,N_8598);
or U8759 (N_8759,N_8514,N_8479);
nor U8760 (N_8760,N_8559,N_8454);
and U8761 (N_8761,N_8545,N_8505);
nor U8762 (N_8762,N_8540,N_8517);
and U8763 (N_8763,N_8533,N_8432);
nand U8764 (N_8764,N_8501,N_8484);
or U8765 (N_8765,N_8502,N_8507);
nor U8766 (N_8766,N_8581,N_8449);
nand U8767 (N_8767,N_8575,N_8531);
nand U8768 (N_8768,N_8519,N_8530);
nand U8769 (N_8769,N_8576,N_8456);
and U8770 (N_8770,N_8529,N_8544);
or U8771 (N_8771,N_8551,N_8567);
or U8772 (N_8772,N_8589,N_8417);
xor U8773 (N_8773,N_8421,N_8454);
nor U8774 (N_8774,N_8404,N_8552);
or U8775 (N_8775,N_8439,N_8534);
and U8776 (N_8776,N_8521,N_8552);
nor U8777 (N_8777,N_8546,N_8597);
or U8778 (N_8778,N_8528,N_8507);
and U8779 (N_8779,N_8485,N_8473);
nand U8780 (N_8780,N_8422,N_8510);
nor U8781 (N_8781,N_8408,N_8464);
nand U8782 (N_8782,N_8457,N_8544);
nor U8783 (N_8783,N_8475,N_8576);
nand U8784 (N_8784,N_8560,N_8547);
nand U8785 (N_8785,N_8599,N_8570);
nand U8786 (N_8786,N_8537,N_8509);
or U8787 (N_8787,N_8451,N_8493);
and U8788 (N_8788,N_8411,N_8529);
and U8789 (N_8789,N_8579,N_8452);
and U8790 (N_8790,N_8433,N_8521);
and U8791 (N_8791,N_8563,N_8506);
and U8792 (N_8792,N_8462,N_8472);
or U8793 (N_8793,N_8509,N_8570);
nor U8794 (N_8794,N_8411,N_8425);
and U8795 (N_8795,N_8500,N_8461);
or U8796 (N_8796,N_8401,N_8534);
or U8797 (N_8797,N_8404,N_8511);
or U8798 (N_8798,N_8536,N_8409);
or U8799 (N_8799,N_8481,N_8455);
nand U8800 (N_8800,N_8741,N_8780);
nor U8801 (N_8801,N_8688,N_8687);
and U8802 (N_8802,N_8743,N_8718);
or U8803 (N_8803,N_8632,N_8785);
and U8804 (N_8804,N_8639,N_8710);
nor U8805 (N_8805,N_8626,N_8774);
and U8806 (N_8806,N_8674,N_8649);
and U8807 (N_8807,N_8647,N_8735);
or U8808 (N_8808,N_8650,N_8756);
nand U8809 (N_8809,N_8662,N_8724);
or U8810 (N_8810,N_8702,N_8779);
and U8811 (N_8811,N_8704,N_8744);
or U8812 (N_8812,N_8624,N_8675);
xor U8813 (N_8813,N_8748,N_8792);
nand U8814 (N_8814,N_8691,N_8602);
nand U8815 (N_8815,N_8765,N_8752);
nor U8816 (N_8816,N_8750,N_8689);
nand U8817 (N_8817,N_8660,N_8726);
nor U8818 (N_8818,N_8755,N_8673);
nand U8819 (N_8819,N_8793,N_8746);
nand U8820 (N_8820,N_8676,N_8708);
and U8821 (N_8821,N_8606,N_8664);
nand U8822 (N_8822,N_8628,N_8754);
nand U8823 (N_8823,N_8728,N_8715);
xnor U8824 (N_8824,N_8607,N_8737);
nor U8825 (N_8825,N_8617,N_8681);
nor U8826 (N_8826,N_8643,N_8663);
nand U8827 (N_8827,N_8712,N_8731);
or U8828 (N_8828,N_8751,N_8781);
nor U8829 (N_8829,N_8618,N_8783);
or U8830 (N_8830,N_8727,N_8686);
and U8831 (N_8831,N_8763,N_8776);
and U8832 (N_8832,N_8659,N_8740);
nor U8833 (N_8833,N_8625,N_8680);
nor U8834 (N_8834,N_8622,N_8711);
nand U8835 (N_8835,N_8614,N_8690);
xor U8836 (N_8836,N_8729,N_8609);
nand U8837 (N_8837,N_8794,N_8720);
nand U8838 (N_8838,N_8600,N_8719);
or U8839 (N_8839,N_8697,N_8788);
and U8840 (N_8840,N_8767,N_8653);
nor U8841 (N_8841,N_8722,N_8616);
and U8842 (N_8842,N_8782,N_8739);
nand U8843 (N_8843,N_8668,N_8766);
or U8844 (N_8844,N_8636,N_8642);
or U8845 (N_8845,N_8667,N_8613);
nand U8846 (N_8846,N_8623,N_8683);
and U8847 (N_8847,N_8665,N_8631);
nor U8848 (N_8848,N_8634,N_8648);
and U8849 (N_8849,N_8682,N_8661);
and U8850 (N_8850,N_8797,N_8699);
nand U8851 (N_8851,N_8714,N_8604);
nand U8852 (N_8852,N_8758,N_8684);
xnor U8853 (N_8853,N_8620,N_8685);
nor U8854 (N_8854,N_8700,N_8799);
nand U8855 (N_8855,N_8753,N_8723);
and U8856 (N_8856,N_8656,N_8669);
nand U8857 (N_8857,N_8627,N_8645);
or U8858 (N_8858,N_8693,N_8610);
and U8859 (N_8859,N_8694,N_8789);
or U8860 (N_8860,N_8621,N_8764);
nand U8861 (N_8861,N_8678,N_8601);
nor U8862 (N_8862,N_8725,N_8679);
and U8863 (N_8863,N_8701,N_8612);
nor U8864 (N_8864,N_8611,N_8760);
or U8865 (N_8865,N_8773,N_8732);
or U8866 (N_8866,N_8745,N_8705);
or U8867 (N_8867,N_8778,N_8658);
nand U8868 (N_8868,N_8670,N_8641);
or U8869 (N_8869,N_8777,N_8768);
nor U8870 (N_8870,N_8757,N_8698);
nor U8871 (N_8871,N_8784,N_8619);
nor U8872 (N_8872,N_8646,N_8605);
or U8873 (N_8873,N_8798,N_8791);
or U8874 (N_8874,N_8706,N_8721);
nand U8875 (N_8875,N_8703,N_8787);
nor U8876 (N_8876,N_8672,N_8652);
nor U8877 (N_8877,N_8654,N_8738);
nand U8878 (N_8878,N_8759,N_8769);
xnor U8879 (N_8879,N_8651,N_8695);
and U8880 (N_8880,N_8709,N_8742);
and U8881 (N_8881,N_8657,N_8644);
or U8882 (N_8882,N_8630,N_8635);
nor U8883 (N_8883,N_8655,N_8638);
xnor U8884 (N_8884,N_8696,N_8747);
and U8885 (N_8885,N_8749,N_8671);
nand U8886 (N_8886,N_8713,N_8603);
xnor U8887 (N_8887,N_8796,N_8771);
and U8888 (N_8888,N_8707,N_8629);
nand U8889 (N_8889,N_8730,N_8716);
nor U8890 (N_8890,N_8666,N_8733);
nor U8891 (N_8891,N_8790,N_8786);
nor U8892 (N_8892,N_8795,N_8608);
nor U8893 (N_8893,N_8736,N_8615);
nor U8894 (N_8894,N_8692,N_8772);
nand U8895 (N_8895,N_8717,N_8633);
nand U8896 (N_8896,N_8734,N_8775);
nor U8897 (N_8897,N_8677,N_8761);
or U8898 (N_8898,N_8762,N_8770);
nor U8899 (N_8899,N_8637,N_8640);
or U8900 (N_8900,N_8704,N_8721);
nand U8901 (N_8901,N_8667,N_8648);
or U8902 (N_8902,N_8614,N_8629);
xnor U8903 (N_8903,N_8756,N_8753);
or U8904 (N_8904,N_8671,N_8665);
nand U8905 (N_8905,N_8729,N_8735);
or U8906 (N_8906,N_8709,N_8697);
and U8907 (N_8907,N_8632,N_8735);
or U8908 (N_8908,N_8619,N_8666);
and U8909 (N_8909,N_8638,N_8699);
or U8910 (N_8910,N_8692,N_8687);
nor U8911 (N_8911,N_8608,N_8600);
or U8912 (N_8912,N_8668,N_8779);
nand U8913 (N_8913,N_8641,N_8613);
or U8914 (N_8914,N_8660,N_8655);
xnor U8915 (N_8915,N_8681,N_8762);
nor U8916 (N_8916,N_8781,N_8694);
nand U8917 (N_8917,N_8691,N_8657);
or U8918 (N_8918,N_8658,N_8794);
nand U8919 (N_8919,N_8727,N_8648);
and U8920 (N_8920,N_8618,N_8660);
nand U8921 (N_8921,N_8667,N_8682);
nand U8922 (N_8922,N_8674,N_8684);
and U8923 (N_8923,N_8604,N_8638);
nor U8924 (N_8924,N_8745,N_8702);
or U8925 (N_8925,N_8687,N_8713);
nor U8926 (N_8926,N_8610,N_8736);
nand U8927 (N_8927,N_8656,N_8714);
or U8928 (N_8928,N_8769,N_8770);
or U8929 (N_8929,N_8621,N_8685);
nor U8930 (N_8930,N_8614,N_8713);
nand U8931 (N_8931,N_8621,N_8700);
or U8932 (N_8932,N_8675,N_8797);
or U8933 (N_8933,N_8742,N_8761);
or U8934 (N_8934,N_8756,N_8667);
nor U8935 (N_8935,N_8756,N_8653);
nand U8936 (N_8936,N_8643,N_8684);
xor U8937 (N_8937,N_8788,N_8620);
nor U8938 (N_8938,N_8716,N_8775);
or U8939 (N_8939,N_8785,N_8617);
xnor U8940 (N_8940,N_8755,N_8780);
or U8941 (N_8941,N_8681,N_8730);
nor U8942 (N_8942,N_8788,N_8682);
nor U8943 (N_8943,N_8766,N_8667);
nor U8944 (N_8944,N_8672,N_8697);
nand U8945 (N_8945,N_8672,N_8701);
nor U8946 (N_8946,N_8736,N_8777);
or U8947 (N_8947,N_8671,N_8766);
nor U8948 (N_8948,N_8618,N_8706);
nand U8949 (N_8949,N_8790,N_8774);
and U8950 (N_8950,N_8663,N_8622);
or U8951 (N_8951,N_8756,N_8725);
or U8952 (N_8952,N_8749,N_8753);
and U8953 (N_8953,N_8681,N_8717);
and U8954 (N_8954,N_8619,N_8706);
or U8955 (N_8955,N_8798,N_8785);
nand U8956 (N_8956,N_8710,N_8600);
and U8957 (N_8957,N_8619,N_8690);
or U8958 (N_8958,N_8756,N_8733);
and U8959 (N_8959,N_8706,N_8676);
nand U8960 (N_8960,N_8616,N_8799);
or U8961 (N_8961,N_8636,N_8673);
and U8962 (N_8962,N_8739,N_8757);
nor U8963 (N_8963,N_8624,N_8780);
or U8964 (N_8964,N_8605,N_8798);
and U8965 (N_8965,N_8774,N_8605);
or U8966 (N_8966,N_8769,N_8603);
or U8967 (N_8967,N_8669,N_8771);
xnor U8968 (N_8968,N_8740,N_8614);
and U8969 (N_8969,N_8765,N_8727);
nor U8970 (N_8970,N_8611,N_8722);
and U8971 (N_8971,N_8607,N_8621);
nand U8972 (N_8972,N_8762,N_8767);
and U8973 (N_8973,N_8713,N_8628);
nor U8974 (N_8974,N_8621,N_8684);
or U8975 (N_8975,N_8674,N_8781);
nand U8976 (N_8976,N_8793,N_8785);
and U8977 (N_8977,N_8704,N_8688);
or U8978 (N_8978,N_8739,N_8623);
nand U8979 (N_8979,N_8617,N_8604);
or U8980 (N_8980,N_8607,N_8657);
nand U8981 (N_8981,N_8604,N_8716);
nor U8982 (N_8982,N_8619,N_8664);
and U8983 (N_8983,N_8796,N_8669);
nand U8984 (N_8984,N_8727,N_8732);
nor U8985 (N_8985,N_8718,N_8678);
or U8986 (N_8986,N_8666,N_8737);
nor U8987 (N_8987,N_8770,N_8673);
nor U8988 (N_8988,N_8639,N_8793);
or U8989 (N_8989,N_8766,N_8664);
and U8990 (N_8990,N_8736,N_8627);
and U8991 (N_8991,N_8708,N_8652);
nand U8992 (N_8992,N_8767,N_8638);
and U8993 (N_8993,N_8731,N_8720);
and U8994 (N_8994,N_8672,N_8771);
or U8995 (N_8995,N_8689,N_8773);
nor U8996 (N_8996,N_8777,N_8636);
and U8997 (N_8997,N_8771,N_8621);
or U8998 (N_8998,N_8655,N_8746);
or U8999 (N_8999,N_8772,N_8790);
nand U9000 (N_9000,N_8841,N_8993);
nor U9001 (N_9001,N_8970,N_8980);
nand U9002 (N_9002,N_8804,N_8948);
or U9003 (N_9003,N_8937,N_8801);
or U9004 (N_9004,N_8976,N_8820);
nor U9005 (N_9005,N_8928,N_8811);
nor U9006 (N_9006,N_8886,N_8973);
and U9007 (N_9007,N_8918,N_8956);
and U9008 (N_9008,N_8812,N_8895);
nor U9009 (N_9009,N_8942,N_8991);
nor U9010 (N_9010,N_8892,N_8962);
or U9011 (N_9011,N_8999,N_8995);
nor U9012 (N_9012,N_8822,N_8990);
or U9013 (N_9013,N_8908,N_8974);
or U9014 (N_9014,N_8919,N_8836);
or U9015 (N_9015,N_8925,N_8816);
and U9016 (N_9016,N_8959,N_8866);
nor U9017 (N_9017,N_8882,N_8870);
nand U9018 (N_9018,N_8968,N_8874);
or U9019 (N_9019,N_8901,N_8992);
nand U9020 (N_9020,N_8861,N_8864);
and U9021 (N_9021,N_8950,N_8899);
nand U9022 (N_9022,N_8851,N_8808);
and U9023 (N_9023,N_8817,N_8967);
nand U9024 (N_9024,N_8881,N_8979);
xnor U9025 (N_9025,N_8977,N_8885);
and U9026 (N_9026,N_8805,N_8878);
nand U9027 (N_9027,N_8880,N_8989);
and U9028 (N_9028,N_8825,N_8888);
and U9029 (N_9029,N_8807,N_8982);
nand U9030 (N_9030,N_8813,N_8802);
and U9031 (N_9031,N_8868,N_8850);
nand U9032 (N_9032,N_8855,N_8871);
and U9033 (N_9033,N_8815,N_8943);
nand U9034 (N_9034,N_8897,N_8912);
xnor U9035 (N_9035,N_8876,N_8969);
and U9036 (N_9036,N_8883,N_8831);
or U9037 (N_9037,N_8837,N_8852);
nand U9038 (N_9038,N_8997,N_8875);
or U9039 (N_9039,N_8856,N_8862);
and U9040 (N_9040,N_8860,N_8921);
and U9041 (N_9041,N_8954,N_8859);
or U9042 (N_9042,N_8940,N_8915);
or U9043 (N_9043,N_8927,N_8975);
nand U9044 (N_9044,N_8857,N_8909);
and U9045 (N_9045,N_8828,N_8971);
nor U9046 (N_9046,N_8834,N_8939);
nor U9047 (N_9047,N_8947,N_8966);
nand U9048 (N_9048,N_8846,N_8863);
and U9049 (N_9049,N_8934,N_8920);
xnor U9050 (N_9050,N_8889,N_8877);
nand U9051 (N_9051,N_8917,N_8903);
or U9052 (N_9052,N_8938,N_8838);
nor U9053 (N_9053,N_8929,N_8931);
and U9054 (N_9054,N_8945,N_8823);
nor U9055 (N_9055,N_8824,N_8902);
xor U9056 (N_9056,N_8844,N_8910);
and U9057 (N_9057,N_8981,N_8978);
nor U9058 (N_9058,N_8849,N_8935);
or U9059 (N_9059,N_8905,N_8854);
or U9060 (N_9060,N_8869,N_8826);
or U9061 (N_9061,N_8906,N_8930);
nor U9062 (N_9062,N_8964,N_8800);
or U9063 (N_9063,N_8946,N_8996);
and U9064 (N_9064,N_8830,N_8998);
nand U9065 (N_9065,N_8806,N_8893);
xnor U9066 (N_9066,N_8818,N_8933);
and U9067 (N_9067,N_8814,N_8944);
nor U9068 (N_9068,N_8907,N_8847);
and U9069 (N_9069,N_8986,N_8858);
or U9070 (N_9070,N_8941,N_8953);
and U9071 (N_9071,N_8911,N_8809);
nand U9072 (N_9072,N_8924,N_8922);
or U9073 (N_9073,N_8916,N_8865);
nand U9074 (N_9074,N_8960,N_8821);
and U9075 (N_9075,N_8987,N_8972);
xnor U9076 (N_9076,N_8835,N_8872);
nand U9077 (N_9077,N_8949,N_8988);
nor U9078 (N_9078,N_8810,N_8951);
nor U9079 (N_9079,N_8845,N_8884);
and U9080 (N_9080,N_8963,N_8985);
and U9081 (N_9081,N_8879,N_8955);
and U9082 (N_9082,N_8913,N_8848);
or U9083 (N_9083,N_8819,N_8961);
nor U9084 (N_9084,N_8891,N_8914);
and U9085 (N_9085,N_8894,N_8896);
xor U9086 (N_9086,N_8890,N_8952);
nor U9087 (N_9087,N_8873,N_8867);
nor U9088 (N_9088,N_8994,N_8965);
nor U9089 (N_9089,N_8958,N_8829);
or U9090 (N_9090,N_8843,N_8887);
or U9091 (N_9091,N_8842,N_8803);
and U9092 (N_9092,N_8957,N_8900);
and U9093 (N_9093,N_8833,N_8926);
and U9094 (N_9094,N_8832,N_8983);
or U9095 (N_9095,N_8827,N_8839);
nand U9096 (N_9096,N_8853,N_8984);
nor U9097 (N_9097,N_8840,N_8936);
nand U9098 (N_9098,N_8904,N_8932);
nor U9099 (N_9099,N_8898,N_8923);
nand U9100 (N_9100,N_8962,N_8996);
and U9101 (N_9101,N_8962,N_8870);
nor U9102 (N_9102,N_8955,N_8843);
xnor U9103 (N_9103,N_8800,N_8947);
nor U9104 (N_9104,N_8983,N_8988);
nor U9105 (N_9105,N_8856,N_8962);
xnor U9106 (N_9106,N_8852,N_8913);
and U9107 (N_9107,N_8812,N_8821);
nand U9108 (N_9108,N_8830,N_8953);
or U9109 (N_9109,N_8910,N_8911);
nor U9110 (N_9110,N_8935,N_8900);
and U9111 (N_9111,N_8955,N_8903);
nor U9112 (N_9112,N_8866,N_8981);
nor U9113 (N_9113,N_8846,N_8892);
or U9114 (N_9114,N_8857,N_8809);
nand U9115 (N_9115,N_8914,N_8876);
or U9116 (N_9116,N_8874,N_8948);
nand U9117 (N_9117,N_8936,N_8984);
and U9118 (N_9118,N_8820,N_8915);
nor U9119 (N_9119,N_8881,N_8954);
or U9120 (N_9120,N_8849,N_8941);
xor U9121 (N_9121,N_8963,N_8834);
and U9122 (N_9122,N_8915,N_8807);
or U9123 (N_9123,N_8833,N_8891);
nand U9124 (N_9124,N_8937,N_8837);
or U9125 (N_9125,N_8870,N_8975);
nor U9126 (N_9126,N_8993,N_8933);
and U9127 (N_9127,N_8987,N_8973);
nand U9128 (N_9128,N_8899,N_8998);
and U9129 (N_9129,N_8923,N_8999);
or U9130 (N_9130,N_8870,N_8808);
and U9131 (N_9131,N_8870,N_8833);
nor U9132 (N_9132,N_8975,N_8885);
and U9133 (N_9133,N_8876,N_8853);
and U9134 (N_9134,N_8967,N_8873);
nand U9135 (N_9135,N_8938,N_8848);
xor U9136 (N_9136,N_8819,N_8812);
and U9137 (N_9137,N_8840,N_8835);
nor U9138 (N_9138,N_8949,N_8999);
or U9139 (N_9139,N_8835,N_8980);
nor U9140 (N_9140,N_8953,N_8969);
nor U9141 (N_9141,N_8864,N_8986);
or U9142 (N_9142,N_8823,N_8904);
and U9143 (N_9143,N_8848,N_8991);
or U9144 (N_9144,N_8993,N_8966);
and U9145 (N_9145,N_8919,N_8873);
or U9146 (N_9146,N_8963,N_8933);
nand U9147 (N_9147,N_8934,N_8846);
nand U9148 (N_9148,N_8926,N_8966);
or U9149 (N_9149,N_8940,N_8862);
and U9150 (N_9150,N_8992,N_8971);
nor U9151 (N_9151,N_8896,N_8885);
or U9152 (N_9152,N_8963,N_8951);
nor U9153 (N_9153,N_8806,N_8830);
and U9154 (N_9154,N_8981,N_8982);
nand U9155 (N_9155,N_8975,N_8849);
or U9156 (N_9156,N_8934,N_8928);
nand U9157 (N_9157,N_8974,N_8886);
or U9158 (N_9158,N_8996,N_8972);
and U9159 (N_9159,N_8997,N_8854);
or U9160 (N_9160,N_8897,N_8964);
and U9161 (N_9161,N_8842,N_8941);
nor U9162 (N_9162,N_8980,N_8888);
and U9163 (N_9163,N_8860,N_8943);
nand U9164 (N_9164,N_8878,N_8809);
and U9165 (N_9165,N_8855,N_8839);
nor U9166 (N_9166,N_8963,N_8865);
nand U9167 (N_9167,N_8866,N_8882);
and U9168 (N_9168,N_8844,N_8903);
nand U9169 (N_9169,N_8846,N_8830);
nor U9170 (N_9170,N_8956,N_8946);
and U9171 (N_9171,N_8935,N_8844);
nand U9172 (N_9172,N_8843,N_8929);
or U9173 (N_9173,N_8820,N_8917);
and U9174 (N_9174,N_8918,N_8846);
or U9175 (N_9175,N_8902,N_8903);
nor U9176 (N_9176,N_8871,N_8880);
and U9177 (N_9177,N_8908,N_8984);
nand U9178 (N_9178,N_8806,N_8894);
and U9179 (N_9179,N_8853,N_8923);
and U9180 (N_9180,N_8844,N_8800);
or U9181 (N_9181,N_8846,N_8857);
nor U9182 (N_9182,N_8978,N_8922);
or U9183 (N_9183,N_8870,N_8822);
nand U9184 (N_9184,N_8835,N_8903);
nand U9185 (N_9185,N_8915,N_8894);
nand U9186 (N_9186,N_8980,N_8889);
and U9187 (N_9187,N_8928,N_8959);
nand U9188 (N_9188,N_8883,N_8899);
nor U9189 (N_9189,N_8848,N_8823);
or U9190 (N_9190,N_8814,N_8989);
xnor U9191 (N_9191,N_8948,N_8969);
nor U9192 (N_9192,N_8924,N_8916);
nor U9193 (N_9193,N_8864,N_8936);
or U9194 (N_9194,N_8981,N_8892);
nor U9195 (N_9195,N_8940,N_8959);
and U9196 (N_9196,N_8978,N_8874);
or U9197 (N_9197,N_8944,N_8809);
and U9198 (N_9198,N_8817,N_8829);
and U9199 (N_9199,N_8964,N_8884);
nor U9200 (N_9200,N_9005,N_9026);
nor U9201 (N_9201,N_9154,N_9173);
and U9202 (N_9202,N_9188,N_9126);
nor U9203 (N_9203,N_9025,N_9053);
nor U9204 (N_9204,N_9009,N_9054);
and U9205 (N_9205,N_9168,N_9052);
and U9206 (N_9206,N_9020,N_9091);
nor U9207 (N_9207,N_9004,N_9112);
or U9208 (N_9208,N_9031,N_9055);
nor U9209 (N_9209,N_9122,N_9124);
and U9210 (N_9210,N_9043,N_9133);
or U9211 (N_9211,N_9002,N_9199);
or U9212 (N_9212,N_9178,N_9103);
or U9213 (N_9213,N_9129,N_9150);
or U9214 (N_9214,N_9073,N_9061);
and U9215 (N_9215,N_9085,N_9182);
and U9216 (N_9216,N_9138,N_9159);
and U9217 (N_9217,N_9108,N_9177);
or U9218 (N_9218,N_9015,N_9065);
or U9219 (N_9219,N_9058,N_9117);
nand U9220 (N_9220,N_9046,N_9088);
and U9221 (N_9221,N_9139,N_9048);
and U9222 (N_9222,N_9006,N_9111);
and U9223 (N_9223,N_9045,N_9120);
and U9224 (N_9224,N_9060,N_9092);
xor U9225 (N_9225,N_9110,N_9038);
nand U9226 (N_9226,N_9102,N_9194);
or U9227 (N_9227,N_9127,N_9080);
nand U9228 (N_9228,N_9014,N_9049);
or U9229 (N_9229,N_9077,N_9161);
nor U9230 (N_9230,N_9130,N_9185);
nor U9231 (N_9231,N_9074,N_9098);
nor U9232 (N_9232,N_9059,N_9144);
and U9233 (N_9233,N_9198,N_9165);
nor U9234 (N_9234,N_9001,N_9034);
xnor U9235 (N_9235,N_9149,N_9121);
xor U9236 (N_9236,N_9099,N_9036);
or U9237 (N_9237,N_9067,N_9042);
nand U9238 (N_9238,N_9101,N_9145);
and U9239 (N_9239,N_9131,N_9084);
nor U9240 (N_9240,N_9003,N_9094);
and U9241 (N_9241,N_9082,N_9051);
nand U9242 (N_9242,N_9176,N_9013);
nor U9243 (N_9243,N_9100,N_9024);
and U9244 (N_9244,N_9156,N_9057);
nand U9245 (N_9245,N_9000,N_9087);
nand U9246 (N_9246,N_9093,N_9105);
and U9247 (N_9247,N_9187,N_9118);
nand U9248 (N_9248,N_9019,N_9151);
or U9249 (N_9249,N_9070,N_9010);
nor U9250 (N_9250,N_9146,N_9181);
and U9251 (N_9251,N_9134,N_9028);
nor U9252 (N_9252,N_9116,N_9189);
nand U9253 (N_9253,N_9170,N_9090);
nand U9254 (N_9254,N_9160,N_9180);
and U9255 (N_9255,N_9022,N_9172);
nand U9256 (N_9256,N_9029,N_9078);
or U9257 (N_9257,N_9039,N_9135);
and U9258 (N_9258,N_9196,N_9106);
and U9259 (N_9259,N_9197,N_9007);
and U9260 (N_9260,N_9119,N_9179);
xnor U9261 (N_9261,N_9140,N_9018);
and U9262 (N_9262,N_9083,N_9164);
nor U9263 (N_9263,N_9132,N_9183);
xnor U9264 (N_9264,N_9012,N_9066);
or U9265 (N_9265,N_9040,N_9044);
nand U9266 (N_9266,N_9047,N_9153);
or U9267 (N_9267,N_9050,N_9008);
nor U9268 (N_9268,N_9089,N_9192);
or U9269 (N_9269,N_9107,N_9123);
or U9270 (N_9270,N_9104,N_9142);
nor U9271 (N_9271,N_9041,N_9157);
nand U9272 (N_9272,N_9021,N_9075);
nor U9273 (N_9273,N_9023,N_9064);
nand U9274 (N_9274,N_9175,N_9072);
nand U9275 (N_9275,N_9186,N_9136);
xor U9276 (N_9276,N_9033,N_9195);
nor U9277 (N_9277,N_9163,N_9056);
nand U9278 (N_9278,N_9171,N_9086);
xnor U9279 (N_9279,N_9147,N_9069);
and U9280 (N_9280,N_9162,N_9193);
or U9281 (N_9281,N_9096,N_9016);
and U9282 (N_9282,N_9063,N_9062);
nand U9283 (N_9283,N_9191,N_9109);
and U9284 (N_9284,N_9037,N_9114);
or U9285 (N_9285,N_9167,N_9027);
or U9286 (N_9286,N_9068,N_9143);
nand U9287 (N_9287,N_9184,N_9095);
and U9288 (N_9288,N_9032,N_9071);
nor U9289 (N_9289,N_9125,N_9190);
nor U9290 (N_9290,N_9115,N_9079);
and U9291 (N_9291,N_9076,N_9011);
xor U9292 (N_9292,N_9137,N_9081);
nand U9293 (N_9293,N_9166,N_9097);
nand U9294 (N_9294,N_9128,N_9035);
nor U9295 (N_9295,N_9113,N_9148);
and U9296 (N_9296,N_9155,N_9017);
nor U9297 (N_9297,N_9152,N_9174);
or U9298 (N_9298,N_9141,N_9158);
nand U9299 (N_9299,N_9169,N_9030);
or U9300 (N_9300,N_9037,N_9143);
or U9301 (N_9301,N_9107,N_9118);
nand U9302 (N_9302,N_9090,N_9167);
and U9303 (N_9303,N_9108,N_9002);
or U9304 (N_9304,N_9027,N_9110);
and U9305 (N_9305,N_9030,N_9170);
and U9306 (N_9306,N_9160,N_9144);
nand U9307 (N_9307,N_9099,N_9005);
nand U9308 (N_9308,N_9199,N_9046);
nor U9309 (N_9309,N_9177,N_9080);
and U9310 (N_9310,N_9083,N_9188);
or U9311 (N_9311,N_9115,N_9043);
and U9312 (N_9312,N_9146,N_9111);
or U9313 (N_9313,N_9176,N_9177);
and U9314 (N_9314,N_9176,N_9038);
or U9315 (N_9315,N_9040,N_9148);
nand U9316 (N_9316,N_9109,N_9031);
and U9317 (N_9317,N_9197,N_9160);
nor U9318 (N_9318,N_9049,N_9151);
nor U9319 (N_9319,N_9107,N_9000);
nor U9320 (N_9320,N_9159,N_9080);
or U9321 (N_9321,N_9125,N_9072);
nor U9322 (N_9322,N_9040,N_9143);
or U9323 (N_9323,N_9197,N_9021);
nand U9324 (N_9324,N_9078,N_9113);
xor U9325 (N_9325,N_9094,N_9136);
nor U9326 (N_9326,N_9092,N_9162);
nand U9327 (N_9327,N_9111,N_9187);
or U9328 (N_9328,N_9006,N_9081);
and U9329 (N_9329,N_9029,N_9059);
nand U9330 (N_9330,N_9057,N_9199);
nand U9331 (N_9331,N_9185,N_9036);
and U9332 (N_9332,N_9060,N_9090);
nor U9333 (N_9333,N_9189,N_9110);
nor U9334 (N_9334,N_9025,N_9082);
nor U9335 (N_9335,N_9002,N_9122);
or U9336 (N_9336,N_9010,N_9195);
and U9337 (N_9337,N_9151,N_9146);
and U9338 (N_9338,N_9060,N_9134);
and U9339 (N_9339,N_9071,N_9049);
and U9340 (N_9340,N_9148,N_9155);
nor U9341 (N_9341,N_9008,N_9047);
and U9342 (N_9342,N_9104,N_9075);
nand U9343 (N_9343,N_9057,N_9101);
nor U9344 (N_9344,N_9199,N_9062);
and U9345 (N_9345,N_9185,N_9046);
nor U9346 (N_9346,N_9121,N_9154);
nor U9347 (N_9347,N_9025,N_9107);
and U9348 (N_9348,N_9023,N_9165);
or U9349 (N_9349,N_9150,N_9163);
nand U9350 (N_9350,N_9114,N_9040);
xnor U9351 (N_9351,N_9099,N_9162);
nand U9352 (N_9352,N_9172,N_9071);
nor U9353 (N_9353,N_9054,N_9192);
nand U9354 (N_9354,N_9154,N_9055);
nor U9355 (N_9355,N_9136,N_9141);
nor U9356 (N_9356,N_9053,N_9113);
xor U9357 (N_9357,N_9181,N_9023);
and U9358 (N_9358,N_9164,N_9111);
or U9359 (N_9359,N_9191,N_9022);
nand U9360 (N_9360,N_9009,N_9136);
xnor U9361 (N_9361,N_9026,N_9154);
nand U9362 (N_9362,N_9079,N_9124);
nand U9363 (N_9363,N_9074,N_9102);
nor U9364 (N_9364,N_9110,N_9039);
or U9365 (N_9365,N_9107,N_9002);
or U9366 (N_9366,N_9048,N_9125);
nor U9367 (N_9367,N_9106,N_9167);
nand U9368 (N_9368,N_9013,N_9157);
nand U9369 (N_9369,N_9188,N_9185);
or U9370 (N_9370,N_9096,N_9074);
nand U9371 (N_9371,N_9094,N_9008);
nand U9372 (N_9372,N_9092,N_9015);
and U9373 (N_9373,N_9176,N_9144);
and U9374 (N_9374,N_9128,N_9198);
nand U9375 (N_9375,N_9127,N_9192);
or U9376 (N_9376,N_9182,N_9190);
nand U9377 (N_9377,N_9049,N_9163);
and U9378 (N_9378,N_9173,N_9050);
nor U9379 (N_9379,N_9030,N_9174);
or U9380 (N_9380,N_9040,N_9164);
and U9381 (N_9381,N_9055,N_9174);
nand U9382 (N_9382,N_9042,N_9041);
or U9383 (N_9383,N_9166,N_9168);
and U9384 (N_9384,N_9098,N_9073);
or U9385 (N_9385,N_9073,N_9063);
and U9386 (N_9386,N_9037,N_9096);
or U9387 (N_9387,N_9166,N_9080);
and U9388 (N_9388,N_9112,N_9196);
nand U9389 (N_9389,N_9062,N_9067);
and U9390 (N_9390,N_9194,N_9018);
nor U9391 (N_9391,N_9070,N_9125);
or U9392 (N_9392,N_9100,N_9176);
and U9393 (N_9393,N_9141,N_9155);
nand U9394 (N_9394,N_9184,N_9186);
nand U9395 (N_9395,N_9147,N_9148);
and U9396 (N_9396,N_9107,N_9091);
nand U9397 (N_9397,N_9135,N_9104);
nand U9398 (N_9398,N_9099,N_9089);
and U9399 (N_9399,N_9186,N_9162);
or U9400 (N_9400,N_9212,N_9360);
nand U9401 (N_9401,N_9391,N_9206);
nand U9402 (N_9402,N_9389,N_9256);
nor U9403 (N_9403,N_9383,N_9232);
nor U9404 (N_9404,N_9203,N_9373);
nor U9405 (N_9405,N_9320,N_9324);
nor U9406 (N_9406,N_9245,N_9376);
and U9407 (N_9407,N_9322,N_9319);
or U9408 (N_9408,N_9267,N_9372);
or U9409 (N_9409,N_9381,N_9233);
or U9410 (N_9410,N_9226,N_9299);
nor U9411 (N_9411,N_9279,N_9303);
or U9412 (N_9412,N_9328,N_9239);
nor U9413 (N_9413,N_9315,N_9323);
nand U9414 (N_9414,N_9207,N_9399);
or U9415 (N_9415,N_9358,N_9254);
nor U9416 (N_9416,N_9326,N_9241);
or U9417 (N_9417,N_9227,N_9384);
nand U9418 (N_9418,N_9396,N_9393);
and U9419 (N_9419,N_9240,N_9243);
or U9420 (N_9420,N_9348,N_9269);
nand U9421 (N_9421,N_9223,N_9255);
and U9422 (N_9422,N_9283,N_9215);
xnor U9423 (N_9423,N_9337,N_9209);
or U9424 (N_9424,N_9306,N_9282);
or U9425 (N_9425,N_9347,N_9247);
nor U9426 (N_9426,N_9350,N_9296);
or U9427 (N_9427,N_9275,N_9272);
and U9428 (N_9428,N_9260,N_9330);
and U9429 (N_9429,N_9355,N_9268);
nand U9430 (N_9430,N_9369,N_9302);
nand U9431 (N_9431,N_9365,N_9221);
and U9432 (N_9432,N_9329,N_9379);
and U9433 (N_9433,N_9352,N_9375);
nand U9434 (N_9434,N_9325,N_9335);
nor U9435 (N_9435,N_9366,N_9292);
and U9436 (N_9436,N_9300,N_9368);
nand U9437 (N_9437,N_9289,N_9297);
or U9438 (N_9438,N_9343,N_9200);
and U9439 (N_9439,N_9367,N_9346);
or U9440 (N_9440,N_9353,N_9310);
or U9441 (N_9441,N_9261,N_9334);
or U9442 (N_9442,N_9257,N_9287);
or U9443 (N_9443,N_9208,N_9242);
nand U9444 (N_9444,N_9246,N_9238);
nand U9445 (N_9445,N_9371,N_9231);
or U9446 (N_9446,N_9249,N_9204);
or U9447 (N_9447,N_9362,N_9293);
nor U9448 (N_9448,N_9284,N_9307);
or U9449 (N_9449,N_9210,N_9363);
nor U9450 (N_9450,N_9201,N_9395);
xnor U9451 (N_9451,N_9225,N_9354);
nor U9452 (N_9452,N_9316,N_9332);
nor U9453 (N_9453,N_9341,N_9280);
and U9454 (N_9454,N_9370,N_9276);
or U9455 (N_9455,N_9274,N_9244);
or U9456 (N_9456,N_9202,N_9258);
and U9457 (N_9457,N_9342,N_9277);
and U9458 (N_9458,N_9305,N_9235);
nand U9459 (N_9459,N_9288,N_9333);
nand U9460 (N_9460,N_9278,N_9290);
and U9461 (N_9461,N_9217,N_9327);
nand U9462 (N_9462,N_9291,N_9224);
or U9463 (N_9463,N_9228,N_9252);
nor U9464 (N_9464,N_9382,N_9222);
nor U9465 (N_9465,N_9359,N_9364);
or U9466 (N_9466,N_9378,N_9294);
or U9467 (N_9467,N_9351,N_9309);
nor U9468 (N_9468,N_9308,N_9220);
nor U9469 (N_9469,N_9229,N_9285);
nor U9470 (N_9470,N_9286,N_9321);
nor U9471 (N_9471,N_9219,N_9253);
or U9472 (N_9472,N_9312,N_9356);
nand U9473 (N_9473,N_9234,N_9218);
or U9474 (N_9474,N_9345,N_9394);
nor U9475 (N_9475,N_9349,N_9301);
or U9476 (N_9476,N_9344,N_9398);
or U9477 (N_9477,N_9390,N_9317);
and U9478 (N_9478,N_9265,N_9237);
nand U9479 (N_9479,N_9262,N_9388);
and U9480 (N_9480,N_9281,N_9338);
and U9481 (N_9481,N_9271,N_9250);
nand U9482 (N_9482,N_9213,N_9386);
or U9483 (N_9483,N_9251,N_9211);
or U9484 (N_9484,N_9318,N_9331);
nor U9485 (N_9485,N_9214,N_9339);
nand U9486 (N_9486,N_9236,N_9298);
and U9487 (N_9487,N_9304,N_9264);
nand U9488 (N_9488,N_9385,N_9216);
nand U9489 (N_9489,N_9295,N_9311);
nand U9490 (N_9490,N_9313,N_9380);
nor U9491 (N_9491,N_9374,N_9263);
nor U9492 (N_9492,N_9361,N_9270);
and U9493 (N_9493,N_9314,N_9392);
or U9494 (N_9494,N_9266,N_9377);
nand U9495 (N_9495,N_9340,N_9205);
or U9496 (N_9496,N_9397,N_9230);
nand U9497 (N_9497,N_9273,N_9336);
nor U9498 (N_9498,N_9357,N_9387);
xor U9499 (N_9499,N_9248,N_9259);
nand U9500 (N_9500,N_9229,N_9276);
and U9501 (N_9501,N_9333,N_9398);
nand U9502 (N_9502,N_9342,N_9265);
nand U9503 (N_9503,N_9212,N_9338);
nand U9504 (N_9504,N_9316,N_9217);
xnor U9505 (N_9505,N_9230,N_9359);
or U9506 (N_9506,N_9315,N_9362);
and U9507 (N_9507,N_9374,N_9339);
or U9508 (N_9508,N_9258,N_9377);
or U9509 (N_9509,N_9315,N_9294);
and U9510 (N_9510,N_9312,N_9309);
and U9511 (N_9511,N_9244,N_9321);
nor U9512 (N_9512,N_9215,N_9301);
or U9513 (N_9513,N_9392,N_9363);
nor U9514 (N_9514,N_9208,N_9372);
and U9515 (N_9515,N_9306,N_9346);
or U9516 (N_9516,N_9315,N_9322);
or U9517 (N_9517,N_9312,N_9360);
nand U9518 (N_9518,N_9264,N_9310);
and U9519 (N_9519,N_9337,N_9233);
and U9520 (N_9520,N_9327,N_9302);
and U9521 (N_9521,N_9371,N_9284);
nor U9522 (N_9522,N_9356,N_9352);
or U9523 (N_9523,N_9350,N_9355);
nor U9524 (N_9524,N_9234,N_9341);
nor U9525 (N_9525,N_9258,N_9271);
nor U9526 (N_9526,N_9395,N_9295);
nand U9527 (N_9527,N_9344,N_9288);
and U9528 (N_9528,N_9396,N_9308);
and U9529 (N_9529,N_9350,N_9235);
and U9530 (N_9530,N_9331,N_9330);
or U9531 (N_9531,N_9324,N_9371);
nand U9532 (N_9532,N_9295,N_9372);
or U9533 (N_9533,N_9284,N_9273);
nand U9534 (N_9534,N_9346,N_9249);
nand U9535 (N_9535,N_9255,N_9258);
and U9536 (N_9536,N_9313,N_9246);
xnor U9537 (N_9537,N_9394,N_9208);
or U9538 (N_9538,N_9312,N_9334);
or U9539 (N_9539,N_9278,N_9354);
nor U9540 (N_9540,N_9343,N_9262);
or U9541 (N_9541,N_9386,N_9395);
and U9542 (N_9542,N_9300,N_9336);
or U9543 (N_9543,N_9392,N_9359);
nor U9544 (N_9544,N_9219,N_9345);
and U9545 (N_9545,N_9394,N_9303);
or U9546 (N_9546,N_9202,N_9383);
nor U9547 (N_9547,N_9376,N_9345);
and U9548 (N_9548,N_9363,N_9290);
nand U9549 (N_9549,N_9359,N_9328);
and U9550 (N_9550,N_9333,N_9290);
and U9551 (N_9551,N_9381,N_9316);
or U9552 (N_9552,N_9362,N_9297);
nor U9553 (N_9553,N_9399,N_9383);
and U9554 (N_9554,N_9206,N_9357);
or U9555 (N_9555,N_9287,N_9253);
nor U9556 (N_9556,N_9353,N_9271);
and U9557 (N_9557,N_9201,N_9249);
nor U9558 (N_9558,N_9274,N_9261);
nand U9559 (N_9559,N_9322,N_9350);
nand U9560 (N_9560,N_9361,N_9249);
and U9561 (N_9561,N_9224,N_9320);
and U9562 (N_9562,N_9322,N_9251);
or U9563 (N_9563,N_9202,N_9322);
and U9564 (N_9564,N_9376,N_9332);
and U9565 (N_9565,N_9316,N_9394);
nor U9566 (N_9566,N_9311,N_9215);
nand U9567 (N_9567,N_9370,N_9281);
and U9568 (N_9568,N_9325,N_9276);
nand U9569 (N_9569,N_9342,N_9369);
nand U9570 (N_9570,N_9251,N_9242);
and U9571 (N_9571,N_9245,N_9204);
nand U9572 (N_9572,N_9319,N_9221);
and U9573 (N_9573,N_9240,N_9309);
nand U9574 (N_9574,N_9231,N_9328);
nand U9575 (N_9575,N_9337,N_9399);
or U9576 (N_9576,N_9215,N_9356);
nand U9577 (N_9577,N_9249,N_9357);
nand U9578 (N_9578,N_9225,N_9215);
and U9579 (N_9579,N_9268,N_9361);
nand U9580 (N_9580,N_9333,N_9211);
nor U9581 (N_9581,N_9272,N_9372);
nand U9582 (N_9582,N_9221,N_9354);
nor U9583 (N_9583,N_9305,N_9333);
or U9584 (N_9584,N_9321,N_9200);
nor U9585 (N_9585,N_9204,N_9275);
or U9586 (N_9586,N_9219,N_9225);
nor U9587 (N_9587,N_9299,N_9329);
and U9588 (N_9588,N_9361,N_9328);
nand U9589 (N_9589,N_9213,N_9334);
nand U9590 (N_9590,N_9370,N_9257);
nand U9591 (N_9591,N_9339,N_9305);
xor U9592 (N_9592,N_9220,N_9274);
nor U9593 (N_9593,N_9389,N_9307);
nor U9594 (N_9594,N_9373,N_9226);
and U9595 (N_9595,N_9392,N_9212);
or U9596 (N_9596,N_9314,N_9260);
nor U9597 (N_9597,N_9320,N_9365);
or U9598 (N_9598,N_9262,N_9321);
nor U9599 (N_9599,N_9232,N_9352);
nand U9600 (N_9600,N_9506,N_9440);
nor U9601 (N_9601,N_9590,N_9500);
or U9602 (N_9602,N_9429,N_9553);
and U9603 (N_9603,N_9594,N_9464);
nand U9604 (N_9604,N_9486,N_9520);
and U9605 (N_9605,N_9472,N_9593);
and U9606 (N_9606,N_9544,N_9411);
and U9607 (N_9607,N_9438,N_9400);
and U9608 (N_9608,N_9416,N_9564);
and U9609 (N_9609,N_9445,N_9537);
or U9610 (N_9610,N_9530,N_9574);
and U9611 (N_9611,N_9424,N_9521);
or U9612 (N_9612,N_9460,N_9423);
nand U9613 (N_9613,N_9453,N_9558);
nor U9614 (N_9614,N_9485,N_9596);
and U9615 (N_9615,N_9437,N_9465);
nand U9616 (N_9616,N_9417,N_9497);
nand U9617 (N_9617,N_9470,N_9552);
nand U9618 (N_9618,N_9508,N_9478);
and U9619 (N_9619,N_9538,N_9403);
nand U9620 (N_9620,N_9413,N_9414);
and U9621 (N_9621,N_9581,N_9597);
or U9622 (N_9622,N_9511,N_9480);
nor U9623 (N_9623,N_9525,N_9426);
nor U9624 (N_9624,N_9582,N_9519);
nor U9625 (N_9625,N_9473,N_9536);
or U9626 (N_9626,N_9512,N_9551);
nor U9627 (N_9627,N_9563,N_9522);
nand U9628 (N_9628,N_9458,N_9436);
and U9629 (N_9629,N_9573,N_9578);
xnor U9630 (N_9630,N_9496,N_9557);
or U9631 (N_9631,N_9404,N_9481);
nor U9632 (N_9632,N_9570,N_9586);
nor U9633 (N_9633,N_9584,N_9535);
nand U9634 (N_9634,N_9408,N_9444);
nand U9635 (N_9635,N_9533,N_9556);
or U9636 (N_9636,N_9412,N_9523);
and U9637 (N_9637,N_9490,N_9483);
and U9638 (N_9638,N_9554,N_9461);
or U9639 (N_9639,N_9524,N_9569);
and U9640 (N_9640,N_9505,N_9503);
nor U9641 (N_9641,N_9442,N_9431);
and U9642 (N_9642,N_9587,N_9491);
nand U9643 (N_9643,N_9409,N_9542);
nand U9644 (N_9644,N_9441,N_9539);
nor U9645 (N_9645,N_9459,N_9540);
nand U9646 (N_9646,N_9532,N_9526);
nand U9647 (N_9647,N_9567,N_9531);
and U9648 (N_9648,N_9430,N_9572);
nor U9649 (N_9649,N_9418,N_9422);
or U9650 (N_9650,N_9467,N_9488);
nand U9651 (N_9651,N_9468,N_9580);
or U9652 (N_9652,N_9575,N_9501);
nand U9653 (N_9653,N_9498,N_9562);
nand U9654 (N_9654,N_9433,N_9543);
nand U9655 (N_9655,N_9446,N_9439);
nor U9656 (N_9656,N_9482,N_9469);
nor U9657 (N_9657,N_9518,N_9517);
nand U9658 (N_9658,N_9528,N_9415);
or U9659 (N_9659,N_9583,N_9435);
nor U9660 (N_9660,N_9476,N_9443);
and U9661 (N_9661,N_9571,N_9555);
nand U9662 (N_9662,N_9502,N_9549);
and U9663 (N_9663,N_9509,N_9595);
and U9664 (N_9664,N_9499,N_9577);
and U9665 (N_9665,N_9471,N_9487);
and U9666 (N_9666,N_9420,N_9515);
or U9667 (N_9667,N_9579,N_9454);
nor U9668 (N_9668,N_9492,N_9489);
nor U9669 (N_9669,N_9545,N_9585);
xor U9670 (N_9670,N_9462,N_9566);
nand U9671 (N_9671,N_9541,N_9548);
nand U9672 (N_9672,N_9402,N_9463);
and U9673 (N_9673,N_9547,N_9434);
and U9674 (N_9674,N_9504,N_9516);
nor U9675 (N_9675,N_9419,N_9527);
or U9676 (N_9676,N_9477,N_9568);
or U9677 (N_9677,N_9410,N_9427);
or U9678 (N_9678,N_9450,N_9455);
nand U9679 (N_9679,N_9428,N_9457);
nor U9680 (N_9680,N_9565,N_9561);
nand U9681 (N_9681,N_9510,N_9546);
and U9682 (N_9682,N_9449,N_9447);
and U9683 (N_9683,N_9550,N_9592);
xor U9684 (N_9684,N_9495,N_9448);
nand U9685 (N_9685,N_9475,N_9466);
or U9686 (N_9686,N_9452,N_9591);
or U9687 (N_9687,N_9598,N_9589);
or U9688 (N_9688,N_9507,N_9484);
and U9689 (N_9689,N_9534,N_9493);
and U9690 (N_9690,N_9599,N_9529);
nand U9691 (N_9691,N_9425,N_9513);
nand U9692 (N_9692,N_9559,N_9421);
nor U9693 (N_9693,N_9401,N_9479);
and U9694 (N_9694,N_9456,N_9474);
or U9695 (N_9695,N_9451,N_9494);
nand U9696 (N_9696,N_9405,N_9576);
and U9697 (N_9697,N_9514,N_9432);
or U9698 (N_9698,N_9407,N_9588);
and U9699 (N_9699,N_9560,N_9406);
nor U9700 (N_9700,N_9421,N_9476);
or U9701 (N_9701,N_9525,N_9537);
or U9702 (N_9702,N_9431,N_9469);
or U9703 (N_9703,N_9501,N_9567);
nand U9704 (N_9704,N_9431,N_9566);
nor U9705 (N_9705,N_9485,N_9597);
and U9706 (N_9706,N_9594,N_9442);
and U9707 (N_9707,N_9521,N_9524);
nand U9708 (N_9708,N_9462,N_9576);
and U9709 (N_9709,N_9439,N_9558);
nor U9710 (N_9710,N_9559,N_9570);
nand U9711 (N_9711,N_9516,N_9491);
nand U9712 (N_9712,N_9538,N_9508);
nand U9713 (N_9713,N_9447,N_9402);
and U9714 (N_9714,N_9501,N_9581);
nand U9715 (N_9715,N_9455,N_9460);
or U9716 (N_9716,N_9490,N_9509);
nor U9717 (N_9717,N_9453,N_9499);
nand U9718 (N_9718,N_9510,N_9500);
nand U9719 (N_9719,N_9496,N_9592);
nor U9720 (N_9720,N_9475,N_9438);
nor U9721 (N_9721,N_9441,N_9491);
nand U9722 (N_9722,N_9587,N_9467);
or U9723 (N_9723,N_9453,N_9583);
and U9724 (N_9724,N_9422,N_9419);
or U9725 (N_9725,N_9418,N_9513);
and U9726 (N_9726,N_9592,N_9492);
and U9727 (N_9727,N_9465,N_9414);
nand U9728 (N_9728,N_9475,N_9459);
or U9729 (N_9729,N_9442,N_9482);
or U9730 (N_9730,N_9541,N_9511);
and U9731 (N_9731,N_9431,N_9471);
nand U9732 (N_9732,N_9410,N_9429);
and U9733 (N_9733,N_9533,N_9512);
nand U9734 (N_9734,N_9530,N_9432);
nand U9735 (N_9735,N_9576,N_9553);
or U9736 (N_9736,N_9476,N_9439);
and U9737 (N_9737,N_9567,N_9504);
and U9738 (N_9738,N_9495,N_9451);
or U9739 (N_9739,N_9485,N_9498);
and U9740 (N_9740,N_9483,N_9484);
or U9741 (N_9741,N_9543,N_9535);
nand U9742 (N_9742,N_9599,N_9474);
and U9743 (N_9743,N_9469,N_9566);
and U9744 (N_9744,N_9580,N_9535);
xnor U9745 (N_9745,N_9483,N_9520);
or U9746 (N_9746,N_9489,N_9584);
nor U9747 (N_9747,N_9497,N_9491);
and U9748 (N_9748,N_9408,N_9592);
nor U9749 (N_9749,N_9465,N_9481);
nand U9750 (N_9750,N_9440,N_9548);
or U9751 (N_9751,N_9401,N_9597);
and U9752 (N_9752,N_9407,N_9458);
nand U9753 (N_9753,N_9420,N_9455);
and U9754 (N_9754,N_9459,N_9439);
and U9755 (N_9755,N_9542,N_9557);
nor U9756 (N_9756,N_9484,N_9520);
and U9757 (N_9757,N_9598,N_9472);
and U9758 (N_9758,N_9420,N_9491);
nor U9759 (N_9759,N_9597,N_9413);
nor U9760 (N_9760,N_9498,N_9450);
nor U9761 (N_9761,N_9443,N_9470);
and U9762 (N_9762,N_9517,N_9549);
nor U9763 (N_9763,N_9522,N_9499);
xor U9764 (N_9764,N_9483,N_9494);
nand U9765 (N_9765,N_9405,N_9554);
nand U9766 (N_9766,N_9526,N_9405);
or U9767 (N_9767,N_9449,N_9561);
nand U9768 (N_9768,N_9523,N_9539);
and U9769 (N_9769,N_9555,N_9430);
nand U9770 (N_9770,N_9506,N_9416);
nor U9771 (N_9771,N_9432,N_9479);
nor U9772 (N_9772,N_9404,N_9418);
nor U9773 (N_9773,N_9522,N_9419);
or U9774 (N_9774,N_9421,N_9429);
nand U9775 (N_9775,N_9405,N_9482);
and U9776 (N_9776,N_9454,N_9419);
and U9777 (N_9777,N_9548,N_9453);
nand U9778 (N_9778,N_9446,N_9488);
or U9779 (N_9779,N_9508,N_9541);
nor U9780 (N_9780,N_9503,N_9513);
and U9781 (N_9781,N_9517,N_9487);
or U9782 (N_9782,N_9526,N_9400);
and U9783 (N_9783,N_9536,N_9577);
xnor U9784 (N_9784,N_9501,N_9444);
nand U9785 (N_9785,N_9504,N_9507);
and U9786 (N_9786,N_9454,N_9513);
nor U9787 (N_9787,N_9533,N_9537);
nor U9788 (N_9788,N_9451,N_9589);
nand U9789 (N_9789,N_9447,N_9423);
or U9790 (N_9790,N_9497,N_9532);
and U9791 (N_9791,N_9459,N_9420);
nand U9792 (N_9792,N_9494,N_9531);
and U9793 (N_9793,N_9424,N_9460);
nor U9794 (N_9794,N_9538,N_9414);
and U9795 (N_9795,N_9588,N_9503);
nand U9796 (N_9796,N_9542,N_9571);
and U9797 (N_9797,N_9432,N_9509);
or U9798 (N_9798,N_9463,N_9554);
nand U9799 (N_9799,N_9448,N_9569);
nand U9800 (N_9800,N_9794,N_9677);
nor U9801 (N_9801,N_9661,N_9695);
or U9802 (N_9802,N_9699,N_9714);
nor U9803 (N_9803,N_9624,N_9748);
nand U9804 (N_9804,N_9747,N_9608);
and U9805 (N_9805,N_9731,N_9739);
or U9806 (N_9806,N_9724,N_9766);
nand U9807 (N_9807,N_9735,N_9637);
and U9808 (N_9808,N_9723,N_9701);
nor U9809 (N_9809,N_9795,N_9689);
and U9810 (N_9810,N_9643,N_9705);
or U9811 (N_9811,N_9706,N_9660);
nand U9812 (N_9812,N_9619,N_9653);
and U9813 (N_9813,N_9712,N_9767);
nor U9814 (N_9814,N_9763,N_9617);
or U9815 (N_9815,N_9764,N_9671);
and U9816 (N_9816,N_9725,N_9758);
xnor U9817 (N_9817,N_9652,N_9776);
or U9818 (N_9818,N_9721,N_9741);
nor U9819 (N_9819,N_9734,N_9663);
nor U9820 (N_9820,N_9761,N_9788);
and U9821 (N_9821,N_9680,N_9785);
or U9822 (N_9822,N_9631,N_9717);
or U9823 (N_9823,N_9782,N_9676);
or U9824 (N_9824,N_9772,N_9683);
nand U9825 (N_9825,N_9698,N_9799);
and U9826 (N_9826,N_9623,N_9633);
nor U9827 (N_9827,N_9786,N_9783);
and U9828 (N_9828,N_9716,N_9679);
or U9829 (N_9829,N_9726,N_9736);
and U9830 (N_9830,N_9727,N_9757);
nor U9831 (N_9831,N_9775,N_9635);
and U9832 (N_9832,N_9667,N_9669);
nand U9833 (N_9833,N_9618,N_9729);
nand U9834 (N_9834,N_9611,N_9632);
or U9835 (N_9835,N_9605,N_9681);
or U9836 (N_9836,N_9774,N_9620);
nor U9837 (N_9837,N_9642,N_9700);
nor U9838 (N_9838,N_9659,N_9609);
nor U9839 (N_9839,N_9606,N_9627);
nand U9840 (N_9840,N_9746,N_9665);
nor U9841 (N_9841,N_9674,N_9645);
and U9842 (N_9842,N_9696,N_9670);
nor U9843 (N_9843,N_9648,N_9773);
or U9844 (N_9844,N_9733,N_9797);
nor U9845 (N_9845,N_9730,N_9644);
or U9846 (N_9846,N_9654,N_9762);
or U9847 (N_9847,N_9778,N_9749);
nand U9848 (N_9848,N_9787,N_9702);
nand U9849 (N_9849,N_9718,N_9621);
or U9850 (N_9850,N_9612,N_9668);
nor U9851 (N_9851,N_9742,N_9745);
and U9852 (N_9852,N_9607,N_9708);
and U9853 (N_9853,N_9754,N_9770);
and U9854 (N_9854,N_9602,N_9710);
and U9855 (N_9855,N_9751,N_9780);
nor U9856 (N_9856,N_9629,N_9655);
or U9857 (N_9857,N_9638,N_9771);
or U9858 (N_9858,N_9744,N_9634);
nor U9859 (N_9859,N_9672,N_9636);
nand U9860 (N_9860,N_9688,N_9792);
and U9861 (N_9861,N_9759,N_9651);
nor U9862 (N_9862,N_9686,N_9781);
and U9863 (N_9863,N_9719,N_9639);
or U9864 (N_9864,N_9715,N_9707);
nand U9865 (N_9865,N_9650,N_9791);
nor U9866 (N_9866,N_9685,N_9768);
or U9867 (N_9867,N_9760,N_9709);
xor U9868 (N_9868,N_9697,N_9750);
nor U9869 (N_9869,N_9711,N_9647);
nand U9870 (N_9870,N_9666,N_9640);
nor U9871 (N_9871,N_9658,N_9704);
nor U9872 (N_9872,N_9613,N_9601);
or U9873 (N_9873,N_9690,N_9755);
and U9874 (N_9874,N_9678,N_9614);
nand U9875 (N_9875,N_9692,N_9684);
nand U9876 (N_9876,N_9682,N_9779);
nor U9877 (N_9877,N_9693,N_9740);
nand U9878 (N_9878,N_9790,N_9649);
or U9879 (N_9879,N_9784,N_9756);
and U9880 (N_9880,N_9752,N_9722);
nand U9881 (N_9881,N_9662,N_9641);
nand U9882 (N_9882,N_9600,N_9753);
nor U9883 (N_9883,N_9656,N_9616);
or U9884 (N_9884,N_9675,N_9604);
nor U9885 (N_9885,N_9694,N_9728);
or U9886 (N_9886,N_9687,N_9673);
nor U9887 (N_9887,N_9789,N_9664);
and U9888 (N_9888,N_9703,N_9765);
or U9889 (N_9889,N_9738,N_9646);
or U9890 (N_9890,N_9628,N_9691);
nand U9891 (N_9891,N_9732,N_9769);
nand U9892 (N_9892,N_9798,N_9777);
and U9893 (N_9893,N_9713,N_9625);
xnor U9894 (N_9894,N_9622,N_9720);
xor U9895 (N_9895,N_9793,N_9657);
nor U9896 (N_9896,N_9603,N_9796);
nor U9897 (N_9897,N_9615,N_9626);
nor U9898 (N_9898,N_9737,N_9610);
nor U9899 (N_9899,N_9630,N_9743);
nand U9900 (N_9900,N_9716,N_9774);
nor U9901 (N_9901,N_9610,N_9745);
or U9902 (N_9902,N_9626,N_9749);
nand U9903 (N_9903,N_9649,N_9701);
nor U9904 (N_9904,N_9654,N_9616);
nor U9905 (N_9905,N_9729,N_9642);
nor U9906 (N_9906,N_9750,N_9649);
and U9907 (N_9907,N_9683,N_9704);
or U9908 (N_9908,N_9776,N_9737);
nor U9909 (N_9909,N_9680,N_9609);
or U9910 (N_9910,N_9737,N_9653);
nand U9911 (N_9911,N_9671,N_9664);
and U9912 (N_9912,N_9642,N_9735);
xor U9913 (N_9913,N_9681,N_9632);
nor U9914 (N_9914,N_9668,N_9678);
or U9915 (N_9915,N_9715,N_9772);
and U9916 (N_9916,N_9781,N_9683);
and U9917 (N_9917,N_9729,N_9759);
and U9918 (N_9918,N_9664,N_9712);
nand U9919 (N_9919,N_9747,N_9643);
nor U9920 (N_9920,N_9651,N_9683);
or U9921 (N_9921,N_9650,N_9615);
and U9922 (N_9922,N_9715,N_9659);
nor U9923 (N_9923,N_9664,N_9713);
nand U9924 (N_9924,N_9739,N_9637);
or U9925 (N_9925,N_9651,N_9649);
nand U9926 (N_9926,N_9756,N_9787);
or U9927 (N_9927,N_9778,N_9617);
nor U9928 (N_9928,N_9791,N_9642);
and U9929 (N_9929,N_9761,N_9648);
nor U9930 (N_9930,N_9654,N_9712);
nand U9931 (N_9931,N_9793,N_9654);
nor U9932 (N_9932,N_9779,N_9620);
and U9933 (N_9933,N_9647,N_9757);
or U9934 (N_9934,N_9768,N_9660);
nor U9935 (N_9935,N_9713,N_9695);
and U9936 (N_9936,N_9715,N_9699);
nand U9937 (N_9937,N_9642,N_9685);
nor U9938 (N_9938,N_9626,N_9772);
or U9939 (N_9939,N_9660,N_9796);
or U9940 (N_9940,N_9701,N_9637);
and U9941 (N_9941,N_9648,N_9691);
nand U9942 (N_9942,N_9619,N_9782);
or U9943 (N_9943,N_9649,N_9603);
nand U9944 (N_9944,N_9737,N_9682);
or U9945 (N_9945,N_9779,N_9649);
nand U9946 (N_9946,N_9700,N_9684);
nand U9947 (N_9947,N_9653,N_9606);
and U9948 (N_9948,N_9767,N_9719);
or U9949 (N_9949,N_9766,N_9776);
nor U9950 (N_9950,N_9652,N_9778);
nand U9951 (N_9951,N_9749,N_9732);
or U9952 (N_9952,N_9688,N_9683);
nand U9953 (N_9953,N_9704,N_9680);
nor U9954 (N_9954,N_9734,N_9632);
and U9955 (N_9955,N_9794,N_9724);
and U9956 (N_9956,N_9755,N_9735);
nor U9957 (N_9957,N_9652,N_9617);
or U9958 (N_9958,N_9666,N_9682);
nor U9959 (N_9959,N_9640,N_9732);
or U9960 (N_9960,N_9628,N_9718);
nor U9961 (N_9961,N_9794,N_9789);
nor U9962 (N_9962,N_9706,N_9694);
and U9963 (N_9963,N_9682,N_9647);
or U9964 (N_9964,N_9673,N_9738);
nand U9965 (N_9965,N_9703,N_9751);
or U9966 (N_9966,N_9778,N_9774);
nor U9967 (N_9967,N_9782,N_9646);
and U9968 (N_9968,N_9753,N_9779);
nand U9969 (N_9969,N_9773,N_9691);
and U9970 (N_9970,N_9611,N_9775);
nor U9971 (N_9971,N_9707,N_9629);
nand U9972 (N_9972,N_9645,N_9735);
or U9973 (N_9973,N_9783,N_9670);
or U9974 (N_9974,N_9614,N_9699);
nand U9975 (N_9975,N_9687,N_9647);
and U9976 (N_9976,N_9681,N_9680);
and U9977 (N_9977,N_9686,N_9739);
nor U9978 (N_9978,N_9647,N_9654);
and U9979 (N_9979,N_9680,N_9615);
nor U9980 (N_9980,N_9775,N_9689);
or U9981 (N_9981,N_9606,N_9746);
xnor U9982 (N_9982,N_9648,N_9766);
nor U9983 (N_9983,N_9632,N_9743);
or U9984 (N_9984,N_9778,N_9683);
and U9985 (N_9985,N_9628,N_9609);
or U9986 (N_9986,N_9626,N_9675);
or U9987 (N_9987,N_9635,N_9652);
or U9988 (N_9988,N_9764,N_9608);
nand U9989 (N_9989,N_9761,N_9681);
and U9990 (N_9990,N_9778,N_9698);
and U9991 (N_9991,N_9611,N_9648);
nand U9992 (N_9992,N_9724,N_9740);
and U9993 (N_9993,N_9617,N_9601);
or U9994 (N_9994,N_9692,N_9660);
nand U9995 (N_9995,N_9603,N_9748);
nand U9996 (N_9996,N_9733,N_9650);
nor U9997 (N_9997,N_9767,N_9666);
nor U9998 (N_9998,N_9746,N_9661);
nor U9999 (N_9999,N_9635,N_9644);
nor UO_0 (O_0,N_9958,N_9923);
nand UO_1 (O_1,N_9881,N_9905);
or UO_2 (O_2,N_9828,N_9993);
nand UO_3 (O_3,N_9877,N_9863);
or UO_4 (O_4,N_9812,N_9996);
and UO_5 (O_5,N_9896,N_9949);
or UO_6 (O_6,N_9891,N_9983);
and UO_7 (O_7,N_9959,N_9872);
and UO_8 (O_8,N_9909,N_9986);
nor UO_9 (O_9,N_9814,N_9928);
or UO_10 (O_10,N_9984,N_9966);
xnor UO_11 (O_11,N_9841,N_9810);
and UO_12 (O_12,N_9851,N_9803);
or UO_13 (O_13,N_9951,N_9939);
nand UO_14 (O_14,N_9957,N_9809);
or UO_15 (O_15,N_9871,N_9906);
nand UO_16 (O_16,N_9802,N_9947);
nand UO_17 (O_17,N_9974,N_9965);
and UO_18 (O_18,N_9852,N_9825);
and UO_19 (O_19,N_9945,N_9840);
xor UO_20 (O_20,N_9930,N_9824);
nand UO_21 (O_21,N_9969,N_9913);
and UO_22 (O_22,N_9893,N_9873);
and UO_23 (O_23,N_9833,N_9992);
or UO_24 (O_24,N_9808,N_9875);
and UO_25 (O_25,N_9937,N_9995);
nand UO_26 (O_26,N_9925,N_9817);
nand UO_27 (O_27,N_9868,N_9832);
or UO_28 (O_28,N_9910,N_9922);
and UO_29 (O_29,N_9862,N_9861);
nand UO_30 (O_30,N_9933,N_9929);
and UO_31 (O_31,N_9813,N_9914);
nand UO_32 (O_32,N_9811,N_9853);
or UO_33 (O_33,N_9847,N_9952);
nor UO_34 (O_34,N_9890,N_9882);
nand UO_35 (O_35,N_9846,N_9934);
nor UO_36 (O_36,N_9878,N_9834);
or UO_37 (O_37,N_9935,N_9854);
nand UO_38 (O_38,N_9999,N_9936);
and UO_39 (O_39,N_9982,N_9956);
nor UO_40 (O_40,N_9979,N_9997);
nor UO_41 (O_41,N_9860,N_9902);
and UO_42 (O_42,N_9917,N_9908);
or UO_43 (O_43,N_9822,N_9980);
nor UO_44 (O_44,N_9887,N_9816);
nand UO_45 (O_45,N_9911,N_9850);
nor UO_46 (O_46,N_9801,N_9831);
and UO_47 (O_47,N_9838,N_9904);
nand UO_48 (O_48,N_9848,N_9892);
and UO_49 (O_49,N_9968,N_9955);
nor UO_50 (O_50,N_9823,N_9869);
or UO_51 (O_51,N_9919,N_9954);
and UO_52 (O_52,N_9827,N_9895);
and UO_53 (O_53,N_9843,N_9883);
nand UO_54 (O_54,N_9973,N_9916);
and UO_55 (O_55,N_9830,N_9855);
nor UO_56 (O_56,N_9888,N_9865);
or UO_57 (O_57,N_9907,N_9899);
nand UO_58 (O_58,N_9804,N_9960);
nor UO_59 (O_59,N_9915,N_9978);
or UO_60 (O_60,N_9839,N_9900);
nand UO_61 (O_61,N_9963,N_9876);
nor UO_62 (O_62,N_9858,N_9931);
and UO_63 (O_63,N_9867,N_9800);
or UO_64 (O_64,N_9807,N_9857);
nand UO_65 (O_65,N_9806,N_9856);
nor UO_66 (O_66,N_9912,N_9964);
nor UO_67 (O_67,N_9970,N_9897);
nand UO_68 (O_68,N_9805,N_9998);
and UO_69 (O_69,N_9961,N_9938);
or UO_70 (O_70,N_9987,N_9829);
or UO_71 (O_71,N_9866,N_9981);
nor UO_72 (O_72,N_9874,N_9837);
or UO_73 (O_73,N_9818,N_9880);
or UO_74 (O_74,N_9835,N_9942);
nor UO_75 (O_75,N_9977,N_9884);
nand UO_76 (O_76,N_9924,N_9948);
nand UO_77 (O_77,N_9889,N_9953);
and UO_78 (O_78,N_9920,N_9901);
and UO_79 (O_79,N_9826,N_9990);
and UO_80 (O_80,N_9821,N_9971);
nor UO_81 (O_81,N_9972,N_9836);
xnor UO_82 (O_82,N_9940,N_9849);
nand UO_83 (O_83,N_9815,N_9976);
and UO_84 (O_84,N_9932,N_9989);
and UO_85 (O_85,N_9926,N_9941);
nand UO_86 (O_86,N_9898,N_9921);
or UO_87 (O_87,N_9943,N_9985);
nor UO_88 (O_88,N_9886,N_9975);
nand UO_89 (O_89,N_9946,N_9842);
and UO_90 (O_90,N_9988,N_9864);
or UO_91 (O_91,N_9944,N_9885);
nand UO_92 (O_92,N_9903,N_9950);
nor UO_93 (O_93,N_9820,N_9962);
nor UO_94 (O_94,N_9894,N_9859);
nand UO_95 (O_95,N_9918,N_9967);
and UO_96 (O_96,N_9819,N_9927);
or UO_97 (O_97,N_9844,N_9994);
or UO_98 (O_98,N_9870,N_9879);
and UO_99 (O_99,N_9845,N_9991);
and UO_100 (O_100,N_9840,N_9815);
and UO_101 (O_101,N_9834,N_9858);
or UO_102 (O_102,N_9836,N_9890);
and UO_103 (O_103,N_9989,N_9905);
nand UO_104 (O_104,N_9928,N_9877);
or UO_105 (O_105,N_9940,N_9918);
and UO_106 (O_106,N_9889,N_9924);
nor UO_107 (O_107,N_9902,N_9937);
and UO_108 (O_108,N_9815,N_9912);
and UO_109 (O_109,N_9965,N_9908);
and UO_110 (O_110,N_9975,N_9835);
or UO_111 (O_111,N_9935,N_9887);
nand UO_112 (O_112,N_9825,N_9815);
and UO_113 (O_113,N_9834,N_9911);
or UO_114 (O_114,N_9884,N_9910);
or UO_115 (O_115,N_9886,N_9994);
nor UO_116 (O_116,N_9870,N_9912);
and UO_117 (O_117,N_9916,N_9921);
nand UO_118 (O_118,N_9851,N_9998);
nand UO_119 (O_119,N_9832,N_9909);
and UO_120 (O_120,N_9829,N_9973);
nor UO_121 (O_121,N_9886,N_9992);
nor UO_122 (O_122,N_9854,N_9856);
nand UO_123 (O_123,N_9922,N_9903);
nor UO_124 (O_124,N_9807,N_9956);
nand UO_125 (O_125,N_9819,N_9833);
and UO_126 (O_126,N_9926,N_9831);
nand UO_127 (O_127,N_9891,N_9893);
and UO_128 (O_128,N_9875,N_9851);
or UO_129 (O_129,N_9849,N_9818);
and UO_130 (O_130,N_9817,N_9998);
and UO_131 (O_131,N_9947,N_9904);
nand UO_132 (O_132,N_9906,N_9802);
and UO_133 (O_133,N_9880,N_9951);
nor UO_134 (O_134,N_9982,N_9939);
nor UO_135 (O_135,N_9800,N_9943);
nand UO_136 (O_136,N_9868,N_9817);
and UO_137 (O_137,N_9906,N_9927);
nor UO_138 (O_138,N_9810,N_9831);
nand UO_139 (O_139,N_9897,N_9916);
nor UO_140 (O_140,N_9806,N_9966);
nand UO_141 (O_141,N_9888,N_9922);
or UO_142 (O_142,N_9824,N_9810);
nand UO_143 (O_143,N_9908,N_9976);
and UO_144 (O_144,N_9925,N_9866);
or UO_145 (O_145,N_9942,N_9891);
nand UO_146 (O_146,N_9876,N_9861);
and UO_147 (O_147,N_9988,N_9984);
or UO_148 (O_148,N_9958,N_9814);
xnor UO_149 (O_149,N_9853,N_9983);
or UO_150 (O_150,N_9834,N_9825);
and UO_151 (O_151,N_9846,N_9862);
nand UO_152 (O_152,N_9934,N_9938);
nand UO_153 (O_153,N_9832,N_9930);
nand UO_154 (O_154,N_9957,N_9893);
nor UO_155 (O_155,N_9909,N_9908);
and UO_156 (O_156,N_9839,N_9943);
nand UO_157 (O_157,N_9987,N_9808);
nand UO_158 (O_158,N_9803,N_9971);
and UO_159 (O_159,N_9866,N_9822);
and UO_160 (O_160,N_9948,N_9975);
or UO_161 (O_161,N_9938,N_9984);
and UO_162 (O_162,N_9811,N_9920);
nand UO_163 (O_163,N_9831,N_9936);
or UO_164 (O_164,N_9828,N_9967);
nand UO_165 (O_165,N_9929,N_9830);
or UO_166 (O_166,N_9951,N_9901);
nor UO_167 (O_167,N_9919,N_9935);
nor UO_168 (O_168,N_9951,N_9820);
nand UO_169 (O_169,N_9818,N_9907);
nand UO_170 (O_170,N_9886,N_9802);
and UO_171 (O_171,N_9808,N_9961);
or UO_172 (O_172,N_9875,N_9853);
and UO_173 (O_173,N_9947,N_9889);
or UO_174 (O_174,N_9872,N_9804);
nor UO_175 (O_175,N_9960,N_9996);
or UO_176 (O_176,N_9949,N_9826);
nand UO_177 (O_177,N_9861,N_9986);
nor UO_178 (O_178,N_9877,N_9887);
and UO_179 (O_179,N_9981,N_9943);
or UO_180 (O_180,N_9935,N_9993);
nor UO_181 (O_181,N_9953,N_9912);
and UO_182 (O_182,N_9967,N_9826);
or UO_183 (O_183,N_9973,N_9835);
xnor UO_184 (O_184,N_9820,N_9965);
and UO_185 (O_185,N_9819,N_9948);
and UO_186 (O_186,N_9806,N_9984);
or UO_187 (O_187,N_9997,N_9851);
and UO_188 (O_188,N_9824,N_9992);
nor UO_189 (O_189,N_9801,N_9829);
and UO_190 (O_190,N_9976,N_9866);
and UO_191 (O_191,N_9801,N_9949);
nor UO_192 (O_192,N_9974,N_9903);
nand UO_193 (O_193,N_9858,N_9924);
xor UO_194 (O_194,N_9809,N_9990);
or UO_195 (O_195,N_9989,N_9826);
or UO_196 (O_196,N_9917,N_9986);
nand UO_197 (O_197,N_9928,N_9955);
nand UO_198 (O_198,N_9801,N_9915);
nand UO_199 (O_199,N_9943,N_9820);
nand UO_200 (O_200,N_9864,N_9924);
nand UO_201 (O_201,N_9872,N_9846);
nor UO_202 (O_202,N_9899,N_9875);
and UO_203 (O_203,N_9834,N_9853);
nor UO_204 (O_204,N_9835,N_9950);
or UO_205 (O_205,N_9901,N_9954);
nor UO_206 (O_206,N_9813,N_9898);
or UO_207 (O_207,N_9807,N_9945);
nand UO_208 (O_208,N_9902,N_9943);
nand UO_209 (O_209,N_9830,N_9883);
nor UO_210 (O_210,N_9874,N_9984);
or UO_211 (O_211,N_9819,N_9848);
and UO_212 (O_212,N_9911,N_9856);
xor UO_213 (O_213,N_9850,N_9943);
or UO_214 (O_214,N_9845,N_9803);
nor UO_215 (O_215,N_9930,N_9878);
or UO_216 (O_216,N_9918,N_9943);
nor UO_217 (O_217,N_9821,N_9935);
nand UO_218 (O_218,N_9916,N_9977);
or UO_219 (O_219,N_9831,N_9835);
xor UO_220 (O_220,N_9885,N_9895);
or UO_221 (O_221,N_9803,N_9957);
nor UO_222 (O_222,N_9934,N_9843);
or UO_223 (O_223,N_9837,N_9878);
nor UO_224 (O_224,N_9878,N_9915);
nor UO_225 (O_225,N_9886,N_9921);
and UO_226 (O_226,N_9880,N_9976);
and UO_227 (O_227,N_9986,N_9961);
nand UO_228 (O_228,N_9806,N_9842);
or UO_229 (O_229,N_9994,N_9869);
or UO_230 (O_230,N_9968,N_9980);
nor UO_231 (O_231,N_9876,N_9996);
nand UO_232 (O_232,N_9974,N_9838);
nand UO_233 (O_233,N_9916,N_9938);
nor UO_234 (O_234,N_9977,N_9807);
and UO_235 (O_235,N_9852,N_9872);
nor UO_236 (O_236,N_9945,N_9854);
or UO_237 (O_237,N_9936,N_9872);
nor UO_238 (O_238,N_9865,N_9891);
or UO_239 (O_239,N_9873,N_9945);
nand UO_240 (O_240,N_9826,N_9834);
and UO_241 (O_241,N_9957,N_9845);
and UO_242 (O_242,N_9819,N_9811);
and UO_243 (O_243,N_9837,N_9903);
and UO_244 (O_244,N_9911,N_9994);
or UO_245 (O_245,N_9803,N_9904);
and UO_246 (O_246,N_9866,N_9853);
and UO_247 (O_247,N_9840,N_9914);
or UO_248 (O_248,N_9814,N_9907);
and UO_249 (O_249,N_9826,N_9999);
nand UO_250 (O_250,N_9899,N_9844);
xor UO_251 (O_251,N_9928,N_9996);
and UO_252 (O_252,N_9912,N_9892);
or UO_253 (O_253,N_9913,N_9804);
and UO_254 (O_254,N_9825,N_9828);
nor UO_255 (O_255,N_9884,N_9897);
and UO_256 (O_256,N_9836,N_9842);
and UO_257 (O_257,N_9875,N_9984);
xor UO_258 (O_258,N_9924,N_9822);
and UO_259 (O_259,N_9885,N_9981);
nor UO_260 (O_260,N_9906,N_9970);
and UO_261 (O_261,N_9915,N_9989);
nand UO_262 (O_262,N_9977,N_9967);
and UO_263 (O_263,N_9876,N_9923);
nor UO_264 (O_264,N_9853,N_9817);
nand UO_265 (O_265,N_9955,N_9858);
or UO_266 (O_266,N_9812,N_9818);
nor UO_267 (O_267,N_9867,N_9809);
nor UO_268 (O_268,N_9845,N_9835);
or UO_269 (O_269,N_9839,N_9827);
or UO_270 (O_270,N_9803,N_9974);
nand UO_271 (O_271,N_9882,N_9866);
nand UO_272 (O_272,N_9854,N_9961);
and UO_273 (O_273,N_9815,N_9880);
and UO_274 (O_274,N_9943,N_9920);
nand UO_275 (O_275,N_9906,N_9931);
nor UO_276 (O_276,N_9963,N_9936);
and UO_277 (O_277,N_9810,N_9855);
nand UO_278 (O_278,N_9839,N_9859);
nand UO_279 (O_279,N_9840,N_9866);
or UO_280 (O_280,N_9975,N_9910);
nand UO_281 (O_281,N_9893,N_9941);
nand UO_282 (O_282,N_9937,N_9825);
nor UO_283 (O_283,N_9839,N_9887);
or UO_284 (O_284,N_9854,N_9825);
nor UO_285 (O_285,N_9956,N_9843);
nand UO_286 (O_286,N_9810,N_9936);
nor UO_287 (O_287,N_9994,N_9852);
or UO_288 (O_288,N_9812,N_9848);
and UO_289 (O_289,N_9989,N_9805);
and UO_290 (O_290,N_9957,N_9829);
or UO_291 (O_291,N_9962,N_9982);
and UO_292 (O_292,N_9939,N_9911);
nand UO_293 (O_293,N_9928,N_9904);
or UO_294 (O_294,N_9991,N_9812);
nand UO_295 (O_295,N_9889,N_9913);
and UO_296 (O_296,N_9949,N_9811);
or UO_297 (O_297,N_9820,N_9934);
nor UO_298 (O_298,N_9866,N_9966);
or UO_299 (O_299,N_9805,N_9876);
or UO_300 (O_300,N_9874,N_9944);
and UO_301 (O_301,N_9890,N_9866);
nor UO_302 (O_302,N_9833,N_9893);
nor UO_303 (O_303,N_9946,N_9886);
or UO_304 (O_304,N_9979,N_9807);
nand UO_305 (O_305,N_9981,N_9830);
nand UO_306 (O_306,N_9818,N_9870);
and UO_307 (O_307,N_9805,N_9841);
or UO_308 (O_308,N_9857,N_9949);
nand UO_309 (O_309,N_9834,N_9827);
nor UO_310 (O_310,N_9945,N_9894);
nand UO_311 (O_311,N_9953,N_9846);
and UO_312 (O_312,N_9884,N_9816);
xor UO_313 (O_313,N_9862,N_9911);
nor UO_314 (O_314,N_9847,N_9822);
nand UO_315 (O_315,N_9921,N_9889);
and UO_316 (O_316,N_9991,N_9969);
or UO_317 (O_317,N_9971,N_9891);
or UO_318 (O_318,N_9832,N_9841);
or UO_319 (O_319,N_9925,N_9997);
and UO_320 (O_320,N_9801,N_9875);
nor UO_321 (O_321,N_9842,N_9916);
or UO_322 (O_322,N_9805,N_9945);
or UO_323 (O_323,N_9923,N_9947);
nand UO_324 (O_324,N_9933,N_9942);
and UO_325 (O_325,N_9832,N_9967);
or UO_326 (O_326,N_9836,N_9908);
or UO_327 (O_327,N_9922,N_9919);
or UO_328 (O_328,N_9890,N_9876);
or UO_329 (O_329,N_9810,N_9926);
nand UO_330 (O_330,N_9979,N_9922);
or UO_331 (O_331,N_9837,N_9827);
nor UO_332 (O_332,N_9940,N_9821);
xor UO_333 (O_333,N_9881,N_9982);
or UO_334 (O_334,N_9821,N_9888);
nor UO_335 (O_335,N_9999,N_9884);
nor UO_336 (O_336,N_9823,N_9961);
and UO_337 (O_337,N_9875,N_9989);
or UO_338 (O_338,N_9825,N_9935);
and UO_339 (O_339,N_9891,N_9989);
or UO_340 (O_340,N_9983,N_9972);
nor UO_341 (O_341,N_9873,N_9899);
or UO_342 (O_342,N_9806,N_9898);
nor UO_343 (O_343,N_9910,N_9846);
and UO_344 (O_344,N_9819,N_9895);
and UO_345 (O_345,N_9902,N_9809);
or UO_346 (O_346,N_9843,N_9878);
nand UO_347 (O_347,N_9869,N_9914);
or UO_348 (O_348,N_9958,N_9983);
nor UO_349 (O_349,N_9993,N_9807);
nand UO_350 (O_350,N_9983,N_9874);
and UO_351 (O_351,N_9887,N_9820);
or UO_352 (O_352,N_9834,N_9892);
nor UO_353 (O_353,N_9983,N_9861);
nor UO_354 (O_354,N_9997,N_9836);
nor UO_355 (O_355,N_9938,N_9940);
and UO_356 (O_356,N_9944,N_9835);
nand UO_357 (O_357,N_9955,N_9954);
or UO_358 (O_358,N_9928,N_9819);
nand UO_359 (O_359,N_9960,N_9982);
nor UO_360 (O_360,N_9859,N_9824);
nor UO_361 (O_361,N_9825,N_9958);
and UO_362 (O_362,N_9813,N_9828);
nor UO_363 (O_363,N_9894,N_9992);
or UO_364 (O_364,N_9843,N_9960);
or UO_365 (O_365,N_9952,N_9817);
and UO_366 (O_366,N_9967,N_9880);
and UO_367 (O_367,N_9854,N_9857);
xor UO_368 (O_368,N_9850,N_9803);
and UO_369 (O_369,N_9849,N_9980);
nor UO_370 (O_370,N_9981,N_9857);
nand UO_371 (O_371,N_9966,N_9955);
or UO_372 (O_372,N_9841,N_9944);
or UO_373 (O_373,N_9817,N_9861);
and UO_374 (O_374,N_9941,N_9876);
nand UO_375 (O_375,N_9914,N_9841);
or UO_376 (O_376,N_9934,N_9920);
nor UO_377 (O_377,N_9951,N_9923);
nor UO_378 (O_378,N_9897,N_9937);
nor UO_379 (O_379,N_9848,N_9886);
nand UO_380 (O_380,N_9956,N_9965);
and UO_381 (O_381,N_9867,N_9848);
nand UO_382 (O_382,N_9942,N_9842);
nor UO_383 (O_383,N_9953,N_9837);
nand UO_384 (O_384,N_9857,N_9847);
or UO_385 (O_385,N_9975,N_9878);
or UO_386 (O_386,N_9931,N_9989);
nand UO_387 (O_387,N_9990,N_9898);
and UO_388 (O_388,N_9865,N_9940);
or UO_389 (O_389,N_9925,N_9999);
nand UO_390 (O_390,N_9860,N_9868);
or UO_391 (O_391,N_9892,N_9929);
nand UO_392 (O_392,N_9847,N_9920);
and UO_393 (O_393,N_9984,N_9952);
or UO_394 (O_394,N_9995,N_9901);
or UO_395 (O_395,N_9870,N_9980);
or UO_396 (O_396,N_9919,N_9998);
nor UO_397 (O_397,N_9961,N_9829);
or UO_398 (O_398,N_9928,N_9803);
nand UO_399 (O_399,N_9806,N_9988);
nor UO_400 (O_400,N_9966,N_9832);
nand UO_401 (O_401,N_9849,N_9858);
nand UO_402 (O_402,N_9842,N_9804);
and UO_403 (O_403,N_9874,N_9860);
and UO_404 (O_404,N_9934,N_9900);
nor UO_405 (O_405,N_9819,N_9834);
nand UO_406 (O_406,N_9869,N_9825);
or UO_407 (O_407,N_9955,N_9997);
or UO_408 (O_408,N_9880,N_9809);
and UO_409 (O_409,N_9800,N_9951);
or UO_410 (O_410,N_9941,N_9886);
and UO_411 (O_411,N_9911,N_9962);
nor UO_412 (O_412,N_9884,N_9838);
xnor UO_413 (O_413,N_9865,N_9821);
nor UO_414 (O_414,N_9823,N_9839);
or UO_415 (O_415,N_9867,N_9913);
or UO_416 (O_416,N_9849,N_9851);
or UO_417 (O_417,N_9941,N_9868);
and UO_418 (O_418,N_9954,N_9970);
nand UO_419 (O_419,N_9923,N_9901);
and UO_420 (O_420,N_9874,N_9934);
and UO_421 (O_421,N_9837,N_9889);
nor UO_422 (O_422,N_9905,N_9857);
nor UO_423 (O_423,N_9879,N_9802);
and UO_424 (O_424,N_9822,N_9856);
and UO_425 (O_425,N_9943,N_9986);
and UO_426 (O_426,N_9999,N_9957);
nor UO_427 (O_427,N_9998,N_9880);
nor UO_428 (O_428,N_9984,N_9956);
or UO_429 (O_429,N_9968,N_9936);
or UO_430 (O_430,N_9917,N_9812);
nand UO_431 (O_431,N_9829,N_9870);
nand UO_432 (O_432,N_9941,N_9997);
or UO_433 (O_433,N_9979,N_9849);
and UO_434 (O_434,N_9925,N_9958);
xnor UO_435 (O_435,N_9850,N_9818);
and UO_436 (O_436,N_9872,N_9853);
nor UO_437 (O_437,N_9957,N_9989);
or UO_438 (O_438,N_9928,N_9908);
and UO_439 (O_439,N_9923,N_9849);
or UO_440 (O_440,N_9850,N_9815);
and UO_441 (O_441,N_9871,N_9818);
nand UO_442 (O_442,N_9807,N_9874);
or UO_443 (O_443,N_9899,N_9874);
and UO_444 (O_444,N_9987,N_9831);
nand UO_445 (O_445,N_9902,N_9843);
and UO_446 (O_446,N_9945,N_9869);
nor UO_447 (O_447,N_9940,N_9979);
or UO_448 (O_448,N_9993,N_9803);
nand UO_449 (O_449,N_9808,N_9995);
or UO_450 (O_450,N_9955,N_9949);
or UO_451 (O_451,N_9901,N_9983);
or UO_452 (O_452,N_9887,N_9993);
or UO_453 (O_453,N_9871,N_9845);
xnor UO_454 (O_454,N_9893,N_9943);
or UO_455 (O_455,N_9985,N_9987);
nor UO_456 (O_456,N_9855,N_9877);
and UO_457 (O_457,N_9812,N_9995);
nor UO_458 (O_458,N_9947,N_9852);
nand UO_459 (O_459,N_9814,N_9891);
nand UO_460 (O_460,N_9805,N_9826);
and UO_461 (O_461,N_9833,N_9887);
or UO_462 (O_462,N_9880,N_9930);
xor UO_463 (O_463,N_9809,N_9992);
and UO_464 (O_464,N_9946,N_9952);
nor UO_465 (O_465,N_9811,N_9934);
and UO_466 (O_466,N_9888,N_9926);
and UO_467 (O_467,N_9930,N_9934);
nand UO_468 (O_468,N_9825,N_9988);
or UO_469 (O_469,N_9949,N_9944);
nor UO_470 (O_470,N_9914,N_9812);
and UO_471 (O_471,N_9896,N_9863);
or UO_472 (O_472,N_9972,N_9995);
or UO_473 (O_473,N_9924,N_9839);
or UO_474 (O_474,N_9941,N_9923);
and UO_475 (O_475,N_9900,N_9919);
or UO_476 (O_476,N_9871,N_9827);
and UO_477 (O_477,N_9858,N_9801);
nand UO_478 (O_478,N_9831,N_9971);
nor UO_479 (O_479,N_9868,N_9965);
nand UO_480 (O_480,N_9912,N_9952);
and UO_481 (O_481,N_9838,N_9890);
and UO_482 (O_482,N_9974,N_9943);
nor UO_483 (O_483,N_9952,N_9937);
and UO_484 (O_484,N_9986,N_9815);
and UO_485 (O_485,N_9974,N_9884);
and UO_486 (O_486,N_9976,N_9998);
nor UO_487 (O_487,N_9956,N_9961);
nor UO_488 (O_488,N_9919,N_9880);
and UO_489 (O_489,N_9903,N_9814);
nor UO_490 (O_490,N_9844,N_9859);
nand UO_491 (O_491,N_9915,N_9962);
and UO_492 (O_492,N_9924,N_9998);
or UO_493 (O_493,N_9974,N_9830);
nor UO_494 (O_494,N_9817,N_9836);
and UO_495 (O_495,N_9842,N_9801);
or UO_496 (O_496,N_9956,N_9889);
nand UO_497 (O_497,N_9919,N_9938);
nand UO_498 (O_498,N_9869,N_9929);
nor UO_499 (O_499,N_9970,N_9857);
and UO_500 (O_500,N_9885,N_9916);
or UO_501 (O_501,N_9800,N_9868);
nand UO_502 (O_502,N_9984,N_9949);
nand UO_503 (O_503,N_9862,N_9857);
or UO_504 (O_504,N_9817,N_9876);
nand UO_505 (O_505,N_9855,N_9923);
nand UO_506 (O_506,N_9889,N_9940);
or UO_507 (O_507,N_9959,N_9932);
nand UO_508 (O_508,N_9975,N_9991);
nor UO_509 (O_509,N_9967,N_9893);
nor UO_510 (O_510,N_9955,N_9800);
and UO_511 (O_511,N_9862,N_9878);
nand UO_512 (O_512,N_9941,N_9883);
xnor UO_513 (O_513,N_9941,N_9994);
or UO_514 (O_514,N_9885,N_9811);
and UO_515 (O_515,N_9989,N_9956);
and UO_516 (O_516,N_9827,N_9987);
nor UO_517 (O_517,N_9886,N_9991);
or UO_518 (O_518,N_9946,N_9972);
xor UO_519 (O_519,N_9854,N_9917);
or UO_520 (O_520,N_9862,N_9821);
or UO_521 (O_521,N_9813,N_9809);
nor UO_522 (O_522,N_9836,N_9850);
nor UO_523 (O_523,N_9865,N_9833);
or UO_524 (O_524,N_9873,N_9993);
nand UO_525 (O_525,N_9911,N_9831);
or UO_526 (O_526,N_9968,N_9926);
nand UO_527 (O_527,N_9942,N_9808);
nand UO_528 (O_528,N_9822,N_9800);
or UO_529 (O_529,N_9817,N_9825);
or UO_530 (O_530,N_9947,N_9936);
nor UO_531 (O_531,N_9800,N_9999);
and UO_532 (O_532,N_9972,N_9951);
and UO_533 (O_533,N_9820,N_9941);
nand UO_534 (O_534,N_9941,N_9882);
nor UO_535 (O_535,N_9895,N_9944);
nor UO_536 (O_536,N_9945,N_9991);
or UO_537 (O_537,N_9959,N_9803);
or UO_538 (O_538,N_9825,N_9924);
xor UO_539 (O_539,N_9957,N_9896);
nand UO_540 (O_540,N_9864,N_9906);
nor UO_541 (O_541,N_9830,N_9823);
and UO_542 (O_542,N_9813,N_9939);
nor UO_543 (O_543,N_9800,N_9801);
or UO_544 (O_544,N_9944,N_9935);
and UO_545 (O_545,N_9804,N_9929);
or UO_546 (O_546,N_9819,N_9858);
nor UO_547 (O_547,N_9878,N_9833);
nand UO_548 (O_548,N_9880,N_9924);
and UO_549 (O_549,N_9916,N_9866);
or UO_550 (O_550,N_9971,N_9983);
nor UO_551 (O_551,N_9830,N_9844);
and UO_552 (O_552,N_9979,N_9851);
or UO_553 (O_553,N_9834,N_9808);
or UO_554 (O_554,N_9928,N_9989);
or UO_555 (O_555,N_9833,N_9930);
nor UO_556 (O_556,N_9849,N_9892);
or UO_557 (O_557,N_9964,N_9956);
and UO_558 (O_558,N_9830,N_9908);
xnor UO_559 (O_559,N_9958,N_9984);
and UO_560 (O_560,N_9963,N_9934);
or UO_561 (O_561,N_9802,N_9966);
nand UO_562 (O_562,N_9950,N_9857);
and UO_563 (O_563,N_9828,N_9802);
and UO_564 (O_564,N_9975,N_9885);
nor UO_565 (O_565,N_9828,N_9946);
nor UO_566 (O_566,N_9968,N_9993);
and UO_567 (O_567,N_9827,N_9916);
or UO_568 (O_568,N_9826,N_9960);
nand UO_569 (O_569,N_9833,N_9913);
nand UO_570 (O_570,N_9932,N_9832);
nand UO_571 (O_571,N_9960,N_9993);
or UO_572 (O_572,N_9996,N_9847);
and UO_573 (O_573,N_9864,N_9877);
nand UO_574 (O_574,N_9814,N_9973);
nand UO_575 (O_575,N_9910,N_9946);
and UO_576 (O_576,N_9896,N_9837);
or UO_577 (O_577,N_9837,N_9818);
nor UO_578 (O_578,N_9898,N_9989);
nor UO_579 (O_579,N_9844,N_9956);
nand UO_580 (O_580,N_9996,N_9932);
and UO_581 (O_581,N_9815,N_9823);
or UO_582 (O_582,N_9878,N_9972);
nand UO_583 (O_583,N_9918,N_9964);
and UO_584 (O_584,N_9803,N_9830);
xor UO_585 (O_585,N_9871,N_9883);
or UO_586 (O_586,N_9835,N_9918);
nand UO_587 (O_587,N_9926,N_9805);
and UO_588 (O_588,N_9980,N_9806);
nor UO_589 (O_589,N_9858,N_9936);
nor UO_590 (O_590,N_9869,N_9981);
and UO_591 (O_591,N_9929,N_9896);
or UO_592 (O_592,N_9843,N_9907);
nand UO_593 (O_593,N_9991,N_9866);
and UO_594 (O_594,N_9887,N_9856);
nor UO_595 (O_595,N_9857,N_9815);
nand UO_596 (O_596,N_9804,N_9833);
and UO_597 (O_597,N_9837,N_9864);
nand UO_598 (O_598,N_9821,N_9960);
or UO_599 (O_599,N_9831,N_9849);
nand UO_600 (O_600,N_9999,N_9995);
and UO_601 (O_601,N_9899,N_9863);
nand UO_602 (O_602,N_9883,N_9913);
or UO_603 (O_603,N_9883,N_9926);
nor UO_604 (O_604,N_9994,N_9814);
nand UO_605 (O_605,N_9901,N_9985);
nand UO_606 (O_606,N_9911,N_9923);
nor UO_607 (O_607,N_9873,N_9889);
nand UO_608 (O_608,N_9958,N_9932);
nor UO_609 (O_609,N_9989,N_9930);
nor UO_610 (O_610,N_9943,N_9931);
nand UO_611 (O_611,N_9961,N_9998);
and UO_612 (O_612,N_9928,N_9932);
or UO_613 (O_613,N_9885,N_9801);
or UO_614 (O_614,N_9885,N_9873);
nand UO_615 (O_615,N_9825,N_9802);
nand UO_616 (O_616,N_9845,N_9997);
or UO_617 (O_617,N_9960,N_9895);
xor UO_618 (O_618,N_9985,N_9993);
xor UO_619 (O_619,N_9936,N_9893);
nor UO_620 (O_620,N_9943,N_9975);
nand UO_621 (O_621,N_9957,N_9816);
nand UO_622 (O_622,N_9803,N_9909);
nor UO_623 (O_623,N_9979,N_9928);
nor UO_624 (O_624,N_9947,N_9935);
or UO_625 (O_625,N_9906,N_9903);
nand UO_626 (O_626,N_9989,N_9883);
or UO_627 (O_627,N_9939,N_9909);
nand UO_628 (O_628,N_9820,N_9991);
or UO_629 (O_629,N_9896,N_9931);
and UO_630 (O_630,N_9903,N_9860);
nand UO_631 (O_631,N_9928,N_9905);
or UO_632 (O_632,N_9804,N_9900);
nor UO_633 (O_633,N_9988,N_9866);
nor UO_634 (O_634,N_9852,N_9877);
nor UO_635 (O_635,N_9886,N_9832);
nand UO_636 (O_636,N_9830,N_9834);
or UO_637 (O_637,N_9867,N_9878);
or UO_638 (O_638,N_9900,N_9925);
and UO_639 (O_639,N_9848,N_9858);
or UO_640 (O_640,N_9971,N_9937);
nand UO_641 (O_641,N_9829,N_9931);
and UO_642 (O_642,N_9983,N_9826);
or UO_643 (O_643,N_9908,N_9801);
or UO_644 (O_644,N_9864,N_9996);
and UO_645 (O_645,N_9865,N_9904);
nand UO_646 (O_646,N_9925,N_9991);
or UO_647 (O_647,N_9998,N_9946);
and UO_648 (O_648,N_9849,N_9857);
nor UO_649 (O_649,N_9983,N_9912);
nand UO_650 (O_650,N_9936,N_9828);
or UO_651 (O_651,N_9905,N_9910);
or UO_652 (O_652,N_9959,N_9867);
nand UO_653 (O_653,N_9881,N_9841);
nand UO_654 (O_654,N_9968,N_9848);
and UO_655 (O_655,N_9949,N_9923);
nor UO_656 (O_656,N_9972,N_9877);
or UO_657 (O_657,N_9864,N_9831);
nand UO_658 (O_658,N_9881,N_9803);
nor UO_659 (O_659,N_9933,N_9802);
nand UO_660 (O_660,N_9942,N_9965);
or UO_661 (O_661,N_9806,N_9885);
and UO_662 (O_662,N_9843,N_9951);
nand UO_663 (O_663,N_9999,N_9852);
nor UO_664 (O_664,N_9869,N_9897);
nor UO_665 (O_665,N_9996,N_9955);
and UO_666 (O_666,N_9893,N_9827);
nor UO_667 (O_667,N_9806,N_9873);
and UO_668 (O_668,N_9997,N_9957);
nand UO_669 (O_669,N_9925,N_9980);
nor UO_670 (O_670,N_9810,N_9866);
or UO_671 (O_671,N_9871,N_9936);
or UO_672 (O_672,N_9803,N_9839);
and UO_673 (O_673,N_9804,N_9899);
and UO_674 (O_674,N_9863,N_9885);
and UO_675 (O_675,N_9905,N_9963);
or UO_676 (O_676,N_9932,N_9893);
nor UO_677 (O_677,N_9951,N_9967);
and UO_678 (O_678,N_9828,N_9990);
nor UO_679 (O_679,N_9805,N_9856);
nand UO_680 (O_680,N_9818,N_9817);
nor UO_681 (O_681,N_9956,N_9913);
nand UO_682 (O_682,N_9953,N_9900);
and UO_683 (O_683,N_9865,N_9923);
and UO_684 (O_684,N_9882,N_9928);
or UO_685 (O_685,N_9834,N_9951);
or UO_686 (O_686,N_9833,N_9937);
or UO_687 (O_687,N_9810,N_9869);
nor UO_688 (O_688,N_9822,N_9898);
or UO_689 (O_689,N_9830,N_9954);
nand UO_690 (O_690,N_9867,N_9876);
or UO_691 (O_691,N_9880,N_9938);
nand UO_692 (O_692,N_9812,N_9908);
nor UO_693 (O_693,N_9854,N_9816);
or UO_694 (O_694,N_9984,N_9933);
nor UO_695 (O_695,N_9882,N_9847);
and UO_696 (O_696,N_9835,N_9899);
nand UO_697 (O_697,N_9966,N_9891);
and UO_698 (O_698,N_9864,N_9959);
or UO_699 (O_699,N_9922,N_9915);
nor UO_700 (O_700,N_9932,N_9927);
and UO_701 (O_701,N_9889,N_9899);
and UO_702 (O_702,N_9838,N_9854);
and UO_703 (O_703,N_9899,N_9955);
or UO_704 (O_704,N_9836,N_9925);
and UO_705 (O_705,N_9861,N_9804);
nand UO_706 (O_706,N_9861,N_9844);
xor UO_707 (O_707,N_9882,N_9978);
nor UO_708 (O_708,N_9939,N_9802);
and UO_709 (O_709,N_9969,N_9908);
and UO_710 (O_710,N_9949,N_9893);
nor UO_711 (O_711,N_9909,N_9960);
and UO_712 (O_712,N_9887,N_9957);
and UO_713 (O_713,N_9834,N_9860);
nor UO_714 (O_714,N_9905,N_9931);
and UO_715 (O_715,N_9924,N_9847);
nand UO_716 (O_716,N_9895,N_9890);
nand UO_717 (O_717,N_9845,N_9978);
nor UO_718 (O_718,N_9889,N_9957);
and UO_719 (O_719,N_9920,N_9964);
xnor UO_720 (O_720,N_9802,N_9868);
nand UO_721 (O_721,N_9929,N_9842);
nand UO_722 (O_722,N_9984,N_9858);
or UO_723 (O_723,N_9821,N_9813);
nor UO_724 (O_724,N_9987,N_9837);
or UO_725 (O_725,N_9886,N_9987);
nand UO_726 (O_726,N_9835,N_9982);
or UO_727 (O_727,N_9939,N_9821);
nor UO_728 (O_728,N_9934,N_9895);
nand UO_729 (O_729,N_9991,N_9973);
nand UO_730 (O_730,N_9957,N_9879);
or UO_731 (O_731,N_9841,N_9912);
nor UO_732 (O_732,N_9936,N_9970);
nor UO_733 (O_733,N_9870,N_9887);
and UO_734 (O_734,N_9837,N_9990);
nor UO_735 (O_735,N_9814,N_9849);
and UO_736 (O_736,N_9919,N_9962);
or UO_737 (O_737,N_9944,N_9891);
nand UO_738 (O_738,N_9927,N_9934);
or UO_739 (O_739,N_9841,N_9975);
nor UO_740 (O_740,N_9865,N_9899);
and UO_741 (O_741,N_9874,N_9943);
and UO_742 (O_742,N_9867,N_9995);
xnor UO_743 (O_743,N_9858,N_9892);
or UO_744 (O_744,N_9917,N_9901);
nor UO_745 (O_745,N_9996,N_9892);
nor UO_746 (O_746,N_9869,N_9802);
or UO_747 (O_747,N_9860,N_9839);
nand UO_748 (O_748,N_9906,N_9943);
and UO_749 (O_749,N_9831,N_9814);
and UO_750 (O_750,N_9957,N_9865);
and UO_751 (O_751,N_9894,N_9936);
nand UO_752 (O_752,N_9882,N_9833);
nand UO_753 (O_753,N_9800,N_9898);
nor UO_754 (O_754,N_9992,N_9895);
and UO_755 (O_755,N_9897,N_9881);
nor UO_756 (O_756,N_9868,N_9859);
nor UO_757 (O_757,N_9950,N_9832);
nand UO_758 (O_758,N_9819,N_9999);
or UO_759 (O_759,N_9995,N_9843);
and UO_760 (O_760,N_9871,N_9875);
or UO_761 (O_761,N_9819,N_9931);
nand UO_762 (O_762,N_9882,N_9889);
and UO_763 (O_763,N_9819,N_9974);
nand UO_764 (O_764,N_9953,N_9832);
or UO_765 (O_765,N_9870,N_9988);
nor UO_766 (O_766,N_9951,N_9919);
and UO_767 (O_767,N_9990,N_9859);
or UO_768 (O_768,N_9973,N_9912);
or UO_769 (O_769,N_9959,N_9886);
nor UO_770 (O_770,N_9890,N_9894);
and UO_771 (O_771,N_9939,N_9967);
and UO_772 (O_772,N_9911,N_9929);
nand UO_773 (O_773,N_9988,N_9840);
nor UO_774 (O_774,N_9933,N_9871);
and UO_775 (O_775,N_9872,N_9843);
and UO_776 (O_776,N_9962,N_9858);
nand UO_777 (O_777,N_9840,N_9908);
nand UO_778 (O_778,N_9888,N_9859);
nor UO_779 (O_779,N_9844,N_9870);
and UO_780 (O_780,N_9837,N_9989);
nand UO_781 (O_781,N_9832,N_9995);
nor UO_782 (O_782,N_9981,N_9982);
or UO_783 (O_783,N_9995,N_9980);
nand UO_784 (O_784,N_9911,N_9936);
and UO_785 (O_785,N_9959,N_9968);
and UO_786 (O_786,N_9908,N_9809);
and UO_787 (O_787,N_9884,N_9953);
and UO_788 (O_788,N_9979,N_9886);
nor UO_789 (O_789,N_9992,N_9936);
or UO_790 (O_790,N_9804,N_9967);
nor UO_791 (O_791,N_9819,N_9838);
nor UO_792 (O_792,N_9875,N_9810);
or UO_793 (O_793,N_9952,N_9813);
and UO_794 (O_794,N_9997,N_9989);
nand UO_795 (O_795,N_9886,N_9950);
and UO_796 (O_796,N_9836,N_9806);
xnor UO_797 (O_797,N_9849,N_9802);
or UO_798 (O_798,N_9814,N_9860);
nor UO_799 (O_799,N_9904,N_9820);
nand UO_800 (O_800,N_9932,N_9864);
nand UO_801 (O_801,N_9805,N_9949);
or UO_802 (O_802,N_9958,N_9951);
nand UO_803 (O_803,N_9885,N_9838);
nand UO_804 (O_804,N_9961,N_9876);
and UO_805 (O_805,N_9933,N_9853);
and UO_806 (O_806,N_9910,N_9864);
and UO_807 (O_807,N_9870,N_9916);
or UO_808 (O_808,N_9894,N_9843);
nand UO_809 (O_809,N_9999,N_9941);
nor UO_810 (O_810,N_9985,N_9910);
or UO_811 (O_811,N_9915,N_9806);
nor UO_812 (O_812,N_9933,N_9930);
nor UO_813 (O_813,N_9924,N_9896);
and UO_814 (O_814,N_9996,N_9843);
nor UO_815 (O_815,N_9835,N_9814);
nor UO_816 (O_816,N_9811,N_9825);
and UO_817 (O_817,N_9820,N_9816);
and UO_818 (O_818,N_9944,N_9862);
or UO_819 (O_819,N_9896,N_9840);
nor UO_820 (O_820,N_9887,N_9939);
or UO_821 (O_821,N_9910,N_9802);
nor UO_822 (O_822,N_9888,N_9923);
and UO_823 (O_823,N_9855,N_9859);
or UO_824 (O_824,N_9858,N_9976);
or UO_825 (O_825,N_9847,N_9861);
nand UO_826 (O_826,N_9913,N_9879);
or UO_827 (O_827,N_9838,N_9965);
nand UO_828 (O_828,N_9836,N_9823);
nor UO_829 (O_829,N_9941,N_9946);
nand UO_830 (O_830,N_9812,N_9898);
nor UO_831 (O_831,N_9957,N_9948);
nor UO_832 (O_832,N_9881,N_9957);
nand UO_833 (O_833,N_9951,N_9860);
nor UO_834 (O_834,N_9905,N_9952);
and UO_835 (O_835,N_9846,N_9800);
or UO_836 (O_836,N_9831,N_9800);
nor UO_837 (O_837,N_9882,N_9910);
or UO_838 (O_838,N_9872,N_9940);
nor UO_839 (O_839,N_9874,N_9901);
nand UO_840 (O_840,N_9833,N_9809);
and UO_841 (O_841,N_9916,N_9928);
or UO_842 (O_842,N_9993,N_9920);
nor UO_843 (O_843,N_9945,N_9986);
and UO_844 (O_844,N_9822,N_9903);
nand UO_845 (O_845,N_9922,N_9868);
or UO_846 (O_846,N_9824,N_9853);
nor UO_847 (O_847,N_9899,N_9842);
nor UO_848 (O_848,N_9961,N_9983);
nand UO_849 (O_849,N_9958,N_9933);
and UO_850 (O_850,N_9838,N_9989);
nor UO_851 (O_851,N_9878,N_9872);
or UO_852 (O_852,N_9802,N_9979);
nand UO_853 (O_853,N_9810,N_9986);
nand UO_854 (O_854,N_9946,N_9951);
nor UO_855 (O_855,N_9872,N_9860);
nor UO_856 (O_856,N_9956,N_9812);
nor UO_857 (O_857,N_9859,N_9901);
xor UO_858 (O_858,N_9957,N_9819);
nand UO_859 (O_859,N_9950,N_9834);
or UO_860 (O_860,N_9965,N_9904);
nand UO_861 (O_861,N_9991,N_9894);
and UO_862 (O_862,N_9870,N_9981);
or UO_863 (O_863,N_9948,N_9908);
nor UO_864 (O_864,N_9854,N_9904);
and UO_865 (O_865,N_9959,N_9920);
and UO_866 (O_866,N_9978,N_9926);
nand UO_867 (O_867,N_9861,N_9913);
and UO_868 (O_868,N_9851,N_9820);
and UO_869 (O_869,N_9806,N_9829);
and UO_870 (O_870,N_9933,N_9869);
or UO_871 (O_871,N_9972,N_9892);
nor UO_872 (O_872,N_9928,N_9896);
nand UO_873 (O_873,N_9826,N_9866);
or UO_874 (O_874,N_9920,N_9832);
nand UO_875 (O_875,N_9871,N_9917);
and UO_876 (O_876,N_9830,N_9973);
nand UO_877 (O_877,N_9924,N_9985);
or UO_878 (O_878,N_9951,N_9982);
nand UO_879 (O_879,N_9998,N_9905);
nand UO_880 (O_880,N_9892,N_9814);
xor UO_881 (O_881,N_9813,N_9941);
and UO_882 (O_882,N_9940,N_9869);
and UO_883 (O_883,N_9868,N_9820);
nor UO_884 (O_884,N_9936,N_9940);
or UO_885 (O_885,N_9866,N_9987);
or UO_886 (O_886,N_9876,N_9933);
nand UO_887 (O_887,N_9932,N_9985);
or UO_888 (O_888,N_9887,N_9879);
and UO_889 (O_889,N_9966,N_9905);
or UO_890 (O_890,N_9962,N_9801);
or UO_891 (O_891,N_9986,N_9850);
nor UO_892 (O_892,N_9922,N_9800);
nor UO_893 (O_893,N_9912,N_9911);
or UO_894 (O_894,N_9942,N_9995);
nor UO_895 (O_895,N_9991,N_9942);
nand UO_896 (O_896,N_9904,N_9915);
nor UO_897 (O_897,N_9952,N_9866);
and UO_898 (O_898,N_9804,N_9823);
and UO_899 (O_899,N_9821,N_9907);
nor UO_900 (O_900,N_9866,N_9847);
nand UO_901 (O_901,N_9917,N_9820);
nor UO_902 (O_902,N_9901,N_9857);
or UO_903 (O_903,N_9935,N_9994);
nor UO_904 (O_904,N_9897,N_9834);
and UO_905 (O_905,N_9840,N_9990);
nand UO_906 (O_906,N_9948,N_9967);
or UO_907 (O_907,N_9954,N_9994);
or UO_908 (O_908,N_9923,N_9817);
and UO_909 (O_909,N_9807,N_9946);
nand UO_910 (O_910,N_9805,N_9934);
nor UO_911 (O_911,N_9964,N_9952);
and UO_912 (O_912,N_9804,N_9864);
and UO_913 (O_913,N_9842,N_9881);
nand UO_914 (O_914,N_9806,N_9962);
and UO_915 (O_915,N_9821,N_9913);
nor UO_916 (O_916,N_9964,N_9951);
or UO_917 (O_917,N_9815,N_9830);
and UO_918 (O_918,N_9997,N_9911);
or UO_919 (O_919,N_9981,N_9935);
nor UO_920 (O_920,N_9841,N_9947);
nand UO_921 (O_921,N_9876,N_9839);
and UO_922 (O_922,N_9932,N_9909);
or UO_923 (O_923,N_9822,N_9817);
nor UO_924 (O_924,N_9924,N_9877);
or UO_925 (O_925,N_9985,N_9966);
nand UO_926 (O_926,N_9815,N_9940);
nand UO_927 (O_927,N_9928,N_9912);
nand UO_928 (O_928,N_9900,N_9856);
or UO_929 (O_929,N_9870,N_9815);
xnor UO_930 (O_930,N_9881,N_9997);
or UO_931 (O_931,N_9808,N_9873);
nor UO_932 (O_932,N_9825,N_9930);
nor UO_933 (O_933,N_9810,N_9865);
nor UO_934 (O_934,N_9825,N_9912);
and UO_935 (O_935,N_9841,N_9970);
and UO_936 (O_936,N_9981,N_9901);
or UO_937 (O_937,N_9930,N_9907);
nor UO_938 (O_938,N_9807,N_9937);
nand UO_939 (O_939,N_9885,N_9953);
and UO_940 (O_940,N_9896,N_9997);
nand UO_941 (O_941,N_9826,N_9929);
nor UO_942 (O_942,N_9837,N_9895);
or UO_943 (O_943,N_9888,N_9881);
and UO_944 (O_944,N_9849,N_9950);
nand UO_945 (O_945,N_9887,N_9889);
or UO_946 (O_946,N_9850,N_9823);
nand UO_947 (O_947,N_9863,N_9806);
nand UO_948 (O_948,N_9838,N_9836);
nand UO_949 (O_949,N_9994,N_9914);
nand UO_950 (O_950,N_9824,N_9857);
or UO_951 (O_951,N_9840,N_9946);
xor UO_952 (O_952,N_9941,N_9810);
or UO_953 (O_953,N_9802,N_9985);
nor UO_954 (O_954,N_9968,N_9852);
nand UO_955 (O_955,N_9933,N_9962);
nand UO_956 (O_956,N_9814,N_9921);
and UO_957 (O_957,N_9901,N_9816);
and UO_958 (O_958,N_9837,N_9801);
nand UO_959 (O_959,N_9984,N_9813);
or UO_960 (O_960,N_9915,N_9985);
nor UO_961 (O_961,N_9975,N_9868);
xor UO_962 (O_962,N_9900,N_9950);
and UO_963 (O_963,N_9876,N_9930);
nor UO_964 (O_964,N_9832,N_9859);
and UO_965 (O_965,N_9870,N_9955);
nand UO_966 (O_966,N_9869,N_9827);
xor UO_967 (O_967,N_9823,N_9930);
or UO_968 (O_968,N_9934,N_9819);
and UO_969 (O_969,N_9810,N_9888);
nand UO_970 (O_970,N_9943,N_9843);
or UO_971 (O_971,N_9892,N_9853);
and UO_972 (O_972,N_9991,N_9801);
nand UO_973 (O_973,N_9925,N_9975);
nand UO_974 (O_974,N_9800,N_9921);
and UO_975 (O_975,N_9983,N_9889);
nand UO_976 (O_976,N_9912,N_9804);
nand UO_977 (O_977,N_9953,N_9940);
nor UO_978 (O_978,N_9929,N_9980);
and UO_979 (O_979,N_9825,N_9933);
nor UO_980 (O_980,N_9938,N_9854);
nand UO_981 (O_981,N_9894,N_9870);
nor UO_982 (O_982,N_9852,N_9977);
xnor UO_983 (O_983,N_9935,N_9964);
nand UO_984 (O_984,N_9829,N_9943);
and UO_985 (O_985,N_9813,N_9991);
nor UO_986 (O_986,N_9986,N_9831);
nor UO_987 (O_987,N_9945,N_9872);
nand UO_988 (O_988,N_9948,N_9916);
nand UO_989 (O_989,N_9973,N_9834);
nor UO_990 (O_990,N_9949,N_9958);
or UO_991 (O_991,N_9840,N_9897);
and UO_992 (O_992,N_9843,N_9858);
nor UO_993 (O_993,N_9874,N_9954);
or UO_994 (O_994,N_9934,N_9923);
and UO_995 (O_995,N_9900,N_9926);
nand UO_996 (O_996,N_9831,N_9833);
nand UO_997 (O_997,N_9942,N_9987);
nor UO_998 (O_998,N_9932,N_9994);
nand UO_999 (O_999,N_9994,N_9995);
or UO_1000 (O_1000,N_9904,N_9835);
or UO_1001 (O_1001,N_9975,N_9825);
nor UO_1002 (O_1002,N_9995,N_9903);
nor UO_1003 (O_1003,N_9800,N_9860);
nand UO_1004 (O_1004,N_9956,N_9803);
nand UO_1005 (O_1005,N_9914,N_9881);
nor UO_1006 (O_1006,N_9862,N_9892);
nor UO_1007 (O_1007,N_9801,N_9916);
and UO_1008 (O_1008,N_9963,N_9816);
or UO_1009 (O_1009,N_9853,N_9855);
or UO_1010 (O_1010,N_9963,N_9935);
nand UO_1011 (O_1011,N_9980,N_9964);
nand UO_1012 (O_1012,N_9909,N_9868);
nand UO_1013 (O_1013,N_9904,N_9878);
nor UO_1014 (O_1014,N_9968,N_9983);
and UO_1015 (O_1015,N_9910,N_9831);
or UO_1016 (O_1016,N_9911,N_9930);
or UO_1017 (O_1017,N_9916,N_9867);
or UO_1018 (O_1018,N_9895,N_9897);
nand UO_1019 (O_1019,N_9855,N_9947);
nand UO_1020 (O_1020,N_9922,N_9891);
or UO_1021 (O_1021,N_9801,N_9845);
nor UO_1022 (O_1022,N_9835,N_9974);
or UO_1023 (O_1023,N_9818,N_9963);
nor UO_1024 (O_1024,N_9989,N_9809);
and UO_1025 (O_1025,N_9963,N_9849);
and UO_1026 (O_1026,N_9906,N_9921);
nor UO_1027 (O_1027,N_9881,N_9929);
and UO_1028 (O_1028,N_9921,N_9849);
and UO_1029 (O_1029,N_9928,N_9874);
or UO_1030 (O_1030,N_9982,N_9940);
and UO_1031 (O_1031,N_9845,N_9847);
nor UO_1032 (O_1032,N_9986,N_9930);
nand UO_1033 (O_1033,N_9836,N_9956);
and UO_1034 (O_1034,N_9926,N_9849);
and UO_1035 (O_1035,N_9818,N_9951);
nor UO_1036 (O_1036,N_9920,N_9823);
nand UO_1037 (O_1037,N_9827,N_9838);
or UO_1038 (O_1038,N_9998,N_9830);
nor UO_1039 (O_1039,N_9804,N_9860);
or UO_1040 (O_1040,N_9967,N_9844);
nand UO_1041 (O_1041,N_9834,N_9995);
nor UO_1042 (O_1042,N_9961,N_9923);
xnor UO_1043 (O_1043,N_9885,N_9850);
nand UO_1044 (O_1044,N_9887,N_9936);
or UO_1045 (O_1045,N_9979,N_9910);
and UO_1046 (O_1046,N_9833,N_9916);
nand UO_1047 (O_1047,N_9936,N_9852);
nor UO_1048 (O_1048,N_9984,N_9898);
and UO_1049 (O_1049,N_9908,N_9803);
nor UO_1050 (O_1050,N_9930,N_9938);
and UO_1051 (O_1051,N_9895,N_9974);
or UO_1052 (O_1052,N_9990,N_9833);
nand UO_1053 (O_1053,N_9876,N_9842);
nor UO_1054 (O_1054,N_9994,N_9879);
and UO_1055 (O_1055,N_9939,N_9870);
and UO_1056 (O_1056,N_9916,N_9950);
and UO_1057 (O_1057,N_9987,N_9848);
or UO_1058 (O_1058,N_9940,N_9891);
or UO_1059 (O_1059,N_9869,N_9805);
nor UO_1060 (O_1060,N_9886,N_9985);
and UO_1061 (O_1061,N_9968,N_9896);
nand UO_1062 (O_1062,N_9980,N_9974);
and UO_1063 (O_1063,N_9938,N_9942);
nand UO_1064 (O_1064,N_9884,N_9878);
nand UO_1065 (O_1065,N_9920,N_9908);
or UO_1066 (O_1066,N_9890,N_9981);
nor UO_1067 (O_1067,N_9869,N_9955);
nand UO_1068 (O_1068,N_9983,N_9934);
and UO_1069 (O_1069,N_9811,N_9923);
nor UO_1070 (O_1070,N_9816,N_9903);
nand UO_1071 (O_1071,N_9930,N_9870);
nor UO_1072 (O_1072,N_9858,N_9891);
or UO_1073 (O_1073,N_9948,N_9839);
nor UO_1074 (O_1074,N_9966,N_9995);
or UO_1075 (O_1075,N_9948,N_9808);
xnor UO_1076 (O_1076,N_9934,N_9998);
nor UO_1077 (O_1077,N_9891,N_9975);
or UO_1078 (O_1078,N_9853,N_9936);
nor UO_1079 (O_1079,N_9830,N_9924);
or UO_1080 (O_1080,N_9936,N_9827);
and UO_1081 (O_1081,N_9902,N_9983);
or UO_1082 (O_1082,N_9815,N_9871);
xnor UO_1083 (O_1083,N_9878,N_9999);
nor UO_1084 (O_1084,N_9812,N_9934);
nor UO_1085 (O_1085,N_9863,N_9941);
nand UO_1086 (O_1086,N_9823,N_9828);
nor UO_1087 (O_1087,N_9984,N_9831);
nand UO_1088 (O_1088,N_9936,N_9988);
nand UO_1089 (O_1089,N_9980,N_9976);
nand UO_1090 (O_1090,N_9845,N_9951);
and UO_1091 (O_1091,N_9942,N_9968);
nand UO_1092 (O_1092,N_9906,N_9852);
nand UO_1093 (O_1093,N_9963,N_9874);
or UO_1094 (O_1094,N_9843,N_9835);
nor UO_1095 (O_1095,N_9812,N_9855);
nand UO_1096 (O_1096,N_9914,N_9906);
or UO_1097 (O_1097,N_9864,N_9872);
nand UO_1098 (O_1098,N_9811,N_9977);
nand UO_1099 (O_1099,N_9844,N_9917);
and UO_1100 (O_1100,N_9913,N_9839);
and UO_1101 (O_1101,N_9957,N_9939);
and UO_1102 (O_1102,N_9960,N_9904);
or UO_1103 (O_1103,N_9872,N_9806);
nand UO_1104 (O_1104,N_9953,N_9976);
nor UO_1105 (O_1105,N_9984,N_9884);
or UO_1106 (O_1106,N_9901,N_9829);
and UO_1107 (O_1107,N_9989,N_9848);
and UO_1108 (O_1108,N_9971,N_9805);
or UO_1109 (O_1109,N_9929,N_9807);
nand UO_1110 (O_1110,N_9973,N_9887);
nor UO_1111 (O_1111,N_9907,N_9835);
nor UO_1112 (O_1112,N_9867,N_9940);
and UO_1113 (O_1113,N_9989,N_9984);
nor UO_1114 (O_1114,N_9829,N_9882);
nand UO_1115 (O_1115,N_9825,N_9830);
xor UO_1116 (O_1116,N_9902,N_9964);
and UO_1117 (O_1117,N_9982,N_9814);
nand UO_1118 (O_1118,N_9947,N_9884);
or UO_1119 (O_1119,N_9935,N_9911);
or UO_1120 (O_1120,N_9891,N_9825);
nand UO_1121 (O_1121,N_9936,N_9833);
and UO_1122 (O_1122,N_9833,N_9822);
nor UO_1123 (O_1123,N_9981,N_9875);
nand UO_1124 (O_1124,N_9937,N_9875);
nor UO_1125 (O_1125,N_9823,N_9912);
and UO_1126 (O_1126,N_9972,N_9976);
or UO_1127 (O_1127,N_9866,N_9807);
nor UO_1128 (O_1128,N_9867,N_9899);
nor UO_1129 (O_1129,N_9866,N_9823);
nor UO_1130 (O_1130,N_9972,N_9829);
and UO_1131 (O_1131,N_9868,N_9930);
or UO_1132 (O_1132,N_9841,N_9811);
nand UO_1133 (O_1133,N_9858,N_9878);
nor UO_1134 (O_1134,N_9856,N_9884);
or UO_1135 (O_1135,N_9935,N_9921);
and UO_1136 (O_1136,N_9918,N_9929);
nor UO_1137 (O_1137,N_9958,N_9959);
or UO_1138 (O_1138,N_9973,N_9923);
nand UO_1139 (O_1139,N_9883,N_9997);
and UO_1140 (O_1140,N_9996,N_9874);
nor UO_1141 (O_1141,N_9818,N_9833);
nand UO_1142 (O_1142,N_9912,N_9811);
or UO_1143 (O_1143,N_9829,N_9835);
nand UO_1144 (O_1144,N_9974,N_9801);
nand UO_1145 (O_1145,N_9999,N_9972);
nor UO_1146 (O_1146,N_9976,N_9821);
nor UO_1147 (O_1147,N_9925,N_9963);
nor UO_1148 (O_1148,N_9901,N_9975);
or UO_1149 (O_1149,N_9884,N_9959);
and UO_1150 (O_1150,N_9964,N_9954);
and UO_1151 (O_1151,N_9948,N_9925);
nand UO_1152 (O_1152,N_9957,N_9909);
nand UO_1153 (O_1153,N_9894,N_9979);
nor UO_1154 (O_1154,N_9893,N_9933);
nor UO_1155 (O_1155,N_9924,N_9837);
nand UO_1156 (O_1156,N_9850,N_9860);
nand UO_1157 (O_1157,N_9989,N_9911);
or UO_1158 (O_1158,N_9803,N_9857);
and UO_1159 (O_1159,N_9928,N_9965);
or UO_1160 (O_1160,N_9997,N_9811);
nor UO_1161 (O_1161,N_9912,N_9889);
nand UO_1162 (O_1162,N_9852,N_9871);
nor UO_1163 (O_1163,N_9830,N_9939);
nor UO_1164 (O_1164,N_9808,N_9973);
nor UO_1165 (O_1165,N_9868,N_9963);
nor UO_1166 (O_1166,N_9818,N_9988);
and UO_1167 (O_1167,N_9886,N_9845);
and UO_1168 (O_1168,N_9965,N_9858);
and UO_1169 (O_1169,N_9853,N_9928);
or UO_1170 (O_1170,N_9866,N_9995);
or UO_1171 (O_1171,N_9992,N_9810);
xnor UO_1172 (O_1172,N_9886,N_9891);
or UO_1173 (O_1173,N_9885,N_9816);
or UO_1174 (O_1174,N_9968,N_9972);
nor UO_1175 (O_1175,N_9875,N_9954);
nor UO_1176 (O_1176,N_9949,N_9809);
and UO_1177 (O_1177,N_9833,N_9928);
xnor UO_1178 (O_1178,N_9943,N_9956);
nor UO_1179 (O_1179,N_9919,N_9867);
and UO_1180 (O_1180,N_9862,N_9839);
nor UO_1181 (O_1181,N_9853,N_9939);
or UO_1182 (O_1182,N_9922,N_9863);
nor UO_1183 (O_1183,N_9817,N_9981);
and UO_1184 (O_1184,N_9945,N_9950);
and UO_1185 (O_1185,N_9912,N_9910);
nand UO_1186 (O_1186,N_9915,N_9894);
nand UO_1187 (O_1187,N_9983,N_9800);
xor UO_1188 (O_1188,N_9850,N_9984);
and UO_1189 (O_1189,N_9897,N_9887);
or UO_1190 (O_1190,N_9874,N_9870);
and UO_1191 (O_1191,N_9842,N_9995);
nor UO_1192 (O_1192,N_9970,N_9817);
and UO_1193 (O_1193,N_9927,N_9866);
or UO_1194 (O_1194,N_9945,N_9841);
xor UO_1195 (O_1195,N_9881,N_9850);
and UO_1196 (O_1196,N_9889,N_9830);
or UO_1197 (O_1197,N_9916,N_9840);
nand UO_1198 (O_1198,N_9885,N_9957);
or UO_1199 (O_1199,N_9920,N_9904);
nand UO_1200 (O_1200,N_9847,N_9981);
nand UO_1201 (O_1201,N_9901,N_9887);
nor UO_1202 (O_1202,N_9931,N_9902);
or UO_1203 (O_1203,N_9852,N_9811);
and UO_1204 (O_1204,N_9921,N_9937);
and UO_1205 (O_1205,N_9816,N_9898);
and UO_1206 (O_1206,N_9902,N_9851);
nor UO_1207 (O_1207,N_9845,N_9851);
or UO_1208 (O_1208,N_9969,N_9985);
nand UO_1209 (O_1209,N_9889,N_9811);
and UO_1210 (O_1210,N_9824,N_9888);
or UO_1211 (O_1211,N_9907,N_9925);
xnor UO_1212 (O_1212,N_9926,N_9838);
or UO_1213 (O_1213,N_9832,N_9977);
nor UO_1214 (O_1214,N_9872,N_9827);
or UO_1215 (O_1215,N_9970,N_9840);
nor UO_1216 (O_1216,N_9822,N_9932);
nand UO_1217 (O_1217,N_9963,N_9945);
and UO_1218 (O_1218,N_9904,N_9840);
xor UO_1219 (O_1219,N_9814,N_9953);
or UO_1220 (O_1220,N_9874,N_9856);
nand UO_1221 (O_1221,N_9988,N_9803);
nor UO_1222 (O_1222,N_9889,N_9986);
and UO_1223 (O_1223,N_9823,N_9814);
nor UO_1224 (O_1224,N_9831,N_9980);
nand UO_1225 (O_1225,N_9958,N_9924);
nor UO_1226 (O_1226,N_9843,N_9939);
nor UO_1227 (O_1227,N_9805,N_9888);
nand UO_1228 (O_1228,N_9853,N_9972);
nor UO_1229 (O_1229,N_9981,N_9842);
nand UO_1230 (O_1230,N_9958,N_9827);
and UO_1231 (O_1231,N_9918,N_9968);
or UO_1232 (O_1232,N_9827,N_9862);
nand UO_1233 (O_1233,N_9812,N_9823);
and UO_1234 (O_1234,N_9904,N_9817);
nand UO_1235 (O_1235,N_9854,N_9873);
nand UO_1236 (O_1236,N_9958,N_9965);
or UO_1237 (O_1237,N_9873,N_9866);
nor UO_1238 (O_1238,N_9934,N_9940);
nor UO_1239 (O_1239,N_9938,N_9879);
or UO_1240 (O_1240,N_9928,N_9892);
and UO_1241 (O_1241,N_9905,N_9811);
and UO_1242 (O_1242,N_9816,N_9934);
nand UO_1243 (O_1243,N_9867,N_9845);
nand UO_1244 (O_1244,N_9840,N_9899);
nand UO_1245 (O_1245,N_9925,N_9822);
or UO_1246 (O_1246,N_9890,N_9943);
nand UO_1247 (O_1247,N_9805,N_9908);
or UO_1248 (O_1248,N_9946,N_9869);
or UO_1249 (O_1249,N_9905,N_9861);
nand UO_1250 (O_1250,N_9948,N_9923);
and UO_1251 (O_1251,N_9898,N_9838);
and UO_1252 (O_1252,N_9944,N_9850);
and UO_1253 (O_1253,N_9854,N_9865);
nor UO_1254 (O_1254,N_9819,N_9919);
nor UO_1255 (O_1255,N_9867,N_9991);
or UO_1256 (O_1256,N_9919,N_9889);
nor UO_1257 (O_1257,N_9936,N_9870);
nor UO_1258 (O_1258,N_9819,N_9855);
nand UO_1259 (O_1259,N_9805,N_9916);
or UO_1260 (O_1260,N_9964,N_9874);
or UO_1261 (O_1261,N_9804,N_9980);
nand UO_1262 (O_1262,N_9906,N_9940);
xnor UO_1263 (O_1263,N_9882,N_9870);
xor UO_1264 (O_1264,N_9848,N_9869);
nor UO_1265 (O_1265,N_9882,N_9851);
or UO_1266 (O_1266,N_9856,N_9843);
or UO_1267 (O_1267,N_9914,N_9806);
or UO_1268 (O_1268,N_9923,N_9886);
nor UO_1269 (O_1269,N_9949,N_9960);
nor UO_1270 (O_1270,N_9904,N_9806);
nor UO_1271 (O_1271,N_9986,N_9813);
nor UO_1272 (O_1272,N_9913,N_9903);
nor UO_1273 (O_1273,N_9976,N_9999);
and UO_1274 (O_1274,N_9989,N_9800);
nand UO_1275 (O_1275,N_9845,N_9902);
and UO_1276 (O_1276,N_9978,N_9966);
nand UO_1277 (O_1277,N_9897,N_9911);
nand UO_1278 (O_1278,N_9958,N_9867);
xnor UO_1279 (O_1279,N_9803,N_9887);
and UO_1280 (O_1280,N_9991,N_9997);
nand UO_1281 (O_1281,N_9892,N_9816);
and UO_1282 (O_1282,N_9944,N_9965);
and UO_1283 (O_1283,N_9851,N_9811);
and UO_1284 (O_1284,N_9914,N_9969);
or UO_1285 (O_1285,N_9836,N_9905);
nor UO_1286 (O_1286,N_9904,N_9864);
and UO_1287 (O_1287,N_9814,N_9810);
or UO_1288 (O_1288,N_9860,N_9895);
or UO_1289 (O_1289,N_9902,N_9981);
or UO_1290 (O_1290,N_9951,N_9887);
nor UO_1291 (O_1291,N_9858,N_9930);
and UO_1292 (O_1292,N_9977,N_9897);
nor UO_1293 (O_1293,N_9949,N_9864);
and UO_1294 (O_1294,N_9858,N_9846);
and UO_1295 (O_1295,N_9837,N_9904);
nor UO_1296 (O_1296,N_9888,N_9905);
xnor UO_1297 (O_1297,N_9974,N_9899);
and UO_1298 (O_1298,N_9946,N_9850);
or UO_1299 (O_1299,N_9987,N_9962);
or UO_1300 (O_1300,N_9974,N_9881);
nor UO_1301 (O_1301,N_9864,N_9884);
nor UO_1302 (O_1302,N_9836,N_9860);
and UO_1303 (O_1303,N_9978,N_9836);
and UO_1304 (O_1304,N_9867,N_9834);
nand UO_1305 (O_1305,N_9855,N_9901);
or UO_1306 (O_1306,N_9887,N_9964);
nor UO_1307 (O_1307,N_9985,N_9904);
nand UO_1308 (O_1308,N_9910,N_9828);
nand UO_1309 (O_1309,N_9918,N_9978);
and UO_1310 (O_1310,N_9840,N_9972);
or UO_1311 (O_1311,N_9839,N_9843);
and UO_1312 (O_1312,N_9917,N_9968);
nand UO_1313 (O_1313,N_9925,N_9916);
and UO_1314 (O_1314,N_9839,N_9939);
and UO_1315 (O_1315,N_9889,N_9869);
or UO_1316 (O_1316,N_9881,N_9937);
nand UO_1317 (O_1317,N_9888,N_9841);
nor UO_1318 (O_1318,N_9822,N_9888);
nand UO_1319 (O_1319,N_9804,N_9954);
nor UO_1320 (O_1320,N_9801,N_9860);
nor UO_1321 (O_1321,N_9869,N_9913);
and UO_1322 (O_1322,N_9803,N_9982);
or UO_1323 (O_1323,N_9869,N_9910);
or UO_1324 (O_1324,N_9925,N_9843);
nor UO_1325 (O_1325,N_9890,N_9804);
xor UO_1326 (O_1326,N_9836,N_9957);
or UO_1327 (O_1327,N_9948,N_9911);
and UO_1328 (O_1328,N_9971,N_9865);
nand UO_1329 (O_1329,N_9991,N_9985);
or UO_1330 (O_1330,N_9862,N_9966);
and UO_1331 (O_1331,N_9920,N_9940);
nor UO_1332 (O_1332,N_9830,N_9984);
xnor UO_1333 (O_1333,N_9857,N_9904);
nand UO_1334 (O_1334,N_9987,N_9833);
nand UO_1335 (O_1335,N_9811,N_9981);
nand UO_1336 (O_1336,N_9932,N_9885);
and UO_1337 (O_1337,N_9898,N_9814);
and UO_1338 (O_1338,N_9892,N_9909);
or UO_1339 (O_1339,N_9882,N_9809);
nand UO_1340 (O_1340,N_9950,N_9958);
or UO_1341 (O_1341,N_9881,N_9852);
and UO_1342 (O_1342,N_9823,N_9848);
nor UO_1343 (O_1343,N_9990,N_9880);
or UO_1344 (O_1344,N_9978,N_9911);
or UO_1345 (O_1345,N_9959,N_9831);
nand UO_1346 (O_1346,N_9807,N_9894);
nand UO_1347 (O_1347,N_9906,N_9987);
nor UO_1348 (O_1348,N_9865,N_9838);
nand UO_1349 (O_1349,N_9896,N_9866);
or UO_1350 (O_1350,N_9958,N_9971);
nand UO_1351 (O_1351,N_9844,N_9879);
nand UO_1352 (O_1352,N_9987,N_9951);
nand UO_1353 (O_1353,N_9973,N_9849);
xor UO_1354 (O_1354,N_9965,N_9946);
nand UO_1355 (O_1355,N_9871,N_9980);
and UO_1356 (O_1356,N_9996,N_9925);
and UO_1357 (O_1357,N_9928,N_9956);
nand UO_1358 (O_1358,N_9950,N_9988);
and UO_1359 (O_1359,N_9954,N_9987);
nor UO_1360 (O_1360,N_9975,N_9843);
or UO_1361 (O_1361,N_9891,N_9861);
or UO_1362 (O_1362,N_9999,N_9898);
or UO_1363 (O_1363,N_9999,N_9848);
xor UO_1364 (O_1364,N_9933,N_9943);
nand UO_1365 (O_1365,N_9997,N_9823);
and UO_1366 (O_1366,N_9878,N_9913);
and UO_1367 (O_1367,N_9914,N_9802);
and UO_1368 (O_1368,N_9880,N_9839);
or UO_1369 (O_1369,N_9958,N_9911);
or UO_1370 (O_1370,N_9928,N_9969);
nor UO_1371 (O_1371,N_9979,N_9930);
and UO_1372 (O_1372,N_9882,N_9899);
and UO_1373 (O_1373,N_9955,N_9935);
or UO_1374 (O_1374,N_9930,N_9961);
nand UO_1375 (O_1375,N_9829,N_9979);
and UO_1376 (O_1376,N_9956,N_9968);
nand UO_1377 (O_1377,N_9806,N_9877);
nor UO_1378 (O_1378,N_9924,N_9915);
nand UO_1379 (O_1379,N_9820,N_9926);
nor UO_1380 (O_1380,N_9896,N_9903);
or UO_1381 (O_1381,N_9899,N_9936);
or UO_1382 (O_1382,N_9930,N_9805);
nand UO_1383 (O_1383,N_9966,N_9808);
or UO_1384 (O_1384,N_9804,N_9974);
and UO_1385 (O_1385,N_9906,N_9825);
nand UO_1386 (O_1386,N_9902,N_9891);
nor UO_1387 (O_1387,N_9935,N_9848);
or UO_1388 (O_1388,N_9950,N_9897);
and UO_1389 (O_1389,N_9808,N_9922);
or UO_1390 (O_1390,N_9952,N_9907);
and UO_1391 (O_1391,N_9813,N_9824);
and UO_1392 (O_1392,N_9864,N_9800);
nor UO_1393 (O_1393,N_9880,N_9804);
nor UO_1394 (O_1394,N_9994,N_9917);
nand UO_1395 (O_1395,N_9822,N_9920);
nand UO_1396 (O_1396,N_9911,N_9967);
and UO_1397 (O_1397,N_9891,N_9881);
nand UO_1398 (O_1398,N_9831,N_9851);
nand UO_1399 (O_1399,N_9927,N_9945);
nor UO_1400 (O_1400,N_9856,N_9810);
nand UO_1401 (O_1401,N_9963,N_9977);
and UO_1402 (O_1402,N_9935,N_9892);
nand UO_1403 (O_1403,N_9818,N_9940);
nand UO_1404 (O_1404,N_9961,N_9911);
and UO_1405 (O_1405,N_9943,N_9882);
and UO_1406 (O_1406,N_9997,N_9809);
nor UO_1407 (O_1407,N_9839,N_9981);
or UO_1408 (O_1408,N_9910,N_9874);
or UO_1409 (O_1409,N_9817,N_9950);
or UO_1410 (O_1410,N_9892,N_9967);
nand UO_1411 (O_1411,N_9831,N_9832);
or UO_1412 (O_1412,N_9824,N_9884);
nand UO_1413 (O_1413,N_9931,N_9930);
nand UO_1414 (O_1414,N_9961,N_9931);
nor UO_1415 (O_1415,N_9939,N_9881);
or UO_1416 (O_1416,N_9879,N_9819);
nand UO_1417 (O_1417,N_9818,N_9989);
nor UO_1418 (O_1418,N_9945,N_9926);
nor UO_1419 (O_1419,N_9872,N_9840);
or UO_1420 (O_1420,N_9818,N_9892);
nand UO_1421 (O_1421,N_9898,N_9841);
nand UO_1422 (O_1422,N_9955,N_9839);
nor UO_1423 (O_1423,N_9819,N_9870);
nor UO_1424 (O_1424,N_9876,N_9854);
nand UO_1425 (O_1425,N_9986,N_9893);
nand UO_1426 (O_1426,N_9844,N_9985);
or UO_1427 (O_1427,N_9976,N_9834);
nor UO_1428 (O_1428,N_9913,N_9926);
nand UO_1429 (O_1429,N_9837,N_9892);
or UO_1430 (O_1430,N_9964,N_9978);
and UO_1431 (O_1431,N_9833,N_9896);
and UO_1432 (O_1432,N_9978,N_9938);
and UO_1433 (O_1433,N_9899,N_9826);
or UO_1434 (O_1434,N_9929,N_9921);
xor UO_1435 (O_1435,N_9811,N_9900);
and UO_1436 (O_1436,N_9891,N_9896);
nand UO_1437 (O_1437,N_9885,N_9831);
or UO_1438 (O_1438,N_9876,N_9936);
nand UO_1439 (O_1439,N_9970,N_9989);
nand UO_1440 (O_1440,N_9878,N_9997);
nand UO_1441 (O_1441,N_9985,N_9874);
or UO_1442 (O_1442,N_9810,N_9800);
or UO_1443 (O_1443,N_9933,N_9982);
and UO_1444 (O_1444,N_9803,N_9983);
nand UO_1445 (O_1445,N_9867,N_9812);
or UO_1446 (O_1446,N_9870,N_9899);
or UO_1447 (O_1447,N_9872,N_9932);
nor UO_1448 (O_1448,N_9964,N_9859);
and UO_1449 (O_1449,N_9987,N_9976);
and UO_1450 (O_1450,N_9932,N_9935);
nor UO_1451 (O_1451,N_9881,N_9909);
and UO_1452 (O_1452,N_9967,N_9857);
and UO_1453 (O_1453,N_9967,N_9996);
and UO_1454 (O_1454,N_9949,N_9902);
nand UO_1455 (O_1455,N_9915,N_9845);
nor UO_1456 (O_1456,N_9860,N_9954);
xnor UO_1457 (O_1457,N_9936,N_9846);
and UO_1458 (O_1458,N_9929,N_9841);
and UO_1459 (O_1459,N_9891,N_9880);
or UO_1460 (O_1460,N_9913,N_9938);
or UO_1461 (O_1461,N_9803,N_9808);
xor UO_1462 (O_1462,N_9877,N_9962);
nor UO_1463 (O_1463,N_9809,N_9836);
nand UO_1464 (O_1464,N_9804,N_9914);
xnor UO_1465 (O_1465,N_9836,N_9816);
or UO_1466 (O_1466,N_9858,N_9867);
or UO_1467 (O_1467,N_9921,N_9862);
nand UO_1468 (O_1468,N_9980,N_9966);
or UO_1469 (O_1469,N_9878,N_9808);
nor UO_1470 (O_1470,N_9857,N_9913);
and UO_1471 (O_1471,N_9806,N_9935);
nand UO_1472 (O_1472,N_9939,N_9910);
nand UO_1473 (O_1473,N_9926,N_9804);
nand UO_1474 (O_1474,N_9826,N_9894);
nor UO_1475 (O_1475,N_9906,N_9881);
nor UO_1476 (O_1476,N_9916,N_9961);
nor UO_1477 (O_1477,N_9966,N_9821);
nor UO_1478 (O_1478,N_9876,N_9950);
or UO_1479 (O_1479,N_9849,N_9970);
xor UO_1480 (O_1480,N_9927,N_9987);
and UO_1481 (O_1481,N_9868,N_9950);
or UO_1482 (O_1482,N_9864,N_9897);
and UO_1483 (O_1483,N_9957,N_9852);
or UO_1484 (O_1484,N_9857,N_9809);
nor UO_1485 (O_1485,N_9896,N_9850);
nor UO_1486 (O_1486,N_9816,N_9814);
and UO_1487 (O_1487,N_9896,N_9995);
nand UO_1488 (O_1488,N_9869,N_9804);
nand UO_1489 (O_1489,N_9947,N_9909);
and UO_1490 (O_1490,N_9838,N_9810);
or UO_1491 (O_1491,N_9880,N_9973);
or UO_1492 (O_1492,N_9984,N_9863);
nor UO_1493 (O_1493,N_9821,N_9979);
nor UO_1494 (O_1494,N_9907,N_9961);
or UO_1495 (O_1495,N_9987,N_9907);
nand UO_1496 (O_1496,N_9826,N_9817);
or UO_1497 (O_1497,N_9850,N_9955);
nor UO_1498 (O_1498,N_9859,N_9821);
or UO_1499 (O_1499,N_9867,N_9853);
endmodule