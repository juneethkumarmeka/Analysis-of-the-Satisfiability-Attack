module basic_500_3000_500_30_levels_2xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_365,In_157);
and U1 (N_1,In_297,In_282);
and U2 (N_2,In_433,In_107);
nand U3 (N_3,In_411,In_179);
nor U4 (N_4,In_221,In_419);
nor U5 (N_5,In_210,In_177);
and U6 (N_6,In_215,In_286);
and U7 (N_7,In_133,In_130);
and U8 (N_8,In_61,In_67);
nor U9 (N_9,In_431,In_92);
and U10 (N_10,In_327,In_322);
or U11 (N_11,In_277,In_229);
and U12 (N_12,In_190,In_479);
or U13 (N_13,In_474,In_470);
and U14 (N_14,In_156,In_112);
or U15 (N_15,In_460,In_63);
or U16 (N_16,In_427,In_87);
or U17 (N_17,In_298,In_422);
nor U18 (N_18,In_99,In_90);
nor U19 (N_19,In_234,In_262);
and U20 (N_20,In_96,In_165);
nor U21 (N_21,In_18,In_22);
or U22 (N_22,In_467,In_402);
nand U23 (N_23,In_345,In_310);
nor U24 (N_24,In_155,In_247);
nor U25 (N_25,In_239,In_26);
nand U26 (N_26,In_136,In_129);
or U27 (N_27,In_464,In_14);
nor U28 (N_28,In_104,In_97);
nor U29 (N_29,In_28,In_123);
or U30 (N_30,In_366,In_252);
nor U31 (N_31,In_226,In_225);
nor U32 (N_32,In_486,In_321);
or U33 (N_33,In_75,In_421);
or U34 (N_34,In_280,In_455);
and U35 (N_35,In_95,In_152);
and U36 (N_36,In_200,In_43);
nand U37 (N_37,In_176,In_432);
or U38 (N_38,In_42,In_77);
and U39 (N_39,In_415,In_16);
xor U40 (N_40,In_472,In_466);
and U41 (N_41,In_450,In_407);
or U42 (N_42,In_162,In_287);
nand U43 (N_43,In_265,In_72);
nand U44 (N_44,In_238,In_307);
and U45 (N_45,In_167,In_308);
and U46 (N_46,In_144,In_41);
or U47 (N_47,In_424,In_279);
and U48 (N_48,In_168,In_369);
nor U49 (N_49,In_246,In_304);
nor U50 (N_50,In_7,In_219);
or U51 (N_51,In_64,In_438);
and U52 (N_52,In_484,In_452);
nor U53 (N_53,In_164,In_45);
nor U54 (N_54,In_120,In_326);
nor U55 (N_55,In_70,In_59);
nor U56 (N_56,In_413,In_55);
or U57 (N_57,In_426,In_334);
xnor U58 (N_58,In_150,In_111);
nor U59 (N_59,In_311,In_122);
and U60 (N_60,In_254,In_249);
xor U61 (N_61,In_335,In_357);
nor U62 (N_62,In_390,In_121);
nand U63 (N_63,In_51,In_347);
nor U64 (N_64,In_272,In_53);
or U65 (N_65,In_232,In_209);
or U66 (N_66,In_73,In_355);
nor U67 (N_67,In_275,In_456);
nand U68 (N_68,In_493,In_263);
and U69 (N_69,In_278,In_217);
nand U70 (N_70,In_463,In_399);
and U71 (N_71,In_199,In_159);
or U72 (N_72,In_137,In_291);
or U73 (N_73,In_416,In_346);
or U74 (N_74,In_370,In_425);
nor U75 (N_75,In_480,In_344);
xor U76 (N_76,In_141,In_441);
or U77 (N_77,In_256,In_13);
and U78 (N_78,In_206,In_68);
nand U79 (N_79,In_227,In_294);
or U80 (N_80,In_5,In_231);
or U81 (N_81,In_188,In_32);
nand U82 (N_82,In_267,In_330);
nor U83 (N_83,In_158,In_193);
and U84 (N_84,In_273,In_264);
nand U85 (N_85,In_350,In_66);
nand U86 (N_86,In_269,In_353);
and U87 (N_87,In_482,In_380);
nand U88 (N_88,In_12,In_409);
and U89 (N_89,In_69,In_180);
nor U90 (N_90,In_125,In_172);
nand U91 (N_91,In_250,In_197);
and U92 (N_92,In_235,In_203);
nor U93 (N_93,In_471,In_317);
nor U94 (N_94,In_338,In_309);
or U95 (N_95,In_389,In_285);
xnor U96 (N_96,In_6,In_196);
nor U97 (N_97,In_11,In_363);
nand U98 (N_98,In_377,In_174);
or U99 (N_99,In_305,In_316);
xor U100 (N_100,In_497,In_270);
nand U101 (N_101,N_54,In_436);
nor U102 (N_102,N_46,N_9);
and U103 (N_103,In_27,N_65);
and U104 (N_104,N_25,In_336);
and U105 (N_105,In_34,In_251);
or U106 (N_106,In_313,N_21);
nor U107 (N_107,In_443,In_85);
nor U108 (N_108,N_24,In_284);
and U109 (N_109,N_6,N_97);
nand U110 (N_110,In_56,N_29);
nand U111 (N_111,In_373,In_154);
or U112 (N_112,In_105,N_58);
nor U113 (N_113,N_2,In_82);
or U114 (N_114,In_428,N_93);
and U115 (N_115,N_37,In_364);
and U116 (N_116,In_83,In_406);
and U117 (N_117,In_352,In_478);
nor U118 (N_118,In_183,In_116);
nand U119 (N_119,N_57,In_359);
or U120 (N_120,N_32,In_462);
nand U121 (N_121,In_400,In_376);
or U122 (N_122,In_106,In_417);
and U123 (N_123,In_477,In_114);
or U124 (N_124,In_451,In_283);
nor U125 (N_125,In_496,N_27);
or U126 (N_126,N_16,In_429);
and U127 (N_127,In_381,In_31);
nor U128 (N_128,In_76,In_185);
nor U129 (N_129,In_405,In_367);
nor U130 (N_130,N_60,In_461);
nor U131 (N_131,In_362,In_86);
nor U132 (N_132,N_22,In_198);
nor U133 (N_133,N_80,In_19);
or U134 (N_134,In_457,In_333);
nand U135 (N_135,N_91,In_81);
and U136 (N_136,In_170,In_361);
and U137 (N_137,N_59,In_356);
or U138 (N_138,In_1,In_341);
and U139 (N_139,In_138,N_1);
and U140 (N_140,In_93,In_224);
nor U141 (N_141,In_54,In_212);
nand U142 (N_142,In_292,In_3);
and U143 (N_143,In_50,N_67);
or U144 (N_144,In_384,N_64);
or U145 (N_145,In_147,In_368);
and U146 (N_146,In_74,In_483);
or U147 (N_147,N_85,In_192);
and U148 (N_148,In_499,In_204);
nand U149 (N_149,N_39,In_293);
or U150 (N_150,In_266,In_258);
nor U151 (N_151,In_145,N_53);
or U152 (N_152,In_329,In_8);
nor U153 (N_153,In_323,In_160);
and U154 (N_154,In_488,In_469);
nor U155 (N_155,In_211,N_13);
nand U156 (N_156,In_371,In_20);
nor U157 (N_157,In_260,In_140);
and U158 (N_158,N_95,N_87);
or U159 (N_159,N_56,In_49);
nand U160 (N_160,In_171,In_0);
or U161 (N_161,In_281,In_442);
nand U162 (N_162,In_358,In_349);
or U163 (N_163,In_60,N_88);
nand U164 (N_164,In_240,In_79);
or U165 (N_165,N_12,In_98);
or U166 (N_166,In_414,In_91);
nor U167 (N_167,In_388,In_117);
nand U168 (N_168,In_102,In_430);
nand U169 (N_169,In_223,In_103);
nand U170 (N_170,In_386,In_408);
nand U171 (N_171,In_119,In_303);
or U172 (N_172,In_444,In_131);
or U173 (N_173,In_135,In_395);
and U174 (N_174,In_412,In_184);
or U175 (N_175,In_374,In_447);
and U176 (N_176,In_261,In_134);
or U177 (N_177,In_44,In_300);
or U178 (N_178,N_61,In_448);
nor U179 (N_179,In_65,In_236);
and U180 (N_180,In_276,In_40);
nand U181 (N_181,In_161,In_47);
nor U182 (N_182,In_126,In_392);
or U183 (N_183,In_299,N_99);
or U184 (N_184,In_393,In_437);
nand U185 (N_185,In_30,N_82);
nand U186 (N_186,N_49,In_271);
or U187 (N_187,In_481,In_268);
nand U188 (N_188,In_473,In_84);
nor U189 (N_189,N_47,In_385);
or U190 (N_190,In_195,In_494);
and U191 (N_191,In_397,In_314);
and U192 (N_192,In_255,In_398);
and U193 (N_193,In_301,N_41);
nand U194 (N_194,In_110,In_453);
and U195 (N_195,In_495,In_324);
and U196 (N_196,N_90,In_78);
and U197 (N_197,In_319,N_31);
nand U198 (N_198,In_108,N_69);
nor U199 (N_199,In_80,N_98);
and U200 (N_200,N_113,N_159);
nor U201 (N_201,In_245,In_387);
nand U202 (N_202,N_23,In_4);
nor U203 (N_203,In_342,N_40);
xnor U204 (N_204,N_156,In_169);
nand U205 (N_205,In_476,In_289);
nor U206 (N_206,N_5,N_134);
or U207 (N_207,In_194,In_205);
nand U208 (N_208,N_4,In_446);
or U209 (N_209,N_194,N_78);
nand U210 (N_210,In_343,N_100);
and U211 (N_211,In_24,N_74);
nand U212 (N_212,N_119,In_382);
or U213 (N_213,In_38,N_62);
and U214 (N_214,In_331,N_193);
and U215 (N_215,N_50,N_136);
or U216 (N_216,N_186,N_187);
xnor U217 (N_217,In_290,N_20);
nand U218 (N_218,N_188,N_36);
and U219 (N_219,N_73,In_318);
xnor U220 (N_220,N_123,N_181);
nor U221 (N_221,N_28,N_109);
nand U222 (N_222,N_7,In_378);
and U223 (N_223,In_202,In_62);
and U224 (N_224,N_125,In_306);
nor U225 (N_225,N_140,N_26);
or U226 (N_226,In_148,In_52);
nor U227 (N_227,N_104,N_155);
and U228 (N_228,In_36,N_81);
or U229 (N_229,In_458,N_35);
or U230 (N_230,N_169,In_187);
nand U231 (N_231,In_492,N_124);
or U232 (N_232,N_160,N_105);
nor U233 (N_233,N_101,N_161);
or U234 (N_234,N_14,In_244);
nor U235 (N_235,In_325,N_177);
and U236 (N_236,In_153,In_296);
and U237 (N_237,N_146,N_55);
nor U238 (N_238,In_25,In_89);
or U239 (N_239,In_23,N_107);
nor U240 (N_240,In_348,N_185);
nand U241 (N_241,In_253,In_113);
or U242 (N_242,In_401,N_128);
nor U243 (N_243,In_259,N_66);
nor U244 (N_244,N_8,N_17);
nand U245 (N_245,In_201,In_394);
nor U246 (N_246,In_332,In_178);
or U247 (N_247,N_96,In_465);
or U248 (N_248,In_146,N_71);
and U249 (N_249,N_130,In_71);
or U250 (N_250,N_77,In_186);
or U251 (N_251,In_491,In_487);
and U252 (N_252,In_320,N_48);
nor U253 (N_253,N_148,In_128);
nand U254 (N_254,N_189,In_37);
and U255 (N_255,N_166,N_103);
xnor U256 (N_256,In_57,In_21);
nor U257 (N_257,In_340,N_131);
nand U258 (N_258,N_84,In_100);
nand U259 (N_259,In_191,N_122);
and U260 (N_260,In_94,In_449);
nand U261 (N_261,N_30,In_439);
nor U262 (N_262,N_102,N_115);
nor U263 (N_263,In_454,N_197);
or U264 (N_264,In_208,In_295);
and U265 (N_265,N_150,N_11);
nand U266 (N_266,In_46,N_68);
nor U267 (N_267,In_132,N_129);
and U268 (N_268,N_138,In_109);
nor U269 (N_269,In_88,In_2);
or U270 (N_270,In_173,N_142);
nor U271 (N_271,In_127,In_337);
and U272 (N_272,N_10,N_72);
nand U273 (N_273,In_29,N_149);
and U274 (N_274,N_157,N_89);
nand U275 (N_275,N_120,In_383);
nand U276 (N_276,N_170,N_154);
xnor U277 (N_277,N_164,N_162);
and U278 (N_278,In_207,In_149);
xnor U279 (N_279,In_118,In_339);
or U280 (N_280,N_151,N_174);
and U281 (N_281,In_391,N_141);
nand U282 (N_282,N_165,In_403);
or U283 (N_283,N_94,N_179);
nor U284 (N_284,In_248,In_175);
nor U285 (N_285,In_9,N_118);
and U286 (N_286,N_171,N_191);
nor U287 (N_287,N_175,In_15);
or U288 (N_288,N_38,In_166);
xnor U289 (N_289,N_127,In_48);
nand U290 (N_290,In_485,In_163);
and U291 (N_291,N_135,N_192);
nand U292 (N_292,In_139,N_83);
or U293 (N_293,N_19,In_151);
and U294 (N_294,In_257,In_423);
nor U295 (N_295,In_233,In_230);
nor U296 (N_296,In_17,N_108);
and U297 (N_297,In_475,N_183);
or U298 (N_298,In_143,N_112);
or U299 (N_299,In_490,N_117);
or U300 (N_300,N_152,N_266);
and U301 (N_301,N_255,N_292);
nand U302 (N_302,N_121,N_208);
nor U303 (N_303,N_147,N_239);
nor U304 (N_304,In_396,In_182);
xnor U305 (N_305,N_264,N_280);
and U306 (N_306,N_110,N_220);
nand U307 (N_307,N_45,In_375);
or U308 (N_308,N_290,N_275);
nor U309 (N_309,N_281,N_213);
nor U310 (N_310,N_285,N_202);
nor U311 (N_311,N_261,In_115);
nor U312 (N_312,N_215,N_258);
nor U313 (N_313,N_182,N_145);
nand U314 (N_314,In_35,N_274);
or U315 (N_315,N_268,N_296);
nor U316 (N_316,In_241,In_288);
xor U317 (N_317,N_229,In_214);
or U318 (N_318,N_240,In_468);
or U319 (N_319,N_252,In_379);
or U320 (N_320,N_263,N_70);
or U321 (N_321,N_201,In_498);
and U322 (N_322,N_206,In_243);
and U323 (N_323,N_250,N_75);
and U324 (N_324,In_237,N_257);
and U325 (N_325,N_176,In_302);
nand U326 (N_326,N_277,In_440);
nor U327 (N_327,N_288,N_256);
xor U328 (N_328,N_86,N_294);
or U329 (N_329,In_181,N_111);
nand U330 (N_330,N_249,N_163);
and U331 (N_331,N_34,N_198);
and U332 (N_332,N_224,In_372);
or U333 (N_333,N_259,In_459);
nand U334 (N_334,N_52,N_242);
nor U335 (N_335,N_247,N_298);
or U336 (N_336,N_295,In_39);
nor U337 (N_337,In_328,In_434);
or U338 (N_338,N_293,N_238);
nor U339 (N_339,N_279,In_312);
nand U340 (N_340,N_204,N_219);
or U341 (N_341,N_212,In_274);
and U342 (N_342,N_214,N_217);
nor U343 (N_343,N_271,In_220);
nand U344 (N_344,N_172,In_445);
nand U345 (N_345,In_420,N_272);
nor U346 (N_346,N_203,N_3);
and U347 (N_347,N_235,In_58);
and U348 (N_348,N_251,N_63);
nand U349 (N_349,N_0,N_18);
nor U350 (N_350,N_195,N_253);
nand U351 (N_351,In_216,N_196);
nor U352 (N_352,N_178,N_269);
or U353 (N_353,N_237,In_489);
nor U354 (N_354,N_278,N_221);
and U355 (N_355,N_289,N_116);
nand U356 (N_356,N_43,N_51);
or U357 (N_357,In_228,N_218);
nor U358 (N_358,N_207,In_242);
nand U359 (N_359,N_106,N_245);
nand U360 (N_360,In_218,N_225);
nand U361 (N_361,N_243,N_33);
or U362 (N_362,N_291,In_418);
nand U363 (N_363,N_92,N_228);
or U364 (N_364,N_132,N_137);
or U365 (N_365,N_114,N_234);
and U366 (N_366,In_213,In_410);
nand U367 (N_367,N_158,N_227);
or U368 (N_368,N_230,In_10);
nor U369 (N_369,N_233,In_360);
or U370 (N_370,In_404,N_254);
nor U371 (N_371,In_315,In_101);
nor U372 (N_372,N_173,In_33);
and U373 (N_373,N_297,N_284);
nand U374 (N_374,N_262,N_283);
or U375 (N_375,N_209,N_270);
and U376 (N_376,N_236,N_210);
or U377 (N_377,N_15,N_246);
nor U378 (N_378,N_126,N_222);
nand U379 (N_379,N_241,N_190);
xor U380 (N_380,N_44,N_139);
and U381 (N_381,In_189,N_180);
nand U382 (N_382,In_142,N_287);
nor U383 (N_383,N_205,N_232);
and U384 (N_384,In_354,N_276);
nand U385 (N_385,N_133,N_79);
nor U386 (N_386,N_244,N_144);
nor U387 (N_387,N_231,N_168);
nor U388 (N_388,N_184,N_267);
and U389 (N_389,N_282,In_222);
or U390 (N_390,N_299,N_42);
nor U391 (N_391,N_211,N_286);
and U392 (N_392,N_248,N_199);
and U393 (N_393,In_435,N_273);
xnor U394 (N_394,In_351,N_260);
nor U395 (N_395,In_124,N_216);
nand U396 (N_396,N_153,N_143);
and U397 (N_397,N_226,N_167);
or U398 (N_398,N_223,N_76);
and U399 (N_399,N_200,N_265);
nor U400 (N_400,N_395,N_306);
nor U401 (N_401,N_366,N_307);
nand U402 (N_402,N_360,N_375);
nand U403 (N_403,N_354,N_319);
nor U404 (N_404,N_342,N_330);
xor U405 (N_405,N_368,N_304);
nand U406 (N_406,N_383,N_387);
and U407 (N_407,N_370,N_337);
nand U408 (N_408,N_334,N_318);
nand U409 (N_409,N_321,N_324);
or U410 (N_410,N_372,N_333);
and U411 (N_411,N_388,N_393);
nor U412 (N_412,N_301,N_351);
or U413 (N_413,N_399,N_384);
xnor U414 (N_414,N_377,N_317);
nor U415 (N_415,N_339,N_356);
or U416 (N_416,N_331,N_320);
nand U417 (N_417,N_350,N_359);
nor U418 (N_418,N_346,N_323);
or U419 (N_419,N_345,N_397);
and U420 (N_420,N_313,N_363);
nor U421 (N_421,N_344,N_325);
or U422 (N_422,N_396,N_343);
and U423 (N_423,N_381,N_322);
or U424 (N_424,N_362,N_327);
nor U425 (N_425,N_314,N_326);
and U426 (N_426,N_300,N_385);
or U427 (N_427,N_335,N_308);
nand U428 (N_428,N_391,N_392);
nor U429 (N_429,N_336,N_365);
nor U430 (N_430,N_376,N_340);
nand U431 (N_431,N_382,N_390);
nor U432 (N_432,N_394,N_303);
nor U433 (N_433,N_374,N_373);
nor U434 (N_434,N_309,N_302);
and U435 (N_435,N_332,N_364);
nand U436 (N_436,N_305,N_347);
or U437 (N_437,N_311,N_371);
or U438 (N_438,N_386,N_310);
or U439 (N_439,N_389,N_338);
or U440 (N_440,N_367,N_348);
nor U441 (N_441,N_315,N_312);
nand U442 (N_442,N_379,N_328);
nand U443 (N_443,N_358,N_316);
or U444 (N_444,N_329,N_349);
nor U445 (N_445,N_353,N_380);
nand U446 (N_446,N_341,N_357);
and U447 (N_447,N_398,N_378);
or U448 (N_448,N_361,N_352);
nand U449 (N_449,N_369,N_355);
and U450 (N_450,N_379,N_398);
or U451 (N_451,N_314,N_360);
nor U452 (N_452,N_328,N_394);
and U453 (N_453,N_323,N_313);
nor U454 (N_454,N_327,N_353);
nor U455 (N_455,N_390,N_303);
nand U456 (N_456,N_386,N_343);
nand U457 (N_457,N_376,N_341);
or U458 (N_458,N_361,N_316);
nor U459 (N_459,N_313,N_394);
or U460 (N_460,N_394,N_382);
nor U461 (N_461,N_310,N_329);
nor U462 (N_462,N_370,N_397);
nand U463 (N_463,N_357,N_327);
nand U464 (N_464,N_348,N_312);
nor U465 (N_465,N_327,N_346);
or U466 (N_466,N_324,N_320);
and U467 (N_467,N_358,N_352);
and U468 (N_468,N_390,N_362);
or U469 (N_469,N_318,N_353);
or U470 (N_470,N_349,N_379);
nand U471 (N_471,N_383,N_318);
or U472 (N_472,N_333,N_326);
nor U473 (N_473,N_381,N_323);
xnor U474 (N_474,N_305,N_337);
and U475 (N_475,N_361,N_302);
nor U476 (N_476,N_352,N_338);
or U477 (N_477,N_331,N_347);
nor U478 (N_478,N_334,N_347);
or U479 (N_479,N_305,N_384);
and U480 (N_480,N_320,N_373);
or U481 (N_481,N_362,N_373);
nand U482 (N_482,N_344,N_380);
nor U483 (N_483,N_367,N_376);
or U484 (N_484,N_369,N_316);
or U485 (N_485,N_308,N_392);
or U486 (N_486,N_345,N_306);
or U487 (N_487,N_302,N_320);
nor U488 (N_488,N_370,N_378);
and U489 (N_489,N_339,N_303);
and U490 (N_490,N_306,N_355);
or U491 (N_491,N_390,N_398);
nor U492 (N_492,N_345,N_312);
and U493 (N_493,N_318,N_328);
and U494 (N_494,N_325,N_326);
nand U495 (N_495,N_389,N_350);
or U496 (N_496,N_394,N_374);
and U497 (N_497,N_306,N_374);
xor U498 (N_498,N_343,N_389);
and U499 (N_499,N_350,N_339);
and U500 (N_500,N_498,N_443);
nand U501 (N_501,N_462,N_427);
xnor U502 (N_502,N_473,N_464);
nor U503 (N_503,N_480,N_422);
or U504 (N_504,N_490,N_433);
nor U505 (N_505,N_456,N_405);
nor U506 (N_506,N_447,N_485);
or U507 (N_507,N_486,N_482);
or U508 (N_508,N_469,N_442);
nor U509 (N_509,N_403,N_411);
nor U510 (N_510,N_439,N_489);
or U511 (N_511,N_444,N_496);
nand U512 (N_512,N_476,N_459);
and U513 (N_513,N_461,N_457);
nor U514 (N_514,N_413,N_423);
nand U515 (N_515,N_432,N_475);
or U516 (N_516,N_468,N_494);
nand U517 (N_517,N_492,N_401);
and U518 (N_518,N_402,N_463);
and U519 (N_519,N_415,N_429);
and U520 (N_520,N_418,N_438);
xnor U521 (N_521,N_460,N_408);
nor U522 (N_522,N_410,N_488);
or U523 (N_523,N_493,N_421);
and U524 (N_524,N_449,N_465);
or U525 (N_525,N_434,N_416);
xnor U526 (N_526,N_420,N_441);
and U527 (N_527,N_454,N_446);
and U528 (N_528,N_471,N_499);
and U529 (N_529,N_445,N_406);
and U530 (N_530,N_470,N_497);
nand U531 (N_531,N_478,N_453);
nor U532 (N_532,N_412,N_440);
nand U533 (N_533,N_409,N_477);
nand U534 (N_534,N_437,N_466);
nand U535 (N_535,N_414,N_404);
or U536 (N_536,N_431,N_495);
xnor U537 (N_537,N_483,N_430);
or U538 (N_538,N_487,N_450);
or U539 (N_539,N_417,N_448);
nor U540 (N_540,N_491,N_400);
or U541 (N_541,N_426,N_435);
and U542 (N_542,N_451,N_425);
xor U543 (N_543,N_452,N_419);
nor U544 (N_544,N_481,N_407);
nor U545 (N_545,N_424,N_474);
or U546 (N_546,N_428,N_484);
nand U547 (N_547,N_458,N_472);
or U548 (N_548,N_455,N_436);
or U549 (N_549,N_467,N_479);
and U550 (N_550,N_445,N_462);
and U551 (N_551,N_425,N_424);
nor U552 (N_552,N_445,N_479);
or U553 (N_553,N_419,N_425);
nor U554 (N_554,N_498,N_414);
and U555 (N_555,N_442,N_436);
and U556 (N_556,N_412,N_434);
or U557 (N_557,N_499,N_430);
nor U558 (N_558,N_463,N_440);
and U559 (N_559,N_429,N_421);
nor U560 (N_560,N_442,N_476);
and U561 (N_561,N_460,N_431);
and U562 (N_562,N_406,N_483);
nand U563 (N_563,N_472,N_477);
nand U564 (N_564,N_406,N_436);
nand U565 (N_565,N_465,N_432);
nor U566 (N_566,N_493,N_492);
and U567 (N_567,N_455,N_470);
nand U568 (N_568,N_416,N_405);
nand U569 (N_569,N_493,N_406);
or U570 (N_570,N_440,N_447);
nor U571 (N_571,N_478,N_432);
nor U572 (N_572,N_438,N_454);
or U573 (N_573,N_447,N_431);
nand U574 (N_574,N_417,N_437);
nor U575 (N_575,N_468,N_435);
and U576 (N_576,N_414,N_418);
or U577 (N_577,N_436,N_419);
or U578 (N_578,N_437,N_406);
nor U579 (N_579,N_496,N_479);
nor U580 (N_580,N_490,N_402);
nor U581 (N_581,N_499,N_443);
xnor U582 (N_582,N_415,N_437);
and U583 (N_583,N_422,N_427);
or U584 (N_584,N_411,N_409);
and U585 (N_585,N_422,N_406);
nor U586 (N_586,N_492,N_454);
nand U587 (N_587,N_498,N_452);
and U588 (N_588,N_471,N_457);
or U589 (N_589,N_435,N_420);
or U590 (N_590,N_450,N_420);
nand U591 (N_591,N_456,N_445);
and U592 (N_592,N_490,N_438);
nand U593 (N_593,N_490,N_453);
nand U594 (N_594,N_425,N_410);
and U595 (N_595,N_447,N_477);
nor U596 (N_596,N_496,N_487);
nor U597 (N_597,N_417,N_456);
or U598 (N_598,N_459,N_454);
nor U599 (N_599,N_477,N_431);
nor U600 (N_600,N_567,N_584);
nor U601 (N_601,N_528,N_576);
and U602 (N_602,N_583,N_589);
xor U603 (N_603,N_562,N_557);
nand U604 (N_604,N_526,N_530);
nand U605 (N_605,N_599,N_561);
nand U606 (N_606,N_553,N_534);
nor U607 (N_607,N_594,N_560);
and U608 (N_608,N_596,N_586);
or U609 (N_609,N_558,N_598);
nand U610 (N_610,N_537,N_552);
and U611 (N_611,N_542,N_536);
nand U612 (N_612,N_521,N_554);
or U613 (N_613,N_514,N_535);
or U614 (N_614,N_590,N_538);
or U615 (N_615,N_506,N_578);
nor U616 (N_616,N_579,N_540);
nor U617 (N_617,N_575,N_585);
or U618 (N_618,N_597,N_513);
nand U619 (N_619,N_520,N_593);
and U620 (N_620,N_518,N_574);
nand U621 (N_621,N_570,N_588);
nand U622 (N_622,N_551,N_582);
or U623 (N_623,N_500,N_503);
nor U624 (N_624,N_523,N_507);
and U625 (N_625,N_501,N_572);
or U626 (N_626,N_529,N_548);
nand U627 (N_627,N_512,N_546);
nor U628 (N_628,N_522,N_533);
nor U629 (N_629,N_564,N_510);
and U630 (N_630,N_580,N_527);
nor U631 (N_631,N_541,N_504);
nand U632 (N_632,N_563,N_555);
and U633 (N_633,N_524,N_559);
nand U634 (N_634,N_544,N_549);
or U635 (N_635,N_550,N_566);
or U636 (N_636,N_505,N_509);
nand U637 (N_637,N_543,N_591);
nand U638 (N_638,N_515,N_532);
nand U639 (N_639,N_545,N_569);
nand U640 (N_640,N_519,N_508);
and U641 (N_641,N_573,N_577);
or U642 (N_642,N_565,N_568);
nand U643 (N_643,N_516,N_592);
and U644 (N_644,N_502,N_581);
or U645 (N_645,N_556,N_595);
and U646 (N_646,N_539,N_531);
and U647 (N_647,N_547,N_587);
or U648 (N_648,N_525,N_517);
or U649 (N_649,N_511,N_571);
or U650 (N_650,N_568,N_503);
and U651 (N_651,N_565,N_544);
nor U652 (N_652,N_574,N_508);
nor U653 (N_653,N_576,N_561);
nor U654 (N_654,N_556,N_536);
or U655 (N_655,N_546,N_534);
or U656 (N_656,N_524,N_567);
and U657 (N_657,N_586,N_574);
and U658 (N_658,N_550,N_575);
and U659 (N_659,N_580,N_551);
nand U660 (N_660,N_568,N_537);
nor U661 (N_661,N_541,N_536);
or U662 (N_662,N_506,N_552);
nand U663 (N_663,N_505,N_586);
and U664 (N_664,N_553,N_596);
nand U665 (N_665,N_588,N_549);
and U666 (N_666,N_516,N_570);
or U667 (N_667,N_540,N_560);
or U668 (N_668,N_598,N_574);
nor U669 (N_669,N_546,N_547);
or U670 (N_670,N_532,N_581);
nand U671 (N_671,N_583,N_529);
and U672 (N_672,N_553,N_514);
nor U673 (N_673,N_585,N_518);
or U674 (N_674,N_518,N_510);
or U675 (N_675,N_527,N_591);
nand U676 (N_676,N_574,N_562);
nand U677 (N_677,N_581,N_539);
and U678 (N_678,N_563,N_588);
nor U679 (N_679,N_557,N_554);
nand U680 (N_680,N_520,N_565);
nand U681 (N_681,N_597,N_598);
nand U682 (N_682,N_599,N_522);
nor U683 (N_683,N_564,N_532);
nand U684 (N_684,N_500,N_596);
and U685 (N_685,N_594,N_534);
nor U686 (N_686,N_591,N_530);
nor U687 (N_687,N_557,N_580);
nand U688 (N_688,N_548,N_579);
nor U689 (N_689,N_551,N_563);
and U690 (N_690,N_522,N_574);
nand U691 (N_691,N_558,N_570);
and U692 (N_692,N_580,N_546);
or U693 (N_693,N_595,N_500);
xnor U694 (N_694,N_599,N_542);
nor U695 (N_695,N_534,N_501);
and U696 (N_696,N_555,N_539);
nor U697 (N_697,N_554,N_504);
and U698 (N_698,N_558,N_599);
nand U699 (N_699,N_544,N_587);
nand U700 (N_700,N_648,N_680);
nor U701 (N_701,N_691,N_692);
nor U702 (N_702,N_687,N_670);
or U703 (N_703,N_686,N_678);
nand U704 (N_704,N_662,N_673);
nor U705 (N_705,N_654,N_649);
nor U706 (N_706,N_682,N_659);
and U707 (N_707,N_628,N_675);
and U708 (N_708,N_631,N_641);
and U709 (N_709,N_634,N_650);
nor U710 (N_710,N_610,N_636);
nand U711 (N_711,N_617,N_685);
xor U712 (N_712,N_644,N_665);
nand U713 (N_713,N_616,N_622);
and U714 (N_714,N_602,N_653);
or U715 (N_715,N_656,N_619);
or U716 (N_716,N_633,N_642);
or U717 (N_717,N_613,N_611);
and U718 (N_718,N_698,N_629);
and U719 (N_719,N_626,N_679);
nand U720 (N_720,N_647,N_690);
nor U721 (N_721,N_621,N_651);
nand U722 (N_722,N_681,N_620);
nand U723 (N_723,N_693,N_625);
or U724 (N_724,N_661,N_612);
nor U725 (N_725,N_601,N_624);
and U726 (N_726,N_676,N_614);
and U727 (N_727,N_635,N_606);
and U728 (N_728,N_605,N_689);
nand U729 (N_729,N_630,N_674);
or U730 (N_730,N_639,N_655);
nand U731 (N_731,N_652,N_669);
and U732 (N_732,N_668,N_608);
nand U733 (N_733,N_677,N_632);
or U734 (N_734,N_618,N_696);
and U735 (N_735,N_640,N_663);
or U736 (N_736,N_609,N_615);
and U737 (N_737,N_660,N_695);
nor U738 (N_738,N_688,N_643);
or U739 (N_739,N_694,N_667);
nand U740 (N_740,N_666,N_684);
nor U741 (N_741,N_657,N_646);
nor U742 (N_742,N_683,N_623);
nand U743 (N_743,N_627,N_645);
or U744 (N_744,N_672,N_638);
and U745 (N_745,N_600,N_637);
and U746 (N_746,N_658,N_603);
and U747 (N_747,N_697,N_699);
nand U748 (N_748,N_604,N_607);
nor U749 (N_749,N_664,N_671);
and U750 (N_750,N_629,N_675);
or U751 (N_751,N_623,N_636);
or U752 (N_752,N_633,N_690);
or U753 (N_753,N_679,N_692);
and U754 (N_754,N_692,N_662);
or U755 (N_755,N_688,N_604);
xor U756 (N_756,N_608,N_629);
nor U757 (N_757,N_672,N_656);
xor U758 (N_758,N_621,N_608);
nor U759 (N_759,N_677,N_636);
nand U760 (N_760,N_653,N_624);
or U761 (N_761,N_651,N_697);
and U762 (N_762,N_685,N_615);
nor U763 (N_763,N_650,N_637);
or U764 (N_764,N_690,N_695);
nand U765 (N_765,N_646,N_679);
nor U766 (N_766,N_609,N_638);
or U767 (N_767,N_601,N_637);
or U768 (N_768,N_688,N_611);
or U769 (N_769,N_662,N_682);
nand U770 (N_770,N_621,N_668);
nand U771 (N_771,N_670,N_603);
or U772 (N_772,N_671,N_654);
and U773 (N_773,N_685,N_690);
or U774 (N_774,N_627,N_654);
nor U775 (N_775,N_625,N_682);
nor U776 (N_776,N_639,N_651);
nor U777 (N_777,N_622,N_620);
nor U778 (N_778,N_672,N_614);
or U779 (N_779,N_669,N_662);
or U780 (N_780,N_660,N_611);
nand U781 (N_781,N_614,N_621);
or U782 (N_782,N_623,N_628);
or U783 (N_783,N_614,N_646);
and U784 (N_784,N_641,N_642);
nand U785 (N_785,N_687,N_626);
and U786 (N_786,N_657,N_639);
nand U787 (N_787,N_667,N_665);
and U788 (N_788,N_698,N_628);
or U789 (N_789,N_608,N_637);
nand U790 (N_790,N_661,N_665);
nor U791 (N_791,N_688,N_629);
nand U792 (N_792,N_604,N_662);
and U793 (N_793,N_604,N_682);
or U794 (N_794,N_665,N_606);
nor U795 (N_795,N_622,N_688);
nor U796 (N_796,N_610,N_658);
nor U797 (N_797,N_607,N_628);
and U798 (N_798,N_668,N_674);
and U799 (N_799,N_614,N_620);
nor U800 (N_800,N_740,N_792);
nand U801 (N_801,N_758,N_736);
and U802 (N_802,N_782,N_733);
and U803 (N_803,N_716,N_788);
nand U804 (N_804,N_710,N_738);
nor U805 (N_805,N_720,N_722);
or U806 (N_806,N_790,N_791);
nor U807 (N_807,N_754,N_727);
nand U808 (N_808,N_701,N_771);
nor U809 (N_809,N_753,N_730);
or U810 (N_810,N_703,N_770);
or U811 (N_811,N_749,N_763);
nor U812 (N_812,N_746,N_717);
and U813 (N_813,N_793,N_715);
nor U814 (N_814,N_704,N_728);
or U815 (N_815,N_748,N_724);
and U816 (N_816,N_777,N_744);
nor U817 (N_817,N_797,N_712);
nand U818 (N_818,N_775,N_789);
nand U819 (N_819,N_751,N_762);
and U820 (N_820,N_774,N_742);
nand U821 (N_821,N_784,N_734);
nand U822 (N_822,N_713,N_798);
nor U823 (N_823,N_769,N_708);
nor U824 (N_824,N_706,N_779);
and U825 (N_825,N_781,N_709);
nand U826 (N_826,N_755,N_757);
or U827 (N_827,N_761,N_765);
xor U828 (N_828,N_783,N_795);
nand U829 (N_829,N_756,N_707);
nor U830 (N_830,N_787,N_747);
and U831 (N_831,N_726,N_773);
and U832 (N_832,N_731,N_711);
nand U833 (N_833,N_718,N_776);
and U834 (N_834,N_772,N_786);
nand U835 (N_835,N_767,N_741);
nor U836 (N_836,N_732,N_725);
or U837 (N_837,N_729,N_745);
or U838 (N_838,N_737,N_723);
and U839 (N_839,N_735,N_760);
or U840 (N_840,N_794,N_785);
nor U841 (N_841,N_764,N_721);
and U842 (N_842,N_768,N_799);
and U843 (N_843,N_766,N_705);
or U844 (N_844,N_743,N_759);
nand U845 (N_845,N_739,N_778);
or U846 (N_846,N_700,N_752);
nor U847 (N_847,N_796,N_780);
or U848 (N_848,N_702,N_714);
and U849 (N_849,N_719,N_750);
and U850 (N_850,N_760,N_759);
nand U851 (N_851,N_736,N_720);
and U852 (N_852,N_763,N_772);
nor U853 (N_853,N_705,N_715);
nor U854 (N_854,N_742,N_795);
or U855 (N_855,N_709,N_741);
and U856 (N_856,N_732,N_703);
nor U857 (N_857,N_706,N_799);
nor U858 (N_858,N_758,N_711);
nand U859 (N_859,N_788,N_770);
nand U860 (N_860,N_763,N_755);
nand U861 (N_861,N_769,N_707);
xnor U862 (N_862,N_738,N_705);
xnor U863 (N_863,N_777,N_738);
nand U864 (N_864,N_774,N_701);
and U865 (N_865,N_737,N_731);
nor U866 (N_866,N_772,N_729);
and U867 (N_867,N_704,N_772);
or U868 (N_868,N_726,N_779);
nand U869 (N_869,N_729,N_715);
or U870 (N_870,N_774,N_770);
or U871 (N_871,N_755,N_782);
or U872 (N_872,N_702,N_746);
nand U873 (N_873,N_708,N_794);
and U874 (N_874,N_777,N_724);
nand U875 (N_875,N_795,N_734);
or U876 (N_876,N_779,N_782);
nor U877 (N_877,N_714,N_734);
nor U878 (N_878,N_771,N_715);
nor U879 (N_879,N_725,N_723);
nor U880 (N_880,N_769,N_780);
nand U881 (N_881,N_787,N_715);
nor U882 (N_882,N_734,N_716);
xnor U883 (N_883,N_752,N_717);
and U884 (N_884,N_732,N_724);
nand U885 (N_885,N_746,N_727);
nand U886 (N_886,N_710,N_773);
and U887 (N_887,N_798,N_799);
and U888 (N_888,N_706,N_736);
or U889 (N_889,N_730,N_739);
and U890 (N_890,N_717,N_765);
nand U891 (N_891,N_768,N_797);
and U892 (N_892,N_783,N_706);
nand U893 (N_893,N_761,N_778);
nand U894 (N_894,N_707,N_736);
xnor U895 (N_895,N_787,N_768);
nand U896 (N_896,N_755,N_788);
nand U897 (N_897,N_769,N_702);
and U898 (N_898,N_739,N_776);
and U899 (N_899,N_781,N_765);
nor U900 (N_900,N_841,N_808);
nand U901 (N_901,N_804,N_839);
or U902 (N_902,N_857,N_848);
nor U903 (N_903,N_893,N_881);
or U904 (N_904,N_856,N_896);
nor U905 (N_905,N_803,N_878);
and U906 (N_906,N_880,N_888);
and U907 (N_907,N_897,N_860);
and U908 (N_908,N_817,N_879);
nor U909 (N_909,N_894,N_832);
nor U910 (N_910,N_821,N_886);
or U911 (N_911,N_852,N_871);
nor U912 (N_912,N_830,N_831);
or U913 (N_913,N_868,N_887);
nor U914 (N_914,N_835,N_855);
and U915 (N_915,N_874,N_800);
nand U916 (N_916,N_849,N_838);
nor U917 (N_917,N_812,N_809);
or U918 (N_918,N_826,N_869);
nor U919 (N_919,N_811,N_819);
or U920 (N_920,N_890,N_864);
and U921 (N_921,N_867,N_847);
nand U922 (N_922,N_820,N_875);
or U923 (N_923,N_845,N_814);
or U924 (N_924,N_873,N_810);
nor U925 (N_925,N_807,N_805);
nand U926 (N_926,N_863,N_854);
nand U927 (N_927,N_824,N_823);
and U928 (N_928,N_891,N_840);
or U929 (N_929,N_844,N_843);
or U930 (N_930,N_883,N_859);
nor U931 (N_931,N_895,N_815);
nor U932 (N_932,N_806,N_861);
or U933 (N_933,N_837,N_850);
nor U934 (N_934,N_889,N_884);
nor U935 (N_935,N_834,N_828);
nand U936 (N_936,N_829,N_892);
nor U937 (N_937,N_899,N_872);
nand U938 (N_938,N_825,N_836);
or U939 (N_939,N_862,N_818);
and U940 (N_940,N_816,N_802);
or U941 (N_941,N_877,N_822);
nor U942 (N_942,N_898,N_882);
nor U943 (N_943,N_851,N_858);
xnor U944 (N_944,N_801,N_846);
nand U945 (N_945,N_833,N_813);
and U946 (N_946,N_866,N_876);
and U947 (N_947,N_865,N_885);
nand U948 (N_948,N_842,N_827);
and U949 (N_949,N_853,N_870);
nand U950 (N_950,N_874,N_811);
nand U951 (N_951,N_847,N_814);
or U952 (N_952,N_871,N_886);
and U953 (N_953,N_870,N_806);
nor U954 (N_954,N_828,N_868);
nor U955 (N_955,N_865,N_857);
or U956 (N_956,N_845,N_883);
nor U957 (N_957,N_855,N_850);
or U958 (N_958,N_808,N_844);
or U959 (N_959,N_809,N_893);
nor U960 (N_960,N_857,N_809);
nand U961 (N_961,N_849,N_815);
nand U962 (N_962,N_863,N_820);
and U963 (N_963,N_874,N_872);
nor U964 (N_964,N_835,N_881);
nand U965 (N_965,N_839,N_888);
or U966 (N_966,N_842,N_894);
and U967 (N_967,N_809,N_890);
or U968 (N_968,N_834,N_887);
nand U969 (N_969,N_874,N_879);
and U970 (N_970,N_876,N_865);
and U971 (N_971,N_888,N_831);
and U972 (N_972,N_801,N_805);
nand U973 (N_973,N_804,N_820);
xnor U974 (N_974,N_830,N_879);
or U975 (N_975,N_804,N_816);
or U976 (N_976,N_841,N_847);
nand U977 (N_977,N_819,N_820);
nand U978 (N_978,N_824,N_825);
xnor U979 (N_979,N_890,N_842);
nor U980 (N_980,N_892,N_834);
or U981 (N_981,N_864,N_828);
xor U982 (N_982,N_821,N_875);
nor U983 (N_983,N_880,N_884);
nand U984 (N_984,N_862,N_864);
or U985 (N_985,N_814,N_840);
nor U986 (N_986,N_861,N_886);
and U987 (N_987,N_881,N_840);
nand U988 (N_988,N_850,N_892);
and U989 (N_989,N_803,N_823);
nor U990 (N_990,N_858,N_883);
or U991 (N_991,N_818,N_883);
or U992 (N_992,N_881,N_858);
or U993 (N_993,N_817,N_877);
nand U994 (N_994,N_843,N_840);
or U995 (N_995,N_852,N_806);
nor U996 (N_996,N_860,N_853);
nand U997 (N_997,N_832,N_841);
and U998 (N_998,N_860,N_868);
and U999 (N_999,N_811,N_844);
or U1000 (N_1000,N_920,N_923);
and U1001 (N_1001,N_903,N_970);
and U1002 (N_1002,N_961,N_984);
and U1003 (N_1003,N_988,N_940);
and U1004 (N_1004,N_965,N_992);
nand U1005 (N_1005,N_939,N_932);
nand U1006 (N_1006,N_927,N_914);
and U1007 (N_1007,N_929,N_958);
nor U1008 (N_1008,N_919,N_987);
and U1009 (N_1009,N_971,N_983);
nand U1010 (N_1010,N_900,N_922);
or U1011 (N_1011,N_933,N_948);
and U1012 (N_1012,N_925,N_980);
or U1013 (N_1013,N_996,N_935);
nand U1014 (N_1014,N_915,N_976);
nand U1015 (N_1015,N_989,N_964);
nor U1016 (N_1016,N_957,N_966);
or U1017 (N_1017,N_978,N_917);
nand U1018 (N_1018,N_951,N_913);
or U1019 (N_1019,N_930,N_934);
or U1020 (N_1020,N_959,N_902);
or U1021 (N_1021,N_931,N_995);
and U1022 (N_1022,N_991,N_999);
or U1023 (N_1023,N_946,N_904);
nand U1024 (N_1024,N_993,N_955);
or U1025 (N_1025,N_928,N_985);
xor U1026 (N_1026,N_936,N_977);
or U1027 (N_1027,N_947,N_963);
or U1028 (N_1028,N_906,N_938);
nor U1029 (N_1029,N_911,N_990);
or U1030 (N_1030,N_979,N_908);
or U1031 (N_1031,N_944,N_952);
or U1032 (N_1032,N_973,N_907);
nand U1033 (N_1033,N_997,N_975);
nor U1034 (N_1034,N_972,N_954);
and U1035 (N_1035,N_967,N_960);
and U1036 (N_1036,N_945,N_998);
nor U1037 (N_1037,N_937,N_916);
or U1038 (N_1038,N_969,N_949);
nand U1039 (N_1039,N_943,N_912);
nand U1040 (N_1040,N_981,N_909);
nor U1041 (N_1041,N_910,N_921);
or U1042 (N_1042,N_982,N_926);
or U1043 (N_1043,N_942,N_974);
nand U1044 (N_1044,N_924,N_901);
or U1045 (N_1045,N_994,N_941);
and U1046 (N_1046,N_956,N_905);
nand U1047 (N_1047,N_918,N_986);
and U1048 (N_1048,N_968,N_950);
and U1049 (N_1049,N_953,N_962);
nand U1050 (N_1050,N_945,N_994);
nand U1051 (N_1051,N_936,N_906);
and U1052 (N_1052,N_974,N_997);
or U1053 (N_1053,N_959,N_929);
or U1054 (N_1054,N_925,N_991);
or U1055 (N_1055,N_984,N_915);
nor U1056 (N_1056,N_961,N_930);
nor U1057 (N_1057,N_909,N_928);
nor U1058 (N_1058,N_911,N_949);
nand U1059 (N_1059,N_903,N_926);
nand U1060 (N_1060,N_907,N_948);
nor U1061 (N_1061,N_952,N_984);
or U1062 (N_1062,N_933,N_978);
nand U1063 (N_1063,N_965,N_963);
and U1064 (N_1064,N_961,N_901);
nor U1065 (N_1065,N_965,N_948);
and U1066 (N_1066,N_992,N_908);
nor U1067 (N_1067,N_990,N_922);
nor U1068 (N_1068,N_924,N_932);
nor U1069 (N_1069,N_966,N_920);
or U1070 (N_1070,N_919,N_938);
nand U1071 (N_1071,N_966,N_931);
and U1072 (N_1072,N_977,N_970);
nand U1073 (N_1073,N_963,N_967);
nand U1074 (N_1074,N_967,N_968);
nor U1075 (N_1075,N_951,N_996);
and U1076 (N_1076,N_954,N_926);
or U1077 (N_1077,N_998,N_926);
or U1078 (N_1078,N_979,N_916);
and U1079 (N_1079,N_929,N_985);
nor U1080 (N_1080,N_945,N_926);
nand U1081 (N_1081,N_934,N_920);
and U1082 (N_1082,N_967,N_932);
nor U1083 (N_1083,N_939,N_968);
or U1084 (N_1084,N_995,N_939);
and U1085 (N_1085,N_908,N_924);
or U1086 (N_1086,N_912,N_971);
and U1087 (N_1087,N_909,N_919);
or U1088 (N_1088,N_966,N_982);
or U1089 (N_1089,N_960,N_959);
nor U1090 (N_1090,N_974,N_923);
or U1091 (N_1091,N_939,N_983);
and U1092 (N_1092,N_904,N_976);
nand U1093 (N_1093,N_963,N_979);
and U1094 (N_1094,N_975,N_967);
nor U1095 (N_1095,N_914,N_972);
or U1096 (N_1096,N_925,N_985);
nor U1097 (N_1097,N_900,N_907);
or U1098 (N_1098,N_987,N_932);
nor U1099 (N_1099,N_945,N_962);
nand U1100 (N_1100,N_1055,N_1006);
nand U1101 (N_1101,N_1079,N_1018);
and U1102 (N_1102,N_1014,N_1071);
and U1103 (N_1103,N_1099,N_1066);
or U1104 (N_1104,N_1052,N_1035);
nor U1105 (N_1105,N_1008,N_1026);
or U1106 (N_1106,N_1027,N_1067);
nor U1107 (N_1107,N_1029,N_1019);
or U1108 (N_1108,N_1059,N_1046);
xnor U1109 (N_1109,N_1047,N_1017);
or U1110 (N_1110,N_1013,N_1085);
and U1111 (N_1111,N_1009,N_1070);
nand U1112 (N_1112,N_1075,N_1060);
and U1113 (N_1113,N_1022,N_1076);
and U1114 (N_1114,N_1012,N_1042);
nand U1115 (N_1115,N_1041,N_1040);
and U1116 (N_1116,N_1084,N_1053);
nor U1117 (N_1117,N_1010,N_1030);
nand U1118 (N_1118,N_1078,N_1034);
or U1119 (N_1119,N_1000,N_1096);
and U1120 (N_1120,N_1045,N_1043);
or U1121 (N_1121,N_1083,N_1089);
nand U1122 (N_1122,N_1048,N_1033);
or U1123 (N_1123,N_1069,N_1001);
nand U1124 (N_1124,N_1011,N_1020);
nand U1125 (N_1125,N_1028,N_1090);
nor U1126 (N_1126,N_1056,N_1050);
nand U1127 (N_1127,N_1088,N_1098);
nor U1128 (N_1128,N_1072,N_1038);
nand U1129 (N_1129,N_1080,N_1095);
or U1130 (N_1130,N_1016,N_1062);
nand U1131 (N_1131,N_1074,N_1064);
and U1132 (N_1132,N_1049,N_1024);
nand U1133 (N_1133,N_1073,N_1002);
nand U1134 (N_1134,N_1093,N_1086);
nor U1135 (N_1135,N_1058,N_1021);
nand U1136 (N_1136,N_1054,N_1032);
and U1137 (N_1137,N_1007,N_1057);
and U1138 (N_1138,N_1051,N_1077);
and U1139 (N_1139,N_1094,N_1023);
nand U1140 (N_1140,N_1036,N_1063);
nor U1141 (N_1141,N_1039,N_1081);
nor U1142 (N_1142,N_1015,N_1092);
nor U1143 (N_1143,N_1097,N_1044);
and U1144 (N_1144,N_1025,N_1037);
nand U1145 (N_1145,N_1087,N_1004);
nor U1146 (N_1146,N_1065,N_1061);
or U1147 (N_1147,N_1031,N_1068);
or U1148 (N_1148,N_1091,N_1005);
and U1149 (N_1149,N_1082,N_1003);
nor U1150 (N_1150,N_1068,N_1008);
or U1151 (N_1151,N_1040,N_1061);
nor U1152 (N_1152,N_1096,N_1002);
or U1153 (N_1153,N_1049,N_1019);
or U1154 (N_1154,N_1032,N_1047);
nand U1155 (N_1155,N_1084,N_1018);
and U1156 (N_1156,N_1045,N_1071);
nand U1157 (N_1157,N_1062,N_1083);
nand U1158 (N_1158,N_1027,N_1031);
nor U1159 (N_1159,N_1066,N_1064);
and U1160 (N_1160,N_1075,N_1017);
or U1161 (N_1161,N_1090,N_1042);
nor U1162 (N_1162,N_1032,N_1024);
nand U1163 (N_1163,N_1087,N_1082);
nand U1164 (N_1164,N_1057,N_1081);
nor U1165 (N_1165,N_1064,N_1008);
or U1166 (N_1166,N_1079,N_1068);
and U1167 (N_1167,N_1015,N_1035);
or U1168 (N_1168,N_1020,N_1071);
xor U1169 (N_1169,N_1081,N_1085);
nor U1170 (N_1170,N_1095,N_1083);
and U1171 (N_1171,N_1030,N_1027);
nand U1172 (N_1172,N_1038,N_1069);
nor U1173 (N_1173,N_1016,N_1054);
nor U1174 (N_1174,N_1027,N_1066);
and U1175 (N_1175,N_1093,N_1097);
or U1176 (N_1176,N_1061,N_1006);
or U1177 (N_1177,N_1074,N_1072);
nand U1178 (N_1178,N_1014,N_1021);
nor U1179 (N_1179,N_1047,N_1050);
and U1180 (N_1180,N_1029,N_1079);
and U1181 (N_1181,N_1008,N_1017);
and U1182 (N_1182,N_1005,N_1067);
nor U1183 (N_1183,N_1050,N_1035);
or U1184 (N_1184,N_1047,N_1065);
and U1185 (N_1185,N_1042,N_1071);
xnor U1186 (N_1186,N_1031,N_1029);
nand U1187 (N_1187,N_1041,N_1096);
and U1188 (N_1188,N_1071,N_1007);
nand U1189 (N_1189,N_1001,N_1007);
or U1190 (N_1190,N_1002,N_1072);
nor U1191 (N_1191,N_1051,N_1014);
nor U1192 (N_1192,N_1074,N_1019);
or U1193 (N_1193,N_1088,N_1077);
and U1194 (N_1194,N_1017,N_1003);
nor U1195 (N_1195,N_1073,N_1030);
and U1196 (N_1196,N_1087,N_1083);
nand U1197 (N_1197,N_1060,N_1016);
nor U1198 (N_1198,N_1044,N_1096);
and U1199 (N_1199,N_1006,N_1012);
and U1200 (N_1200,N_1186,N_1155);
and U1201 (N_1201,N_1184,N_1181);
nor U1202 (N_1202,N_1172,N_1177);
nor U1203 (N_1203,N_1183,N_1118);
xor U1204 (N_1204,N_1126,N_1137);
or U1205 (N_1205,N_1125,N_1180);
nand U1206 (N_1206,N_1107,N_1197);
or U1207 (N_1207,N_1147,N_1112);
nor U1208 (N_1208,N_1193,N_1136);
nand U1209 (N_1209,N_1129,N_1100);
and U1210 (N_1210,N_1128,N_1162);
nand U1211 (N_1211,N_1161,N_1166);
or U1212 (N_1212,N_1171,N_1173);
nand U1213 (N_1213,N_1108,N_1159);
or U1214 (N_1214,N_1116,N_1148);
and U1215 (N_1215,N_1157,N_1160);
or U1216 (N_1216,N_1105,N_1185);
nor U1217 (N_1217,N_1135,N_1110);
and U1218 (N_1218,N_1111,N_1130);
nor U1219 (N_1219,N_1153,N_1131);
xor U1220 (N_1220,N_1187,N_1117);
xnor U1221 (N_1221,N_1182,N_1124);
and U1222 (N_1222,N_1199,N_1164);
nor U1223 (N_1223,N_1127,N_1134);
and U1224 (N_1224,N_1119,N_1176);
nor U1225 (N_1225,N_1150,N_1158);
or U1226 (N_1226,N_1138,N_1156);
and U1227 (N_1227,N_1152,N_1190);
or U1228 (N_1228,N_1188,N_1175);
nand U1229 (N_1229,N_1149,N_1146);
and U1230 (N_1230,N_1192,N_1113);
nor U1231 (N_1231,N_1103,N_1106);
nand U1232 (N_1232,N_1168,N_1114);
or U1233 (N_1233,N_1109,N_1133);
nor U1234 (N_1234,N_1196,N_1169);
and U1235 (N_1235,N_1179,N_1121);
nand U1236 (N_1236,N_1154,N_1143);
or U1237 (N_1237,N_1115,N_1151);
and U1238 (N_1238,N_1123,N_1189);
nand U1239 (N_1239,N_1167,N_1198);
nand U1240 (N_1240,N_1191,N_1163);
or U1241 (N_1241,N_1140,N_1165);
nand U1242 (N_1242,N_1144,N_1122);
or U1243 (N_1243,N_1195,N_1101);
nor U1244 (N_1244,N_1102,N_1178);
nand U1245 (N_1245,N_1174,N_1120);
or U1246 (N_1246,N_1145,N_1139);
and U1247 (N_1247,N_1104,N_1142);
nor U1248 (N_1248,N_1132,N_1141);
and U1249 (N_1249,N_1170,N_1194);
nand U1250 (N_1250,N_1102,N_1188);
nor U1251 (N_1251,N_1187,N_1156);
or U1252 (N_1252,N_1103,N_1151);
nor U1253 (N_1253,N_1196,N_1127);
and U1254 (N_1254,N_1161,N_1132);
and U1255 (N_1255,N_1126,N_1123);
or U1256 (N_1256,N_1181,N_1105);
nand U1257 (N_1257,N_1193,N_1156);
nor U1258 (N_1258,N_1159,N_1100);
nor U1259 (N_1259,N_1181,N_1192);
nand U1260 (N_1260,N_1155,N_1178);
or U1261 (N_1261,N_1120,N_1109);
and U1262 (N_1262,N_1158,N_1160);
nor U1263 (N_1263,N_1195,N_1178);
xnor U1264 (N_1264,N_1131,N_1190);
nand U1265 (N_1265,N_1104,N_1148);
nand U1266 (N_1266,N_1100,N_1162);
nor U1267 (N_1267,N_1101,N_1149);
nand U1268 (N_1268,N_1179,N_1150);
nand U1269 (N_1269,N_1149,N_1197);
or U1270 (N_1270,N_1111,N_1138);
nand U1271 (N_1271,N_1122,N_1197);
nor U1272 (N_1272,N_1155,N_1100);
nor U1273 (N_1273,N_1128,N_1115);
nor U1274 (N_1274,N_1150,N_1168);
nor U1275 (N_1275,N_1120,N_1106);
or U1276 (N_1276,N_1143,N_1128);
nand U1277 (N_1277,N_1181,N_1107);
nor U1278 (N_1278,N_1143,N_1119);
and U1279 (N_1279,N_1195,N_1189);
nand U1280 (N_1280,N_1140,N_1102);
and U1281 (N_1281,N_1115,N_1167);
xor U1282 (N_1282,N_1196,N_1149);
nand U1283 (N_1283,N_1149,N_1133);
xor U1284 (N_1284,N_1132,N_1138);
and U1285 (N_1285,N_1129,N_1165);
and U1286 (N_1286,N_1154,N_1108);
nand U1287 (N_1287,N_1155,N_1142);
or U1288 (N_1288,N_1142,N_1149);
and U1289 (N_1289,N_1175,N_1153);
nand U1290 (N_1290,N_1190,N_1166);
nand U1291 (N_1291,N_1186,N_1113);
and U1292 (N_1292,N_1127,N_1132);
xor U1293 (N_1293,N_1199,N_1125);
or U1294 (N_1294,N_1157,N_1178);
nor U1295 (N_1295,N_1142,N_1160);
nand U1296 (N_1296,N_1109,N_1100);
nand U1297 (N_1297,N_1121,N_1196);
xnor U1298 (N_1298,N_1141,N_1144);
and U1299 (N_1299,N_1119,N_1179);
nand U1300 (N_1300,N_1260,N_1206);
nor U1301 (N_1301,N_1249,N_1225);
or U1302 (N_1302,N_1282,N_1229);
and U1303 (N_1303,N_1236,N_1237);
or U1304 (N_1304,N_1240,N_1241);
nand U1305 (N_1305,N_1271,N_1273);
or U1306 (N_1306,N_1264,N_1278);
or U1307 (N_1307,N_1294,N_1275);
and U1308 (N_1308,N_1297,N_1277);
nand U1309 (N_1309,N_1286,N_1285);
or U1310 (N_1310,N_1203,N_1268);
and U1311 (N_1311,N_1212,N_1270);
and U1312 (N_1312,N_1215,N_1257);
or U1313 (N_1313,N_1214,N_1258);
nor U1314 (N_1314,N_1266,N_1228);
or U1315 (N_1315,N_1205,N_1287);
or U1316 (N_1316,N_1247,N_1265);
or U1317 (N_1317,N_1243,N_1220);
or U1318 (N_1318,N_1224,N_1256);
nor U1319 (N_1319,N_1250,N_1289);
nor U1320 (N_1320,N_1202,N_1284);
nand U1321 (N_1321,N_1218,N_1252);
nand U1322 (N_1322,N_1255,N_1232);
nor U1323 (N_1323,N_1242,N_1292);
and U1324 (N_1324,N_1269,N_1295);
and U1325 (N_1325,N_1227,N_1239);
nor U1326 (N_1326,N_1245,N_1204);
xnor U1327 (N_1327,N_1274,N_1261);
or U1328 (N_1328,N_1222,N_1221);
or U1329 (N_1329,N_1230,N_1235);
nand U1330 (N_1330,N_1234,N_1290);
nand U1331 (N_1331,N_1226,N_1211);
and U1332 (N_1332,N_1254,N_1251);
or U1333 (N_1333,N_1219,N_1281);
nor U1334 (N_1334,N_1248,N_1207);
and U1335 (N_1335,N_1210,N_1262);
and U1336 (N_1336,N_1208,N_1213);
nand U1337 (N_1337,N_1296,N_1209);
nor U1338 (N_1338,N_1231,N_1216);
nor U1339 (N_1339,N_1233,N_1246);
or U1340 (N_1340,N_1223,N_1291);
xor U1341 (N_1341,N_1280,N_1272);
nor U1342 (N_1342,N_1283,N_1298);
and U1343 (N_1343,N_1244,N_1238);
nand U1344 (N_1344,N_1263,N_1267);
or U1345 (N_1345,N_1201,N_1299);
and U1346 (N_1346,N_1217,N_1200);
nor U1347 (N_1347,N_1288,N_1276);
nand U1348 (N_1348,N_1259,N_1253);
nand U1349 (N_1349,N_1279,N_1293);
nor U1350 (N_1350,N_1213,N_1283);
nand U1351 (N_1351,N_1255,N_1226);
and U1352 (N_1352,N_1271,N_1266);
or U1353 (N_1353,N_1298,N_1225);
and U1354 (N_1354,N_1275,N_1254);
or U1355 (N_1355,N_1291,N_1265);
xnor U1356 (N_1356,N_1248,N_1282);
or U1357 (N_1357,N_1286,N_1202);
or U1358 (N_1358,N_1211,N_1288);
or U1359 (N_1359,N_1264,N_1288);
nor U1360 (N_1360,N_1201,N_1210);
or U1361 (N_1361,N_1223,N_1298);
nor U1362 (N_1362,N_1261,N_1255);
or U1363 (N_1363,N_1271,N_1235);
or U1364 (N_1364,N_1237,N_1243);
and U1365 (N_1365,N_1222,N_1278);
and U1366 (N_1366,N_1273,N_1269);
nor U1367 (N_1367,N_1278,N_1219);
nor U1368 (N_1368,N_1289,N_1277);
nor U1369 (N_1369,N_1227,N_1266);
or U1370 (N_1370,N_1214,N_1206);
nor U1371 (N_1371,N_1296,N_1232);
nor U1372 (N_1372,N_1286,N_1233);
or U1373 (N_1373,N_1203,N_1274);
nand U1374 (N_1374,N_1267,N_1210);
and U1375 (N_1375,N_1283,N_1235);
or U1376 (N_1376,N_1286,N_1215);
and U1377 (N_1377,N_1202,N_1238);
and U1378 (N_1378,N_1212,N_1296);
nand U1379 (N_1379,N_1239,N_1217);
and U1380 (N_1380,N_1250,N_1230);
nor U1381 (N_1381,N_1248,N_1201);
and U1382 (N_1382,N_1231,N_1272);
nor U1383 (N_1383,N_1232,N_1259);
xnor U1384 (N_1384,N_1277,N_1233);
nor U1385 (N_1385,N_1281,N_1265);
nand U1386 (N_1386,N_1202,N_1268);
nor U1387 (N_1387,N_1233,N_1231);
and U1388 (N_1388,N_1222,N_1257);
and U1389 (N_1389,N_1210,N_1244);
and U1390 (N_1390,N_1200,N_1285);
and U1391 (N_1391,N_1215,N_1221);
or U1392 (N_1392,N_1254,N_1202);
nand U1393 (N_1393,N_1213,N_1271);
or U1394 (N_1394,N_1256,N_1297);
nor U1395 (N_1395,N_1243,N_1251);
nor U1396 (N_1396,N_1230,N_1229);
and U1397 (N_1397,N_1278,N_1217);
nand U1398 (N_1398,N_1221,N_1228);
xor U1399 (N_1399,N_1278,N_1205);
or U1400 (N_1400,N_1370,N_1394);
nand U1401 (N_1401,N_1380,N_1321);
nand U1402 (N_1402,N_1353,N_1342);
or U1403 (N_1403,N_1304,N_1301);
nor U1404 (N_1404,N_1373,N_1322);
nor U1405 (N_1405,N_1302,N_1311);
nand U1406 (N_1406,N_1378,N_1361);
or U1407 (N_1407,N_1379,N_1360);
xnor U1408 (N_1408,N_1317,N_1344);
and U1409 (N_1409,N_1318,N_1372);
nor U1410 (N_1410,N_1399,N_1309);
nand U1411 (N_1411,N_1312,N_1364);
nor U1412 (N_1412,N_1307,N_1326);
or U1413 (N_1413,N_1382,N_1366);
nand U1414 (N_1414,N_1349,N_1384);
nor U1415 (N_1415,N_1306,N_1357);
and U1416 (N_1416,N_1333,N_1335);
nor U1417 (N_1417,N_1354,N_1392);
nor U1418 (N_1418,N_1351,N_1397);
nor U1419 (N_1419,N_1336,N_1352);
nor U1420 (N_1420,N_1377,N_1355);
or U1421 (N_1421,N_1303,N_1369);
and U1422 (N_1422,N_1389,N_1345);
and U1423 (N_1423,N_1359,N_1362);
or U1424 (N_1424,N_1356,N_1385);
xor U1425 (N_1425,N_1327,N_1347);
nor U1426 (N_1426,N_1371,N_1319);
and U1427 (N_1427,N_1325,N_1334);
and U1428 (N_1428,N_1320,N_1396);
nand U1429 (N_1429,N_1337,N_1315);
and U1430 (N_1430,N_1365,N_1300);
nor U1431 (N_1431,N_1330,N_1340);
or U1432 (N_1432,N_1310,N_1329);
or U1433 (N_1433,N_1341,N_1367);
and U1434 (N_1434,N_1374,N_1393);
and U1435 (N_1435,N_1308,N_1358);
or U1436 (N_1436,N_1398,N_1395);
xnor U1437 (N_1437,N_1314,N_1331);
nand U1438 (N_1438,N_1387,N_1305);
or U1439 (N_1439,N_1313,N_1332);
nor U1440 (N_1440,N_1323,N_1343);
or U1441 (N_1441,N_1376,N_1338);
or U1442 (N_1442,N_1381,N_1339);
and U1443 (N_1443,N_1388,N_1348);
and U1444 (N_1444,N_1346,N_1350);
and U1445 (N_1445,N_1316,N_1328);
xor U1446 (N_1446,N_1375,N_1368);
and U1447 (N_1447,N_1363,N_1324);
or U1448 (N_1448,N_1383,N_1386);
or U1449 (N_1449,N_1391,N_1390);
nand U1450 (N_1450,N_1321,N_1337);
nor U1451 (N_1451,N_1318,N_1347);
and U1452 (N_1452,N_1357,N_1339);
nand U1453 (N_1453,N_1301,N_1371);
or U1454 (N_1454,N_1334,N_1358);
xor U1455 (N_1455,N_1371,N_1339);
and U1456 (N_1456,N_1350,N_1331);
or U1457 (N_1457,N_1312,N_1335);
nand U1458 (N_1458,N_1326,N_1387);
nor U1459 (N_1459,N_1339,N_1373);
or U1460 (N_1460,N_1301,N_1368);
and U1461 (N_1461,N_1368,N_1398);
nand U1462 (N_1462,N_1380,N_1392);
and U1463 (N_1463,N_1304,N_1370);
nor U1464 (N_1464,N_1390,N_1384);
nand U1465 (N_1465,N_1372,N_1382);
xnor U1466 (N_1466,N_1384,N_1373);
or U1467 (N_1467,N_1356,N_1380);
or U1468 (N_1468,N_1396,N_1309);
and U1469 (N_1469,N_1368,N_1386);
nor U1470 (N_1470,N_1397,N_1354);
nor U1471 (N_1471,N_1319,N_1325);
nand U1472 (N_1472,N_1375,N_1312);
nand U1473 (N_1473,N_1338,N_1334);
nand U1474 (N_1474,N_1386,N_1313);
and U1475 (N_1475,N_1326,N_1371);
and U1476 (N_1476,N_1357,N_1390);
or U1477 (N_1477,N_1364,N_1388);
and U1478 (N_1478,N_1363,N_1326);
and U1479 (N_1479,N_1322,N_1366);
nand U1480 (N_1480,N_1363,N_1399);
nand U1481 (N_1481,N_1352,N_1339);
or U1482 (N_1482,N_1354,N_1349);
or U1483 (N_1483,N_1320,N_1342);
xor U1484 (N_1484,N_1319,N_1331);
nor U1485 (N_1485,N_1377,N_1372);
or U1486 (N_1486,N_1338,N_1305);
nand U1487 (N_1487,N_1329,N_1314);
and U1488 (N_1488,N_1374,N_1300);
nand U1489 (N_1489,N_1386,N_1339);
and U1490 (N_1490,N_1392,N_1315);
and U1491 (N_1491,N_1368,N_1333);
and U1492 (N_1492,N_1325,N_1399);
nor U1493 (N_1493,N_1362,N_1355);
or U1494 (N_1494,N_1303,N_1371);
nand U1495 (N_1495,N_1355,N_1371);
xnor U1496 (N_1496,N_1391,N_1314);
nand U1497 (N_1497,N_1396,N_1385);
nand U1498 (N_1498,N_1365,N_1353);
and U1499 (N_1499,N_1360,N_1326);
nand U1500 (N_1500,N_1448,N_1403);
nand U1501 (N_1501,N_1437,N_1485);
nand U1502 (N_1502,N_1474,N_1410);
nor U1503 (N_1503,N_1496,N_1484);
or U1504 (N_1504,N_1458,N_1452);
xor U1505 (N_1505,N_1427,N_1411);
nor U1506 (N_1506,N_1473,N_1483);
nand U1507 (N_1507,N_1438,N_1447);
xor U1508 (N_1508,N_1424,N_1497);
and U1509 (N_1509,N_1444,N_1493);
and U1510 (N_1510,N_1453,N_1482);
or U1511 (N_1511,N_1480,N_1412);
and U1512 (N_1512,N_1429,N_1471);
or U1513 (N_1513,N_1460,N_1494);
and U1514 (N_1514,N_1416,N_1434);
nor U1515 (N_1515,N_1407,N_1446);
or U1516 (N_1516,N_1409,N_1408);
nand U1517 (N_1517,N_1487,N_1405);
or U1518 (N_1518,N_1454,N_1415);
nand U1519 (N_1519,N_1422,N_1441);
nand U1520 (N_1520,N_1426,N_1462);
nor U1521 (N_1521,N_1461,N_1490);
or U1522 (N_1522,N_1435,N_1449);
and U1523 (N_1523,N_1450,N_1489);
and U1524 (N_1524,N_1498,N_1423);
nor U1525 (N_1525,N_1457,N_1421);
nor U1526 (N_1526,N_1451,N_1466);
nor U1527 (N_1527,N_1430,N_1463);
nor U1528 (N_1528,N_1414,N_1445);
xnor U1529 (N_1529,N_1433,N_1400);
and U1530 (N_1530,N_1459,N_1443);
nor U1531 (N_1531,N_1425,N_1499);
nand U1532 (N_1532,N_1455,N_1468);
nor U1533 (N_1533,N_1440,N_1432);
xor U1534 (N_1534,N_1418,N_1479);
xor U1535 (N_1535,N_1488,N_1404);
and U1536 (N_1536,N_1476,N_1481);
or U1537 (N_1537,N_1428,N_1492);
nor U1538 (N_1538,N_1470,N_1456);
nand U1539 (N_1539,N_1419,N_1465);
or U1540 (N_1540,N_1401,N_1413);
nor U1541 (N_1541,N_1417,N_1491);
or U1542 (N_1542,N_1469,N_1442);
nor U1543 (N_1543,N_1475,N_1467);
and U1544 (N_1544,N_1478,N_1439);
and U1545 (N_1545,N_1472,N_1431);
nand U1546 (N_1546,N_1402,N_1464);
or U1547 (N_1547,N_1477,N_1406);
nor U1548 (N_1548,N_1486,N_1495);
nor U1549 (N_1549,N_1420,N_1436);
nand U1550 (N_1550,N_1419,N_1447);
or U1551 (N_1551,N_1415,N_1440);
nor U1552 (N_1552,N_1474,N_1446);
and U1553 (N_1553,N_1492,N_1404);
nor U1554 (N_1554,N_1469,N_1418);
nor U1555 (N_1555,N_1489,N_1453);
and U1556 (N_1556,N_1460,N_1448);
and U1557 (N_1557,N_1408,N_1462);
and U1558 (N_1558,N_1486,N_1404);
and U1559 (N_1559,N_1419,N_1494);
nand U1560 (N_1560,N_1423,N_1415);
or U1561 (N_1561,N_1421,N_1406);
and U1562 (N_1562,N_1446,N_1440);
nor U1563 (N_1563,N_1423,N_1404);
or U1564 (N_1564,N_1473,N_1460);
nand U1565 (N_1565,N_1405,N_1437);
nand U1566 (N_1566,N_1411,N_1497);
or U1567 (N_1567,N_1469,N_1459);
and U1568 (N_1568,N_1494,N_1478);
nor U1569 (N_1569,N_1455,N_1446);
and U1570 (N_1570,N_1493,N_1468);
or U1571 (N_1571,N_1472,N_1457);
nand U1572 (N_1572,N_1426,N_1463);
nor U1573 (N_1573,N_1435,N_1488);
and U1574 (N_1574,N_1457,N_1407);
nor U1575 (N_1575,N_1421,N_1412);
and U1576 (N_1576,N_1478,N_1472);
nand U1577 (N_1577,N_1403,N_1418);
xor U1578 (N_1578,N_1477,N_1473);
or U1579 (N_1579,N_1473,N_1422);
nand U1580 (N_1580,N_1432,N_1452);
and U1581 (N_1581,N_1411,N_1466);
nor U1582 (N_1582,N_1492,N_1484);
xor U1583 (N_1583,N_1454,N_1420);
or U1584 (N_1584,N_1484,N_1478);
nand U1585 (N_1585,N_1428,N_1445);
and U1586 (N_1586,N_1487,N_1456);
and U1587 (N_1587,N_1476,N_1457);
and U1588 (N_1588,N_1495,N_1472);
and U1589 (N_1589,N_1429,N_1452);
nor U1590 (N_1590,N_1446,N_1465);
and U1591 (N_1591,N_1429,N_1453);
or U1592 (N_1592,N_1464,N_1477);
and U1593 (N_1593,N_1442,N_1488);
or U1594 (N_1594,N_1401,N_1457);
or U1595 (N_1595,N_1468,N_1435);
nor U1596 (N_1596,N_1432,N_1400);
or U1597 (N_1597,N_1462,N_1400);
nor U1598 (N_1598,N_1489,N_1414);
or U1599 (N_1599,N_1463,N_1418);
nor U1600 (N_1600,N_1544,N_1596);
and U1601 (N_1601,N_1565,N_1550);
or U1602 (N_1602,N_1527,N_1514);
nand U1603 (N_1603,N_1589,N_1532);
nand U1604 (N_1604,N_1512,N_1516);
nand U1605 (N_1605,N_1554,N_1560);
or U1606 (N_1606,N_1526,N_1521);
and U1607 (N_1607,N_1592,N_1585);
and U1608 (N_1608,N_1510,N_1599);
xor U1609 (N_1609,N_1530,N_1506);
xnor U1610 (N_1610,N_1597,N_1534);
and U1611 (N_1611,N_1561,N_1549);
nor U1612 (N_1612,N_1517,N_1531);
xor U1613 (N_1613,N_1564,N_1522);
nand U1614 (N_1614,N_1518,N_1537);
nand U1615 (N_1615,N_1547,N_1573);
or U1616 (N_1616,N_1502,N_1567);
or U1617 (N_1617,N_1538,N_1587);
and U1618 (N_1618,N_1576,N_1548);
and U1619 (N_1619,N_1511,N_1507);
or U1620 (N_1620,N_1571,N_1594);
or U1621 (N_1621,N_1591,N_1568);
nor U1622 (N_1622,N_1569,N_1528);
nor U1623 (N_1623,N_1582,N_1581);
or U1624 (N_1624,N_1553,N_1543);
nand U1625 (N_1625,N_1579,N_1551);
nor U1626 (N_1626,N_1577,N_1586);
nand U1627 (N_1627,N_1513,N_1555);
or U1628 (N_1628,N_1529,N_1590);
or U1629 (N_1629,N_1520,N_1578);
and U1630 (N_1630,N_1524,N_1557);
and U1631 (N_1631,N_1535,N_1580);
and U1632 (N_1632,N_1588,N_1509);
nand U1633 (N_1633,N_1563,N_1552);
nor U1634 (N_1634,N_1542,N_1508);
xnor U1635 (N_1635,N_1546,N_1583);
and U1636 (N_1636,N_1541,N_1566);
nor U1637 (N_1637,N_1540,N_1584);
nor U1638 (N_1638,N_1505,N_1572);
and U1639 (N_1639,N_1501,N_1559);
or U1640 (N_1640,N_1558,N_1562);
nor U1641 (N_1641,N_1539,N_1556);
and U1642 (N_1642,N_1525,N_1536);
nand U1643 (N_1643,N_1545,N_1574);
nand U1644 (N_1644,N_1570,N_1575);
or U1645 (N_1645,N_1598,N_1503);
and U1646 (N_1646,N_1519,N_1593);
and U1647 (N_1647,N_1515,N_1500);
and U1648 (N_1648,N_1523,N_1504);
nand U1649 (N_1649,N_1533,N_1595);
nand U1650 (N_1650,N_1585,N_1558);
nor U1651 (N_1651,N_1565,N_1561);
and U1652 (N_1652,N_1569,N_1507);
nand U1653 (N_1653,N_1580,N_1500);
or U1654 (N_1654,N_1571,N_1550);
or U1655 (N_1655,N_1524,N_1512);
or U1656 (N_1656,N_1544,N_1573);
nand U1657 (N_1657,N_1588,N_1533);
nor U1658 (N_1658,N_1563,N_1550);
nor U1659 (N_1659,N_1540,N_1594);
nand U1660 (N_1660,N_1580,N_1562);
or U1661 (N_1661,N_1525,N_1583);
and U1662 (N_1662,N_1564,N_1537);
nand U1663 (N_1663,N_1599,N_1535);
or U1664 (N_1664,N_1572,N_1591);
or U1665 (N_1665,N_1501,N_1500);
and U1666 (N_1666,N_1597,N_1501);
or U1667 (N_1667,N_1510,N_1557);
and U1668 (N_1668,N_1584,N_1549);
and U1669 (N_1669,N_1585,N_1537);
nand U1670 (N_1670,N_1575,N_1587);
and U1671 (N_1671,N_1566,N_1536);
nand U1672 (N_1672,N_1545,N_1523);
xor U1673 (N_1673,N_1573,N_1532);
or U1674 (N_1674,N_1528,N_1562);
or U1675 (N_1675,N_1572,N_1523);
nand U1676 (N_1676,N_1549,N_1509);
or U1677 (N_1677,N_1569,N_1510);
or U1678 (N_1678,N_1583,N_1581);
nor U1679 (N_1679,N_1577,N_1563);
or U1680 (N_1680,N_1503,N_1555);
nand U1681 (N_1681,N_1555,N_1584);
and U1682 (N_1682,N_1513,N_1540);
nand U1683 (N_1683,N_1546,N_1519);
nor U1684 (N_1684,N_1593,N_1581);
nor U1685 (N_1685,N_1540,N_1553);
nor U1686 (N_1686,N_1576,N_1541);
nand U1687 (N_1687,N_1500,N_1569);
nand U1688 (N_1688,N_1549,N_1513);
nor U1689 (N_1689,N_1523,N_1528);
and U1690 (N_1690,N_1518,N_1557);
or U1691 (N_1691,N_1562,N_1541);
nand U1692 (N_1692,N_1507,N_1598);
or U1693 (N_1693,N_1593,N_1536);
nand U1694 (N_1694,N_1545,N_1543);
or U1695 (N_1695,N_1575,N_1562);
xor U1696 (N_1696,N_1513,N_1536);
and U1697 (N_1697,N_1528,N_1537);
or U1698 (N_1698,N_1529,N_1546);
or U1699 (N_1699,N_1559,N_1541);
and U1700 (N_1700,N_1616,N_1646);
nand U1701 (N_1701,N_1681,N_1603);
and U1702 (N_1702,N_1625,N_1657);
nor U1703 (N_1703,N_1649,N_1620);
and U1704 (N_1704,N_1634,N_1697);
or U1705 (N_1705,N_1654,N_1656);
and U1706 (N_1706,N_1624,N_1675);
or U1707 (N_1707,N_1651,N_1636);
or U1708 (N_1708,N_1672,N_1685);
or U1709 (N_1709,N_1638,N_1680);
xor U1710 (N_1710,N_1650,N_1668);
or U1711 (N_1711,N_1683,N_1658);
nor U1712 (N_1712,N_1660,N_1631);
and U1713 (N_1713,N_1663,N_1615);
nor U1714 (N_1714,N_1679,N_1659);
and U1715 (N_1715,N_1676,N_1623);
and U1716 (N_1716,N_1619,N_1647);
nor U1717 (N_1717,N_1629,N_1641);
nand U1718 (N_1718,N_1667,N_1653);
nand U1719 (N_1719,N_1648,N_1682);
nor U1720 (N_1720,N_1644,N_1696);
or U1721 (N_1721,N_1639,N_1677);
nor U1722 (N_1722,N_1662,N_1628);
nand U1723 (N_1723,N_1607,N_1614);
nand U1724 (N_1724,N_1602,N_1652);
xnor U1725 (N_1725,N_1608,N_1635);
or U1726 (N_1726,N_1694,N_1609);
and U1727 (N_1727,N_1626,N_1643);
or U1728 (N_1728,N_1687,N_1633);
or U1729 (N_1729,N_1673,N_1655);
or U1730 (N_1730,N_1665,N_1613);
and U1731 (N_1731,N_1671,N_1605);
or U1732 (N_1732,N_1640,N_1617);
nor U1733 (N_1733,N_1604,N_1693);
nand U1734 (N_1734,N_1611,N_1601);
and U1735 (N_1735,N_1688,N_1678);
or U1736 (N_1736,N_1692,N_1686);
nand U1737 (N_1737,N_1674,N_1690);
nand U1738 (N_1738,N_1698,N_1670);
nand U1739 (N_1739,N_1642,N_1666);
and U1740 (N_1740,N_1618,N_1627);
nor U1741 (N_1741,N_1689,N_1695);
nor U1742 (N_1742,N_1637,N_1691);
and U1743 (N_1743,N_1632,N_1621);
and U1744 (N_1744,N_1622,N_1645);
nand U1745 (N_1745,N_1612,N_1630);
nor U1746 (N_1746,N_1664,N_1684);
xor U1747 (N_1747,N_1600,N_1699);
and U1748 (N_1748,N_1610,N_1606);
and U1749 (N_1749,N_1669,N_1661);
or U1750 (N_1750,N_1669,N_1635);
nor U1751 (N_1751,N_1686,N_1616);
or U1752 (N_1752,N_1663,N_1671);
nor U1753 (N_1753,N_1645,N_1690);
nand U1754 (N_1754,N_1661,N_1636);
or U1755 (N_1755,N_1647,N_1681);
nor U1756 (N_1756,N_1692,N_1667);
nand U1757 (N_1757,N_1670,N_1607);
or U1758 (N_1758,N_1637,N_1624);
nand U1759 (N_1759,N_1601,N_1682);
nor U1760 (N_1760,N_1642,N_1669);
nand U1761 (N_1761,N_1658,N_1640);
or U1762 (N_1762,N_1677,N_1615);
and U1763 (N_1763,N_1654,N_1691);
and U1764 (N_1764,N_1662,N_1634);
or U1765 (N_1765,N_1633,N_1659);
or U1766 (N_1766,N_1652,N_1682);
or U1767 (N_1767,N_1624,N_1668);
nand U1768 (N_1768,N_1607,N_1640);
or U1769 (N_1769,N_1628,N_1699);
and U1770 (N_1770,N_1639,N_1670);
or U1771 (N_1771,N_1652,N_1662);
nor U1772 (N_1772,N_1663,N_1680);
or U1773 (N_1773,N_1670,N_1675);
nand U1774 (N_1774,N_1646,N_1668);
and U1775 (N_1775,N_1696,N_1699);
nand U1776 (N_1776,N_1646,N_1645);
and U1777 (N_1777,N_1630,N_1642);
and U1778 (N_1778,N_1674,N_1646);
or U1779 (N_1779,N_1614,N_1696);
nor U1780 (N_1780,N_1653,N_1669);
and U1781 (N_1781,N_1631,N_1652);
nor U1782 (N_1782,N_1653,N_1641);
nor U1783 (N_1783,N_1641,N_1638);
nor U1784 (N_1784,N_1629,N_1695);
and U1785 (N_1785,N_1612,N_1676);
or U1786 (N_1786,N_1623,N_1696);
and U1787 (N_1787,N_1602,N_1674);
xor U1788 (N_1788,N_1690,N_1636);
and U1789 (N_1789,N_1646,N_1613);
nor U1790 (N_1790,N_1605,N_1692);
and U1791 (N_1791,N_1618,N_1615);
and U1792 (N_1792,N_1678,N_1650);
nand U1793 (N_1793,N_1698,N_1657);
nor U1794 (N_1794,N_1670,N_1649);
nor U1795 (N_1795,N_1669,N_1643);
nor U1796 (N_1796,N_1607,N_1601);
and U1797 (N_1797,N_1658,N_1650);
xor U1798 (N_1798,N_1649,N_1622);
and U1799 (N_1799,N_1656,N_1604);
nor U1800 (N_1800,N_1796,N_1775);
or U1801 (N_1801,N_1771,N_1715);
or U1802 (N_1802,N_1763,N_1780);
nand U1803 (N_1803,N_1766,N_1779);
nor U1804 (N_1804,N_1791,N_1738);
nand U1805 (N_1805,N_1750,N_1739);
or U1806 (N_1806,N_1751,N_1765);
and U1807 (N_1807,N_1713,N_1749);
and U1808 (N_1808,N_1769,N_1770);
nor U1809 (N_1809,N_1781,N_1795);
and U1810 (N_1810,N_1708,N_1764);
nand U1811 (N_1811,N_1716,N_1797);
nor U1812 (N_1812,N_1798,N_1777);
xnor U1813 (N_1813,N_1754,N_1740);
nand U1814 (N_1814,N_1788,N_1761);
nand U1815 (N_1815,N_1755,N_1790);
nor U1816 (N_1816,N_1747,N_1792);
and U1817 (N_1817,N_1735,N_1700);
nand U1818 (N_1818,N_1701,N_1785);
nand U1819 (N_1819,N_1722,N_1772);
and U1820 (N_1820,N_1794,N_1727);
or U1821 (N_1821,N_1767,N_1752);
and U1822 (N_1822,N_1724,N_1707);
and U1823 (N_1823,N_1784,N_1718);
and U1824 (N_1824,N_1744,N_1723);
xor U1825 (N_1825,N_1732,N_1733);
or U1826 (N_1826,N_1710,N_1717);
and U1827 (N_1827,N_1737,N_1799);
or U1828 (N_1828,N_1730,N_1745);
and U1829 (N_1829,N_1725,N_1789);
and U1830 (N_1830,N_1711,N_1793);
nand U1831 (N_1831,N_1703,N_1762);
nor U1832 (N_1832,N_1776,N_1712);
or U1833 (N_1833,N_1702,N_1786);
nand U1834 (N_1834,N_1758,N_1714);
nand U1835 (N_1835,N_1736,N_1753);
nor U1836 (N_1836,N_1741,N_1782);
nand U1837 (N_1837,N_1729,N_1774);
nor U1838 (N_1838,N_1757,N_1759);
nor U1839 (N_1839,N_1768,N_1726);
or U1840 (N_1840,N_1719,N_1787);
nor U1841 (N_1841,N_1748,N_1756);
xor U1842 (N_1842,N_1760,N_1728);
nand U1843 (N_1843,N_1705,N_1743);
and U1844 (N_1844,N_1778,N_1706);
and U1845 (N_1845,N_1783,N_1773);
nand U1846 (N_1846,N_1742,N_1721);
nor U1847 (N_1847,N_1704,N_1720);
nor U1848 (N_1848,N_1731,N_1746);
and U1849 (N_1849,N_1709,N_1734);
or U1850 (N_1850,N_1768,N_1740);
or U1851 (N_1851,N_1749,N_1725);
or U1852 (N_1852,N_1783,N_1723);
nor U1853 (N_1853,N_1764,N_1773);
or U1854 (N_1854,N_1771,N_1755);
and U1855 (N_1855,N_1762,N_1713);
and U1856 (N_1856,N_1741,N_1772);
nand U1857 (N_1857,N_1705,N_1700);
and U1858 (N_1858,N_1728,N_1776);
or U1859 (N_1859,N_1705,N_1759);
nor U1860 (N_1860,N_1774,N_1731);
nand U1861 (N_1861,N_1754,N_1722);
nor U1862 (N_1862,N_1792,N_1755);
nor U1863 (N_1863,N_1784,N_1723);
nand U1864 (N_1864,N_1736,N_1791);
nor U1865 (N_1865,N_1776,N_1757);
nand U1866 (N_1866,N_1767,N_1711);
and U1867 (N_1867,N_1797,N_1790);
and U1868 (N_1868,N_1780,N_1776);
and U1869 (N_1869,N_1797,N_1735);
nor U1870 (N_1870,N_1700,N_1771);
nand U1871 (N_1871,N_1759,N_1782);
nand U1872 (N_1872,N_1746,N_1709);
nor U1873 (N_1873,N_1719,N_1751);
nor U1874 (N_1874,N_1747,N_1771);
nor U1875 (N_1875,N_1740,N_1719);
or U1876 (N_1876,N_1792,N_1795);
or U1877 (N_1877,N_1747,N_1783);
nand U1878 (N_1878,N_1757,N_1725);
nor U1879 (N_1879,N_1723,N_1737);
nand U1880 (N_1880,N_1712,N_1798);
or U1881 (N_1881,N_1762,N_1712);
nand U1882 (N_1882,N_1704,N_1726);
or U1883 (N_1883,N_1789,N_1799);
nand U1884 (N_1884,N_1769,N_1717);
nand U1885 (N_1885,N_1733,N_1729);
and U1886 (N_1886,N_1737,N_1774);
nor U1887 (N_1887,N_1739,N_1780);
nor U1888 (N_1888,N_1728,N_1744);
nand U1889 (N_1889,N_1789,N_1701);
and U1890 (N_1890,N_1733,N_1746);
nor U1891 (N_1891,N_1778,N_1725);
or U1892 (N_1892,N_1760,N_1739);
nor U1893 (N_1893,N_1711,N_1766);
and U1894 (N_1894,N_1707,N_1747);
and U1895 (N_1895,N_1782,N_1713);
nor U1896 (N_1896,N_1795,N_1703);
nand U1897 (N_1897,N_1722,N_1764);
nor U1898 (N_1898,N_1700,N_1702);
or U1899 (N_1899,N_1764,N_1721);
nand U1900 (N_1900,N_1882,N_1817);
and U1901 (N_1901,N_1870,N_1819);
or U1902 (N_1902,N_1852,N_1875);
and U1903 (N_1903,N_1814,N_1830);
nor U1904 (N_1904,N_1856,N_1897);
and U1905 (N_1905,N_1807,N_1826);
or U1906 (N_1906,N_1805,N_1858);
and U1907 (N_1907,N_1801,N_1891);
and U1908 (N_1908,N_1868,N_1827);
and U1909 (N_1909,N_1816,N_1825);
nand U1910 (N_1910,N_1836,N_1876);
nor U1911 (N_1911,N_1832,N_1899);
nor U1912 (N_1912,N_1828,N_1895);
nand U1913 (N_1913,N_1885,N_1839);
or U1914 (N_1914,N_1883,N_1874);
and U1915 (N_1915,N_1802,N_1811);
or U1916 (N_1916,N_1845,N_1887);
or U1917 (N_1917,N_1840,N_1831);
and U1918 (N_1918,N_1892,N_1808);
or U1919 (N_1919,N_1823,N_1859);
or U1920 (N_1920,N_1829,N_1851);
xnor U1921 (N_1921,N_1824,N_1857);
and U1922 (N_1922,N_1860,N_1869);
nand U1923 (N_1923,N_1820,N_1848);
nand U1924 (N_1924,N_1833,N_1893);
nand U1925 (N_1925,N_1862,N_1881);
nand U1926 (N_1926,N_1879,N_1880);
and U1927 (N_1927,N_1803,N_1873);
nand U1928 (N_1928,N_1884,N_1834);
nand U1929 (N_1929,N_1867,N_1864);
or U1930 (N_1930,N_1872,N_1898);
and U1931 (N_1931,N_1821,N_1877);
nand U1932 (N_1932,N_1854,N_1813);
nor U1933 (N_1933,N_1865,N_1837);
or U1934 (N_1934,N_1835,N_1866);
or U1935 (N_1935,N_1846,N_1855);
xnor U1936 (N_1936,N_1804,N_1809);
nor U1937 (N_1937,N_1818,N_1822);
nand U1938 (N_1938,N_1815,N_1842);
and U1939 (N_1939,N_1853,N_1838);
or U1940 (N_1940,N_1890,N_1878);
nor U1941 (N_1941,N_1894,N_1850);
xor U1942 (N_1942,N_1871,N_1888);
nand U1943 (N_1943,N_1844,N_1861);
xnor U1944 (N_1944,N_1843,N_1806);
and U1945 (N_1945,N_1849,N_1889);
and U1946 (N_1946,N_1886,N_1810);
nor U1947 (N_1947,N_1841,N_1896);
nor U1948 (N_1948,N_1800,N_1863);
nor U1949 (N_1949,N_1812,N_1847);
nor U1950 (N_1950,N_1831,N_1865);
or U1951 (N_1951,N_1810,N_1865);
and U1952 (N_1952,N_1836,N_1816);
or U1953 (N_1953,N_1875,N_1868);
nor U1954 (N_1954,N_1868,N_1858);
or U1955 (N_1955,N_1849,N_1857);
nor U1956 (N_1956,N_1870,N_1841);
nor U1957 (N_1957,N_1838,N_1837);
and U1958 (N_1958,N_1842,N_1862);
nand U1959 (N_1959,N_1837,N_1831);
and U1960 (N_1960,N_1879,N_1828);
nor U1961 (N_1961,N_1872,N_1874);
or U1962 (N_1962,N_1891,N_1892);
nor U1963 (N_1963,N_1800,N_1840);
nand U1964 (N_1964,N_1831,N_1828);
or U1965 (N_1965,N_1886,N_1833);
nor U1966 (N_1966,N_1836,N_1838);
and U1967 (N_1967,N_1811,N_1896);
nand U1968 (N_1968,N_1838,N_1885);
nor U1969 (N_1969,N_1839,N_1874);
or U1970 (N_1970,N_1800,N_1862);
and U1971 (N_1971,N_1862,N_1816);
nand U1972 (N_1972,N_1882,N_1853);
or U1973 (N_1973,N_1806,N_1809);
or U1974 (N_1974,N_1812,N_1894);
or U1975 (N_1975,N_1850,N_1837);
and U1976 (N_1976,N_1840,N_1876);
or U1977 (N_1977,N_1818,N_1815);
or U1978 (N_1978,N_1879,N_1806);
or U1979 (N_1979,N_1820,N_1840);
nor U1980 (N_1980,N_1867,N_1875);
and U1981 (N_1981,N_1818,N_1839);
and U1982 (N_1982,N_1800,N_1898);
and U1983 (N_1983,N_1828,N_1842);
and U1984 (N_1984,N_1879,N_1860);
and U1985 (N_1985,N_1886,N_1800);
and U1986 (N_1986,N_1821,N_1831);
nand U1987 (N_1987,N_1852,N_1867);
or U1988 (N_1988,N_1877,N_1864);
nor U1989 (N_1989,N_1892,N_1865);
and U1990 (N_1990,N_1867,N_1822);
and U1991 (N_1991,N_1878,N_1811);
nand U1992 (N_1992,N_1879,N_1830);
nand U1993 (N_1993,N_1834,N_1842);
nor U1994 (N_1994,N_1847,N_1885);
nand U1995 (N_1995,N_1813,N_1899);
nand U1996 (N_1996,N_1840,N_1846);
xor U1997 (N_1997,N_1838,N_1827);
xnor U1998 (N_1998,N_1800,N_1893);
nor U1999 (N_1999,N_1863,N_1827);
and U2000 (N_2000,N_1919,N_1958);
nand U2001 (N_2001,N_1941,N_1976);
nor U2002 (N_2002,N_1930,N_1921);
nor U2003 (N_2003,N_1943,N_1945);
nor U2004 (N_2004,N_1999,N_1906);
and U2005 (N_2005,N_1988,N_1974);
and U2006 (N_2006,N_1992,N_1965);
nand U2007 (N_2007,N_1951,N_1911);
and U2008 (N_2008,N_1953,N_1915);
and U2009 (N_2009,N_1980,N_1957);
or U2010 (N_2010,N_1912,N_1972);
nor U2011 (N_2011,N_1914,N_1990);
or U2012 (N_2012,N_1966,N_1998);
nand U2013 (N_2013,N_1926,N_1996);
and U2014 (N_2014,N_1969,N_1936);
nor U2015 (N_2015,N_1918,N_1993);
and U2016 (N_2016,N_1978,N_1922);
nand U2017 (N_2017,N_1916,N_1944);
or U2018 (N_2018,N_1970,N_1937);
nand U2019 (N_2019,N_1907,N_1931);
or U2020 (N_2020,N_1994,N_1977);
nor U2021 (N_2021,N_1927,N_1934);
or U2022 (N_2022,N_1960,N_1963);
nand U2023 (N_2023,N_1932,N_1955);
nor U2024 (N_2024,N_1971,N_1956);
and U2025 (N_2025,N_1905,N_1952);
or U2026 (N_2026,N_1908,N_1986);
nor U2027 (N_2027,N_1962,N_1964);
or U2028 (N_2028,N_1910,N_1920);
and U2029 (N_2029,N_1902,N_1961);
and U2030 (N_2030,N_1967,N_1950);
nor U2031 (N_2031,N_1925,N_1929);
or U2032 (N_2032,N_1987,N_1989);
and U2033 (N_2033,N_1903,N_1983);
nand U2034 (N_2034,N_1979,N_1924);
nand U2035 (N_2035,N_1968,N_1948);
or U2036 (N_2036,N_1995,N_1973);
nand U2037 (N_2037,N_1923,N_1933);
and U2038 (N_2038,N_1917,N_1909);
nor U2039 (N_2039,N_1985,N_1981);
and U2040 (N_2040,N_1901,N_1947);
nor U2041 (N_2041,N_1928,N_1913);
or U2042 (N_2042,N_1942,N_1940);
and U2043 (N_2043,N_1939,N_1904);
or U2044 (N_2044,N_1949,N_1982);
nor U2045 (N_2045,N_1975,N_1946);
nand U2046 (N_2046,N_1984,N_1991);
nand U2047 (N_2047,N_1959,N_1938);
or U2048 (N_2048,N_1954,N_1900);
or U2049 (N_2049,N_1997,N_1935);
or U2050 (N_2050,N_1984,N_1988);
nor U2051 (N_2051,N_1900,N_1987);
nand U2052 (N_2052,N_1934,N_1912);
or U2053 (N_2053,N_1955,N_1926);
nor U2054 (N_2054,N_1978,N_1939);
and U2055 (N_2055,N_1999,N_1997);
nand U2056 (N_2056,N_1975,N_1992);
and U2057 (N_2057,N_1964,N_1926);
or U2058 (N_2058,N_1975,N_1930);
nor U2059 (N_2059,N_1904,N_1923);
and U2060 (N_2060,N_1988,N_1977);
or U2061 (N_2061,N_1903,N_1904);
nand U2062 (N_2062,N_1948,N_1945);
nand U2063 (N_2063,N_1924,N_1975);
or U2064 (N_2064,N_1919,N_1978);
and U2065 (N_2065,N_1960,N_1957);
nand U2066 (N_2066,N_1996,N_1950);
nor U2067 (N_2067,N_1916,N_1910);
nand U2068 (N_2068,N_1963,N_1911);
nand U2069 (N_2069,N_1908,N_1975);
or U2070 (N_2070,N_1975,N_1915);
nor U2071 (N_2071,N_1914,N_1960);
nand U2072 (N_2072,N_1985,N_1928);
nor U2073 (N_2073,N_1987,N_1938);
or U2074 (N_2074,N_1926,N_1930);
and U2075 (N_2075,N_1944,N_1932);
nor U2076 (N_2076,N_1941,N_1986);
nand U2077 (N_2077,N_1982,N_1965);
and U2078 (N_2078,N_1985,N_1970);
nor U2079 (N_2079,N_1921,N_1986);
or U2080 (N_2080,N_1942,N_1922);
and U2081 (N_2081,N_1988,N_1986);
nor U2082 (N_2082,N_1982,N_1959);
nor U2083 (N_2083,N_1908,N_1906);
and U2084 (N_2084,N_1973,N_1925);
and U2085 (N_2085,N_1979,N_1997);
or U2086 (N_2086,N_1906,N_1939);
and U2087 (N_2087,N_1924,N_1974);
or U2088 (N_2088,N_1968,N_1933);
nor U2089 (N_2089,N_1978,N_1932);
nand U2090 (N_2090,N_1917,N_1958);
or U2091 (N_2091,N_1950,N_1909);
nand U2092 (N_2092,N_1941,N_1960);
and U2093 (N_2093,N_1961,N_1934);
nand U2094 (N_2094,N_1956,N_1900);
or U2095 (N_2095,N_1939,N_1971);
or U2096 (N_2096,N_1983,N_1986);
or U2097 (N_2097,N_1968,N_1940);
or U2098 (N_2098,N_1909,N_1921);
nor U2099 (N_2099,N_1907,N_1964);
and U2100 (N_2100,N_2058,N_2024);
and U2101 (N_2101,N_2088,N_2007);
nor U2102 (N_2102,N_2032,N_2084);
nor U2103 (N_2103,N_2054,N_2001);
nand U2104 (N_2104,N_2057,N_2051);
nor U2105 (N_2105,N_2042,N_2046);
nor U2106 (N_2106,N_2029,N_2006);
nand U2107 (N_2107,N_2022,N_2049);
and U2108 (N_2108,N_2099,N_2016);
or U2109 (N_2109,N_2033,N_2078);
or U2110 (N_2110,N_2098,N_2056);
and U2111 (N_2111,N_2060,N_2004);
or U2112 (N_2112,N_2081,N_2059);
nand U2113 (N_2113,N_2030,N_2068);
or U2114 (N_2114,N_2095,N_2025);
or U2115 (N_2115,N_2093,N_2074);
and U2116 (N_2116,N_2070,N_2066);
nand U2117 (N_2117,N_2013,N_2036);
xnor U2118 (N_2118,N_2005,N_2003);
nand U2119 (N_2119,N_2079,N_2062);
and U2120 (N_2120,N_2052,N_2034);
nand U2121 (N_2121,N_2094,N_2086);
nand U2122 (N_2122,N_2087,N_2065);
and U2123 (N_2123,N_2020,N_2077);
nand U2124 (N_2124,N_2080,N_2053);
nor U2125 (N_2125,N_2083,N_2055);
or U2126 (N_2126,N_2035,N_2072);
and U2127 (N_2127,N_2028,N_2012);
or U2128 (N_2128,N_2043,N_2031);
nand U2129 (N_2129,N_2085,N_2039);
or U2130 (N_2130,N_2082,N_2009);
and U2131 (N_2131,N_2040,N_2096);
or U2132 (N_2132,N_2075,N_2045);
or U2133 (N_2133,N_2002,N_2014);
nor U2134 (N_2134,N_2092,N_2027);
or U2135 (N_2135,N_2018,N_2008);
or U2136 (N_2136,N_2017,N_2048);
nor U2137 (N_2137,N_2061,N_2091);
nand U2138 (N_2138,N_2090,N_2050);
or U2139 (N_2139,N_2026,N_2071);
nor U2140 (N_2140,N_2011,N_2089);
or U2141 (N_2141,N_2063,N_2044);
and U2142 (N_2142,N_2021,N_2069);
and U2143 (N_2143,N_2047,N_2023);
and U2144 (N_2144,N_2076,N_2041);
nand U2145 (N_2145,N_2097,N_2000);
and U2146 (N_2146,N_2010,N_2038);
nand U2147 (N_2147,N_2067,N_2019);
nand U2148 (N_2148,N_2064,N_2073);
nor U2149 (N_2149,N_2015,N_2037);
and U2150 (N_2150,N_2018,N_2059);
or U2151 (N_2151,N_2049,N_2017);
and U2152 (N_2152,N_2082,N_2094);
or U2153 (N_2153,N_2079,N_2016);
nand U2154 (N_2154,N_2029,N_2099);
and U2155 (N_2155,N_2072,N_2013);
or U2156 (N_2156,N_2012,N_2018);
nand U2157 (N_2157,N_2033,N_2093);
nand U2158 (N_2158,N_2090,N_2073);
nor U2159 (N_2159,N_2063,N_2011);
or U2160 (N_2160,N_2002,N_2008);
nand U2161 (N_2161,N_2093,N_2061);
xor U2162 (N_2162,N_2009,N_2012);
nor U2163 (N_2163,N_2021,N_2038);
nor U2164 (N_2164,N_2050,N_2004);
and U2165 (N_2165,N_2002,N_2085);
nor U2166 (N_2166,N_2018,N_2054);
nor U2167 (N_2167,N_2093,N_2064);
nand U2168 (N_2168,N_2019,N_2078);
nand U2169 (N_2169,N_2061,N_2095);
or U2170 (N_2170,N_2077,N_2031);
or U2171 (N_2171,N_2053,N_2050);
nor U2172 (N_2172,N_2025,N_2030);
nor U2173 (N_2173,N_2055,N_2007);
or U2174 (N_2174,N_2020,N_2027);
nand U2175 (N_2175,N_2056,N_2052);
nor U2176 (N_2176,N_2080,N_2040);
nor U2177 (N_2177,N_2014,N_2065);
or U2178 (N_2178,N_2043,N_2016);
nand U2179 (N_2179,N_2041,N_2027);
nand U2180 (N_2180,N_2050,N_2013);
xor U2181 (N_2181,N_2020,N_2068);
or U2182 (N_2182,N_2006,N_2037);
and U2183 (N_2183,N_2006,N_2081);
nor U2184 (N_2184,N_2059,N_2003);
and U2185 (N_2185,N_2055,N_2085);
or U2186 (N_2186,N_2009,N_2046);
nand U2187 (N_2187,N_2078,N_2008);
and U2188 (N_2188,N_2018,N_2040);
or U2189 (N_2189,N_2037,N_2046);
nor U2190 (N_2190,N_2090,N_2057);
nand U2191 (N_2191,N_2044,N_2018);
nand U2192 (N_2192,N_2023,N_2055);
or U2193 (N_2193,N_2088,N_2041);
nand U2194 (N_2194,N_2098,N_2061);
or U2195 (N_2195,N_2053,N_2023);
nand U2196 (N_2196,N_2042,N_2025);
and U2197 (N_2197,N_2086,N_2097);
nand U2198 (N_2198,N_2071,N_2082);
or U2199 (N_2199,N_2019,N_2042);
or U2200 (N_2200,N_2121,N_2161);
nand U2201 (N_2201,N_2188,N_2194);
nor U2202 (N_2202,N_2107,N_2136);
and U2203 (N_2203,N_2189,N_2168);
or U2204 (N_2204,N_2135,N_2182);
nor U2205 (N_2205,N_2142,N_2150);
xor U2206 (N_2206,N_2124,N_2164);
and U2207 (N_2207,N_2127,N_2193);
and U2208 (N_2208,N_2122,N_2172);
nor U2209 (N_2209,N_2184,N_2113);
and U2210 (N_2210,N_2165,N_2133);
nand U2211 (N_2211,N_2171,N_2128);
nor U2212 (N_2212,N_2139,N_2178);
and U2213 (N_2213,N_2167,N_2195);
nor U2214 (N_2214,N_2112,N_2160);
or U2215 (N_2215,N_2180,N_2166);
and U2216 (N_2216,N_2163,N_2109);
nand U2217 (N_2217,N_2173,N_2162);
or U2218 (N_2218,N_2108,N_2192);
and U2219 (N_2219,N_2196,N_2151);
nor U2220 (N_2220,N_2132,N_2104);
and U2221 (N_2221,N_2197,N_2126);
or U2222 (N_2222,N_2141,N_2100);
nand U2223 (N_2223,N_2181,N_2103);
nor U2224 (N_2224,N_2138,N_2152);
nor U2225 (N_2225,N_2156,N_2147);
or U2226 (N_2226,N_2199,N_2140);
and U2227 (N_2227,N_2123,N_2191);
or U2228 (N_2228,N_2110,N_2118);
and U2229 (N_2229,N_2179,N_2105);
nor U2230 (N_2230,N_2176,N_2169);
nand U2231 (N_2231,N_2143,N_2117);
or U2232 (N_2232,N_2157,N_2198);
and U2233 (N_2233,N_2116,N_2134);
and U2234 (N_2234,N_2185,N_2129);
nand U2235 (N_2235,N_2120,N_2145);
nor U2236 (N_2236,N_2190,N_2153);
or U2237 (N_2237,N_2102,N_2170);
nor U2238 (N_2238,N_2125,N_2158);
or U2239 (N_2239,N_2114,N_2175);
xnor U2240 (N_2240,N_2174,N_2187);
and U2241 (N_2241,N_2183,N_2106);
or U2242 (N_2242,N_2146,N_2148);
nand U2243 (N_2243,N_2154,N_2177);
or U2244 (N_2244,N_2131,N_2186);
or U2245 (N_2245,N_2111,N_2130);
or U2246 (N_2246,N_2149,N_2155);
and U2247 (N_2247,N_2119,N_2101);
and U2248 (N_2248,N_2159,N_2137);
nand U2249 (N_2249,N_2144,N_2115);
or U2250 (N_2250,N_2129,N_2160);
and U2251 (N_2251,N_2116,N_2124);
nand U2252 (N_2252,N_2162,N_2161);
nor U2253 (N_2253,N_2147,N_2198);
nor U2254 (N_2254,N_2123,N_2133);
and U2255 (N_2255,N_2144,N_2104);
nor U2256 (N_2256,N_2121,N_2174);
nor U2257 (N_2257,N_2115,N_2142);
and U2258 (N_2258,N_2198,N_2171);
or U2259 (N_2259,N_2187,N_2144);
nand U2260 (N_2260,N_2124,N_2102);
nand U2261 (N_2261,N_2101,N_2112);
or U2262 (N_2262,N_2111,N_2146);
or U2263 (N_2263,N_2131,N_2133);
nor U2264 (N_2264,N_2156,N_2131);
and U2265 (N_2265,N_2104,N_2180);
xnor U2266 (N_2266,N_2156,N_2198);
nand U2267 (N_2267,N_2106,N_2169);
nand U2268 (N_2268,N_2165,N_2127);
nand U2269 (N_2269,N_2188,N_2187);
nor U2270 (N_2270,N_2143,N_2100);
or U2271 (N_2271,N_2112,N_2164);
nor U2272 (N_2272,N_2132,N_2159);
and U2273 (N_2273,N_2174,N_2178);
nand U2274 (N_2274,N_2178,N_2187);
and U2275 (N_2275,N_2159,N_2196);
and U2276 (N_2276,N_2125,N_2175);
nor U2277 (N_2277,N_2110,N_2107);
or U2278 (N_2278,N_2116,N_2194);
nor U2279 (N_2279,N_2134,N_2175);
nor U2280 (N_2280,N_2111,N_2124);
nand U2281 (N_2281,N_2155,N_2195);
or U2282 (N_2282,N_2175,N_2139);
nor U2283 (N_2283,N_2139,N_2137);
and U2284 (N_2284,N_2161,N_2191);
nand U2285 (N_2285,N_2153,N_2150);
and U2286 (N_2286,N_2133,N_2136);
nor U2287 (N_2287,N_2147,N_2111);
nand U2288 (N_2288,N_2157,N_2181);
nor U2289 (N_2289,N_2145,N_2195);
or U2290 (N_2290,N_2192,N_2170);
and U2291 (N_2291,N_2164,N_2159);
or U2292 (N_2292,N_2132,N_2174);
nor U2293 (N_2293,N_2165,N_2157);
and U2294 (N_2294,N_2160,N_2183);
or U2295 (N_2295,N_2125,N_2180);
nand U2296 (N_2296,N_2154,N_2178);
nand U2297 (N_2297,N_2118,N_2172);
and U2298 (N_2298,N_2178,N_2164);
and U2299 (N_2299,N_2132,N_2130);
nor U2300 (N_2300,N_2299,N_2219);
and U2301 (N_2301,N_2222,N_2289);
and U2302 (N_2302,N_2238,N_2239);
or U2303 (N_2303,N_2267,N_2251);
and U2304 (N_2304,N_2201,N_2210);
or U2305 (N_2305,N_2232,N_2207);
or U2306 (N_2306,N_2216,N_2298);
xor U2307 (N_2307,N_2259,N_2255);
nor U2308 (N_2308,N_2233,N_2212);
nand U2309 (N_2309,N_2221,N_2261);
and U2310 (N_2310,N_2294,N_2230);
nand U2311 (N_2311,N_2269,N_2264);
and U2312 (N_2312,N_2217,N_2228);
and U2313 (N_2313,N_2257,N_2290);
nand U2314 (N_2314,N_2260,N_2211);
or U2315 (N_2315,N_2287,N_2253);
or U2316 (N_2316,N_2248,N_2205);
and U2317 (N_2317,N_2295,N_2273);
and U2318 (N_2318,N_2213,N_2263);
nor U2319 (N_2319,N_2292,N_2277);
and U2320 (N_2320,N_2202,N_2256);
nand U2321 (N_2321,N_2225,N_2250);
and U2322 (N_2322,N_2271,N_2258);
nand U2323 (N_2323,N_2226,N_2242);
and U2324 (N_2324,N_2281,N_2284);
and U2325 (N_2325,N_2234,N_2275);
and U2326 (N_2326,N_2262,N_2272);
and U2327 (N_2327,N_2285,N_2246);
nand U2328 (N_2328,N_2245,N_2209);
nor U2329 (N_2329,N_2265,N_2231);
nor U2330 (N_2330,N_2244,N_2282);
nor U2331 (N_2331,N_2240,N_2243);
nor U2332 (N_2332,N_2279,N_2237);
and U2333 (N_2333,N_2220,N_2236);
and U2334 (N_2334,N_2278,N_2200);
xnor U2335 (N_2335,N_2204,N_2208);
and U2336 (N_2336,N_2247,N_2296);
nor U2337 (N_2337,N_2283,N_2218);
or U2338 (N_2338,N_2214,N_2270);
nand U2339 (N_2339,N_2286,N_2268);
or U2340 (N_2340,N_2276,N_2223);
nand U2341 (N_2341,N_2206,N_2252);
or U2342 (N_2342,N_2291,N_2235);
nand U2343 (N_2343,N_2215,N_2203);
and U2344 (N_2344,N_2266,N_2224);
nand U2345 (N_2345,N_2254,N_2274);
nand U2346 (N_2346,N_2288,N_2241);
or U2347 (N_2347,N_2229,N_2227);
and U2348 (N_2348,N_2293,N_2249);
nor U2349 (N_2349,N_2280,N_2297);
nand U2350 (N_2350,N_2237,N_2225);
nand U2351 (N_2351,N_2240,N_2297);
nand U2352 (N_2352,N_2270,N_2261);
nand U2353 (N_2353,N_2241,N_2275);
nor U2354 (N_2354,N_2283,N_2251);
nor U2355 (N_2355,N_2203,N_2232);
nor U2356 (N_2356,N_2255,N_2210);
nand U2357 (N_2357,N_2227,N_2252);
or U2358 (N_2358,N_2205,N_2283);
nor U2359 (N_2359,N_2209,N_2216);
and U2360 (N_2360,N_2219,N_2298);
and U2361 (N_2361,N_2202,N_2294);
and U2362 (N_2362,N_2262,N_2293);
xor U2363 (N_2363,N_2270,N_2213);
nor U2364 (N_2364,N_2279,N_2272);
nand U2365 (N_2365,N_2263,N_2203);
nor U2366 (N_2366,N_2262,N_2274);
nor U2367 (N_2367,N_2291,N_2281);
nand U2368 (N_2368,N_2212,N_2232);
nor U2369 (N_2369,N_2285,N_2240);
and U2370 (N_2370,N_2236,N_2234);
nand U2371 (N_2371,N_2245,N_2239);
and U2372 (N_2372,N_2204,N_2262);
nand U2373 (N_2373,N_2299,N_2287);
nor U2374 (N_2374,N_2273,N_2203);
nand U2375 (N_2375,N_2277,N_2255);
nand U2376 (N_2376,N_2228,N_2206);
nand U2377 (N_2377,N_2206,N_2214);
nand U2378 (N_2378,N_2274,N_2278);
and U2379 (N_2379,N_2276,N_2212);
nor U2380 (N_2380,N_2239,N_2264);
nor U2381 (N_2381,N_2254,N_2256);
or U2382 (N_2382,N_2232,N_2264);
nand U2383 (N_2383,N_2257,N_2200);
or U2384 (N_2384,N_2297,N_2239);
or U2385 (N_2385,N_2263,N_2270);
and U2386 (N_2386,N_2221,N_2256);
nor U2387 (N_2387,N_2223,N_2267);
nand U2388 (N_2388,N_2258,N_2264);
nor U2389 (N_2389,N_2200,N_2213);
nor U2390 (N_2390,N_2205,N_2265);
nor U2391 (N_2391,N_2200,N_2228);
nor U2392 (N_2392,N_2208,N_2224);
or U2393 (N_2393,N_2222,N_2217);
nor U2394 (N_2394,N_2215,N_2212);
or U2395 (N_2395,N_2235,N_2241);
nor U2396 (N_2396,N_2250,N_2267);
or U2397 (N_2397,N_2248,N_2273);
and U2398 (N_2398,N_2288,N_2227);
or U2399 (N_2399,N_2273,N_2210);
and U2400 (N_2400,N_2342,N_2300);
or U2401 (N_2401,N_2377,N_2324);
xor U2402 (N_2402,N_2304,N_2371);
nor U2403 (N_2403,N_2370,N_2332);
nor U2404 (N_2404,N_2350,N_2380);
xnor U2405 (N_2405,N_2310,N_2399);
nand U2406 (N_2406,N_2303,N_2348);
or U2407 (N_2407,N_2361,N_2356);
nand U2408 (N_2408,N_2372,N_2369);
nand U2409 (N_2409,N_2390,N_2393);
and U2410 (N_2410,N_2338,N_2365);
and U2411 (N_2411,N_2351,N_2381);
nor U2412 (N_2412,N_2373,N_2317);
nor U2413 (N_2413,N_2382,N_2345);
nor U2414 (N_2414,N_2321,N_2320);
nand U2415 (N_2415,N_2314,N_2398);
and U2416 (N_2416,N_2397,N_2347);
nand U2417 (N_2417,N_2319,N_2343);
nand U2418 (N_2418,N_2341,N_2383);
nor U2419 (N_2419,N_2374,N_2305);
nor U2420 (N_2420,N_2353,N_2302);
nor U2421 (N_2421,N_2379,N_2316);
or U2422 (N_2422,N_2311,N_2395);
nor U2423 (N_2423,N_2375,N_2359);
or U2424 (N_2424,N_2307,N_2354);
or U2425 (N_2425,N_2312,N_2362);
nor U2426 (N_2426,N_2318,N_2309);
nand U2427 (N_2427,N_2308,N_2364);
or U2428 (N_2428,N_2325,N_2367);
nor U2429 (N_2429,N_2330,N_2394);
nand U2430 (N_2430,N_2355,N_2386);
and U2431 (N_2431,N_2328,N_2327);
or U2432 (N_2432,N_2385,N_2336);
nand U2433 (N_2433,N_2352,N_2323);
nor U2434 (N_2434,N_2389,N_2363);
nor U2435 (N_2435,N_2376,N_2360);
nand U2436 (N_2436,N_2340,N_2358);
and U2437 (N_2437,N_2301,N_2391);
or U2438 (N_2438,N_2326,N_2396);
nand U2439 (N_2439,N_2331,N_2392);
or U2440 (N_2440,N_2366,N_2334);
or U2441 (N_2441,N_2335,N_2322);
nor U2442 (N_2442,N_2306,N_2378);
xor U2443 (N_2443,N_2329,N_2313);
and U2444 (N_2444,N_2388,N_2349);
nor U2445 (N_2445,N_2339,N_2384);
nor U2446 (N_2446,N_2337,N_2387);
or U2447 (N_2447,N_2315,N_2368);
nand U2448 (N_2448,N_2344,N_2346);
or U2449 (N_2449,N_2333,N_2357);
nand U2450 (N_2450,N_2316,N_2354);
and U2451 (N_2451,N_2320,N_2328);
nand U2452 (N_2452,N_2321,N_2396);
or U2453 (N_2453,N_2308,N_2397);
nand U2454 (N_2454,N_2381,N_2316);
nor U2455 (N_2455,N_2379,N_2330);
nand U2456 (N_2456,N_2312,N_2329);
nor U2457 (N_2457,N_2304,N_2395);
nor U2458 (N_2458,N_2310,N_2391);
or U2459 (N_2459,N_2300,N_2329);
and U2460 (N_2460,N_2331,N_2369);
and U2461 (N_2461,N_2387,N_2384);
nor U2462 (N_2462,N_2357,N_2343);
nor U2463 (N_2463,N_2346,N_2361);
nand U2464 (N_2464,N_2340,N_2327);
nand U2465 (N_2465,N_2365,N_2360);
or U2466 (N_2466,N_2333,N_2359);
xor U2467 (N_2467,N_2361,N_2379);
nor U2468 (N_2468,N_2321,N_2387);
and U2469 (N_2469,N_2304,N_2340);
nand U2470 (N_2470,N_2362,N_2318);
or U2471 (N_2471,N_2381,N_2333);
nand U2472 (N_2472,N_2377,N_2351);
nor U2473 (N_2473,N_2324,N_2387);
or U2474 (N_2474,N_2371,N_2311);
nor U2475 (N_2475,N_2365,N_2381);
nand U2476 (N_2476,N_2358,N_2365);
and U2477 (N_2477,N_2317,N_2352);
nand U2478 (N_2478,N_2390,N_2322);
nand U2479 (N_2479,N_2304,N_2302);
nand U2480 (N_2480,N_2319,N_2373);
nand U2481 (N_2481,N_2320,N_2345);
nand U2482 (N_2482,N_2369,N_2354);
and U2483 (N_2483,N_2391,N_2304);
nand U2484 (N_2484,N_2397,N_2349);
and U2485 (N_2485,N_2369,N_2382);
and U2486 (N_2486,N_2387,N_2375);
or U2487 (N_2487,N_2328,N_2337);
and U2488 (N_2488,N_2339,N_2362);
nand U2489 (N_2489,N_2399,N_2309);
xnor U2490 (N_2490,N_2379,N_2348);
xor U2491 (N_2491,N_2355,N_2317);
or U2492 (N_2492,N_2351,N_2320);
and U2493 (N_2493,N_2377,N_2325);
or U2494 (N_2494,N_2339,N_2320);
nand U2495 (N_2495,N_2347,N_2333);
nor U2496 (N_2496,N_2369,N_2368);
nor U2497 (N_2497,N_2358,N_2317);
or U2498 (N_2498,N_2318,N_2324);
and U2499 (N_2499,N_2397,N_2329);
or U2500 (N_2500,N_2483,N_2444);
and U2501 (N_2501,N_2476,N_2497);
nor U2502 (N_2502,N_2450,N_2431);
or U2503 (N_2503,N_2409,N_2470);
or U2504 (N_2504,N_2477,N_2414);
nor U2505 (N_2505,N_2469,N_2462);
or U2506 (N_2506,N_2495,N_2482);
nand U2507 (N_2507,N_2423,N_2425);
nor U2508 (N_2508,N_2465,N_2438);
nand U2509 (N_2509,N_2479,N_2400);
or U2510 (N_2510,N_2481,N_2485);
and U2511 (N_2511,N_2448,N_2416);
nor U2512 (N_2512,N_2418,N_2430);
nand U2513 (N_2513,N_2486,N_2466);
nor U2514 (N_2514,N_2421,N_2492);
and U2515 (N_2515,N_2432,N_2426);
or U2516 (N_2516,N_2403,N_2467);
nor U2517 (N_2517,N_2422,N_2457);
nand U2518 (N_2518,N_2474,N_2419);
or U2519 (N_2519,N_2491,N_2455);
or U2520 (N_2520,N_2412,N_2446);
nor U2521 (N_2521,N_2440,N_2460);
or U2522 (N_2522,N_2480,N_2461);
nor U2523 (N_2523,N_2445,N_2439);
nand U2524 (N_2524,N_2402,N_2452);
and U2525 (N_2525,N_2442,N_2493);
nor U2526 (N_2526,N_2428,N_2443);
or U2527 (N_2527,N_2463,N_2484);
or U2528 (N_2528,N_2478,N_2475);
or U2529 (N_2529,N_2454,N_2449);
and U2530 (N_2530,N_2489,N_2464);
or U2531 (N_2531,N_2406,N_2401);
xnor U2532 (N_2532,N_2415,N_2499);
nand U2533 (N_2533,N_2427,N_2411);
xnor U2534 (N_2534,N_2413,N_2408);
nor U2535 (N_2535,N_2451,N_2410);
and U2536 (N_2536,N_2472,N_2434);
and U2537 (N_2537,N_2459,N_2404);
nand U2538 (N_2538,N_2498,N_2433);
and U2539 (N_2539,N_2490,N_2429);
nand U2540 (N_2540,N_2494,N_2496);
nand U2541 (N_2541,N_2468,N_2488);
and U2542 (N_2542,N_2458,N_2407);
and U2543 (N_2543,N_2447,N_2473);
nor U2544 (N_2544,N_2471,N_2435);
nor U2545 (N_2545,N_2441,N_2453);
and U2546 (N_2546,N_2405,N_2420);
xor U2547 (N_2547,N_2487,N_2456);
or U2548 (N_2548,N_2424,N_2437);
nor U2549 (N_2549,N_2417,N_2436);
or U2550 (N_2550,N_2429,N_2487);
xnor U2551 (N_2551,N_2432,N_2486);
nand U2552 (N_2552,N_2496,N_2402);
or U2553 (N_2553,N_2481,N_2461);
and U2554 (N_2554,N_2442,N_2482);
and U2555 (N_2555,N_2403,N_2465);
nand U2556 (N_2556,N_2400,N_2430);
or U2557 (N_2557,N_2441,N_2498);
and U2558 (N_2558,N_2473,N_2402);
and U2559 (N_2559,N_2422,N_2499);
and U2560 (N_2560,N_2436,N_2428);
or U2561 (N_2561,N_2413,N_2456);
nor U2562 (N_2562,N_2491,N_2428);
nor U2563 (N_2563,N_2468,N_2440);
nand U2564 (N_2564,N_2418,N_2474);
or U2565 (N_2565,N_2487,N_2410);
and U2566 (N_2566,N_2400,N_2426);
nand U2567 (N_2567,N_2437,N_2489);
nand U2568 (N_2568,N_2430,N_2480);
and U2569 (N_2569,N_2438,N_2430);
nand U2570 (N_2570,N_2415,N_2479);
nand U2571 (N_2571,N_2499,N_2475);
or U2572 (N_2572,N_2472,N_2448);
and U2573 (N_2573,N_2450,N_2425);
or U2574 (N_2574,N_2470,N_2450);
and U2575 (N_2575,N_2450,N_2411);
and U2576 (N_2576,N_2474,N_2433);
nand U2577 (N_2577,N_2406,N_2477);
and U2578 (N_2578,N_2472,N_2423);
and U2579 (N_2579,N_2431,N_2423);
nor U2580 (N_2580,N_2469,N_2415);
nor U2581 (N_2581,N_2499,N_2496);
or U2582 (N_2582,N_2460,N_2426);
nand U2583 (N_2583,N_2475,N_2490);
and U2584 (N_2584,N_2479,N_2410);
nand U2585 (N_2585,N_2401,N_2400);
nand U2586 (N_2586,N_2444,N_2488);
and U2587 (N_2587,N_2433,N_2488);
nand U2588 (N_2588,N_2479,N_2447);
nand U2589 (N_2589,N_2426,N_2434);
nor U2590 (N_2590,N_2461,N_2497);
or U2591 (N_2591,N_2411,N_2484);
and U2592 (N_2592,N_2465,N_2497);
or U2593 (N_2593,N_2484,N_2430);
nand U2594 (N_2594,N_2414,N_2480);
or U2595 (N_2595,N_2445,N_2484);
or U2596 (N_2596,N_2491,N_2473);
nor U2597 (N_2597,N_2443,N_2497);
nand U2598 (N_2598,N_2417,N_2458);
and U2599 (N_2599,N_2483,N_2493);
and U2600 (N_2600,N_2520,N_2539);
nor U2601 (N_2601,N_2558,N_2513);
and U2602 (N_2602,N_2588,N_2505);
or U2603 (N_2603,N_2529,N_2582);
nor U2604 (N_2604,N_2564,N_2543);
and U2605 (N_2605,N_2548,N_2569);
nand U2606 (N_2606,N_2554,N_2518);
and U2607 (N_2607,N_2589,N_2523);
nor U2608 (N_2608,N_2590,N_2593);
and U2609 (N_2609,N_2591,N_2573);
or U2610 (N_2610,N_2521,N_2598);
nor U2611 (N_2611,N_2572,N_2580);
and U2612 (N_2612,N_2549,N_2544);
or U2613 (N_2613,N_2501,N_2510);
nand U2614 (N_2614,N_2537,N_2579);
and U2615 (N_2615,N_2528,N_2542);
nor U2616 (N_2616,N_2547,N_2565);
or U2617 (N_2617,N_2538,N_2571);
or U2618 (N_2618,N_2545,N_2534);
and U2619 (N_2619,N_2568,N_2541);
and U2620 (N_2620,N_2522,N_2524);
or U2621 (N_2621,N_2532,N_2578);
nand U2622 (N_2622,N_2574,N_2540);
nand U2623 (N_2623,N_2566,N_2546);
xnor U2624 (N_2624,N_2507,N_2504);
nor U2625 (N_2625,N_2581,N_2506);
or U2626 (N_2626,N_2515,N_2527);
nand U2627 (N_2627,N_2557,N_2530);
xor U2628 (N_2628,N_2595,N_2587);
or U2629 (N_2629,N_2551,N_2511);
nor U2630 (N_2630,N_2519,N_2550);
nand U2631 (N_2631,N_2585,N_2500);
and U2632 (N_2632,N_2576,N_2526);
nor U2633 (N_2633,N_2503,N_2525);
nand U2634 (N_2634,N_2594,N_2556);
nand U2635 (N_2635,N_2559,N_2517);
or U2636 (N_2636,N_2583,N_2555);
and U2637 (N_2637,N_2570,N_2592);
or U2638 (N_2638,N_2516,N_2508);
nor U2639 (N_2639,N_2514,N_2563);
and U2640 (N_2640,N_2575,N_2553);
and U2641 (N_2641,N_2509,N_2562);
and U2642 (N_2642,N_2531,N_2577);
or U2643 (N_2643,N_2533,N_2560);
nor U2644 (N_2644,N_2561,N_2536);
nor U2645 (N_2645,N_2584,N_2599);
nand U2646 (N_2646,N_2502,N_2535);
nand U2647 (N_2647,N_2597,N_2596);
nor U2648 (N_2648,N_2586,N_2512);
and U2649 (N_2649,N_2552,N_2567);
nor U2650 (N_2650,N_2517,N_2516);
or U2651 (N_2651,N_2523,N_2505);
nand U2652 (N_2652,N_2563,N_2585);
nand U2653 (N_2653,N_2509,N_2525);
nand U2654 (N_2654,N_2515,N_2581);
and U2655 (N_2655,N_2514,N_2512);
nand U2656 (N_2656,N_2567,N_2509);
or U2657 (N_2657,N_2590,N_2563);
or U2658 (N_2658,N_2513,N_2504);
or U2659 (N_2659,N_2589,N_2583);
nor U2660 (N_2660,N_2567,N_2514);
nor U2661 (N_2661,N_2589,N_2510);
and U2662 (N_2662,N_2545,N_2569);
and U2663 (N_2663,N_2554,N_2571);
nand U2664 (N_2664,N_2572,N_2585);
and U2665 (N_2665,N_2592,N_2534);
or U2666 (N_2666,N_2520,N_2518);
nor U2667 (N_2667,N_2594,N_2543);
nand U2668 (N_2668,N_2542,N_2561);
nand U2669 (N_2669,N_2583,N_2525);
nand U2670 (N_2670,N_2509,N_2515);
or U2671 (N_2671,N_2563,N_2523);
or U2672 (N_2672,N_2584,N_2553);
or U2673 (N_2673,N_2545,N_2598);
nand U2674 (N_2674,N_2585,N_2578);
or U2675 (N_2675,N_2537,N_2503);
and U2676 (N_2676,N_2500,N_2567);
nand U2677 (N_2677,N_2531,N_2551);
and U2678 (N_2678,N_2566,N_2596);
or U2679 (N_2679,N_2589,N_2537);
nor U2680 (N_2680,N_2594,N_2502);
or U2681 (N_2681,N_2512,N_2505);
and U2682 (N_2682,N_2547,N_2556);
and U2683 (N_2683,N_2571,N_2596);
nand U2684 (N_2684,N_2532,N_2550);
xor U2685 (N_2685,N_2575,N_2501);
nor U2686 (N_2686,N_2584,N_2549);
xnor U2687 (N_2687,N_2551,N_2507);
nand U2688 (N_2688,N_2562,N_2556);
nor U2689 (N_2689,N_2571,N_2599);
and U2690 (N_2690,N_2520,N_2551);
nand U2691 (N_2691,N_2563,N_2522);
or U2692 (N_2692,N_2569,N_2582);
nand U2693 (N_2693,N_2572,N_2582);
nand U2694 (N_2694,N_2515,N_2543);
nor U2695 (N_2695,N_2503,N_2574);
nor U2696 (N_2696,N_2508,N_2509);
nand U2697 (N_2697,N_2576,N_2578);
or U2698 (N_2698,N_2559,N_2529);
nand U2699 (N_2699,N_2564,N_2549);
or U2700 (N_2700,N_2647,N_2681);
nor U2701 (N_2701,N_2642,N_2661);
and U2702 (N_2702,N_2627,N_2674);
nor U2703 (N_2703,N_2600,N_2630);
or U2704 (N_2704,N_2695,N_2654);
or U2705 (N_2705,N_2698,N_2628);
nand U2706 (N_2706,N_2685,N_2631);
or U2707 (N_2707,N_2646,N_2610);
nor U2708 (N_2708,N_2617,N_2684);
nor U2709 (N_2709,N_2613,N_2633);
and U2710 (N_2710,N_2687,N_2608);
or U2711 (N_2711,N_2667,N_2686);
or U2712 (N_2712,N_2620,N_2621);
nor U2713 (N_2713,N_2657,N_2699);
nor U2714 (N_2714,N_2672,N_2673);
or U2715 (N_2715,N_2625,N_2644);
and U2716 (N_2716,N_2622,N_2659);
and U2717 (N_2717,N_2609,N_2656);
nand U2718 (N_2718,N_2648,N_2639);
and U2719 (N_2719,N_2612,N_2655);
or U2720 (N_2720,N_2670,N_2663);
or U2721 (N_2721,N_2650,N_2679);
nor U2722 (N_2722,N_2669,N_2696);
nand U2723 (N_2723,N_2693,N_2616);
nand U2724 (N_2724,N_2615,N_2626);
and U2725 (N_2725,N_2602,N_2692);
or U2726 (N_2726,N_2607,N_2682);
nor U2727 (N_2727,N_2651,N_2605);
and U2728 (N_2728,N_2629,N_2688);
or U2729 (N_2729,N_2694,N_2678);
nand U2730 (N_2730,N_2652,N_2603);
or U2731 (N_2731,N_2689,N_2604);
and U2732 (N_2732,N_2635,N_2614);
and U2733 (N_2733,N_2606,N_2691);
nor U2734 (N_2734,N_2637,N_2690);
nor U2735 (N_2735,N_2664,N_2666);
or U2736 (N_2736,N_2640,N_2643);
or U2737 (N_2737,N_2618,N_2671);
and U2738 (N_2738,N_2601,N_2619);
nor U2739 (N_2739,N_2680,N_2675);
nor U2740 (N_2740,N_2677,N_2636);
nand U2741 (N_2741,N_2649,N_2645);
xnor U2742 (N_2742,N_2638,N_2624);
xor U2743 (N_2743,N_2623,N_2653);
nand U2744 (N_2744,N_2662,N_2665);
and U2745 (N_2745,N_2660,N_2697);
or U2746 (N_2746,N_2658,N_2641);
or U2747 (N_2747,N_2634,N_2632);
and U2748 (N_2748,N_2676,N_2668);
or U2749 (N_2749,N_2683,N_2611);
nand U2750 (N_2750,N_2672,N_2675);
or U2751 (N_2751,N_2602,N_2690);
nand U2752 (N_2752,N_2674,N_2606);
and U2753 (N_2753,N_2692,N_2632);
and U2754 (N_2754,N_2666,N_2616);
or U2755 (N_2755,N_2695,N_2638);
xor U2756 (N_2756,N_2697,N_2608);
nand U2757 (N_2757,N_2690,N_2643);
nand U2758 (N_2758,N_2632,N_2660);
nand U2759 (N_2759,N_2645,N_2634);
or U2760 (N_2760,N_2615,N_2611);
xor U2761 (N_2761,N_2687,N_2694);
nand U2762 (N_2762,N_2634,N_2693);
xnor U2763 (N_2763,N_2634,N_2624);
nand U2764 (N_2764,N_2666,N_2601);
or U2765 (N_2765,N_2657,N_2677);
nor U2766 (N_2766,N_2644,N_2646);
nor U2767 (N_2767,N_2628,N_2694);
nor U2768 (N_2768,N_2629,N_2694);
nor U2769 (N_2769,N_2600,N_2693);
and U2770 (N_2770,N_2690,N_2681);
nand U2771 (N_2771,N_2679,N_2621);
nor U2772 (N_2772,N_2648,N_2625);
nor U2773 (N_2773,N_2689,N_2656);
nand U2774 (N_2774,N_2629,N_2699);
nor U2775 (N_2775,N_2691,N_2659);
nand U2776 (N_2776,N_2699,N_2625);
nor U2777 (N_2777,N_2627,N_2621);
nand U2778 (N_2778,N_2690,N_2644);
nor U2779 (N_2779,N_2632,N_2672);
nor U2780 (N_2780,N_2664,N_2601);
nor U2781 (N_2781,N_2660,N_2651);
xor U2782 (N_2782,N_2622,N_2625);
nor U2783 (N_2783,N_2653,N_2647);
nor U2784 (N_2784,N_2695,N_2600);
nand U2785 (N_2785,N_2620,N_2632);
nor U2786 (N_2786,N_2625,N_2676);
and U2787 (N_2787,N_2604,N_2602);
and U2788 (N_2788,N_2644,N_2654);
or U2789 (N_2789,N_2672,N_2656);
nor U2790 (N_2790,N_2638,N_2660);
nor U2791 (N_2791,N_2665,N_2688);
nor U2792 (N_2792,N_2623,N_2670);
and U2793 (N_2793,N_2643,N_2672);
or U2794 (N_2794,N_2675,N_2697);
nor U2795 (N_2795,N_2672,N_2693);
nor U2796 (N_2796,N_2611,N_2696);
and U2797 (N_2797,N_2632,N_2655);
nand U2798 (N_2798,N_2696,N_2646);
and U2799 (N_2799,N_2663,N_2616);
nor U2800 (N_2800,N_2703,N_2744);
nand U2801 (N_2801,N_2728,N_2787);
nor U2802 (N_2802,N_2705,N_2711);
nor U2803 (N_2803,N_2791,N_2790);
and U2804 (N_2804,N_2724,N_2739);
nor U2805 (N_2805,N_2707,N_2710);
nand U2806 (N_2806,N_2749,N_2795);
or U2807 (N_2807,N_2723,N_2733);
and U2808 (N_2808,N_2721,N_2784);
and U2809 (N_2809,N_2709,N_2731);
and U2810 (N_2810,N_2727,N_2768);
nor U2811 (N_2811,N_2777,N_2746);
nand U2812 (N_2812,N_2718,N_2798);
and U2813 (N_2813,N_2756,N_2748);
nand U2814 (N_2814,N_2747,N_2719);
or U2815 (N_2815,N_2704,N_2759);
or U2816 (N_2816,N_2706,N_2708);
xnor U2817 (N_2817,N_2794,N_2714);
nor U2818 (N_2818,N_2765,N_2781);
nor U2819 (N_2819,N_2751,N_2778);
and U2820 (N_2820,N_2782,N_2775);
or U2821 (N_2821,N_2793,N_2783);
or U2822 (N_2822,N_2729,N_2773);
or U2823 (N_2823,N_2761,N_2702);
and U2824 (N_2824,N_2713,N_2779);
or U2825 (N_2825,N_2750,N_2742);
and U2826 (N_2826,N_2796,N_2754);
and U2827 (N_2827,N_2722,N_2720);
or U2828 (N_2828,N_2752,N_2738);
or U2829 (N_2829,N_2730,N_2717);
nand U2830 (N_2830,N_2762,N_2772);
nor U2831 (N_2831,N_2786,N_2701);
or U2832 (N_2832,N_2757,N_2741);
nand U2833 (N_2833,N_2774,N_2771);
xor U2834 (N_2834,N_2769,N_2789);
or U2835 (N_2835,N_2732,N_2737);
nand U2836 (N_2836,N_2726,N_2760);
or U2837 (N_2837,N_2797,N_2788);
nand U2838 (N_2838,N_2776,N_2715);
or U2839 (N_2839,N_2766,N_2716);
nor U2840 (N_2840,N_2770,N_2735);
or U2841 (N_2841,N_2745,N_2753);
or U2842 (N_2842,N_2740,N_2725);
nand U2843 (N_2843,N_2755,N_2743);
or U2844 (N_2844,N_2763,N_2764);
nand U2845 (N_2845,N_2799,N_2736);
and U2846 (N_2846,N_2767,N_2700);
or U2847 (N_2847,N_2785,N_2712);
and U2848 (N_2848,N_2758,N_2792);
and U2849 (N_2849,N_2734,N_2780);
and U2850 (N_2850,N_2766,N_2775);
and U2851 (N_2851,N_2700,N_2783);
nor U2852 (N_2852,N_2783,N_2799);
nand U2853 (N_2853,N_2792,N_2702);
nor U2854 (N_2854,N_2792,N_2770);
or U2855 (N_2855,N_2729,N_2730);
nand U2856 (N_2856,N_2729,N_2784);
nor U2857 (N_2857,N_2713,N_2789);
or U2858 (N_2858,N_2730,N_2739);
nand U2859 (N_2859,N_2789,N_2732);
nor U2860 (N_2860,N_2745,N_2783);
nor U2861 (N_2861,N_2756,N_2743);
or U2862 (N_2862,N_2725,N_2776);
or U2863 (N_2863,N_2727,N_2792);
and U2864 (N_2864,N_2775,N_2767);
or U2865 (N_2865,N_2769,N_2779);
or U2866 (N_2866,N_2790,N_2797);
and U2867 (N_2867,N_2787,N_2720);
nand U2868 (N_2868,N_2726,N_2778);
nor U2869 (N_2869,N_2709,N_2720);
or U2870 (N_2870,N_2729,N_2725);
or U2871 (N_2871,N_2731,N_2786);
and U2872 (N_2872,N_2710,N_2772);
and U2873 (N_2873,N_2743,N_2784);
and U2874 (N_2874,N_2733,N_2762);
nor U2875 (N_2875,N_2765,N_2707);
nor U2876 (N_2876,N_2720,N_2753);
or U2877 (N_2877,N_2797,N_2779);
nor U2878 (N_2878,N_2749,N_2796);
or U2879 (N_2879,N_2731,N_2764);
or U2880 (N_2880,N_2780,N_2754);
and U2881 (N_2881,N_2750,N_2712);
nor U2882 (N_2882,N_2744,N_2755);
nor U2883 (N_2883,N_2748,N_2765);
nor U2884 (N_2884,N_2783,N_2767);
and U2885 (N_2885,N_2757,N_2781);
nor U2886 (N_2886,N_2731,N_2742);
or U2887 (N_2887,N_2752,N_2746);
nor U2888 (N_2888,N_2772,N_2795);
nor U2889 (N_2889,N_2737,N_2730);
or U2890 (N_2890,N_2772,N_2754);
nor U2891 (N_2891,N_2717,N_2714);
and U2892 (N_2892,N_2707,N_2751);
or U2893 (N_2893,N_2778,N_2707);
or U2894 (N_2894,N_2777,N_2740);
nand U2895 (N_2895,N_2772,N_2748);
or U2896 (N_2896,N_2743,N_2747);
nand U2897 (N_2897,N_2725,N_2787);
or U2898 (N_2898,N_2787,N_2785);
or U2899 (N_2899,N_2735,N_2761);
nand U2900 (N_2900,N_2856,N_2816);
nand U2901 (N_2901,N_2837,N_2862);
and U2902 (N_2902,N_2885,N_2899);
and U2903 (N_2903,N_2882,N_2825);
and U2904 (N_2904,N_2845,N_2841);
nand U2905 (N_2905,N_2817,N_2807);
or U2906 (N_2906,N_2839,N_2827);
or U2907 (N_2907,N_2851,N_2811);
nor U2908 (N_2908,N_2838,N_2879);
and U2909 (N_2909,N_2888,N_2855);
nor U2910 (N_2910,N_2819,N_2868);
nand U2911 (N_2911,N_2832,N_2896);
nor U2912 (N_2912,N_2874,N_2818);
nand U2913 (N_2913,N_2828,N_2835);
nand U2914 (N_2914,N_2860,N_2826);
nand U2915 (N_2915,N_2808,N_2800);
and U2916 (N_2916,N_2806,N_2842);
nor U2917 (N_2917,N_2865,N_2840);
and U2918 (N_2918,N_2857,N_2802);
nor U2919 (N_2919,N_2813,N_2804);
or U2920 (N_2920,N_2815,N_2872);
nor U2921 (N_2921,N_2847,N_2834);
nor U2922 (N_2922,N_2854,N_2869);
nor U2923 (N_2923,N_2891,N_2880);
or U2924 (N_2924,N_2803,N_2820);
nor U2925 (N_2925,N_2805,N_2853);
and U2926 (N_2926,N_2846,N_2873);
and U2927 (N_2927,N_2875,N_2887);
nor U2928 (N_2928,N_2889,N_2894);
nor U2929 (N_2929,N_2881,N_2823);
or U2930 (N_2930,N_2878,N_2850);
nor U2931 (N_2931,N_2890,N_2836);
and U2932 (N_2932,N_2843,N_2892);
nor U2933 (N_2933,N_2895,N_2876);
nand U2934 (N_2934,N_2814,N_2884);
xor U2935 (N_2935,N_2822,N_2859);
nand U2936 (N_2936,N_2809,N_2877);
or U2937 (N_2937,N_2866,N_2870);
or U2938 (N_2938,N_2833,N_2858);
or U2939 (N_2939,N_2829,N_2848);
or U2940 (N_2940,N_2863,N_2824);
or U2941 (N_2941,N_2844,N_2830);
nand U2942 (N_2942,N_2852,N_2871);
and U2943 (N_2943,N_2810,N_2849);
nand U2944 (N_2944,N_2861,N_2898);
nand U2945 (N_2945,N_2893,N_2812);
or U2946 (N_2946,N_2831,N_2897);
or U2947 (N_2947,N_2801,N_2883);
nand U2948 (N_2948,N_2886,N_2867);
and U2949 (N_2949,N_2864,N_2821);
and U2950 (N_2950,N_2809,N_2813);
and U2951 (N_2951,N_2882,N_2890);
and U2952 (N_2952,N_2829,N_2883);
nor U2953 (N_2953,N_2816,N_2820);
and U2954 (N_2954,N_2892,N_2837);
nor U2955 (N_2955,N_2830,N_2821);
nor U2956 (N_2956,N_2895,N_2860);
nor U2957 (N_2957,N_2800,N_2827);
and U2958 (N_2958,N_2800,N_2833);
and U2959 (N_2959,N_2817,N_2875);
or U2960 (N_2960,N_2838,N_2804);
or U2961 (N_2961,N_2847,N_2856);
nand U2962 (N_2962,N_2827,N_2886);
and U2963 (N_2963,N_2859,N_2841);
and U2964 (N_2964,N_2827,N_2890);
xnor U2965 (N_2965,N_2841,N_2815);
nor U2966 (N_2966,N_2800,N_2822);
nand U2967 (N_2967,N_2816,N_2888);
nand U2968 (N_2968,N_2802,N_2826);
or U2969 (N_2969,N_2841,N_2824);
nor U2970 (N_2970,N_2882,N_2879);
or U2971 (N_2971,N_2838,N_2836);
nor U2972 (N_2972,N_2842,N_2819);
nor U2973 (N_2973,N_2873,N_2864);
or U2974 (N_2974,N_2832,N_2895);
and U2975 (N_2975,N_2848,N_2889);
and U2976 (N_2976,N_2897,N_2869);
nor U2977 (N_2977,N_2855,N_2823);
nand U2978 (N_2978,N_2819,N_2880);
nand U2979 (N_2979,N_2804,N_2808);
nand U2980 (N_2980,N_2824,N_2870);
nand U2981 (N_2981,N_2813,N_2862);
nor U2982 (N_2982,N_2818,N_2830);
and U2983 (N_2983,N_2814,N_2820);
nor U2984 (N_2984,N_2854,N_2803);
nand U2985 (N_2985,N_2808,N_2836);
and U2986 (N_2986,N_2833,N_2839);
or U2987 (N_2987,N_2853,N_2897);
or U2988 (N_2988,N_2879,N_2812);
or U2989 (N_2989,N_2886,N_2850);
and U2990 (N_2990,N_2870,N_2872);
xor U2991 (N_2991,N_2864,N_2809);
nand U2992 (N_2992,N_2813,N_2895);
nand U2993 (N_2993,N_2873,N_2862);
nand U2994 (N_2994,N_2833,N_2813);
and U2995 (N_2995,N_2825,N_2808);
nor U2996 (N_2996,N_2815,N_2800);
nor U2997 (N_2997,N_2868,N_2865);
nand U2998 (N_2998,N_2895,N_2872);
nor U2999 (N_2999,N_2813,N_2818);
or UO_0 (O_0,N_2930,N_2989);
and UO_1 (O_1,N_2957,N_2909);
nand UO_2 (O_2,N_2984,N_2900);
nor UO_3 (O_3,N_2991,N_2977);
or UO_4 (O_4,N_2958,N_2922);
or UO_5 (O_5,N_2965,N_2905);
nand UO_6 (O_6,N_2968,N_2927);
or UO_7 (O_7,N_2911,N_2975);
nand UO_8 (O_8,N_2962,N_2960);
nor UO_9 (O_9,N_2908,N_2994);
and UO_10 (O_10,N_2997,N_2938);
and UO_11 (O_11,N_2929,N_2954);
or UO_12 (O_12,N_2952,N_2933);
nand UO_13 (O_13,N_2966,N_2972);
or UO_14 (O_14,N_2967,N_2974);
or UO_15 (O_15,N_2919,N_2979);
or UO_16 (O_16,N_2928,N_2941);
xnor UO_17 (O_17,N_2982,N_2987);
or UO_18 (O_18,N_2901,N_2980);
nand UO_19 (O_19,N_2992,N_2990);
and UO_20 (O_20,N_2945,N_2963);
and UO_21 (O_21,N_2935,N_2912);
nor UO_22 (O_22,N_2946,N_2902);
and UO_23 (O_23,N_2924,N_2981);
nor UO_24 (O_24,N_2995,N_2955);
and UO_25 (O_25,N_2937,N_2988);
and UO_26 (O_26,N_2993,N_2978);
and UO_27 (O_27,N_2986,N_2916);
xor UO_28 (O_28,N_2910,N_2961);
nor UO_29 (O_29,N_2959,N_2914);
or UO_30 (O_30,N_2926,N_2904);
nor UO_31 (O_31,N_2971,N_2932);
nor UO_32 (O_32,N_2999,N_2903);
nor UO_33 (O_33,N_2944,N_2920);
and UO_34 (O_34,N_2906,N_2950);
or UO_35 (O_35,N_2947,N_2948);
nor UO_36 (O_36,N_2917,N_2996);
or UO_37 (O_37,N_2923,N_2939);
or UO_38 (O_38,N_2956,N_2931);
nor UO_39 (O_39,N_2943,N_2951);
nand UO_40 (O_40,N_2949,N_2940);
or UO_41 (O_41,N_2925,N_2998);
or UO_42 (O_42,N_2969,N_2936);
or UO_43 (O_43,N_2921,N_2983);
nor UO_44 (O_44,N_2953,N_2934);
nand UO_45 (O_45,N_2985,N_2942);
nor UO_46 (O_46,N_2913,N_2973);
nor UO_47 (O_47,N_2915,N_2918);
nor UO_48 (O_48,N_2976,N_2970);
and UO_49 (O_49,N_2964,N_2907);
nor UO_50 (O_50,N_2956,N_2990);
nand UO_51 (O_51,N_2989,N_2906);
nor UO_52 (O_52,N_2994,N_2947);
or UO_53 (O_53,N_2905,N_2981);
and UO_54 (O_54,N_2978,N_2922);
nand UO_55 (O_55,N_2981,N_2961);
nand UO_56 (O_56,N_2907,N_2959);
nor UO_57 (O_57,N_2922,N_2914);
nand UO_58 (O_58,N_2979,N_2903);
xnor UO_59 (O_59,N_2903,N_2918);
or UO_60 (O_60,N_2901,N_2933);
nand UO_61 (O_61,N_2964,N_2908);
nor UO_62 (O_62,N_2903,N_2990);
and UO_63 (O_63,N_2973,N_2999);
nand UO_64 (O_64,N_2923,N_2924);
and UO_65 (O_65,N_2927,N_2914);
nand UO_66 (O_66,N_2970,N_2927);
or UO_67 (O_67,N_2909,N_2931);
or UO_68 (O_68,N_2947,N_2920);
and UO_69 (O_69,N_2980,N_2913);
nor UO_70 (O_70,N_2917,N_2941);
nor UO_71 (O_71,N_2910,N_2978);
xor UO_72 (O_72,N_2903,N_2993);
or UO_73 (O_73,N_2978,N_2958);
or UO_74 (O_74,N_2982,N_2932);
nor UO_75 (O_75,N_2954,N_2992);
nor UO_76 (O_76,N_2981,N_2955);
or UO_77 (O_77,N_2909,N_2980);
or UO_78 (O_78,N_2929,N_2969);
nand UO_79 (O_79,N_2984,N_2920);
xor UO_80 (O_80,N_2941,N_2985);
and UO_81 (O_81,N_2978,N_2906);
nor UO_82 (O_82,N_2941,N_2977);
nand UO_83 (O_83,N_2982,N_2901);
nand UO_84 (O_84,N_2968,N_2971);
or UO_85 (O_85,N_2934,N_2937);
and UO_86 (O_86,N_2980,N_2959);
and UO_87 (O_87,N_2995,N_2926);
or UO_88 (O_88,N_2902,N_2908);
and UO_89 (O_89,N_2929,N_2948);
and UO_90 (O_90,N_2904,N_2960);
nor UO_91 (O_91,N_2901,N_2936);
nor UO_92 (O_92,N_2963,N_2954);
or UO_93 (O_93,N_2972,N_2980);
or UO_94 (O_94,N_2954,N_2922);
nor UO_95 (O_95,N_2919,N_2951);
nand UO_96 (O_96,N_2977,N_2932);
nand UO_97 (O_97,N_2961,N_2926);
nor UO_98 (O_98,N_2950,N_2946);
nor UO_99 (O_99,N_2999,N_2957);
or UO_100 (O_100,N_2901,N_2967);
nor UO_101 (O_101,N_2949,N_2902);
and UO_102 (O_102,N_2917,N_2968);
nand UO_103 (O_103,N_2946,N_2962);
nand UO_104 (O_104,N_2996,N_2968);
or UO_105 (O_105,N_2970,N_2914);
and UO_106 (O_106,N_2971,N_2961);
and UO_107 (O_107,N_2929,N_2979);
nor UO_108 (O_108,N_2983,N_2925);
nor UO_109 (O_109,N_2931,N_2938);
nor UO_110 (O_110,N_2980,N_2927);
and UO_111 (O_111,N_2954,N_2984);
nand UO_112 (O_112,N_2991,N_2946);
nand UO_113 (O_113,N_2914,N_2947);
nor UO_114 (O_114,N_2980,N_2954);
nand UO_115 (O_115,N_2944,N_2993);
nor UO_116 (O_116,N_2999,N_2926);
or UO_117 (O_117,N_2953,N_2900);
or UO_118 (O_118,N_2989,N_2944);
or UO_119 (O_119,N_2984,N_2934);
or UO_120 (O_120,N_2933,N_2927);
nor UO_121 (O_121,N_2954,N_2917);
nand UO_122 (O_122,N_2999,N_2946);
nor UO_123 (O_123,N_2931,N_2990);
and UO_124 (O_124,N_2939,N_2974);
nor UO_125 (O_125,N_2923,N_2932);
nand UO_126 (O_126,N_2936,N_2945);
or UO_127 (O_127,N_2900,N_2945);
nand UO_128 (O_128,N_2986,N_2961);
nor UO_129 (O_129,N_2915,N_2904);
nand UO_130 (O_130,N_2924,N_2961);
and UO_131 (O_131,N_2947,N_2942);
and UO_132 (O_132,N_2923,N_2947);
or UO_133 (O_133,N_2981,N_2920);
and UO_134 (O_134,N_2939,N_2900);
and UO_135 (O_135,N_2905,N_2915);
or UO_136 (O_136,N_2957,N_2917);
and UO_137 (O_137,N_2951,N_2912);
nand UO_138 (O_138,N_2944,N_2981);
nand UO_139 (O_139,N_2977,N_2947);
xor UO_140 (O_140,N_2924,N_2952);
or UO_141 (O_141,N_2900,N_2955);
nor UO_142 (O_142,N_2988,N_2963);
nand UO_143 (O_143,N_2978,N_2955);
or UO_144 (O_144,N_2963,N_2946);
nor UO_145 (O_145,N_2954,N_2919);
and UO_146 (O_146,N_2931,N_2973);
nand UO_147 (O_147,N_2994,N_2927);
or UO_148 (O_148,N_2997,N_2985);
nand UO_149 (O_149,N_2960,N_2947);
nor UO_150 (O_150,N_2998,N_2929);
nand UO_151 (O_151,N_2925,N_2928);
or UO_152 (O_152,N_2933,N_2937);
nor UO_153 (O_153,N_2904,N_2929);
or UO_154 (O_154,N_2982,N_2900);
and UO_155 (O_155,N_2997,N_2987);
nand UO_156 (O_156,N_2921,N_2964);
nand UO_157 (O_157,N_2931,N_2942);
nor UO_158 (O_158,N_2981,N_2911);
or UO_159 (O_159,N_2907,N_2917);
or UO_160 (O_160,N_2974,N_2920);
or UO_161 (O_161,N_2927,N_2989);
nor UO_162 (O_162,N_2951,N_2923);
or UO_163 (O_163,N_2910,N_2927);
and UO_164 (O_164,N_2921,N_2938);
nor UO_165 (O_165,N_2944,N_2913);
nand UO_166 (O_166,N_2966,N_2985);
xnor UO_167 (O_167,N_2959,N_2909);
xnor UO_168 (O_168,N_2951,N_2942);
or UO_169 (O_169,N_2981,N_2945);
and UO_170 (O_170,N_2908,N_2943);
and UO_171 (O_171,N_2991,N_2925);
nor UO_172 (O_172,N_2922,N_2976);
and UO_173 (O_173,N_2924,N_2938);
nor UO_174 (O_174,N_2993,N_2994);
nor UO_175 (O_175,N_2995,N_2921);
nor UO_176 (O_176,N_2973,N_2917);
nand UO_177 (O_177,N_2918,N_2943);
and UO_178 (O_178,N_2999,N_2978);
nor UO_179 (O_179,N_2964,N_2971);
nor UO_180 (O_180,N_2919,N_2942);
and UO_181 (O_181,N_2923,N_2957);
and UO_182 (O_182,N_2990,N_2968);
or UO_183 (O_183,N_2908,N_2982);
or UO_184 (O_184,N_2985,N_2915);
and UO_185 (O_185,N_2947,N_2906);
nor UO_186 (O_186,N_2959,N_2934);
and UO_187 (O_187,N_2996,N_2904);
nor UO_188 (O_188,N_2978,N_2900);
and UO_189 (O_189,N_2986,N_2967);
and UO_190 (O_190,N_2946,N_2931);
or UO_191 (O_191,N_2970,N_2984);
or UO_192 (O_192,N_2932,N_2902);
nor UO_193 (O_193,N_2939,N_2919);
xnor UO_194 (O_194,N_2901,N_2985);
and UO_195 (O_195,N_2939,N_2986);
nor UO_196 (O_196,N_2918,N_2926);
and UO_197 (O_197,N_2980,N_2905);
or UO_198 (O_198,N_2985,N_2926);
and UO_199 (O_199,N_2939,N_2978);
or UO_200 (O_200,N_2966,N_2939);
nor UO_201 (O_201,N_2940,N_2901);
nand UO_202 (O_202,N_2937,N_2993);
nand UO_203 (O_203,N_2902,N_2940);
and UO_204 (O_204,N_2931,N_2929);
or UO_205 (O_205,N_2915,N_2924);
nor UO_206 (O_206,N_2984,N_2964);
nand UO_207 (O_207,N_2924,N_2934);
nand UO_208 (O_208,N_2978,N_2988);
or UO_209 (O_209,N_2923,N_2933);
and UO_210 (O_210,N_2929,N_2961);
nand UO_211 (O_211,N_2974,N_2963);
or UO_212 (O_212,N_2911,N_2936);
and UO_213 (O_213,N_2996,N_2964);
nand UO_214 (O_214,N_2941,N_2959);
nor UO_215 (O_215,N_2939,N_2933);
or UO_216 (O_216,N_2980,N_2973);
or UO_217 (O_217,N_2990,N_2991);
nand UO_218 (O_218,N_2997,N_2942);
nor UO_219 (O_219,N_2984,N_2940);
or UO_220 (O_220,N_2925,N_2964);
nand UO_221 (O_221,N_2956,N_2908);
or UO_222 (O_222,N_2951,N_2945);
nand UO_223 (O_223,N_2948,N_2989);
and UO_224 (O_224,N_2988,N_2952);
and UO_225 (O_225,N_2999,N_2977);
nor UO_226 (O_226,N_2977,N_2931);
and UO_227 (O_227,N_2990,N_2909);
or UO_228 (O_228,N_2950,N_2985);
or UO_229 (O_229,N_2952,N_2979);
nand UO_230 (O_230,N_2992,N_2941);
or UO_231 (O_231,N_2976,N_2913);
and UO_232 (O_232,N_2992,N_2914);
nand UO_233 (O_233,N_2925,N_2987);
nor UO_234 (O_234,N_2953,N_2994);
or UO_235 (O_235,N_2990,N_2978);
and UO_236 (O_236,N_2936,N_2977);
or UO_237 (O_237,N_2983,N_2958);
nand UO_238 (O_238,N_2963,N_2952);
nor UO_239 (O_239,N_2992,N_2907);
or UO_240 (O_240,N_2905,N_2959);
and UO_241 (O_241,N_2998,N_2909);
or UO_242 (O_242,N_2934,N_2956);
or UO_243 (O_243,N_2945,N_2970);
or UO_244 (O_244,N_2926,N_2917);
nand UO_245 (O_245,N_2916,N_2928);
and UO_246 (O_246,N_2934,N_2936);
and UO_247 (O_247,N_2906,N_2960);
or UO_248 (O_248,N_2974,N_2930);
or UO_249 (O_249,N_2956,N_2948);
or UO_250 (O_250,N_2935,N_2910);
or UO_251 (O_251,N_2962,N_2914);
and UO_252 (O_252,N_2991,N_2921);
or UO_253 (O_253,N_2944,N_2972);
or UO_254 (O_254,N_2940,N_2982);
and UO_255 (O_255,N_2923,N_2964);
nor UO_256 (O_256,N_2967,N_2960);
or UO_257 (O_257,N_2968,N_2993);
nand UO_258 (O_258,N_2988,N_2916);
nor UO_259 (O_259,N_2996,N_2912);
or UO_260 (O_260,N_2967,N_2998);
nand UO_261 (O_261,N_2910,N_2939);
and UO_262 (O_262,N_2942,N_2972);
nand UO_263 (O_263,N_2903,N_2967);
or UO_264 (O_264,N_2955,N_2972);
nor UO_265 (O_265,N_2959,N_2935);
nor UO_266 (O_266,N_2926,N_2929);
xnor UO_267 (O_267,N_2903,N_2923);
nor UO_268 (O_268,N_2935,N_2907);
nor UO_269 (O_269,N_2907,N_2926);
nor UO_270 (O_270,N_2915,N_2967);
or UO_271 (O_271,N_2922,N_2998);
or UO_272 (O_272,N_2966,N_2988);
nor UO_273 (O_273,N_2949,N_2926);
and UO_274 (O_274,N_2938,N_2905);
nor UO_275 (O_275,N_2957,N_2905);
and UO_276 (O_276,N_2949,N_2953);
nand UO_277 (O_277,N_2959,N_2962);
nand UO_278 (O_278,N_2986,N_2979);
and UO_279 (O_279,N_2906,N_2911);
nor UO_280 (O_280,N_2904,N_2905);
and UO_281 (O_281,N_2917,N_2913);
nor UO_282 (O_282,N_2983,N_2904);
nand UO_283 (O_283,N_2929,N_2946);
nor UO_284 (O_284,N_2989,N_2935);
nor UO_285 (O_285,N_2912,N_2910);
and UO_286 (O_286,N_2981,N_2959);
or UO_287 (O_287,N_2951,N_2946);
nand UO_288 (O_288,N_2902,N_2971);
or UO_289 (O_289,N_2982,N_2978);
nand UO_290 (O_290,N_2987,N_2986);
and UO_291 (O_291,N_2994,N_2921);
or UO_292 (O_292,N_2961,N_2953);
nand UO_293 (O_293,N_2925,N_2920);
and UO_294 (O_294,N_2932,N_2993);
nor UO_295 (O_295,N_2964,N_2986);
nand UO_296 (O_296,N_2977,N_2913);
and UO_297 (O_297,N_2907,N_2900);
and UO_298 (O_298,N_2985,N_2932);
nor UO_299 (O_299,N_2973,N_2930);
nor UO_300 (O_300,N_2928,N_2924);
nor UO_301 (O_301,N_2915,N_2961);
nor UO_302 (O_302,N_2921,N_2989);
or UO_303 (O_303,N_2901,N_2974);
and UO_304 (O_304,N_2990,N_2970);
nand UO_305 (O_305,N_2996,N_2934);
nand UO_306 (O_306,N_2925,N_2901);
nand UO_307 (O_307,N_2935,N_2932);
nor UO_308 (O_308,N_2928,N_2934);
and UO_309 (O_309,N_2921,N_2905);
nor UO_310 (O_310,N_2992,N_2920);
and UO_311 (O_311,N_2966,N_2997);
nand UO_312 (O_312,N_2975,N_2971);
nor UO_313 (O_313,N_2932,N_2922);
xor UO_314 (O_314,N_2911,N_2972);
xnor UO_315 (O_315,N_2985,N_2964);
or UO_316 (O_316,N_2911,N_2980);
nand UO_317 (O_317,N_2936,N_2980);
nor UO_318 (O_318,N_2900,N_2986);
nand UO_319 (O_319,N_2966,N_2950);
nand UO_320 (O_320,N_2957,N_2941);
or UO_321 (O_321,N_2959,N_2939);
or UO_322 (O_322,N_2942,N_2970);
and UO_323 (O_323,N_2978,N_2923);
nand UO_324 (O_324,N_2930,N_2995);
and UO_325 (O_325,N_2971,N_2946);
nand UO_326 (O_326,N_2961,N_2979);
nand UO_327 (O_327,N_2983,N_2939);
nor UO_328 (O_328,N_2913,N_2987);
and UO_329 (O_329,N_2945,N_2947);
nor UO_330 (O_330,N_2951,N_2917);
or UO_331 (O_331,N_2942,N_2941);
or UO_332 (O_332,N_2927,N_2981);
nand UO_333 (O_333,N_2992,N_2947);
nand UO_334 (O_334,N_2917,N_2909);
and UO_335 (O_335,N_2910,N_2907);
or UO_336 (O_336,N_2991,N_2922);
xor UO_337 (O_337,N_2982,N_2911);
and UO_338 (O_338,N_2943,N_2942);
and UO_339 (O_339,N_2942,N_2963);
or UO_340 (O_340,N_2923,N_2928);
or UO_341 (O_341,N_2995,N_2915);
and UO_342 (O_342,N_2938,N_2907);
nor UO_343 (O_343,N_2985,N_2998);
or UO_344 (O_344,N_2929,N_2999);
and UO_345 (O_345,N_2914,N_2928);
or UO_346 (O_346,N_2953,N_2915);
nand UO_347 (O_347,N_2989,N_2982);
nor UO_348 (O_348,N_2968,N_2982);
nor UO_349 (O_349,N_2950,N_2941);
or UO_350 (O_350,N_2922,N_2941);
xor UO_351 (O_351,N_2953,N_2996);
and UO_352 (O_352,N_2984,N_2917);
and UO_353 (O_353,N_2981,N_2999);
nand UO_354 (O_354,N_2900,N_2948);
and UO_355 (O_355,N_2914,N_2940);
or UO_356 (O_356,N_2952,N_2982);
or UO_357 (O_357,N_2955,N_2997);
or UO_358 (O_358,N_2922,N_2953);
nand UO_359 (O_359,N_2974,N_2962);
or UO_360 (O_360,N_2999,N_2906);
and UO_361 (O_361,N_2975,N_2987);
nand UO_362 (O_362,N_2953,N_2979);
nand UO_363 (O_363,N_2996,N_2928);
and UO_364 (O_364,N_2942,N_2915);
or UO_365 (O_365,N_2985,N_2927);
nor UO_366 (O_366,N_2926,N_2953);
or UO_367 (O_367,N_2953,N_2998);
nor UO_368 (O_368,N_2911,N_2977);
or UO_369 (O_369,N_2942,N_2964);
xnor UO_370 (O_370,N_2905,N_2998);
nand UO_371 (O_371,N_2954,N_2982);
and UO_372 (O_372,N_2907,N_2962);
or UO_373 (O_373,N_2908,N_2960);
and UO_374 (O_374,N_2907,N_2966);
or UO_375 (O_375,N_2955,N_2988);
nand UO_376 (O_376,N_2909,N_2949);
and UO_377 (O_377,N_2978,N_2965);
nor UO_378 (O_378,N_2919,N_2918);
nand UO_379 (O_379,N_2936,N_2941);
and UO_380 (O_380,N_2984,N_2988);
or UO_381 (O_381,N_2983,N_2963);
nor UO_382 (O_382,N_2918,N_2994);
nand UO_383 (O_383,N_2909,N_2964);
nor UO_384 (O_384,N_2930,N_2996);
or UO_385 (O_385,N_2945,N_2966);
and UO_386 (O_386,N_2914,N_2983);
nor UO_387 (O_387,N_2939,N_2957);
xnor UO_388 (O_388,N_2904,N_2969);
nand UO_389 (O_389,N_2980,N_2953);
nor UO_390 (O_390,N_2983,N_2970);
nand UO_391 (O_391,N_2981,N_2919);
nand UO_392 (O_392,N_2924,N_2905);
and UO_393 (O_393,N_2996,N_2907);
or UO_394 (O_394,N_2989,N_2995);
nand UO_395 (O_395,N_2910,N_2928);
xor UO_396 (O_396,N_2928,N_2944);
nand UO_397 (O_397,N_2981,N_2985);
nor UO_398 (O_398,N_2904,N_2940);
and UO_399 (O_399,N_2952,N_2901);
nor UO_400 (O_400,N_2905,N_2988);
nand UO_401 (O_401,N_2943,N_2986);
and UO_402 (O_402,N_2905,N_2991);
nand UO_403 (O_403,N_2985,N_2963);
or UO_404 (O_404,N_2935,N_2992);
or UO_405 (O_405,N_2966,N_2981);
nor UO_406 (O_406,N_2975,N_2973);
nand UO_407 (O_407,N_2961,N_2916);
or UO_408 (O_408,N_2902,N_2989);
and UO_409 (O_409,N_2991,N_2951);
and UO_410 (O_410,N_2976,N_2968);
or UO_411 (O_411,N_2931,N_2919);
nor UO_412 (O_412,N_2946,N_2998);
and UO_413 (O_413,N_2937,N_2928);
or UO_414 (O_414,N_2955,N_2914);
or UO_415 (O_415,N_2960,N_2969);
xor UO_416 (O_416,N_2925,N_2929);
nor UO_417 (O_417,N_2984,N_2948);
and UO_418 (O_418,N_2937,N_2965);
and UO_419 (O_419,N_2993,N_2973);
and UO_420 (O_420,N_2976,N_2929);
or UO_421 (O_421,N_2925,N_2902);
nor UO_422 (O_422,N_2932,N_2931);
or UO_423 (O_423,N_2904,N_2956);
nand UO_424 (O_424,N_2961,N_2968);
or UO_425 (O_425,N_2905,N_2941);
nand UO_426 (O_426,N_2965,N_2963);
nor UO_427 (O_427,N_2966,N_2965);
nor UO_428 (O_428,N_2917,N_2944);
nand UO_429 (O_429,N_2907,N_2945);
or UO_430 (O_430,N_2957,N_2956);
and UO_431 (O_431,N_2939,N_2903);
or UO_432 (O_432,N_2921,N_2929);
nor UO_433 (O_433,N_2969,N_2910);
nor UO_434 (O_434,N_2938,N_2965);
nand UO_435 (O_435,N_2985,N_2957);
or UO_436 (O_436,N_2991,N_2924);
and UO_437 (O_437,N_2950,N_2927);
nor UO_438 (O_438,N_2942,N_2956);
or UO_439 (O_439,N_2955,N_2951);
and UO_440 (O_440,N_2969,N_2974);
nand UO_441 (O_441,N_2963,N_2931);
nor UO_442 (O_442,N_2982,N_2934);
and UO_443 (O_443,N_2951,N_2924);
xor UO_444 (O_444,N_2937,N_2972);
nand UO_445 (O_445,N_2930,N_2991);
or UO_446 (O_446,N_2911,N_2948);
or UO_447 (O_447,N_2951,N_2953);
and UO_448 (O_448,N_2907,N_2995);
nand UO_449 (O_449,N_2942,N_2929);
and UO_450 (O_450,N_2992,N_2908);
and UO_451 (O_451,N_2951,N_2927);
nand UO_452 (O_452,N_2952,N_2906);
and UO_453 (O_453,N_2931,N_2908);
nor UO_454 (O_454,N_2921,N_2978);
or UO_455 (O_455,N_2975,N_2946);
xnor UO_456 (O_456,N_2943,N_2978);
and UO_457 (O_457,N_2993,N_2908);
nand UO_458 (O_458,N_2923,N_2927);
nor UO_459 (O_459,N_2995,N_2977);
nand UO_460 (O_460,N_2992,N_2956);
and UO_461 (O_461,N_2954,N_2935);
and UO_462 (O_462,N_2962,N_2963);
nor UO_463 (O_463,N_2928,N_2915);
nand UO_464 (O_464,N_2954,N_2939);
or UO_465 (O_465,N_2946,N_2919);
nand UO_466 (O_466,N_2947,N_2934);
nor UO_467 (O_467,N_2968,N_2941);
and UO_468 (O_468,N_2955,N_2938);
nor UO_469 (O_469,N_2903,N_2927);
and UO_470 (O_470,N_2900,N_2924);
and UO_471 (O_471,N_2912,N_2946);
xor UO_472 (O_472,N_2921,N_2912);
or UO_473 (O_473,N_2977,N_2904);
and UO_474 (O_474,N_2949,N_2903);
nor UO_475 (O_475,N_2996,N_2915);
or UO_476 (O_476,N_2910,N_2985);
and UO_477 (O_477,N_2957,N_2961);
and UO_478 (O_478,N_2905,N_2973);
nor UO_479 (O_479,N_2945,N_2967);
nand UO_480 (O_480,N_2943,N_2904);
and UO_481 (O_481,N_2914,N_2984);
and UO_482 (O_482,N_2919,N_2911);
nand UO_483 (O_483,N_2936,N_2949);
nand UO_484 (O_484,N_2900,N_2910);
nand UO_485 (O_485,N_2989,N_2936);
nor UO_486 (O_486,N_2906,N_2984);
nor UO_487 (O_487,N_2958,N_2935);
and UO_488 (O_488,N_2901,N_2906);
or UO_489 (O_489,N_2985,N_2918);
or UO_490 (O_490,N_2997,N_2995);
or UO_491 (O_491,N_2952,N_2915);
nor UO_492 (O_492,N_2999,N_2974);
nand UO_493 (O_493,N_2906,N_2959);
or UO_494 (O_494,N_2916,N_2979);
xor UO_495 (O_495,N_2909,N_2932);
or UO_496 (O_496,N_2994,N_2904);
or UO_497 (O_497,N_2980,N_2996);
and UO_498 (O_498,N_2977,N_2950);
xnor UO_499 (O_499,N_2978,N_2980);
endmodule