module basic_1000_10000_1500_5_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
xor U0 (N_0,In_210,In_156);
xor U1 (N_1,In_652,In_57);
or U2 (N_2,In_322,In_546);
and U3 (N_3,In_208,In_551);
and U4 (N_4,In_158,In_130);
xnor U5 (N_5,In_377,In_820);
and U6 (N_6,In_785,In_771);
xor U7 (N_7,In_943,In_618);
or U8 (N_8,In_650,In_687);
and U9 (N_9,In_343,In_327);
nor U10 (N_10,In_522,In_659);
or U11 (N_11,In_113,In_341);
or U12 (N_12,In_96,In_630);
or U13 (N_13,In_969,In_38);
and U14 (N_14,In_90,In_972);
nor U15 (N_15,In_892,In_496);
nand U16 (N_16,In_243,In_231);
xnor U17 (N_17,In_64,In_398);
and U18 (N_18,In_980,In_635);
xor U19 (N_19,In_338,In_395);
or U20 (N_20,In_403,In_601);
nand U21 (N_21,In_662,In_484);
nand U22 (N_22,In_886,In_281);
or U23 (N_23,In_367,In_29);
nor U24 (N_24,In_437,In_445);
xnor U25 (N_25,In_248,In_187);
or U26 (N_26,In_951,In_444);
xor U27 (N_27,In_100,In_110);
or U28 (N_28,In_720,In_303);
xor U29 (N_29,In_106,In_236);
nand U30 (N_30,In_238,In_558);
xnor U31 (N_31,In_518,In_702);
nor U32 (N_32,In_595,In_179);
xnor U33 (N_33,In_548,In_901);
xor U34 (N_34,In_394,In_351);
nand U35 (N_35,In_942,In_731);
and U36 (N_36,In_469,In_487);
nor U37 (N_37,In_644,In_597);
nand U38 (N_38,In_319,In_378);
xor U39 (N_39,In_946,In_163);
nand U40 (N_40,In_555,In_762);
and U41 (N_41,In_312,In_468);
or U42 (N_42,In_258,In_71);
nor U43 (N_43,In_107,In_693);
or U44 (N_44,In_356,In_973);
nand U45 (N_45,In_389,In_227);
and U46 (N_46,In_30,In_714);
nand U47 (N_47,In_162,In_837);
nor U48 (N_48,In_470,In_909);
nand U49 (N_49,In_218,In_192);
and U50 (N_50,In_481,In_178);
xnor U51 (N_51,In_70,In_845);
nor U52 (N_52,In_896,In_744);
and U53 (N_53,In_184,In_862);
and U54 (N_54,In_751,In_212);
nand U55 (N_55,In_968,In_617);
or U56 (N_56,In_126,In_274);
nor U57 (N_57,In_439,In_596);
nand U58 (N_58,In_455,In_554);
or U59 (N_59,In_682,In_935);
nand U60 (N_60,In_72,In_825);
xnor U61 (N_61,In_423,In_786);
or U62 (N_62,In_602,In_261);
nand U63 (N_63,In_399,In_414);
or U64 (N_64,In_703,In_260);
and U65 (N_65,In_730,In_373);
nand U66 (N_66,In_142,In_755);
nor U67 (N_67,In_957,In_342);
and U68 (N_68,In_902,In_707);
xnor U69 (N_69,In_194,In_51);
and U70 (N_70,In_308,In_473);
nand U71 (N_71,In_141,In_323);
xor U72 (N_72,In_748,In_987);
or U73 (N_73,In_257,In_101);
or U74 (N_74,In_18,In_516);
or U75 (N_75,In_19,In_76);
xnor U76 (N_76,In_186,In_801);
nor U77 (N_77,In_524,In_463);
xnor U78 (N_78,In_369,In_198);
or U79 (N_79,In_294,In_583);
and U80 (N_80,In_858,In_346);
nor U81 (N_81,In_893,In_181);
or U82 (N_82,In_937,In_0);
nand U83 (N_83,In_854,In_514);
and U84 (N_84,In_355,In_247);
xnor U85 (N_85,In_643,In_42);
nor U86 (N_86,In_229,In_796);
nand U87 (N_87,In_520,In_33);
or U88 (N_88,In_170,In_196);
xnor U89 (N_89,In_930,In_734);
nand U90 (N_90,In_872,In_784);
and U91 (N_91,In_381,In_613);
or U92 (N_92,In_759,In_647);
nor U93 (N_93,In_138,In_35);
xnor U94 (N_94,In_8,In_875);
and U95 (N_95,In_767,In_449);
or U96 (N_96,In_207,In_125);
or U97 (N_97,In_9,In_4);
nor U98 (N_98,In_637,In_807);
or U99 (N_99,In_663,In_136);
xnor U100 (N_100,In_692,In_954);
and U101 (N_101,In_386,In_735);
xor U102 (N_102,In_624,In_698);
or U103 (N_103,In_235,In_545);
or U104 (N_104,In_499,In_894);
and U105 (N_105,In_161,In_990);
and U106 (N_106,In_649,In_500);
and U107 (N_107,In_574,In_572);
nor U108 (N_108,In_953,In_855);
and U109 (N_109,In_453,In_22);
nand U110 (N_110,In_272,In_740);
nand U111 (N_111,In_92,In_991);
nand U112 (N_112,In_180,In_971);
or U113 (N_113,In_259,In_239);
and U114 (N_114,In_77,In_139);
or U115 (N_115,In_541,In_310);
xnor U116 (N_116,In_945,In_612);
nor U117 (N_117,In_674,In_465);
nor U118 (N_118,In_733,In_651);
nor U119 (N_119,In_360,In_581);
and U120 (N_120,In_315,In_653);
or U121 (N_121,In_561,In_93);
and U122 (N_122,In_223,In_599);
nand U123 (N_123,In_678,In_262);
nand U124 (N_124,In_409,In_864);
xnor U125 (N_125,In_82,In_17);
nor U126 (N_126,In_966,In_457);
nand U127 (N_127,In_506,In_590);
or U128 (N_128,In_150,In_411);
nand U129 (N_129,In_515,In_859);
or U130 (N_130,In_593,In_427);
or U131 (N_131,In_120,In_182);
or U132 (N_132,In_103,In_321);
nand U133 (N_133,In_206,In_47);
nand U134 (N_134,In_654,In_115);
nor U135 (N_135,In_448,In_766);
nor U136 (N_136,In_814,In_202);
or U137 (N_137,In_757,In_763);
xor U138 (N_138,In_401,In_527);
nor U139 (N_139,In_986,In_592);
nand U140 (N_140,In_298,In_293);
xnor U141 (N_141,In_795,In_52);
xor U142 (N_142,In_509,In_533);
or U143 (N_143,In_565,In_328);
or U144 (N_144,In_376,In_277);
nor U145 (N_145,In_970,In_679);
and U146 (N_146,In_668,In_419);
and U147 (N_147,In_627,In_1);
and U148 (N_148,In_94,In_721);
nand U149 (N_149,In_230,In_610);
nor U150 (N_150,In_958,In_454);
and U151 (N_151,In_718,In_523);
nor U152 (N_152,In_12,In_694);
xor U153 (N_153,In_648,In_62);
nand U154 (N_154,In_938,In_529);
nor U155 (N_155,In_217,In_812);
xor U156 (N_156,In_537,In_920);
nor U157 (N_157,In_884,In_406);
and U158 (N_158,In_21,In_549);
nand U159 (N_159,In_677,In_878);
nor U160 (N_160,In_568,In_646);
nand U161 (N_161,In_818,In_340);
and U162 (N_162,In_276,In_388);
or U163 (N_163,In_750,In_963);
nand U164 (N_164,In_225,In_889);
nor U165 (N_165,In_949,In_95);
xor U166 (N_166,In_686,In_24);
or U167 (N_167,In_810,In_80);
nor U168 (N_168,In_841,In_615);
nor U169 (N_169,In_540,In_416);
xnor U170 (N_170,In_768,In_944);
nand U171 (N_171,In_782,In_37);
xnor U172 (N_172,In_567,In_778);
nand U173 (N_173,In_984,In_933);
nand U174 (N_174,In_753,In_461);
nor U175 (N_175,In_111,In_405);
nor U176 (N_176,In_737,In_267);
and U177 (N_177,In_526,In_587);
nand U178 (N_178,In_667,In_263);
or U179 (N_179,In_370,In_988);
and U180 (N_180,In_904,In_844);
nand U181 (N_181,In_209,In_288);
or U182 (N_182,In_831,In_636);
and U183 (N_183,In_888,In_362);
xnor U184 (N_184,In_2,In_426);
xor U185 (N_185,In_477,In_255);
nor U186 (N_186,In_553,In_626);
or U187 (N_187,In_983,In_440);
xnor U188 (N_188,In_603,In_964);
or U189 (N_189,In_271,In_337);
or U190 (N_190,In_508,In_715);
or U191 (N_191,In_604,In_569);
or U192 (N_192,In_738,In_947);
nor U193 (N_193,In_912,In_234);
xnor U194 (N_194,In_726,In_577);
nand U195 (N_195,In_123,In_640);
or U196 (N_196,In_907,In_656);
nand U197 (N_197,In_25,In_49);
nand U198 (N_198,In_924,In_788);
and U199 (N_199,In_591,In_350);
nor U200 (N_200,In_368,In_169);
xor U201 (N_201,In_586,In_874);
nand U202 (N_202,In_332,In_127);
or U203 (N_203,In_780,In_977);
and U204 (N_204,In_998,In_89);
and U205 (N_205,In_512,In_366);
nor U206 (N_206,In_270,In_632);
nor U207 (N_207,In_441,In_460);
nor U208 (N_208,In_926,In_279);
xnor U209 (N_209,In_672,In_645);
xnor U210 (N_210,In_999,In_756);
and U211 (N_211,In_608,In_213);
or U212 (N_212,In_550,In_482);
xnor U213 (N_213,In_390,In_464);
xor U214 (N_214,In_916,In_564);
or U215 (N_215,In_16,In_189);
xor U216 (N_216,In_195,In_26);
nand U217 (N_217,In_976,In_530);
and U218 (N_218,In_879,In_598);
or U219 (N_219,In_696,In_299);
xnor U220 (N_220,In_869,In_559);
and U221 (N_221,In_917,In_794);
nand U222 (N_222,In_772,In_361);
and U223 (N_223,In_639,In_5);
nor U224 (N_224,In_900,In_83);
or U225 (N_225,In_291,In_839);
nand U226 (N_226,In_655,In_848);
or U227 (N_227,In_365,In_252);
or U228 (N_228,In_928,In_517);
or U229 (N_229,In_164,In_621);
or U230 (N_230,In_664,In_956);
and U231 (N_231,In_447,In_292);
xor U232 (N_232,In_967,In_224);
nor U233 (N_233,In_925,In_838);
nand U234 (N_234,In_249,In_326);
nor U235 (N_235,In_934,In_69);
xor U236 (N_236,In_456,In_697);
and U237 (N_237,In_681,In_675);
or U238 (N_238,In_191,In_266);
nor U239 (N_239,In_557,In_81);
nor U240 (N_240,In_725,In_713);
nor U241 (N_241,In_438,In_420);
nor U242 (N_242,In_396,In_826);
nand U243 (N_243,In_421,In_860);
or U244 (N_244,In_134,In_585);
xnor U245 (N_245,In_153,In_345);
and U246 (N_246,In_932,In_168);
nor U247 (N_247,In_695,In_352);
nor U248 (N_248,In_594,In_53);
xor U249 (N_249,In_711,In_578);
nand U250 (N_250,In_275,In_410);
nor U251 (N_251,In_467,In_485);
or U252 (N_252,In_190,In_579);
nor U253 (N_253,In_307,In_851);
or U254 (N_254,In_61,In_413);
and U255 (N_255,In_940,In_948);
nor U256 (N_256,In_962,In_774);
xnor U257 (N_257,In_911,In_472);
xor U258 (N_258,In_297,In_978);
nor U259 (N_259,In_769,In_129);
xnor U260 (N_260,In_392,In_98);
xor U261 (N_261,In_15,In_535);
nor U262 (N_262,In_54,In_65);
nand U263 (N_263,In_619,In_850);
and U264 (N_264,In_939,In_538);
or U265 (N_265,In_241,In_614);
xnor U266 (N_266,In_203,In_442);
nand U267 (N_267,In_105,In_741);
or U268 (N_268,In_324,In_348);
nor U269 (N_269,In_289,In_27);
nand U270 (N_270,In_85,In_489);
xnor U271 (N_271,In_880,In_278);
and U272 (N_272,In_840,In_476);
nand U273 (N_273,In_488,In_822);
or U274 (N_274,In_708,In_3);
xor U275 (N_275,In_211,In_435);
nand U276 (N_276,In_634,In_462);
and U277 (N_277,In_871,In_354);
xor U278 (N_278,In_995,In_913);
or U279 (N_279,In_919,In_14);
xor U280 (N_280,In_580,In_743);
xor U281 (N_281,In_495,In_765);
xor U282 (N_282,In_334,In_616);
and U283 (N_283,In_525,In_91);
nor U284 (N_284,In_317,In_719);
or U285 (N_285,In_480,In_511);
xnor U286 (N_286,In_959,In_283);
or U287 (N_287,In_867,In_996);
xor U288 (N_288,In_576,In_861);
nand U289 (N_289,In_280,In_295);
or U290 (N_290,In_330,In_539);
and U291 (N_291,In_177,In_6);
nand U292 (N_292,In_251,In_821);
xnor U293 (N_293,In_335,In_402);
xor U294 (N_294,In_269,In_805);
or U295 (N_295,In_357,In_287);
or U296 (N_296,In_471,In_185);
xor U297 (N_297,In_706,In_528);
nand U298 (N_298,In_232,In_952);
or U299 (N_299,In_791,In_119);
xor U300 (N_300,In_363,In_745);
nor U301 (N_301,In_443,In_176);
and U302 (N_302,In_400,In_23);
nor U303 (N_303,In_505,In_915);
and U304 (N_304,In_811,In_296);
or U305 (N_305,In_575,In_709);
and U306 (N_306,In_353,In_760);
xor U307 (N_307,In_46,In_143);
nand U308 (N_308,In_922,In_197);
nand U309 (N_309,In_974,In_620);
or U310 (N_310,In_333,In_781);
xor U311 (N_311,In_364,In_459);
and U312 (N_312,In_799,In_501);
nor U313 (N_313,In_797,In_425);
or U314 (N_314,In_7,In_905);
xor U315 (N_315,In_793,In_374);
nor U316 (N_316,In_382,In_131);
and U317 (N_317,In_84,In_975);
and U318 (N_318,In_140,In_710);
and U319 (N_319,In_857,In_723);
nand U320 (N_320,In_193,In_347);
nand U321 (N_321,In_237,In_205);
and U322 (N_322,In_918,In_490);
and U323 (N_323,In_10,In_349);
and U324 (N_324,In_955,In_493);
xor U325 (N_325,In_773,In_344);
or U326 (N_326,In_588,In_242);
and U327 (N_327,In_31,In_830);
or U328 (N_328,In_570,In_404);
xor U329 (N_329,In_228,In_44);
or U330 (N_330,In_633,In_43);
and U331 (N_331,In_311,In_746);
nor U332 (N_332,In_989,In_359);
nand U333 (N_333,In_384,In_834);
xor U334 (N_334,In_40,In_927);
xor U335 (N_335,In_117,In_669);
nor U336 (N_336,In_536,In_56);
and U337 (N_337,In_623,In_543);
nand U338 (N_338,In_318,In_770);
nand U339 (N_339,In_776,In_642);
or U340 (N_340,In_824,In_273);
and U341 (N_341,In_379,In_188);
nand U342 (N_342,In_430,In_846);
and U343 (N_343,In_112,In_104);
or U344 (N_344,In_705,In_124);
nor U345 (N_345,In_304,In_732);
or U346 (N_346,In_284,In_758);
or U347 (N_347,In_629,In_817);
nor U348 (N_348,In_658,In_552);
and U349 (N_349,In_775,In_547);
or U350 (N_350,In_865,In_563);
or U351 (N_351,In_691,In_246);
and U352 (N_352,In_700,In_183);
nor U353 (N_353,In_39,In_200);
nor U354 (N_354,In_50,In_783);
nor U355 (N_355,In_657,In_466);
xor U356 (N_356,In_428,In_132);
nand U357 (N_357,In_842,In_412);
nand U358 (N_358,In_531,In_173);
nand U359 (N_359,In_717,In_779);
xnor U360 (N_360,In_898,In_638);
nand U361 (N_361,In_78,In_336);
xor U362 (N_362,In_887,In_589);
or U363 (N_363,In_175,In_88);
nor U364 (N_364,In_159,In_128);
and U365 (N_365,In_285,In_899);
or U366 (N_366,In_253,In_240);
or U367 (N_367,In_148,In_739);
nand U368 (N_368,In_73,In_498);
and U369 (N_369,In_121,In_313);
or U370 (N_370,In_302,In_329);
xor U371 (N_371,In_316,In_923);
and U372 (N_372,In_729,In_849);
nand U373 (N_373,In_372,In_478);
nor U374 (N_374,In_688,In_155);
nand U375 (N_375,In_300,In_157);
xnor U376 (N_376,In_670,In_165);
nand U377 (N_377,In_600,In_789);
and U378 (N_378,In_813,In_254);
nor U379 (N_379,In_556,In_221);
xnor U380 (N_380,In_866,In_754);
and U381 (N_381,In_305,In_122);
and U382 (N_382,In_133,In_87);
nand U383 (N_383,In_256,In_172);
and U384 (N_384,In_97,In_214);
xor U385 (N_385,In_268,In_605);
xor U386 (N_386,In_60,In_408);
and U387 (N_387,In_167,In_146);
nand U388 (N_388,In_802,In_787);
and U389 (N_389,In_301,In_582);
and U390 (N_390,In_941,In_997);
nor U391 (N_391,In_245,In_680);
and U392 (N_392,In_833,In_808);
or U393 (N_393,In_532,In_562);
nand U394 (N_394,In_873,In_67);
nand U395 (N_395,In_171,In_827);
and U396 (N_396,In_75,In_761);
xnor U397 (N_397,In_936,In_513);
and U398 (N_398,In_339,In_566);
nand U399 (N_399,In_11,In_174);
xnor U400 (N_400,In_929,In_118);
and U401 (N_401,In_371,In_504);
nand U402 (N_402,In_832,In_204);
and U403 (N_403,In_145,In_584);
or U404 (N_404,In_79,In_885);
nor U405 (N_405,In_36,In_747);
or U406 (N_406,In_264,In_417);
nor U407 (N_407,In_137,In_41);
nor U408 (N_408,In_66,In_806);
or U409 (N_409,In_507,In_151);
and U410 (N_410,In_960,In_876);
nor U411 (N_411,In_607,In_154);
and U412 (N_412,In_828,In_676);
nor U413 (N_413,In_544,In_883);
xor U414 (N_414,In_809,In_109);
xnor U415 (N_415,In_432,In_314);
xor U416 (N_416,In_631,In_961);
xnor U417 (N_417,In_521,In_451);
or U418 (N_418,In_483,In_407);
nand U419 (N_419,In_752,In_215);
nand U420 (N_420,In_742,In_542);
xnor U421 (N_421,In_816,In_331);
nand U422 (N_422,In_910,In_931);
and U423 (N_423,In_147,In_994);
or U424 (N_424,In_309,In_503);
or U425 (N_425,In_397,In_868);
nand U426 (N_426,In_863,In_777);
nor U427 (N_427,In_474,In_68);
nand U428 (N_428,In_908,In_86);
nor U429 (N_429,In_573,In_375);
nor U430 (N_430,In_433,In_222);
xnor U431 (N_431,In_492,In_981);
xor U432 (N_432,In_722,In_727);
nor U433 (N_433,In_992,In_226);
and U434 (N_434,In_611,In_34);
or U435 (N_435,In_199,In_391);
nor U436 (N_436,In_690,In_114);
or U437 (N_437,In_728,In_571);
xnor U438 (N_438,In_422,In_149);
and U439 (N_439,In_244,In_921);
or U440 (N_440,In_479,In_829);
or U441 (N_441,In_689,In_877);
xnor U442 (N_442,In_99,In_673);
nand U443 (N_443,In_63,In_622);
and U444 (N_444,In_306,In_800);
xnor U445 (N_445,In_803,In_250);
and U446 (N_446,In_282,In_59);
nand U447 (N_447,In_666,In_609);
xnor U448 (N_448,In_606,In_393);
nor U449 (N_449,In_704,In_415);
xnor U450 (N_450,In_965,In_233);
or U451 (N_451,In_219,In_424);
and U452 (N_452,In_387,In_882);
nor U453 (N_453,In_431,In_950);
and U454 (N_454,In_665,In_320);
nor U455 (N_455,In_641,In_660);
and U456 (N_456,In_724,In_870);
or U457 (N_457,In_560,In_819);
nand U458 (N_458,In_475,In_993);
nand U459 (N_459,In_325,In_486);
nor U460 (N_460,In_661,In_701);
nor U461 (N_461,In_502,In_684);
and U462 (N_462,In_890,In_843);
or U463 (N_463,In_497,In_446);
or U464 (N_464,In_881,In_28);
and U465 (N_465,In_815,In_853);
xor U466 (N_466,In_856,In_804);
and U467 (N_467,In_903,In_358);
xnor U468 (N_468,In_20,In_982);
and U469 (N_469,In_434,In_102);
xor U470 (N_470,In_683,In_290);
nand U471 (N_471,In_716,In_792);
and U472 (N_472,In_286,In_450);
nor U473 (N_473,In_836,In_55);
nor U474 (N_474,In_265,In_625);
or U475 (N_475,In_510,In_895);
or U476 (N_476,In_380,In_458);
nand U477 (N_477,In_628,In_491);
nor U478 (N_478,In_45,In_13);
xnor U479 (N_479,In_429,In_534);
and U480 (N_480,In_712,In_736);
or U481 (N_481,In_852,In_914);
or U482 (N_482,In_452,In_671);
nand U483 (N_483,In_906,In_220);
and U484 (N_484,In_48,In_201);
xor U485 (N_485,In_798,In_823);
or U486 (N_486,In_383,In_74);
or U487 (N_487,In_160,In_436);
or U488 (N_488,In_152,In_699);
and U489 (N_489,In_764,In_32);
xnor U490 (N_490,In_144,In_135);
nand U491 (N_491,In_685,In_116);
and U492 (N_492,In_216,In_58);
or U493 (N_493,In_418,In_897);
and U494 (N_494,In_847,In_790);
or U495 (N_495,In_519,In_891);
and U496 (N_496,In_494,In_985);
nand U497 (N_497,In_979,In_108);
xor U498 (N_498,In_166,In_835);
nor U499 (N_499,In_385,In_749);
xnor U500 (N_500,In_296,In_605);
and U501 (N_501,In_36,In_782);
nand U502 (N_502,In_91,In_818);
and U503 (N_503,In_376,In_931);
or U504 (N_504,In_133,In_304);
xor U505 (N_505,In_261,In_140);
nor U506 (N_506,In_69,In_415);
nand U507 (N_507,In_540,In_553);
xor U508 (N_508,In_398,In_811);
or U509 (N_509,In_691,In_381);
nand U510 (N_510,In_747,In_324);
nand U511 (N_511,In_324,In_145);
and U512 (N_512,In_637,In_342);
or U513 (N_513,In_121,In_893);
xnor U514 (N_514,In_488,In_121);
or U515 (N_515,In_91,In_224);
nand U516 (N_516,In_934,In_989);
nor U517 (N_517,In_628,In_208);
nor U518 (N_518,In_256,In_461);
nor U519 (N_519,In_660,In_314);
nand U520 (N_520,In_114,In_861);
and U521 (N_521,In_13,In_465);
and U522 (N_522,In_544,In_630);
nand U523 (N_523,In_1,In_979);
and U524 (N_524,In_338,In_73);
nand U525 (N_525,In_157,In_778);
nand U526 (N_526,In_315,In_482);
and U527 (N_527,In_625,In_81);
xnor U528 (N_528,In_137,In_761);
and U529 (N_529,In_444,In_675);
nor U530 (N_530,In_863,In_64);
and U531 (N_531,In_605,In_21);
nand U532 (N_532,In_540,In_637);
xnor U533 (N_533,In_740,In_973);
xnor U534 (N_534,In_792,In_419);
xnor U535 (N_535,In_122,In_954);
xor U536 (N_536,In_152,In_22);
xor U537 (N_537,In_402,In_504);
nand U538 (N_538,In_69,In_391);
xor U539 (N_539,In_667,In_733);
nand U540 (N_540,In_136,In_479);
and U541 (N_541,In_135,In_168);
and U542 (N_542,In_145,In_466);
nor U543 (N_543,In_559,In_397);
nand U544 (N_544,In_334,In_326);
and U545 (N_545,In_4,In_892);
nand U546 (N_546,In_594,In_212);
and U547 (N_547,In_303,In_316);
nor U548 (N_548,In_719,In_33);
and U549 (N_549,In_134,In_963);
xnor U550 (N_550,In_860,In_426);
nor U551 (N_551,In_435,In_20);
nand U552 (N_552,In_10,In_176);
and U553 (N_553,In_227,In_799);
and U554 (N_554,In_83,In_532);
nor U555 (N_555,In_109,In_377);
nand U556 (N_556,In_648,In_199);
nand U557 (N_557,In_695,In_439);
xor U558 (N_558,In_662,In_258);
xor U559 (N_559,In_660,In_515);
nand U560 (N_560,In_169,In_628);
xor U561 (N_561,In_292,In_625);
nor U562 (N_562,In_848,In_482);
nand U563 (N_563,In_128,In_745);
and U564 (N_564,In_221,In_126);
nor U565 (N_565,In_79,In_637);
or U566 (N_566,In_762,In_725);
xor U567 (N_567,In_613,In_679);
nand U568 (N_568,In_75,In_137);
or U569 (N_569,In_515,In_673);
nand U570 (N_570,In_435,In_967);
and U571 (N_571,In_612,In_625);
nand U572 (N_572,In_52,In_305);
nor U573 (N_573,In_884,In_837);
xor U574 (N_574,In_385,In_936);
nor U575 (N_575,In_67,In_639);
nand U576 (N_576,In_268,In_909);
and U577 (N_577,In_221,In_733);
or U578 (N_578,In_361,In_419);
xnor U579 (N_579,In_778,In_915);
or U580 (N_580,In_814,In_842);
nand U581 (N_581,In_878,In_427);
nor U582 (N_582,In_66,In_187);
and U583 (N_583,In_60,In_627);
xor U584 (N_584,In_474,In_377);
nand U585 (N_585,In_370,In_201);
or U586 (N_586,In_439,In_824);
xor U587 (N_587,In_334,In_379);
nand U588 (N_588,In_691,In_273);
nor U589 (N_589,In_39,In_980);
and U590 (N_590,In_719,In_815);
nor U591 (N_591,In_145,In_648);
xnor U592 (N_592,In_552,In_698);
or U593 (N_593,In_814,In_55);
or U594 (N_594,In_274,In_898);
and U595 (N_595,In_441,In_759);
or U596 (N_596,In_145,In_797);
nor U597 (N_597,In_663,In_413);
nand U598 (N_598,In_189,In_870);
nand U599 (N_599,In_166,In_814);
and U600 (N_600,In_519,In_840);
nor U601 (N_601,In_522,In_314);
nor U602 (N_602,In_941,In_86);
and U603 (N_603,In_659,In_607);
xnor U604 (N_604,In_244,In_228);
nand U605 (N_605,In_536,In_633);
nor U606 (N_606,In_692,In_924);
or U607 (N_607,In_829,In_51);
nor U608 (N_608,In_643,In_793);
nor U609 (N_609,In_860,In_36);
xor U610 (N_610,In_326,In_292);
xor U611 (N_611,In_94,In_906);
and U612 (N_612,In_533,In_758);
nand U613 (N_613,In_330,In_205);
nand U614 (N_614,In_941,In_12);
xnor U615 (N_615,In_662,In_42);
nor U616 (N_616,In_553,In_189);
xor U617 (N_617,In_751,In_608);
nand U618 (N_618,In_77,In_417);
xnor U619 (N_619,In_21,In_759);
nor U620 (N_620,In_867,In_325);
nand U621 (N_621,In_33,In_545);
nand U622 (N_622,In_83,In_943);
nor U623 (N_623,In_266,In_988);
and U624 (N_624,In_793,In_110);
nand U625 (N_625,In_554,In_388);
nand U626 (N_626,In_767,In_592);
nor U627 (N_627,In_920,In_568);
nor U628 (N_628,In_282,In_924);
nor U629 (N_629,In_631,In_954);
or U630 (N_630,In_365,In_92);
xor U631 (N_631,In_476,In_98);
nor U632 (N_632,In_118,In_315);
xor U633 (N_633,In_72,In_972);
xnor U634 (N_634,In_39,In_539);
and U635 (N_635,In_698,In_908);
nor U636 (N_636,In_363,In_344);
nor U637 (N_637,In_661,In_468);
nand U638 (N_638,In_903,In_110);
and U639 (N_639,In_429,In_814);
and U640 (N_640,In_295,In_885);
and U641 (N_641,In_688,In_599);
and U642 (N_642,In_550,In_542);
nor U643 (N_643,In_170,In_23);
nand U644 (N_644,In_971,In_159);
or U645 (N_645,In_145,In_475);
xnor U646 (N_646,In_858,In_294);
nor U647 (N_647,In_856,In_629);
nor U648 (N_648,In_611,In_643);
nor U649 (N_649,In_163,In_43);
xor U650 (N_650,In_361,In_182);
xor U651 (N_651,In_718,In_16);
and U652 (N_652,In_382,In_865);
and U653 (N_653,In_83,In_824);
nand U654 (N_654,In_663,In_987);
nor U655 (N_655,In_130,In_864);
xnor U656 (N_656,In_818,In_845);
nand U657 (N_657,In_690,In_390);
or U658 (N_658,In_392,In_557);
nor U659 (N_659,In_960,In_867);
or U660 (N_660,In_299,In_596);
or U661 (N_661,In_910,In_259);
or U662 (N_662,In_825,In_517);
nand U663 (N_663,In_234,In_787);
and U664 (N_664,In_964,In_47);
xor U665 (N_665,In_363,In_512);
or U666 (N_666,In_530,In_868);
or U667 (N_667,In_929,In_121);
nand U668 (N_668,In_186,In_393);
nor U669 (N_669,In_330,In_588);
or U670 (N_670,In_222,In_976);
and U671 (N_671,In_84,In_613);
nor U672 (N_672,In_907,In_221);
or U673 (N_673,In_418,In_823);
nand U674 (N_674,In_543,In_754);
nor U675 (N_675,In_451,In_363);
nand U676 (N_676,In_152,In_934);
nand U677 (N_677,In_909,In_780);
nand U678 (N_678,In_993,In_716);
and U679 (N_679,In_92,In_173);
or U680 (N_680,In_942,In_297);
xnor U681 (N_681,In_571,In_599);
nor U682 (N_682,In_571,In_967);
or U683 (N_683,In_686,In_949);
and U684 (N_684,In_338,In_867);
nand U685 (N_685,In_725,In_73);
or U686 (N_686,In_977,In_884);
nor U687 (N_687,In_330,In_123);
xor U688 (N_688,In_783,In_897);
xor U689 (N_689,In_871,In_380);
and U690 (N_690,In_207,In_846);
xor U691 (N_691,In_41,In_926);
nor U692 (N_692,In_483,In_962);
or U693 (N_693,In_792,In_519);
nor U694 (N_694,In_44,In_831);
or U695 (N_695,In_725,In_570);
or U696 (N_696,In_970,In_764);
xor U697 (N_697,In_530,In_679);
and U698 (N_698,In_735,In_633);
nand U699 (N_699,In_543,In_498);
nor U700 (N_700,In_438,In_933);
xnor U701 (N_701,In_148,In_532);
nand U702 (N_702,In_406,In_324);
or U703 (N_703,In_55,In_121);
or U704 (N_704,In_630,In_601);
nand U705 (N_705,In_793,In_353);
nand U706 (N_706,In_270,In_698);
nand U707 (N_707,In_905,In_718);
or U708 (N_708,In_914,In_175);
xnor U709 (N_709,In_693,In_810);
or U710 (N_710,In_297,In_575);
or U711 (N_711,In_388,In_55);
nand U712 (N_712,In_785,In_451);
nor U713 (N_713,In_368,In_265);
or U714 (N_714,In_239,In_173);
or U715 (N_715,In_873,In_102);
and U716 (N_716,In_969,In_57);
or U717 (N_717,In_255,In_891);
nor U718 (N_718,In_381,In_621);
or U719 (N_719,In_730,In_275);
nand U720 (N_720,In_78,In_140);
or U721 (N_721,In_79,In_29);
and U722 (N_722,In_929,In_59);
and U723 (N_723,In_227,In_10);
nor U724 (N_724,In_819,In_675);
nand U725 (N_725,In_914,In_844);
xor U726 (N_726,In_896,In_826);
xnor U727 (N_727,In_896,In_938);
xor U728 (N_728,In_345,In_793);
and U729 (N_729,In_764,In_73);
or U730 (N_730,In_829,In_244);
xnor U731 (N_731,In_770,In_589);
and U732 (N_732,In_423,In_974);
or U733 (N_733,In_316,In_117);
nor U734 (N_734,In_260,In_75);
nor U735 (N_735,In_912,In_711);
or U736 (N_736,In_224,In_570);
or U737 (N_737,In_713,In_295);
and U738 (N_738,In_87,In_853);
xor U739 (N_739,In_150,In_8);
and U740 (N_740,In_973,In_828);
and U741 (N_741,In_297,In_891);
nor U742 (N_742,In_347,In_473);
nand U743 (N_743,In_790,In_139);
xnor U744 (N_744,In_494,In_310);
nor U745 (N_745,In_859,In_920);
and U746 (N_746,In_483,In_686);
nor U747 (N_747,In_487,In_228);
or U748 (N_748,In_841,In_824);
nor U749 (N_749,In_871,In_277);
xor U750 (N_750,In_740,In_805);
xor U751 (N_751,In_59,In_906);
xnor U752 (N_752,In_753,In_985);
xor U753 (N_753,In_457,In_168);
nor U754 (N_754,In_397,In_36);
or U755 (N_755,In_469,In_877);
or U756 (N_756,In_736,In_487);
nand U757 (N_757,In_894,In_834);
nor U758 (N_758,In_0,In_561);
and U759 (N_759,In_448,In_664);
or U760 (N_760,In_162,In_183);
and U761 (N_761,In_427,In_701);
or U762 (N_762,In_961,In_219);
xor U763 (N_763,In_107,In_365);
xor U764 (N_764,In_285,In_161);
nor U765 (N_765,In_14,In_573);
nand U766 (N_766,In_64,In_412);
and U767 (N_767,In_838,In_56);
nor U768 (N_768,In_973,In_108);
nor U769 (N_769,In_737,In_568);
nor U770 (N_770,In_586,In_199);
xnor U771 (N_771,In_644,In_692);
nand U772 (N_772,In_703,In_159);
and U773 (N_773,In_603,In_904);
or U774 (N_774,In_400,In_84);
nand U775 (N_775,In_109,In_868);
nand U776 (N_776,In_399,In_145);
xnor U777 (N_777,In_84,In_804);
nor U778 (N_778,In_371,In_279);
or U779 (N_779,In_686,In_699);
xnor U780 (N_780,In_933,In_340);
xor U781 (N_781,In_181,In_95);
xor U782 (N_782,In_466,In_574);
xnor U783 (N_783,In_474,In_25);
and U784 (N_784,In_359,In_345);
nand U785 (N_785,In_669,In_613);
nand U786 (N_786,In_380,In_192);
nand U787 (N_787,In_891,In_735);
nand U788 (N_788,In_759,In_654);
nand U789 (N_789,In_663,In_288);
xor U790 (N_790,In_530,In_238);
xnor U791 (N_791,In_864,In_796);
xnor U792 (N_792,In_921,In_395);
and U793 (N_793,In_289,In_511);
and U794 (N_794,In_156,In_529);
or U795 (N_795,In_171,In_444);
xnor U796 (N_796,In_72,In_299);
xnor U797 (N_797,In_519,In_174);
and U798 (N_798,In_965,In_498);
nor U799 (N_799,In_890,In_93);
nand U800 (N_800,In_873,In_833);
or U801 (N_801,In_442,In_801);
or U802 (N_802,In_447,In_708);
nand U803 (N_803,In_980,In_910);
nand U804 (N_804,In_97,In_45);
nand U805 (N_805,In_395,In_835);
nor U806 (N_806,In_689,In_7);
xor U807 (N_807,In_550,In_510);
or U808 (N_808,In_885,In_377);
or U809 (N_809,In_367,In_250);
and U810 (N_810,In_712,In_516);
or U811 (N_811,In_203,In_129);
or U812 (N_812,In_240,In_881);
or U813 (N_813,In_656,In_763);
nor U814 (N_814,In_544,In_606);
nand U815 (N_815,In_974,In_334);
and U816 (N_816,In_294,In_432);
xor U817 (N_817,In_295,In_58);
nand U818 (N_818,In_16,In_334);
nand U819 (N_819,In_5,In_709);
or U820 (N_820,In_614,In_77);
and U821 (N_821,In_233,In_207);
nor U822 (N_822,In_248,In_794);
and U823 (N_823,In_998,In_510);
xnor U824 (N_824,In_383,In_624);
and U825 (N_825,In_661,In_526);
xnor U826 (N_826,In_60,In_269);
or U827 (N_827,In_921,In_716);
xor U828 (N_828,In_731,In_963);
nand U829 (N_829,In_198,In_714);
nor U830 (N_830,In_627,In_932);
xor U831 (N_831,In_654,In_553);
or U832 (N_832,In_448,In_157);
nor U833 (N_833,In_920,In_452);
nand U834 (N_834,In_480,In_91);
nor U835 (N_835,In_829,In_590);
xor U836 (N_836,In_162,In_314);
nor U837 (N_837,In_231,In_726);
or U838 (N_838,In_718,In_135);
nand U839 (N_839,In_310,In_179);
nor U840 (N_840,In_465,In_129);
or U841 (N_841,In_67,In_827);
xnor U842 (N_842,In_668,In_494);
or U843 (N_843,In_70,In_521);
or U844 (N_844,In_711,In_239);
nand U845 (N_845,In_650,In_644);
nor U846 (N_846,In_877,In_504);
xnor U847 (N_847,In_942,In_273);
or U848 (N_848,In_690,In_293);
or U849 (N_849,In_418,In_46);
nor U850 (N_850,In_87,In_325);
and U851 (N_851,In_432,In_5);
and U852 (N_852,In_289,In_553);
or U853 (N_853,In_253,In_822);
and U854 (N_854,In_361,In_162);
xor U855 (N_855,In_938,In_922);
nor U856 (N_856,In_249,In_474);
and U857 (N_857,In_734,In_156);
and U858 (N_858,In_235,In_697);
and U859 (N_859,In_601,In_535);
nand U860 (N_860,In_521,In_315);
nor U861 (N_861,In_282,In_10);
nor U862 (N_862,In_306,In_59);
or U863 (N_863,In_590,In_63);
xnor U864 (N_864,In_769,In_167);
xor U865 (N_865,In_680,In_5);
or U866 (N_866,In_812,In_506);
and U867 (N_867,In_112,In_63);
or U868 (N_868,In_94,In_592);
or U869 (N_869,In_260,In_550);
nand U870 (N_870,In_987,In_937);
or U871 (N_871,In_596,In_433);
or U872 (N_872,In_202,In_437);
xnor U873 (N_873,In_556,In_56);
xnor U874 (N_874,In_213,In_760);
and U875 (N_875,In_933,In_915);
and U876 (N_876,In_579,In_410);
nor U877 (N_877,In_285,In_293);
nor U878 (N_878,In_860,In_48);
or U879 (N_879,In_138,In_240);
xnor U880 (N_880,In_580,In_15);
xnor U881 (N_881,In_731,In_584);
or U882 (N_882,In_584,In_630);
xnor U883 (N_883,In_517,In_572);
or U884 (N_884,In_763,In_874);
and U885 (N_885,In_642,In_495);
or U886 (N_886,In_661,In_223);
or U887 (N_887,In_954,In_2);
nand U888 (N_888,In_764,In_601);
or U889 (N_889,In_127,In_79);
nand U890 (N_890,In_246,In_433);
nor U891 (N_891,In_124,In_364);
xor U892 (N_892,In_373,In_640);
xnor U893 (N_893,In_574,In_236);
nor U894 (N_894,In_843,In_129);
nor U895 (N_895,In_313,In_895);
nor U896 (N_896,In_106,In_57);
nor U897 (N_897,In_442,In_923);
nand U898 (N_898,In_311,In_74);
nand U899 (N_899,In_516,In_525);
or U900 (N_900,In_56,In_640);
nand U901 (N_901,In_441,In_37);
nand U902 (N_902,In_545,In_865);
nor U903 (N_903,In_761,In_38);
nor U904 (N_904,In_483,In_287);
nand U905 (N_905,In_140,In_197);
or U906 (N_906,In_900,In_246);
nand U907 (N_907,In_772,In_369);
or U908 (N_908,In_790,In_62);
nor U909 (N_909,In_792,In_933);
nand U910 (N_910,In_398,In_700);
nor U911 (N_911,In_842,In_343);
nor U912 (N_912,In_133,In_169);
xor U913 (N_913,In_313,In_761);
nand U914 (N_914,In_284,In_445);
xnor U915 (N_915,In_4,In_396);
xor U916 (N_916,In_992,In_814);
nand U917 (N_917,In_187,In_166);
nand U918 (N_918,In_99,In_983);
or U919 (N_919,In_405,In_141);
nand U920 (N_920,In_198,In_69);
xnor U921 (N_921,In_648,In_592);
or U922 (N_922,In_777,In_284);
and U923 (N_923,In_166,In_624);
xor U924 (N_924,In_719,In_300);
nor U925 (N_925,In_988,In_703);
and U926 (N_926,In_958,In_427);
nand U927 (N_927,In_90,In_803);
and U928 (N_928,In_938,In_594);
xor U929 (N_929,In_759,In_961);
xnor U930 (N_930,In_940,In_7);
nor U931 (N_931,In_703,In_463);
or U932 (N_932,In_782,In_773);
nor U933 (N_933,In_991,In_395);
or U934 (N_934,In_521,In_368);
nor U935 (N_935,In_223,In_711);
or U936 (N_936,In_55,In_108);
nand U937 (N_937,In_856,In_204);
nand U938 (N_938,In_629,In_534);
and U939 (N_939,In_980,In_178);
nand U940 (N_940,In_778,In_667);
nand U941 (N_941,In_556,In_105);
xor U942 (N_942,In_305,In_956);
nor U943 (N_943,In_717,In_5);
nand U944 (N_944,In_453,In_975);
nand U945 (N_945,In_845,In_174);
or U946 (N_946,In_899,In_516);
xnor U947 (N_947,In_863,In_25);
or U948 (N_948,In_284,In_867);
nor U949 (N_949,In_726,In_522);
nand U950 (N_950,In_500,In_710);
and U951 (N_951,In_835,In_557);
nor U952 (N_952,In_761,In_327);
xor U953 (N_953,In_172,In_589);
nor U954 (N_954,In_477,In_276);
or U955 (N_955,In_882,In_806);
or U956 (N_956,In_573,In_474);
and U957 (N_957,In_144,In_874);
xor U958 (N_958,In_502,In_60);
xor U959 (N_959,In_397,In_808);
xor U960 (N_960,In_482,In_407);
xnor U961 (N_961,In_919,In_953);
and U962 (N_962,In_344,In_604);
and U963 (N_963,In_429,In_484);
or U964 (N_964,In_877,In_56);
nor U965 (N_965,In_433,In_789);
nor U966 (N_966,In_435,In_86);
nor U967 (N_967,In_773,In_299);
xnor U968 (N_968,In_98,In_517);
xnor U969 (N_969,In_907,In_321);
and U970 (N_970,In_0,In_621);
nand U971 (N_971,In_839,In_877);
nand U972 (N_972,In_118,In_993);
xor U973 (N_973,In_787,In_169);
or U974 (N_974,In_530,In_620);
nand U975 (N_975,In_816,In_537);
nand U976 (N_976,In_908,In_493);
or U977 (N_977,In_33,In_983);
xnor U978 (N_978,In_342,In_627);
xor U979 (N_979,In_834,In_366);
nor U980 (N_980,In_782,In_290);
nor U981 (N_981,In_967,In_41);
or U982 (N_982,In_11,In_595);
and U983 (N_983,In_687,In_635);
or U984 (N_984,In_16,In_963);
nand U985 (N_985,In_771,In_354);
and U986 (N_986,In_228,In_261);
nand U987 (N_987,In_799,In_347);
xnor U988 (N_988,In_686,In_928);
xor U989 (N_989,In_903,In_679);
and U990 (N_990,In_265,In_684);
xnor U991 (N_991,In_284,In_493);
and U992 (N_992,In_864,In_902);
and U993 (N_993,In_104,In_576);
nor U994 (N_994,In_549,In_29);
nand U995 (N_995,In_756,In_853);
nand U996 (N_996,In_247,In_689);
xor U997 (N_997,In_309,In_546);
nor U998 (N_998,In_127,In_314);
xor U999 (N_999,In_224,In_111);
nor U1000 (N_1000,In_106,In_659);
and U1001 (N_1001,In_114,In_200);
nand U1002 (N_1002,In_135,In_232);
xnor U1003 (N_1003,In_478,In_724);
and U1004 (N_1004,In_754,In_642);
nor U1005 (N_1005,In_990,In_79);
or U1006 (N_1006,In_909,In_348);
nor U1007 (N_1007,In_259,In_877);
and U1008 (N_1008,In_375,In_904);
or U1009 (N_1009,In_932,In_859);
xnor U1010 (N_1010,In_119,In_870);
or U1011 (N_1011,In_734,In_746);
xnor U1012 (N_1012,In_356,In_491);
xor U1013 (N_1013,In_344,In_253);
nor U1014 (N_1014,In_422,In_992);
nand U1015 (N_1015,In_764,In_517);
nand U1016 (N_1016,In_366,In_952);
xnor U1017 (N_1017,In_581,In_345);
or U1018 (N_1018,In_727,In_451);
and U1019 (N_1019,In_62,In_622);
nor U1020 (N_1020,In_632,In_10);
and U1021 (N_1021,In_47,In_222);
nand U1022 (N_1022,In_89,In_418);
or U1023 (N_1023,In_468,In_698);
xor U1024 (N_1024,In_944,In_234);
nor U1025 (N_1025,In_539,In_356);
and U1026 (N_1026,In_198,In_258);
nor U1027 (N_1027,In_322,In_407);
nor U1028 (N_1028,In_825,In_801);
xor U1029 (N_1029,In_373,In_556);
xnor U1030 (N_1030,In_614,In_856);
and U1031 (N_1031,In_509,In_824);
or U1032 (N_1032,In_643,In_26);
xor U1033 (N_1033,In_390,In_995);
nand U1034 (N_1034,In_794,In_242);
and U1035 (N_1035,In_609,In_899);
or U1036 (N_1036,In_484,In_711);
and U1037 (N_1037,In_166,In_64);
nor U1038 (N_1038,In_411,In_658);
nor U1039 (N_1039,In_966,In_471);
nor U1040 (N_1040,In_872,In_994);
nand U1041 (N_1041,In_32,In_579);
xnor U1042 (N_1042,In_363,In_384);
nor U1043 (N_1043,In_847,In_931);
and U1044 (N_1044,In_212,In_956);
and U1045 (N_1045,In_211,In_758);
or U1046 (N_1046,In_34,In_539);
or U1047 (N_1047,In_473,In_644);
nand U1048 (N_1048,In_626,In_804);
nand U1049 (N_1049,In_448,In_544);
nand U1050 (N_1050,In_822,In_256);
or U1051 (N_1051,In_85,In_108);
and U1052 (N_1052,In_743,In_549);
xnor U1053 (N_1053,In_604,In_722);
or U1054 (N_1054,In_567,In_507);
nor U1055 (N_1055,In_539,In_826);
xnor U1056 (N_1056,In_120,In_49);
xor U1057 (N_1057,In_561,In_373);
and U1058 (N_1058,In_28,In_96);
and U1059 (N_1059,In_740,In_112);
xor U1060 (N_1060,In_590,In_443);
xor U1061 (N_1061,In_617,In_909);
xnor U1062 (N_1062,In_393,In_922);
nor U1063 (N_1063,In_507,In_308);
or U1064 (N_1064,In_22,In_41);
xor U1065 (N_1065,In_847,In_806);
and U1066 (N_1066,In_555,In_597);
nand U1067 (N_1067,In_187,In_793);
and U1068 (N_1068,In_375,In_129);
xnor U1069 (N_1069,In_236,In_427);
nand U1070 (N_1070,In_332,In_578);
and U1071 (N_1071,In_933,In_337);
or U1072 (N_1072,In_111,In_900);
and U1073 (N_1073,In_598,In_114);
nor U1074 (N_1074,In_495,In_718);
or U1075 (N_1075,In_804,In_507);
or U1076 (N_1076,In_478,In_98);
or U1077 (N_1077,In_610,In_381);
and U1078 (N_1078,In_918,In_266);
and U1079 (N_1079,In_676,In_948);
xor U1080 (N_1080,In_215,In_232);
nand U1081 (N_1081,In_608,In_598);
xnor U1082 (N_1082,In_64,In_196);
nand U1083 (N_1083,In_105,In_340);
or U1084 (N_1084,In_695,In_932);
nand U1085 (N_1085,In_611,In_463);
nor U1086 (N_1086,In_527,In_692);
nand U1087 (N_1087,In_249,In_544);
and U1088 (N_1088,In_468,In_72);
nand U1089 (N_1089,In_113,In_500);
xor U1090 (N_1090,In_405,In_14);
nand U1091 (N_1091,In_218,In_897);
or U1092 (N_1092,In_667,In_302);
and U1093 (N_1093,In_488,In_878);
nor U1094 (N_1094,In_286,In_3);
or U1095 (N_1095,In_851,In_547);
nand U1096 (N_1096,In_810,In_289);
xor U1097 (N_1097,In_434,In_851);
and U1098 (N_1098,In_268,In_37);
and U1099 (N_1099,In_96,In_140);
nor U1100 (N_1100,In_496,In_928);
nand U1101 (N_1101,In_960,In_986);
xor U1102 (N_1102,In_100,In_463);
xor U1103 (N_1103,In_820,In_923);
xnor U1104 (N_1104,In_712,In_324);
or U1105 (N_1105,In_924,In_605);
nor U1106 (N_1106,In_295,In_162);
and U1107 (N_1107,In_192,In_947);
nand U1108 (N_1108,In_946,In_854);
nand U1109 (N_1109,In_656,In_780);
xnor U1110 (N_1110,In_427,In_590);
nor U1111 (N_1111,In_898,In_442);
and U1112 (N_1112,In_195,In_692);
or U1113 (N_1113,In_658,In_320);
and U1114 (N_1114,In_682,In_832);
nor U1115 (N_1115,In_25,In_547);
and U1116 (N_1116,In_446,In_325);
and U1117 (N_1117,In_428,In_745);
nor U1118 (N_1118,In_533,In_285);
or U1119 (N_1119,In_183,In_400);
nor U1120 (N_1120,In_858,In_792);
nor U1121 (N_1121,In_933,In_168);
and U1122 (N_1122,In_347,In_420);
xnor U1123 (N_1123,In_553,In_697);
xor U1124 (N_1124,In_485,In_938);
or U1125 (N_1125,In_639,In_162);
or U1126 (N_1126,In_884,In_448);
xnor U1127 (N_1127,In_77,In_89);
nor U1128 (N_1128,In_218,In_709);
xor U1129 (N_1129,In_579,In_970);
nand U1130 (N_1130,In_370,In_407);
and U1131 (N_1131,In_242,In_297);
nand U1132 (N_1132,In_678,In_379);
and U1133 (N_1133,In_154,In_943);
nor U1134 (N_1134,In_976,In_516);
nor U1135 (N_1135,In_454,In_31);
or U1136 (N_1136,In_23,In_295);
nor U1137 (N_1137,In_396,In_370);
and U1138 (N_1138,In_317,In_841);
or U1139 (N_1139,In_148,In_491);
xor U1140 (N_1140,In_509,In_337);
xor U1141 (N_1141,In_425,In_958);
and U1142 (N_1142,In_230,In_684);
and U1143 (N_1143,In_267,In_939);
or U1144 (N_1144,In_194,In_359);
or U1145 (N_1145,In_43,In_534);
nand U1146 (N_1146,In_142,In_434);
nand U1147 (N_1147,In_181,In_271);
and U1148 (N_1148,In_206,In_510);
and U1149 (N_1149,In_4,In_45);
nand U1150 (N_1150,In_601,In_50);
or U1151 (N_1151,In_869,In_34);
and U1152 (N_1152,In_26,In_843);
nor U1153 (N_1153,In_198,In_879);
or U1154 (N_1154,In_807,In_386);
or U1155 (N_1155,In_509,In_426);
xnor U1156 (N_1156,In_666,In_118);
nor U1157 (N_1157,In_323,In_686);
or U1158 (N_1158,In_611,In_766);
nor U1159 (N_1159,In_768,In_518);
nor U1160 (N_1160,In_571,In_477);
nor U1161 (N_1161,In_959,In_965);
xnor U1162 (N_1162,In_480,In_958);
xnor U1163 (N_1163,In_21,In_668);
or U1164 (N_1164,In_342,In_771);
nor U1165 (N_1165,In_871,In_861);
xor U1166 (N_1166,In_883,In_585);
or U1167 (N_1167,In_482,In_72);
or U1168 (N_1168,In_960,In_498);
and U1169 (N_1169,In_274,In_823);
xor U1170 (N_1170,In_728,In_809);
nand U1171 (N_1171,In_355,In_864);
nor U1172 (N_1172,In_324,In_868);
nand U1173 (N_1173,In_795,In_259);
and U1174 (N_1174,In_453,In_832);
and U1175 (N_1175,In_363,In_772);
and U1176 (N_1176,In_450,In_716);
and U1177 (N_1177,In_567,In_948);
or U1178 (N_1178,In_459,In_832);
nor U1179 (N_1179,In_964,In_192);
nor U1180 (N_1180,In_520,In_1);
nor U1181 (N_1181,In_774,In_240);
and U1182 (N_1182,In_252,In_805);
nand U1183 (N_1183,In_850,In_326);
xor U1184 (N_1184,In_246,In_878);
and U1185 (N_1185,In_630,In_400);
xnor U1186 (N_1186,In_641,In_576);
xnor U1187 (N_1187,In_478,In_371);
and U1188 (N_1188,In_595,In_684);
nor U1189 (N_1189,In_356,In_14);
and U1190 (N_1190,In_826,In_563);
xor U1191 (N_1191,In_43,In_751);
xor U1192 (N_1192,In_596,In_2);
nor U1193 (N_1193,In_489,In_232);
or U1194 (N_1194,In_94,In_875);
or U1195 (N_1195,In_860,In_492);
or U1196 (N_1196,In_217,In_467);
nor U1197 (N_1197,In_370,In_631);
nor U1198 (N_1198,In_755,In_537);
or U1199 (N_1199,In_883,In_274);
nor U1200 (N_1200,In_170,In_283);
or U1201 (N_1201,In_481,In_950);
and U1202 (N_1202,In_746,In_870);
xnor U1203 (N_1203,In_483,In_23);
and U1204 (N_1204,In_408,In_320);
xor U1205 (N_1205,In_11,In_766);
or U1206 (N_1206,In_667,In_702);
xor U1207 (N_1207,In_266,In_774);
or U1208 (N_1208,In_222,In_395);
nand U1209 (N_1209,In_926,In_994);
xnor U1210 (N_1210,In_215,In_412);
or U1211 (N_1211,In_426,In_982);
nand U1212 (N_1212,In_377,In_485);
and U1213 (N_1213,In_692,In_718);
and U1214 (N_1214,In_791,In_722);
nand U1215 (N_1215,In_383,In_250);
xnor U1216 (N_1216,In_860,In_275);
xor U1217 (N_1217,In_751,In_298);
xor U1218 (N_1218,In_711,In_772);
nor U1219 (N_1219,In_580,In_933);
nand U1220 (N_1220,In_752,In_316);
and U1221 (N_1221,In_208,In_552);
or U1222 (N_1222,In_443,In_753);
and U1223 (N_1223,In_920,In_183);
nor U1224 (N_1224,In_902,In_535);
nand U1225 (N_1225,In_192,In_753);
or U1226 (N_1226,In_95,In_327);
nand U1227 (N_1227,In_361,In_362);
nand U1228 (N_1228,In_430,In_183);
and U1229 (N_1229,In_327,In_188);
nand U1230 (N_1230,In_238,In_863);
and U1231 (N_1231,In_619,In_164);
nand U1232 (N_1232,In_392,In_871);
and U1233 (N_1233,In_764,In_204);
or U1234 (N_1234,In_205,In_720);
nand U1235 (N_1235,In_214,In_306);
xnor U1236 (N_1236,In_66,In_947);
or U1237 (N_1237,In_250,In_833);
and U1238 (N_1238,In_312,In_53);
or U1239 (N_1239,In_817,In_781);
xor U1240 (N_1240,In_59,In_238);
nand U1241 (N_1241,In_769,In_540);
or U1242 (N_1242,In_636,In_848);
xnor U1243 (N_1243,In_423,In_200);
xor U1244 (N_1244,In_837,In_552);
and U1245 (N_1245,In_840,In_795);
nor U1246 (N_1246,In_765,In_469);
or U1247 (N_1247,In_386,In_831);
xor U1248 (N_1248,In_49,In_826);
and U1249 (N_1249,In_169,In_170);
nor U1250 (N_1250,In_208,In_134);
and U1251 (N_1251,In_468,In_63);
xor U1252 (N_1252,In_336,In_527);
nand U1253 (N_1253,In_139,In_192);
and U1254 (N_1254,In_777,In_723);
or U1255 (N_1255,In_264,In_961);
nand U1256 (N_1256,In_659,In_325);
or U1257 (N_1257,In_522,In_340);
nor U1258 (N_1258,In_854,In_174);
xor U1259 (N_1259,In_504,In_191);
nor U1260 (N_1260,In_531,In_450);
nand U1261 (N_1261,In_541,In_551);
or U1262 (N_1262,In_433,In_272);
xor U1263 (N_1263,In_384,In_805);
and U1264 (N_1264,In_30,In_194);
and U1265 (N_1265,In_367,In_856);
or U1266 (N_1266,In_713,In_931);
nor U1267 (N_1267,In_247,In_623);
nand U1268 (N_1268,In_706,In_411);
nand U1269 (N_1269,In_740,In_704);
xnor U1270 (N_1270,In_622,In_572);
nor U1271 (N_1271,In_247,In_174);
nand U1272 (N_1272,In_146,In_505);
or U1273 (N_1273,In_671,In_555);
or U1274 (N_1274,In_610,In_199);
nor U1275 (N_1275,In_198,In_407);
or U1276 (N_1276,In_723,In_254);
xor U1277 (N_1277,In_93,In_400);
nor U1278 (N_1278,In_115,In_329);
xor U1279 (N_1279,In_442,In_661);
nor U1280 (N_1280,In_815,In_825);
nor U1281 (N_1281,In_91,In_970);
nand U1282 (N_1282,In_530,In_222);
nand U1283 (N_1283,In_824,In_449);
nor U1284 (N_1284,In_457,In_333);
or U1285 (N_1285,In_97,In_672);
nand U1286 (N_1286,In_599,In_562);
nand U1287 (N_1287,In_807,In_256);
and U1288 (N_1288,In_917,In_54);
and U1289 (N_1289,In_267,In_206);
or U1290 (N_1290,In_478,In_844);
nand U1291 (N_1291,In_382,In_927);
xor U1292 (N_1292,In_894,In_520);
or U1293 (N_1293,In_184,In_63);
nor U1294 (N_1294,In_440,In_836);
nand U1295 (N_1295,In_454,In_641);
nand U1296 (N_1296,In_258,In_363);
xnor U1297 (N_1297,In_734,In_383);
nand U1298 (N_1298,In_979,In_125);
and U1299 (N_1299,In_539,In_723);
nor U1300 (N_1300,In_704,In_568);
nand U1301 (N_1301,In_151,In_349);
xnor U1302 (N_1302,In_182,In_393);
or U1303 (N_1303,In_697,In_64);
nor U1304 (N_1304,In_41,In_123);
xnor U1305 (N_1305,In_351,In_845);
nor U1306 (N_1306,In_589,In_562);
and U1307 (N_1307,In_894,In_714);
nand U1308 (N_1308,In_869,In_799);
nand U1309 (N_1309,In_335,In_103);
or U1310 (N_1310,In_275,In_979);
nor U1311 (N_1311,In_49,In_83);
nand U1312 (N_1312,In_120,In_331);
xor U1313 (N_1313,In_251,In_231);
xnor U1314 (N_1314,In_826,In_395);
or U1315 (N_1315,In_143,In_204);
and U1316 (N_1316,In_286,In_435);
and U1317 (N_1317,In_968,In_626);
and U1318 (N_1318,In_197,In_892);
or U1319 (N_1319,In_366,In_567);
nor U1320 (N_1320,In_990,In_151);
or U1321 (N_1321,In_446,In_575);
or U1322 (N_1322,In_132,In_415);
or U1323 (N_1323,In_867,In_499);
nand U1324 (N_1324,In_268,In_892);
and U1325 (N_1325,In_425,In_459);
and U1326 (N_1326,In_301,In_944);
or U1327 (N_1327,In_935,In_906);
nand U1328 (N_1328,In_308,In_981);
and U1329 (N_1329,In_761,In_446);
xor U1330 (N_1330,In_71,In_842);
and U1331 (N_1331,In_698,In_36);
nor U1332 (N_1332,In_649,In_973);
and U1333 (N_1333,In_201,In_847);
nand U1334 (N_1334,In_774,In_628);
or U1335 (N_1335,In_450,In_800);
nand U1336 (N_1336,In_975,In_846);
xnor U1337 (N_1337,In_596,In_718);
nor U1338 (N_1338,In_777,In_124);
nor U1339 (N_1339,In_617,In_805);
nand U1340 (N_1340,In_654,In_539);
xnor U1341 (N_1341,In_931,In_969);
nor U1342 (N_1342,In_932,In_317);
or U1343 (N_1343,In_408,In_87);
xnor U1344 (N_1344,In_824,In_223);
and U1345 (N_1345,In_113,In_136);
or U1346 (N_1346,In_967,In_25);
and U1347 (N_1347,In_820,In_768);
nor U1348 (N_1348,In_804,In_316);
or U1349 (N_1349,In_295,In_599);
nand U1350 (N_1350,In_562,In_282);
nor U1351 (N_1351,In_308,In_164);
xnor U1352 (N_1352,In_609,In_51);
nand U1353 (N_1353,In_352,In_643);
or U1354 (N_1354,In_801,In_214);
or U1355 (N_1355,In_852,In_82);
xor U1356 (N_1356,In_318,In_125);
nor U1357 (N_1357,In_536,In_250);
nor U1358 (N_1358,In_379,In_328);
or U1359 (N_1359,In_81,In_366);
nor U1360 (N_1360,In_85,In_678);
nor U1361 (N_1361,In_367,In_255);
nor U1362 (N_1362,In_562,In_383);
nand U1363 (N_1363,In_98,In_137);
nand U1364 (N_1364,In_499,In_822);
or U1365 (N_1365,In_841,In_66);
and U1366 (N_1366,In_280,In_698);
xor U1367 (N_1367,In_76,In_306);
or U1368 (N_1368,In_262,In_515);
and U1369 (N_1369,In_489,In_274);
nor U1370 (N_1370,In_886,In_680);
xor U1371 (N_1371,In_618,In_638);
or U1372 (N_1372,In_599,In_548);
and U1373 (N_1373,In_881,In_779);
nand U1374 (N_1374,In_541,In_165);
xor U1375 (N_1375,In_728,In_758);
nand U1376 (N_1376,In_678,In_559);
or U1377 (N_1377,In_37,In_550);
and U1378 (N_1378,In_711,In_158);
and U1379 (N_1379,In_751,In_18);
nand U1380 (N_1380,In_93,In_391);
nor U1381 (N_1381,In_265,In_767);
xor U1382 (N_1382,In_966,In_930);
nand U1383 (N_1383,In_597,In_993);
and U1384 (N_1384,In_927,In_771);
nor U1385 (N_1385,In_192,In_125);
xnor U1386 (N_1386,In_223,In_935);
nor U1387 (N_1387,In_674,In_566);
nor U1388 (N_1388,In_547,In_692);
nand U1389 (N_1389,In_685,In_529);
xor U1390 (N_1390,In_580,In_826);
and U1391 (N_1391,In_515,In_606);
xnor U1392 (N_1392,In_605,In_220);
and U1393 (N_1393,In_861,In_898);
xor U1394 (N_1394,In_7,In_904);
nor U1395 (N_1395,In_353,In_945);
nand U1396 (N_1396,In_840,In_468);
nor U1397 (N_1397,In_102,In_787);
and U1398 (N_1398,In_669,In_522);
or U1399 (N_1399,In_429,In_821);
or U1400 (N_1400,In_964,In_864);
nand U1401 (N_1401,In_316,In_865);
xor U1402 (N_1402,In_113,In_946);
or U1403 (N_1403,In_240,In_444);
nand U1404 (N_1404,In_690,In_284);
and U1405 (N_1405,In_53,In_893);
nand U1406 (N_1406,In_692,In_858);
nand U1407 (N_1407,In_694,In_731);
and U1408 (N_1408,In_524,In_862);
nor U1409 (N_1409,In_522,In_140);
or U1410 (N_1410,In_260,In_795);
nand U1411 (N_1411,In_613,In_859);
nand U1412 (N_1412,In_368,In_419);
nand U1413 (N_1413,In_375,In_932);
xnor U1414 (N_1414,In_16,In_683);
and U1415 (N_1415,In_127,In_425);
xor U1416 (N_1416,In_301,In_430);
xnor U1417 (N_1417,In_712,In_863);
nand U1418 (N_1418,In_339,In_271);
xnor U1419 (N_1419,In_617,In_9);
nand U1420 (N_1420,In_66,In_702);
nand U1421 (N_1421,In_992,In_577);
nand U1422 (N_1422,In_960,In_938);
nand U1423 (N_1423,In_967,In_874);
xnor U1424 (N_1424,In_626,In_832);
nor U1425 (N_1425,In_762,In_988);
nand U1426 (N_1426,In_646,In_201);
xor U1427 (N_1427,In_554,In_608);
xnor U1428 (N_1428,In_921,In_625);
or U1429 (N_1429,In_456,In_788);
and U1430 (N_1430,In_441,In_474);
and U1431 (N_1431,In_51,In_221);
or U1432 (N_1432,In_201,In_356);
nor U1433 (N_1433,In_280,In_366);
and U1434 (N_1434,In_473,In_285);
and U1435 (N_1435,In_15,In_566);
or U1436 (N_1436,In_704,In_926);
or U1437 (N_1437,In_618,In_774);
and U1438 (N_1438,In_271,In_617);
nor U1439 (N_1439,In_37,In_741);
xnor U1440 (N_1440,In_241,In_542);
nand U1441 (N_1441,In_177,In_221);
and U1442 (N_1442,In_145,In_353);
or U1443 (N_1443,In_419,In_590);
xor U1444 (N_1444,In_92,In_873);
nand U1445 (N_1445,In_805,In_180);
nor U1446 (N_1446,In_126,In_252);
or U1447 (N_1447,In_114,In_365);
xor U1448 (N_1448,In_841,In_649);
or U1449 (N_1449,In_46,In_694);
and U1450 (N_1450,In_735,In_938);
nor U1451 (N_1451,In_438,In_753);
nand U1452 (N_1452,In_662,In_829);
nand U1453 (N_1453,In_557,In_0);
xor U1454 (N_1454,In_984,In_423);
nor U1455 (N_1455,In_591,In_77);
nand U1456 (N_1456,In_157,In_873);
nor U1457 (N_1457,In_697,In_780);
nor U1458 (N_1458,In_75,In_835);
xor U1459 (N_1459,In_184,In_579);
nor U1460 (N_1460,In_745,In_890);
nor U1461 (N_1461,In_150,In_550);
nor U1462 (N_1462,In_653,In_962);
nor U1463 (N_1463,In_291,In_110);
and U1464 (N_1464,In_281,In_831);
nor U1465 (N_1465,In_989,In_727);
or U1466 (N_1466,In_44,In_501);
xor U1467 (N_1467,In_338,In_68);
xor U1468 (N_1468,In_69,In_545);
nor U1469 (N_1469,In_540,In_554);
nor U1470 (N_1470,In_576,In_39);
or U1471 (N_1471,In_577,In_281);
nand U1472 (N_1472,In_935,In_386);
and U1473 (N_1473,In_777,In_228);
nand U1474 (N_1474,In_193,In_215);
and U1475 (N_1475,In_784,In_287);
nand U1476 (N_1476,In_914,In_768);
nor U1477 (N_1477,In_740,In_882);
xnor U1478 (N_1478,In_397,In_189);
nor U1479 (N_1479,In_190,In_92);
nand U1480 (N_1480,In_907,In_903);
nand U1481 (N_1481,In_984,In_995);
or U1482 (N_1482,In_433,In_923);
and U1483 (N_1483,In_871,In_262);
nor U1484 (N_1484,In_569,In_480);
nand U1485 (N_1485,In_14,In_125);
and U1486 (N_1486,In_940,In_201);
nor U1487 (N_1487,In_896,In_666);
and U1488 (N_1488,In_508,In_385);
and U1489 (N_1489,In_460,In_128);
xor U1490 (N_1490,In_774,In_136);
xnor U1491 (N_1491,In_433,In_893);
or U1492 (N_1492,In_501,In_79);
and U1493 (N_1493,In_599,In_690);
or U1494 (N_1494,In_791,In_755);
nand U1495 (N_1495,In_874,In_143);
nor U1496 (N_1496,In_164,In_778);
and U1497 (N_1497,In_803,In_62);
nand U1498 (N_1498,In_26,In_913);
nor U1499 (N_1499,In_582,In_435);
nor U1500 (N_1500,In_10,In_669);
or U1501 (N_1501,In_483,In_239);
nor U1502 (N_1502,In_246,In_256);
nor U1503 (N_1503,In_669,In_360);
nor U1504 (N_1504,In_720,In_128);
and U1505 (N_1505,In_507,In_997);
xnor U1506 (N_1506,In_254,In_60);
nor U1507 (N_1507,In_851,In_822);
nor U1508 (N_1508,In_651,In_606);
nand U1509 (N_1509,In_229,In_331);
nand U1510 (N_1510,In_435,In_397);
nor U1511 (N_1511,In_703,In_692);
or U1512 (N_1512,In_30,In_443);
xnor U1513 (N_1513,In_573,In_620);
xnor U1514 (N_1514,In_296,In_987);
or U1515 (N_1515,In_787,In_754);
or U1516 (N_1516,In_746,In_915);
or U1517 (N_1517,In_80,In_437);
xnor U1518 (N_1518,In_398,In_280);
and U1519 (N_1519,In_887,In_325);
nor U1520 (N_1520,In_250,In_749);
nor U1521 (N_1521,In_355,In_671);
xnor U1522 (N_1522,In_152,In_48);
xor U1523 (N_1523,In_369,In_322);
and U1524 (N_1524,In_860,In_718);
and U1525 (N_1525,In_648,In_801);
nand U1526 (N_1526,In_130,In_769);
or U1527 (N_1527,In_902,In_592);
nor U1528 (N_1528,In_380,In_966);
nor U1529 (N_1529,In_562,In_315);
or U1530 (N_1530,In_287,In_324);
nand U1531 (N_1531,In_921,In_452);
and U1532 (N_1532,In_642,In_292);
nand U1533 (N_1533,In_105,In_407);
nand U1534 (N_1534,In_880,In_518);
and U1535 (N_1535,In_682,In_345);
and U1536 (N_1536,In_139,In_854);
or U1537 (N_1537,In_657,In_956);
or U1538 (N_1538,In_520,In_719);
and U1539 (N_1539,In_606,In_375);
nor U1540 (N_1540,In_952,In_107);
nand U1541 (N_1541,In_448,In_290);
nand U1542 (N_1542,In_184,In_724);
xor U1543 (N_1543,In_11,In_219);
and U1544 (N_1544,In_295,In_242);
and U1545 (N_1545,In_785,In_535);
nand U1546 (N_1546,In_505,In_112);
xor U1547 (N_1547,In_261,In_133);
xor U1548 (N_1548,In_558,In_222);
xor U1549 (N_1549,In_659,In_196);
and U1550 (N_1550,In_645,In_554);
xnor U1551 (N_1551,In_360,In_464);
or U1552 (N_1552,In_651,In_760);
nand U1553 (N_1553,In_611,In_282);
or U1554 (N_1554,In_507,In_867);
nor U1555 (N_1555,In_449,In_642);
nor U1556 (N_1556,In_750,In_622);
xor U1557 (N_1557,In_706,In_746);
nor U1558 (N_1558,In_867,In_931);
nand U1559 (N_1559,In_64,In_609);
or U1560 (N_1560,In_913,In_341);
or U1561 (N_1561,In_988,In_543);
nand U1562 (N_1562,In_403,In_795);
nand U1563 (N_1563,In_291,In_187);
nor U1564 (N_1564,In_906,In_767);
nand U1565 (N_1565,In_530,In_997);
and U1566 (N_1566,In_300,In_68);
nor U1567 (N_1567,In_177,In_492);
xor U1568 (N_1568,In_397,In_358);
or U1569 (N_1569,In_672,In_4);
nand U1570 (N_1570,In_590,In_279);
xnor U1571 (N_1571,In_85,In_343);
nor U1572 (N_1572,In_654,In_116);
or U1573 (N_1573,In_324,In_294);
nor U1574 (N_1574,In_366,In_285);
nor U1575 (N_1575,In_671,In_845);
and U1576 (N_1576,In_869,In_121);
and U1577 (N_1577,In_124,In_941);
nand U1578 (N_1578,In_272,In_962);
nand U1579 (N_1579,In_442,In_984);
nand U1580 (N_1580,In_149,In_431);
and U1581 (N_1581,In_61,In_889);
and U1582 (N_1582,In_918,In_841);
and U1583 (N_1583,In_604,In_299);
nand U1584 (N_1584,In_688,In_630);
xor U1585 (N_1585,In_138,In_653);
nand U1586 (N_1586,In_472,In_295);
and U1587 (N_1587,In_918,In_188);
xor U1588 (N_1588,In_330,In_209);
nand U1589 (N_1589,In_273,In_731);
or U1590 (N_1590,In_237,In_577);
or U1591 (N_1591,In_458,In_57);
or U1592 (N_1592,In_6,In_613);
xnor U1593 (N_1593,In_157,In_651);
nor U1594 (N_1594,In_909,In_636);
nand U1595 (N_1595,In_33,In_68);
or U1596 (N_1596,In_45,In_6);
and U1597 (N_1597,In_455,In_258);
nor U1598 (N_1598,In_262,In_207);
nand U1599 (N_1599,In_281,In_721);
xnor U1600 (N_1600,In_17,In_151);
nand U1601 (N_1601,In_870,In_804);
xor U1602 (N_1602,In_372,In_886);
nor U1603 (N_1603,In_969,In_819);
nand U1604 (N_1604,In_896,In_506);
xnor U1605 (N_1605,In_385,In_390);
or U1606 (N_1606,In_962,In_779);
or U1607 (N_1607,In_379,In_826);
nand U1608 (N_1608,In_533,In_821);
or U1609 (N_1609,In_7,In_900);
xor U1610 (N_1610,In_145,In_320);
xor U1611 (N_1611,In_20,In_913);
nor U1612 (N_1612,In_105,In_782);
nor U1613 (N_1613,In_702,In_752);
nand U1614 (N_1614,In_409,In_661);
nand U1615 (N_1615,In_145,In_925);
nand U1616 (N_1616,In_968,In_584);
or U1617 (N_1617,In_854,In_992);
or U1618 (N_1618,In_235,In_405);
or U1619 (N_1619,In_537,In_76);
and U1620 (N_1620,In_552,In_434);
or U1621 (N_1621,In_510,In_661);
xor U1622 (N_1622,In_209,In_849);
xnor U1623 (N_1623,In_2,In_543);
and U1624 (N_1624,In_924,In_971);
xor U1625 (N_1625,In_624,In_750);
nand U1626 (N_1626,In_602,In_664);
nor U1627 (N_1627,In_604,In_478);
nand U1628 (N_1628,In_418,In_185);
nor U1629 (N_1629,In_263,In_185);
and U1630 (N_1630,In_821,In_358);
and U1631 (N_1631,In_723,In_989);
and U1632 (N_1632,In_821,In_733);
nand U1633 (N_1633,In_802,In_740);
nand U1634 (N_1634,In_660,In_723);
nor U1635 (N_1635,In_477,In_716);
nor U1636 (N_1636,In_251,In_966);
xor U1637 (N_1637,In_800,In_945);
nor U1638 (N_1638,In_723,In_396);
xor U1639 (N_1639,In_148,In_740);
or U1640 (N_1640,In_476,In_670);
nor U1641 (N_1641,In_933,In_584);
and U1642 (N_1642,In_425,In_614);
xnor U1643 (N_1643,In_320,In_383);
nor U1644 (N_1644,In_205,In_247);
nor U1645 (N_1645,In_737,In_861);
or U1646 (N_1646,In_783,In_592);
or U1647 (N_1647,In_206,In_525);
nand U1648 (N_1648,In_657,In_350);
or U1649 (N_1649,In_106,In_13);
or U1650 (N_1650,In_18,In_819);
or U1651 (N_1651,In_429,In_964);
xnor U1652 (N_1652,In_696,In_266);
nor U1653 (N_1653,In_200,In_177);
nand U1654 (N_1654,In_917,In_202);
xnor U1655 (N_1655,In_527,In_197);
or U1656 (N_1656,In_986,In_925);
nor U1657 (N_1657,In_824,In_106);
xnor U1658 (N_1658,In_627,In_404);
xor U1659 (N_1659,In_18,In_3);
nand U1660 (N_1660,In_445,In_819);
and U1661 (N_1661,In_47,In_497);
nand U1662 (N_1662,In_195,In_556);
or U1663 (N_1663,In_113,In_266);
nor U1664 (N_1664,In_101,In_255);
nand U1665 (N_1665,In_542,In_660);
and U1666 (N_1666,In_805,In_543);
xnor U1667 (N_1667,In_156,In_145);
or U1668 (N_1668,In_214,In_28);
or U1669 (N_1669,In_105,In_260);
and U1670 (N_1670,In_658,In_246);
nand U1671 (N_1671,In_750,In_484);
or U1672 (N_1672,In_569,In_615);
and U1673 (N_1673,In_756,In_770);
nor U1674 (N_1674,In_122,In_900);
and U1675 (N_1675,In_979,In_935);
nor U1676 (N_1676,In_331,In_467);
or U1677 (N_1677,In_631,In_160);
and U1678 (N_1678,In_93,In_710);
nor U1679 (N_1679,In_942,In_709);
nor U1680 (N_1680,In_29,In_270);
and U1681 (N_1681,In_978,In_998);
nand U1682 (N_1682,In_438,In_920);
and U1683 (N_1683,In_286,In_251);
and U1684 (N_1684,In_527,In_486);
nor U1685 (N_1685,In_596,In_315);
nor U1686 (N_1686,In_106,In_191);
nor U1687 (N_1687,In_188,In_155);
xnor U1688 (N_1688,In_248,In_172);
xor U1689 (N_1689,In_958,In_350);
nor U1690 (N_1690,In_515,In_227);
and U1691 (N_1691,In_539,In_317);
xor U1692 (N_1692,In_498,In_617);
nand U1693 (N_1693,In_400,In_221);
nor U1694 (N_1694,In_904,In_563);
and U1695 (N_1695,In_227,In_633);
nand U1696 (N_1696,In_73,In_547);
nor U1697 (N_1697,In_745,In_232);
or U1698 (N_1698,In_196,In_295);
nor U1699 (N_1699,In_730,In_210);
xor U1700 (N_1700,In_466,In_147);
nor U1701 (N_1701,In_807,In_26);
nor U1702 (N_1702,In_671,In_786);
nor U1703 (N_1703,In_140,In_587);
nand U1704 (N_1704,In_941,In_293);
nand U1705 (N_1705,In_237,In_929);
nor U1706 (N_1706,In_923,In_25);
xnor U1707 (N_1707,In_712,In_819);
nand U1708 (N_1708,In_77,In_102);
or U1709 (N_1709,In_208,In_364);
xnor U1710 (N_1710,In_766,In_688);
and U1711 (N_1711,In_293,In_567);
or U1712 (N_1712,In_227,In_883);
and U1713 (N_1713,In_702,In_365);
xnor U1714 (N_1714,In_292,In_56);
nor U1715 (N_1715,In_445,In_258);
and U1716 (N_1716,In_184,In_294);
and U1717 (N_1717,In_423,In_504);
or U1718 (N_1718,In_827,In_157);
nand U1719 (N_1719,In_877,In_722);
xnor U1720 (N_1720,In_957,In_456);
or U1721 (N_1721,In_384,In_307);
nor U1722 (N_1722,In_789,In_260);
xor U1723 (N_1723,In_781,In_25);
nand U1724 (N_1724,In_214,In_614);
and U1725 (N_1725,In_75,In_161);
and U1726 (N_1726,In_853,In_498);
nand U1727 (N_1727,In_781,In_173);
xor U1728 (N_1728,In_138,In_374);
xnor U1729 (N_1729,In_319,In_185);
nand U1730 (N_1730,In_389,In_376);
and U1731 (N_1731,In_300,In_530);
nand U1732 (N_1732,In_344,In_126);
nand U1733 (N_1733,In_74,In_188);
xor U1734 (N_1734,In_401,In_956);
xnor U1735 (N_1735,In_198,In_545);
nor U1736 (N_1736,In_294,In_877);
nand U1737 (N_1737,In_690,In_895);
and U1738 (N_1738,In_539,In_846);
and U1739 (N_1739,In_341,In_81);
nand U1740 (N_1740,In_487,In_285);
and U1741 (N_1741,In_365,In_510);
or U1742 (N_1742,In_826,In_148);
or U1743 (N_1743,In_456,In_471);
nand U1744 (N_1744,In_994,In_418);
xnor U1745 (N_1745,In_106,In_27);
and U1746 (N_1746,In_505,In_654);
nand U1747 (N_1747,In_899,In_719);
and U1748 (N_1748,In_961,In_660);
or U1749 (N_1749,In_971,In_583);
nor U1750 (N_1750,In_443,In_637);
nand U1751 (N_1751,In_995,In_482);
or U1752 (N_1752,In_777,In_562);
nor U1753 (N_1753,In_772,In_246);
and U1754 (N_1754,In_960,In_996);
or U1755 (N_1755,In_306,In_47);
xor U1756 (N_1756,In_445,In_30);
xnor U1757 (N_1757,In_91,In_821);
xor U1758 (N_1758,In_939,In_820);
or U1759 (N_1759,In_332,In_171);
and U1760 (N_1760,In_31,In_970);
or U1761 (N_1761,In_627,In_786);
nor U1762 (N_1762,In_316,In_732);
and U1763 (N_1763,In_374,In_824);
nand U1764 (N_1764,In_539,In_686);
nor U1765 (N_1765,In_448,In_846);
nand U1766 (N_1766,In_347,In_126);
xor U1767 (N_1767,In_109,In_332);
nor U1768 (N_1768,In_885,In_713);
xor U1769 (N_1769,In_418,In_278);
or U1770 (N_1770,In_859,In_84);
nand U1771 (N_1771,In_457,In_336);
nor U1772 (N_1772,In_72,In_310);
or U1773 (N_1773,In_332,In_683);
and U1774 (N_1774,In_862,In_208);
and U1775 (N_1775,In_660,In_872);
xor U1776 (N_1776,In_425,In_653);
or U1777 (N_1777,In_868,In_291);
or U1778 (N_1778,In_847,In_455);
and U1779 (N_1779,In_665,In_261);
xnor U1780 (N_1780,In_742,In_584);
nor U1781 (N_1781,In_330,In_873);
xnor U1782 (N_1782,In_920,In_382);
or U1783 (N_1783,In_112,In_481);
nor U1784 (N_1784,In_729,In_735);
or U1785 (N_1785,In_938,In_111);
xor U1786 (N_1786,In_16,In_896);
nor U1787 (N_1787,In_193,In_755);
or U1788 (N_1788,In_965,In_45);
and U1789 (N_1789,In_642,In_883);
or U1790 (N_1790,In_527,In_298);
nand U1791 (N_1791,In_45,In_253);
xnor U1792 (N_1792,In_698,In_402);
nand U1793 (N_1793,In_851,In_316);
nand U1794 (N_1794,In_717,In_555);
or U1795 (N_1795,In_491,In_327);
or U1796 (N_1796,In_551,In_376);
nand U1797 (N_1797,In_349,In_227);
and U1798 (N_1798,In_855,In_62);
nor U1799 (N_1799,In_98,In_963);
xnor U1800 (N_1800,In_330,In_114);
or U1801 (N_1801,In_44,In_843);
or U1802 (N_1802,In_502,In_133);
nor U1803 (N_1803,In_656,In_55);
or U1804 (N_1804,In_273,In_782);
xnor U1805 (N_1805,In_708,In_95);
nor U1806 (N_1806,In_95,In_503);
xnor U1807 (N_1807,In_515,In_188);
xor U1808 (N_1808,In_847,In_434);
nand U1809 (N_1809,In_966,In_259);
xnor U1810 (N_1810,In_324,In_450);
and U1811 (N_1811,In_455,In_180);
nand U1812 (N_1812,In_859,In_413);
nand U1813 (N_1813,In_810,In_96);
and U1814 (N_1814,In_374,In_480);
nand U1815 (N_1815,In_746,In_940);
or U1816 (N_1816,In_933,In_703);
xnor U1817 (N_1817,In_445,In_577);
or U1818 (N_1818,In_192,In_382);
xnor U1819 (N_1819,In_863,In_97);
or U1820 (N_1820,In_973,In_730);
or U1821 (N_1821,In_273,In_688);
nor U1822 (N_1822,In_268,In_893);
or U1823 (N_1823,In_120,In_71);
nand U1824 (N_1824,In_587,In_697);
xnor U1825 (N_1825,In_312,In_567);
nand U1826 (N_1826,In_321,In_52);
nand U1827 (N_1827,In_211,In_824);
nor U1828 (N_1828,In_419,In_812);
and U1829 (N_1829,In_189,In_79);
and U1830 (N_1830,In_949,In_960);
and U1831 (N_1831,In_759,In_663);
or U1832 (N_1832,In_242,In_938);
and U1833 (N_1833,In_688,In_266);
and U1834 (N_1834,In_161,In_446);
nor U1835 (N_1835,In_188,In_85);
nand U1836 (N_1836,In_276,In_986);
xnor U1837 (N_1837,In_2,In_730);
xor U1838 (N_1838,In_683,In_204);
nor U1839 (N_1839,In_680,In_973);
or U1840 (N_1840,In_854,In_455);
or U1841 (N_1841,In_990,In_27);
or U1842 (N_1842,In_420,In_583);
or U1843 (N_1843,In_298,In_211);
or U1844 (N_1844,In_751,In_371);
or U1845 (N_1845,In_14,In_235);
and U1846 (N_1846,In_851,In_104);
nand U1847 (N_1847,In_950,In_544);
and U1848 (N_1848,In_266,In_494);
or U1849 (N_1849,In_246,In_102);
nor U1850 (N_1850,In_368,In_405);
nand U1851 (N_1851,In_406,In_901);
and U1852 (N_1852,In_424,In_645);
and U1853 (N_1853,In_280,In_198);
xor U1854 (N_1854,In_653,In_473);
nand U1855 (N_1855,In_864,In_826);
nor U1856 (N_1856,In_306,In_428);
nand U1857 (N_1857,In_769,In_442);
nand U1858 (N_1858,In_6,In_851);
or U1859 (N_1859,In_808,In_92);
nand U1860 (N_1860,In_966,In_686);
nand U1861 (N_1861,In_641,In_158);
xor U1862 (N_1862,In_578,In_431);
xnor U1863 (N_1863,In_271,In_532);
nor U1864 (N_1864,In_16,In_137);
and U1865 (N_1865,In_885,In_273);
nand U1866 (N_1866,In_695,In_606);
nor U1867 (N_1867,In_569,In_446);
nor U1868 (N_1868,In_609,In_578);
xnor U1869 (N_1869,In_660,In_264);
nand U1870 (N_1870,In_225,In_902);
nand U1871 (N_1871,In_916,In_280);
and U1872 (N_1872,In_379,In_549);
or U1873 (N_1873,In_217,In_170);
xor U1874 (N_1874,In_848,In_861);
and U1875 (N_1875,In_74,In_760);
or U1876 (N_1876,In_426,In_246);
nor U1877 (N_1877,In_687,In_394);
or U1878 (N_1878,In_863,In_988);
xnor U1879 (N_1879,In_226,In_703);
nand U1880 (N_1880,In_714,In_343);
or U1881 (N_1881,In_398,In_296);
and U1882 (N_1882,In_131,In_518);
xnor U1883 (N_1883,In_899,In_186);
nand U1884 (N_1884,In_392,In_753);
nor U1885 (N_1885,In_872,In_760);
nand U1886 (N_1886,In_644,In_908);
and U1887 (N_1887,In_992,In_656);
nor U1888 (N_1888,In_730,In_111);
nand U1889 (N_1889,In_801,In_723);
or U1890 (N_1890,In_773,In_330);
xor U1891 (N_1891,In_103,In_467);
nor U1892 (N_1892,In_910,In_189);
nor U1893 (N_1893,In_622,In_821);
and U1894 (N_1894,In_365,In_69);
nor U1895 (N_1895,In_281,In_247);
nand U1896 (N_1896,In_295,In_881);
and U1897 (N_1897,In_880,In_423);
nand U1898 (N_1898,In_393,In_543);
and U1899 (N_1899,In_557,In_854);
or U1900 (N_1900,In_243,In_118);
nand U1901 (N_1901,In_985,In_274);
or U1902 (N_1902,In_639,In_680);
or U1903 (N_1903,In_489,In_102);
nand U1904 (N_1904,In_282,In_741);
or U1905 (N_1905,In_578,In_32);
and U1906 (N_1906,In_212,In_439);
nor U1907 (N_1907,In_828,In_208);
nor U1908 (N_1908,In_767,In_537);
xor U1909 (N_1909,In_905,In_731);
nor U1910 (N_1910,In_120,In_240);
xor U1911 (N_1911,In_672,In_695);
nor U1912 (N_1912,In_349,In_230);
xnor U1913 (N_1913,In_417,In_643);
xnor U1914 (N_1914,In_42,In_917);
xnor U1915 (N_1915,In_873,In_427);
or U1916 (N_1916,In_634,In_881);
and U1917 (N_1917,In_438,In_267);
nor U1918 (N_1918,In_548,In_90);
and U1919 (N_1919,In_854,In_738);
or U1920 (N_1920,In_626,In_652);
and U1921 (N_1921,In_29,In_93);
nand U1922 (N_1922,In_878,In_586);
and U1923 (N_1923,In_790,In_117);
nor U1924 (N_1924,In_889,In_851);
or U1925 (N_1925,In_640,In_981);
and U1926 (N_1926,In_312,In_746);
and U1927 (N_1927,In_984,In_629);
or U1928 (N_1928,In_642,In_62);
xor U1929 (N_1929,In_987,In_189);
nor U1930 (N_1930,In_343,In_491);
nor U1931 (N_1931,In_892,In_466);
xnor U1932 (N_1932,In_118,In_534);
or U1933 (N_1933,In_268,In_155);
nand U1934 (N_1934,In_808,In_530);
or U1935 (N_1935,In_438,In_444);
nor U1936 (N_1936,In_289,In_224);
nor U1937 (N_1937,In_788,In_305);
and U1938 (N_1938,In_380,In_115);
or U1939 (N_1939,In_199,In_483);
xnor U1940 (N_1940,In_516,In_72);
or U1941 (N_1941,In_289,In_236);
or U1942 (N_1942,In_285,In_916);
and U1943 (N_1943,In_394,In_440);
nor U1944 (N_1944,In_471,In_923);
nor U1945 (N_1945,In_484,In_574);
xnor U1946 (N_1946,In_772,In_165);
nand U1947 (N_1947,In_656,In_466);
xnor U1948 (N_1948,In_406,In_83);
and U1949 (N_1949,In_883,In_690);
and U1950 (N_1950,In_167,In_808);
or U1951 (N_1951,In_659,In_678);
or U1952 (N_1952,In_662,In_840);
nand U1953 (N_1953,In_760,In_661);
xor U1954 (N_1954,In_360,In_184);
and U1955 (N_1955,In_630,In_174);
or U1956 (N_1956,In_241,In_801);
nand U1957 (N_1957,In_845,In_523);
xnor U1958 (N_1958,In_733,In_831);
xor U1959 (N_1959,In_842,In_439);
xor U1960 (N_1960,In_41,In_542);
nor U1961 (N_1961,In_27,In_49);
and U1962 (N_1962,In_559,In_805);
nand U1963 (N_1963,In_415,In_371);
nor U1964 (N_1964,In_180,In_130);
nand U1965 (N_1965,In_31,In_294);
nand U1966 (N_1966,In_202,In_795);
or U1967 (N_1967,In_901,In_668);
nor U1968 (N_1968,In_529,In_475);
nor U1969 (N_1969,In_523,In_321);
and U1970 (N_1970,In_223,In_53);
nand U1971 (N_1971,In_645,In_707);
and U1972 (N_1972,In_520,In_280);
nor U1973 (N_1973,In_615,In_915);
nor U1974 (N_1974,In_428,In_57);
nand U1975 (N_1975,In_601,In_589);
nand U1976 (N_1976,In_843,In_624);
and U1977 (N_1977,In_884,In_45);
xnor U1978 (N_1978,In_6,In_789);
and U1979 (N_1979,In_303,In_38);
and U1980 (N_1980,In_432,In_346);
or U1981 (N_1981,In_401,In_979);
xnor U1982 (N_1982,In_270,In_749);
nand U1983 (N_1983,In_413,In_353);
nor U1984 (N_1984,In_126,In_377);
and U1985 (N_1985,In_439,In_942);
or U1986 (N_1986,In_247,In_897);
nand U1987 (N_1987,In_994,In_703);
xor U1988 (N_1988,In_948,In_719);
or U1989 (N_1989,In_476,In_941);
xor U1990 (N_1990,In_141,In_795);
or U1991 (N_1991,In_354,In_415);
nor U1992 (N_1992,In_674,In_650);
nand U1993 (N_1993,In_732,In_271);
or U1994 (N_1994,In_144,In_4);
xor U1995 (N_1995,In_515,In_78);
nand U1996 (N_1996,In_899,In_570);
and U1997 (N_1997,In_568,In_664);
nand U1998 (N_1998,In_591,In_458);
or U1999 (N_1999,In_880,In_693);
nand U2000 (N_2000,N_1723,N_1215);
nor U2001 (N_2001,N_1677,N_345);
nand U2002 (N_2002,N_711,N_31);
xor U2003 (N_2003,N_503,N_1347);
xnor U2004 (N_2004,N_626,N_212);
nand U2005 (N_2005,N_397,N_1120);
or U2006 (N_2006,N_1407,N_1065);
nor U2007 (N_2007,N_1443,N_587);
xor U2008 (N_2008,N_1115,N_260);
nand U2009 (N_2009,N_716,N_1283);
or U2010 (N_2010,N_771,N_1359);
or U2011 (N_2011,N_1782,N_285);
nand U2012 (N_2012,N_1094,N_1924);
nand U2013 (N_2013,N_1531,N_1621);
xor U2014 (N_2014,N_1456,N_960);
nor U2015 (N_2015,N_532,N_250);
xor U2016 (N_2016,N_1327,N_1976);
nor U2017 (N_2017,N_1282,N_1229);
nor U2018 (N_2018,N_1995,N_986);
xor U2019 (N_2019,N_1756,N_1616);
or U2020 (N_2020,N_1653,N_976);
xnor U2021 (N_2021,N_984,N_978);
nand U2022 (N_2022,N_147,N_1838);
xnor U2023 (N_2023,N_1242,N_1608);
and U2024 (N_2024,N_1295,N_735);
nand U2025 (N_2025,N_144,N_1592);
nand U2026 (N_2026,N_138,N_574);
xnor U2027 (N_2027,N_604,N_1418);
nor U2028 (N_2028,N_1564,N_766);
and U2029 (N_2029,N_371,N_824);
nand U2030 (N_2030,N_1854,N_21);
xor U2031 (N_2031,N_996,N_394);
or U2032 (N_2032,N_183,N_554);
or U2033 (N_2033,N_615,N_846);
nor U2034 (N_2034,N_1644,N_1364);
or U2035 (N_2035,N_1532,N_1139);
nor U2036 (N_2036,N_1469,N_1461);
or U2037 (N_2037,N_1222,N_1167);
nand U2038 (N_2038,N_1866,N_608);
and U2039 (N_2039,N_1553,N_1472);
nor U2040 (N_2040,N_1414,N_1107);
and U2041 (N_2041,N_569,N_498);
xnor U2042 (N_2042,N_1983,N_1780);
or U2043 (N_2043,N_1864,N_733);
and U2044 (N_2044,N_1547,N_651);
xnor U2045 (N_2045,N_1626,N_1596);
and U2046 (N_2046,N_1758,N_1422);
and U2047 (N_2047,N_1615,N_1966);
and U2048 (N_2048,N_769,N_1234);
nand U2049 (N_2049,N_507,N_92);
or U2050 (N_2050,N_1795,N_1668);
xnor U2051 (N_2051,N_642,N_232);
or U2052 (N_2052,N_1829,N_848);
or U2053 (N_2053,N_1951,N_449);
nor U2054 (N_2054,N_739,N_1606);
xnor U2055 (N_2055,N_188,N_1190);
xnor U2056 (N_2056,N_1991,N_1240);
nor U2057 (N_2057,N_481,N_1509);
nor U2058 (N_2058,N_415,N_886);
or U2059 (N_2059,N_1238,N_1427);
or U2060 (N_2060,N_1146,N_827);
and U2061 (N_2061,N_513,N_737);
and U2062 (N_2062,N_1058,N_1535);
nor U2063 (N_2063,N_516,N_68);
and U2064 (N_2064,N_1464,N_1661);
or U2065 (N_2065,N_77,N_1145);
nor U2066 (N_2066,N_1467,N_145);
nor U2067 (N_2067,N_1105,N_1322);
and U2068 (N_2068,N_1377,N_1800);
nand U2069 (N_2069,N_688,N_1223);
nand U2070 (N_2070,N_1882,N_81);
or U2071 (N_2071,N_1049,N_1702);
or U2072 (N_2072,N_849,N_1417);
and U2073 (N_2073,N_57,N_381);
or U2074 (N_2074,N_1940,N_1557);
and U2075 (N_2075,N_946,N_1008);
nor U2076 (N_2076,N_814,N_152);
xor U2077 (N_2077,N_1281,N_1013);
nor U2078 (N_2078,N_1595,N_672);
nor U2079 (N_2079,N_1929,N_1409);
nor U2080 (N_2080,N_1163,N_1586);
or U2081 (N_2081,N_1818,N_1540);
nor U2082 (N_2082,N_1019,N_1286);
or U2083 (N_2083,N_116,N_1368);
and U2084 (N_2084,N_247,N_197);
and U2085 (N_2085,N_139,N_957);
nand U2086 (N_2086,N_1772,N_23);
or U2087 (N_2087,N_1266,N_1278);
and U2088 (N_2088,N_550,N_1884);
nand U2089 (N_2089,N_885,N_1620);
or U2090 (N_2090,N_15,N_895);
nor U2091 (N_2091,N_476,N_231);
and U2092 (N_2092,N_246,N_1518);
nor U2093 (N_2093,N_515,N_326);
and U2094 (N_2094,N_1219,N_162);
and U2095 (N_2095,N_1545,N_1381);
nor U2096 (N_2096,N_202,N_531);
or U2097 (N_2097,N_8,N_359);
nor U2098 (N_2098,N_1396,N_1771);
xnor U2099 (N_2099,N_88,N_971);
and U2100 (N_2100,N_1397,N_5);
or U2101 (N_2101,N_56,N_1906);
xnor U2102 (N_2102,N_1089,N_338);
nor U2103 (N_2103,N_1994,N_1346);
nand U2104 (N_2104,N_434,N_683);
or U2105 (N_2105,N_485,N_668);
nor U2106 (N_2106,N_82,N_664);
xnor U2107 (N_2107,N_395,N_727);
xnor U2108 (N_2108,N_1707,N_977);
or U2109 (N_2109,N_795,N_640);
nor U2110 (N_2110,N_75,N_703);
and U2111 (N_2111,N_883,N_952);
or U2112 (N_2112,N_1257,N_210);
nand U2113 (N_2113,N_19,N_256);
or U2114 (N_2114,N_1842,N_1949);
and U2115 (N_2115,N_1999,N_951);
or U2116 (N_2116,N_621,N_1431);
xor U2117 (N_2117,N_176,N_1872);
and U2118 (N_2118,N_1528,N_189);
nand U2119 (N_2119,N_204,N_1189);
nor U2120 (N_2120,N_979,N_455);
nand U2121 (N_2121,N_1850,N_844);
xnor U2122 (N_2122,N_709,N_288);
or U2123 (N_2123,N_1688,N_362);
and U2124 (N_2124,N_900,N_251);
nand U2125 (N_2125,N_1142,N_837);
nor U2126 (N_2126,N_266,N_165);
nand U2127 (N_2127,N_760,N_489);
or U2128 (N_2128,N_500,N_659);
nor U2129 (N_2129,N_612,N_881);
or U2130 (N_2130,N_1114,N_1293);
or U2131 (N_2131,N_514,N_872);
xnor U2132 (N_2132,N_1767,N_859);
nor U2133 (N_2133,N_323,N_1098);
nor U2134 (N_2134,N_573,N_106);
nand U2135 (N_2135,N_1869,N_599);
or U2136 (N_2136,N_1127,N_1053);
and U2137 (N_2137,N_1235,N_815);
nor U2138 (N_2138,N_1815,N_1965);
and U2139 (N_2139,N_1077,N_1710);
and U2140 (N_2140,N_776,N_1214);
nand U2141 (N_2141,N_1916,N_1218);
or U2142 (N_2142,N_25,N_1319);
nor U2143 (N_2143,N_29,N_1311);
and U2144 (N_2144,N_322,N_566);
nand U2145 (N_2145,N_1665,N_861);
xor U2146 (N_2146,N_1640,N_1154);
nand U2147 (N_2147,N_80,N_217);
nand U2148 (N_2148,N_1173,N_1663);
xor U2149 (N_2149,N_765,N_959);
nand U2150 (N_2150,N_1100,N_1224);
and U2151 (N_2151,N_400,N_1759);
nor U2152 (N_2152,N_72,N_1880);
nor U2153 (N_2153,N_1982,N_619);
nor U2154 (N_2154,N_1434,N_1268);
nor U2155 (N_2155,N_101,N_1591);
and U2156 (N_2156,N_836,N_1205);
nor U2157 (N_2157,N_1790,N_829);
nand U2158 (N_2158,N_1534,N_517);
nand U2159 (N_2159,N_882,N_1079);
nand U2160 (N_2160,N_274,N_1097);
xor U2161 (N_2161,N_1122,N_1367);
nor U2162 (N_2162,N_843,N_1111);
xor U2163 (N_2163,N_834,N_1221);
nor U2164 (N_2164,N_333,N_511);
or U2165 (N_2165,N_54,N_693);
and U2166 (N_2166,N_756,N_598);
nand U2167 (N_2167,N_1910,N_1216);
nand U2168 (N_2168,N_389,N_32);
or U2169 (N_2169,N_463,N_170);
nor U2170 (N_2170,N_1743,N_1823);
xor U2171 (N_2171,N_1303,N_732);
and U2172 (N_2172,N_1104,N_1739);
or U2173 (N_2173,N_1188,N_1898);
nand U2174 (N_2174,N_1753,N_304);
nor U2175 (N_2175,N_1550,N_105);
or U2176 (N_2176,N_1323,N_537);
nor U2177 (N_2177,N_893,N_789);
xor U2178 (N_2178,N_99,N_412);
and U2179 (N_2179,N_891,N_1162);
and U2180 (N_2180,N_1061,N_956);
and U2181 (N_2181,N_67,N_751);
and U2182 (N_2182,N_1404,N_1953);
xor U2183 (N_2183,N_1783,N_1131);
nand U2184 (N_2184,N_1348,N_108);
nor U2185 (N_2185,N_613,N_1475);
nand U2186 (N_2186,N_527,N_1984);
xor U2187 (N_2187,N_665,N_1284);
nor U2188 (N_2188,N_1370,N_1204);
and U2189 (N_2189,N_1683,N_1070);
nor U2190 (N_2190,N_1119,N_1042);
nor U2191 (N_2191,N_1371,N_1958);
xnor U2192 (N_2192,N_1876,N_1671);
and U2193 (N_2193,N_953,N_1987);
nor U2194 (N_2194,N_1751,N_264);
nand U2195 (N_2195,N_1117,N_1393);
xor U2196 (N_2196,N_1867,N_282);
or U2197 (N_2197,N_966,N_968);
or U2198 (N_2198,N_1044,N_1598);
nand U2199 (N_2199,N_1401,N_1352);
or U2200 (N_2200,N_1629,N_1438);
and U2201 (N_2201,N_1667,N_945);
nand U2202 (N_2202,N_821,N_1571);
xnor U2203 (N_2203,N_435,N_617);
xor U2204 (N_2204,N_1436,N_1811);
and U2205 (N_2205,N_1091,N_261);
or U2206 (N_2206,N_1263,N_244);
nand U2207 (N_2207,N_1384,N_1847);
or U2208 (N_2208,N_559,N_1600);
xnor U2209 (N_2209,N_1833,N_563);
xor U2210 (N_2210,N_923,N_832);
and U2211 (N_2211,N_1118,N_850);
or U2212 (N_2212,N_905,N_257);
nand U2213 (N_2213,N_191,N_319);
and U2214 (N_2214,N_1925,N_1904);
and U2215 (N_2215,N_1195,N_1985);
or U2216 (N_2216,N_199,N_925);
or U2217 (N_2217,N_1330,N_1428);
xnor U2218 (N_2218,N_487,N_896);
or U2219 (N_2219,N_444,N_1186);
xnor U2220 (N_2220,N_1307,N_1279);
nor U2221 (N_2221,N_1481,N_548);
nor U2222 (N_2222,N_1074,N_1781);
xor U2223 (N_2223,N_1064,N_1354);
or U2224 (N_2224,N_787,N_792);
or U2225 (N_2225,N_207,N_1237);
nor U2226 (N_2226,N_1010,N_1959);
nor U2227 (N_2227,N_512,N_1918);
and U2228 (N_2228,N_989,N_1236);
nand U2229 (N_2229,N_480,N_186);
and U2230 (N_2230,N_1580,N_1106);
nor U2231 (N_2231,N_1516,N_393);
xor U2232 (N_2232,N_1349,N_1478);
nand U2233 (N_2233,N_1172,N_1124);
nand U2234 (N_2234,N_680,N_590);
and U2235 (N_2235,N_94,N_1932);
xor U2236 (N_2236,N_1792,N_1726);
or U2237 (N_2237,N_662,N_1968);
xor U2238 (N_2238,N_293,N_1433);
nand U2239 (N_2239,N_1298,N_1155);
xnor U2240 (N_2240,N_1344,N_851);
and U2241 (N_2241,N_375,N_1619);
nor U2242 (N_2242,N_666,N_1669);
xor U2243 (N_2243,N_761,N_911);
or U2244 (N_2244,N_1684,N_1423);
xnor U2245 (N_2245,N_3,N_858);
xor U2246 (N_2246,N_1652,N_459);
xor U2247 (N_2247,N_343,N_1902);
and U2248 (N_2248,N_234,N_1259);
xor U2249 (N_2249,N_215,N_483);
nand U2250 (N_2250,N_1389,N_1868);
and U2251 (N_2251,N_682,N_1177);
xnor U2252 (N_2252,N_320,N_1921);
xor U2253 (N_2253,N_1225,N_519);
and U2254 (N_2254,N_1241,N_1757);
nor U2255 (N_2255,N_1329,N_1841);
and U2256 (N_2256,N_1416,N_1583);
and U2257 (N_2257,N_562,N_864);
or U2258 (N_2258,N_628,N_1861);
and U2259 (N_2259,N_700,N_1442);
nand U2260 (N_2260,N_991,N_630);
or U2261 (N_2261,N_892,N_830);
or U2262 (N_2262,N_1696,N_1007);
nor U2263 (N_2263,N_1562,N_213);
or U2264 (N_2264,N_639,N_114);
xor U2265 (N_2265,N_692,N_115);
xnor U2266 (N_2266,N_706,N_1769);
xor U2267 (N_2267,N_1400,N_1803);
nand U2268 (N_2268,N_280,N_539);
and U2269 (N_2269,N_1623,N_522);
or U2270 (N_2270,N_1137,N_647);
nand U2271 (N_2271,N_930,N_271);
nand U2272 (N_2272,N_904,N_1067);
or U2273 (N_2273,N_79,N_391);
xnor U2274 (N_2274,N_744,N_1128);
xor U2275 (N_2275,N_658,N_1836);
nand U2276 (N_2276,N_1862,N_1379);
or U2277 (N_2277,N_1785,N_1316);
or U2278 (N_2278,N_1385,N_1479);
nand U2279 (N_2279,N_1102,N_360);
and U2280 (N_2280,N_1365,N_1650);
nand U2281 (N_2281,N_1280,N_710);
nand U2282 (N_2282,N_1140,N_1825);
nand U2283 (N_2283,N_90,N_1402);
xor U2284 (N_2284,N_1037,N_1088);
nor U2285 (N_2285,N_652,N_1308);
nor U2286 (N_2286,N_1814,N_113);
nor U2287 (N_2287,N_1915,N_1713);
and U2288 (N_2288,N_73,N_1301);
xor U2289 (N_2289,N_646,N_1946);
or U2290 (N_2290,N_425,N_1063);
and U2291 (N_2291,N_1943,N_799);
nor U2292 (N_2292,N_1476,N_1788);
or U2293 (N_2293,N_134,N_1444);
and U2294 (N_2294,N_1967,N_158);
xor U2295 (N_2295,N_812,N_1527);
or U2296 (N_2296,N_1605,N_629);
nand U2297 (N_2297,N_1181,N_1043);
nor U2298 (N_2298,N_942,N_89);
and U2299 (N_2299,N_985,N_1326);
nand U2300 (N_2300,N_1599,N_1699);
nor U2301 (N_2301,N_1666,N_1273);
or U2302 (N_2302,N_436,N_1116);
nor U2303 (N_2303,N_1143,N_1858);
nand U2304 (N_2304,N_913,N_964);
nor U2305 (N_2305,N_635,N_1016);
and U2306 (N_2306,N_1253,N_417);
and U2307 (N_2307,N_277,N_720);
and U2308 (N_2308,N_1636,N_1733);
nor U2309 (N_2309,N_1911,N_356);
nand U2310 (N_2310,N_185,N_774);
and U2311 (N_2311,N_1152,N_1210);
nand U2312 (N_2312,N_1700,N_1731);
xnor U2313 (N_2313,N_332,N_482);
nand U2314 (N_2314,N_867,N_1863);
nor U2315 (N_2315,N_722,N_564);
and U2316 (N_2316,N_967,N_1536);
nand U2317 (N_2317,N_30,N_875);
or U2318 (N_2318,N_1170,N_376);
or U2319 (N_2319,N_1698,N_494);
nor U2320 (N_2320,N_778,N_1108);
xor U2321 (N_2321,N_1813,N_1579);
nand U2322 (N_2322,N_1093,N_1763);
or U2323 (N_2323,N_1530,N_263);
nor U2324 (N_2324,N_1694,N_1617);
or U2325 (N_2325,N_508,N_1185);
nand U2326 (N_2326,N_1541,N_386);
nand U2327 (N_2327,N_1986,N_1310);
nor U2328 (N_2328,N_1738,N_1337);
or U2329 (N_2329,N_130,N_346);
nand U2330 (N_2330,N_794,N_506);
xor U2331 (N_2331,N_173,N_1200);
or U2332 (N_2332,N_785,N_216);
and U2333 (N_2333,N_768,N_1026);
and U2334 (N_2334,N_51,N_818);
or U2335 (N_2335,N_337,N_1069);
nand U2336 (N_2336,N_718,N_616);
or U2337 (N_2337,N_603,N_61);
nand U2338 (N_2338,N_1048,N_1632);
nor U2339 (N_2339,N_1761,N_678);
and U2340 (N_2340,N_762,N_715);
xnor U2341 (N_2341,N_1522,N_353);
xnor U2342 (N_2342,N_1657,N_705);
nand U2343 (N_2343,N_1908,N_1597);
or U2344 (N_2344,N_650,N_1339);
xnor U2345 (N_2345,N_473,N_1046);
nor U2346 (N_2346,N_1740,N_1486);
nor U2347 (N_2347,N_198,N_1470);
nand U2348 (N_2348,N_1488,N_1055);
and U2349 (N_2349,N_1821,N_748);
and U2350 (N_2350,N_312,N_1826);
and U2351 (N_2351,N_97,N_1161);
xnor U2352 (N_2352,N_1913,N_177);
xnor U2353 (N_2353,N_262,N_1820);
nor U2354 (N_2354,N_1960,N_1554);
and U2355 (N_2355,N_783,N_1618);
nor U2356 (N_2356,N_20,N_1299);
nand U2357 (N_2357,N_1395,N_384);
nand U2358 (N_2358,N_679,N_63);
or U2359 (N_2359,N_1141,N_1747);
and U2360 (N_2360,N_1449,N_1670);
xnor U2361 (N_2361,N_888,N_754);
nand U2362 (N_2362,N_746,N_270);
nor U2363 (N_2363,N_845,N_1012);
nand U2364 (N_2364,N_1483,N_728);
or U2365 (N_2365,N_249,N_567);
xnor U2366 (N_2366,N_1972,N_477);
or U2367 (N_2367,N_1935,N_1148);
nor U2368 (N_2368,N_59,N_396);
and U2369 (N_2369,N_348,N_1062);
nand U2370 (N_2370,N_1712,N_1080);
or U2371 (N_2371,N_1745,N_214);
or U2372 (N_2372,N_65,N_802);
and U2373 (N_2373,N_973,N_518);
nand U2374 (N_2374,N_758,N_767);
and U2375 (N_2375,N_1722,N_1865);
or U2376 (N_2376,N_1926,N_935);
xnor U2377 (N_2377,N_1555,N_1584);
nand U2378 (N_2378,N_1812,N_1027);
xor U2379 (N_2379,N_1799,N_1403);
nand U2380 (N_2380,N_1315,N_1827);
xor U2381 (N_2381,N_1388,N_1581);
nand U2382 (N_2382,N_690,N_1998);
nor U2383 (N_2383,N_1228,N_1432);
or U2384 (N_2384,N_790,N_1052);
nor U2385 (N_2385,N_600,N_934);
nor U2386 (N_2386,N_431,N_1643);
or U2387 (N_2387,N_1614,N_1627);
xor U2388 (N_2388,N_1593,N_299);
xor U2389 (N_2389,N_1970,N_602);
nand U2390 (N_2390,N_1511,N_1568);
nor U2391 (N_2391,N_1230,N_1659);
xnor U2392 (N_2392,N_1538,N_331);
nor U2393 (N_2393,N_1828,N_685);
xnor U2394 (N_2394,N_1804,N_1355);
xnor U2395 (N_2395,N_865,N_404);
nor U2396 (N_2396,N_1260,N_451);
and U2397 (N_2397,N_1888,N_644);
xor U2398 (N_2398,N_1543,N_643);
nand U2399 (N_2399,N_41,N_909);
nor U2400 (N_2400,N_993,N_579);
xnor U2401 (N_2401,N_970,N_1086);
nor U2402 (N_2402,N_1500,N_912);
or U2403 (N_2403,N_297,N_458);
and U2404 (N_2404,N_142,N_281);
or U2405 (N_2405,N_1363,N_857);
xnor U2406 (N_2406,N_529,N_1891);
nand U2407 (N_2407,N_126,N_982);
nor U2408 (N_2408,N_770,N_1822);
or U2409 (N_2409,N_1539,N_920);
xor U2410 (N_2410,N_11,N_1497);
nor U2411 (N_2411,N_9,N_536);
nand U2412 (N_2412,N_520,N_1879);
or U2413 (N_2413,N_910,N_466);
and U2414 (N_2414,N_943,N_364);
xnor U2415 (N_2415,N_995,N_929);
or U2416 (N_2416,N_580,N_1957);
nor U2417 (N_2417,N_1025,N_190);
nor U2418 (N_2418,N_1660,N_314);
nor U2419 (N_2419,N_1424,N_1682);
or U2420 (N_2420,N_1937,N_622);
and U2421 (N_2421,N_205,N_1981);
or U2422 (N_2422,N_1437,N_479);
or U2423 (N_2423,N_1135,N_318);
or U2424 (N_2424,N_804,N_38);
nand U2425 (N_2425,N_474,N_1252);
nand U2426 (N_2426,N_149,N_491);
nor U2427 (N_2427,N_545,N_443);
and U2428 (N_2428,N_437,N_1594);
or U2429 (N_2429,N_1714,N_1033);
xnor U2430 (N_2430,N_983,N_1749);
and U2431 (N_2431,N_1578,N_1351);
or U2432 (N_2432,N_1770,N_187);
nand U2433 (N_2433,N_416,N_120);
xor U2434 (N_2434,N_161,N_1291);
and U2435 (N_2435,N_1206,N_488);
nand U2436 (N_2436,N_1523,N_307);
nor U2437 (N_2437,N_847,N_1830);
nand U2438 (N_2438,N_1466,N_1947);
or U2439 (N_2439,N_660,N_606);
nand U2440 (N_2440,N_1732,N_691);
or U2441 (N_2441,N_334,N_1729);
xor U2442 (N_2442,N_1474,N_842);
xnor U2443 (N_2443,N_1798,N_44);
nor U2444 (N_2444,N_245,N_26);
nand U2445 (N_2445,N_1011,N_136);
or U2446 (N_2446,N_505,N_1290);
xor U2447 (N_2447,N_1076,N_366);
xnor U2448 (N_2448,N_889,N_914);
or U2449 (N_2449,N_184,N_310);
or U2450 (N_2450,N_1101,N_1881);
xnor U2451 (N_2451,N_296,N_424);
or U2452 (N_2452,N_83,N_1589);
and U2453 (N_2453,N_1569,N_1680);
and U2454 (N_2454,N_833,N_1328);
nand U2455 (N_2455,N_69,N_571);
and U2456 (N_2456,N_538,N_325);
nor U2457 (N_2457,N_267,N_1917);
nor U2458 (N_2458,N_713,N_1159);
xnor U2459 (N_2459,N_556,N_1103);
nor U2460 (N_2460,N_1174,N_1171);
and U2461 (N_2461,N_440,N_524);
nor U2462 (N_2462,N_1369,N_1649);
or U2463 (N_2463,N_1576,N_676);
and U2464 (N_2464,N_962,N_1964);
xnor U2465 (N_2465,N_1247,N_290);
and U2466 (N_2466,N_753,N_209);
and U2467 (N_2467,N_95,N_1398);
nand U2468 (N_2468,N_1572,N_194);
nor U2469 (N_2469,N_1718,N_454);
and U2470 (N_2470,N_122,N_1524);
or U2471 (N_2471,N_997,N_1233);
or U2472 (N_2472,N_269,N_645);
or U2473 (N_2473,N_551,N_49);
xnor U2474 (N_2474,N_1824,N_7);
or U2475 (N_2475,N_582,N_1877);
and U2476 (N_2476,N_1460,N_430);
and U2477 (N_2477,N_357,N_46);
xnor U2478 (N_2478,N_1501,N_620);
nor U2479 (N_2479,N_388,N_1207);
xnor U2480 (N_2480,N_641,N_1232);
or U2481 (N_2481,N_530,N_798);
nor U2482 (N_2482,N_1493,N_862);
xor U2483 (N_2483,N_408,N_329);
nor U2484 (N_2484,N_1386,N_648);
xnor U2485 (N_2485,N_1948,N_241);
nor U2486 (N_2486,N_558,N_1387);
xnor U2487 (N_2487,N_379,N_510);
and U2488 (N_2488,N_1256,N_390);
nor U2489 (N_2489,N_1023,N_368);
xnor U2490 (N_2490,N_1341,N_1945);
and U2491 (N_2491,N_933,N_1848);
xor U2492 (N_2492,N_1192,N_1036);
nor U2493 (N_2493,N_475,N_866);
or U2494 (N_2494,N_907,N_526);
or U2495 (N_2495,N_70,N_696);
nand U2496 (N_2496,N_1262,N_961);
xor U2497 (N_2497,N_610,N_1860);
xnor U2498 (N_2498,N_1647,N_1936);
nor U2499 (N_2499,N_433,N_819);
nand U2500 (N_2500,N_1655,N_66);
nand U2501 (N_2501,N_221,N_697);
xnor U2502 (N_2502,N_614,N_1575);
xor U2503 (N_2503,N_1519,N_1897);
or U2504 (N_2504,N_1907,N_1040);
or U2505 (N_2505,N_1988,N_1574);
nand U2506 (N_2506,N_839,N_1941);
and U2507 (N_2507,N_156,N_140);
nand U2508 (N_2508,N_726,N_1243);
xnor U2509 (N_2509,N_764,N_1704);
xor U2510 (N_2510,N_1017,N_1944);
or U2511 (N_2511,N_632,N_1664);
nand U2512 (N_2512,N_1021,N_738);
xnor U2513 (N_2513,N_649,N_1213);
nor U2514 (N_2514,N_86,N_980);
or U2515 (N_2515,N_53,N_1508);
nor U2516 (N_2516,N_1565,N_465);
xor U2517 (N_2517,N_940,N_1577);
and U2518 (N_2518,N_1166,N_887);
nor U2519 (N_2519,N_1582,N_1809);
xnor U2520 (N_2520,N_1727,N_1275);
nand U2521 (N_2521,N_171,N_695);
xor U2522 (N_2522,N_1198,N_34);
nand U2523 (N_2523,N_655,N_759);
and U2524 (N_2524,N_1646,N_111);
nand U2525 (N_2525,N_1755,N_1885);
and U2526 (N_2526,N_560,N_181);
nand U2527 (N_2527,N_1933,N_1005);
and U2528 (N_2528,N_1954,N_1276);
nand U2529 (N_2529,N_1413,N_1612);
nand U2530 (N_2530,N_219,N_1246);
and U2531 (N_2531,N_240,N_823);
xor U2532 (N_2532,N_1975,N_484);
or U2533 (N_2533,N_1150,N_924);
xor U2534 (N_2534,N_349,N_1734);
xnor U2535 (N_2535,N_607,N_392);
nor U2536 (N_2536,N_699,N_1720);
or U2537 (N_2537,N_965,N_736);
and U2538 (N_2538,N_1893,N_1874);
or U2539 (N_2539,N_383,N_1);
xor U2540 (N_2540,N_813,N_1032);
nor U2541 (N_2541,N_1133,N_638);
and U2542 (N_2542,N_975,N_1542);
nand U2543 (N_2543,N_1797,N_107);
or U2544 (N_2544,N_284,N_917);
xnor U2545 (N_2545,N_552,N_1366);
nor U2546 (N_2546,N_1429,N_561);
nand U2547 (N_2547,N_275,N_64);
xnor U2548 (N_2548,N_1689,N_1134);
nor U2549 (N_2549,N_211,N_1638);
xnor U2550 (N_2550,N_1990,N_445);
nor U2551 (N_2551,N_1635,N_1373);
nand U2552 (N_2552,N_1791,N_1009);
xor U2553 (N_2553,N_265,N_1183);
xnor U2554 (N_2554,N_1845,N_1029);
nand U2555 (N_2555,N_1742,N_298);
xor U2556 (N_2556,N_373,N_193);
nor U2557 (N_2557,N_1394,N_1526);
nand U2558 (N_2558,N_493,N_135);
nor U2559 (N_2559,N_243,N_1165);
nor U2560 (N_2560,N_835,N_1306);
nand U2561 (N_2561,N_1686,N_330);
or U2562 (N_2562,N_1325,N_1197);
nor U2563 (N_2563,N_572,N_441);
nor U2564 (N_2564,N_174,N_1996);
xor U2565 (N_2565,N_549,N_654);
or U2566 (N_2566,N_788,N_1441);
and U2567 (N_2567,N_1989,N_763);
nand U2568 (N_2568,N_1651,N_1226);
or U2569 (N_2569,N_1485,N_981);
nand U2570 (N_2570,N_1047,N_1840);
or U2571 (N_2571,N_286,N_1559);
nand U2572 (N_2572,N_963,N_1302);
xnor U2573 (N_2573,N_87,N_916);
xnor U2574 (N_2574,N_1735,N_793);
nor U2575 (N_2575,N_22,N_39);
nand U2576 (N_2576,N_1774,N_1695);
or U2577 (N_2577,N_1628,N_36);
nor U2578 (N_2578,N_380,N_1144);
and U2579 (N_2579,N_1835,N_1923);
and U2580 (N_2580,N_1212,N_674);
or U2581 (N_2581,N_208,N_1336);
xor U2582 (N_2582,N_110,N_14);
nor U2583 (N_2583,N_220,N_119);
or U2584 (N_2584,N_1002,N_1673);
and U2585 (N_2585,N_1873,N_201);
and U2586 (N_2586,N_826,N_777);
and U2587 (N_2587,N_1178,N_1078);
xnor U2588 (N_2588,N_399,N_906);
nand U2589 (N_2589,N_1992,N_1126);
xor U2590 (N_2590,N_1611,N_228);
nor U2591 (N_2591,N_595,N_729);
or U2592 (N_2592,N_372,N_352);
and U2593 (N_2593,N_1430,N_1969);
xor U2594 (N_2594,N_1786,N_743);
xnor U2595 (N_2595,N_1928,N_1560);
and U2596 (N_2596,N_1859,N_1147);
nand U2597 (N_2597,N_222,N_1457);
xnor U2598 (N_2598,N_1709,N_501);
and U2599 (N_2599,N_303,N_592);
nor U2600 (N_2600,N_10,N_341);
xnor U2601 (N_2601,N_570,N_1853);
xnor U2602 (N_2602,N_248,N_12);
nand U2603 (N_2603,N_1513,N_663);
and U2604 (N_2604,N_1624,N_1503);
nor U2605 (N_2605,N_611,N_259);
nand U2606 (N_2606,N_1030,N_157);
xor U2607 (N_2607,N_460,N_1766);
xnor U2608 (N_2608,N_884,N_405);
and U2609 (N_2609,N_631,N_922);
xor U2610 (N_2610,N_1496,N_1978);
nand U2611 (N_2611,N_702,N_258);
nand U2612 (N_2612,N_447,N_1412);
nand U2613 (N_2613,N_1744,N_1201);
and U2614 (N_2614,N_146,N_1209);
and U2615 (N_2615,N_1020,N_1909);
and U2616 (N_2616,N_594,N_62);
and U2617 (N_2617,N_327,N_1455);
nand U2618 (N_2618,N_27,N_591);
xnor U2619 (N_2619,N_137,N_1631);
nand U2620 (N_2620,N_164,N_167);
nand U2621 (N_2621,N_1028,N_1110);
and U2622 (N_2622,N_880,N_673);
nor U2623 (N_2623,N_1050,N_238);
nand U2624 (N_2624,N_370,N_461);
nor U2625 (N_2625,N_927,N_969);
nor U2626 (N_2626,N_869,N_1834);
or U2627 (N_2627,N_653,N_1024);
nor U2628 (N_2628,N_1269,N_1549);
and U2629 (N_2629,N_1132,N_670);
nand U2630 (N_2630,N_1979,N_1317);
nor U2631 (N_2631,N_1123,N_1789);
nor U2632 (N_2632,N_557,N_1473);
nor U2633 (N_2633,N_37,N_998);
or U2634 (N_2634,N_583,N_24);
nor U2635 (N_2635,N_1802,N_701);
or U2636 (N_2636,N_1272,N_428);
nand U2637 (N_2637,N_575,N_593);
xnor U2638 (N_2638,N_1125,N_523);
and U2639 (N_2639,N_528,N_987);
and U2640 (N_2640,N_1625,N_351);
nand U2641 (N_2641,N_1318,N_407);
nor U2642 (N_2642,N_235,N_1191);
xnor U2643 (N_2643,N_229,N_1852);
or U2644 (N_2644,N_13,N_276);
xor U2645 (N_2645,N_525,N_1018);
or U2646 (N_2646,N_741,N_1899);
xnor U2647 (N_2647,N_100,N_192);
xnor U2648 (N_2648,N_47,N_1419);
nor U2649 (N_2649,N_1736,N_1320);
nand U2650 (N_2650,N_123,N_1312);
xor U2651 (N_2651,N_1006,N_1831);
nor U2652 (N_2652,N_955,N_1741);
and U2653 (N_2653,N_470,N_1525);
nand U2654 (N_2654,N_398,N_901);
nand U2655 (N_2655,N_239,N_1410);
xor U2656 (N_2656,N_1687,N_1776);
nor U2657 (N_2657,N_1529,N_1459);
nand U2658 (N_2658,N_806,N_492);
nor U2659 (N_2659,N_684,N_800);
xor U2660 (N_2660,N_1265,N_175);
xnor U2661 (N_2661,N_919,N_742);
nor U2662 (N_2662,N_321,N_410);
nand U2663 (N_2663,N_401,N_254);
xnor U2664 (N_2664,N_1435,N_1477);
or U2665 (N_2665,N_1446,N_853);
and U2666 (N_2666,N_1639,N_876);
nor U2667 (N_2667,N_71,N_747);
nor U2668 (N_2668,N_1793,N_1294);
or U2669 (N_2669,N_377,N_414);
xnor U2670 (N_2670,N_1440,N_350);
and U2671 (N_2671,N_374,N_1066);
xor U2672 (N_2672,N_45,N_58);
or U2673 (N_2673,N_1685,N_301);
nor U2674 (N_2674,N_486,N_1645);
nor U2675 (N_2675,N_1708,N_1296);
and U2676 (N_2676,N_1544,N_1807);
nor U2677 (N_2677,N_863,N_504);
xnor U2678 (N_2678,N_809,N_808);
nand U2679 (N_2679,N_93,N_385);
and U2680 (N_2680,N_347,N_151);
nor U2681 (N_2681,N_1633,N_1180);
xnor U2682 (N_2682,N_1051,N_870);
and U2683 (N_2683,N_1199,N_195);
and U2684 (N_2684,N_1164,N_1701);
nand U2685 (N_2685,N_1775,N_403);
xor U2686 (N_2686,N_132,N_994);
nand U2687 (N_2687,N_1843,N_1658);
xnor U2688 (N_2688,N_1563,N_1378);
xnor U2689 (N_2689,N_1087,N_1622);
or U2690 (N_2690,N_292,N_1249);
nand U2691 (N_2691,N_816,N_1587);
nor U2692 (N_2692,N_898,N_1060);
nand U2693 (N_2693,N_1690,N_387);
or U2694 (N_2694,N_365,N_342);
xor U2695 (N_2695,N_1453,N_1892);
nor U2696 (N_2696,N_936,N_1956);
nor U2697 (N_2697,N_128,N_1642);
or U2698 (N_2698,N_723,N_1353);
or U2699 (N_2699,N_1514,N_1851);
xor U2700 (N_2700,N_677,N_203);
or U2701 (N_2701,N_1692,N_543);
nand U2702 (N_2702,N_453,N_1168);
and U2703 (N_2703,N_1250,N_854);
nand U2704 (N_2704,N_811,N_1193);
nand U2705 (N_2705,N_1090,N_206);
nand U2706 (N_2706,N_1468,N_938);
xnor U2707 (N_2707,N_1112,N_1334);
nand U2708 (N_2708,N_634,N_18);
nand U2709 (N_2709,N_1160,N_1465);
nor U2710 (N_2710,N_1561,N_1919);
nand U2711 (N_2711,N_1520,N_1129);
nand U2712 (N_2712,N_233,N_497);
and U2713 (N_2713,N_1920,N_1071);
or U2714 (N_2714,N_731,N_1490);
nor U2715 (N_2715,N_585,N_1716);
nor U2716 (N_2716,N_1654,N_1674);
or U2717 (N_2717,N_4,N_309);
or U2718 (N_2718,N_422,N_698);
or U2719 (N_2719,N_878,N_17);
and U2720 (N_2720,N_681,N_471);
nand U2721 (N_2721,N_686,N_1955);
and U2722 (N_2722,N_1085,N_1405);
xnor U2723 (N_2723,N_1175,N_502);
nand U2724 (N_2724,N_1383,N_1778);
nand U2725 (N_2725,N_418,N_947);
xnor U2726 (N_2726,N_926,N_801);
nor U2727 (N_2727,N_196,N_1784);
or U2728 (N_2728,N_578,N_825);
xnor U2729 (N_2729,N_1169,N_1721);
nand U2730 (N_2730,N_1927,N_227);
nor U2731 (N_2731,N_1084,N_35);
nor U2732 (N_2732,N_102,N_1054);
nor U2733 (N_2733,N_1973,N_1289);
nor U2734 (N_2734,N_1041,N_1156);
xnor U2735 (N_2735,N_948,N_1816);
or U2736 (N_2736,N_409,N_1507);
and U2737 (N_2737,N_745,N_344);
and U2738 (N_2738,N_1332,N_180);
and U2739 (N_2739,N_1487,N_1340);
and U2740 (N_2740,N_1149,N_462);
nor U2741 (N_2741,N_1896,N_1271);
and U2742 (N_2742,N_1426,N_775);
nand U2743 (N_2743,N_568,N_730);
and U2744 (N_2744,N_225,N_1258);
nor U2745 (N_2745,N_1121,N_406);
or U2746 (N_2746,N_822,N_439);
nand U2747 (N_2747,N_1245,N_1895);
nor U2748 (N_2748,N_1779,N_218);
nor U2749 (N_2749,N_717,N_553);
xnor U2750 (N_2750,N_546,N_589);
xor U2751 (N_2751,N_179,N_1408);
xor U2752 (N_2752,N_1875,N_1138);
nand U2753 (N_2753,N_1676,N_317);
nor U2754 (N_2754,N_780,N_316);
nor U2755 (N_2755,N_534,N_1447);
or U2756 (N_2756,N_294,N_1796);
nand U2757 (N_2757,N_784,N_1420);
or U2758 (N_2758,N_992,N_1566);
nor U2759 (N_2759,N_78,N_28);
nand U2760 (N_2760,N_103,N_1350);
and U2761 (N_2761,N_1136,N_1015);
xnor U2762 (N_2762,N_154,N_1392);
or U2763 (N_2763,N_456,N_496);
nand U2764 (N_2764,N_1971,N_1411);
or U2765 (N_2765,N_335,N_521);
nand U2766 (N_2766,N_1962,N_1463);
xor U2767 (N_2767,N_1450,N_230);
xnor U2768 (N_2768,N_1375,N_725);
xor U2769 (N_2769,N_868,N_724);
nand U2770 (N_2770,N_1839,N_719);
nand U2771 (N_2771,N_124,N_1374);
nor U2772 (N_2772,N_915,N_1151);
nand U2773 (N_2773,N_118,N_694);
or U2774 (N_2774,N_1448,N_988);
xor U2775 (N_2775,N_1570,N_469);
or U2776 (N_2776,N_1938,N_1130);
nand U2777 (N_2777,N_1343,N_1934);
nor U2778 (N_2778,N_1773,N_609);
or U2779 (N_2779,N_1244,N_242);
or U2780 (N_2780,N_541,N_1691);
xor U2781 (N_2781,N_1672,N_1601);
or U2782 (N_2782,N_166,N_1251);
xor U2783 (N_2783,N_1314,N_155);
nand U2784 (N_2784,N_291,N_712);
or U2785 (N_2785,N_1517,N_6);
and U2786 (N_2786,N_311,N_1590);
nor U2787 (N_2787,N_43,N_60);
and U2788 (N_2788,N_874,N_1693);
nor U2789 (N_2789,N_1335,N_1264);
and U2790 (N_2790,N_757,N_1662);
nand U2791 (N_2791,N_1602,N_1887);
nor U2792 (N_2792,N_1656,N_1801);
and U2793 (N_2793,N_856,N_1338);
nor U2794 (N_2794,N_1305,N_457);
nor U2795 (N_2795,N_540,N_168);
xor U2796 (N_2796,N_1754,N_1499);
and U2797 (N_2797,N_734,N_1096);
and U2798 (N_2798,N_1380,N_1997);
and U2799 (N_2799,N_340,N_1552);
or U2800 (N_2800,N_671,N_918);
or U2801 (N_2801,N_283,N_369);
and U2802 (N_2802,N_1719,N_1886);
nor U2803 (N_2803,N_586,N_421);
and U2804 (N_2804,N_1765,N_597);
and U2805 (N_2805,N_464,N_1182);
nand U2806 (N_2806,N_1176,N_1415);
or U2807 (N_2807,N_1609,N_1748);
xnor U2808 (N_2808,N_0,N_1505);
nand U2809 (N_2809,N_873,N_1610);
nand U2810 (N_2810,N_1202,N_1890);
xor U2811 (N_2811,N_226,N_1309);
nor U2812 (N_2812,N_289,N_1095);
nor U2813 (N_2813,N_1752,N_450);
xor U2814 (N_2814,N_1889,N_1082);
and U2815 (N_2815,N_1521,N_313);
and U2816 (N_2816,N_1484,N_1399);
or U2817 (N_2817,N_1494,N_1855);
xnor U2818 (N_2818,N_1031,N_831);
nand U2819 (N_2819,N_1678,N_223);
or U2820 (N_2820,N_1728,N_361);
nand U2821 (N_2821,N_336,N_805);
xor U2822 (N_2822,N_949,N_478);
nor U2823 (N_2823,N_860,N_98);
xnor U2824 (N_2824,N_1267,N_278);
nand U2825 (N_2825,N_797,N_420);
or U2826 (N_2826,N_305,N_958);
or U2827 (N_2827,N_1194,N_40);
or U2828 (N_2828,N_623,N_596);
nor U2829 (N_2829,N_287,N_637);
nand U2830 (N_2830,N_109,N_339);
and U2831 (N_2831,N_786,N_1750);
nand U2832 (N_2832,N_921,N_1158);
nor U2833 (N_2833,N_1292,N_939);
nor U2834 (N_2834,N_490,N_1425);
nor U2835 (N_2835,N_576,N_1922);
or U2836 (N_2836,N_1157,N_894);
and U2837 (N_2837,N_1059,N_669);
xnor U2838 (N_2838,N_752,N_581);
and U2839 (N_2839,N_1894,N_1075);
nor U2840 (N_2840,N_413,N_841);
and U2841 (N_2841,N_1762,N_499);
and U2842 (N_2842,N_1717,N_112);
xor U2843 (N_2843,N_1537,N_627);
xnor U2844 (N_2844,N_1313,N_1548);
and U2845 (N_2845,N_1324,N_1607);
or U2846 (N_2846,N_253,N_791);
xor U2847 (N_2847,N_542,N_131);
xor U2848 (N_2848,N_1333,N_268);
nor U2849 (N_2849,N_328,N_1556);
nand U2850 (N_2850,N_1056,N_1452);
nand U2851 (N_2851,N_772,N_1705);
xnor U2852 (N_2852,N_1035,N_1724);
nor U2853 (N_2853,N_411,N_1604);
xnor U2854 (N_2854,N_601,N_605);
and U2855 (N_2855,N_302,N_1361);
nand U2856 (N_2856,N_1613,N_1255);
or U2857 (N_2857,N_1637,N_796);
and U2858 (N_2858,N_143,N_279);
nand U2859 (N_2859,N_355,N_495);
or U2860 (N_2860,N_1360,N_509);
or U2861 (N_2861,N_1506,N_781);
nand U2862 (N_2862,N_272,N_1900);
or U2863 (N_2863,N_1254,N_1003);
nor U2864 (N_2864,N_452,N_159);
and U2865 (N_2865,N_172,N_1342);
and U2866 (N_2866,N_1764,N_902);
nand U2867 (N_2867,N_779,N_1039);
or U2868 (N_2868,N_687,N_1573);
nand U2869 (N_2869,N_1358,N_1211);
xnor U2870 (N_2870,N_1285,N_148);
xnor U2871 (N_2871,N_169,N_1376);
nor U2872 (N_2872,N_1382,N_153);
xor U2873 (N_2873,N_1471,N_1321);
xnor U2874 (N_2874,N_1304,N_1288);
nand U2875 (N_2875,N_1648,N_1227);
and U2876 (N_2876,N_1492,N_255);
xor U2877 (N_2877,N_1489,N_295);
and U2878 (N_2878,N_1832,N_879);
and U2879 (N_2879,N_438,N_1715);
and U2880 (N_2880,N_96,N_656);
nand U2881 (N_2881,N_178,N_1808);
and U2882 (N_2882,N_533,N_1787);
nor U2883 (N_2883,N_160,N_315);
nand U2884 (N_2884,N_708,N_899);
or U2885 (N_2885,N_1277,N_990);
nor U2886 (N_2886,N_1099,N_714);
or U2887 (N_2887,N_1357,N_1711);
nand U2888 (N_2888,N_588,N_1974);
and U2889 (N_2889,N_52,N_1184);
or U2890 (N_2890,N_1870,N_820);
nand U2891 (N_2891,N_306,N_1196);
nor U2892 (N_2892,N_807,N_224);
nand U2893 (N_2893,N_1794,N_127);
or U2894 (N_2894,N_1551,N_42);
or U2895 (N_2895,N_429,N_1533);
xnor U2896 (N_2896,N_117,N_1630);
xor U2897 (N_2897,N_828,N_1546);
nand U2898 (N_2898,N_50,N_402);
nand U2899 (N_2899,N_1153,N_1239);
nor U2900 (N_2900,N_1372,N_1034);
or U2901 (N_2901,N_1641,N_85);
nand U2902 (N_2902,N_1510,N_721);
xnor U2903 (N_2903,N_1073,N_427);
or U2904 (N_2904,N_446,N_378);
xor U2905 (N_2905,N_1462,N_1806);
nand U2906 (N_2906,N_1345,N_1439);
nor U2907 (N_2907,N_931,N_354);
and U2908 (N_2908,N_1482,N_448);
nand U2909 (N_2909,N_121,N_1871);
or U2910 (N_2910,N_1512,N_467);
nand U2911 (N_2911,N_782,N_750);
nor U2912 (N_2912,N_1297,N_74);
or U2913 (N_2913,N_2,N_1567);
or U2914 (N_2914,N_1849,N_1445);
nand U2915 (N_2915,N_300,N_544);
nand U2916 (N_2916,N_133,N_273);
and U2917 (N_2917,N_1817,N_675);
xnor U2918 (N_2918,N_624,N_367);
or U2919 (N_2919,N_1057,N_1001);
or U2920 (N_2920,N_252,N_633);
and U2921 (N_2921,N_937,N_1458);
nor U2922 (N_2922,N_636,N_1952);
and U2923 (N_2923,N_1914,N_16);
nand U2924 (N_2924,N_897,N_200);
xnor U2925 (N_2925,N_1931,N_1846);
nand U2926 (N_2926,N_954,N_1081);
or U2927 (N_2927,N_1942,N_749);
nand U2928 (N_2928,N_150,N_1421);
and U2929 (N_2929,N_855,N_810);
xor U2930 (N_2930,N_1068,N_877);
and U2931 (N_2931,N_141,N_1950);
nand U2932 (N_2932,N_657,N_468);
nand U2933 (N_2933,N_908,N_1495);
or U2934 (N_2934,N_472,N_1980);
nor U2935 (N_2935,N_974,N_1022);
and U2936 (N_2936,N_1498,N_584);
nor U2937 (N_2937,N_1406,N_803);
nor U2938 (N_2938,N_1603,N_1287);
nand U2939 (N_2939,N_33,N_1912);
xnor U2940 (N_2940,N_928,N_1588);
xor U2941 (N_2941,N_1220,N_104);
or U2942 (N_2942,N_1737,N_1977);
and U2943 (N_2943,N_1480,N_1109);
and U2944 (N_2944,N_1217,N_817);
nor U2945 (N_2945,N_1113,N_1356);
nor U2946 (N_2946,N_1504,N_1706);
and U2947 (N_2947,N_1768,N_1883);
xor U2948 (N_2948,N_1634,N_1092);
nand U2949 (N_2949,N_972,N_1362);
or U2950 (N_2950,N_950,N_618);
or U2951 (N_2951,N_1930,N_903);
nor U2952 (N_2952,N_1679,N_1274);
or U2953 (N_2953,N_1905,N_308);
nor U2954 (N_2954,N_1004,N_941);
nor U2955 (N_2955,N_1810,N_1857);
and U2956 (N_2956,N_1451,N_547);
and U2957 (N_2957,N_76,N_1901);
xnor U2958 (N_2958,N_125,N_535);
nand U2959 (N_2959,N_1856,N_1703);
nand U2960 (N_2960,N_565,N_1878);
xor U2961 (N_2961,N_163,N_1083);
nand U2962 (N_2962,N_1585,N_689);
nand U2963 (N_2963,N_1777,N_426);
and U2964 (N_2964,N_555,N_1746);
xnor U2965 (N_2965,N_1270,N_423);
xor U2966 (N_2966,N_1515,N_1903);
xnor U2967 (N_2967,N_999,N_363);
and U2968 (N_2968,N_324,N_577);
xor U2969 (N_2969,N_358,N_1697);
or U2970 (N_2970,N_740,N_1837);
nor U2971 (N_2971,N_419,N_1045);
and U2972 (N_2972,N_1681,N_442);
and U2973 (N_2973,N_704,N_667);
and U2974 (N_2974,N_1963,N_1187);
and U2975 (N_2975,N_1730,N_707);
xor U2976 (N_2976,N_1203,N_91);
xnor U2977 (N_2977,N_182,N_1844);
nand U2978 (N_2978,N_1961,N_1725);
nand U2979 (N_2979,N_773,N_890);
xnor U2980 (N_2980,N_838,N_1819);
xnor U2981 (N_2981,N_1502,N_382);
nand U2982 (N_2982,N_1000,N_1805);
and U2983 (N_2983,N_1331,N_237);
or U2984 (N_2984,N_1939,N_1038);
nand U2985 (N_2985,N_1760,N_661);
and U2986 (N_2986,N_1390,N_1208);
or U2987 (N_2987,N_1248,N_852);
or U2988 (N_2988,N_432,N_1300);
nor U2989 (N_2989,N_55,N_1391);
nor U2990 (N_2990,N_1993,N_840);
nor U2991 (N_2991,N_1014,N_1072);
or U2992 (N_2992,N_129,N_1454);
xor U2993 (N_2993,N_84,N_1675);
nand U2994 (N_2994,N_871,N_236);
xor U2995 (N_2995,N_932,N_625);
xor U2996 (N_2996,N_48,N_1179);
xor U2997 (N_2997,N_1261,N_1558);
nor U2998 (N_2998,N_944,N_1231);
nor U2999 (N_2999,N_1491,N_755);
nand U3000 (N_3000,N_371,N_233);
nand U3001 (N_3001,N_358,N_1830);
or U3002 (N_3002,N_1966,N_1246);
nor U3003 (N_3003,N_8,N_552);
nand U3004 (N_3004,N_1718,N_1061);
and U3005 (N_3005,N_1734,N_379);
and U3006 (N_3006,N_348,N_527);
or U3007 (N_3007,N_904,N_1831);
and U3008 (N_3008,N_1401,N_1569);
or U3009 (N_3009,N_175,N_1685);
nor U3010 (N_3010,N_1404,N_794);
or U3011 (N_3011,N_121,N_179);
nand U3012 (N_3012,N_1415,N_482);
nor U3013 (N_3013,N_154,N_1179);
xor U3014 (N_3014,N_1517,N_160);
xor U3015 (N_3015,N_1526,N_1649);
nand U3016 (N_3016,N_156,N_903);
and U3017 (N_3017,N_1385,N_1225);
and U3018 (N_3018,N_1466,N_1097);
nand U3019 (N_3019,N_1567,N_1432);
nand U3020 (N_3020,N_1808,N_769);
nor U3021 (N_3021,N_1858,N_752);
and U3022 (N_3022,N_1891,N_198);
and U3023 (N_3023,N_1256,N_1009);
xnor U3024 (N_3024,N_71,N_563);
nor U3025 (N_3025,N_1625,N_1909);
or U3026 (N_3026,N_1449,N_1211);
nand U3027 (N_3027,N_198,N_1668);
and U3028 (N_3028,N_622,N_944);
nand U3029 (N_3029,N_323,N_1811);
xnor U3030 (N_3030,N_1837,N_1128);
xnor U3031 (N_3031,N_1583,N_601);
xnor U3032 (N_3032,N_542,N_1770);
nor U3033 (N_3033,N_888,N_410);
or U3034 (N_3034,N_334,N_1302);
nor U3035 (N_3035,N_914,N_1106);
or U3036 (N_3036,N_1202,N_510);
nor U3037 (N_3037,N_115,N_124);
nor U3038 (N_3038,N_977,N_29);
nor U3039 (N_3039,N_104,N_1942);
nand U3040 (N_3040,N_1901,N_1355);
nand U3041 (N_3041,N_609,N_1142);
nand U3042 (N_3042,N_225,N_1134);
or U3043 (N_3043,N_1598,N_1609);
nand U3044 (N_3044,N_1423,N_1139);
nand U3045 (N_3045,N_1925,N_47);
or U3046 (N_3046,N_327,N_1336);
nor U3047 (N_3047,N_321,N_1351);
nor U3048 (N_3048,N_1201,N_509);
nand U3049 (N_3049,N_794,N_1958);
and U3050 (N_3050,N_557,N_866);
or U3051 (N_3051,N_139,N_677);
xor U3052 (N_3052,N_1726,N_1280);
or U3053 (N_3053,N_42,N_1834);
or U3054 (N_3054,N_259,N_1227);
nand U3055 (N_3055,N_1597,N_265);
nor U3056 (N_3056,N_1298,N_1529);
nor U3057 (N_3057,N_861,N_1021);
or U3058 (N_3058,N_382,N_992);
or U3059 (N_3059,N_46,N_72);
or U3060 (N_3060,N_1011,N_907);
and U3061 (N_3061,N_264,N_1808);
nand U3062 (N_3062,N_774,N_385);
nor U3063 (N_3063,N_58,N_1282);
nor U3064 (N_3064,N_1665,N_967);
nor U3065 (N_3065,N_1840,N_1277);
or U3066 (N_3066,N_1559,N_1027);
and U3067 (N_3067,N_138,N_1924);
xor U3068 (N_3068,N_703,N_240);
xnor U3069 (N_3069,N_335,N_1217);
or U3070 (N_3070,N_377,N_1811);
or U3071 (N_3071,N_1750,N_1146);
and U3072 (N_3072,N_1070,N_445);
xor U3073 (N_3073,N_410,N_196);
and U3074 (N_3074,N_1543,N_726);
nor U3075 (N_3075,N_1188,N_13);
and U3076 (N_3076,N_1763,N_586);
nor U3077 (N_3077,N_395,N_1545);
nand U3078 (N_3078,N_1570,N_959);
nor U3079 (N_3079,N_1046,N_966);
xor U3080 (N_3080,N_1130,N_1768);
nor U3081 (N_3081,N_161,N_800);
and U3082 (N_3082,N_223,N_1406);
and U3083 (N_3083,N_1869,N_1351);
xor U3084 (N_3084,N_1912,N_152);
and U3085 (N_3085,N_50,N_1572);
nor U3086 (N_3086,N_1364,N_1724);
and U3087 (N_3087,N_320,N_305);
nor U3088 (N_3088,N_977,N_1956);
nand U3089 (N_3089,N_512,N_1971);
or U3090 (N_3090,N_1455,N_1165);
nand U3091 (N_3091,N_1252,N_1535);
nand U3092 (N_3092,N_440,N_1715);
nor U3093 (N_3093,N_986,N_137);
nand U3094 (N_3094,N_630,N_1919);
and U3095 (N_3095,N_1686,N_10);
nor U3096 (N_3096,N_1363,N_839);
xnor U3097 (N_3097,N_961,N_758);
or U3098 (N_3098,N_989,N_1690);
xnor U3099 (N_3099,N_1833,N_357);
nand U3100 (N_3100,N_36,N_1346);
xnor U3101 (N_3101,N_391,N_542);
or U3102 (N_3102,N_696,N_448);
or U3103 (N_3103,N_822,N_1292);
or U3104 (N_3104,N_1406,N_1538);
xor U3105 (N_3105,N_351,N_1504);
nand U3106 (N_3106,N_1652,N_1535);
nor U3107 (N_3107,N_957,N_1138);
nor U3108 (N_3108,N_486,N_1926);
nor U3109 (N_3109,N_1044,N_300);
nor U3110 (N_3110,N_1081,N_1350);
xor U3111 (N_3111,N_1412,N_1976);
xor U3112 (N_3112,N_416,N_1140);
nor U3113 (N_3113,N_1864,N_21);
nand U3114 (N_3114,N_513,N_1447);
nor U3115 (N_3115,N_1550,N_107);
nand U3116 (N_3116,N_1640,N_1180);
and U3117 (N_3117,N_1031,N_321);
nand U3118 (N_3118,N_735,N_129);
xor U3119 (N_3119,N_1472,N_1410);
xor U3120 (N_3120,N_393,N_1957);
nand U3121 (N_3121,N_602,N_1863);
nor U3122 (N_3122,N_411,N_1162);
nor U3123 (N_3123,N_435,N_1648);
or U3124 (N_3124,N_168,N_1924);
nand U3125 (N_3125,N_1512,N_361);
nor U3126 (N_3126,N_226,N_951);
or U3127 (N_3127,N_1581,N_267);
nand U3128 (N_3128,N_456,N_842);
or U3129 (N_3129,N_613,N_1851);
xnor U3130 (N_3130,N_1989,N_1194);
xor U3131 (N_3131,N_1372,N_805);
or U3132 (N_3132,N_1742,N_496);
nand U3133 (N_3133,N_1562,N_1757);
and U3134 (N_3134,N_1141,N_1097);
xnor U3135 (N_3135,N_1295,N_710);
nand U3136 (N_3136,N_385,N_1892);
nand U3137 (N_3137,N_133,N_425);
xor U3138 (N_3138,N_1439,N_1142);
xnor U3139 (N_3139,N_589,N_1357);
nand U3140 (N_3140,N_1856,N_215);
nor U3141 (N_3141,N_1893,N_60);
and U3142 (N_3142,N_333,N_899);
xnor U3143 (N_3143,N_1762,N_110);
nor U3144 (N_3144,N_67,N_1115);
nand U3145 (N_3145,N_1559,N_183);
or U3146 (N_3146,N_1433,N_1477);
nor U3147 (N_3147,N_171,N_1498);
nand U3148 (N_3148,N_845,N_1098);
nand U3149 (N_3149,N_870,N_1200);
nor U3150 (N_3150,N_506,N_979);
nand U3151 (N_3151,N_600,N_1521);
nor U3152 (N_3152,N_1793,N_1428);
nor U3153 (N_3153,N_498,N_1318);
nor U3154 (N_3154,N_1566,N_303);
nor U3155 (N_3155,N_1958,N_1197);
xnor U3156 (N_3156,N_922,N_815);
nor U3157 (N_3157,N_347,N_876);
xor U3158 (N_3158,N_126,N_1848);
nor U3159 (N_3159,N_1531,N_1616);
xor U3160 (N_3160,N_1307,N_351);
nand U3161 (N_3161,N_134,N_986);
xnor U3162 (N_3162,N_1911,N_1720);
xnor U3163 (N_3163,N_1653,N_359);
nor U3164 (N_3164,N_1212,N_1210);
nand U3165 (N_3165,N_273,N_1600);
nand U3166 (N_3166,N_732,N_962);
nand U3167 (N_3167,N_256,N_1416);
or U3168 (N_3168,N_890,N_481);
nor U3169 (N_3169,N_345,N_1932);
nand U3170 (N_3170,N_1670,N_1576);
and U3171 (N_3171,N_1536,N_716);
or U3172 (N_3172,N_1428,N_1253);
or U3173 (N_3173,N_1390,N_30);
nor U3174 (N_3174,N_1426,N_1414);
xnor U3175 (N_3175,N_1101,N_1686);
xnor U3176 (N_3176,N_1439,N_142);
xnor U3177 (N_3177,N_24,N_549);
nor U3178 (N_3178,N_1520,N_1249);
xnor U3179 (N_3179,N_472,N_1348);
xor U3180 (N_3180,N_1817,N_1123);
or U3181 (N_3181,N_1274,N_1826);
xnor U3182 (N_3182,N_1924,N_1415);
and U3183 (N_3183,N_1245,N_180);
xor U3184 (N_3184,N_1760,N_1702);
or U3185 (N_3185,N_807,N_119);
xnor U3186 (N_3186,N_1116,N_1263);
nor U3187 (N_3187,N_1947,N_246);
xnor U3188 (N_3188,N_991,N_1872);
xor U3189 (N_3189,N_610,N_1550);
and U3190 (N_3190,N_1984,N_1717);
nor U3191 (N_3191,N_733,N_1489);
and U3192 (N_3192,N_1338,N_932);
or U3193 (N_3193,N_940,N_1362);
xnor U3194 (N_3194,N_1931,N_1765);
nor U3195 (N_3195,N_469,N_1715);
nor U3196 (N_3196,N_1621,N_412);
or U3197 (N_3197,N_1753,N_383);
nand U3198 (N_3198,N_506,N_1042);
xor U3199 (N_3199,N_687,N_802);
or U3200 (N_3200,N_208,N_764);
xor U3201 (N_3201,N_310,N_242);
nor U3202 (N_3202,N_1633,N_764);
xor U3203 (N_3203,N_1813,N_502);
or U3204 (N_3204,N_1180,N_72);
nor U3205 (N_3205,N_1012,N_334);
nand U3206 (N_3206,N_1691,N_381);
and U3207 (N_3207,N_1203,N_1285);
nand U3208 (N_3208,N_925,N_1371);
xnor U3209 (N_3209,N_1565,N_1691);
xor U3210 (N_3210,N_667,N_1442);
nor U3211 (N_3211,N_1951,N_1593);
nor U3212 (N_3212,N_465,N_793);
or U3213 (N_3213,N_566,N_710);
nand U3214 (N_3214,N_1939,N_1081);
and U3215 (N_3215,N_1200,N_1179);
and U3216 (N_3216,N_1215,N_1932);
and U3217 (N_3217,N_742,N_905);
nor U3218 (N_3218,N_392,N_1336);
and U3219 (N_3219,N_1587,N_864);
and U3220 (N_3220,N_218,N_1227);
xor U3221 (N_3221,N_401,N_41);
nand U3222 (N_3222,N_358,N_385);
nand U3223 (N_3223,N_1519,N_1487);
or U3224 (N_3224,N_1049,N_1363);
nor U3225 (N_3225,N_94,N_838);
xor U3226 (N_3226,N_1802,N_1872);
or U3227 (N_3227,N_1001,N_1186);
nor U3228 (N_3228,N_544,N_1668);
and U3229 (N_3229,N_1873,N_782);
and U3230 (N_3230,N_0,N_412);
nand U3231 (N_3231,N_640,N_723);
and U3232 (N_3232,N_878,N_178);
nor U3233 (N_3233,N_1437,N_1812);
or U3234 (N_3234,N_483,N_678);
nand U3235 (N_3235,N_1624,N_1092);
nand U3236 (N_3236,N_1619,N_1093);
or U3237 (N_3237,N_762,N_1197);
nor U3238 (N_3238,N_1796,N_682);
xnor U3239 (N_3239,N_1611,N_840);
xnor U3240 (N_3240,N_248,N_1890);
and U3241 (N_3241,N_524,N_431);
and U3242 (N_3242,N_878,N_1240);
and U3243 (N_3243,N_1397,N_422);
nor U3244 (N_3244,N_332,N_1104);
or U3245 (N_3245,N_1500,N_411);
or U3246 (N_3246,N_1208,N_1721);
nand U3247 (N_3247,N_1567,N_1940);
xor U3248 (N_3248,N_1144,N_177);
nor U3249 (N_3249,N_1148,N_1617);
nand U3250 (N_3250,N_700,N_1924);
xor U3251 (N_3251,N_1929,N_1730);
xor U3252 (N_3252,N_1238,N_335);
or U3253 (N_3253,N_241,N_1897);
and U3254 (N_3254,N_1123,N_267);
xnor U3255 (N_3255,N_246,N_1366);
and U3256 (N_3256,N_1722,N_1095);
nor U3257 (N_3257,N_48,N_289);
and U3258 (N_3258,N_1681,N_501);
or U3259 (N_3259,N_697,N_913);
or U3260 (N_3260,N_211,N_1980);
and U3261 (N_3261,N_187,N_275);
or U3262 (N_3262,N_28,N_155);
nand U3263 (N_3263,N_989,N_1848);
or U3264 (N_3264,N_41,N_409);
nand U3265 (N_3265,N_845,N_1500);
xnor U3266 (N_3266,N_1564,N_1014);
xor U3267 (N_3267,N_893,N_1905);
nor U3268 (N_3268,N_713,N_322);
nor U3269 (N_3269,N_706,N_9);
nand U3270 (N_3270,N_1626,N_914);
and U3271 (N_3271,N_331,N_1547);
or U3272 (N_3272,N_791,N_44);
nand U3273 (N_3273,N_764,N_473);
nor U3274 (N_3274,N_188,N_706);
nor U3275 (N_3275,N_1808,N_1124);
xor U3276 (N_3276,N_1848,N_1814);
nor U3277 (N_3277,N_212,N_1222);
nand U3278 (N_3278,N_1352,N_1685);
nand U3279 (N_3279,N_357,N_625);
nor U3280 (N_3280,N_1941,N_1676);
or U3281 (N_3281,N_982,N_1707);
nor U3282 (N_3282,N_1845,N_50);
nor U3283 (N_3283,N_1584,N_309);
and U3284 (N_3284,N_655,N_806);
or U3285 (N_3285,N_811,N_1770);
nand U3286 (N_3286,N_1764,N_1330);
nor U3287 (N_3287,N_1922,N_321);
nand U3288 (N_3288,N_1930,N_1931);
nand U3289 (N_3289,N_897,N_824);
or U3290 (N_3290,N_266,N_1672);
and U3291 (N_3291,N_204,N_428);
xnor U3292 (N_3292,N_1228,N_1663);
nand U3293 (N_3293,N_1086,N_584);
and U3294 (N_3294,N_632,N_1819);
and U3295 (N_3295,N_1381,N_543);
nor U3296 (N_3296,N_506,N_1100);
nand U3297 (N_3297,N_417,N_295);
nand U3298 (N_3298,N_206,N_563);
or U3299 (N_3299,N_768,N_1060);
nor U3300 (N_3300,N_366,N_199);
or U3301 (N_3301,N_461,N_1406);
and U3302 (N_3302,N_1039,N_533);
and U3303 (N_3303,N_1542,N_665);
nand U3304 (N_3304,N_291,N_605);
nand U3305 (N_3305,N_1152,N_1372);
nor U3306 (N_3306,N_494,N_615);
xnor U3307 (N_3307,N_168,N_332);
nand U3308 (N_3308,N_326,N_480);
xor U3309 (N_3309,N_1997,N_903);
or U3310 (N_3310,N_674,N_365);
xnor U3311 (N_3311,N_1084,N_1082);
and U3312 (N_3312,N_1398,N_467);
or U3313 (N_3313,N_1545,N_747);
or U3314 (N_3314,N_1547,N_849);
and U3315 (N_3315,N_1255,N_1110);
and U3316 (N_3316,N_1110,N_1652);
xnor U3317 (N_3317,N_1054,N_1488);
xor U3318 (N_3318,N_918,N_50);
xor U3319 (N_3319,N_1709,N_1548);
nor U3320 (N_3320,N_778,N_1053);
nand U3321 (N_3321,N_395,N_1588);
nor U3322 (N_3322,N_1783,N_1100);
nand U3323 (N_3323,N_969,N_1310);
nor U3324 (N_3324,N_601,N_1662);
or U3325 (N_3325,N_1797,N_1726);
and U3326 (N_3326,N_1127,N_1374);
or U3327 (N_3327,N_535,N_148);
or U3328 (N_3328,N_1915,N_643);
nand U3329 (N_3329,N_997,N_482);
xnor U3330 (N_3330,N_376,N_779);
and U3331 (N_3331,N_1238,N_585);
xor U3332 (N_3332,N_425,N_494);
nand U3333 (N_3333,N_895,N_1231);
nand U3334 (N_3334,N_1483,N_853);
or U3335 (N_3335,N_1929,N_1026);
nor U3336 (N_3336,N_380,N_1763);
or U3337 (N_3337,N_1095,N_320);
and U3338 (N_3338,N_895,N_531);
nand U3339 (N_3339,N_629,N_1606);
nor U3340 (N_3340,N_1909,N_1781);
or U3341 (N_3341,N_939,N_676);
xor U3342 (N_3342,N_407,N_465);
and U3343 (N_3343,N_807,N_1915);
xnor U3344 (N_3344,N_459,N_321);
xor U3345 (N_3345,N_1409,N_1639);
or U3346 (N_3346,N_105,N_1446);
xor U3347 (N_3347,N_771,N_1933);
or U3348 (N_3348,N_644,N_565);
nor U3349 (N_3349,N_1302,N_350);
xnor U3350 (N_3350,N_317,N_658);
or U3351 (N_3351,N_294,N_947);
nand U3352 (N_3352,N_952,N_1269);
nand U3353 (N_3353,N_804,N_576);
xnor U3354 (N_3354,N_1172,N_1267);
nor U3355 (N_3355,N_778,N_1690);
nor U3356 (N_3356,N_1279,N_891);
or U3357 (N_3357,N_527,N_1348);
nor U3358 (N_3358,N_741,N_1443);
nor U3359 (N_3359,N_1979,N_799);
nor U3360 (N_3360,N_558,N_1860);
and U3361 (N_3361,N_1017,N_1564);
xnor U3362 (N_3362,N_1491,N_747);
xnor U3363 (N_3363,N_606,N_1554);
or U3364 (N_3364,N_1162,N_952);
nor U3365 (N_3365,N_1266,N_439);
nand U3366 (N_3366,N_762,N_919);
and U3367 (N_3367,N_793,N_383);
or U3368 (N_3368,N_1823,N_1942);
nor U3369 (N_3369,N_678,N_271);
nand U3370 (N_3370,N_901,N_182);
nor U3371 (N_3371,N_1419,N_1007);
nor U3372 (N_3372,N_604,N_17);
xnor U3373 (N_3373,N_1069,N_1024);
xnor U3374 (N_3374,N_1508,N_1189);
and U3375 (N_3375,N_1764,N_274);
xnor U3376 (N_3376,N_283,N_929);
nand U3377 (N_3377,N_677,N_689);
xor U3378 (N_3378,N_1182,N_1917);
or U3379 (N_3379,N_1383,N_412);
nor U3380 (N_3380,N_1925,N_820);
nor U3381 (N_3381,N_999,N_1531);
and U3382 (N_3382,N_1110,N_961);
and U3383 (N_3383,N_1808,N_531);
or U3384 (N_3384,N_1120,N_1727);
nor U3385 (N_3385,N_966,N_1631);
nand U3386 (N_3386,N_1742,N_1723);
and U3387 (N_3387,N_1909,N_419);
xnor U3388 (N_3388,N_504,N_236);
xor U3389 (N_3389,N_179,N_1997);
and U3390 (N_3390,N_489,N_577);
nand U3391 (N_3391,N_653,N_1618);
or U3392 (N_3392,N_1516,N_1855);
and U3393 (N_3393,N_1891,N_141);
nor U3394 (N_3394,N_791,N_716);
xnor U3395 (N_3395,N_1150,N_55);
nand U3396 (N_3396,N_1693,N_1605);
or U3397 (N_3397,N_1426,N_1898);
nand U3398 (N_3398,N_278,N_756);
nand U3399 (N_3399,N_1731,N_950);
or U3400 (N_3400,N_58,N_1001);
or U3401 (N_3401,N_1329,N_1842);
or U3402 (N_3402,N_1967,N_1293);
nand U3403 (N_3403,N_606,N_965);
nor U3404 (N_3404,N_474,N_1802);
xnor U3405 (N_3405,N_898,N_1499);
nor U3406 (N_3406,N_1820,N_125);
or U3407 (N_3407,N_1144,N_266);
or U3408 (N_3408,N_1203,N_1762);
and U3409 (N_3409,N_227,N_516);
and U3410 (N_3410,N_706,N_1549);
or U3411 (N_3411,N_415,N_1464);
nand U3412 (N_3412,N_219,N_1631);
or U3413 (N_3413,N_722,N_454);
nand U3414 (N_3414,N_721,N_1760);
xor U3415 (N_3415,N_643,N_388);
nor U3416 (N_3416,N_909,N_390);
xor U3417 (N_3417,N_651,N_174);
and U3418 (N_3418,N_429,N_66);
and U3419 (N_3419,N_781,N_1118);
nor U3420 (N_3420,N_1868,N_1576);
and U3421 (N_3421,N_1870,N_867);
nand U3422 (N_3422,N_1153,N_1377);
and U3423 (N_3423,N_1327,N_190);
and U3424 (N_3424,N_404,N_1487);
nand U3425 (N_3425,N_1707,N_184);
or U3426 (N_3426,N_200,N_1039);
nor U3427 (N_3427,N_1615,N_1775);
or U3428 (N_3428,N_47,N_774);
and U3429 (N_3429,N_866,N_118);
or U3430 (N_3430,N_1983,N_151);
or U3431 (N_3431,N_64,N_494);
or U3432 (N_3432,N_846,N_1599);
xnor U3433 (N_3433,N_1302,N_1195);
and U3434 (N_3434,N_1593,N_1342);
xnor U3435 (N_3435,N_1872,N_887);
or U3436 (N_3436,N_1444,N_795);
or U3437 (N_3437,N_748,N_435);
nand U3438 (N_3438,N_785,N_670);
nor U3439 (N_3439,N_997,N_1665);
or U3440 (N_3440,N_406,N_1984);
nor U3441 (N_3441,N_86,N_1338);
or U3442 (N_3442,N_1685,N_297);
nand U3443 (N_3443,N_1360,N_1488);
nand U3444 (N_3444,N_226,N_1415);
nand U3445 (N_3445,N_1970,N_350);
or U3446 (N_3446,N_1623,N_123);
xnor U3447 (N_3447,N_580,N_1683);
or U3448 (N_3448,N_1834,N_382);
xor U3449 (N_3449,N_1248,N_1220);
nor U3450 (N_3450,N_1903,N_179);
xor U3451 (N_3451,N_784,N_846);
nand U3452 (N_3452,N_255,N_1651);
and U3453 (N_3453,N_1116,N_749);
nand U3454 (N_3454,N_1931,N_522);
or U3455 (N_3455,N_194,N_978);
nor U3456 (N_3456,N_1717,N_775);
and U3457 (N_3457,N_53,N_431);
nand U3458 (N_3458,N_1791,N_1087);
nand U3459 (N_3459,N_52,N_1253);
and U3460 (N_3460,N_780,N_791);
nand U3461 (N_3461,N_206,N_375);
or U3462 (N_3462,N_257,N_753);
nor U3463 (N_3463,N_959,N_23);
nor U3464 (N_3464,N_207,N_1134);
nand U3465 (N_3465,N_1684,N_1673);
xor U3466 (N_3466,N_1653,N_1389);
or U3467 (N_3467,N_1450,N_689);
nor U3468 (N_3468,N_1239,N_1875);
nand U3469 (N_3469,N_51,N_1556);
xnor U3470 (N_3470,N_1316,N_1044);
or U3471 (N_3471,N_1597,N_1015);
xnor U3472 (N_3472,N_845,N_1367);
xor U3473 (N_3473,N_153,N_1069);
nor U3474 (N_3474,N_266,N_182);
and U3475 (N_3475,N_282,N_1929);
and U3476 (N_3476,N_988,N_1756);
and U3477 (N_3477,N_566,N_632);
or U3478 (N_3478,N_232,N_1471);
nor U3479 (N_3479,N_999,N_240);
and U3480 (N_3480,N_230,N_1598);
nor U3481 (N_3481,N_128,N_1727);
nor U3482 (N_3482,N_1208,N_1911);
and U3483 (N_3483,N_19,N_1167);
xor U3484 (N_3484,N_892,N_1611);
or U3485 (N_3485,N_52,N_362);
or U3486 (N_3486,N_1502,N_1507);
or U3487 (N_3487,N_171,N_1457);
and U3488 (N_3488,N_755,N_29);
nor U3489 (N_3489,N_1037,N_283);
nand U3490 (N_3490,N_1631,N_459);
xor U3491 (N_3491,N_1650,N_1838);
nand U3492 (N_3492,N_473,N_404);
or U3493 (N_3493,N_720,N_1479);
xor U3494 (N_3494,N_1319,N_1133);
nand U3495 (N_3495,N_1623,N_779);
or U3496 (N_3496,N_389,N_1871);
or U3497 (N_3497,N_925,N_837);
and U3498 (N_3498,N_446,N_1296);
and U3499 (N_3499,N_1812,N_1944);
or U3500 (N_3500,N_582,N_208);
nor U3501 (N_3501,N_1394,N_1909);
nor U3502 (N_3502,N_956,N_1707);
or U3503 (N_3503,N_363,N_647);
nor U3504 (N_3504,N_1429,N_1068);
xnor U3505 (N_3505,N_273,N_142);
or U3506 (N_3506,N_1999,N_694);
nor U3507 (N_3507,N_1847,N_1886);
nand U3508 (N_3508,N_841,N_666);
xor U3509 (N_3509,N_1675,N_7);
nor U3510 (N_3510,N_1402,N_1297);
and U3511 (N_3511,N_1408,N_1779);
nand U3512 (N_3512,N_943,N_431);
and U3513 (N_3513,N_184,N_379);
nand U3514 (N_3514,N_1036,N_1156);
and U3515 (N_3515,N_1075,N_749);
nor U3516 (N_3516,N_616,N_827);
nor U3517 (N_3517,N_355,N_1764);
nor U3518 (N_3518,N_1891,N_1089);
and U3519 (N_3519,N_417,N_1177);
xor U3520 (N_3520,N_514,N_1306);
and U3521 (N_3521,N_1799,N_1212);
and U3522 (N_3522,N_670,N_823);
nand U3523 (N_3523,N_1435,N_216);
or U3524 (N_3524,N_104,N_1850);
xor U3525 (N_3525,N_1455,N_365);
or U3526 (N_3526,N_328,N_96);
nor U3527 (N_3527,N_1724,N_657);
or U3528 (N_3528,N_1524,N_1482);
xnor U3529 (N_3529,N_260,N_839);
nand U3530 (N_3530,N_758,N_1643);
and U3531 (N_3531,N_1380,N_1115);
or U3532 (N_3532,N_185,N_872);
and U3533 (N_3533,N_1912,N_1256);
nand U3534 (N_3534,N_441,N_1142);
or U3535 (N_3535,N_1416,N_1894);
nor U3536 (N_3536,N_978,N_1974);
and U3537 (N_3537,N_1522,N_1126);
nor U3538 (N_3538,N_1593,N_1298);
xnor U3539 (N_3539,N_332,N_817);
and U3540 (N_3540,N_1587,N_380);
nand U3541 (N_3541,N_1951,N_673);
xor U3542 (N_3542,N_1370,N_88);
or U3543 (N_3543,N_1903,N_1446);
nor U3544 (N_3544,N_1250,N_1493);
and U3545 (N_3545,N_1056,N_822);
xnor U3546 (N_3546,N_1955,N_540);
and U3547 (N_3547,N_1797,N_883);
nand U3548 (N_3548,N_818,N_525);
nand U3549 (N_3549,N_389,N_1492);
xnor U3550 (N_3550,N_690,N_514);
nand U3551 (N_3551,N_937,N_816);
or U3552 (N_3552,N_83,N_98);
nor U3553 (N_3553,N_873,N_121);
nand U3554 (N_3554,N_476,N_1843);
or U3555 (N_3555,N_1009,N_1934);
xor U3556 (N_3556,N_932,N_1009);
and U3557 (N_3557,N_300,N_122);
nand U3558 (N_3558,N_41,N_1511);
nor U3559 (N_3559,N_42,N_104);
xnor U3560 (N_3560,N_1063,N_1927);
or U3561 (N_3561,N_689,N_274);
and U3562 (N_3562,N_7,N_1119);
nor U3563 (N_3563,N_498,N_465);
nand U3564 (N_3564,N_891,N_1272);
nand U3565 (N_3565,N_1800,N_558);
xnor U3566 (N_3566,N_1793,N_1448);
or U3567 (N_3567,N_1210,N_893);
nand U3568 (N_3568,N_1830,N_192);
or U3569 (N_3569,N_187,N_777);
nor U3570 (N_3570,N_1789,N_1350);
xor U3571 (N_3571,N_1453,N_1377);
nand U3572 (N_3572,N_149,N_976);
nor U3573 (N_3573,N_1482,N_487);
or U3574 (N_3574,N_1576,N_1903);
or U3575 (N_3575,N_544,N_850);
xor U3576 (N_3576,N_1348,N_163);
and U3577 (N_3577,N_1266,N_528);
and U3578 (N_3578,N_805,N_1298);
and U3579 (N_3579,N_470,N_594);
nand U3580 (N_3580,N_388,N_1409);
xnor U3581 (N_3581,N_752,N_331);
xor U3582 (N_3582,N_442,N_273);
or U3583 (N_3583,N_1202,N_264);
nor U3584 (N_3584,N_1178,N_1021);
or U3585 (N_3585,N_1716,N_191);
nand U3586 (N_3586,N_866,N_1960);
nand U3587 (N_3587,N_1891,N_1655);
or U3588 (N_3588,N_152,N_1239);
nor U3589 (N_3589,N_177,N_1161);
xor U3590 (N_3590,N_833,N_869);
or U3591 (N_3591,N_44,N_317);
nor U3592 (N_3592,N_463,N_1477);
nand U3593 (N_3593,N_1673,N_170);
xor U3594 (N_3594,N_1134,N_584);
nor U3595 (N_3595,N_1147,N_1369);
nand U3596 (N_3596,N_1273,N_1144);
or U3597 (N_3597,N_39,N_19);
xnor U3598 (N_3598,N_774,N_1065);
or U3599 (N_3599,N_516,N_1239);
nand U3600 (N_3600,N_890,N_697);
xnor U3601 (N_3601,N_1641,N_334);
and U3602 (N_3602,N_643,N_839);
or U3603 (N_3603,N_1079,N_1104);
nand U3604 (N_3604,N_1157,N_1667);
nand U3605 (N_3605,N_1724,N_725);
nor U3606 (N_3606,N_1195,N_869);
or U3607 (N_3607,N_1212,N_1160);
nand U3608 (N_3608,N_1424,N_692);
nor U3609 (N_3609,N_1631,N_1943);
xor U3610 (N_3610,N_662,N_790);
and U3611 (N_3611,N_1721,N_1931);
or U3612 (N_3612,N_1956,N_1248);
and U3613 (N_3613,N_1589,N_1844);
or U3614 (N_3614,N_1538,N_651);
xor U3615 (N_3615,N_1622,N_1537);
or U3616 (N_3616,N_1665,N_1431);
xnor U3617 (N_3617,N_1111,N_323);
nor U3618 (N_3618,N_1143,N_1830);
or U3619 (N_3619,N_1281,N_1026);
and U3620 (N_3620,N_1110,N_281);
and U3621 (N_3621,N_1603,N_842);
or U3622 (N_3622,N_633,N_551);
and U3623 (N_3623,N_1756,N_332);
and U3624 (N_3624,N_804,N_461);
xnor U3625 (N_3625,N_1345,N_1755);
nor U3626 (N_3626,N_1371,N_1412);
or U3627 (N_3627,N_1928,N_1440);
and U3628 (N_3628,N_1199,N_881);
or U3629 (N_3629,N_1036,N_1590);
nand U3630 (N_3630,N_1193,N_1404);
nand U3631 (N_3631,N_1993,N_1682);
and U3632 (N_3632,N_367,N_1212);
xor U3633 (N_3633,N_1219,N_183);
xnor U3634 (N_3634,N_1273,N_515);
nor U3635 (N_3635,N_1315,N_1117);
xor U3636 (N_3636,N_1810,N_1912);
or U3637 (N_3637,N_628,N_1413);
nand U3638 (N_3638,N_895,N_1267);
xor U3639 (N_3639,N_1358,N_1103);
xnor U3640 (N_3640,N_1386,N_186);
or U3641 (N_3641,N_1729,N_1050);
or U3642 (N_3642,N_1515,N_959);
nor U3643 (N_3643,N_1391,N_1406);
xnor U3644 (N_3644,N_355,N_1399);
and U3645 (N_3645,N_877,N_1071);
or U3646 (N_3646,N_1328,N_1584);
nor U3647 (N_3647,N_354,N_449);
xor U3648 (N_3648,N_730,N_1124);
or U3649 (N_3649,N_920,N_1522);
nor U3650 (N_3650,N_1048,N_529);
xnor U3651 (N_3651,N_1517,N_1226);
and U3652 (N_3652,N_633,N_1439);
xnor U3653 (N_3653,N_1192,N_1607);
and U3654 (N_3654,N_1165,N_49);
nor U3655 (N_3655,N_1458,N_1920);
and U3656 (N_3656,N_657,N_121);
and U3657 (N_3657,N_1325,N_1665);
and U3658 (N_3658,N_1407,N_1885);
or U3659 (N_3659,N_1917,N_441);
xor U3660 (N_3660,N_1314,N_525);
or U3661 (N_3661,N_1483,N_1101);
and U3662 (N_3662,N_1194,N_889);
nand U3663 (N_3663,N_544,N_1608);
or U3664 (N_3664,N_1224,N_887);
and U3665 (N_3665,N_453,N_1213);
and U3666 (N_3666,N_1058,N_627);
and U3667 (N_3667,N_213,N_496);
xnor U3668 (N_3668,N_1873,N_1666);
xor U3669 (N_3669,N_1679,N_1924);
nand U3670 (N_3670,N_1194,N_1359);
and U3671 (N_3671,N_136,N_1209);
or U3672 (N_3672,N_1206,N_328);
xnor U3673 (N_3673,N_1710,N_907);
or U3674 (N_3674,N_336,N_296);
and U3675 (N_3675,N_391,N_184);
xnor U3676 (N_3676,N_1921,N_1050);
nand U3677 (N_3677,N_1368,N_686);
or U3678 (N_3678,N_1090,N_1914);
nor U3679 (N_3679,N_1686,N_1216);
nor U3680 (N_3680,N_786,N_141);
nor U3681 (N_3681,N_760,N_1959);
and U3682 (N_3682,N_679,N_222);
xor U3683 (N_3683,N_1071,N_1452);
nor U3684 (N_3684,N_657,N_546);
or U3685 (N_3685,N_1293,N_6);
nor U3686 (N_3686,N_1939,N_936);
nor U3687 (N_3687,N_270,N_1136);
xor U3688 (N_3688,N_1445,N_1912);
nand U3689 (N_3689,N_1119,N_803);
or U3690 (N_3690,N_1060,N_1079);
or U3691 (N_3691,N_682,N_1750);
nand U3692 (N_3692,N_723,N_945);
or U3693 (N_3693,N_1795,N_165);
and U3694 (N_3694,N_1923,N_99);
nor U3695 (N_3695,N_912,N_278);
or U3696 (N_3696,N_1972,N_1751);
nor U3697 (N_3697,N_871,N_471);
and U3698 (N_3698,N_122,N_771);
nor U3699 (N_3699,N_1249,N_1789);
nor U3700 (N_3700,N_416,N_545);
or U3701 (N_3701,N_673,N_983);
or U3702 (N_3702,N_1671,N_581);
and U3703 (N_3703,N_1110,N_1185);
xnor U3704 (N_3704,N_112,N_139);
xor U3705 (N_3705,N_1437,N_1403);
nand U3706 (N_3706,N_1682,N_1174);
xnor U3707 (N_3707,N_1030,N_1208);
xnor U3708 (N_3708,N_266,N_473);
nor U3709 (N_3709,N_662,N_1213);
nand U3710 (N_3710,N_681,N_692);
nor U3711 (N_3711,N_1853,N_826);
and U3712 (N_3712,N_1805,N_1913);
or U3713 (N_3713,N_542,N_1151);
nor U3714 (N_3714,N_840,N_1386);
nor U3715 (N_3715,N_759,N_476);
nor U3716 (N_3716,N_1256,N_70);
or U3717 (N_3717,N_1323,N_979);
nor U3718 (N_3718,N_390,N_465);
and U3719 (N_3719,N_1893,N_1671);
and U3720 (N_3720,N_359,N_1563);
nor U3721 (N_3721,N_1029,N_49);
and U3722 (N_3722,N_563,N_487);
xnor U3723 (N_3723,N_916,N_1469);
and U3724 (N_3724,N_793,N_800);
nor U3725 (N_3725,N_1397,N_1166);
nand U3726 (N_3726,N_227,N_1329);
and U3727 (N_3727,N_1463,N_322);
nor U3728 (N_3728,N_132,N_479);
xnor U3729 (N_3729,N_1809,N_314);
or U3730 (N_3730,N_1694,N_1505);
or U3731 (N_3731,N_1633,N_1834);
nor U3732 (N_3732,N_1513,N_726);
nand U3733 (N_3733,N_1593,N_986);
nor U3734 (N_3734,N_1124,N_475);
or U3735 (N_3735,N_1471,N_1783);
or U3736 (N_3736,N_1310,N_1651);
xnor U3737 (N_3737,N_709,N_1188);
xor U3738 (N_3738,N_1773,N_266);
or U3739 (N_3739,N_1980,N_1307);
xnor U3740 (N_3740,N_1420,N_554);
and U3741 (N_3741,N_114,N_905);
or U3742 (N_3742,N_1576,N_351);
or U3743 (N_3743,N_726,N_1155);
nand U3744 (N_3744,N_707,N_168);
and U3745 (N_3745,N_1659,N_1618);
and U3746 (N_3746,N_1800,N_1116);
or U3747 (N_3747,N_5,N_1099);
and U3748 (N_3748,N_1459,N_1330);
and U3749 (N_3749,N_420,N_1284);
or U3750 (N_3750,N_796,N_1794);
nand U3751 (N_3751,N_1294,N_85);
xnor U3752 (N_3752,N_1766,N_991);
xor U3753 (N_3753,N_1942,N_1852);
or U3754 (N_3754,N_1122,N_79);
nand U3755 (N_3755,N_1047,N_1776);
xor U3756 (N_3756,N_1101,N_1741);
nand U3757 (N_3757,N_524,N_369);
xnor U3758 (N_3758,N_1456,N_1661);
nor U3759 (N_3759,N_1582,N_302);
xor U3760 (N_3760,N_1540,N_1517);
nor U3761 (N_3761,N_1940,N_949);
and U3762 (N_3762,N_78,N_13);
and U3763 (N_3763,N_1061,N_391);
and U3764 (N_3764,N_310,N_800);
and U3765 (N_3765,N_1427,N_560);
or U3766 (N_3766,N_1796,N_719);
xor U3767 (N_3767,N_1849,N_771);
nand U3768 (N_3768,N_86,N_284);
or U3769 (N_3769,N_813,N_144);
nor U3770 (N_3770,N_1621,N_160);
and U3771 (N_3771,N_20,N_363);
xor U3772 (N_3772,N_1178,N_802);
or U3773 (N_3773,N_1741,N_1007);
and U3774 (N_3774,N_217,N_1163);
nand U3775 (N_3775,N_1355,N_1119);
xor U3776 (N_3776,N_690,N_1903);
nand U3777 (N_3777,N_1014,N_1786);
or U3778 (N_3778,N_262,N_1502);
nand U3779 (N_3779,N_737,N_798);
nand U3780 (N_3780,N_669,N_995);
or U3781 (N_3781,N_1665,N_1536);
nor U3782 (N_3782,N_1958,N_1244);
nand U3783 (N_3783,N_1417,N_662);
nand U3784 (N_3784,N_796,N_441);
nor U3785 (N_3785,N_1936,N_1177);
nor U3786 (N_3786,N_1770,N_21);
nand U3787 (N_3787,N_1143,N_473);
or U3788 (N_3788,N_1665,N_896);
nand U3789 (N_3789,N_903,N_1105);
or U3790 (N_3790,N_108,N_1536);
xor U3791 (N_3791,N_1037,N_1707);
nand U3792 (N_3792,N_367,N_87);
and U3793 (N_3793,N_1787,N_1629);
nor U3794 (N_3794,N_1247,N_621);
nand U3795 (N_3795,N_700,N_327);
nor U3796 (N_3796,N_932,N_161);
xnor U3797 (N_3797,N_1388,N_725);
and U3798 (N_3798,N_921,N_1462);
xnor U3799 (N_3799,N_1460,N_204);
or U3800 (N_3800,N_1721,N_1403);
and U3801 (N_3801,N_479,N_197);
xnor U3802 (N_3802,N_350,N_1112);
nand U3803 (N_3803,N_192,N_142);
xor U3804 (N_3804,N_778,N_38);
and U3805 (N_3805,N_571,N_23);
or U3806 (N_3806,N_1951,N_369);
or U3807 (N_3807,N_1272,N_321);
xnor U3808 (N_3808,N_819,N_513);
nand U3809 (N_3809,N_307,N_449);
xor U3810 (N_3810,N_883,N_1363);
nand U3811 (N_3811,N_1499,N_1485);
nand U3812 (N_3812,N_1896,N_1794);
nor U3813 (N_3813,N_1256,N_1056);
xnor U3814 (N_3814,N_626,N_14);
xnor U3815 (N_3815,N_1545,N_1768);
xnor U3816 (N_3816,N_689,N_1117);
nor U3817 (N_3817,N_487,N_1001);
nand U3818 (N_3818,N_308,N_1960);
or U3819 (N_3819,N_441,N_1181);
xnor U3820 (N_3820,N_274,N_952);
nand U3821 (N_3821,N_1078,N_1869);
nand U3822 (N_3822,N_927,N_941);
nand U3823 (N_3823,N_1968,N_1054);
nand U3824 (N_3824,N_1262,N_968);
nor U3825 (N_3825,N_253,N_852);
nand U3826 (N_3826,N_765,N_147);
nor U3827 (N_3827,N_450,N_1888);
nand U3828 (N_3828,N_315,N_557);
xor U3829 (N_3829,N_1214,N_1388);
nor U3830 (N_3830,N_1791,N_1820);
nor U3831 (N_3831,N_1649,N_570);
or U3832 (N_3832,N_51,N_1253);
xor U3833 (N_3833,N_1609,N_569);
nand U3834 (N_3834,N_1711,N_440);
nand U3835 (N_3835,N_1958,N_957);
xor U3836 (N_3836,N_1612,N_1590);
xnor U3837 (N_3837,N_1168,N_187);
xnor U3838 (N_3838,N_512,N_135);
nor U3839 (N_3839,N_789,N_806);
xor U3840 (N_3840,N_1218,N_1649);
xor U3841 (N_3841,N_1271,N_936);
nor U3842 (N_3842,N_11,N_1332);
or U3843 (N_3843,N_1054,N_1801);
nor U3844 (N_3844,N_366,N_50);
nand U3845 (N_3845,N_1328,N_570);
or U3846 (N_3846,N_355,N_783);
and U3847 (N_3847,N_1870,N_206);
and U3848 (N_3848,N_800,N_359);
and U3849 (N_3849,N_86,N_1380);
or U3850 (N_3850,N_1719,N_660);
nand U3851 (N_3851,N_661,N_641);
nor U3852 (N_3852,N_1124,N_184);
nor U3853 (N_3853,N_239,N_214);
nor U3854 (N_3854,N_1975,N_466);
nand U3855 (N_3855,N_1332,N_238);
nand U3856 (N_3856,N_1641,N_36);
or U3857 (N_3857,N_1781,N_60);
xnor U3858 (N_3858,N_1208,N_540);
or U3859 (N_3859,N_1995,N_152);
nand U3860 (N_3860,N_836,N_761);
or U3861 (N_3861,N_1821,N_818);
nor U3862 (N_3862,N_701,N_1457);
xor U3863 (N_3863,N_1468,N_685);
xor U3864 (N_3864,N_534,N_101);
nor U3865 (N_3865,N_542,N_183);
and U3866 (N_3866,N_1038,N_1532);
or U3867 (N_3867,N_1430,N_340);
and U3868 (N_3868,N_1161,N_823);
nor U3869 (N_3869,N_447,N_125);
and U3870 (N_3870,N_1546,N_1944);
and U3871 (N_3871,N_1455,N_1913);
xor U3872 (N_3872,N_1314,N_99);
nand U3873 (N_3873,N_1006,N_1222);
xnor U3874 (N_3874,N_1562,N_989);
or U3875 (N_3875,N_1833,N_531);
nor U3876 (N_3876,N_1192,N_384);
or U3877 (N_3877,N_507,N_1824);
xor U3878 (N_3878,N_818,N_791);
xor U3879 (N_3879,N_194,N_877);
or U3880 (N_3880,N_1653,N_1962);
nand U3881 (N_3881,N_17,N_1786);
or U3882 (N_3882,N_6,N_48);
or U3883 (N_3883,N_621,N_1315);
xor U3884 (N_3884,N_1559,N_1897);
nand U3885 (N_3885,N_733,N_258);
and U3886 (N_3886,N_1114,N_577);
xnor U3887 (N_3887,N_1167,N_141);
nor U3888 (N_3888,N_1725,N_56);
or U3889 (N_3889,N_1124,N_1566);
nand U3890 (N_3890,N_1292,N_882);
xnor U3891 (N_3891,N_1462,N_1167);
or U3892 (N_3892,N_159,N_1550);
or U3893 (N_3893,N_540,N_1228);
or U3894 (N_3894,N_641,N_667);
xor U3895 (N_3895,N_1915,N_1968);
or U3896 (N_3896,N_1898,N_1833);
xor U3897 (N_3897,N_1996,N_206);
nor U3898 (N_3898,N_990,N_1551);
nand U3899 (N_3899,N_1233,N_1496);
or U3900 (N_3900,N_231,N_1144);
xnor U3901 (N_3901,N_825,N_18);
and U3902 (N_3902,N_1429,N_1446);
xor U3903 (N_3903,N_376,N_728);
nand U3904 (N_3904,N_412,N_1161);
and U3905 (N_3905,N_1551,N_1402);
xor U3906 (N_3906,N_43,N_778);
nand U3907 (N_3907,N_1094,N_1357);
or U3908 (N_3908,N_1702,N_48);
nand U3909 (N_3909,N_811,N_204);
nor U3910 (N_3910,N_1914,N_671);
nor U3911 (N_3911,N_1905,N_769);
xnor U3912 (N_3912,N_1311,N_1902);
nand U3913 (N_3913,N_166,N_1250);
and U3914 (N_3914,N_891,N_592);
xnor U3915 (N_3915,N_478,N_1175);
xnor U3916 (N_3916,N_1247,N_204);
nor U3917 (N_3917,N_1286,N_1108);
xor U3918 (N_3918,N_1417,N_1685);
or U3919 (N_3919,N_585,N_1252);
and U3920 (N_3920,N_240,N_1576);
nand U3921 (N_3921,N_60,N_1060);
xnor U3922 (N_3922,N_1358,N_1671);
xor U3923 (N_3923,N_231,N_1670);
xor U3924 (N_3924,N_363,N_1366);
and U3925 (N_3925,N_422,N_749);
xnor U3926 (N_3926,N_421,N_153);
or U3927 (N_3927,N_283,N_142);
nand U3928 (N_3928,N_1780,N_450);
and U3929 (N_3929,N_1371,N_1462);
nand U3930 (N_3930,N_681,N_50);
xnor U3931 (N_3931,N_1757,N_61);
nor U3932 (N_3932,N_1798,N_293);
nor U3933 (N_3933,N_1460,N_1347);
nor U3934 (N_3934,N_175,N_1264);
nor U3935 (N_3935,N_1123,N_248);
and U3936 (N_3936,N_660,N_1458);
or U3937 (N_3937,N_805,N_264);
nor U3938 (N_3938,N_1126,N_1764);
nand U3939 (N_3939,N_989,N_319);
or U3940 (N_3940,N_1318,N_1895);
and U3941 (N_3941,N_1434,N_1398);
nor U3942 (N_3942,N_1146,N_519);
nor U3943 (N_3943,N_1129,N_1169);
nand U3944 (N_3944,N_1398,N_169);
nand U3945 (N_3945,N_122,N_1430);
nor U3946 (N_3946,N_1579,N_1269);
nand U3947 (N_3947,N_360,N_543);
or U3948 (N_3948,N_1624,N_18);
nand U3949 (N_3949,N_468,N_842);
nor U3950 (N_3950,N_960,N_1291);
or U3951 (N_3951,N_1349,N_1427);
or U3952 (N_3952,N_784,N_1726);
nand U3953 (N_3953,N_507,N_412);
xnor U3954 (N_3954,N_378,N_729);
nand U3955 (N_3955,N_1928,N_429);
and U3956 (N_3956,N_1614,N_817);
nor U3957 (N_3957,N_1230,N_1297);
xnor U3958 (N_3958,N_807,N_446);
nand U3959 (N_3959,N_504,N_1936);
xnor U3960 (N_3960,N_1678,N_1692);
nor U3961 (N_3961,N_1508,N_84);
xnor U3962 (N_3962,N_120,N_1025);
and U3963 (N_3963,N_591,N_736);
or U3964 (N_3964,N_556,N_679);
xor U3965 (N_3965,N_1420,N_1012);
nand U3966 (N_3966,N_966,N_831);
nor U3967 (N_3967,N_112,N_551);
nor U3968 (N_3968,N_1817,N_743);
nor U3969 (N_3969,N_901,N_1792);
nand U3970 (N_3970,N_1910,N_1177);
nand U3971 (N_3971,N_1311,N_1592);
xnor U3972 (N_3972,N_1139,N_1542);
nand U3973 (N_3973,N_934,N_266);
xnor U3974 (N_3974,N_1727,N_1464);
nand U3975 (N_3975,N_266,N_255);
or U3976 (N_3976,N_620,N_114);
or U3977 (N_3977,N_231,N_1884);
xor U3978 (N_3978,N_636,N_1188);
and U3979 (N_3979,N_1212,N_416);
nand U3980 (N_3980,N_160,N_710);
xor U3981 (N_3981,N_1856,N_234);
or U3982 (N_3982,N_343,N_1003);
nor U3983 (N_3983,N_615,N_266);
nand U3984 (N_3984,N_793,N_557);
or U3985 (N_3985,N_302,N_520);
or U3986 (N_3986,N_1326,N_214);
nand U3987 (N_3987,N_37,N_1259);
or U3988 (N_3988,N_694,N_350);
nand U3989 (N_3989,N_318,N_1282);
xor U3990 (N_3990,N_66,N_1070);
nor U3991 (N_3991,N_819,N_1175);
nand U3992 (N_3992,N_1214,N_191);
nand U3993 (N_3993,N_1295,N_1208);
and U3994 (N_3994,N_189,N_541);
nand U3995 (N_3995,N_1189,N_414);
nor U3996 (N_3996,N_1758,N_583);
and U3997 (N_3997,N_924,N_1488);
nor U3998 (N_3998,N_1366,N_1504);
nor U3999 (N_3999,N_661,N_12);
and U4000 (N_4000,N_3401,N_2803);
or U4001 (N_4001,N_2578,N_3053);
nand U4002 (N_4002,N_2430,N_3506);
xor U4003 (N_4003,N_2846,N_2157);
nand U4004 (N_4004,N_2964,N_3125);
nor U4005 (N_4005,N_2884,N_3021);
nand U4006 (N_4006,N_3067,N_3636);
xor U4007 (N_4007,N_2877,N_2092);
xnor U4008 (N_4008,N_3480,N_3490);
xnor U4009 (N_4009,N_2439,N_2188);
and U4010 (N_4010,N_2571,N_2232);
nor U4011 (N_4011,N_2815,N_2647);
nor U4012 (N_4012,N_2348,N_2245);
nand U4013 (N_4013,N_2498,N_2548);
and U4014 (N_4014,N_3303,N_3664);
nor U4015 (N_4015,N_2648,N_3827);
xnor U4016 (N_4016,N_2804,N_3041);
nand U4017 (N_4017,N_2431,N_3859);
or U4018 (N_4018,N_3049,N_2611);
xor U4019 (N_4019,N_2701,N_3014);
nor U4020 (N_4020,N_3114,N_2851);
nand U4021 (N_4021,N_3946,N_2483);
nor U4022 (N_4022,N_3126,N_3682);
and U4023 (N_4023,N_2110,N_2546);
xor U4024 (N_4024,N_2321,N_3189);
xnor U4025 (N_4025,N_2067,N_3085);
nor U4026 (N_4026,N_3503,N_3860);
nand U4027 (N_4027,N_2264,N_2443);
xor U4028 (N_4028,N_2454,N_3420);
nand U4029 (N_4029,N_3479,N_2784);
or U4030 (N_4030,N_2202,N_3591);
xnor U4031 (N_4031,N_3839,N_3108);
and U4032 (N_4032,N_3246,N_2146);
or U4033 (N_4033,N_3079,N_2458);
nor U4034 (N_4034,N_3528,N_2751);
and U4035 (N_4035,N_3484,N_3803);
and U4036 (N_4036,N_2780,N_3549);
xor U4037 (N_4037,N_3375,N_3144);
nor U4038 (N_4038,N_3317,N_3704);
and U4039 (N_4039,N_3716,N_3386);
and U4040 (N_4040,N_3550,N_2073);
xnor U4041 (N_4041,N_3987,N_2604);
xnor U4042 (N_4042,N_2984,N_2995);
xor U4043 (N_4043,N_3045,N_2520);
nand U4044 (N_4044,N_3133,N_3361);
nor U4045 (N_4045,N_2745,N_2494);
nand U4046 (N_4046,N_2526,N_2470);
and U4047 (N_4047,N_2683,N_3834);
nand U4048 (N_4048,N_2818,N_2510);
nor U4049 (N_4049,N_3651,N_3540);
xnor U4050 (N_4050,N_3618,N_2425);
or U4051 (N_4051,N_3501,N_2136);
nor U4052 (N_4052,N_3134,N_3997);
or U4053 (N_4053,N_2983,N_2326);
nand U4054 (N_4054,N_2918,N_2887);
or U4055 (N_4055,N_2435,N_2889);
or U4056 (N_4056,N_2120,N_2222);
nor U4057 (N_4057,N_3828,N_3790);
xnor U4058 (N_4058,N_3263,N_3287);
nand U4059 (N_4059,N_3293,N_2580);
and U4060 (N_4060,N_3387,N_3989);
nand U4061 (N_4061,N_2457,N_2640);
or U4062 (N_4062,N_2852,N_2947);
nor U4063 (N_4063,N_2065,N_3445);
xnor U4064 (N_4064,N_2069,N_2699);
or U4065 (N_4065,N_3695,N_2729);
and U4066 (N_4066,N_3260,N_3933);
or U4067 (N_4067,N_3944,N_2821);
nor U4068 (N_4068,N_2644,N_2697);
xor U4069 (N_4069,N_3015,N_3917);
nand U4070 (N_4070,N_2968,N_3872);
xor U4071 (N_4071,N_2128,N_2632);
xor U4072 (N_4072,N_3782,N_3147);
xnor U4073 (N_4073,N_3368,N_2527);
or U4074 (N_4074,N_3336,N_2933);
nand U4075 (N_4075,N_2709,N_2035);
or U4076 (N_4076,N_3269,N_3177);
nand U4077 (N_4077,N_2170,N_2047);
nand U4078 (N_4078,N_3635,N_2779);
xor U4079 (N_4079,N_3692,N_3927);
xnor U4080 (N_4080,N_3493,N_3883);
nor U4081 (N_4081,N_2456,N_2667);
and U4082 (N_4082,N_3697,N_3814);
nor U4083 (N_4083,N_3728,N_3504);
xnor U4084 (N_4084,N_2337,N_3072);
nor U4085 (N_4085,N_3237,N_3005);
or U4086 (N_4086,N_2684,N_2738);
nor U4087 (N_4087,N_3693,N_3849);
nand U4088 (N_4088,N_3775,N_3888);
nor U4089 (N_4089,N_2545,N_2369);
nand U4090 (N_4090,N_2340,N_2514);
nor U4091 (N_4091,N_2599,N_3345);
and U4092 (N_4092,N_2936,N_2014);
nor U4093 (N_4093,N_3453,N_2086);
nor U4094 (N_4094,N_2612,N_3720);
xnor U4095 (N_4095,N_3901,N_3390);
or U4096 (N_4096,N_2842,N_2975);
or U4097 (N_4097,N_2841,N_2763);
and U4098 (N_4098,N_3384,N_3877);
and U4099 (N_4099,N_3907,N_3809);
and U4100 (N_4100,N_3095,N_2433);
nor U4101 (N_4101,N_3857,N_3261);
or U4102 (N_4102,N_2614,N_3936);
or U4103 (N_4103,N_2140,N_3127);
and U4104 (N_4104,N_2346,N_2728);
and U4105 (N_4105,N_3753,N_3942);
xor U4106 (N_4106,N_3296,N_3130);
xor U4107 (N_4107,N_3934,N_3898);
xor U4108 (N_4108,N_3574,N_2270);
xnor U4109 (N_4109,N_3110,N_2972);
nor U4110 (N_4110,N_2316,N_2556);
and U4111 (N_4111,N_2799,N_3982);
nand U4112 (N_4112,N_3205,N_3713);
nand U4113 (N_4113,N_3895,N_2777);
nand U4114 (N_4114,N_2859,N_2950);
and U4115 (N_4115,N_2455,N_3525);
nor U4116 (N_4116,N_3090,N_2523);
nor U4117 (N_4117,N_3688,N_3176);
nand U4118 (N_4118,N_3168,N_3197);
xor U4119 (N_4119,N_2398,N_3924);
or U4120 (N_4120,N_3326,N_2323);
nor U4121 (N_4121,N_3832,N_3033);
or U4122 (N_4122,N_2331,N_2334);
and U4123 (N_4123,N_2702,N_2001);
or U4124 (N_4124,N_3173,N_2583);
nor U4125 (N_4125,N_2080,N_3430);
and U4126 (N_4126,N_3031,N_2265);
xnor U4127 (N_4127,N_2093,N_3150);
or U4128 (N_4128,N_2218,N_3351);
and U4129 (N_4129,N_3109,N_3171);
nor U4130 (N_4130,N_3707,N_2186);
nand U4131 (N_4131,N_2797,N_3265);
nand U4132 (N_4132,N_2078,N_3084);
and U4133 (N_4133,N_2289,N_3210);
or U4134 (N_4134,N_3628,N_2707);
and U4135 (N_4135,N_2206,N_2999);
nand U4136 (N_4136,N_2113,N_2967);
nor U4137 (N_4137,N_2448,N_2676);
and U4138 (N_4138,N_2848,N_2282);
and U4139 (N_4139,N_2541,N_3402);
nand U4140 (N_4140,N_2630,N_2229);
or U4141 (N_4141,N_2085,N_3904);
or U4142 (N_4142,N_2938,N_3039);
nand U4143 (N_4143,N_3137,N_3494);
nor U4144 (N_4144,N_3873,N_2150);
xnor U4145 (N_4145,N_2307,N_3449);
or U4146 (N_4146,N_3411,N_2173);
and U4147 (N_4147,N_2244,N_3773);
or U4148 (N_4148,N_3458,N_2782);
xnor U4149 (N_4149,N_3481,N_3091);
and U4150 (N_4150,N_2932,N_3460);
and U4151 (N_4151,N_2725,N_2072);
xor U4152 (N_4152,N_2695,N_2847);
nand U4153 (N_4153,N_3363,N_2872);
nand U4154 (N_4154,N_3755,N_2063);
or U4155 (N_4155,N_3560,N_2060);
nor U4156 (N_4156,N_2377,N_3365);
and U4157 (N_4157,N_3209,N_3925);
nand U4158 (N_4158,N_3649,N_2646);
nor U4159 (N_4159,N_2205,N_3185);
xor U4160 (N_4160,N_2837,N_2260);
or U4161 (N_4161,N_2518,N_3149);
nand U4162 (N_4162,N_3155,N_3588);
nor U4163 (N_4163,N_2033,N_2434);
xor U4164 (N_4164,N_3040,N_3739);
nor U4165 (N_4165,N_2084,N_3370);
nor U4166 (N_4166,N_3940,N_2594);
nand U4167 (N_4167,N_2502,N_2896);
nand U4168 (N_4168,N_2207,N_2749);
nand U4169 (N_4169,N_2391,N_2905);
nor U4170 (N_4170,N_3663,N_2511);
nor U4171 (N_4171,N_3271,N_2241);
xor U4172 (N_4172,N_3097,N_3615);
and U4173 (N_4173,N_3322,N_2744);
and U4174 (N_4174,N_3554,N_2512);
nand U4175 (N_4175,N_2558,N_2164);
nand U4176 (N_4176,N_3212,N_3333);
nor U4177 (N_4177,N_2094,N_2517);
nand U4178 (N_4178,N_3879,N_2243);
or U4179 (N_4179,N_3026,N_2951);
nand U4180 (N_4180,N_2757,N_3561);
xor U4181 (N_4181,N_3448,N_2703);
xnor U4182 (N_4182,N_3641,N_2655);
nand U4183 (N_4183,N_3511,N_3488);
or U4184 (N_4184,N_2990,N_2131);
xor U4185 (N_4185,N_3037,N_3431);
xnor U4186 (N_4186,N_2902,N_2184);
nand U4187 (N_4187,N_2592,N_3829);
xnor U4188 (N_4188,N_2772,N_2192);
nor U4189 (N_4189,N_3714,N_2867);
nor U4190 (N_4190,N_3413,N_2774);
xnor U4191 (N_4191,N_3225,N_2389);
xor U4192 (N_4192,N_3586,N_3964);
or U4193 (N_4193,N_2500,N_3359);
nor U4194 (N_4194,N_2183,N_3699);
nand U4195 (N_4195,N_2906,N_2343);
or U4196 (N_4196,N_2758,N_3616);
xor U4197 (N_4197,N_2026,N_3227);
or U4198 (N_4198,N_3966,N_2269);
nor U4199 (N_4199,N_3062,N_2978);
nand U4200 (N_4200,N_3056,N_3065);
nor U4201 (N_4201,N_2096,N_3558);
nor U4202 (N_4202,N_2166,N_2004);
and U4203 (N_4203,N_3017,N_3280);
xor U4204 (N_4204,N_2690,N_3406);
nor U4205 (N_4205,N_3242,N_2620);
or U4206 (N_4206,N_3585,N_2428);
nor U4207 (N_4207,N_3519,N_2020);
nor U4208 (N_4208,N_2883,N_3186);
and U4209 (N_4209,N_3949,N_3043);
xnor U4210 (N_4210,N_2602,N_2634);
and U4211 (N_4211,N_3107,N_2373);
or U4212 (N_4212,N_3566,N_3310);
xor U4213 (N_4213,N_2165,N_2567);
nand U4214 (N_4214,N_2252,N_3443);
nand U4215 (N_4215,N_2739,N_2145);
and U4216 (N_4216,N_3959,N_3148);
nor U4217 (N_4217,N_2985,N_3187);
xnor U4218 (N_4218,N_3643,N_2149);
or U4219 (N_4219,N_3258,N_3248);
and U4220 (N_4220,N_2625,N_3824);
xor U4221 (N_4221,N_2721,N_2045);
nand U4222 (N_4222,N_2616,N_3767);
or U4223 (N_4223,N_2402,N_3512);
or U4224 (N_4224,N_2897,N_2813);
or U4225 (N_4225,N_3305,N_3470);
nand U4226 (N_4226,N_3820,N_2475);
and U4227 (N_4227,N_2608,N_2360);
or U4228 (N_4228,N_3590,N_3247);
and U4229 (N_4229,N_2862,N_2037);
nor U4230 (N_4230,N_2296,N_3852);
or U4231 (N_4231,N_3668,N_2687);
xor U4232 (N_4232,N_3250,N_3798);
nand U4233 (N_4233,N_3234,N_3658);
nand U4234 (N_4234,N_2006,N_3099);
or U4235 (N_4235,N_2624,N_2319);
xor U4236 (N_4236,N_3462,N_2327);
nand U4237 (N_4237,N_2794,N_3805);
nor U4238 (N_4238,N_2816,N_3734);
or U4239 (N_4239,N_3853,N_2935);
nor U4240 (N_4240,N_2099,N_3123);
nor U4241 (N_4241,N_3815,N_2062);
nand U4242 (N_4242,N_2419,N_2079);
xor U4243 (N_4243,N_3662,N_3776);
and U4244 (N_4244,N_2759,N_2970);
xor U4245 (N_4245,N_2529,N_2503);
nand U4246 (N_4246,N_3657,N_2349);
nor U4247 (N_4247,N_2266,N_3266);
nand U4248 (N_4248,N_3429,N_3241);
nand U4249 (N_4249,N_3508,N_2781);
or U4250 (N_4250,N_3471,N_3701);
nand U4251 (N_4251,N_2288,N_3948);
xnor U4252 (N_4252,N_3995,N_3112);
and U4253 (N_4253,N_3388,N_3821);
or U4254 (N_4254,N_2743,N_3275);
nor U4255 (N_4255,N_3098,N_2141);
nand U4256 (N_4256,N_3800,N_2314);
and U4257 (N_4257,N_3432,N_2581);
nor U4258 (N_4258,N_2176,N_3403);
or U4259 (N_4259,N_3028,N_3956);
and U4260 (N_4260,N_2665,N_2808);
nand U4261 (N_4261,N_2607,N_3928);
or U4262 (N_4262,N_2521,N_2250);
or U4263 (N_4263,N_3335,N_2557);
nand U4264 (N_4264,N_2524,N_2054);
xnor U4265 (N_4265,N_3178,N_2290);
nor U4266 (N_4266,N_2027,N_3788);
nor U4267 (N_4267,N_3467,N_2915);
and U4268 (N_4268,N_2203,N_3353);
and U4269 (N_4269,N_3524,N_2538);
or U4270 (N_4270,N_2858,N_2273);
or U4271 (N_4271,N_3954,N_2427);
or U4272 (N_4272,N_3415,N_3138);
and U4273 (N_4273,N_3279,N_2098);
and U4274 (N_4274,N_2497,N_2650);
or U4275 (N_4275,N_2300,N_3224);
nor U4276 (N_4276,N_3219,N_3795);
xor U4277 (N_4277,N_3145,N_2249);
and U4278 (N_4278,N_2645,N_3141);
or U4279 (N_4279,N_3094,N_2301);
or U4280 (N_4280,N_2267,N_3520);
nor U4281 (N_4281,N_3004,N_2764);
nor U4282 (N_4282,N_2585,N_3182);
and U4283 (N_4283,N_3887,N_2432);
and U4284 (N_4284,N_3876,N_2075);
xnor U4285 (N_4285,N_3089,N_3491);
and U4286 (N_4286,N_3906,N_3654);
nor U4287 (N_4287,N_2182,N_3179);
xor U4288 (N_4288,N_2766,N_2801);
and U4289 (N_4289,N_3745,N_2168);
xor U4290 (N_4290,N_3121,N_3850);
nand U4291 (N_4291,N_3536,N_3496);
and U4292 (N_4292,N_3772,N_2187);
xor U4293 (N_4293,N_2181,N_2417);
nand U4294 (N_4294,N_3529,N_3742);
or U4295 (N_4295,N_3796,N_3162);
nor U4296 (N_4296,N_2677,N_2765);
xnor U4297 (N_4297,N_2942,N_3958);
xnor U4298 (N_4298,N_3301,N_2750);
and U4299 (N_4299,N_2733,N_3607);
xnor U4300 (N_4300,N_2394,N_3077);
nand U4301 (N_4301,N_2390,N_3088);
nand U4302 (N_4302,N_2835,N_3507);
nor U4303 (N_4303,N_2226,N_2582);
and U4304 (N_4304,N_3215,N_3660);
xnor U4305 (N_4305,N_3639,N_2212);
nor U4306 (N_4306,N_3486,N_3671);
xor U4307 (N_4307,N_2961,N_2597);
nand U4308 (N_4308,N_2540,N_2937);
xnor U4309 (N_4309,N_3295,N_3913);
nor U4310 (N_4310,N_2383,N_3256);
nand U4311 (N_4311,N_2871,N_2934);
and U4312 (N_4312,N_3223,N_3882);
nand U4313 (N_4313,N_3547,N_3749);
and U4314 (N_4314,N_3836,N_3063);
and U4315 (N_4315,N_3765,N_3578);
or U4316 (N_4316,N_3804,N_3139);
or U4317 (N_4317,N_2482,N_3841);
xnor U4318 (N_4318,N_2991,N_2798);
and U4319 (N_4319,N_2253,N_3546);
and U4320 (N_4320,N_2275,N_2753);
and U4321 (N_4321,N_3947,N_2901);
nor U4322 (N_4322,N_3309,N_2834);
nor U4323 (N_4323,N_3597,N_2124);
nand U4324 (N_4324,N_2572,N_3249);
xor U4325 (N_4325,N_2303,N_3835);
nand U4326 (N_4326,N_2949,N_2324);
nand U4327 (N_4327,N_2351,N_3854);
or U4328 (N_4328,N_2863,N_2643);
nand U4329 (N_4329,N_3397,N_3457);
xor U4330 (N_4330,N_3357,N_2076);
nor U4331 (N_4331,N_2022,N_2484);
and U4332 (N_4332,N_3622,N_3569);
xnor U4333 (N_4333,N_2663,N_3802);
xor U4334 (N_4334,N_3096,N_3344);
nor U4335 (N_4335,N_2587,N_3381);
or U4336 (N_4336,N_2486,N_2742);
or U4337 (N_4337,N_2588,N_2230);
or U4338 (N_4338,N_2603,N_2686);
nand U4339 (N_4339,N_3347,N_2513);
xor U4340 (N_4340,N_3659,N_3777);
nand U4341 (N_4341,N_3489,N_2706);
or U4342 (N_4342,N_2057,N_2393);
nor U4343 (N_4343,N_2345,N_2447);
nor U4344 (N_4344,N_3427,N_3456);
or U4345 (N_4345,N_2409,N_2998);
nand U4346 (N_4346,N_3086,N_2297);
nand U4347 (N_4347,N_2771,N_3153);
or U4348 (N_4348,N_3637,N_2410);
or U4349 (N_4349,N_2473,N_3408);
nand U4350 (N_4350,N_2059,N_2566);
nand U4351 (N_4351,N_2962,N_3999);
and U4352 (N_4352,N_2910,N_3196);
or U4353 (N_4353,N_2441,N_3025);
nor U4354 (N_4354,N_3230,N_3410);
nor U4355 (N_4355,N_2444,N_2095);
nor U4356 (N_4356,N_2672,N_3372);
nand U4357 (N_4357,N_2106,N_2864);
xnor U4358 (N_4358,N_3497,N_2921);
nor U4359 (N_4359,N_2914,N_3579);
nand U4360 (N_4360,N_2235,N_3444);
and U4361 (N_4361,N_3629,N_2944);
and U4362 (N_4362,N_3619,N_3181);
or U4363 (N_4363,N_2237,N_3527);
and U4364 (N_4364,N_3421,N_2913);
xor U4365 (N_4365,N_2704,N_3042);
nand U4366 (N_4366,N_2421,N_2948);
xnor U4367 (N_4367,N_2287,N_3848);
nand U4368 (N_4368,N_2822,N_2617);
nor U4369 (N_4369,N_2380,N_3012);
nor U4370 (N_4370,N_3104,N_2652);
nand U4371 (N_4371,N_3455,N_2108);
and U4372 (N_4372,N_3424,N_3568);
or U4373 (N_4373,N_3758,N_2474);
or U4374 (N_4374,N_2776,N_3981);
nand U4375 (N_4375,N_2722,N_3594);
nand U4376 (N_4376,N_2416,N_3653);
nor U4377 (N_4377,N_3239,N_2216);
nand U4378 (N_4378,N_2280,N_3143);
nor U4379 (N_4379,N_3548,N_2878);
nand U4380 (N_4380,N_2525,N_2680);
nor U4381 (N_4381,N_2401,N_2870);
nor U4382 (N_4382,N_2268,N_2274);
or U4383 (N_4383,N_2584,N_2112);
xnor U4384 (N_4384,N_3447,N_2016);
or U4385 (N_4385,N_2693,N_3975);
nor U4386 (N_4386,N_3757,N_3433);
nand U4387 (N_4387,N_3195,N_3953);
xor U4388 (N_4388,N_2081,N_3346);
xor U4389 (N_4389,N_3926,N_2442);
nand U4390 (N_4390,N_3101,N_3087);
or U4391 (N_4391,N_3052,N_3294);
nor U4392 (N_4392,N_3010,N_3469);
nand U4393 (N_4393,N_3977,N_2760);
xor U4394 (N_4394,N_3786,N_3608);
xnor U4395 (N_4395,N_2819,N_2853);
xor U4396 (N_4396,N_3683,N_2626);
and U4397 (N_4397,N_3499,N_2681);
and U4398 (N_4398,N_2692,N_2362);
xor U4399 (N_4399,N_2281,N_2609);
xnor U4400 (N_4400,N_2762,N_3330);
or U4401 (N_4401,N_2860,N_3845);
xor U4402 (N_4402,N_3535,N_3166);
or U4403 (N_4403,N_2214,N_2152);
nand U4404 (N_4404,N_2365,N_3756);
and U4405 (N_4405,N_3793,N_2668);
and U4406 (N_4406,N_3685,N_3779);
or U4407 (N_4407,N_2775,N_3277);
or U4408 (N_4408,N_2976,N_2796);
or U4409 (N_4409,N_3816,N_3575);
nand U4410 (N_4410,N_3694,N_3071);
and U4411 (N_4411,N_2489,N_2811);
xnor U4412 (N_4412,N_3655,N_3932);
nor U4413 (N_4413,N_2589,N_3899);
nand U4414 (N_4414,N_2234,N_3875);
nor U4415 (N_4415,N_3703,N_2028);
and U4416 (N_4416,N_2143,N_2137);
or U4417 (N_4417,N_2255,N_3702);
nor U4418 (N_4418,N_2988,N_2213);
nor U4419 (N_4419,N_2747,N_2658);
nor U4420 (N_4420,N_3285,N_2077);
or U4421 (N_4421,N_2082,N_2973);
nand U4422 (N_4422,N_2411,N_2941);
or U4423 (N_4423,N_3632,N_2940);
xnor U4424 (N_4424,N_3656,N_2685);
xor U4425 (N_4425,N_3863,N_3487);
or U4426 (N_4426,N_2987,N_2159);
nand U4427 (N_4427,N_3730,N_3044);
nor U4428 (N_4428,N_2403,N_3909);
or U4429 (N_4429,N_2189,N_2151);
xor U4430 (N_4430,N_3349,N_2283);
xor U4431 (N_4431,N_2515,N_2087);
nor U4432 (N_4432,N_3624,N_3510);
nand U4433 (N_4433,N_2516,N_3232);
and U4434 (N_4434,N_3438,N_3170);
nand U4435 (N_4435,N_3961,N_2126);
nor U4436 (N_4436,N_2109,N_2310);
and U4437 (N_4437,N_2012,N_3286);
and U4438 (N_4438,N_2412,N_2056);
and U4439 (N_4439,N_3640,N_2649);
and U4440 (N_4440,N_2317,N_2298);
nor U4441 (N_4441,N_2735,N_3823);
and U4442 (N_4442,N_3289,N_2844);
nand U4443 (N_4443,N_3951,N_3567);
xnor U4444 (N_4444,N_2927,N_2277);
nand U4445 (N_4445,N_2008,N_2386);
nand U4446 (N_4446,N_3665,N_3360);
or U4447 (N_4447,N_3319,N_2633);
xnor U4448 (N_4448,N_2736,N_3416);
or U4449 (N_4449,N_2036,N_3348);
and U4450 (N_4450,N_2487,N_3874);
and U4451 (N_4451,N_3825,N_3589);
or U4452 (N_4452,N_2179,N_2734);
and U4453 (N_4453,N_2946,N_2138);
nor U4454 (N_4454,N_2271,N_3818);
xor U4455 (N_4455,N_3962,N_3473);
or U4456 (N_4456,N_3032,N_3020);
and U4457 (N_4457,N_2127,N_2619);
and U4458 (N_4458,N_3157,N_2342);
and U4459 (N_4459,N_2424,N_3395);
xnor U4460 (N_4460,N_2825,N_3255);
and U4461 (N_4461,N_2392,N_3974);
nand U4462 (N_4462,N_2537,N_2261);
nor U4463 (N_4463,N_2278,N_3007);
nor U4464 (N_4464,N_3968,N_3175);
nor U4465 (N_4465,N_2900,N_2160);
nor U4466 (N_4466,N_2909,N_2330);
xor U4467 (N_4467,N_3036,N_2468);
nand U4468 (N_4468,N_3712,N_3744);
nor U4469 (N_4469,N_3931,N_2810);
xor U4470 (N_4470,N_2175,N_3115);
or U4471 (N_4471,N_3680,N_2364);
nand U4472 (N_4472,N_2460,N_3748);
nor U4473 (N_4473,N_2357,N_2038);
nand U4474 (N_4474,N_3016,N_3812);
nor U4475 (N_4475,N_2769,N_2178);
nor U4476 (N_4476,N_3254,N_3791);
and U4477 (N_4477,N_2452,N_3617);
nand U4478 (N_4478,N_2294,N_2162);
nor U4479 (N_4479,N_3355,N_3316);
or U4480 (N_4480,N_3136,N_3935);
xnor U4481 (N_4481,N_2544,N_3035);
xor U4482 (N_4482,N_2097,N_3912);
xnor U4483 (N_4483,N_3477,N_2705);
nand U4484 (N_4484,N_2332,N_2814);
nand U4485 (N_4485,N_3743,N_3038);
and U4486 (N_4486,N_3452,N_2132);
and U4487 (N_4487,N_2845,N_2856);
and U4488 (N_4488,N_3172,N_2730);
or U4489 (N_4489,N_3251,N_2247);
nand U4490 (N_4490,N_2215,N_3866);
xnor U4491 (N_4491,N_3746,N_2122);
or U4492 (N_4492,N_2148,N_2091);
nor U4493 (N_4493,N_2596,N_3978);
nand U4494 (N_4494,N_2700,N_3700);
xor U4495 (N_4495,N_2726,N_2509);
and U4496 (N_4496,N_3274,N_2358);
xnor U4497 (N_4497,N_3612,N_2134);
nor U4498 (N_4498,N_2642,N_3174);
xor U4499 (N_4499,N_2040,N_3572);
nand U4500 (N_4500,N_2211,N_2963);
nand U4501 (N_4501,N_2339,N_3288);
and U4502 (N_4502,N_2675,N_2694);
nand U4503 (N_4503,N_2103,N_2039);
nor U4504 (N_4504,N_3302,N_2133);
nor U4505 (N_4505,N_2501,N_2955);
nand U4506 (N_4506,N_2490,N_2233);
nor U4507 (N_4507,N_2083,N_3270);
nand U4508 (N_4508,N_3609,N_2359);
xnor U4509 (N_4509,N_2368,N_3379);
nor U4510 (N_4510,N_2718,N_3783);
xor U4511 (N_4511,N_3583,N_3634);
nand U4512 (N_4512,N_2875,N_3314);
xor U4513 (N_4513,N_2032,N_2719);
nor U4514 (N_4514,N_3321,N_2154);
and U4515 (N_4515,N_2019,N_3690);
or U4516 (N_4516,N_3435,N_3669);
xor U4517 (N_4517,N_2836,N_2220);
or U4518 (N_4518,N_2904,N_3061);
nor U4519 (N_4519,N_2737,N_2768);
and U4520 (N_4520,N_3436,N_3320);
or U4521 (N_4521,N_3910,N_2024);
or U4522 (N_4522,N_2868,N_3723);
nor U4523 (N_4523,N_3941,N_2239);
or U4524 (N_4524,N_2849,N_2741);
nor U4525 (N_4525,N_2259,N_3523);
nor U4526 (N_4526,N_2381,N_3441);
nor U4527 (N_4527,N_3552,N_3516);
xnor U4528 (N_4528,N_2873,N_2208);
and U4529 (N_4529,N_3563,N_2886);
or U4530 (N_4530,N_3204,N_3290);
or U4531 (N_4531,N_3454,N_3377);
nand U4532 (N_4532,N_3582,N_2903);
xnor U4533 (N_4533,N_2881,N_2009);
nand U4534 (N_4534,N_3916,N_2713);
nand U4535 (N_4535,N_2256,N_3509);
nor U4536 (N_4536,N_3792,N_3218);
nand U4537 (N_4537,N_3811,N_3404);
nor U4538 (N_4538,N_2400,N_3394);
or U4539 (N_4539,N_2329,N_3750);
nand U4540 (N_4540,N_2285,N_3761);
or U4541 (N_4541,N_3240,N_3214);
nand U4542 (N_4542,N_3472,N_2792);
and U4543 (N_4543,N_3216,N_2654);
or U4544 (N_4544,N_3865,N_2171);
and U4545 (N_4545,N_3434,N_2785);
nand U4546 (N_4546,N_3389,N_2002);
xnor U4547 (N_4547,N_2958,N_2174);
nor U4548 (N_4548,N_3323,N_2879);
nor U4549 (N_4549,N_3542,N_3667);
nand U4550 (N_4550,N_2820,N_2943);
and U4551 (N_4551,N_3715,N_3092);
nor U4552 (N_4552,N_2313,N_3885);
and U4553 (N_4553,N_3760,N_3869);
nor U4554 (N_4554,N_3190,N_3681);
or U4555 (N_4555,N_2636,N_2552);
nand U4556 (N_4556,N_2418,N_2341);
and U4557 (N_4557,N_3485,N_2451);
xor U4558 (N_4558,N_2013,N_3847);
or U4559 (N_4559,N_3054,N_2445);
or U4560 (N_4560,N_3778,N_2590);
xor U4561 (N_4561,N_3238,N_3521);
or U4562 (N_4562,N_3268,N_3362);
nor U4563 (N_4563,N_2440,N_3596);
xnor U4564 (N_4564,N_3437,N_2894);
xor U4565 (N_4565,N_2015,N_3192);
or U4566 (N_4566,N_2191,N_3896);
or U4567 (N_4567,N_3000,N_2347);
nor U4568 (N_4568,N_2052,N_2003);
or U4569 (N_4569,N_2917,N_3708);
or U4570 (N_4570,N_3211,N_2574);
nor U4571 (N_4571,N_3526,N_3500);
and U4572 (N_4572,N_2217,N_2299);
nor U4573 (N_4573,N_3337,N_3220);
or U4574 (N_4574,N_3605,N_3930);
xnor U4575 (N_4575,N_2854,N_3281);
nor U4576 (N_4576,N_2420,N_2046);
xor U4577 (N_4577,N_3893,N_3180);
nor U4578 (N_4578,N_3794,N_3915);
nor U4579 (N_4579,N_2292,N_2561);
and U4580 (N_4580,N_3724,N_3644);
xor U4581 (N_4581,N_2049,N_2591);
and U4582 (N_4582,N_2459,N_3291);
nor U4583 (N_4583,N_2831,N_2279);
or U4584 (N_4584,N_3614,N_2387);
nand U4585 (N_4585,N_2336,N_3638);
or U4586 (N_4586,N_2029,N_3008);
nand U4587 (N_4587,N_3856,N_3556);
and U4588 (N_4588,N_3952,N_2531);
or U4589 (N_4589,N_2823,N_3705);
nor U4590 (N_4590,N_3955,N_3019);
or U4591 (N_4591,N_2125,N_3741);
and U4592 (N_4592,N_3601,N_2320);
or U4593 (N_4593,N_2481,N_2050);
and U4594 (N_4594,N_3851,N_3376);
xor U4595 (N_4595,N_2928,N_3003);
and U4596 (N_4596,N_2564,N_2070);
nor U4597 (N_4597,N_3297,N_3001);
nand U4598 (N_4598,N_3459,N_3892);
nor U4599 (N_4599,N_3980,N_2472);
xnor U4600 (N_4600,N_2671,N_3029);
and U4601 (N_4601,N_3562,N_3891);
nor U4602 (N_4602,N_3201,N_3013);
nor U4603 (N_4603,N_2257,N_2492);
xnor U4604 (N_4604,N_2506,N_3996);
nor U4605 (N_4605,N_3979,N_2708);
nor U4606 (N_4606,N_3264,N_2827);
and U4607 (N_4607,N_2374,N_2673);
nand U4608 (N_4608,N_3217,N_3352);
or U4609 (N_4609,N_3844,N_2464);
xor U4610 (N_4610,N_2892,N_3156);
nand U4611 (N_4611,N_3630,N_3709);
and U4612 (N_4612,N_2196,N_3120);
xnor U4613 (N_4613,N_2375,N_2715);
and U4614 (N_4614,N_2338,N_3731);
and U4615 (N_4615,N_2674,N_2710);
or U4616 (N_4616,N_2974,N_2156);
or U4617 (N_4617,N_3862,N_3324);
or U4618 (N_4618,N_2491,N_3371);
and U4619 (N_4619,N_3861,N_2669);
or U4620 (N_4620,N_2577,N_3300);
nand U4621 (N_4621,N_3645,N_3676);
xor U4622 (N_4622,N_2712,N_3082);
and U4623 (N_4623,N_3078,N_3600);
nor U4624 (N_4624,N_2723,N_2994);
and U4625 (N_4625,N_2058,N_2167);
nor U4626 (N_4626,N_2861,N_2388);
nand U4627 (N_4627,N_2788,N_2829);
xnor U4628 (N_4628,N_2982,N_3838);
and U4629 (N_4629,N_3598,N_2479);
xor U4630 (N_4630,N_3897,N_3327);
xnor U4631 (N_4631,N_3972,N_2068);
xor U4632 (N_4632,N_3921,N_3328);
and U4633 (N_4633,N_2600,N_2601);
nor U4634 (N_4634,N_3950,N_3988);
nand U4635 (N_4635,N_2399,N_2147);
or U4636 (N_4636,N_3855,N_3559);
or U4637 (N_4637,N_3945,N_2807);
and U4638 (N_4638,N_2885,N_3100);
and U4639 (N_4639,N_3817,N_3564);
and U4640 (N_4640,N_3830,N_2787);
or U4641 (N_4641,N_3604,N_2965);
and U4642 (N_4642,N_2325,N_2959);
xnor U4643 (N_4643,N_3518,N_2610);
xnor U4644 (N_4644,N_3023,N_3119);
nor U4645 (N_4645,N_3116,N_2924);
nor U4646 (N_4646,N_3339,N_3439);
nor U4647 (N_4647,N_3414,N_2504);
or U4648 (N_4648,N_3729,N_3957);
nand U4649 (N_4649,N_3378,N_3325);
nor U4650 (N_4650,N_2437,N_3551);
or U4651 (N_4651,N_2793,N_3674);
xor U4652 (N_4652,N_3678,N_3846);
xor U4653 (N_4653,N_2312,N_3132);
nor U4654 (N_4654,N_3048,N_2088);
xnor U4655 (N_4655,N_3725,N_3272);
nand U4656 (N_4656,N_2144,N_2406);
nor U4657 (N_4657,N_3199,N_3160);
nor U4658 (N_4658,N_3687,N_2724);
nor U4659 (N_4659,N_2866,N_3152);
or U4660 (N_4660,N_3446,N_2480);
and U4661 (N_4661,N_2221,N_3581);
nor U4662 (N_4662,N_2929,N_2493);
xor U4663 (N_4663,N_2201,N_3131);
nor U4664 (N_4664,N_2539,N_3252);
and U4665 (N_4665,N_2989,N_3024);
nand U4666 (N_4666,N_3733,N_2931);
nor U4667 (N_4667,N_2055,N_2030);
and U4668 (N_4668,N_3412,N_2240);
nor U4669 (N_4669,N_2641,N_2446);
nand U4670 (N_4670,N_2551,N_2865);
nand U4671 (N_4671,N_2135,N_3027);
nand U4672 (N_4672,N_3299,N_2956);
and U4673 (N_4673,N_2767,N_3369);
or U4674 (N_4674,N_2254,N_2074);
xnor U4675 (N_4675,N_2010,N_2363);
or U4676 (N_4676,N_3183,N_2308);
xnor U4677 (N_4677,N_2850,N_3164);
nor U4678 (N_4678,N_2395,N_3919);
nor U4679 (N_4679,N_2017,N_3530);
and U4680 (N_4680,N_2238,N_3986);
and U4681 (N_4681,N_3534,N_2372);
or U4682 (N_4682,N_2121,N_3881);
nand U4683 (N_4683,N_3736,N_3474);
or U4684 (N_4684,N_2107,N_2408);
nand U4685 (N_4685,N_3030,N_2790);
and U4686 (N_4686,N_2882,N_3880);
nor U4687 (N_4687,N_2618,N_2051);
xnor U4688 (N_4688,N_3442,N_2678);
nand U4689 (N_4689,N_2284,N_3801);
xnor U4690 (N_4690,N_2912,N_2089);
or U4691 (N_4691,N_3009,N_3193);
nor U4692 (N_4692,N_3533,N_3960);
nor U4693 (N_4693,N_2463,N_3400);
and U4694 (N_4694,N_3806,N_3482);
and U4695 (N_4695,N_3329,N_3018);
xnor U4696 (N_4696,N_3111,N_3532);
nand U4697 (N_4697,N_3650,N_3647);
xor U4698 (N_4698,N_3341,N_2554);
nand U4699 (N_4699,N_3226,N_3884);
nor U4700 (N_4700,N_2895,N_2100);
and U4701 (N_4701,N_2286,N_2530);
nand U4702 (N_4702,N_3244,N_2370);
xor U4703 (N_4703,N_2945,N_2670);
nand U4704 (N_4704,N_2857,N_2682);
and U4705 (N_4705,N_2800,N_3576);
xor U4706 (N_4706,N_3331,N_2828);
xor U4707 (N_4707,N_2485,N_2429);
nand U4708 (N_4708,N_3113,N_2465);
nor U4709 (N_4709,N_2996,N_2657);
or U4710 (N_4710,N_2809,N_2977);
and U4711 (N_4711,N_3050,N_3356);
xor U4712 (N_4712,N_2880,N_3383);
xnor U4713 (N_4713,N_3398,N_3905);
nand U4714 (N_4714,N_3198,N_3080);
or U4715 (N_4715,N_3666,N_3990);
nand U4716 (N_4716,N_2615,N_3517);
or U4717 (N_4717,N_3840,N_2021);
nand U4718 (N_4718,N_3165,N_2462);
and U4719 (N_4719,N_3184,N_2622);
nand U4720 (N_4720,N_3633,N_3373);
or U4721 (N_4721,N_3573,N_2114);
xor U4722 (N_4722,N_2204,N_2893);
or U4723 (N_4723,N_3762,N_2276);
and U4724 (N_4724,N_2005,N_2379);
and U4725 (N_4725,N_3939,N_3732);
or U4726 (N_4726,N_2385,N_3603);
nand U4727 (N_4727,N_2534,N_2659);
nor U4728 (N_4728,N_2414,N_3466);
nand U4729 (N_4729,N_2595,N_2662);
or U4730 (N_4730,N_2139,N_3235);
or U4731 (N_4731,N_3706,N_3992);
xor U4732 (N_4732,N_3991,N_3652);
and U4733 (N_4733,N_3229,N_3450);
nand U4734 (N_4734,N_3461,N_2223);
nand U4735 (N_4735,N_2923,N_2352);
nand U4736 (N_4736,N_3418,N_3068);
or U4737 (N_4737,N_2773,N_2248);
and U4738 (N_4738,N_2130,N_2888);
and U4739 (N_4739,N_3727,N_3399);
or U4740 (N_4740,N_3721,N_2158);
xnor U4741 (N_4741,N_3200,N_2717);
and U4742 (N_4742,N_3083,N_3231);
and U4743 (N_4743,N_2007,N_2210);
nand U4744 (N_4744,N_2404,N_3595);
and U4745 (N_4745,N_3698,N_3691);
and U4746 (N_4746,N_2382,N_3868);
nor U4747 (N_4747,N_3864,N_2031);
or U4748 (N_4748,N_2505,N_2071);
and U4749 (N_4749,N_2560,N_2466);
or U4750 (N_4750,N_3914,N_2916);
nand U4751 (N_4751,N_3539,N_3871);
or U4752 (N_4752,N_3154,N_2064);
xnor U4753 (N_4753,N_3476,N_2679);
xnor U4754 (N_4754,N_3545,N_2770);
and U4755 (N_4755,N_3451,N_3074);
nand U4756 (N_4756,N_3315,N_2553);
or U4757 (N_4757,N_2405,N_3766);
nand U4758 (N_4758,N_3257,N_3312);
and U4759 (N_4759,N_2315,N_3366);
nand U4760 (N_4760,N_3405,N_3253);
nor U4761 (N_4761,N_2194,N_2025);
nor U4762 (N_4762,N_3826,N_3350);
nor U4763 (N_4763,N_2061,N_3055);
or U4764 (N_4764,N_2090,N_2478);
and U4765 (N_4765,N_3282,N_3970);
nor U4766 (N_4766,N_2041,N_2631);
xor U4767 (N_4767,N_2413,N_3057);
nor U4768 (N_4768,N_3259,N_3059);
nor U4769 (N_4769,N_3502,N_3833);
xnor U4770 (N_4770,N_2740,N_3283);
xor U4771 (N_4771,N_3994,N_3292);
and U4772 (N_4772,N_2101,N_2246);
and U4773 (N_4773,N_2746,N_3677);
and U4774 (N_4774,N_3843,N_3858);
nor U4775 (N_4775,N_3340,N_3738);
or U4776 (N_4776,N_3367,N_3276);
and U4777 (N_4777,N_3675,N_3648);
nand U4778 (N_4778,N_2606,N_3515);
xnor U4779 (N_4779,N_2727,N_3169);
nand U4780 (N_4780,N_3580,N_3969);
and U4781 (N_4781,N_2843,N_2666);
nor U4782 (N_4782,N_3385,N_2251);
and U4783 (N_4783,N_2536,N_3531);
nand U4784 (N_4784,N_3304,N_3831);
and U4785 (N_4785,N_3984,N_3093);
nor U4786 (N_4786,N_2228,N_3722);
nand U4787 (N_4787,N_3122,N_3267);
nor U4788 (N_4788,N_2833,N_2376);
xor U4789 (N_4789,N_3483,N_2922);
nand U4790 (N_4790,N_3513,N_3565);
xnor U4791 (N_4791,N_2605,N_3570);
and U4792 (N_4792,N_2384,N_2543);
or U4793 (N_4793,N_3819,N_2407);
nor U4794 (N_4794,N_3929,N_3354);
or U4795 (N_4795,N_3106,N_2508);
and U4796 (N_4796,N_3407,N_2830);
xor U4797 (N_4797,N_2311,N_3557);
or U4798 (N_4798,N_3419,N_2366);
nand U4799 (N_4799,N_3338,N_3417);
nor U4800 (N_4800,N_2169,N_3543);
and U4801 (N_4801,N_3813,N_2309);
xor U4802 (N_4802,N_2656,N_3606);
and U4803 (N_4803,N_3751,N_3672);
or U4804 (N_4804,N_2789,N_2627);
and U4805 (N_4805,N_2350,N_3425);
or U4806 (N_4806,N_3993,N_3670);
nor U4807 (N_4807,N_3332,N_3673);
or U4808 (N_4808,N_2957,N_3058);
xor U4809 (N_4809,N_3571,N_2302);
xor U4810 (N_4810,N_3047,N_3318);
or U4811 (N_4811,N_2637,N_2356);
xor U4812 (N_4812,N_2532,N_3306);
nor U4813 (N_4813,N_3129,N_2291);
and U4814 (N_4814,N_2477,N_2786);
or U4815 (N_4815,N_2613,N_3142);
and U4816 (N_4816,N_3167,N_2467);
xnor U4817 (N_4817,N_3971,N_2328);
xnor U4818 (N_4818,N_2469,N_3298);
and U4819 (N_4819,N_3918,N_3382);
and U4820 (N_4820,N_2044,N_3696);
xnor U4821 (N_4821,N_3900,N_2190);
nor U4822 (N_4822,N_3752,N_2034);
nor U4823 (N_4823,N_2111,N_3135);
nand U4824 (N_4824,N_2224,N_2986);
nand U4825 (N_4825,N_3621,N_3623);
nor U4826 (N_4826,N_3602,N_3577);
and U4827 (N_4827,N_2305,N_3611);
and U4828 (N_4828,N_3159,N_3492);
nand U4829 (N_4829,N_2570,N_3076);
xnor U4830 (N_4830,N_2397,N_2869);
nand U4831 (N_4831,N_3073,N_2354);
or U4832 (N_4832,N_2195,N_3102);
and U4833 (N_4833,N_2664,N_2731);
nor U4834 (N_4834,N_3207,N_3426);
nor U4835 (N_4835,N_3380,N_2488);
or U4836 (N_4836,N_3105,N_3878);
and U4837 (N_4837,N_3343,N_3051);
xnor U4838 (N_4838,N_2119,N_2979);
and U4839 (N_4839,N_2997,N_3465);
nor U4840 (N_4840,N_3735,N_3726);
or U4841 (N_4841,N_2361,N_2209);
and U4842 (N_4842,N_2198,N_3391);
xnor U4843 (N_4843,N_2550,N_2651);
nand U4844 (N_4844,N_3203,N_3781);
and U4845 (N_4845,N_2118,N_3774);
and U4846 (N_4846,N_3440,N_3464);
nand U4847 (N_4847,N_2102,N_2322);
xnor U4848 (N_4848,N_2898,N_2593);
nor U4849 (N_4849,N_3364,N_3011);
nor U4850 (N_4850,N_3592,N_3075);
xnor U4851 (N_4851,N_3920,N_3938);
or U4852 (N_4852,N_3243,N_3625);
and U4853 (N_4853,N_3422,N_2262);
and U4854 (N_4854,N_3759,N_2911);
xnor U4855 (N_4855,N_2499,N_2011);
nor U4856 (N_4856,N_3837,N_3587);
and U4857 (N_4857,N_3985,N_3151);
or U4858 (N_4858,N_2116,N_2197);
and U4859 (N_4859,N_3768,N_2569);
nor U4860 (N_4860,N_2306,N_2783);
xor U4861 (N_4861,N_3737,N_2528);
and U4862 (N_4862,N_2639,N_3967);
xnor U4863 (N_4863,N_3787,N_3903);
nor U4864 (N_4864,N_3307,N_2225);
nand U4865 (N_4865,N_3902,N_2542);
xor U4866 (N_4866,N_2939,N_3937);
and U4867 (N_4867,N_3771,N_3060);
and U4868 (N_4868,N_3584,N_3228);
nand U4869 (N_4869,N_3889,N_2826);
xor U4870 (N_4870,N_3810,N_2714);
nor U4871 (N_4871,N_3069,N_2471);
and U4872 (N_4872,N_3208,N_3066);
xnor U4873 (N_4873,N_2926,N_3475);
nor U4874 (N_4874,N_3541,N_2438);
and U4875 (N_4875,N_3222,N_2969);
xor U4876 (N_4876,N_3374,N_3593);
nor U4877 (N_4877,N_2344,N_2043);
xor U4878 (N_4878,N_3894,N_2930);
or U4879 (N_4879,N_2199,N_3002);
xor U4880 (N_4880,N_3626,N_3022);
nor U4881 (N_4881,N_2476,N_2754);
xor U4882 (N_4882,N_3423,N_3278);
nand U4883 (N_4883,N_2231,N_2415);
xnor U4884 (N_4884,N_3514,N_2522);
and U4885 (N_4885,N_3555,N_3206);
xor U4886 (N_4886,N_2519,N_2732);
xor U4887 (N_4887,N_3740,N_3717);
xnor U4888 (N_4888,N_3784,N_2272);
nor U4889 (N_4889,N_3785,N_2660);
nor U4890 (N_4890,N_2180,N_3610);
xor U4891 (N_4891,N_2698,N_3613);
nor U4892 (N_4892,N_2163,N_2549);
nor U4893 (N_4893,N_3081,N_2562);
or U4894 (N_4894,N_2422,N_2805);
and U4895 (N_4895,N_2890,N_2689);
xnor U4896 (N_4896,N_3070,N_3599);
nand U4897 (N_4897,N_2547,N_3194);
or U4898 (N_4898,N_2838,N_3923);
nand U4899 (N_4899,N_3191,N_2153);
nor U4900 (N_4900,N_3311,N_2177);
nand U4901 (N_4901,N_2129,N_3334);
xor U4902 (N_4902,N_3468,N_3006);
and U4903 (N_4903,N_3646,N_2586);
xnor U4904 (N_4904,N_3911,N_2185);
or U4905 (N_4905,N_2954,N_2426);
xor U4906 (N_4906,N_2635,N_2142);
and U4907 (N_4907,N_3273,N_2993);
nor U4908 (N_4908,N_3478,N_3789);
xor U4909 (N_4909,N_2755,N_3202);
nor U4910 (N_4910,N_2053,N_3463);
or U4911 (N_4911,N_3963,N_3140);
nand U4912 (N_4912,N_3392,N_2876);
or U4913 (N_4913,N_2691,N_3661);
xnor U4914 (N_4914,N_2333,N_2761);
or U4915 (N_4915,N_2748,N_2752);
nand U4916 (N_4916,N_2623,N_2018);
nor U4917 (N_4917,N_2899,N_2066);
nand U4918 (N_4918,N_2355,N_2396);
and U4919 (N_4919,N_2568,N_3428);
nand U4920 (N_4920,N_3620,N_2453);
nor U4921 (N_4921,N_3908,N_2293);
or U4922 (N_4922,N_2621,N_2802);
nor U4923 (N_4923,N_3245,N_2200);
or U4924 (N_4924,N_3754,N_2628);
nand U4925 (N_4925,N_2778,N_3146);
nor U4926 (N_4926,N_2449,N_3631);
or U4927 (N_4927,N_2123,N_2711);
nand U4928 (N_4928,N_2461,N_3870);
xnor U4929 (N_4929,N_2219,N_2263);
nand U4930 (N_4930,N_3495,N_2000);
nand U4931 (N_4931,N_2840,N_3358);
and U4932 (N_4932,N_2318,N_2371);
nor U4933 (N_4933,N_2688,N_2661);
xnor U4934 (N_4934,N_2716,N_3498);
nor U4935 (N_4935,N_3284,N_2579);
or U4936 (N_4936,N_3342,N_3747);
nor U4937 (N_4937,N_2907,N_2980);
nand U4938 (N_4938,N_3711,N_2795);
xor U4939 (N_4939,N_2161,N_2824);
and U4940 (N_4940,N_3538,N_2258);
and U4941 (N_4941,N_2720,N_3890);
or U4942 (N_4942,N_3867,N_2919);
nor U4943 (N_4943,N_3522,N_3763);
nand U4944 (N_4944,N_2598,N_2367);
and U4945 (N_4945,N_3213,N_2236);
nor U4946 (N_4946,N_3034,N_3221);
and U4947 (N_4947,N_2839,N_3764);
xor U4948 (N_4948,N_2423,N_2891);
xor U4949 (N_4949,N_2193,N_3128);
xnor U4950 (N_4950,N_3396,N_3161);
or U4951 (N_4951,N_2559,N_2981);
nand U4952 (N_4952,N_2696,N_2653);
xnor U4953 (N_4953,N_3393,N_2952);
and U4954 (N_4954,N_3965,N_2925);
xnor U4955 (N_4955,N_3770,N_3808);
nand U4956 (N_4956,N_2104,N_2576);
xnor U4957 (N_4957,N_2495,N_3537);
or U4958 (N_4958,N_2353,N_2563);
or U4959 (N_4959,N_2629,N_3236);
nor U4960 (N_4960,N_3627,N_2992);
xor U4961 (N_4961,N_2295,N_3998);
nand U4962 (N_4962,N_3118,N_3718);
nand U4963 (N_4963,N_3505,N_2812);
nor U4964 (N_4964,N_3188,N_2874);
nand U4965 (N_4965,N_3544,N_2105);
or U4966 (N_4966,N_3797,N_3684);
nand U4967 (N_4967,N_2638,N_2023);
nor U4968 (N_4968,N_2155,N_3117);
or U4969 (N_4969,N_3769,N_2115);
or U4970 (N_4970,N_3233,N_3064);
nand U4971 (N_4971,N_3799,N_3262);
nor U4972 (N_4972,N_2436,N_2953);
nand U4973 (N_4973,N_2335,N_3710);
nand U4974 (N_4974,N_3973,N_2575);
xor U4975 (N_4975,N_2908,N_2533);
xor U4976 (N_4976,N_3409,N_2971);
and U4977 (N_4977,N_2048,N_2806);
or U4978 (N_4978,N_2573,N_2042);
and U4979 (N_4979,N_3842,N_2832);
nand U4980 (N_4980,N_2555,N_3046);
or U4981 (N_4981,N_3103,N_3158);
and U4982 (N_4982,N_3553,N_2855);
or U4983 (N_4983,N_3780,N_3163);
nand U4984 (N_4984,N_3943,N_3822);
nor U4985 (N_4985,N_2172,N_3983);
xnor U4986 (N_4986,N_3976,N_3807);
or U4987 (N_4987,N_2496,N_2920);
xnor U4988 (N_4988,N_2817,N_2535);
xor U4989 (N_4989,N_3679,N_3313);
and U4990 (N_4990,N_3689,N_2117);
and U4991 (N_4991,N_3719,N_2960);
and U4992 (N_4992,N_2378,N_2966);
xnor U4993 (N_4993,N_2507,N_2304);
and U4994 (N_4994,N_3922,N_2242);
or U4995 (N_4995,N_3642,N_2756);
nor U4996 (N_4996,N_3308,N_2565);
nand U4997 (N_4997,N_2450,N_3886);
nor U4998 (N_4998,N_3686,N_2791);
and U4999 (N_4999,N_2227,N_3124);
nor U5000 (N_5000,N_2708,N_3841);
xnor U5001 (N_5001,N_3410,N_3096);
nor U5002 (N_5002,N_3719,N_2338);
xnor U5003 (N_5003,N_2838,N_2002);
xor U5004 (N_5004,N_3391,N_3466);
nor U5005 (N_5005,N_3687,N_3099);
nand U5006 (N_5006,N_2077,N_3573);
nor U5007 (N_5007,N_3941,N_2049);
nor U5008 (N_5008,N_3500,N_3748);
and U5009 (N_5009,N_3199,N_3135);
and U5010 (N_5010,N_2864,N_2859);
xnor U5011 (N_5011,N_2551,N_3092);
nor U5012 (N_5012,N_2973,N_3204);
nand U5013 (N_5013,N_2383,N_3344);
or U5014 (N_5014,N_3548,N_3338);
nand U5015 (N_5015,N_3550,N_2312);
xor U5016 (N_5016,N_2837,N_3326);
or U5017 (N_5017,N_2107,N_3556);
nor U5018 (N_5018,N_3120,N_3920);
nor U5019 (N_5019,N_2783,N_2095);
or U5020 (N_5020,N_3485,N_3150);
or U5021 (N_5021,N_2035,N_3946);
and U5022 (N_5022,N_3003,N_2434);
nand U5023 (N_5023,N_3962,N_2758);
nand U5024 (N_5024,N_3955,N_3263);
xnor U5025 (N_5025,N_3403,N_2846);
and U5026 (N_5026,N_2467,N_3138);
xor U5027 (N_5027,N_3110,N_2866);
xor U5028 (N_5028,N_3793,N_3104);
nand U5029 (N_5029,N_2903,N_2811);
nand U5030 (N_5030,N_2827,N_2630);
or U5031 (N_5031,N_2158,N_2846);
nor U5032 (N_5032,N_3558,N_3207);
and U5033 (N_5033,N_2074,N_2043);
and U5034 (N_5034,N_2033,N_3360);
nand U5035 (N_5035,N_2190,N_3674);
xnor U5036 (N_5036,N_2136,N_3934);
or U5037 (N_5037,N_2578,N_2965);
nor U5038 (N_5038,N_3395,N_2084);
xor U5039 (N_5039,N_3488,N_2498);
nor U5040 (N_5040,N_2874,N_2626);
nand U5041 (N_5041,N_2533,N_2551);
nand U5042 (N_5042,N_3103,N_2048);
and U5043 (N_5043,N_2717,N_2191);
xnor U5044 (N_5044,N_3015,N_2809);
xor U5045 (N_5045,N_2998,N_3739);
xor U5046 (N_5046,N_3023,N_2981);
and U5047 (N_5047,N_2653,N_2475);
nand U5048 (N_5048,N_3851,N_3531);
or U5049 (N_5049,N_3611,N_2860);
nand U5050 (N_5050,N_2558,N_3717);
and U5051 (N_5051,N_3605,N_2193);
and U5052 (N_5052,N_3975,N_3992);
nor U5053 (N_5053,N_3754,N_3738);
or U5054 (N_5054,N_2835,N_2755);
nor U5055 (N_5055,N_2339,N_3696);
or U5056 (N_5056,N_2875,N_2049);
or U5057 (N_5057,N_2029,N_2290);
and U5058 (N_5058,N_3825,N_2415);
or U5059 (N_5059,N_3872,N_2123);
or U5060 (N_5060,N_2351,N_3356);
or U5061 (N_5061,N_3654,N_2577);
and U5062 (N_5062,N_2432,N_3451);
xor U5063 (N_5063,N_2088,N_3348);
or U5064 (N_5064,N_2333,N_2860);
xnor U5065 (N_5065,N_3900,N_2617);
xnor U5066 (N_5066,N_3444,N_3066);
nand U5067 (N_5067,N_2658,N_2769);
nor U5068 (N_5068,N_3986,N_3435);
nand U5069 (N_5069,N_2062,N_3950);
nand U5070 (N_5070,N_3742,N_2012);
and U5071 (N_5071,N_2354,N_3480);
or U5072 (N_5072,N_2245,N_2267);
and U5073 (N_5073,N_2740,N_2892);
and U5074 (N_5074,N_2559,N_2007);
xor U5075 (N_5075,N_3966,N_3637);
and U5076 (N_5076,N_3360,N_3806);
or U5077 (N_5077,N_2631,N_3253);
xor U5078 (N_5078,N_3287,N_3667);
nand U5079 (N_5079,N_3523,N_3119);
or U5080 (N_5080,N_3653,N_3584);
or U5081 (N_5081,N_2398,N_2918);
nand U5082 (N_5082,N_2967,N_2161);
nor U5083 (N_5083,N_2270,N_3565);
or U5084 (N_5084,N_2166,N_3657);
nand U5085 (N_5085,N_2436,N_2901);
or U5086 (N_5086,N_3295,N_3807);
and U5087 (N_5087,N_2450,N_2197);
nor U5088 (N_5088,N_2920,N_3361);
nor U5089 (N_5089,N_3188,N_3271);
and U5090 (N_5090,N_2018,N_3084);
xnor U5091 (N_5091,N_3609,N_3039);
or U5092 (N_5092,N_2531,N_2798);
or U5093 (N_5093,N_2840,N_2942);
nor U5094 (N_5094,N_2264,N_3570);
nor U5095 (N_5095,N_2568,N_3729);
or U5096 (N_5096,N_3976,N_3435);
or U5097 (N_5097,N_3749,N_3492);
nand U5098 (N_5098,N_3820,N_2542);
and U5099 (N_5099,N_3732,N_2347);
and U5100 (N_5100,N_3949,N_3586);
or U5101 (N_5101,N_3731,N_2645);
xnor U5102 (N_5102,N_3003,N_2776);
nand U5103 (N_5103,N_3059,N_3204);
nand U5104 (N_5104,N_3991,N_2100);
nand U5105 (N_5105,N_2311,N_3578);
nor U5106 (N_5106,N_3591,N_2375);
and U5107 (N_5107,N_3802,N_2395);
nor U5108 (N_5108,N_2988,N_3350);
or U5109 (N_5109,N_2607,N_2859);
xnor U5110 (N_5110,N_3114,N_2438);
nor U5111 (N_5111,N_3048,N_2500);
or U5112 (N_5112,N_3937,N_2852);
or U5113 (N_5113,N_2991,N_3467);
nand U5114 (N_5114,N_3613,N_2618);
nand U5115 (N_5115,N_2486,N_2582);
nand U5116 (N_5116,N_2365,N_3305);
and U5117 (N_5117,N_2140,N_2105);
and U5118 (N_5118,N_2366,N_3987);
xnor U5119 (N_5119,N_3466,N_2897);
xnor U5120 (N_5120,N_2382,N_2504);
and U5121 (N_5121,N_2734,N_2320);
and U5122 (N_5122,N_2280,N_2898);
xor U5123 (N_5123,N_3600,N_2341);
or U5124 (N_5124,N_3049,N_3093);
nor U5125 (N_5125,N_3572,N_3345);
or U5126 (N_5126,N_3311,N_3973);
or U5127 (N_5127,N_3973,N_3792);
or U5128 (N_5128,N_2051,N_3870);
and U5129 (N_5129,N_2688,N_2351);
xor U5130 (N_5130,N_3468,N_2328);
xor U5131 (N_5131,N_3326,N_3590);
nand U5132 (N_5132,N_3577,N_2236);
xnor U5133 (N_5133,N_2965,N_3625);
nand U5134 (N_5134,N_2279,N_3525);
xnor U5135 (N_5135,N_2367,N_2122);
xor U5136 (N_5136,N_2121,N_2993);
nor U5137 (N_5137,N_2437,N_3758);
or U5138 (N_5138,N_3028,N_2364);
nand U5139 (N_5139,N_3351,N_3114);
and U5140 (N_5140,N_3517,N_2284);
nand U5141 (N_5141,N_2495,N_3889);
or U5142 (N_5142,N_3546,N_3048);
and U5143 (N_5143,N_3761,N_3254);
or U5144 (N_5144,N_2471,N_3230);
xor U5145 (N_5145,N_3381,N_3423);
xnor U5146 (N_5146,N_3790,N_3837);
and U5147 (N_5147,N_3046,N_2388);
and U5148 (N_5148,N_3308,N_2425);
nor U5149 (N_5149,N_2074,N_2814);
and U5150 (N_5150,N_2850,N_3833);
nor U5151 (N_5151,N_2015,N_3466);
and U5152 (N_5152,N_2410,N_2151);
or U5153 (N_5153,N_3483,N_3954);
or U5154 (N_5154,N_3328,N_3871);
and U5155 (N_5155,N_3535,N_3986);
nor U5156 (N_5156,N_3695,N_3432);
and U5157 (N_5157,N_3953,N_2129);
nor U5158 (N_5158,N_2947,N_2395);
xnor U5159 (N_5159,N_3892,N_2517);
nand U5160 (N_5160,N_3422,N_3262);
xnor U5161 (N_5161,N_3304,N_3072);
nor U5162 (N_5162,N_3268,N_2925);
nor U5163 (N_5163,N_2902,N_3843);
nor U5164 (N_5164,N_2214,N_3357);
nand U5165 (N_5165,N_2297,N_2498);
nor U5166 (N_5166,N_2423,N_2079);
and U5167 (N_5167,N_3088,N_2072);
and U5168 (N_5168,N_3784,N_3854);
nand U5169 (N_5169,N_2982,N_2265);
or U5170 (N_5170,N_3428,N_3983);
and U5171 (N_5171,N_3495,N_3822);
or U5172 (N_5172,N_3741,N_2526);
or U5173 (N_5173,N_2369,N_3280);
nor U5174 (N_5174,N_3082,N_3775);
or U5175 (N_5175,N_3120,N_3266);
or U5176 (N_5176,N_2660,N_2916);
nand U5177 (N_5177,N_2219,N_3509);
nor U5178 (N_5178,N_2907,N_3613);
nand U5179 (N_5179,N_2240,N_3624);
or U5180 (N_5180,N_2531,N_2691);
or U5181 (N_5181,N_2329,N_3320);
nand U5182 (N_5182,N_3473,N_2178);
or U5183 (N_5183,N_3813,N_3843);
xor U5184 (N_5184,N_3636,N_3880);
xnor U5185 (N_5185,N_3207,N_3781);
or U5186 (N_5186,N_3111,N_2656);
xor U5187 (N_5187,N_3134,N_3567);
xor U5188 (N_5188,N_3797,N_3952);
xnor U5189 (N_5189,N_3913,N_3483);
and U5190 (N_5190,N_2965,N_3982);
and U5191 (N_5191,N_3979,N_3492);
or U5192 (N_5192,N_2827,N_2845);
nor U5193 (N_5193,N_3173,N_3241);
and U5194 (N_5194,N_3182,N_2304);
nand U5195 (N_5195,N_3608,N_3717);
or U5196 (N_5196,N_3669,N_2259);
nand U5197 (N_5197,N_2090,N_2553);
and U5198 (N_5198,N_2257,N_2274);
nand U5199 (N_5199,N_3236,N_2411);
xor U5200 (N_5200,N_2983,N_2710);
xnor U5201 (N_5201,N_2850,N_2084);
xnor U5202 (N_5202,N_3317,N_3273);
nor U5203 (N_5203,N_3570,N_2905);
and U5204 (N_5204,N_2971,N_2886);
and U5205 (N_5205,N_2261,N_2105);
nand U5206 (N_5206,N_3677,N_2293);
or U5207 (N_5207,N_2718,N_2831);
xnor U5208 (N_5208,N_2384,N_2275);
or U5209 (N_5209,N_3619,N_3253);
nand U5210 (N_5210,N_2426,N_3715);
nand U5211 (N_5211,N_3932,N_3373);
nor U5212 (N_5212,N_2811,N_3073);
nor U5213 (N_5213,N_3965,N_3007);
and U5214 (N_5214,N_2529,N_2760);
nand U5215 (N_5215,N_3817,N_3230);
nand U5216 (N_5216,N_3095,N_3691);
nand U5217 (N_5217,N_2222,N_2193);
or U5218 (N_5218,N_2086,N_3015);
xor U5219 (N_5219,N_3323,N_2681);
nor U5220 (N_5220,N_3665,N_2637);
nand U5221 (N_5221,N_2115,N_3857);
nand U5222 (N_5222,N_2806,N_3520);
nand U5223 (N_5223,N_2441,N_2270);
xor U5224 (N_5224,N_3993,N_3829);
xor U5225 (N_5225,N_3291,N_2770);
nand U5226 (N_5226,N_3829,N_3796);
nor U5227 (N_5227,N_3818,N_2425);
nand U5228 (N_5228,N_2764,N_3748);
or U5229 (N_5229,N_3519,N_3296);
xnor U5230 (N_5230,N_2353,N_2819);
and U5231 (N_5231,N_2243,N_3986);
nand U5232 (N_5232,N_3825,N_3342);
xnor U5233 (N_5233,N_2201,N_3515);
nand U5234 (N_5234,N_3018,N_2716);
and U5235 (N_5235,N_3002,N_3508);
and U5236 (N_5236,N_2573,N_2190);
nand U5237 (N_5237,N_3790,N_3513);
nor U5238 (N_5238,N_3642,N_2392);
or U5239 (N_5239,N_3441,N_2116);
nand U5240 (N_5240,N_2786,N_3611);
nand U5241 (N_5241,N_3067,N_3403);
nand U5242 (N_5242,N_2325,N_2348);
xor U5243 (N_5243,N_2892,N_3371);
or U5244 (N_5244,N_3134,N_3790);
nor U5245 (N_5245,N_3479,N_3343);
and U5246 (N_5246,N_3482,N_2756);
nor U5247 (N_5247,N_2721,N_3477);
nor U5248 (N_5248,N_2368,N_3949);
or U5249 (N_5249,N_3971,N_2304);
and U5250 (N_5250,N_3016,N_2817);
xor U5251 (N_5251,N_2405,N_3054);
xor U5252 (N_5252,N_2729,N_3343);
or U5253 (N_5253,N_2156,N_2361);
or U5254 (N_5254,N_2038,N_3668);
xor U5255 (N_5255,N_3133,N_2600);
and U5256 (N_5256,N_3476,N_3407);
nor U5257 (N_5257,N_3833,N_3579);
and U5258 (N_5258,N_3867,N_3369);
or U5259 (N_5259,N_2158,N_3426);
nor U5260 (N_5260,N_3429,N_2009);
nor U5261 (N_5261,N_2232,N_2064);
xor U5262 (N_5262,N_2611,N_2237);
xor U5263 (N_5263,N_3491,N_3504);
nand U5264 (N_5264,N_2921,N_2146);
xnor U5265 (N_5265,N_2608,N_3579);
nor U5266 (N_5266,N_3563,N_3958);
nor U5267 (N_5267,N_3062,N_2487);
or U5268 (N_5268,N_2608,N_2785);
nor U5269 (N_5269,N_3472,N_3418);
and U5270 (N_5270,N_3584,N_2500);
or U5271 (N_5271,N_2368,N_3846);
and U5272 (N_5272,N_3173,N_2619);
nor U5273 (N_5273,N_2871,N_3367);
xnor U5274 (N_5274,N_3854,N_2810);
nand U5275 (N_5275,N_2681,N_2677);
and U5276 (N_5276,N_2557,N_3680);
xor U5277 (N_5277,N_3068,N_3460);
nand U5278 (N_5278,N_3197,N_3343);
or U5279 (N_5279,N_3456,N_2828);
xor U5280 (N_5280,N_3100,N_2983);
nor U5281 (N_5281,N_2194,N_3619);
nand U5282 (N_5282,N_2384,N_2342);
xnor U5283 (N_5283,N_3546,N_3274);
nand U5284 (N_5284,N_3776,N_3339);
nand U5285 (N_5285,N_3761,N_2910);
and U5286 (N_5286,N_3429,N_2758);
nand U5287 (N_5287,N_3272,N_3693);
xnor U5288 (N_5288,N_3521,N_3028);
xor U5289 (N_5289,N_3663,N_2071);
xor U5290 (N_5290,N_3318,N_2004);
xor U5291 (N_5291,N_2884,N_2737);
or U5292 (N_5292,N_2790,N_3156);
nor U5293 (N_5293,N_3611,N_2712);
nor U5294 (N_5294,N_3473,N_3913);
or U5295 (N_5295,N_3896,N_3599);
nand U5296 (N_5296,N_2357,N_3556);
xnor U5297 (N_5297,N_2074,N_2405);
and U5298 (N_5298,N_2489,N_2975);
xor U5299 (N_5299,N_3064,N_2636);
nand U5300 (N_5300,N_3613,N_3918);
nand U5301 (N_5301,N_2604,N_3971);
and U5302 (N_5302,N_3869,N_2033);
nand U5303 (N_5303,N_3129,N_2535);
xnor U5304 (N_5304,N_3087,N_2062);
or U5305 (N_5305,N_2499,N_2160);
or U5306 (N_5306,N_2473,N_3350);
nand U5307 (N_5307,N_3290,N_2226);
and U5308 (N_5308,N_2640,N_2205);
or U5309 (N_5309,N_3791,N_3667);
or U5310 (N_5310,N_2192,N_3696);
nor U5311 (N_5311,N_2168,N_2091);
xnor U5312 (N_5312,N_3340,N_2981);
xor U5313 (N_5313,N_3748,N_3626);
nor U5314 (N_5314,N_2850,N_3534);
nand U5315 (N_5315,N_2261,N_2520);
or U5316 (N_5316,N_3559,N_3192);
xnor U5317 (N_5317,N_3759,N_3316);
nor U5318 (N_5318,N_2200,N_2501);
or U5319 (N_5319,N_2452,N_3922);
and U5320 (N_5320,N_3506,N_3973);
nand U5321 (N_5321,N_2993,N_3831);
or U5322 (N_5322,N_2542,N_3547);
nand U5323 (N_5323,N_2942,N_2400);
nand U5324 (N_5324,N_3093,N_2541);
nor U5325 (N_5325,N_2474,N_2373);
nor U5326 (N_5326,N_3659,N_2992);
and U5327 (N_5327,N_3812,N_2964);
nor U5328 (N_5328,N_2125,N_3318);
xor U5329 (N_5329,N_2467,N_3320);
or U5330 (N_5330,N_3039,N_3115);
or U5331 (N_5331,N_2307,N_3952);
and U5332 (N_5332,N_2831,N_3966);
xor U5333 (N_5333,N_2665,N_2829);
xnor U5334 (N_5334,N_2091,N_2075);
nor U5335 (N_5335,N_2158,N_3359);
nor U5336 (N_5336,N_2434,N_2819);
xnor U5337 (N_5337,N_2367,N_3661);
or U5338 (N_5338,N_3183,N_3919);
xnor U5339 (N_5339,N_3866,N_3325);
nor U5340 (N_5340,N_2504,N_2572);
xnor U5341 (N_5341,N_2130,N_3761);
and U5342 (N_5342,N_2511,N_2272);
and U5343 (N_5343,N_3054,N_3314);
xnor U5344 (N_5344,N_3712,N_2078);
nand U5345 (N_5345,N_3378,N_2601);
or U5346 (N_5346,N_2462,N_3199);
nand U5347 (N_5347,N_2650,N_2382);
and U5348 (N_5348,N_2061,N_2311);
or U5349 (N_5349,N_3473,N_3675);
xor U5350 (N_5350,N_3570,N_3338);
xor U5351 (N_5351,N_2861,N_2183);
nand U5352 (N_5352,N_3325,N_3358);
xnor U5353 (N_5353,N_3030,N_3979);
or U5354 (N_5354,N_3436,N_3602);
or U5355 (N_5355,N_3756,N_2606);
and U5356 (N_5356,N_3293,N_2051);
xor U5357 (N_5357,N_2186,N_3714);
or U5358 (N_5358,N_2590,N_2878);
nor U5359 (N_5359,N_3999,N_3571);
nand U5360 (N_5360,N_2999,N_2779);
xor U5361 (N_5361,N_2785,N_2571);
nor U5362 (N_5362,N_3431,N_3849);
and U5363 (N_5363,N_3426,N_3321);
and U5364 (N_5364,N_2566,N_3545);
xor U5365 (N_5365,N_3492,N_2313);
or U5366 (N_5366,N_2883,N_3594);
nand U5367 (N_5367,N_3687,N_2645);
nand U5368 (N_5368,N_2897,N_3930);
and U5369 (N_5369,N_3850,N_2621);
nand U5370 (N_5370,N_2092,N_3182);
nor U5371 (N_5371,N_3097,N_2304);
or U5372 (N_5372,N_3325,N_2213);
or U5373 (N_5373,N_2458,N_2244);
nor U5374 (N_5374,N_2089,N_2082);
nor U5375 (N_5375,N_3237,N_3612);
or U5376 (N_5376,N_2871,N_2466);
xnor U5377 (N_5377,N_2426,N_3550);
and U5378 (N_5378,N_2408,N_2948);
and U5379 (N_5379,N_2659,N_2223);
xor U5380 (N_5380,N_2601,N_3567);
or U5381 (N_5381,N_2185,N_3180);
xor U5382 (N_5382,N_2038,N_2515);
or U5383 (N_5383,N_3429,N_3572);
xnor U5384 (N_5384,N_2177,N_3202);
nor U5385 (N_5385,N_3209,N_2669);
nor U5386 (N_5386,N_3992,N_3072);
nor U5387 (N_5387,N_2463,N_3883);
or U5388 (N_5388,N_3343,N_2671);
xor U5389 (N_5389,N_3979,N_2449);
or U5390 (N_5390,N_3994,N_3387);
nor U5391 (N_5391,N_2003,N_3588);
or U5392 (N_5392,N_2846,N_2627);
nand U5393 (N_5393,N_3969,N_3995);
nor U5394 (N_5394,N_2405,N_2684);
xor U5395 (N_5395,N_2521,N_2813);
nor U5396 (N_5396,N_3648,N_2364);
or U5397 (N_5397,N_3009,N_3441);
xor U5398 (N_5398,N_3304,N_3242);
or U5399 (N_5399,N_2938,N_2719);
nor U5400 (N_5400,N_3665,N_2483);
or U5401 (N_5401,N_3301,N_3026);
and U5402 (N_5402,N_2429,N_3617);
nor U5403 (N_5403,N_2775,N_3267);
xor U5404 (N_5404,N_2730,N_3585);
and U5405 (N_5405,N_2727,N_2333);
nand U5406 (N_5406,N_2935,N_2011);
nor U5407 (N_5407,N_2263,N_3923);
or U5408 (N_5408,N_3457,N_2589);
and U5409 (N_5409,N_3930,N_2511);
nor U5410 (N_5410,N_2745,N_2304);
nand U5411 (N_5411,N_3946,N_3991);
or U5412 (N_5412,N_2911,N_3877);
or U5413 (N_5413,N_2261,N_2396);
nor U5414 (N_5414,N_2458,N_3032);
nor U5415 (N_5415,N_3666,N_3638);
xor U5416 (N_5416,N_2266,N_2587);
nand U5417 (N_5417,N_2364,N_3946);
and U5418 (N_5418,N_2072,N_3148);
nand U5419 (N_5419,N_2732,N_2573);
nor U5420 (N_5420,N_2275,N_3842);
nand U5421 (N_5421,N_3391,N_2898);
and U5422 (N_5422,N_2777,N_2903);
nand U5423 (N_5423,N_2424,N_3112);
and U5424 (N_5424,N_2818,N_3247);
xor U5425 (N_5425,N_2599,N_2320);
or U5426 (N_5426,N_3381,N_2768);
nor U5427 (N_5427,N_3354,N_2255);
or U5428 (N_5428,N_2007,N_2391);
or U5429 (N_5429,N_3980,N_3758);
and U5430 (N_5430,N_3568,N_3246);
nand U5431 (N_5431,N_2841,N_3835);
and U5432 (N_5432,N_2867,N_2585);
nand U5433 (N_5433,N_3316,N_3477);
and U5434 (N_5434,N_2951,N_2542);
and U5435 (N_5435,N_3010,N_2991);
xnor U5436 (N_5436,N_2805,N_3449);
or U5437 (N_5437,N_3553,N_2561);
nor U5438 (N_5438,N_3135,N_2452);
and U5439 (N_5439,N_3422,N_2374);
nand U5440 (N_5440,N_3464,N_2841);
and U5441 (N_5441,N_2557,N_2577);
and U5442 (N_5442,N_2909,N_2720);
xor U5443 (N_5443,N_3710,N_3086);
nand U5444 (N_5444,N_2874,N_2344);
nor U5445 (N_5445,N_3398,N_2916);
nand U5446 (N_5446,N_3879,N_2139);
nor U5447 (N_5447,N_3407,N_2096);
and U5448 (N_5448,N_3256,N_3122);
nand U5449 (N_5449,N_3687,N_2346);
xor U5450 (N_5450,N_3913,N_3146);
xor U5451 (N_5451,N_3946,N_2426);
xor U5452 (N_5452,N_3859,N_2217);
nor U5453 (N_5453,N_3816,N_3024);
and U5454 (N_5454,N_3613,N_3465);
or U5455 (N_5455,N_3023,N_3270);
xnor U5456 (N_5456,N_3394,N_3515);
nor U5457 (N_5457,N_3034,N_2866);
or U5458 (N_5458,N_3425,N_2336);
nor U5459 (N_5459,N_2356,N_2479);
nor U5460 (N_5460,N_3599,N_2924);
and U5461 (N_5461,N_2512,N_3972);
or U5462 (N_5462,N_3668,N_2138);
or U5463 (N_5463,N_3246,N_3939);
nor U5464 (N_5464,N_2417,N_2994);
or U5465 (N_5465,N_2204,N_3327);
and U5466 (N_5466,N_3958,N_2363);
and U5467 (N_5467,N_2253,N_2302);
nor U5468 (N_5468,N_2817,N_2648);
nor U5469 (N_5469,N_2115,N_2245);
nor U5470 (N_5470,N_2925,N_3395);
nand U5471 (N_5471,N_3679,N_3763);
and U5472 (N_5472,N_3916,N_2959);
nand U5473 (N_5473,N_2834,N_2049);
and U5474 (N_5474,N_3339,N_2918);
nand U5475 (N_5475,N_3741,N_2045);
or U5476 (N_5476,N_2890,N_2318);
nor U5477 (N_5477,N_3105,N_2318);
and U5478 (N_5478,N_3174,N_2912);
and U5479 (N_5479,N_3791,N_3145);
nand U5480 (N_5480,N_2766,N_2740);
xnor U5481 (N_5481,N_3459,N_2318);
or U5482 (N_5482,N_2745,N_3970);
xor U5483 (N_5483,N_2390,N_3296);
nand U5484 (N_5484,N_3575,N_3369);
and U5485 (N_5485,N_3075,N_3641);
and U5486 (N_5486,N_2446,N_3738);
and U5487 (N_5487,N_2053,N_3936);
nor U5488 (N_5488,N_3080,N_2416);
or U5489 (N_5489,N_3323,N_2208);
or U5490 (N_5490,N_2064,N_3529);
nor U5491 (N_5491,N_2304,N_2996);
nor U5492 (N_5492,N_3150,N_2394);
or U5493 (N_5493,N_2162,N_3632);
nand U5494 (N_5494,N_3527,N_2242);
and U5495 (N_5495,N_3086,N_2840);
nand U5496 (N_5496,N_2674,N_3259);
nand U5497 (N_5497,N_3400,N_3830);
xor U5498 (N_5498,N_3225,N_2370);
xor U5499 (N_5499,N_2039,N_2343);
nor U5500 (N_5500,N_3494,N_2695);
and U5501 (N_5501,N_3572,N_3640);
or U5502 (N_5502,N_2533,N_3759);
and U5503 (N_5503,N_3579,N_3999);
nand U5504 (N_5504,N_3708,N_2587);
nand U5505 (N_5505,N_2530,N_2235);
xor U5506 (N_5506,N_2077,N_2169);
or U5507 (N_5507,N_2930,N_2351);
xnor U5508 (N_5508,N_2362,N_3047);
nor U5509 (N_5509,N_3191,N_2795);
or U5510 (N_5510,N_3548,N_2194);
or U5511 (N_5511,N_2922,N_3975);
nand U5512 (N_5512,N_2704,N_2991);
or U5513 (N_5513,N_2553,N_2083);
or U5514 (N_5514,N_2815,N_3805);
or U5515 (N_5515,N_2516,N_2003);
and U5516 (N_5516,N_2230,N_2244);
nand U5517 (N_5517,N_2320,N_3152);
nand U5518 (N_5518,N_3313,N_3778);
nand U5519 (N_5519,N_2337,N_3249);
nor U5520 (N_5520,N_2104,N_3374);
and U5521 (N_5521,N_2055,N_2951);
nand U5522 (N_5522,N_2009,N_3948);
xnor U5523 (N_5523,N_3126,N_2653);
xor U5524 (N_5524,N_3104,N_2226);
nand U5525 (N_5525,N_3858,N_3445);
and U5526 (N_5526,N_3037,N_2126);
and U5527 (N_5527,N_2283,N_3502);
nor U5528 (N_5528,N_2645,N_3101);
and U5529 (N_5529,N_3612,N_3221);
nor U5530 (N_5530,N_3567,N_3035);
nand U5531 (N_5531,N_2682,N_2943);
xor U5532 (N_5532,N_2238,N_3611);
nor U5533 (N_5533,N_2916,N_2941);
xnor U5534 (N_5534,N_3684,N_3396);
or U5535 (N_5535,N_3436,N_3173);
xnor U5536 (N_5536,N_2486,N_3330);
and U5537 (N_5537,N_2405,N_3565);
nand U5538 (N_5538,N_3760,N_3227);
nor U5539 (N_5539,N_3500,N_3239);
nand U5540 (N_5540,N_2003,N_3194);
or U5541 (N_5541,N_2213,N_2487);
nand U5542 (N_5542,N_2269,N_3234);
nand U5543 (N_5543,N_2959,N_2408);
xnor U5544 (N_5544,N_2786,N_2668);
xor U5545 (N_5545,N_3987,N_3820);
and U5546 (N_5546,N_2555,N_2643);
and U5547 (N_5547,N_3968,N_3903);
and U5548 (N_5548,N_3177,N_2856);
or U5549 (N_5549,N_2478,N_2968);
nand U5550 (N_5550,N_2385,N_2492);
nand U5551 (N_5551,N_3961,N_3186);
or U5552 (N_5552,N_2565,N_2421);
or U5553 (N_5553,N_3291,N_2836);
nor U5554 (N_5554,N_3777,N_2585);
or U5555 (N_5555,N_3546,N_3267);
nor U5556 (N_5556,N_3636,N_3582);
or U5557 (N_5557,N_3760,N_3091);
nor U5558 (N_5558,N_2073,N_2997);
nand U5559 (N_5559,N_2833,N_3289);
xor U5560 (N_5560,N_2414,N_2689);
or U5561 (N_5561,N_3391,N_3807);
xor U5562 (N_5562,N_3789,N_2046);
or U5563 (N_5563,N_3823,N_2014);
or U5564 (N_5564,N_2473,N_2246);
xor U5565 (N_5565,N_2308,N_3920);
and U5566 (N_5566,N_2704,N_2253);
nand U5567 (N_5567,N_3438,N_3948);
and U5568 (N_5568,N_2811,N_3836);
nand U5569 (N_5569,N_2638,N_2779);
and U5570 (N_5570,N_2696,N_3004);
nand U5571 (N_5571,N_2972,N_2565);
xnor U5572 (N_5572,N_3294,N_3041);
xor U5573 (N_5573,N_3293,N_3342);
xor U5574 (N_5574,N_3694,N_2474);
xnor U5575 (N_5575,N_2720,N_3863);
xnor U5576 (N_5576,N_3450,N_3673);
or U5577 (N_5577,N_3884,N_3427);
or U5578 (N_5578,N_2307,N_2764);
and U5579 (N_5579,N_2407,N_2661);
and U5580 (N_5580,N_2509,N_3713);
nor U5581 (N_5581,N_3967,N_3727);
or U5582 (N_5582,N_2692,N_3616);
or U5583 (N_5583,N_2589,N_2080);
nor U5584 (N_5584,N_2103,N_2667);
and U5585 (N_5585,N_2672,N_3421);
xor U5586 (N_5586,N_3013,N_3088);
or U5587 (N_5587,N_2937,N_2790);
or U5588 (N_5588,N_2922,N_2391);
nor U5589 (N_5589,N_3721,N_3106);
nor U5590 (N_5590,N_3848,N_3924);
nand U5591 (N_5591,N_2167,N_2576);
or U5592 (N_5592,N_3076,N_2942);
xnor U5593 (N_5593,N_2673,N_2100);
or U5594 (N_5594,N_3917,N_3461);
nor U5595 (N_5595,N_2408,N_2793);
xor U5596 (N_5596,N_2234,N_3736);
nand U5597 (N_5597,N_2571,N_2083);
nand U5598 (N_5598,N_2214,N_2615);
and U5599 (N_5599,N_2400,N_2338);
xnor U5600 (N_5600,N_2470,N_2199);
nand U5601 (N_5601,N_2902,N_2573);
xor U5602 (N_5602,N_3178,N_2719);
or U5603 (N_5603,N_3871,N_3382);
nand U5604 (N_5604,N_3059,N_2771);
and U5605 (N_5605,N_2541,N_3397);
nor U5606 (N_5606,N_3377,N_2430);
or U5607 (N_5607,N_2724,N_2534);
or U5608 (N_5608,N_2183,N_3748);
nor U5609 (N_5609,N_3739,N_3780);
nor U5610 (N_5610,N_3424,N_2603);
nor U5611 (N_5611,N_2046,N_2888);
xor U5612 (N_5612,N_2139,N_3746);
nand U5613 (N_5613,N_2268,N_2003);
xnor U5614 (N_5614,N_2557,N_3158);
and U5615 (N_5615,N_3773,N_2180);
or U5616 (N_5616,N_2347,N_2228);
nand U5617 (N_5617,N_3573,N_3623);
or U5618 (N_5618,N_2952,N_2461);
nand U5619 (N_5619,N_3318,N_2884);
nand U5620 (N_5620,N_3470,N_3210);
or U5621 (N_5621,N_2688,N_2753);
nor U5622 (N_5622,N_2931,N_3597);
or U5623 (N_5623,N_3723,N_3325);
or U5624 (N_5624,N_2244,N_2619);
xnor U5625 (N_5625,N_2179,N_3986);
xnor U5626 (N_5626,N_3753,N_2122);
nor U5627 (N_5627,N_3289,N_2416);
and U5628 (N_5628,N_3142,N_2009);
or U5629 (N_5629,N_2874,N_3117);
or U5630 (N_5630,N_2710,N_2279);
xnor U5631 (N_5631,N_2878,N_3309);
and U5632 (N_5632,N_2233,N_3166);
xnor U5633 (N_5633,N_3551,N_2726);
and U5634 (N_5634,N_2769,N_2166);
and U5635 (N_5635,N_2748,N_3793);
or U5636 (N_5636,N_3699,N_2573);
nor U5637 (N_5637,N_3338,N_3265);
and U5638 (N_5638,N_3247,N_3695);
xnor U5639 (N_5639,N_2075,N_2884);
and U5640 (N_5640,N_3527,N_3646);
nand U5641 (N_5641,N_3142,N_2001);
or U5642 (N_5642,N_2370,N_3104);
xor U5643 (N_5643,N_2421,N_3529);
xnor U5644 (N_5644,N_2901,N_2450);
or U5645 (N_5645,N_3546,N_3068);
or U5646 (N_5646,N_2035,N_3273);
xnor U5647 (N_5647,N_2525,N_3232);
and U5648 (N_5648,N_3318,N_3025);
nand U5649 (N_5649,N_3078,N_2991);
nor U5650 (N_5650,N_3996,N_3287);
or U5651 (N_5651,N_3931,N_2918);
xnor U5652 (N_5652,N_2039,N_2063);
or U5653 (N_5653,N_3752,N_2957);
and U5654 (N_5654,N_3858,N_2988);
and U5655 (N_5655,N_2666,N_2766);
xor U5656 (N_5656,N_2069,N_3100);
nand U5657 (N_5657,N_2680,N_2875);
and U5658 (N_5658,N_3960,N_2924);
and U5659 (N_5659,N_2943,N_3046);
or U5660 (N_5660,N_3206,N_2049);
nand U5661 (N_5661,N_3021,N_2656);
and U5662 (N_5662,N_2229,N_3217);
or U5663 (N_5663,N_3922,N_2266);
and U5664 (N_5664,N_2974,N_2490);
nor U5665 (N_5665,N_3247,N_3899);
and U5666 (N_5666,N_2605,N_2925);
nor U5667 (N_5667,N_2338,N_3291);
xnor U5668 (N_5668,N_2435,N_3264);
and U5669 (N_5669,N_2292,N_3146);
nand U5670 (N_5670,N_3795,N_3592);
nor U5671 (N_5671,N_3294,N_3624);
xnor U5672 (N_5672,N_3490,N_2383);
or U5673 (N_5673,N_2043,N_2121);
nor U5674 (N_5674,N_2634,N_2649);
xor U5675 (N_5675,N_3291,N_2640);
or U5676 (N_5676,N_2273,N_2844);
nor U5677 (N_5677,N_2128,N_3994);
nand U5678 (N_5678,N_2880,N_3856);
nand U5679 (N_5679,N_2173,N_2946);
nand U5680 (N_5680,N_3560,N_3242);
nor U5681 (N_5681,N_2768,N_3181);
and U5682 (N_5682,N_2659,N_2081);
or U5683 (N_5683,N_2308,N_3677);
nor U5684 (N_5684,N_2593,N_3407);
and U5685 (N_5685,N_3866,N_2950);
nand U5686 (N_5686,N_3489,N_3622);
nor U5687 (N_5687,N_2709,N_2424);
nand U5688 (N_5688,N_3343,N_2538);
or U5689 (N_5689,N_2052,N_3045);
nor U5690 (N_5690,N_3157,N_3222);
nor U5691 (N_5691,N_3542,N_2106);
nor U5692 (N_5692,N_3904,N_3620);
or U5693 (N_5693,N_2569,N_3894);
nor U5694 (N_5694,N_2775,N_3635);
nor U5695 (N_5695,N_2024,N_3716);
nand U5696 (N_5696,N_3025,N_3261);
xor U5697 (N_5697,N_3781,N_2159);
or U5698 (N_5698,N_3266,N_3698);
nor U5699 (N_5699,N_3799,N_2772);
and U5700 (N_5700,N_2485,N_3965);
and U5701 (N_5701,N_3533,N_2206);
and U5702 (N_5702,N_3871,N_2658);
and U5703 (N_5703,N_2159,N_3974);
xnor U5704 (N_5704,N_3907,N_3680);
nor U5705 (N_5705,N_3818,N_2954);
xnor U5706 (N_5706,N_2190,N_2897);
xnor U5707 (N_5707,N_3367,N_2416);
xor U5708 (N_5708,N_3830,N_3368);
nand U5709 (N_5709,N_2390,N_3231);
or U5710 (N_5710,N_3325,N_3065);
and U5711 (N_5711,N_3322,N_3039);
nand U5712 (N_5712,N_2277,N_3642);
and U5713 (N_5713,N_2098,N_2329);
xor U5714 (N_5714,N_3493,N_3193);
nor U5715 (N_5715,N_2132,N_2778);
xor U5716 (N_5716,N_3616,N_2428);
nand U5717 (N_5717,N_3860,N_3290);
nor U5718 (N_5718,N_2909,N_3487);
nor U5719 (N_5719,N_2167,N_2870);
xor U5720 (N_5720,N_2763,N_2776);
nand U5721 (N_5721,N_2797,N_3280);
nand U5722 (N_5722,N_3171,N_3896);
nor U5723 (N_5723,N_3585,N_3143);
nand U5724 (N_5724,N_3232,N_3020);
xnor U5725 (N_5725,N_2816,N_3184);
xnor U5726 (N_5726,N_3618,N_2833);
and U5727 (N_5727,N_3408,N_3711);
nor U5728 (N_5728,N_2199,N_2710);
and U5729 (N_5729,N_3932,N_2564);
xor U5730 (N_5730,N_3290,N_2462);
nor U5731 (N_5731,N_3880,N_2336);
nand U5732 (N_5732,N_3069,N_2091);
nand U5733 (N_5733,N_2806,N_2340);
and U5734 (N_5734,N_3769,N_2654);
nand U5735 (N_5735,N_2255,N_3767);
xnor U5736 (N_5736,N_3526,N_3960);
nor U5737 (N_5737,N_2720,N_2194);
xor U5738 (N_5738,N_2489,N_3828);
or U5739 (N_5739,N_2509,N_3347);
or U5740 (N_5740,N_2830,N_3025);
nor U5741 (N_5741,N_3890,N_3339);
nand U5742 (N_5742,N_3072,N_3713);
or U5743 (N_5743,N_3660,N_3817);
nor U5744 (N_5744,N_3243,N_2081);
or U5745 (N_5745,N_2153,N_2395);
xor U5746 (N_5746,N_2011,N_2370);
and U5747 (N_5747,N_3017,N_3237);
nor U5748 (N_5748,N_2857,N_2117);
and U5749 (N_5749,N_3604,N_2599);
xor U5750 (N_5750,N_2212,N_3042);
nor U5751 (N_5751,N_3223,N_3970);
or U5752 (N_5752,N_2394,N_2727);
nor U5753 (N_5753,N_3577,N_3467);
and U5754 (N_5754,N_2278,N_2266);
and U5755 (N_5755,N_3237,N_2173);
nor U5756 (N_5756,N_3690,N_3232);
and U5757 (N_5757,N_2858,N_2176);
nand U5758 (N_5758,N_3363,N_3135);
xnor U5759 (N_5759,N_3327,N_2991);
nor U5760 (N_5760,N_3830,N_2828);
nand U5761 (N_5761,N_2011,N_3785);
and U5762 (N_5762,N_3002,N_3444);
and U5763 (N_5763,N_3346,N_3473);
xor U5764 (N_5764,N_3385,N_3766);
xnor U5765 (N_5765,N_2251,N_2854);
or U5766 (N_5766,N_2013,N_3722);
xor U5767 (N_5767,N_2909,N_2144);
nor U5768 (N_5768,N_2485,N_2767);
xor U5769 (N_5769,N_3050,N_2968);
and U5770 (N_5770,N_2311,N_2312);
nor U5771 (N_5771,N_3810,N_2078);
or U5772 (N_5772,N_2970,N_2629);
nand U5773 (N_5773,N_2943,N_2218);
nor U5774 (N_5774,N_2438,N_2317);
xor U5775 (N_5775,N_2852,N_2725);
and U5776 (N_5776,N_3633,N_3217);
or U5777 (N_5777,N_3434,N_2515);
nand U5778 (N_5778,N_2679,N_2895);
nor U5779 (N_5779,N_2763,N_2260);
or U5780 (N_5780,N_2833,N_2846);
nor U5781 (N_5781,N_3207,N_3575);
and U5782 (N_5782,N_2228,N_2767);
nand U5783 (N_5783,N_2385,N_2194);
nand U5784 (N_5784,N_3665,N_2428);
and U5785 (N_5785,N_3361,N_3776);
nand U5786 (N_5786,N_3572,N_2273);
and U5787 (N_5787,N_2364,N_3351);
or U5788 (N_5788,N_3232,N_3209);
nor U5789 (N_5789,N_3812,N_2421);
nor U5790 (N_5790,N_3125,N_3523);
and U5791 (N_5791,N_2083,N_2737);
and U5792 (N_5792,N_2675,N_3568);
xnor U5793 (N_5793,N_2933,N_2013);
nor U5794 (N_5794,N_2412,N_2590);
and U5795 (N_5795,N_3997,N_2437);
or U5796 (N_5796,N_2031,N_3283);
and U5797 (N_5797,N_3251,N_3381);
nor U5798 (N_5798,N_3245,N_3938);
and U5799 (N_5799,N_3305,N_2296);
and U5800 (N_5800,N_3730,N_3032);
or U5801 (N_5801,N_2455,N_3937);
xnor U5802 (N_5802,N_3748,N_3451);
nand U5803 (N_5803,N_3972,N_2967);
and U5804 (N_5804,N_3028,N_2438);
or U5805 (N_5805,N_2497,N_3975);
nor U5806 (N_5806,N_2574,N_2212);
and U5807 (N_5807,N_2980,N_3962);
or U5808 (N_5808,N_3495,N_2123);
and U5809 (N_5809,N_2365,N_2482);
and U5810 (N_5810,N_3840,N_2947);
nor U5811 (N_5811,N_2522,N_3294);
nor U5812 (N_5812,N_2305,N_3836);
xnor U5813 (N_5813,N_3374,N_3770);
nand U5814 (N_5814,N_2211,N_3474);
nor U5815 (N_5815,N_3426,N_3449);
nand U5816 (N_5816,N_3208,N_3573);
xnor U5817 (N_5817,N_3500,N_2549);
or U5818 (N_5818,N_2995,N_3617);
nor U5819 (N_5819,N_2350,N_2826);
and U5820 (N_5820,N_2734,N_2825);
or U5821 (N_5821,N_2409,N_3707);
nor U5822 (N_5822,N_3614,N_2906);
nand U5823 (N_5823,N_2337,N_3293);
xor U5824 (N_5824,N_2706,N_3287);
xnor U5825 (N_5825,N_2661,N_3196);
or U5826 (N_5826,N_2289,N_2773);
nand U5827 (N_5827,N_2142,N_2475);
and U5828 (N_5828,N_3596,N_2320);
and U5829 (N_5829,N_3932,N_3715);
and U5830 (N_5830,N_2365,N_3833);
nand U5831 (N_5831,N_2243,N_2136);
xor U5832 (N_5832,N_2158,N_3461);
nor U5833 (N_5833,N_3321,N_3820);
xnor U5834 (N_5834,N_2226,N_3767);
or U5835 (N_5835,N_3971,N_3407);
and U5836 (N_5836,N_2464,N_3116);
and U5837 (N_5837,N_3653,N_2479);
xnor U5838 (N_5838,N_3879,N_2926);
xnor U5839 (N_5839,N_3155,N_2871);
nand U5840 (N_5840,N_3123,N_2587);
or U5841 (N_5841,N_2288,N_2456);
or U5842 (N_5842,N_3629,N_3961);
nand U5843 (N_5843,N_3960,N_2735);
xnor U5844 (N_5844,N_3613,N_2142);
nor U5845 (N_5845,N_3338,N_2248);
or U5846 (N_5846,N_2770,N_3776);
nor U5847 (N_5847,N_3250,N_2152);
xor U5848 (N_5848,N_3968,N_2780);
or U5849 (N_5849,N_2908,N_3160);
or U5850 (N_5850,N_2531,N_2367);
xor U5851 (N_5851,N_3926,N_2908);
and U5852 (N_5852,N_2654,N_2354);
nand U5853 (N_5853,N_2670,N_2294);
xor U5854 (N_5854,N_3568,N_3554);
or U5855 (N_5855,N_2034,N_2987);
or U5856 (N_5856,N_2652,N_2209);
nor U5857 (N_5857,N_2481,N_3908);
or U5858 (N_5858,N_3482,N_2014);
nor U5859 (N_5859,N_2542,N_3128);
nor U5860 (N_5860,N_3036,N_2136);
xnor U5861 (N_5861,N_2800,N_3780);
nor U5862 (N_5862,N_3528,N_3972);
nand U5863 (N_5863,N_2419,N_2708);
nor U5864 (N_5864,N_3371,N_3612);
and U5865 (N_5865,N_3446,N_2651);
nor U5866 (N_5866,N_2235,N_2971);
nand U5867 (N_5867,N_3043,N_3628);
xnor U5868 (N_5868,N_3785,N_3929);
or U5869 (N_5869,N_3317,N_3373);
xnor U5870 (N_5870,N_3830,N_3349);
and U5871 (N_5871,N_3590,N_3167);
xor U5872 (N_5872,N_2945,N_3952);
or U5873 (N_5873,N_2591,N_3870);
or U5874 (N_5874,N_3069,N_3118);
nor U5875 (N_5875,N_3773,N_3109);
and U5876 (N_5876,N_3495,N_2466);
xor U5877 (N_5877,N_3669,N_2581);
or U5878 (N_5878,N_2508,N_3070);
and U5879 (N_5879,N_2178,N_3763);
and U5880 (N_5880,N_3191,N_3028);
xor U5881 (N_5881,N_2461,N_3408);
or U5882 (N_5882,N_2665,N_2709);
or U5883 (N_5883,N_3979,N_3786);
xor U5884 (N_5884,N_3618,N_3655);
or U5885 (N_5885,N_3114,N_2572);
xor U5886 (N_5886,N_3107,N_2835);
or U5887 (N_5887,N_2121,N_3756);
xor U5888 (N_5888,N_2330,N_3541);
or U5889 (N_5889,N_2661,N_3527);
and U5890 (N_5890,N_3641,N_3676);
nand U5891 (N_5891,N_2128,N_3984);
nand U5892 (N_5892,N_2063,N_2629);
xor U5893 (N_5893,N_2970,N_3388);
and U5894 (N_5894,N_3240,N_3985);
and U5895 (N_5895,N_3733,N_2102);
nor U5896 (N_5896,N_3514,N_3399);
or U5897 (N_5897,N_2328,N_3590);
nor U5898 (N_5898,N_3901,N_2546);
and U5899 (N_5899,N_2544,N_3181);
nand U5900 (N_5900,N_2518,N_3993);
nand U5901 (N_5901,N_3743,N_3437);
nor U5902 (N_5902,N_3766,N_2312);
or U5903 (N_5903,N_3338,N_3206);
nor U5904 (N_5904,N_2879,N_3719);
xnor U5905 (N_5905,N_2905,N_3306);
xnor U5906 (N_5906,N_3283,N_2112);
xor U5907 (N_5907,N_3794,N_3864);
or U5908 (N_5908,N_2424,N_3276);
and U5909 (N_5909,N_2966,N_2420);
nor U5910 (N_5910,N_2947,N_2849);
xor U5911 (N_5911,N_3429,N_3652);
and U5912 (N_5912,N_3358,N_3681);
or U5913 (N_5913,N_2345,N_2806);
nor U5914 (N_5914,N_2936,N_3247);
nor U5915 (N_5915,N_2480,N_2384);
and U5916 (N_5916,N_3848,N_2470);
nor U5917 (N_5917,N_2143,N_3264);
nor U5918 (N_5918,N_3975,N_2608);
nor U5919 (N_5919,N_3810,N_2598);
xnor U5920 (N_5920,N_3995,N_3642);
or U5921 (N_5921,N_2744,N_2572);
or U5922 (N_5922,N_2317,N_3268);
or U5923 (N_5923,N_3948,N_2010);
nor U5924 (N_5924,N_3023,N_3564);
nand U5925 (N_5925,N_3884,N_2651);
xor U5926 (N_5926,N_2130,N_2856);
and U5927 (N_5927,N_2405,N_2544);
nor U5928 (N_5928,N_3566,N_3063);
xnor U5929 (N_5929,N_2514,N_2070);
nor U5930 (N_5930,N_3146,N_3714);
nor U5931 (N_5931,N_3012,N_3123);
nand U5932 (N_5932,N_2702,N_2934);
xor U5933 (N_5933,N_2273,N_3994);
nand U5934 (N_5934,N_3721,N_2968);
and U5935 (N_5935,N_3313,N_3382);
and U5936 (N_5936,N_3206,N_3078);
nor U5937 (N_5937,N_3222,N_2182);
or U5938 (N_5938,N_2095,N_2049);
nand U5939 (N_5939,N_3272,N_3765);
xor U5940 (N_5940,N_2528,N_2416);
nand U5941 (N_5941,N_3366,N_2251);
nor U5942 (N_5942,N_2792,N_2740);
xnor U5943 (N_5943,N_2300,N_2284);
or U5944 (N_5944,N_3702,N_2076);
nand U5945 (N_5945,N_2864,N_2882);
and U5946 (N_5946,N_3307,N_3614);
nor U5947 (N_5947,N_2530,N_2690);
and U5948 (N_5948,N_2747,N_3550);
and U5949 (N_5949,N_3773,N_3610);
and U5950 (N_5950,N_3805,N_2628);
or U5951 (N_5951,N_3704,N_3999);
nor U5952 (N_5952,N_2815,N_2365);
and U5953 (N_5953,N_3273,N_2344);
nand U5954 (N_5954,N_3208,N_3143);
nor U5955 (N_5955,N_3346,N_2258);
nand U5956 (N_5956,N_2702,N_2862);
and U5957 (N_5957,N_3105,N_3563);
nor U5958 (N_5958,N_2541,N_3597);
or U5959 (N_5959,N_3285,N_2443);
and U5960 (N_5960,N_3827,N_3053);
nand U5961 (N_5961,N_2646,N_2621);
xnor U5962 (N_5962,N_3414,N_2047);
nand U5963 (N_5963,N_2427,N_3776);
or U5964 (N_5964,N_3095,N_3105);
nor U5965 (N_5965,N_3789,N_2200);
nand U5966 (N_5966,N_2377,N_2904);
nand U5967 (N_5967,N_3369,N_2124);
nor U5968 (N_5968,N_3151,N_2926);
and U5969 (N_5969,N_2487,N_3658);
xor U5970 (N_5970,N_3486,N_3396);
nor U5971 (N_5971,N_2037,N_2305);
nor U5972 (N_5972,N_2244,N_2067);
and U5973 (N_5973,N_2059,N_3773);
xor U5974 (N_5974,N_3085,N_3413);
xor U5975 (N_5975,N_2794,N_3249);
nor U5976 (N_5976,N_2872,N_2837);
nand U5977 (N_5977,N_3505,N_3587);
or U5978 (N_5978,N_3311,N_2735);
nand U5979 (N_5979,N_3034,N_3237);
xor U5980 (N_5980,N_2073,N_3189);
and U5981 (N_5981,N_2556,N_2389);
nor U5982 (N_5982,N_3357,N_3845);
and U5983 (N_5983,N_2537,N_2483);
xor U5984 (N_5984,N_3631,N_2368);
xor U5985 (N_5985,N_2977,N_3157);
xnor U5986 (N_5986,N_3549,N_3856);
nand U5987 (N_5987,N_3792,N_3881);
nand U5988 (N_5988,N_3106,N_3772);
nor U5989 (N_5989,N_3204,N_3480);
nand U5990 (N_5990,N_3498,N_2766);
nor U5991 (N_5991,N_3311,N_2017);
xor U5992 (N_5992,N_2291,N_3184);
or U5993 (N_5993,N_3965,N_3307);
xor U5994 (N_5994,N_3537,N_2958);
and U5995 (N_5995,N_3281,N_3295);
nor U5996 (N_5996,N_3503,N_2701);
xor U5997 (N_5997,N_2464,N_2490);
or U5998 (N_5998,N_2489,N_3696);
or U5999 (N_5999,N_2442,N_3870);
nor U6000 (N_6000,N_5015,N_4067);
nand U6001 (N_6001,N_4860,N_4702);
xor U6002 (N_6002,N_4989,N_4334);
nor U6003 (N_6003,N_5089,N_4612);
or U6004 (N_6004,N_4752,N_5893);
and U6005 (N_6005,N_4948,N_4920);
xnor U6006 (N_6006,N_4943,N_5624);
xnor U6007 (N_6007,N_4749,N_5457);
nand U6008 (N_6008,N_4834,N_4518);
or U6009 (N_6009,N_4429,N_4293);
xnor U6010 (N_6010,N_5864,N_4157);
and U6011 (N_6011,N_5156,N_5065);
nor U6012 (N_6012,N_4730,N_4022);
xnor U6013 (N_6013,N_5276,N_4999);
xor U6014 (N_6014,N_4421,N_5296);
xor U6015 (N_6015,N_5758,N_5660);
or U6016 (N_6016,N_5066,N_5420);
nor U6017 (N_6017,N_5990,N_4362);
nand U6018 (N_6018,N_5506,N_5687);
xnor U6019 (N_6019,N_5251,N_5847);
nand U6020 (N_6020,N_4300,N_5496);
xnor U6021 (N_6021,N_4212,N_4141);
or U6022 (N_6022,N_4333,N_5837);
xnor U6023 (N_6023,N_5057,N_5610);
nand U6024 (N_6024,N_5832,N_5281);
or U6025 (N_6025,N_5612,N_5862);
xnor U6026 (N_6026,N_4913,N_4604);
and U6027 (N_6027,N_5934,N_4469);
and U6028 (N_6028,N_4205,N_4158);
or U6029 (N_6029,N_4955,N_5717);
or U6030 (N_6030,N_4383,N_5080);
xnor U6031 (N_6031,N_4974,N_5374);
xor U6032 (N_6032,N_4688,N_4657);
nor U6033 (N_6033,N_4084,N_5663);
xnor U6034 (N_6034,N_4886,N_4456);
nand U6035 (N_6035,N_4000,N_4678);
nand U6036 (N_6036,N_4896,N_4583);
and U6037 (N_6037,N_5931,N_5627);
or U6038 (N_6038,N_5779,N_4237);
xor U6039 (N_6039,N_4673,N_5607);
nor U6040 (N_6040,N_5335,N_4203);
or U6041 (N_6041,N_4406,N_4757);
xor U6042 (N_6042,N_5565,N_4168);
xnor U6043 (N_6043,N_5725,N_5407);
nand U6044 (N_6044,N_4751,N_4940);
and U6045 (N_6045,N_4634,N_4545);
xor U6046 (N_6046,N_5652,N_4802);
xor U6047 (N_6047,N_5641,N_5176);
and U6048 (N_6048,N_5812,N_5474);
xnor U6049 (N_6049,N_5170,N_5428);
and U6050 (N_6050,N_5333,N_5291);
nor U6051 (N_6051,N_5962,N_4485);
nand U6052 (N_6052,N_4269,N_5716);
nor U6053 (N_6053,N_4031,N_5897);
nand U6054 (N_6054,N_4180,N_5006);
xor U6055 (N_6055,N_5238,N_5554);
or U6056 (N_6056,N_5707,N_4289);
and U6057 (N_6057,N_5178,N_5871);
nand U6058 (N_6058,N_5194,N_4097);
nand U6059 (N_6059,N_4626,N_4295);
nand U6060 (N_6060,N_4102,N_4761);
nor U6061 (N_6061,N_4987,N_5566);
nor U6062 (N_6062,N_5120,N_5375);
nor U6063 (N_6063,N_4240,N_5372);
nor U6064 (N_6064,N_4239,N_4019);
xnor U6065 (N_6065,N_4575,N_5289);
xor U6066 (N_6066,N_4745,N_4932);
nor U6067 (N_6067,N_5785,N_4951);
xnor U6068 (N_6068,N_4096,N_4428);
and U6069 (N_6069,N_5932,N_4550);
or U6070 (N_6070,N_5094,N_5340);
or U6071 (N_6071,N_5155,N_5219);
or U6072 (N_6072,N_4714,N_4511);
nor U6073 (N_6073,N_5086,N_4907);
nor U6074 (N_6074,N_5090,N_4915);
and U6075 (N_6075,N_5041,N_4361);
or U6076 (N_6076,N_4326,N_4347);
nor U6077 (N_6077,N_4670,N_5043);
nand U6078 (N_6078,N_5682,N_4762);
nand U6079 (N_6079,N_5907,N_4033);
nor U6080 (N_6080,N_4595,N_5757);
nand U6081 (N_6081,N_5708,N_5764);
and U6082 (N_6082,N_4549,N_5952);
nand U6083 (N_6083,N_5227,N_4044);
xor U6084 (N_6084,N_4717,N_5456);
xnor U6085 (N_6085,N_5819,N_4687);
xor U6086 (N_6086,N_4558,N_5298);
and U6087 (N_6087,N_5587,N_4181);
nor U6088 (N_6088,N_4538,N_4863);
nor U6089 (N_6089,N_4779,N_5017);
and U6090 (N_6090,N_4233,N_4439);
xor U6091 (N_6091,N_5772,N_4387);
and U6092 (N_6092,N_5315,N_5339);
nand U6093 (N_6093,N_5911,N_4658);
nor U6094 (N_6094,N_5577,N_5835);
and U6095 (N_6095,N_5891,N_5697);
xnor U6096 (N_6096,N_4872,N_5856);
or U6097 (N_6097,N_4007,N_5834);
xor U6098 (N_6098,N_5811,N_4103);
nand U6099 (N_6099,N_5807,N_4190);
and U6100 (N_6100,N_4804,N_5241);
or U6101 (N_6101,N_4993,N_4458);
or U6102 (N_6102,N_5525,N_5505);
and U6103 (N_6103,N_5489,N_5849);
or U6104 (N_6104,N_5000,N_4394);
nor U6105 (N_6105,N_4153,N_5596);
nor U6106 (N_6106,N_5626,N_4949);
or U6107 (N_6107,N_5396,N_5463);
or U6108 (N_6108,N_4580,N_5154);
nor U6109 (N_6109,N_4013,N_5113);
nor U6110 (N_6110,N_5352,N_5801);
nand U6111 (N_6111,N_4017,N_4480);
and U6112 (N_6112,N_5974,N_4748);
nor U6113 (N_6113,N_4106,N_4507);
nand U6114 (N_6114,N_5752,N_4128);
nand U6115 (N_6115,N_5431,N_4009);
nand U6116 (N_6116,N_4728,N_5160);
xnor U6117 (N_6117,N_5853,N_4194);
nor U6118 (N_6118,N_4668,N_5198);
xor U6119 (N_6119,N_4767,N_4246);
xnor U6120 (N_6120,N_4769,N_4214);
nor U6121 (N_6121,N_4266,N_5132);
or U6122 (N_6122,N_4320,N_4297);
xnor U6123 (N_6123,N_4488,N_5715);
xnor U6124 (N_6124,N_5824,N_5423);
or U6125 (N_6125,N_5693,N_5355);
nor U6126 (N_6126,N_4392,N_5625);
and U6127 (N_6127,N_5747,N_4966);
xnor U6128 (N_6128,N_5207,N_5751);
and U6129 (N_6129,N_4969,N_4746);
xor U6130 (N_6130,N_4837,N_4378);
and U6131 (N_6131,N_4039,N_4897);
nand U6132 (N_6132,N_5531,N_4766);
xor U6133 (N_6133,N_5353,N_4308);
xor U6134 (N_6134,N_5696,N_4003);
nor U6135 (N_6135,N_4491,N_4950);
and U6136 (N_6136,N_5600,N_4072);
or U6137 (N_6137,N_5584,N_4909);
nor U6138 (N_6138,N_5304,N_4736);
and U6139 (N_6139,N_5710,N_5988);
nand U6140 (N_6140,N_5808,N_5426);
nor U6141 (N_6141,N_5754,N_5323);
and U6142 (N_6142,N_4139,N_5368);
and U6143 (N_6143,N_4741,N_4043);
and U6144 (N_6144,N_4747,N_5258);
nor U6145 (N_6145,N_4628,N_5214);
and U6146 (N_6146,N_4083,N_5024);
and U6147 (N_6147,N_5037,N_5597);
and U6148 (N_6148,N_4134,N_4829);
nor U6149 (N_6149,N_5437,N_4119);
or U6150 (N_6150,N_4548,N_4841);
and U6151 (N_6151,N_4881,N_4242);
or U6152 (N_6152,N_5602,N_4880);
or U6153 (N_6153,N_5191,N_4792);
or U6154 (N_6154,N_4245,N_4776);
nor U6155 (N_6155,N_5059,N_4547);
nor U6156 (N_6156,N_4912,N_5616);
xnor U6157 (N_6157,N_5760,N_4529);
xor U6158 (N_6158,N_4322,N_5500);
xor U6159 (N_6159,N_4226,N_4996);
xnor U6160 (N_6160,N_5117,N_5783);
nand U6161 (N_6161,N_4521,N_5071);
nor U6162 (N_6162,N_5076,N_5946);
xor U6163 (N_6163,N_5691,N_5723);
and U6164 (N_6164,N_4182,N_5153);
and U6165 (N_6165,N_5288,N_4539);
or U6166 (N_6166,N_5392,N_4613);
nor U6167 (N_6167,N_5111,N_5999);
xnor U6168 (N_6168,N_5486,N_4086);
nor U6169 (N_6169,N_5308,N_5628);
nand U6170 (N_6170,N_4442,N_5929);
nor U6171 (N_6171,N_4551,N_5414);
and U6172 (N_6172,N_5150,N_4325);
or U6173 (N_6173,N_4016,N_5350);
and U6174 (N_6174,N_5133,N_4928);
nor U6175 (N_6175,N_4389,N_5441);
or U6176 (N_6176,N_4643,N_5380);
nand U6177 (N_6177,N_4649,N_4399);
nor U6178 (N_6178,N_5439,N_4568);
and U6179 (N_6179,N_5875,N_4025);
or U6180 (N_6180,N_4369,N_5800);
xnor U6181 (N_6181,N_5888,N_5885);
nand U6182 (N_6182,N_4419,N_4712);
nand U6183 (N_6183,N_5014,N_5733);
nand U6184 (N_6184,N_4621,N_4506);
xor U6185 (N_6185,N_4965,N_5035);
and U6186 (N_6186,N_5055,N_4532);
xor U6187 (N_6187,N_5249,N_5520);
xor U6188 (N_6188,N_4482,N_5771);
xor U6189 (N_6189,N_4682,N_5346);
or U6190 (N_6190,N_4349,N_5993);
xnor U6191 (N_6191,N_4287,N_4663);
nor U6192 (N_6192,N_5967,N_5432);
nand U6193 (N_6193,N_5937,N_5787);
nand U6194 (N_6194,N_4337,N_4352);
nand U6195 (N_6195,N_4574,N_5164);
nor U6196 (N_6196,N_4081,N_5205);
or U6197 (N_6197,N_4274,N_4785);
nand U6198 (N_6198,N_4567,N_5955);
nor U6199 (N_6199,N_5821,N_4654);
xor U6200 (N_6200,N_4315,N_5539);
nand U6201 (N_6201,N_4402,N_5443);
xor U6202 (N_6202,N_4151,N_5796);
xnor U6203 (N_6203,N_4952,N_5983);
and U6204 (N_6204,N_4534,N_5773);
xor U6205 (N_6205,N_4890,N_4065);
and U6206 (N_6206,N_5215,N_4639);
or U6207 (N_6207,N_4608,N_4184);
xnor U6208 (N_6208,N_4892,N_4027);
nand U6209 (N_6209,N_4939,N_5363);
and U6210 (N_6210,N_4684,N_4887);
and U6211 (N_6211,N_5918,N_5501);
nor U6212 (N_6212,N_5243,N_4998);
nand U6213 (N_6213,N_4201,N_5775);
nand U6214 (N_6214,N_5451,N_5151);
and U6215 (N_6215,N_5868,N_5609);
and U6216 (N_6216,N_5574,N_4859);
xnor U6217 (N_6217,N_5533,N_4962);
and U6218 (N_6218,N_4426,N_5411);
nor U6219 (N_6219,N_4196,N_4244);
or U6220 (N_6220,N_5376,N_5467);
nor U6221 (N_6221,N_5012,N_5662);
xnor U6222 (N_6222,N_4847,N_5157);
and U6223 (N_6223,N_4268,N_4659);
or U6224 (N_6224,N_4319,N_4306);
xnor U6225 (N_6225,N_5804,N_4927);
and U6226 (N_6226,N_5360,N_5831);
or U6227 (N_6227,N_4318,N_4342);
or U6228 (N_6228,N_5973,N_5292);
nand U6229 (N_6229,N_5255,N_4459);
xnor U6230 (N_6230,N_4395,N_5852);
nor U6231 (N_6231,N_4596,N_4795);
and U6232 (N_6232,N_4652,N_4155);
nand U6233 (N_6233,N_5571,N_5594);
and U6234 (N_6234,N_5608,N_4453);
and U6235 (N_6235,N_5985,N_4411);
nor U6236 (N_6236,N_5870,N_4808);
nand U6237 (N_6237,N_4372,N_5913);
and U6238 (N_6238,N_5643,N_4816);
xor U6239 (N_6239,N_4824,N_4270);
nand U6240 (N_6240,N_5809,N_4814);
nand U6241 (N_6241,N_5644,N_4466);
and U6242 (N_6242,N_5667,N_4755);
xor U6243 (N_6243,N_5711,N_5449);
xor U6244 (N_6244,N_4026,N_4450);
nor U6245 (N_6245,N_5138,N_5247);
nand U6246 (N_6246,N_4537,N_4467);
nand U6247 (N_6247,N_4563,N_5568);
nor U6248 (N_6248,N_4137,N_5031);
and U6249 (N_6249,N_5767,N_5382);
nand U6250 (N_6250,N_5455,N_5127);
nor U6251 (N_6251,N_4852,N_5307);
nand U6252 (N_6252,N_4058,N_5054);
xnor U6253 (N_6253,N_5234,N_5873);
and U6254 (N_6254,N_4207,N_4720);
nand U6255 (N_6255,N_5692,N_4844);
nor U6256 (N_6256,N_4777,N_5254);
or U6257 (N_6257,N_5200,N_4475);
or U6258 (N_6258,N_5570,N_5684);
nand U6259 (N_6259,N_4647,N_5422);
nor U6260 (N_6260,N_5393,N_4112);
nor U6261 (N_6261,N_5544,N_4864);
nor U6262 (N_6262,N_4523,N_5399);
and U6263 (N_6263,N_5706,N_5010);
nor U6264 (N_6264,N_5297,N_4407);
nor U6265 (N_6265,N_4803,N_5362);
nor U6266 (N_6266,N_5421,N_5485);
and U6267 (N_6267,N_5397,N_4671);
nand U6268 (N_6268,N_4267,N_4183);
xnor U6269 (N_6269,N_4069,N_5846);
nand U6270 (N_6270,N_5330,N_5105);
nand U6271 (N_6271,N_4020,N_5978);
or U6272 (N_6272,N_5147,N_4206);
nand U6273 (N_6273,N_5598,N_5018);
or U6274 (N_6274,N_5429,N_4447);
nor U6275 (N_6275,N_5734,N_5336);
or U6276 (N_6276,N_4105,N_5188);
nor U6277 (N_6277,N_5620,N_4377);
xor U6278 (N_6278,N_5477,N_4679);
nor U6279 (N_6279,N_5799,N_5528);
or U6280 (N_6280,N_4208,N_4343);
xnor U6281 (N_6281,N_4499,N_4651);
xor U6282 (N_6282,N_5904,N_5475);
or U6283 (N_6283,N_5581,N_5367);
nor U6284 (N_6284,N_5008,N_5886);
xor U6285 (N_6285,N_4142,N_4540);
nand U6286 (N_6286,N_5933,N_5034);
or U6287 (N_6287,N_5369,N_4629);
or U6288 (N_6288,N_4988,N_4937);
and U6289 (N_6289,N_4648,N_4850);
nor U6290 (N_6290,N_5152,N_4577);
or U6291 (N_6291,N_4172,N_5736);
or U6292 (N_6292,N_5948,N_5358);
nor U6293 (N_6293,N_5617,N_4553);
or U6294 (N_6294,N_4030,N_4211);
and U6295 (N_6295,N_5256,N_5269);
nand U6296 (N_6296,N_5550,N_5097);
or U6297 (N_6297,N_5357,N_4616);
and U6298 (N_6298,N_5201,N_5348);
and U6299 (N_6299,N_5469,N_5329);
xor U6300 (N_6300,N_5665,N_4520);
nor U6301 (N_6301,N_5072,N_5067);
nand U6302 (N_6302,N_4484,N_5975);
or U6303 (N_6303,N_5714,N_4771);
and U6304 (N_6304,N_5746,N_5344);
nor U6305 (N_6305,N_4980,N_5877);
and U6306 (N_6306,N_5483,N_4353);
xor U6307 (N_6307,N_5895,N_5497);
nand U6308 (N_6308,N_5592,N_4590);
nor U6309 (N_6309,N_4159,N_4535);
nor U6310 (N_6310,N_5741,N_4432);
nand U6311 (N_6311,N_5239,N_4486);
nand U6312 (N_6312,N_4522,N_5190);
nor U6313 (N_6313,N_5220,N_4586);
and U6314 (N_6314,N_5324,N_5373);
and U6315 (N_6315,N_4059,N_4990);
or U6316 (N_6316,N_4891,N_5248);
xor U6317 (N_6317,N_5670,N_5698);
and U6318 (N_6318,N_5813,N_5939);
and U6319 (N_6319,N_5593,N_5576);
and U6320 (N_6320,N_4440,N_5126);
or U6321 (N_6321,N_5503,N_5518);
and U6322 (N_6322,N_4252,N_5588);
nand U6323 (N_6323,N_5954,N_4686);
or U6324 (N_6324,N_5079,N_5640);
or U6325 (N_6325,N_5022,N_4089);
or U6326 (N_6326,N_4052,N_5078);
and U6327 (N_6327,N_4832,N_5471);
or U6328 (N_6328,N_5106,N_5240);
and U6329 (N_6329,N_5720,N_4276);
or U6330 (N_6330,N_4189,N_4386);
and U6331 (N_6331,N_5996,N_5664);
nor U6332 (N_6332,N_4476,N_5519);
or U6333 (N_6333,N_4519,N_4866);
nand U6334 (N_6334,N_4936,N_4054);
nor U6335 (N_6335,N_5280,N_5135);
nand U6336 (N_6336,N_4725,N_5884);
and U6337 (N_6337,N_5840,N_5514);
xnor U6338 (N_6338,N_4331,N_4781);
and U6339 (N_6339,N_4350,N_4316);
or U6340 (N_6340,N_5211,N_4021);
and U6341 (N_6341,N_4472,N_4517);
nand U6342 (N_6342,N_5305,N_4991);
nand U6343 (N_6343,N_5048,N_5828);
or U6344 (N_6344,N_4994,N_4873);
and U6345 (N_6345,N_5991,N_5633);
xnor U6346 (N_6346,N_4957,N_4820);
nand U6347 (N_6347,N_4130,N_5745);
nor U6348 (N_6348,N_5045,N_5476);
xnor U6349 (N_6349,N_4633,N_4357);
nand U6350 (N_6350,N_5770,N_5964);
nor U6351 (N_6351,N_4774,N_4035);
nand U6352 (N_6352,N_5650,N_5174);
and U6353 (N_6353,N_5653,N_4715);
xnor U6354 (N_6354,N_4301,N_4156);
nor U6355 (N_6355,N_5019,N_4282);
and U6356 (N_6356,N_5074,N_5409);
nor U6357 (N_6357,N_4911,N_4125);
xnor U6358 (N_6358,N_5887,N_5062);
and U6359 (N_6359,N_4573,N_5963);
nor U6360 (N_6360,N_5841,N_5112);
nor U6361 (N_6361,N_5342,N_4840);
or U6362 (N_6362,N_5892,N_4145);
or U6363 (N_6363,N_5548,N_4677);
nand U6364 (N_6364,N_4697,N_5547);
or U6365 (N_6365,N_5534,N_5210);
nor U6366 (N_6366,N_5699,N_5192);
nand U6367 (N_6367,N_5686,N_4006);
nand U6368 (N_6368,N_5642,N_4743);
xnor U6369 (N_6369,N_4216,N_4336);
and U6370 (N_6370,N_5508,N_5825);
xnor U6371 (N_6371,N_5186,N_5002);
or U6372 (N_6372,N_4090,N_5047);
nand U6373 (N_6373,N_4531,N_4129);
nand U6374 (N_6374,N_5246,N_4942);
nor U6375 (N_6375,N_5470,N_5563);
xnor U6376 (N_6376,N_4884,N_5389);
or U6377 (N_6377,N_4764,N_4382);
xnor U6378 (N_6378,N_4505,N_4433);
nor U6379 (N_6379,N_4376,N_4179);
or U6380 (N_6380,N_5977,N_5316);
nor U6381 (N_6381,N_4231,N_4695);
xor U6382 (N_6382,N_4412,N_4441);
nor U6383 (N_6383,N_4265,N_5938);
xnor U6384 (N_6384,N_5599,N_5433);
and U6385 (N_6385,N_4177,N_5016);
nor U6386 (N_6386,N_4722,N_5446);
or U6387 (N_6387,N_5579,N_5004);
and U6388 (N_6388,N_4602,N_4284);
or U6389 (N_6389,N_4676,N_5728);
xor U6390 (N_6390,N_4215,N_4735);
or U6391 (N_6391,N_5143,N_4667);
xnor U6392 (N_6392,N_5702,N_4004);
nand U6393 (N_6393,N_4321,N_5029);
or U6394 (N_6394,N_5386,N_5136);
nand U6395 (N_6395,N_4258,N_5381);
nor U6396 (N_6396,N_5851,N_4838);
or U6397 (N_6397,N_4946,N_5492);
and U6398 (N_6398,N_5666,N_4570);
nand U6399 (N_6399,N_5631,N_5826);
and U6400 (N_6400,N_4597,N_4656);
or U6401 (N_6401,N_5260,N_5553);
nor U6402 (N_6402,N_5349,N_4925);
nor U6403 (N_6403,N_4109,N_5051);
and U6404 (N_6404,N_5790,N_4857);
or U6405 (N_6405,N_5820,N_4554);
xnor U6406 (N_6406,N_5069,N_4191);
nand U6407 (N_6407,N_5134,N_4644);
or U6408 (N_6408,N_4995,N_4446);
xor U6409 (N_6409,N_5253,N_4430);
and U6410 (N_6410,N_5883,N_5119);
nor U6411 (N_6411,N_5647,N_4941);
and U6412 (N_6412,N_4150,N_4147);
or U6413 (N_6413,N_5690,N_4236);
nor U6414 (N_6414,N_4028,N_5959);
nor U6415 (N_6415,N_4904,N_4285);
or U6416 (N_6416,N_5613,N_4960);
xor U6417 (N_6417,N_4140,N_5860);
or U6418 (N_6418,N_5075,N_4977);
or U6419 (N_6419,N_4423,N_5793);
xor U6420 (N_6420,N_5524,N_4826);
nand U6421 (N_6421,N_5654,N_4463);
and U6422 (N_6422,N_5272,N_5591);
xnor U6423 (N_6423,N_5753,N_5992);
nand U6424 (N_6424,N_4010,N_4954);
nor U6425 (N_6425,N_4471,N_4045);
nor U6426 (N_6426,N_5413,N_4351);
xor U6427 (N_6427,N_4641,N_4136);
nor U6428 (N_6428,N_4964,N_4972);
and U6429 (N_6429,N_4217,N_4615);
and U6430 (N_6430,N_5115,N_4403);
and U6431 (N_6431,N_5604,N_5928);
nand U6432 (N_6432,N_4074,N_5614);
or U6433 (N_6433,N_5095,N_5064);
nor U6434 (N_6434,N_5552,N_5096);
nand U6435 (N_6435,N_4229,N_4924);
xnor U6436 (N_6436,N_4259,N_4631);
nand U6437 (N_6437,N_4313,N_5158);
nand U6438 (N_6438,N_4503,N_5264);
xnor U6439 (N_6439,N_5947,N_5081);
and U6440 (N_6440,N_5914,N_5924);
nand U6441 (N_6441,N_5951,N_4302);
nor U6442 (N_6442,N_5021,N_4164);
or U6443 (N_6443,N_5273,N_4510);
or U6444 (N_6444,N_5371,N_5060);
and U6445 (N_6445,N_5347,N_4784);
or U6446 (N_6446,N_4589,N_5123);
and U6447 (N_6447,N_5259,N_5639);
and U6448 (N_6448,N_4711,N_4750);
nand U6449 (N_6449,N_5495,N_5629);
or U6450 (N_6450,N_5365,N_5769);
nand U6451 (N_6451,N_4445,N_4001);
and U6452 (N_6452,N_5848,N_5722);
or U6453 (N_6453,N_5540,N_4359);
nor U6454 (N_6454,N_4899,N_5867);
or U6455 (N_6455,N_5444,N_4740);
and U6456 (N_6456,N_4487,N_4727);
nor U6457 (N_6457,N_4034,N_5791);
nor U6458 (N_6458,N_4257,N_4818);
xor U6459 (N_6459,N_5168,N_5322);
or U6460 (N_6460,N_4650,N_5865);
nand U6461 (N_6461,N_4513,N_5645);
nor U6462 (N_6462,N_5944,N_5318);
and U6463 (N_6463,N_5169,N_5510);
nand U6464 (N_6464,N_4875,N_5965);
nand U6465 (N_6465,N_4794,N_5523);
and U6466 (N_6466,N_4833,N_4390);
xnor U6467 (N_6467,N_5786,N_4391);
or U6468 (N_6468,N_5313,N_5225);
nor U6469 (N_6469,N_4366,N_5843);
nor U6470 (N_6470,N_5245,N_4056);
xor U6471 (N_6471,N_4424,N_4719);
nor U6472 (N_6472,N_5780,N_5181);
xnor U6473 (N_6473,N_4465,N_5649);
xor U6474 (N_6474,N_4489,N_5233);
xor U6475 (N_6475,N_5391,N_4061);
or U6476 (N_6476,N_4296,N_5845);
nor U6477 (N_6477,N_5498,N_5395);
or U6478 (N_6478,N_4576,N_5546);
and U6479 (N_6479,N_5527,N_5726);
and U6480 (N_6480,N_5116,N_5141);
and U6481 (N_6481,N_5104,N_5222);
and U6482 (N_6482,N_5268,N_5310);
and U6483 (N_6483,N_5515,N_5517);
xnor U6484 (N_6484,N_5920,N_5561);
and U6485 (N_6485,N_4425,N_4146);
and U6486 (N_6486,N_5538,N_5634);
nand U6487 (N_6487,N_5761,N_5379);
or U6488 (N_6488,N_5418,N_4883);
nand U6489 (N_6489,N_5674,N_5073);
and U6490 (N_6490,N_4133,N_4638);
nand U6491 (N_6491,N_5208,N_5982);
nand U6492 (N_6492,N_5338,N_4290);
nor U6493 (N_6493,N_5005,N_5481);
nand U6494 (N_6494,N_5301,N_5829);
and U6495 (N_6495,N_4005,N_5989);
and U6496 (N_6496,N_4655,N_4582);
xnor U6497 (N_6497,N_5231,N_4273);
and U6498 (N_6498,N_5488,N_5424);
nor U6499 (N_6499,N_5466,N_5969);
nor U6500 (N_6500,N_5242,N_5712);
or U6501 (N_6501,N_4202,N_5816);
or U6502 (N_6502,N_5774,N_5092);
or U6503 (N_6503,N_4718,N_4514);
and U6504 (N_6504,N_4160,N_4023);
nand U6505 (N_6505,N_4324,N_4032);
nor U6506 (N_6506,N_5167,N_4292);
or U6507 (N_6507,N_4627,N_5854);
and U6508 (N_6508,N_5009,N_5795);
xnor U6509 (N_6509,N_4230,N_5657);
or U6510 (N_6510,N_4552,N_4953);
nor U6511 (N_6511,N_5454,N_4756);
nor U6512 (N_6512,N_5180,N_4232);
nor U6513 (N_6513,N_4219,N_5145);
or U6514 (N_6514,N_5605,N_4490);
xor U6515 (N_6515,N_5257,N_4704);
or U6516 (N_6516,N_5028,N_5209);
nor U6517 (N_6517,N_4477,N_4187);
nand U6518 (N_6518,N_4846,N_4492);
and U6519 (N_6519,N_5619,N_4094);
and U6520 (N_6520,N_4213,N_4874);
nand U6521 (N_6521,N_4599,N_5319);
nor U6522 (N_6522,N_4983,N_5306);
nand U6523 (N_6523,N_4345,N_4801);
and U6524 (N_6524,N_5916,N_4606);
and U6525 (N_6525,N_4787,N_5419);
and U6526 (N_6526,N_4888,N_5683);
xnor U6527 (N_6527,N_4114,N_4311);
nor U6528 (N_6528,N_4858,N_5659);
or U6529 (N_6529,N_4737,N_4481);
and U6530 (N_6530,N_5416,N_4754);
nor U6531 (N_6531,N_4898,N_5270);
and U6532 (N_6532,N_5842,N_4689);
nor U6533 (N_6533,N_5082,N_4922);
nand U6534 (N_6534,N_4821,N_5083);
xor U6535 (N_6535,N_5494,N_5223);
xnor U6536 (N_6536,N_4149,N_4314);
nor U6537 (N_6537,N_5404,N_4468);
xor U6538 (N_6538,N_5695,N_5638);
xor U6539 (N_6539,N_4861,N_5161);
and U6540 (N_6540,N_4600,N_4082);
xnor U6541 (N_6541,N_5427,N_5232);
nand U6542 (N_6542,N_5558,N_4618);
nor U6543 (N_6543,N_4726,N_4504);
xor U6544 (N_6544,N_4380,N_4126);
xnor U6545 (N_6545,N_4339,N_5184);
nor U6546 (N_6546,N_5673,N_5635);
nand U6547 (N_6547,N_4358,N_4209);
nand U6548 (N_6548,N_5994,N_4085);
or U6549 (N_6549,N_4903,N_4981);
nor U6550 (N_6550,N_5880,N_4338);
nor U6551 (N_6551,N_4508,N_4865);
nor U6552 (N_6552,N_4092,N_5900);
nor U6553 (N_6553,N_5855,N_4700);
xnor U6554 (N_6554,N_5675,N_4335);
nor U6555 (N_6555,N_4076,N_4248);
nor U6556 (N_6556,N_5648,N_4780);
and U6557 (N_6557,N_4255,N_4815);
or U6558 (N_6558,N_5142,N_5572);
and U6559 (N_6559,N_4851,N_5926);
or U6560 (N_6560,N_4564,N_4050);
and U6561 (N_6561,N_5910,N_4431);
or U6562 (N_6562,N_4929,N_5742);
xor U6563 (N_6563,N_5468,N_4279);
nor U6564 (N_6564,N_4546,N_4247);
xnor U6565 (N_6565,N_4171,N_4397);
nand U6566 (N_6566,N_4435,N_5956);
and U6567 (N_6567,N_4578,N_4420);
or U6568 (N_6568,N_5630,N_4696);
nand U6569 (N_6569,N_5970,N_4317);
and U6570 (N_6570,N_4976,N_5543);
and U6571 (N_6571,N_4304,N_5925);
nor U6572 (N_6572,N_5244,N_4091);
or U6573 (N_6573,N_5902,N_5440);
nand U6574 (N_6574,N_4323,N_4985);
nand U6575 (N_6575,N_5144,N_4587);
nand U6576 (N_6576,N_5196,N_5729);
nand U6577 (N_6577,N_5114,N_4653);
xor U6578 (N_6578,N_5261,N_5228);
or U6579 (N_6579,N_5903,N_5317);
nor U6580 (N_6580,N_4982,N_5960);
or U6581 (N_6581,N_5011,N_4835);
or U6582 (N_6582,N_4195,N_5309);
or U6583 (N_6583,N_4451,N_4839);
nand U6584 (N_6584,N_5185,N_5236);
nand U6585 (N_6585,N_4854,N_4724);
or U6586 (N_6586,N_5839,N_4227);
nor U6587 (N_6587,N_5882,N_5282);
nand U6588 (N_6588,N_5193,N_5906);
or U6589 (N_6589,N_4734,N_4992);
nor U6590 (N_6590,N_5235,N_5890);
nor U6591 (N_6591,N_5502,N_4410);
and U6592 (N_6592,N_4379,N_5279);
nand U6593 (N_6593,N_5535,N_4415);
and U6594 (N_6594,N_4494,N_4462);
nand U6595 (N_6595,N_4169,N_5398);
nand U6596 (N_6596,N_4895,N_4571);
or U6597 (N_6597,N_4152,N_5575);
and U6598 (N_6598,N_5107,N_5410);
nor U6599 (N_6599,N_4115,N_4685);
xor U6600 (N_6600,N_5345,N_4691);
or U6601 (N_6601,N_4396,N_5504);
and U6602 (N_6602,N_5894,N_5265);
or U6603 (N_6603,N_4642,N_4739);
xor U6604 (N_6604,N_4862,N_5748);
nand U6605 (N_6605,N_4617,N_5285);
or U6606 (N_6606,N_4956,N_4721);
or U6607 (N_6607,N_5312,N_4384);
and U6608 (N_6608,N_4635,N_5480);
or U6609 (N_6609,N_4283,N_4327);
and U6610 (N_6610,N_4303,N_4124);
or U6611 (N_6611,N_5805,N_5266);
nand U6612 (N_6612,N_5122,N_4823);
and U6613 (N_6613,N_5958,N_4278);
and U6614 (N_6614,N_4692,N_5275);
nand U6615 (N_6615,N_4709,N_5321);
xor U6616 (N_6616,N_5300,N_4515);
nand U6617 (N_6617,N_4791,N_5283);
xor U6618 (N_6618,N_4701,N_4370);
nor U6619 (N_6619,N_4099,N_4116);
xnor U6620 (N_6620,N_5402,N_4572);
xnor U6621 (N_6621,N_5464,N_4204);
or U6622 (N_6622,N_5478,N_4805);
or U6623 (N_6623,N_4078,N_4789);
nand U6624 (N_6624,N_4889,N_5703);
xnor U6625 (N_6625,N_4830,N_4607);
or U6626 (N_6626,N_5487,N_5606);
xor U6627 (N_6627,N_4914,N_5859);
nor U6628 (N_6628,N_5085,N_4367);
nor U6629 (N_6629,N_5327,N_5023);
or U6630 (N_6630,N_5130,N_5462);
nor U6631 (N_6631,N_4444,N_5033);
xor U6632 (N_6632,N_4710,N_5103);
or U6633 (N_6633,N_4309,N_5459);
and U6634 (N_6634,N_5953,N_4063);
or U6635 (N_6635,N_4434,N_5452);
and U6636 (N_6636,N_5833,N_4630);
and U6637 (N_6637,N_5632,N_5776);
or U6638 (N_6638,N_5098,N_4048);
or U6639 (N_6639,N_5325,N_4250);
nor U6640 (N_6640,N_5569,N_4664);
nand U6641 (N_6641,N_4132,N_4261);
or U6642 (N_6642,N_4393,N_5125);
xor U6643 (N_6643,N_5197,N_5435);
xor U6644 (N_6644,N_5230,N_4416);
xnor U6645 (N_6645,N_5199,N_5189);
xnor U6646 (N_6646,N_5766,N_5794);
or U6647 (N_6647,N_5149,N_4812);
and U6648 (N_6648,N_5084,N_5915);
nand U6649 (N_6649,N_5968,N_4516);
nor U6650 (N_6650,N_4690,N_4770);
nor U6651 (N_6651,N_5087,N_4388);
or U6652 (N_6652,N_4592,N_4024);
nor U6653 (N_6653,N_4773,N_5252);
xnor U6654 (N_6654,N_5585,N_5896);
nor U6655 (N_6655,N_5936,N_5919);
nand U6656 (N_6656,N_5213,N_4193);
and U6657 (N_6657,N_4111,N_5179);
xor U6658 (N_6658,N_5658,N_5511);
or U6659 (N_6659,N_5961,N_5366);
and U6660 (N_6660,N_5493,N_4849);
nor U6661 (N_6661,N_4249,N_4371);
or U6662 (N_6662,N_4528,N_5159);
nor U6663 (N_6663,N_4694,N_4042);
and U6664 (N_6664,N_4460,N_5430);
xor U6665 (N_6665,N_5830,N_4530);
nand U6666 (N_6666,N_4713,N_5636);
nor U6667 (N_6667,N_4275,N_5930);
or U6668 (N_6668,N_5778,N_4723);
and U6669 (N_6669,N_4055,N_5491);
nor U6670 (N_6670,N_4744,N_5737);
or U6671 (N_6671,N_5986,N_4665);
nand U6672 (N_6672,N_4075,N_5484);
or U6673 (N_6673,N_5957,N_4729);
nand U6674 (N_6674,N_4798,N_5050);
nand U6675 (N_6675,N_4921,N_4144);
nand U6676 (N_6676,N_4107,N_5689);
nor U6677 (N_6677,N_5020,N_4855);
nand U6678 (N_6678,N_5881,N_5063);
or U6679 (N_6679,N_4683,N_4660);
and U6680 (N_6680,N_5204,N_5995);
nand U6681 (N_6681,N_5013,N_5172);
or U6682 (N_6682,N_5128,N_5863);
xor U6683 (N_6683,N_5445,N_4260);
nor U6684 (N_6684,N_4218,N_4108);
nand U6685 (N_6685,N_5718,N_5879);
xnor U6686 (N_6686,N_5530,N_4272);
xnor U6687 (N_6687,N_4401,N_5110);
and U6688 (N_6688,N_5030,N_5387);
or U6689 (N_6689,N_5768,N_4501);
and U6690 (N_6690,N_4186,N_4173);
xnor U6691 (N_6691,N_4011,N_4036);
nand U6692 (N_6692,N_5490,N_4448);
or U6693 (N_6693,N_4280,N_5438);
xor U6694 (N_6694,N_5676,N_4271);
nand U6695 (N_6695,N_4104,N_5756);
xor U6696 (N_6696,N_4541,N_4646);
nand U6697 (N_6697,N_4645,N_5040);
xor U6698 (N_6698,N_5221,N_4672);
and U6699 (N_6699,N_5262,N_4675);
nand U6700 (N_6700,N_4971,N_4931);
nand U6701 (N_6701,N_5042,N_4291);
nor U6702 (N_6702,N_5146,N_4605);
and U6703 (N_6703,N_5583,N_4916);
or U6704 (N_6704,N_4385,N_5278);
xnor U6705 (N_6705,N_5044,N_4251);
xor U6706 (N_6706,N_5226,N_5777);
nor U6707 (N_6707,N_5651,N_4312);
nor U6708 (N_6708,N_4262,N_5595);
nand U6709 (N_6709,N_4356,N_5479);
nor U6710 (N_6710,N_5056,N_5049);
nor U6711 (N_6711,N_5981,N_5731);
and U6712 (N_6712,N_5166,N_5601);
nand U6713 (N_6713,N_5759,N_5331);
nor U6714 (N_6714,N_4422,N_5417);
xor U6715 (N_6715,N_4708,N_4414);
or U6716 (N_6716,N_4329,N_4197);
xor U6717 (N_6717,N_4087,N_5603);
or U6718 (N_6718,N_5537,N_5980);
nand U6719 (N_6719,N_4926,N_5704);
xor U6720 (N_6720,N_4500,N_4871);
nor U6721 (N_6721,N_4527,N_4223);
and U6722 (N_6722,N_5762,N_5137);
xnor U6723 (N_6723,N_5337,N_4167);
nand U6724 (N_6724,N_4161,N_5656);
and U6725 (N_6725,N_5450,N_5898);
xnor U6726 (N_6726,N_4101,N_4967);
or U6727 (N_6727,N_5680,N_5447);
and U6728 (N_6728,N_4536,N_4800);
nor U6729 (N_6729,N_4008,N_5838);
or U6730 (N_6730,N_5412,N_5749);
or U6731 (N_6731,N_4878,N_4581);
or U6732 (N_6732,N_4984,N_5341);
nand U6733 (N_6733,N_5735,N_5987);
and U6734 (N_6734,N_5555,N_4037);
and U6735 (N_6735,N_5343,N_5274);
nor U6736 (N_6736,N_4170,N_5171);
xor U6737 (N_6737,N_4057,N_4228);
or U6738 (N_6738,N_5872,N_4264);
or U6739 (N_6739,N_4680,N_5844);
or U6740 (N_6740,N_5556,N_5303);
nor U6741 (N_6741,N_5070,N_5732);
nand U6742 (N_6742,N_5765,N_5669);
and U6743 (N_6743,N_4224,N_4073);
or U6744 (N_6744,N_4341,N_4963);
or U6745 (N_6745,N_5237,N_4162);
nor U6746 (N_6746,N_5541,N_4122);
xor U6747 (N_6747,N_4666,N_5131);
nand U6748 (N_6748,N_4046,N_5655);
and U6749 (N_6749,N_5763,N_4797);
or U6750 (N_6750,N_5173,N_5425);
xor U6751 (N_6751,N_5782,N_4012);
xnor U6752 (N_6752,N_5562,N_4294);
and U6753 (N_6753,N_5332,N_4930);
and U6754 (N_6754,N_5405,N_4002);
and U6755 (N_6755,N_4944,N_4062);
and U6756 (N_6756,N_5377,N_4917);
xor U6757 (N_6757,N_4533,N_4555);
xor U6758 (N_6758,N_4355,N_4699);
nand U6759 (N_6759,N_5679,N_5293);
nand U6760 (N_6760,N_4934,N_4938);
nand U6761 (N_6761,N_4254,N_5836);
xor U6762 (N_6762,N_5390,N_4765);
nand U6763 (N_6763,N_4457,N_4674);
or U6764 (N_6764,N_5182,N_5077);
nand U6765 (N_6765,N_4298,N_5061);
and U6766 (N_6766,N_4138,N_5351);
nor U6767 (N_6767,N_4768,N_5364);
nor U6768 (N_6768,N_4733,N_4417);
xor U6769 (N_6769,N_4598,N_5195);
and U6770 (N_6770,N_4968,N_5068);
nand U6771 (N_6771,N_4344,N_4763);
or U6772 (N_6772,N_4856,N_4877);
xnor U6773 (N_6773,N_5950,N_4443);
or U6774 (N_6774,N_5806,N_5941);
or U6775 (N_6775,N_5781,N_4093);
nand U6776 (N_6776,N_4070,N_5026);
nand U6777 (N_6777,N_5730,N_5677);
or U6778 (N_6778,N_4121,N_5559);
xor U6779 (N_6779,N_5637,N_4742);
nand U6780 (N_6780,N_4565,N_5250);
and U6781 (N_6781,N_4077,N_4961);
xor U6782 (N_6782,N_5217,N_4788);
nor U6783 (N_6783,N_4263,N_5784);
or U6784 (N_6784,N_4822,N_4619);
or U6785 (N_6785,N_4958,N_5175);
xor U6786 (N_6786,N_5909,N_4330);
or U6787 (N_6787,N_5814,N_5869);
or U6788 (N_6788,N_4758,N_4375);
nand U6789 (N_6789,N_5719,N_4579);
or U6790 (N_6790,N_4610,N_4560);
nand U6791 (N_6791,N_4584,N_5557);
or U6792 (N_6792,N_4174,N_4906);
nand U6793 (N_6793,N_4935,N_5536);
nor U6794 (N_6794,N_4543,N_5388);
and U6795 (N_6795,N_5681,N_4176);
nor U6796 (N_6796,N_4561,N_4188);
xor U6797 (N_6797,N_4409,N_4614);
and U6798 (N_6798,N_5036,N_4902);
or U6799 (N_6799,N_4669,N_5713);
or U6800 (N_6800,N_4436,N_4225);
xor U6801 (N_6801,N_5139,N_4772);
nand U6802 (N_6802,N_4707,N_4894);
nand U6803 (N_6803,N_4848,N_5738);
xor U6804 (N_6804,N_5507,N_4060);
xor U6805 (N_6805,N_5100,N_5453);
xor U6806 (N_6806,N_4845,N_5727);
nor U6807 (N_6807,N_4199,N_4843);
nor U6808 (N_6808,N_4286,N_4277);
nor U6809 (N_6809,N_4398,N_5385);
or U6810 (N_6810,N_4661,N_4810);
or U6811 (N_6811,N_4110,N_4365);
and U6812 (N_6812,N_4256,N_4559);
and U6813 (N_6813,N_4623,N_5979);
nand U6814 (N_6814,N_5688,N_5899);
and U6815 (N_6815,N_5823,N_5046);
and U6816 (N_6816,N_4910,N_5921);
nor U6817 (N_6817,N_4098,N_5586);
and U6818 (N_6818,N_5140,N_5578);
and U6819 (N_6819,N_5685,N_5320);
or U6820 (N_6820,N_4783,N_4842);
nor U6821 (N_6821,N_5740,N_5672);
and U6822 (N_6822,N_4799,N_5943);
xnor U6823 (N_6823,N_4113,N_5984);
nand U6824 (N_6824,N_5827,N_5001);
nor U6825 (N_6825,N_4900,N_5803);
and U6826 (N_6826,N_4310,N_4868);
nand U6827 (N_6827,N_5271,N_5905);
nor U6828 (N_6828,N_4811,N_5750);
nand U6829 (N_6829,N_5705,N_5922);
nor U6830 (N_6830,N_4234,N_4408);
or U6831 (N_6831,N_4876,N_5326);
nor U6832 (N_6832,N_4975,N_4470);
or U6833 (N_6833,N_5545,N_4095);
nor U6834 (N_6834,N_5694,N_4192);
nor U6835 (N_6835,N_4496,N_4238);
and U6836 (N_6836,N_4143,N_4175);
and U6837 (N_6837,N_5917,N_4542);
nor U6838 (N_6838,N_4148,N_4474);
nor U6839 (N_6839,N_4400,N_5560);
xnor U6840 (N_6840,N_5942,N_5165);
or U6841 (N_6841,N_5611,N_4455);
and U6842 (N_6842,N_4901,N_4479);
nand U6843 (N_6843,N_5384,N_5522);
xnor U6844 (N_6844,N_5709,N_5700);
nor U6845 (N_6845,N_4620,N_4100);
and U6846 (N_6846,N_4363,N_5876);
and U6847 (N_6847,N_4636,N_5582);
or U6848 (N_6848,N_5623,N_5277);
nor U6849 (N_6849,N_4703,N_5229);
nand U6850 (N_6850,N_4753,N_5434);
and U6851 (N_6851,N_5148,N_4594);
or U6852 (N_6852,N_5287,N_5889);
nand U6853 (N_6853,N_4716,N_4079);
nor U6854 (N_6854,N_4609,N_4360);
or U6855 (N_6855,N_5908,N_4593);
or U6856 (N_6856,N_5755,N_4637);
nand U6857 (N_6857,N_4569,N_4118);
and U6858 (N_6858,N_4413,N_5526);
nand U6859 (N_6859,N_4908,N_5058);
nand U6860 (N_6860,N_5589,N_4601);
and U6861 (N_6861,N_5436,N_4185);
nand U6862 (N_6862,N_4947,N_4882);
or U6863 (N_6863,N_4705,N_4919);
nand U6864 (N_6864,N_5314,N_4525);
nor U6865 (N_6865,N_5403,N_4893);
or U6866 (N_6866,N_4813,N_5118);
xor U6867 (N_6867,N_5448,N_4698);
xor U6868 (N_6868,N_4123,N_5108);
xnor U6869 (N_6869,N_4869,N_4566);
nor U6870 (N_6870,N_4374,N_4307);
xnor U6871 (N_6871,N_4014,N_5206);
nor U6872 (N_6872,N_4053,N_5797);
or U6873 (N_6873,N_5370,N_4825);
xnor U6874 (N_6874,N_4047,N_5007);
or U6875 (N_6875,N_5949,N_5945);
nor U6876 (N_6876,N_4404,N_5798);
and U6877 (N_6877,N_5003,N_5509);
nor U6878 (N_6878,N_5129,N_5618);
and U6879 (N_6879,N_5512,N_5822);
nand U6880 (N_6880,N_4235,N_5356);
nor U6881 (N_6881,N_5966,N_4624);
or U6882 (N_6882,N_5163,N_5109);
nand U6883 (N_6883,N_4200,N_4979);
xnor U6884 (N_6884,N_4738,N_5311);
nand U6885 (N_6885,N_4632,N_4973);
xor U6886 (N_6886,N_4986,N_5354);
xor U6887 (N_6887,N_4923,N_4557);
nand U6888 (N_6888,N_4782,N_5361);
nor U6889 (N_6889,N_4066,N_5818);
xor U6890 (N_6890,N_4497,N_4163);
xnor U6891 (N_6891,N_4405,N_5549);
xnor U6892 (N_6892,N_5668,N_4870);
and U6893 (N_6893,N_4473,N_5817);
or U6894 (N_6894,N_5458,N_5202);
or U6895 (N_6895,N_4348,N_5590);
or U6896 (N_6896,N_4827,N_4732);
and U6897 (N_6897,N_5721,N_5038);
nor U6898 (N_6898,N_5027,N_4449);
or U6899 (N_6899,N_5216,N_4970);
nor U6900 (N_6900,N_4933,N_4502);
and U6901 (N_6901,N_4340,N_5099);
nor U6902 (N_6902,N_4828,N_5093);
and U6903 (N_6903,N_4556,N_5224);
xor U6904 (N_6904,N_5529,N_4885);
or U6905 (N_6905,N_4018,N_4454);
or U6906 (N_6906,N_5573,N_5460);
nor U6907 (N_6907,N_5861,N_4807);
xnor U6908 (N_6908,N_5461,N_5472);
nor U6909 (N_6909,N_5162,N_5295);
xor U6910 (N_6910,N_5743,N_4222);
nand U6911 (N_6911,N_4905,N_4836);
or U6912 (N_6912,N_5858,N_4038);
nand U6913 (N_6913,N_4706,N_5299);
xnor U6914 (N_6914,N_4127,N_4495);
or U6915 (N_6915,N_4759,N_4373);
or U6916 (N_6916,N_5378,N_5121);
or U6917 (N_6917,N_4281,N_4040);
nor U6918 (N_6918,N_5792,N_4622);
nand U6919 (N_6919,N_4867,N_5499);
and U6920 (N_6920,N_4029,N_5802);
and U6921 (N_6921,N_5328,N_5465);
nor U6922 (N_6922,N_4493,N_4997);
nand U6923 (N_6923,N_4041,N_5923);
or U6924 (N_6924,N_5218,N_5901);
nand U6925 (N_6925,N_4120,N_5971);
or U6926 (N_6926,N_5263,N_4585);
nand U6927 (N_6927,N_5053,N_5187);
or U6928 (N_6928,N_4959,N_5284);
nor U6929 (N_6929,N_4806,N_4945);
and U6930 (N_6930,N_4778,N_5542);
or U6931 (N_6931,N_5935,N_4483);
or U6932 (N_6932,N_5513,N_5940);
and U6933 (N_6933,N_5532,N_5442);
nor U6934 (N_6934,N_4049,N_5815);
nor U6935 (N_6935,N_5408,N_5912);
nand U6936 (N_6936,N_5025,N_5212);
nor U6937 (N_6937,N_4015,N_5622);
or U6938 (N_6938,N_4588,N_5621);
or U6939 (N_6939,N_5302,N_4760);
or U6940 (N_6940,N_5394,N_5032);
and U6941 (N_6941,N_4088,N_4509);
and U6942 (N_6942,N_4512,N_5415);
or U6943 (N_6943,N_5521,N_4731);
xnor U6944 (N_6944,N_4305,N_5580);
nor U6945 (N_6945,N_5088,N_4381);
xnor U6946 (N_6946,N_5091,N_5701);
and U6947 (N_6947,N_4438,N_5567);
or U6948 (N_6948,N_4051,N_5102);
nor U6949 (N_6949,N_4368,N_4221);
nand U6950 (N_6950,N_5646,N_5400);
nor U6951 (N_6951,N_5406,N_5101);
nor U6952 (N_6952,N_5294,N_5052);
xor U6953 (N_6953,N_4819,N_4241);
nand U6954 (N_6954,N_4853,N_5183);
and U6955 (N_6955,N_5177,N_5857);
and U6956 (N_6956,N_5124,N_5850);
nor U6957 (N_6957,N_5516,N_5998);
xor U6958 (N_6958,N_4328,N_4299);
and U6959 (N_6959,N_4131,N_4354);
xor U6960 (N_6960,N_4437,N_4879);
nand U6961 (N_6961,N_4817,N_4544);
nor U6962 (N_6962,N_4524,N_4198);
xnor U6963 (N_6963,N_5874,N_5671);
nand U6964 (N_6964,N_5997,N_4452);
nor U6965 (N_6965,N_5788,N_4693);
nor U6966 (N_6966,N_4253,N_4978);
and U6967 (N_6967,N_4625,N_5789);
nand U6968 (N_6968,N_5866,N_5473);
or U6969 (N_6969,N_5359,N_5927);
and U6970 (N_6970,N_4775,N_4793);
nand U6971 (N_6971,N_4591,N_4498);
nor U6972 (N_6972,N_4166,N_4526);
nand U6973 (N_6973,N_4165,N_5976);
nand U6974 (N_6974,N_4662,N_4332);
or U6975 (N_6975,N_4064,N_4135);
nand U6976 (N_6976,N_4603,N_4918);
nand U6977 (N_6977,N_4831,N_4786);
xor U6978 (N_6978,N_4427,N_4154);
nor U6979 (N_6979,N_5661,N_4178);
and U6980 (N_6980,N_4364,N_5551);
and U6981 (N_6981,N_4346,N_4809);
nand U6982 (N_6982,N_4220,N_5724);
xor U6983 (N_6983,N_5334,N_5615);
nor U6984 (N_6984,N_4796,N_4562);
xor U6985 (N_6985,N_5972,N_4464);
and U6986 (N_6986,N_5564,N_5203);
nor U6987 (N_6987,N_5401,N_4117);
and U6988 (N_6988,N_4640,N_4461);
nor U6989 (N_6989,N_5039,N_5290);
nand U6990 (N_6990,N_4790,N_5878);
nand U6991 (N_6991,N_5383,N_4071);
nand U6992 (N_6992,N_4210,N_4068);
and U6993 (N_6993,N_4080,N_4243);
nand U6994 (N_6994,N_4611,N_5267);
nand U6995 (N_6995,N_4418,N_5678);
nand U6996 (N_6996,N_5744,N_5286);
or U6997 (N_6997,N_5482,N_4288);
nor U6998 (N_6998,N_4681,N_4478);
nand U6999 (N_6999,N_5739,N_5810);
and U7000 (N_7000,N_4076,N_5375);
xnor U7001 (N_7001,N_5038,N_5719);
xor U7002 (N_7002,N_4646,N_4166);
or U7003 (N_7003,N_5485,N_4169);
or U7004 (N_7004,N_4033,N_4637);
or U7005 (N_7005,N_5713,N_5672);
nand U7006 (N_7006,N_4184,N_4491);
and U7007 (N_7007,N_4049,N_5175);
nand U7008 (N_7008,N_4815,N_5325);
nor U7009 (N_7009,N_5679,N_4738);
or U7010 (N_7010,N_4880,N_5206);
xor U7011 (N_7011,N_4573,N_4473);
nand U7012 (N_7012,N_4944,N_5192);
or U7013 (N_7013,N_4983,N_5930);
and U7014 (N_7014,N_5687,N_5931);
nor U7015 (N_7015,N_4892,N_4713);
and U7016 (N_7016,N_5393,N_5816);
nand U7017 (N_7017,N_5390,N_4183);
and U7018 (N_7018,N_5581,N_4592);
nor U7019 (N_7019,N_5874,N_4416);
and U7020 (N_7020,N_5367,N_5248);
nand U7021 (N_7021,N_5052,N_5189);
and U7022 (N_7022,N_5172,N_4435);
or U7023 (N_7023,N_5129,N_4525);
xor U7024 (N_7024,N_5299,N_4579);
and U7025 (N_7025,N_4905,N_5137);
or U7026 (N_7026,N_5215,N_5090);
or U7027 (N_7027,N_4517,N_5504);
nor U7028 (N_7028,N_4215,N_4835);
nor U7029 (N_7029,N_4001,N_5894);
and U7030 (N_7030,N_4340,N_4749);
and U7031 (N_7031,N_4187,N_5518);
xnor U7032 (N_7032,N_4998,N_5941);
nand U7033 (N_7033,N_4555,N_4032);
and U7034 (N_7034,N_4140,N_5214);
nor U7035 (N_7035,N_4244,N_4206);
or U7036 (N_7036,N_4527,N_5330);
nand U7037 (N_7037,N_5529,N_5448);
nand U7038 (N_7038,N_5957,N_4817);
or U7039 (N_7039,N_4880,N_4034);
and U7040 (N_7040,N_4479,N_5071);
or U7041 (N_7041,N_4429,N_5971);
nor U7042 (N_7042,N_4270,N_5303);
and U7043 (N_7043,N_4732,N_4666);
or U7044 (N_7044,N_4328,N_5600);
nor U7045 (N_7045,N_4028,N_5680);
nor U7046 (N_7046,N_5187,N_5972);
nand U7047 (N_7047,N_5241,N_4414);
nand U7048 (N_7048,N_4699,N_4881);
nor U7049 (N_7049,N_4428,N_4508);
nand U7050 (N_7050,N_4798,N_4622);
nor U7051 (N_7051,N_5297,N_5624);
and U7052 (N_7052,N_5233,N_5979);
xnor U7053 (N_7053,N_4618,N_5327);
and U7054 (N_7054,N_4233,N_5921);
or U7055 (N_7055,N_5694,N_5945);
nand U7056 (N_7056,N_4733,N_5031);
nand U7057 (N_7057,N_5919,N_4860);
and U7058 (N_7058,N_4534,N_5831);
xnor U7059 (N_7059,N_4224,N_4760);
nor U7060 (N_7060,N_5487,N_4388);
nor U7061 (N_7061,N_4651,N_4118);
xnor U7062 (N_7062,N_5003,N_4724);
and U7063 (N_7063,N_5073,N_5288);
nor U7064 (N_7064,N_4627,N_5549);
nand U7065 (N_7065,N_4035,N_5917);
and U7066 (N_7066,N_4469,N_5824);
nand U7067 (N_7067,N_5654,N_5797);
xor U7068 (N_7068,N_4482,N_4439);
or U7069 (N_7069,N_4568,N_4708);
nor U7070 (N_7070,N_4715,N_4987);
nor U7071 (N_7071,N_4095,N_5000);
or U7072 (N_7072,N_5950,N_5891);
nor U7073 (N_7073,N_4977,N_4828);
nor U7074 (N_7074,N_4546,N_5753);
xnor U7075 (N_7075,N_5998,N_5652);
or U7076 (N_7076,N_5847,N_5627);
nor U7077 (N_7077,N_4394,N_4836);
nor U7078 (N_7078,N_4033,N_5673);
nand U7079 (N_7079,N_4506,N_5734);
nand U7080 (N_7080,N_5448,N_4726);
xnor U7081 (N_7081,N_5004,N_5596);
nand U7082 (N_7082,N_4077,N_4233);
and U7083 (N_7083,N_5365,N_5991);
xor U7084 (N_7084,N_4931,N_4208);
nand U7085 (N_7085,N_5188,N_5331);
nand U7086 (N_7086,N_5546,N_4625);
nor U7087 (N_7087,N_4550,N_4224);
and U7088 (N_7088,N_5646,N_5067);
and U7089 (N_7089,N_5256,N_4761);
nand U7090 (N_7090,N_4575,N_5535);
nor U7091 (N_7091,N_5363,N_5242);
nand U7092 (N_7092,N_5849,N_4374);
and U7093 (N_7093,N_4483,N_5786);
or U7094 (N_7094,N_5285,N_4239);
nor U7095 (N_7095,N_5309,N_4728);
xnor U7096 (N_7096,N_5216,N_5351);
and U7097 (N_7097,N_4818,N_4292);
and U7098 (N_7098,N_5866,N_4707);
nand U7099 (N_7099,N_4666,N_5861);
nor U7100 (N_7100,N_4237,N_4212);
or U7101 (N_7101,N_4373,N_5933);
and U7102 (N_7102,N_5294,N_5878);
nand U7103 (N_7103,N_4325,N_5360);
and U7104 (N_7104,N_4200,N_4733);
nor U7105 (N_7105,N_4327,N_5224);
or U7106 (N_7106,N_4387,N_5714);
nor U7107 (N_7107,N_4786,N_4031);
nand U7108 (N_7108,N_4242,N_5287);
nand U7109 (N_7109,N_5079,N_4410);
or U7110 (N_7110,N_4341,N_4395);
nor U7111 (N_7111,N_5202,N_4856);
or U7112 (N_7112,N_4242,N_4832);
or U7113 (N_7113,N_5967,N_5796);
nand U7114 (N_7114,N_4782,N_4558);
or U7115 (N_7115,N_5237,N_4380);
or U7116 (N_7116,N_4061,N_4381);
nor U7117 (N_7117,N_5537,N_5044);
xor U7118 (N_7118,N_5730,N_4901);
nand U7119 (N_7119,N_4443,N_5750);
nor U7120 (N_7120,N_5200,N_5528);
nand U7121 (N_7121,N_4807,N_4490);
nand U7122 (N_7122,N_4443,N_5610);
xnor U7123 (N_7123,N_5991,N_5745);
nor U7124 (N_7124,N_4805,N_4409);
or U7125 (N_7125,N_5185,N_5693);
xor U7126 (N_7126,N_5324,N_5853);
nor U7127 (N_7127,N_4779,N_4078);
nand U7128 (N_7128,N_4870,N_4540);
nor U7129 (N_7129,N_5560,N_5319);
or U7130 (N_7130,N_4708,N_5519);
or U7131 (N_7131,N_4258,N_5893);
xnor U7132 (N_7132,N_5394,N_4997);
nand U7133 (N_7133,N_5522,N_4751);
nor U7134 (N_7134,N_4647,N_4616);
or U7135 (N_7135,N_5416,N_4438);
xnor U7136 (N_7136,N_4124,N_4511);
and U7137 (N_7137,N_4249,N_5121);
xor U7138 (N_7138,N_5094,N_5737);
xnor U7139 (N_7139,N_5449,N_4276);
xor U7140 (N_7140,N_5876,N_4633);
or U7141 (N_7141,N_4919,N_4760);
xnor U7142 (N_7142,N_5665,N_5661);
and U7143 (N_7143,N_4980,N_4264);
nor U7144 (N_7144,N_5635,N_5787);
nand U7145 (N_7145,N_4460,N_5253);
nand U7146 (N_7146,N_5935,N_5528);
nor U7147 (N_7147,N_4580,N_4582);
nor U7148 (N_7148,N_5234,N_5862);
xnor U7149 (N_7149,N_5734,N_5430);
nor U7150 (N_7150,N_4834,N_4290);
or U7151 (N_7151,N_4456,N_5449);
xnor U7152 (N_7152,N_5090,N_5576);
nor U7153 (N_7153,N_5697,N_4330);
nand U7154 (N_7154,N_5089,N_5032);
and U7155 (N_7155,N_5932,N_4727);
and U7156 (N_7156,N_5400,N_5337);
and U7157 (N_7157,N_4913,N_4275);
or U7158 (N_7158,N_4184,N_5455);
nand U7159 (N_7159,N_4723,N_4007);
or U7160 (N_7160,N_5644,N_4999);
and U7161 (N_7161,N_5124,N_5213);
or U7162 (N_7162,N_5930,N_4476);
nor U7163 (N_7163,N_5928,N_5183);
or U7164 (N_7164,N_4452,N_5282);
nand U7165 (N_7165,N_5231,N_4885);
and U7166 (N_7166,N_5808,N_4777);
and U7167 (N_7167,N_5798,N_5366);
xnor U7168 (N_7168,N_5551,N_5962);
nand U7169 (N_7169,N_4812,N_5514);
nand U7170 (N_7170,N_5824,N_4497);
xnor U7171 (N_7171,N_5959,N_5803);
and U7172 (N_7172,N_4556,N_4778);
nor U7173 (N_7173,N_4272,N_4971);
nor U7174 (N_7174,N_5622,N_5261);
or U7175 (N_7175,N_4961,N_4028);
or U7176 (N_7176,N_4657,N_4599);
and U7177 (N_7177,N_4743,N_4927);
nand U7178 (N_7178,N_4097,N_4721);
or U7179 (N_7179,N_5733,N_5410);
nand U7180 (N_7180,N_4174,N_4249);
or U7181 (N_7181,N_4236,N_4676);
and U7182 (N_7182,N_5888,N_5648);
or U7183 (N_7183,N_4581,N_4311);
and U7184 (N_7184,N_4299,N_5617);
or U7185 (N_7185,N_4209,N_4660);
nand U7186 (N_7186,N_4350,N_4151);
nor U7187 (N_7187,N_5396,N_5607);
nand U7188 (N_7188,N_4772,N_4296);
and U7189 (N_7189,N_5968,N_5008);
xnor U7190 (N_7190,N_5396,N_4300);
nor U7191 (N_7191,N_5196,N_5122);
xor U7192 (N_7192,N_5639,N_4980);
xor U7193 (N_7193,N_4178,N_4417);
nor U7194 (N_7194,N_4614,N_5180);
and U7195 (N_7195,N_5056,N_4111);
and U7196 (N_7196,N_4151,N_5996);
and U7197 (N_7197,N_4729,N_5728);
xnor U7198 (N_7198,N_5235,N_5383);
nand U7199 (N_7199,N_5553,N_5356);
nor U7200 (N_7200,N_5890,N_4562);
nand U7201 (N_7201,N_5794,N_4839);
nor U7202 (N_7202,N_4525,N_4667);
nor U7203 (N_7203,N_5334,N_4861);
xor U7204 (N_7204,N_4601,N_5594);
xor U7205 (N_7205,N_5830,N_4547);
nor U7206 (N_7206,N_4342,N_5586);
nand U7207 (N_7207,N_4135,N_5657);
or U7208 (N_7208,N_4002,N_4182);
xor U7209 (N_7209,N_4795,N_4995);
xor U7210 (N_7210,N_5596,N_5948);
or U7211 (N_7211,N_4452,N_5075);
xor U7212 (N_7212,N_5863,N_5689);
or U7213 (N_7213,N_4538,N_5992);
and U7214 (N_7214,N_4555,N_4680);
nand U7215 (N_7215,N_4063,N_5941);
nor U7216 (N_7216,N_4474,N_5806);
and U7217 (N_7217,N_4150,N_5987);
xnor U7218 (N_7218,N_5020,N_5669);
nand U7219 (N_7219,N_5477,N_5454);
xnor U7220 (N_7220,N_4550,N_4811);
nand U7221 (N_7221,N_5175,N_5688);
nand U7222 (N_7222,N_4960,N_4426);
or U7223 (N_7223,N_4868,N_4105);
or U7224 (N_7224,N_5115,N_4069);
or U7225 (N_7225,N_5168,N_5375);
xnor U7226 (N_7226,N_4185,N_4681);
xnor U7227 (N_7227,N_4955,N_4315);
nor U7228 (N_7228,N_5394,N_4561);
or U7229 (N_7229,N_4937,N_4712);
or U7230 (N_7230,N_4281,N_4450);
xor U7231 (N_7231,N_4802,N_5371);
or U7232 (N_7232,N_4363,N_4103);
xnor U7233 (N_7233,N_4991,N_4917);
nor U7234 (N_7234,N_4994,N_5436);
nand U7235 (N_7235,N_4302,N_4088);
xnor U7236 (N_7236,N_4962,N_5949);
or U7237 (N_7237,N_5553,N_4446);
or U7238 (N_7238,N_4489,N_5967);
or U7239 (N_7239,N_4534,N_4715);
nor U7240 (N_7240,N_4231,N_5414);
and U7241 (N_7241,N_4665,N_5255);
and U7242 (N_7242,N_4103,N_5370);
nand U7243 (N_7243,N_4537,N_5984);
nor U7244 (N_7244,N_4948,N_5038);
nor U7245 (N_7245,N_4820,N_5928);
nand U7246 (N_7246,N_5308,N_4782);
or U7247 (N_7247,N_5550,N_4966);
or U7248 (N_7248,N_4980,N_4163);
nor U7249 (N_7249,N_5693,N_4361);
nor U7250 (N_7250,N_4879,N_4395);
and U7251 (N_7251,N_5899,N_5173);
or U7252 (N_7252,N_4439,N_5714);
nor U7253 (N_7253,N_4223,N_5860);
and U7254 (N_7254,N_4795,N_4628);
and U7255 (N_7255,N_4532,N_5907);
nand U7256 (N_7256,N_4464,N_4861);
and U7257 (N_7257,N_5000,N_5187);
nor U7258 (N_7258,N_4552,N_4062);
nor U7259 (N_7259,N_5125,N_5628);
nor U7260 (N_7260,N_4130,N_4601);
nand U7261 (N_7261,N_5694,N_4897);
nand U7262 (N_7262,N_4330,N_5208);
or U7263 (N_7263,N_5709,N_4017);
nor U7264 (N_7264,N_4603,N_5598);
nand U7265 (N_7265,N_5847,N_4411);
nand U7266 (N_7266,N_4144,N_4383);
or U7267 (N_7267,N_4189,N_5811);
nand U7268 (N_7268,N_4592,N_5785);
or U7269 (N_7269,N_5701,N_5356);
xor U7270 (N_7270,N_5528,N_4597);
and U7271 (N_7271,N_5611,N_5659);
nand U7272 (N_7272,N_5391,N_4393);
xnor U7273 (N_7273,N_4759,N_5035);
xor U7274 (N_7274,N_4889,N_5892);
xor U7275 (N_7275,N_4304,N_5351);
or U7276 (N_7276,N_4028,N_4693);
nand U7277 (N_7277,N_4264,N_5946);
and U7278 (N_7278,N_4852,N_4203);
nor U7279 (N_7279,N_5079,N_5833);
nor U7280 (N_7280,N_5332,N_4285);
xor U7281 (N_7281,N_4341,N_4667);
xor U7282 (N_7282,N_5862,N_4707);
and U7283 (N_7283,N_5506,N_5632);
xor U7284 (N_7284,N_4323,N_5098);
and U7285 (N_7285,N_5973,N_5877);
or U7286 (N_7286,N_4280,N_5099);
xnor U7287 (N_7287,N_5828,N_4930);
and U7288 (N_7288,N_5030,N_4694);
or U7289 (N_7289,N_5052,N_4132);
nand U7290 (N_7290,N_5406,N_5608);
nor U7291 (N_7291,N_4530,N_5525);
nand U7292 (N_7292,N_4138,N_4510);
nor U7293 (N_7293,N_5204,N_4504);
xor U7294 (N_7294,N_4212,N_5596);
or U7295 (N_7295,N_4299,N_4753);
xnor U7296 (N_7296,N_4580,N_5702);
xnor U7297 (N_7297,N_5151,N_4555);
or U7298 (N_7298,N_4780,N_4982);
nor U7299 (N_7299,N_4554,N_5964);
and U7300 (N_7300,N_5839,N_5574);
nand U7301 (N_7301,N_4961,N_5950);
or U7302 (N_7302,N_4816,N_5882);
xor U7303 (N_7303,N_4613,N_4006);
nand U7304 (N_7304,N_5143,N_4328);
xor U7305 (N_7305,N_4677,N_5194);
and U7306 (N_7306,N_5822,N_5370);
and U7307 (N_7307,N_4056,N_4343);
or U7308 (N_7308,N_5050,N_5590);
xnor U7309 (N_7309,N_4014,N_4480);
xnor U7310 (N_7310,N_4697,N_5662);
or U7311 (N_7311,N_4214,N_4222);
nor U7312 (N_7312,N_4004,N_4378);
xor U7313 (N_7313,N_4193,N_5495);
nor U7314 (N_7314,N_4868,N_4184);
or U7315 (N_7315,N_4233,N_4468);
xor U7316 (N_7316,N_5153,N_5238);
and U7317 (N_7317,N_4559,N_4778);
nand U7318 (N_7318,N_4513,N_4160);
or U7319 (N_7319,N_5890,N_5664);
or U7320 (N_7320,N_4105,N_4635);
nand U7321 (N_7321,N_4044,N_5872);
xor U7322 (N_7322,N_5152,N_4175);
or U7323 (N_7323,N_4286,N_5678);
xnor U7324 (N_7324,N_5459,N_4350);
or U7325 (N_7325,N_4090,N_4478);
xnor U7326 (N_7326,N_5166,N_4458);
nor U7327 (N_7327,N_4943,N_4562);
nand U7328 (N_7328,N_5544,N_5649);
xnor U7329 (N_7329,N_4016,N_5755);
and U7330 (N_7330,N_5709,N_4428);
and U7331 (N_7331,N_5104,N_5395);
nand U7332 (N_7332,N_5208,N_4129);
nor U7333 (N_7333,N_5275,N_4931);
nand U7334 (N_7334,N_4815,N_5548);
or U7335 (N_7335,N_5612,N_5500);
or U7336 (N_7336,N_5942,N_5768);
and U7337 (N_7337,N_4262,N_4109);
or U7338 (N_7338,N_4284,N_5223);
and U7339 (N_7339,N_4904,N_5904);
or U7340 (N_7340,N_4197,N_5642);
or U7341 (N_7341,N_4795,N_4015);
and U7342 (N_7342,N_4397,N_4662);
or U7343 (N_7343,N_4086,N_5953);
xor U7344 (N_7344,N_5672,N_4331);
nand U7345 (N_7345,N_4656,N_5112);
nand U7346 (N_7346,N_4077,N_4740);
or U7347 (N_7347,N_5719,N_4152);
and U7348 (N_7348,N_4831,N_4273);
or U7349 (N_7349,N_5913,N_4596);
and U7350 (N_7350,N_4540,N_5063);
or U7351 (N_7351,N_4850,N_5855);
nor U7352 (N_7352,N_4840,N_4167);
nand U7353 (N_7353,N_4128,N_4480);
or U7354 (N_7354,N_4809,N_5188);
and U7355 (N_7355,N_5648,N_5750);
xnor U7356 (N_7356,N_5664,N_5285);
and U7357 (N_7357,N_4998,N_5239);
nor U7358 (N_7358,N_4012,N_5548);
xor U7359 (N_7359,N_5601,N_5285);
nor U7360 (N_7360,N_5069,N_4924);
xor U7361 (N_7361,N_4988,N_5689);
and U7362 (N_7362,N_4546,N_4739);
nor U7363 (N_7363,N_5526,N_4510);
and U7364 (N_7364,N_5123,N_4145);
and U7365 (N_7365,N_5656,N_4443);
and U7366 (N_7366,N_4214,N_5411);
or U7367 (N_7367,N_5252,N_4181);
nand U7368 (N_7368,N_5807,N_5883);
and U7369 (N_7369,N_5931,N_5911);
nand U7370 (N_7370,N_5520,N_5587);
and U7371 (N_7371,N_4210,N_4027);
xor U7372 (N_7372,N_5704,N_5283);
or U7373 (N_7373,N_4877,N_4553);
xnor U7374 (N_7374,N_5913,N_5927);
and U7375 (N_7375,N_5332,N_4297);
and U7376 (N_7376,N_5562,N_4181);
nor U7377 (N_7377,N_5095,N_5629);
nor U7378 (N_7378,N_4694,N_5608);
nor U7379 (N_7379,N_4829,N_4758);
nand U7380 (N_7380,N_4457,N_5668);
xnor U7381 (N_7381,N_4804,N_4613);
and U7382 (N_7382,N_4207,N_4148);
or U7383 (N_7383,N_4284,N_5142);
xnor U7384 (N_7384,N_5592,N_4327);
nor U7385 (N_7385,N_5915,N_4992);
xor U7386 (N_7386,N_5415,N_4131);
and U7387 (N_7387,N_4587,N_5747);
and U7388 (N_7388,N_4021,N_4266);
nor U7389 (N_7389,N_4304,N_4520);
nor U7390 (N_7390,N_4271,N_4526);
and U7391 (N_7391,N_5397,N_5376);
nor U7392 (N_7392,N_4729,N_5380);
xor U7393 (N_7393,N_4127,N_4039);
nor U7394 (N_7394,N_4876,N_5476);
nand U7395 (N_7395,N_5806,N_5935);
nand U7396 (N_7396,N_5220,N_4885);
xor U7397 (N_7397,N_4135,N_4060);
and U7398 (N_7398,N_5019,N_5399);
and U7399 (N_7399,N_4825,N_4813);
or U7400 (N_7400,N_4027,N_5568);
or U7401 (N_7401,N_5429,N_5337);
nor U7402 (N_7402,N_5447,N_5582);
or U7403 (N_7403,N_4585,N_5923);
nor U7404 (N_7404,N_4654,N_4658);
or U7405 (N_7405,N_5368,N_4533);
and U7406 (N_7406,N_5396,N_5334);
or U7407 (N_7407,N_4218,N_5264);
xor U7408 (N_7408,N_4208,N_5659);
and U7409 (N_7409,N_5286,N_5812);
and U7410 (N_7410,N_4882,N_4215);
and U7411 (N_7411,N_4497,N_4367);
xnor U7412 (N_7412,N_5946,N_5238);
or U7413 (N_7413,N_4849,N_4235);
or U7414 (N_7414,N_4551,N_4068);
and U7415 (N_7415,N_4840,N_5333);
or U7416 (N_7416,N_4554,N_5240);
nand U7417 (N_7417,N_5313,N_5761);
nand U7418 (N_7418,N_4687,N_5486);
nand U7419 (N_7419,N_5609,N_5799);
xnor U7420 (N_7420,N_4726,N_5932);
xor U7421 (N_7421,N_5993,N_4533);
or U7422 (N_7422,N_5895,N_4360);
nor U7423 (N_7423,N_5121,N_5004);
and U7424 (N_7424,N_4674,N_4748);
and U7425 (N_7425,N_4248,N_4380);
or U7426 (N_7426,N_4205,N_4349);
xnor U7427 (N_7427,N_5697,N_4660);
xor U7428 (N_7428,N_5722,N_5200);
nand U7429 (N_7429,N_5685,N_4449);
nor U7430 (N_7430,N_5506,N_5921);
and U7431 (N_7431,N_5563,N_5963);
nor U7432 (N_7432,N_5519,N_5413);
nor U7433 (N_7433,N_4748,N_4495);
nand U7434 (N_7434,N_5262,N_5187);
nand U7435 (N_7435,N_5609,N_4696);
nand U7436 (N_7436,N_4800,N_4249);
and U7437 (N_7437,N_4612,N_5232);
and U7438 (N_7438,N_4074,N_5851);
nand U7439 (N_7439,N_4907,N_4849);
or U7440 (N_7440,N_5688,N_4319);
xor U7441 (N_7441,N_5155,N_4246);
xor U7442 (N_7442,N_4431,N_4288);
nand U7443 (N_7443,N_5202,N_5536);
xor U7444 (N_7444,N_4982,N_5907);
xor U7445 (N_7445,N_5219,N_4402);
xnor U7446 (N_7446,N_4783,N_4808);
nand U7447 (N_7447,N_4053,N_5779);
xor U7448 (N_7448,N_5991,N_5784);
and U7449 (N_7449,N_5928,N_4853);
nor U7450 (N_7450,N_4548,N_5340);
or U7451 (N_7451,N_4896,N_5146);
xor U7452 (N_7452,N_4228,N_4892);
xnor U7453 (N_7453,N_5616,N_5909);
xor U7454 (N_7454,N_4521,N_5193);
nand U7455 (N_7455,N_4727,N_4200);
nand U7456 (N_7456,N_5794,N_5342);
or U7457 (N_7457,N_5421,N_5481);
and U7458 (N_7458,N_4608,N_4429);
and U7459 (N_7459,N_5421,N_5633);
nor U7460 (N_7460,N_4324,N_5984);
nor U7461 (N_7461,N_4346,N_4887);
nor U7462 (N_7462,N_4058,N_4533);
or U7463 (N_7463,N_4478,N_4723);
or U7464 (N_7464,N_4610,N_4083);
nor U7465 (N_7465,N_4228,N_5367);
xnor U7466 (N_7466,N_5448,N_4536);
or U7467 (N_7467,N_5800,N_4112);
nor U7468 (N_7468,N_4816,N_4122);
or U7469 (N_7469,N_4656,N_4984);
nand U7470 (N_7470,N_4687,N_5039);
and U7471 (N_7471,N_4413,N_5256);
and U7472 (N_7472,N_4848,N_5268);
nand U7473 (N_7473,N_5199,N_5647);
nand U7474 (N_7474,N_4973,N_4065);
and U7475 (N_7475,N_5318,N_4380);
nand U7476 (N_7476,N_5860,N_4016);
and U7477 (N_7477,N_5630,N_4893);
or U7478 (N_7478,N_4540,N_4303);
and U7479 (N_7479,N_5208,N_5134);
nand U7480 (N_7480,N_4441,N_4026);
xor U7481 (N_7481,N_5036,N_5446);
nor U7482 (N_7482,N_5092,N_5483);
or U7483 (N_7483,N_4147,N_5460);
or U7484 (N_7484,N_4741,N_5080);
xnor U7485 (N_7485,N_4265,N_4999);
or U7486 (N_7486,N_4854,N_4051);
and U7487 (N_7487,N_5873,N_5332);
nand U7488 (N_7488,N_4474,N_4649);
nor U7489 (N_7489,N_4371,N_4193);
or U7490 (N_7490,N_5868,N_5548);
nor U7491 (N_7491,N_4380,N_4395);
xor U7492 (N_7492,N_4192,N_4328);
and U7493 (N_7493,N_5284,N_4245);
or U7494 (N_7494,N_4546,N_5822);
or U7495 (N_7495,N_4291,N_5272);
nor U7496 (N_7496,N_5122,N_4151);
nor U7497 (N_7497,N_4194,N_5998);
nand U7498 (N_7498,N_5290,N_4107);
nand U7499 (N_7499,N_4615,N_5794);
nand U7500 (N_7500,N_4161,N_4872);
or U7501 (N_7501,N_4020,N_5325);
and U7502 (N_7502,N_5018,N_4608);
nor U7503 (N_7503,N_4627,N_4149);
nor U7504 (N_7504,N_4335,N_5117);
xnor U7505 (N_7505,N_5872,N_5666);
nor U7506 (N_7506,N_5103,N_4090);
nor U7507 (N_7507,N_5629,N_4940);
and U7508 (N_7508,N_4630,N_5891);
nand U7509 (N_7509,N_4960,N_5292);
and U7510 (N_7510,N_5443,N_4894);
or U7511 (N_7511,N_5349,N_5603);
nor U7512 (N_7512,N_5580,N_4280);
nor U7513 (N_7513,N_5870,N_5202);
and U7514 (N_7514,N_5093,N_5824);
or U7515 (N_7515,N_5194,N_5168);
xnor U7516 (N_7516,N_5379,N_4840);
and U7517 (N_7517,N_5865,N_5753);
or U7518 (N_7518,N_5101,N_5401);
xnor U7519 (N_7519,N_4366,N_4895);
nand U7520 (N_7520,N_5483,N_4704);
nor U7521 (N_7521,N_4565,N_4142);
nand U7522 (N_7522,N_5499,N_4675);
or U7523 (N_7523,N_4566,N_5639);
and U7524 (N_7524,N_4757,N_4018);
or U7525 (N_7525,N_5061,N_5411);
nand U7526 (N_7526,N_4336,N_5895);
or U7527 (N_7527,N_5797,N_4004);
nor U7528 (N_7528,N_5849,N_5628);
xor U7529 (N_7529,N_5998,N_4813);
nand U7530 (N_7530,N_4227,N_5505);
nor U7531 (N_7531,N_4485,N_4882);
nand U7532 (N_7532,N_4737,N_5285);
and U7533 (N_7533,N_4390,N_4707);
nand U7534 (N_7534,N_4151,N_4533);
nand U7535 (N_7535,N_4452,N_5756);
nand U7536 (N_7536,N_4806,N_4916);
xor U7537 (N_7537,N_4935,N_5401);
nor U7538 (N_7538,N_5999,N_4458);
nor U7539 (N_7539,N_5074,N_5507);
or U7540 (N_7540,N_5976,N_4758);
and U7541 (N_7541,N_4919,N_4302);
or U7542 (N_7542,N_5491,N_5273);
xor U7543 (N_7543,N_5455,N_5988);
nor U7544 (N_7544,N_5828,N_5788);
or U7545 (N_7545,N_5024,N_5899);
and U7546 (N_7546,N_5580,N_5369);
or U7547 (N_7547,N_4947,N_4865);
nand U7548 (N_7548,N_4460,N_4671);
and U7549 (N_7549,N_5070,N_4274);
nor U7550 (N_7550,N_4724,N_5536);
xnor U7551 (N_7551,N_5904,N_4186);
nand U7552 (N_7552,N_5010,N_5804);
or U7553 (N_7553,N_4942,N_5336);
xnor U7554 (N_7554,N_4992,N_4664);
or U7555 (N_7555,N_5975,N_4064);
and U7556 (N_7556,N_5589,N_5186);
nand U7557 (N_7557,N_4521,N_5062);
or U7558 (N_7558,N_4693,N_5201);
nor U7559 (N_7559,N_5556,N_5347);
nand U7560 (N_7560,N_4968,N_4448);
xor U7561 (N_7561,N_5527,N_4765);
nand U7562 (N_7562,N_5263,N_5411);
xnor U7563 (N_7563,N_4672,N_5260);
or U7564 (N_7564,N_5808,N_5152);
and U7565 (N_7565,N_4717,N_4774);
xor U7566 (N_7566,N_4950,N_5838);
xnor U7567 (N_7567,N_5028,N_4532);
and U7568 (N_7568,N_5721,N_4006);
nor U7569 (N_7569,N_5404,N_5167);
and U7570 (N_7570,N_5979,N_5749);
and U7571 (N_7571,N_4434,N_5330);
and U7572 (N_7572,N_4225,N_4136);
nor U7573 (N_7573,N_4368,N_4241);
nor U7574 (N_7574,N_5062,N_5630);
nand U7575 (N_7575,N_4781,N_5429);
nand U7576 (N_7576,N_5797,N_4244);
xnor U7577 (N_7577,N_4158,N_4574);
xor U7578 (N_7578,N_5583,N_4268);
and U7579 (N_7579,N_4454,N_4317);
and U7580 (N_7580,N_5720,N_4777);
or U7581 (N_7581,N_5964,N_4924);
or U7582 (N_7582,N_4346,N_5115);
xor U7583 (N_7583,N_4163,N_4075);
nor U7584 (N_7584,N_4101,N_4577);
or U7585 (N_7585,N_5890,N_4269);
or U7586 (N_7586,N_4867,N_4085);
and U7587 (N_7587,N_5684,N_4620);
and U7588 (N_7588,N_4502,N_4797);
xor U7589 (N_7589,N_5900,N_5042);
nor U7590 (N_7590,N_5598,N_4415);
nand U7591 (N_7591,N_5130,N_4231);
xnor U7592 (N_7592,N_5969,N_5092);
or U7593 (N_7593,N_5776,N_5980);
xnor U7594 (N_7594,N_4362,N_4253);
or U7595 (N_7595,N_5712,N_5915);
nand U7596 (N_7596,N_5990,N_4673);
nand U7597 (N_7597,N_5632,N_5477);
nor U7598 (N_7598,N_4848,N_4043);
xnor U7599 (N_7599,N_5456,N_5864);
and U7600 (N_7600,N_5536,N_4296);
and U7601 (N_7601,N_4847,N_5689);
xor U7602 (N_7602,N_4871,N_4806);
nor U7603 (N_7603,N_4379,N_5342);
nor U7604 (N_7604,N_5797,N_5984);
xnor U7605 (N_7605,N_5369,N_4971);
and U7606 (N_7606,N_4578,N_4293);
and U7607 (N_7607,N_5163,N_5078);
and U7608 (N_7608,N_4066,N_4242);
or U7609 (N_7609,N_5428,N_5383);
or U7610 (N_7610,N_4912,N_5726);
nor U7611 (N_7611,N_4940,N_4770);
nor U7612 (N_7612,N_4356,N_4787);
or U7613 (N_7613,N_5401,N_4985);
xnor U7614 (N_7614,N_5087,N_4621);
or U7615 (N_7615,N_5939,N_5832);
nor U7616 (N_7616,N_5618,N_5422);
nor U7617 (N_7617,N_4647,N_5254);
nor U7618 (N_7618,N_4914,N_4461);
and U7619 (N_7619,N_4637,N_5357);
nor U7620 (N_7620,N_4293,N_5003);
or U7621 (N_7621,N_5209,N_5203);
nor U7622 (N_7622,N_4552,N_5267);
and U7623 (N_7623,N_5339,N_4917);
nor U7624 (N_7624,N_5278,N_4395);
or U7625 (N_7625,N_4390,N_4341);
nand U7626 (N_7626,N_5403,N_4646);
and U7627 (N_7627,N_4339,N_4859);
and U7628 (N_7628,N_5184,N_5189);
nor U7629 (N_7629,N_4120,N_4167);
and U7630 (N_7630,N_5696,N_5753);
xnor U7631 (N_7631,N_5784,N_5833);
and U7632 (N_7632,N_4304,N_5139);
or U7633 (N_7633,N_4909,N_5885);
nor U7634 (N_7634,N_5124,N_4276);
nand U7635 (N_7635,N_4526,N_4917);
nand U7636 (N_7636,N_5631,N_4855);
and U7637 (N_7637,N_5151,N_5324);
and U7638 (N_7638,N_5546,N_5842);
and U7639 (N_7639,N_4564,N_5515);
xnor U7640 (N_7640,N_5578,N_5559);
and U7641 (N_7641,N_4497,N_4898);
and U7642 (N_7642,N_4048,N_4280);
nor U7643 (N_7643,N_4708,N_5837);
xnor U7644 (N_7644,N_4792,N_4404);
or U7645 (N_7645,N_5175,N_4988);
or U7646 (N_7646,N_4840,N_4617);
xor U7647 (N_7647,N_4027,N_4250);
nor U7648 (N_7648,N_4951,N_5136);
xnor U7649 (N_7649,N_5874,N_4893);
nor U7650 (N_7650,N_4579,N_4256);
and U7651 (N_7651,N_5918,N_5760);
xnor U7652 (N_7652,N_4693,N_5466);
nor U7653 (N_7653,N_5148,N_5428);
nor U7654 (N_7654,N_5900,N_5815);
and U7655 (N_7655,N_4785,N_5423);
or U7656 (N_7656,N_5436,N_5412);
and U7657 (N_7657,N_4019,N_4901);
and U7658 (N_7658,N_5301,N_5248);
nand U7659 (N_7659,N_5094,N_4100);
and U7660 (N_7660,N_5412,N_5405);
or U7661 (N_7661,N_4823,N_5221);
xnor U7662 (N_7662,N_4113,N_4079);
nor U7663 (N_7663,N_4914,N_5736);
nor U7664 (N_7664,N_4595,N_4446);
xor U7665 (N_7665,N_5190,N_5139);
nor U7666 (N_7666,N_5429,N_5671);
or U7667 (N_7667,N_5190,N_4762);
or U7668 (N_7668,N_5273,N_4972);
nor U7669 (N_7669,N_4687,N_4002);
nand U7670 (N_7670,N_5823,N_5763);
nor U7671 (N_7671,N_5613,N_5797);
and U7672 (N_7672,N_4561,N_4741);
nand U7673 (N_7673,N_4453,N_4755);
and U7674 (N_7674,N_5585,N_5323);
nand U7675 (N_7675,N_5238,N_5299);
and U7676 (N_7676,N_4437,N_4141);
nor U7677 (N_7677,N_5536,N_5637);
xor U7678 (N_7678,N_4380,N_5857);
nor U7679 (N_7679,N_4079,N_5123);
xnor U7680 (N_7680,N_5651,N_5822);
or U7681 (N_7681,N_4421,N_4826);
xor U7682 (N_7682,N_5278,N_5026);
nand U7683 (N_7683,N_4382,N_4305);
nor U7684 (N_7684,N_5396,N_5532);
or U7685 (N_7685,N_4179,N_5262);
xnor U7686 (N_7686,N_4782,N_4537);
nor U7687 (N_7687,N_4427,N_5737);
nor U7688 (N_7688,N_4920,N_5861);
nor U7689 (N_7689,N_5427,N_4198);
and U7690 (N_7690,N_5235,N_4426);
nor U7691 (N_7691,N_5561,N_4448);
nor U7692 (N_7692,N_4748,N_5198);
nor U7693 (N_7693,N_5460,N_5523);
nor U7694 (N_7694,N_4600,N_5929);
and U7695 (N_7695,N_4019,N_4121);
nand U7696 (N_7696,N_5012,N_4475);
xor U7697 (N_7697,N_5704,N_4403);
or U7698 (N_7698,N_4902,N_4321);
or U7699 (N_7699,N_5857,N_5151);
nand U7700 (N_7700,N_5825,N_5344);
and U7701 (N_7701,N_4218,N_4420);
and U7702 (N_7702,N_4128,N_4904);
xnor U7703 (N_7703,N_5399,N_5213);
nand U7704 (N_7704,N_4338,N_5390);
nor U7705 (N_7705,N_4618,N_5981);
xor U7706 (N_7706,N_5304,N_4177);
xor U7707 (N_7707,N_4601,N_5917);
nand U7708 (N_7708,N_5638,N_5132);
nand U7709 (N_7709,N_4397,N_5593);
nor U7710 (N_7710,N_4575,N_5925);
xor U7711 (N_7711,N_4049,N_4006);
or U7712 (N_7712,N_4587,N_5382);
or U7713 (N_7713,N_5415,N_5648);
or U7714 (N_7714,N_5300,N_4001);
or U7715 (N_7715,N_4606,N_4736);
or U7716 (N_7716,N_4334,N_4783);
nor U7717 (N_7717,N_4523,N_4207);
or U7718 (N_7718,N_5709,N_4925);
nor U7719 (N_7719,N_5863,N_5444);
and U7720 (N_7720,N_5111,N_4730);
xnor U7721 (N_7721,N_4872,N_4111);
nand U7722 (N_7722,N_4135,N_5922);
or U7723 (N_7723,N_4688,N_4471);
and U7724 (N_7724,N_4618,N_5855);
or U7725 (N_7725,N_4797,N_4179);
nand U7726 (N_7726,N_5118,N_4809);
xnor U7727 (N_7727,N_5917,N_5354);
and U7728 (N_7728,N_4619,N_5408);
xor U7729 (N_7729,N_5979,N_5238);
xor U7730 (N_7730,N_4587,N_5303);
nor U7731 (N_7731,N_4620,N_5194);
nor U7732 (N_7732,N_4786,N_5220);
or U7733 (N_7733,N_4028,N_5837);
or U7734 (N_7734,N_5482,N_4184);
xnor U7735 (N_7735,N_4991,N_5340);
xnor U7736 (N_7736,N_4737,N_5313);
or U7737 (N_7737,N_5929,N_4845);
nor U7738 (N_7738,N_4140,N_5127);
and U7739 (N_7739,N_5154,N_4544);
nor U7740 (N_7740,N_4453,N_5506);
nor U7741 (N_7741,N_5949,N_5594);
xnor U7742 (N_7742,N_4984,N_4722);
and U7743 (N_7743,N_5212,N_4238);
nor U7744 (N_7744,N_5997,N_5938);
and U7745 (N_7745,N_4201,N_4821);
nand U7746 (N_7746,N_5627,N_4124);
or U7747 (N_7747,N_4240,N_4190);
nand U7748 (N_7748,N_5828,N_4935);
or U7749 (N_7749,N_5117,N_4924);
and U7750 (N_7750,N_4086,N_5969);
nor U7751 (N_7751,N_4017,N_4539);
nor U7752 (N_7752,N_4330,N_5020);
xnor U7753 (N_7753,N_4954,N_5272);
or U7754 (N_7754,N_5967,N_4569);
nor U7755 (N_7755,N_5604,N_5369);
nand U7756 (N_7756,N_4776,N_4028);
nor U7757 (N_7757,N_5905,N_5233);
and U7758 (N_7758,N_4360,N_4088);
xnor U7759 (N_7759,N_5265,N_5288);
nor U7760 (N_7760,N_5272,N_5856);
nor U7761 (N_7761,N_4631,N_4140);
xnor U7762 (N_7762,N_4510,N_5119);
nand U7763 (N_7763,N_4819,N_5108);
and U7764 (N_7764,N_4432,N_5961);
xnor U7765 (N_7765,N_5576,N_5220);
and U7766 (N_7766,N_5010,N_5383);
and U7767 (N_7767,N_4385,N_5821);
and U7768 (N_7768,N_5101,N_5464);
xor U7769 (N_7769,N_5095,N_4384);
nor U7770 (N_7770,N_4123,N_4351);
nand U7771 (N_7771,N_4916,N_5412);
nor U7772 (N_7772,N_5714,N_5653);
and U7773 (N_7773,N_4408,N_4850);
nand U7774 (N_7774,N_5150,N_4208);
or U7775 (N_7775,N_4460,N_5139);
nor U7776 (N_7776,N_5184,N_5873);
nand U7777 (N_7777,N_4972,N_5088);
nand U7778 (N_7778,N_4604,N_4236);
nand U7779 (N_7779,N_5341,N_5638);
nor U7780 (N_7780,N_4161,N_4326);
or U7781 (N_7781,N_5136,N_5991);
nor U7782 (N_7782,N_5919,N_4160);
nand U7783 (N_7783,N_5674,N_4523);
xnor U7784 (N_7784,N_4773,N_4270);
and U7785 (N_7785,N_4087,N_4216);
and U7786 (N_7786,N_4576,N_4296);
and U7787 (N_7787,N_5420,N_4916);
and U7788 (N_7788,N_4152,N_5537);
or U7789 (N_7789,N_4394,N_5919);
and U7790 (N_7790,N_5345,N_5574);
nand U7791 (N_7791,N_5329,N_4575);
or U7792 (N_7792,N_4599,N_5247);
nor U7793 (N_7793,N_5002,N_5001);
or U7794 (N_7794,N_4167,N_5473);
nor U7795 (N_7795,N_4112,N_5546);
nor U7796 (N_7796,N_4255,N_4722);
nand U7797 (N_7797,N_4832,N_4991);
nor U7798 (N_7798,N_4789,N_5383);
nor U7799 (N_7799,N_4389,N_4383);
nand U7800 (N_7800,N_5372,N_4503);
or U7801 (N_7801,N_5336,N_4676);
nor U7802 (N_7802,N_4702,N_5012);
nor U7803 (N_7803,N_4053,N_5182);
or U7804 (N_7804,N_4489,N_5311);
nor U7805 (N_7805,N_4799,N_5167);
or U7806 (N_7806,N_5775,N_5087);
and U7807 (N_7807,N_4630,N_5545);
or U7808 (N_7808,N_4867,N_4626);
and U7809 (N_7809,N_4992,N_5666);
or U7810 (N_7810,N_4714,N_4824);
nor U7811 (N_7811,N_4538,N_4711);
and U7812 (N_7812,N_5416,N_4016);
and U7813 (N_7813,N_4693,N_5512);
nor U7814 (N_7814,N_4848,N_5685);
xnor U7815 (N_7815,N_4898,N_5520);
nor U7816 (N_7816,N_4159,N_5739);
xnor U7817 (N_7817,N_5102,N_5889);
nand U7818 (N_7818,N_4180,N_4668);
or U7819 (N_7819,N_4260,N_4785);
or U7820 (N_7820,N_5528,N_5237);
or U7821 (N_7821,N_4025,N_4473);
nor U7822 (N_7822,N_4506,N_5917);
or U7823 (N_7823,N_4720,N_4304);
or U7824 (N_7824,N_5020,N_5772);
nor U7825 (N_7825,N_4566,N_5589);
and U7826 (N_7826,N_4618,N_4414);
nor U7827 (N_7827,N_5500,N_5993);
xnor U7828 (N_7828,N_4834,N_5650);
or U7829 (N_7829,N_4020,N_5918);
xor U7830 (N_7830,N_5160,N_4560);
or U7831 (N_7831,N_4697,N_4099);
and U7832 (N_7832,N_5452,N_5702);
or U7833 (N_7833,N_5812,N_5901);
and U7834 (N_7834,N_4844,N_4502);
and U7835 (N_7835,N_4342,N_4718);
nand U7836 (N_7836,N_5431,N_5018);
nand U7837 (N_7837,N_4456,N_5616);
nand U7838 (N_7838,N_5652,N_5227);
or U7839 (N_7839,N_5428,N_4068);
and U7840 (N_7840,N_4309,N_4462);
nor U7841 (N_7841,N_4967,N_5776);
xnor U7842 (N_7842,N_4216,N_4391);
or U7843 (N_7843,N_4260,N_5960);
and U7844 (N_7844,N_4256,N_5921);
xor U7845 (N_7845,N_5471,N_4871);
xnor U7846 (N_7846,N_4037,N_4859);
and U7847 (N_7847,N_5912,N_4102);
xnor U7848 (N_7848,N_5423,N_4138);
nor U7849 (N_7849,N_4305,N_5670);
nand U7850 (N_7850,N_4002,N_5014);
or U7851 (N_7851,N_5485,N_5720);
nor U7852 (N_7852,N_4373,N_5079);
nand U7853 (N_7853,N_5904,N_5773);
nor U7854 (N_7854,N_5517,N_4729);
xnor U7855 (N_7855,N_4799,N_4858);
or U7856 (N_7856,N_5132,N_5951);
nand U7857 (N_7857,N_5404,N_5656);
nor U7858 (N_7858,N_4003,N_4200);
and U7859 (N_7859,N_5868,N_4287);
or U7860 (N_7860,N_4355,N_5041);
nor U7861 (N_7861,N_4457,N_4440);
nor U7862 (N_7862,N_4417,N_5085);
nand U7863 (N_7863,N_4687,N_4129);
nand U7864 (N_7864,N_4885,N_4150);
nand U7865 (N_7865,N_5622,N_4753);
or U7866 (N_7866,N_4689,N_5436);
nor U7867 (N_7867,N_4628,N_4590);
nand U7868 (N_7868,N_5959,N_5086);
and U7869 (N_7869,N_4734,N_5666);
or U7870 (N_7870,N_5059,N_4627);
and U7871 (N_7871,N_5099,N_5954);
or U7872 (N_7872,N_4280,N_5085);
or U7873 (N_7873,N_4363,N_4685);
or U7874 (N_7874,N_5293,N_4375);
and U7875 (N_7875,N_5655,N_5302);
xnor U7876 (N_7876,N_5351,N_4062);
or U7877 (N_7877,N_4628,N_5244);
nor U7878 (N_7878,N_5682,N_5985);
nor U7879 (N_7879,N_5175,N_5505);
or U7880 (N_7880,N_4765,N_4617);
nand U7881 (N_7881,N_5788,N_5588);
xor U7882 (N_7882,N_4729,N_5738);
nor U7883 (N_7883,N_5508,N_4033);
and U7884 (N_7884,N_5710,N_5586);
and U7885 (N_7885,N_5495,N_5203);
xnor U7886 (N_7886,N_4766,N_4898);
nor U7887 (N_7887,N_5293,N_5709);
xor U7888 (N_7888,N_5928,N_5640);
and U7889 (N_7889,N_4605,N_5012);
xnor U7890 (N_7890,N_5376,N_4149);
nor U7891 (N_7891,N_4990,N_5015);
nand U7892 (N_7892,N_4834,N_5497);
xnor U7893 (N_7893,N_4210,N_5095);
nor U7894 (N_7894,N_5347,N_5665);
and U7895 (N_7895,N_4636,N_5907);
xnor U7896 (N_7896,N_4763,N_4645);
and U7897 (N_7897,N_5214,N_4683);
xnor U7898 (N_7898,N_4419,N_4969);
nand U7899 (N_7899,N_4915,N_5107);
xnor U7900 (N_7900,N_5794,N_4580);
and U7901 (N_7901,N_4381,N_4471);
nor U7902 (N_7902,N_4710,N_5335);
and U7903 (N_7903,N_5139,N_5807);
nor U7904 (N_7904,N_5239,N_4149);
or U7905 (N_7905,N_5574,N_5275);
nand U7906 (N_7906,N_4490,N_5184);
nand U7907 (N_7907,N_5455,N_5752);
and U7908 (N_7908,N_5566,N_5942);
nand U7909 (N_7909,N_4274,N_5975);
or U7910 (N_7910,N_5481,N_5929);
xnor U7911 (N_7911,N_4116,N_5404);
nand U7912 (N_7912,N_4048,N_5835);
xor U7913 (N_7913,N_5135,N_5631);
nand U7914 (N_7914,N_5959,N_4252);
or U7915 (N_7915,N_4628,N_5628);
or U7916 (N_7916,N_5417,N_4392);
nand U7917 (N_7917,N_4005,N_4084);
or U7918 (N_7918,N_4727,N_4959);
or U7919 (N_7919,N_5224,N_5714);
xor U7920 (N_7920,N_4991,N_4175);
and U7921 (N_7921,N_5910,N_5113);
xor U7922 (N_7922,N_4478,N_4246);
and U7923 (N_7923,N_5224,N_4049);
and U7924 (N_7924,N_5355,N_4739);
or U7925 (N_7925,N_4364,N_4426);
nand U7926 (N_7926,N_5198,N_5161);
nor U7927 (N_7927,N_5765,N_5796);
or U7928 (N_7928,N_5495,N_5223);
nand U7929 (N_7929,N_5922,N_4263);
nor U7930 (N_7930,N_4743,N_4688);
and U7931 (N_7931,N_4010,N_4795);
xnor U7932 (N_7932,N_4572,N_4100);
nor U7933 (N_7933,N_5199,N_4980);
and U7934 (N_7934,N_4604,N_5060);
or U7935 (N_7935,N_4981,N_5358);
and U7936 (N_7936,N_5512,N_4115);
nor U7937 (N_7937,N_5542,N_5036);
nor U7938 (N_7938,N_5653,N_4864);
nand U7939 (N_7939,N_4800,N_4961);
nor U7940 (N_7940,N_4384,N_5893);
and U7941 (N_7941,N_5374,N_5237);
xnor U7942 (N_7942,N_4640,N_5878);
and U7943 (N_7943,N_5501,N_5141);
nor U7944 (N_7944,N_4827,N_5353);
and U7945 (N_7945,N_5941,N_4615);
xor U7946 (N_7946,N_4221,N_4127);
or U7947 (N_7947,N_5867,N_4241);
xor U7948 (N_7948,N_5099,N_5104);
and U7949 (N_7949,N_4205,N_4755);
xnor U7950 (N_7950,N_4404,N_4449);
xor U7951 (N_7951,N_5138,N_4281);
and U7952 (N_7952,N_5125,N_5308);
or U7953 (N_7953,N_5385,N_5187);
or U7954 (N_7954,N_5869,N_5693);
or U7955 (N_7955,N_4033,N_4059);
nor U7956 (N_7956,N_4424,N_4613);
nand U7957 (N_7957,N_4560,N_5950);
and U7958 (N_7958,N_4493,N_5113);
nand U7959 (N_7959,N_5534,N_4491);
nand U7960 (N_7960,N_5400,N_4752);
nand U7961 (N_7961,N_4415,N_4531);
nand U7962 (N_7962,N_4025,N_5569);
and U7963 (N_7963,N_4126,N_4619);
and U7964 (N_7964,N_4531,N_4831);
xor U7965 (N_7965,N_5917,N_5116);
xnor U7966 (N_7966,N_5366,N_4443);
nand U7967 (N_7967,N_4715,N_4561);
or U7968 (N_7968,N_5314,N_4212);
nor U7969 (N_7969,N_5680,N_4562);
nand U7970 (N_7970,N_5828,N_5043);
xnor U7971 (N_7971,N_5047,N_4463);
nand U7972 (N_7972,N_5901,N_5447);
and U7973 (N_7973,N_5520,N_5537);
nand U7974 (N_7974,N_5547,N_5465);
or U7975 (N_7975,N_4589,N_4327);
and U7976 (N_7976,N_4479,N_4478);
nand U7977 (N_7977,N_4087,N_5368);
and U7978 (N_7978,N_4559,N_5235);
or U7979 (N_7979,N_4923,N_4037);
nor U7980 (N_7980,N_4865,N_4251);
nor U7981 (N_7981,N_5193,N_4338);
or U7982 (N_7982,N_4006,N_4577);
nor U7983 (N_7983,N_4274,N_4095);
nor U7984 (N_7984,N_5160,N_4507);
xor U7985 (N_7985,N_5574,N_5508);
nand U7986 (N_7986,N_4012,N_5773);
and U7987 (N_7987,N_4578,N_5882);
and U7988 (N_7988,N_4877,N_5651);
or U7989 (N_7989,N_5489,N_5065);
nor U7990 (N_7990,N_5251,N_5225);
xnor U7991 (N_7991,N_4811,N_5175);
nor U7992 (N_7992,N_5638,N_4450);
and U7993 (N_7993,N_5893,N_5889);
nor U7994 (N_7994,N_4938,N_5169);
xor U7995 (N_7995,N_5324,N_5808);
nand U7996 (N_7996,N_4620,N_5571);
or U7997 (N_7997,N_5483,N_5636);
nand U7998 (N_7998,N_5861,N_4911);
or U7999 (N_7999,N_5856,N_4021);
or U8000 (N_8000,N_6316,N_7082);
nor U8001 (N_8001,N_7137,N_7861);
and U8002 (N_8002,N_6141,N_6317);
nand U8003 (N_8003,N_6655,N_6651);
nor U8004 (N_8004,N_7600,N_6627);
or U8005 (N_8005,N_7410,N_7700);
or U8006 (N_8006,N_6348,N_6350);
nor U8007 (N_8007,N_7123,N_6016);
nand U8008 (N_8008,N_7380,N_6387);
xnor U8009 (N_8009,N_6761,N_7807);
or U8010 (N_8010,N_6564,N_6437);
and U8011 (N_8011,N_6704,N_6267);
and U8012 (N_8012,N_6003,N_7844);
nand U8013 (N_8013,N_6413,N_6597);
nor U8014 (N_8014,N_6937,N_6185);
nand U8015 (N_8015,N_7465,N_6057);
nand U8016 (N_8016,N_6219,N_7183);
nor U8017 (N_8017,N_7179,N_7185);
xor U8018 (N_8018,N_7874,N_7783);
nand U8019 (N_8019,N_7502,N_7672);
or U8020 (N_8020,N_7392,N_7097);
xor U8021 (N_8021,N_6904,N_7613);
and U8022 (N_8022,N_6096,N_6641);
nand U8023 (N_8023,N_7327,N_7173);
or U8024 (N_8024,N_7751,N_7412);
nand U8025 (N_8025,N_6766,N_6539);
or U8026 (N_8026,N_7913,N_7681);
nor U8027 (N_8027,N_6553,N_6735);
nor U8028 (N_8028,N_7618,N_6355);
or U8029 (N_8029,N_6980,N_6780);
nor U8030 (N_8030,N_6715,N_7023);
or U8031 (N_8031,N_6441,N_7815);
and U8032 (N_8032,N_6371,N_7761);
nand U8033 (N_8033,N_7974,N_7434);
or U8034 (N_8034,N_7590,N_7586);
and U8035 (N_8035,N_6365,N_7995);
or U8036 (N_8036,N_7743,N_7556);
nor U8037 (N_8037,N_7814,N_6093);
and U8038 (N_8038,N_6943,N_6854);
and U8039 (N_8039,N_6646,N_6726);
nor U8040 (N_8040,N_7071,N_7174);
or U8041 (N_8041,N_7064,N_7947);
xnor U8042 (N_8042,N_6807,N_6446);
nand U8043 (N_8043,N_7225,N_7396);
xor U8044 (N_8044,N_7161,N_6664);
xor U8045 (N_8045,N_7129,N_7357);
nand U8046 (N_8046,N_7841,N_7270);
or U8047 (N_8047,N_7040,N_7448);
or U8048 (N_8048,N_7573,N_7331);
nor U8049 (N_8049,N_6588,N_6910);
xor U8050 (N_8050,N_6543,N_6369);
and U8051 (N_8051,N_7234,N_6128);
nor U8052 (N_8052,N_7541,N_6504);
or U8053 (N_8053,N_7239,N_6952);
or U8054 (N_8054,N_7004,N_7142);
xnor U8055 (N_8055,N_7182,N_7339);
or U8056 (N_8056,N_7926,N_7949);
and U8057 (N_8057,N_6183,N_7208);
nand U8058 (N_8058,N_6823,N_6740);
xnor U8059 (N_8059,N_7829,N_7847);
and U8060 (N_8060,N_6720,N_7468);
nor U8061 (N_8061,N_7399,N_6531);
or U8062 (N_8062,N_6188,N_7732);
or U8063 (N_8063,N_7398,N_7593);
xnor U8064 (N_8064,N_6161,N_7083);
nand U8065 (N_8065,N_7688,N_6940);
nand U8066 (N_8066,N_7450,N_6073);
nor U8067 (N_8067,N_7927,N_7092);
or U8068 (N_8068,N_6784,N_7351);
xor U8069 (N_8069,N_6657,N_7825);
or U8070 (N_8070,N_6024,N_7987);
and U8071 (N_8071,N_6250,N_7726);
xor U8072 (N_8072,N_7988,N_7637);
and U8073 (N_8073,N_7235,N_6748);
xnor U8074 (N_8074,N_7853,N_7858);
xnor U8075 (N_8075,N_7616,N_6861);
nand U8076 (N_8076,N_7651,N_6035);
nand U8077 (N_8077,N_7362,N_7203);
or U8078 (N_8078,N_6060,N_6934);
nand U8079 (N_8079,N_7824,N_6370);
nand U8080 (N_8080,N_6572,N_7155);
or U8081 (N_8081,N_7739,N_7568);
or U8082 (N_8082,N_6618,N_6260);
nand U8083 (N_8083,N_7971,N_6310);
nand U8084 (N_8084,N_6744,N_6044);
nand U8085 (N_8085,N_6589,N_7912);
and U8086 (N_8086,N_7777,N_7831);
or U8087 (N_8087,N_7958,N_6966);
and U8088 (N_8088,N_7966,N_6635);
xor U8089 (N_8089,N_6663,N_6283);
or U8090 (N_8090,N_6661,N_6909);
nor U8091 (N_8091,N_6075,N_7745);
xor U8092 (N_8092,N_6351,N_7017);
or U8093 (N_8093,N_7488,N_6678);
xor U8094 (N_8094,N_6489,N_7285);
and U8095 (N_8095,N_7849,N_7310);
nor U8096 (N_8096,N_6939,N_6319);
and U8097 (N_8097,N_6825,N_7516);
nand U8098 (N_8098,N_7609,N_7854);
or U8099 (N_8099,N_6401,N_7605);
nor U8100 (N_8100,N_7232,N_7051);
xor U8101 (N_8101,N_7445,N_7400);
or U8102 (N_8102,N_7116,N_6047);
nor U8103 (N_8103,N_7812,N_6235);
or U8104 (N_8104,N_6533,N_6237);
nand U8105 (N_8105,N_7126,N_7521);
or U8106 (N_8106,N_6231,N_7774);
or U8107 (N_8107,N_6674,N_6546);
nor U8108 (N_8108,N_6366,N_6195);
xnor U8109 (N_8109,N_6200,N_6066);
and U8110 (N_8110,N_6116,N_7524);
and U8111 (N_8111,N_7619,N_7149);
and U8112 (N_8112,N_6115,N_7319);
xnor U8113 (N_8113,N_7638,N_7081);
nor U8114 (N_8114,N_6711,N_7391);
xor U8115 (N_8115,N_7589,N_6160);
and U8116 (N_8116,N_7134,N_7472);
or U8117 (N_8117,N_6760,N_6942);
nor U8118 (N_8118,N_6957,N_6776);
or U8119 (N_8119,N_7230,N_7295);
or U8120 (N_8120,N_6520,N_6154);
nand U8121 (N_8121,N_6473,N_6841);
nor U8122 (N_8122,N_6261,N_6105);
or U8123 (N_8123,N_7411,N_7715);
and U8124 (N_8124,N_6361,N_7650);
and U8125 (N_8125,N_6425,N_6282);
xor U8126 (N_8126,N_7467,N_7094);
nand U8127 (N_8127,N_6965,N_7705);
or U8128 (N_8128,N_6148,N_6037);
xnor U8129 (N_8129,N_7304,N_6168);
and U8130 (N_8130,N_6835,N_6503);
or U8131 (N_8131,N_7517,N_7397);
xor U8132 (N_8132,N_6617,N_7557);
or U8133 (N_8133,N_6084,N_6118);
and U8134 (N_8134,N_7447,N_6220);
and U8135 (N_8135,N_6969,N_7067);
xnor U8136 (N_8136,N_7390,N_6392);
xor U8137 (N_8137,N_6254,N_6100);
xnor U8138 (N_8138,N_7477,N_7099);
xnor U8139 (N_8139,N_6330,N_7943);
nor U8140 (N_8140,N_6967,N_6038);
nand U8141 (N_8141,N_7163,N_6284);
nand U8142 (N_8142,N_6155,N_7406);
nand U8143 (N_8143,N_7626,N_6376);
or U8144 (N_8144,N_7010,N_6997);
nor U8145 (N_8145,N_6698,N_6029);
or U8146 (N_8146,N_7317,N_6139);
and U8147 (N_8147,N_6872,N_6397);
xor U8148 (N_8148,N_6768,N_6022);
or U8149 (N_8149,N_7654,N_7728);
and U8150 (N_8150,N_6988,N_7003);
xor U8151 (N_8151,N_6332,N_7817);
and U8152 (N_8152,N_7997,N_6307);
xor U8153 (N_8153,N_6810,N_7222);
xnor U8154 (N_8154,N_6290,N_7444);
xor U8155 (N_8155,N_6379,N_7537);
nand U8156 (N_8156,N_6978,N_7627);
nand U8157 (N_8157,N_6121,N_6295);
or U8158 (N_8158,N_6547,N_7454);
and U8159 (N_8159,N_6731,N_6848);
and U8160 (N_8160,N_6492,N_7559);
or U8161 (N_8161,N_7551,N_6245);
or U8162 (N_8162,N_7826,N_7113);
or U8163 (N_8163,N_7522,N_6620);
nor U8164 (N_8164,N_6278,N_7053);
xnor U8165 (N_8165,N_6318,N_6789);
nor U8166 (N_8166,N_7242,N_6710);
and U8167 (N_8167,N_7676,N_7975);
and U8168 (N_8168,N_6189,N_6689);
or U8169 (N_8169,N_6866,N_7429);
or U8170 (N_8170,N_6275,N_6672);
nand U8171 (N_8171,N_6878,N_6706);
nor U8172 (N_8172,N_6686,N_7901);
nand U8173 (N_8173,N_7070,N_6021);
xnor U8174 (N_8174,N_6718,N_7529);
xnor U8175 (N_8175,N_6809,N_6530);
or U8176 (N_8176,N_7560,N_6637);
or U8177 (N_8177,N_7671,N_7254);
or U8178 (N_8178,N_7193,N_7436);
nand U8179 (N_8179,N_7005,N_7819);
or U8180 (N_8180,N_7820,N_6994);
xnor U8181 (N_8181,N_6758,N_6450);
nor U8182 (N_8182,N_7227,N_7439);
or U8183 (N_8183,N_7490,N_7716);
or U8184 (N_8184,N_6174,N_7850);
or U8185 (N_8185,N_6049,N_6683);
or U8186 (N_8186,N_7887,N_7891);
nand U8187 (N_8187,N_6505,N_6347);
nand U8188 (N_8188,N_6578,N_6359);
nand U8189 (N_8189,N_7816,N_6805);
or U8190 (N_8190,N_6039,N_7684);
and U8191 (N_8191,N_7896,N_7701);
nor U8192 (N_8192,N_6565,N_7917);
nand U8193 (N_8193,N_6747,N_7859);
nor U8194 (N_8194,N_6569,N_6729);
or U8195 (N_8195,N_7255,N_7598);
nand U8196 (N_8196,N_7121,N_7367);
nor U8197 (N_8197,N_6325,N_7523);
or U8198 (N_8198,N_7389,N_7508);
and U8199 (N_8199,N_6871,N_7544);
xor U8200 (N_8200,N_7822,N_6822);
and U8201 (N_8201,N_6297,N_7915);
and U8202 (N_8202,N_6728,N_7779);
or U8203 (N_8203,N_7000,N_6570);
nor U8204 (N_8204,N_6793,N_6501);
nor U8205 (N_8205,N_6915,N_6935);
nor U8206 (N_8206,N_6532,N_6490);
nand U8207 (N_8207,N_6333,N_7476);
xor U8208 (N_8208,N_7496,N_6938);
nand U8209 (N_8209,N_6725,N_7888);
nand U8210 (N_8210,N_7109,N_6893);
and U8211 (N_8211,N_7561,N_6309);
nor U8212 (N_8212,N_7757,N_7595);
and U8213 (N_8213,N_6465,N_7018);
nand U8214 (N_8214,N_6455,N_6127);
xor U8215 (N_8215,N_6415,N_6156);
and U8216 (N_8216,N_7525,N_7921);
xor U8217 (N_8217,N_6903,N_6676);
nand U8218 (N_8218,N_6847,N_7355);
xor U8219 (N_8219,N_6454,N_7273);
nor U8220 (N_8220,N_7119,N_7281);
or U8221 (N_8221,N_7002,N_6803);
xor U8222 (N_8222,N_6285,N_6433);
and U8223 (N_8223,N_6767,N_7372);
or U8224 (N_8224,N_6251,N_7827);
nand U8225 (N_8225,N_6920,N_6364);
nand U8226 (N_8226,N_7704,N_7293);
and U8227 (N_8227,N_7167,N_6380);
or U8228 (N_8228,N_6898,N_7275);
and U8229 (N_8229,N_7007,N_6989);
nand U8230 (N_8230,N_6917,N_6403);
or U8231 (N_8231,N_7922,N_7581);
nand U8232 (N_8232,N_7687,N_7625);
and U8233 (N_8233,N_6534,N_6106);
or U8234 (N_8234,N_6449,N_7299);
nor U8235 (N_8235,N_6311,N_6953);
xnor U8236 (N_8236,N_6368,N_7973);
or U8237 (N_8237,N_7001,N_7158);
nor U8238 (N_8238,N_7286,N_6113);
nand U8239 (N_8239,N_7811,N_7706);
or U8240 (N_8240,N_6268,N_6101);
xnor U8241 (N_8241,N_6818,N_7754);
xor U8242 (N_8242,N_7440,N_7152);
nor U8243 (N_8243,N_6613,N_6270);
and U8244 (N_8244,N_7838,N_6973);
or U8245 (N_8245,N_7309,N_7933);
nand U8246 (N_8246,N_7624,N_7146);
nand U8247 (N_8247,N_7311,N_7130);
xnor U8248 (N_8248,N_6352,N_6599);
and U8249 (N_8249,N_7056,N_6070);
and U8250 (N_8250,N_7699,N_7668);
and U8251 (N_8251,N_7878,N_7528);
nor U8252 (N_8252,N_7833,N_6493);
xnor U8253 (N_8253,N_7417,N_6811);
nor U8254 (N_8254,N_7170,N_6480);
or U8255 (N_8255,N_6144,N_6559);
xnor U8256 (N_8256,N_7930,N_6839);
nor U8257 (N_8257,N_6542,N_6552);
nor U8258 (N_8258,N_6193,N_7159);
xnor U8259 (N_8259,N_6315,N_7283);
nor U8260 (N_8260,N_7879,N_6558);
xor U8261 (N_8261,N_6407,N_7897);
xor U8262 (N_8262,N_6293,N_7721);
nor U8263 (N_8263,N_6964,N_7249);
nand U8264 (N_8264,N_6582,N_7652);
xor U8265 (N_8265,N_7553,N_7505);
or U8266 (N_8266,N_7571,N_7967);
nand U8267 (N_8267,N_6344,N_7312);
xnor U8268 (N_8268,N_6264,N_7923);
nand U8269 (N_8269,N_6962,N_7375);
xor U8270 (N_8270,N_6085,N_6630);
or U8271 (N_8271,N_7769,N_7359);
nor U8272 (N_8272,N_6308,N_6305);
and U8273 (N_8273,N_7370,N_7482);
and U8274 (N_8274,N_7512,N_6636);
xnor U8275 (N_8275,N_7122,N_7846);
xnor U8276 (N_8276,N_7938,N_6198);
or U8277 (N_8277,N_6230,N_7431);
and U8278 (N_8278,N_7307,N_6521);
nor U8279 (N_8279,N_6779,N_6502);
xnor U8280 (N_8280,N_7452,N_6701);
nand U8281 (N_8281,N_6573,N_6152);
and U8282 (N_8282,N_6296,N_6723);
nor U8283 (N_8283,N_7368,N_7201);
nand U8284 (N_8284,N_7449,N_6068);
xnor U8285 (N_8285,N_6402,N_6273);
or U8286 (N_8286,N_7025,N_7218);
nand U8287 (N_8287,N_7112,N_7669);
or U8288 (N_8288,N_6363,N_6615);
and U8289 (N_8289,N_6216,N_7114);
and U8290 (N_8290,N_7583,N_6619);
nand U8291 (N_8291,N_6874,N_6142);
or U8292 (N_8292,N_6255,N_7178);
nor U8293 (N_8293,N_7670,N_6336);
and U8294 (N_8294,N_7607,N_6061);
or U8295 (N_8295,N_7451,N_6751);
xor U8296 (N_8296,N_6561,N_7555);
xnor U8297 (N_8297,N_7656,N_6081);
and U8298 (N_8298,N_6287,N_7863);
or U8299 (N_8299,N_6604,N_7379);
and U8300 (N_8300,N_6765,N_6529);
nand U8301 (N_8301,N_6756,N_6467);
nor U8302 (N_8302,N_7291,N_7526);
or U8303 (N_8303,N_7127,N_6932);
or U8304 (N_8304,N_7959,N_6692);
or U8305 (N_8305,N_6399,N_7442);
nor U8306 (N_8306,N_7793,N_7100);
or U8307 (N_8307,N_7383,N_6536);
xor U8308 (N_8308,N_7107,N_6867);
nor U8309 (N_8309,N_6563,N_6643);
or U8310 (N_8310,N_7437,N_6858);
nand U8311 (N_8311,N_7803,N_7903);
nor U8312 (N_8312,N_6968,N_6693);
nand U8313 (N_8313,N_7946,N_7247);
xnor U8314 (N_8314,N_7993,N_6707);
and U8315 (N_8315,N_6474,N_6591);
or U8316 (N_8316,N_7674,N_7347);
and U8317 (N_8317,N_7691,N_6991);
nand U8318 (N_8318,N_6621,N_7510);
and U8319 (N_8319,N_7198,N_7271);
or U8320 (N_8320,N_7998,N_6528);
nor U8321 (N_8321,N_6484,N_6448);
nor U8322 (N_8322,N_7799,N_6451);
nor U8323 (N_8323,N_6659,N_6056);
nor U8324 (N_8324,N_7349,N_7723);
xor U8325 (N_8325,N_7022,N_7519);
and U8326 (N_8326,N_6164,N_7186);
nor U8327 (N_8327,N_7258,N_6120);
xnor U8328 (N_8328,N_7176,N_6009);
and U8329 (N_8329,N_7763,N_6905);
or U8330 (N_8330,N_7322,N_7061);
and U8331 (N_8331,N_6289,N_7033);
nand U8332 (N_8332,N_7895,N_7038);
xor U8333 (N_8333,N_6855,N_7564);
and U8334 (N_8334,N_6713,N_7089);
or U8335 (N_8335,N_6395,N_7032);
nor U8336 (N_8336,N_7160,N_7640);
or U8337 (N_8337,N_7306,N_6705);
nor U8338 (N_8338,N_7765,N_7197);
nand U8339 (N_8339,N_7257,N_7087);
xor U8340 (N_8340,N_6069,N_7011);
or U8341 (N_8341,N_7219,N_7401);
and U8342 (N_8342,N_6236,N_7334);
nor U8343 (N_8343,N_6945,N_7353);
xnor U8344 (N_8344,N_7013,N_6622);
xor U8345 (N_8345,N_7869,N_7288);
xor U8346 (N_8346,N_7981,N_6378);
and U8347 (N_8347,N_6034,N_6721);
xnor U8348 (N_8348,N_6795,N_7382);
or U8349 (N_8349,N_7297,N_6648);
or U8350 (N_8350,N_6986,N_7287);
nor U8351 (N_8351,N_7904,N_6476);
nand U8352 (N_8352,N_7864,N_6125);
xnor U8353 (N_8353,N_6794,N_7366);
nor U8354 (N_8354,N_7026,N_6491);
nor U8355 (N_8355,N_7474,N_7060);
nor U8356 (N_8356,N_7860,N_7683);
and U8357 (N_8357,N_7084,N_6340);
nand U8358 (N_8358,N_7711,N_6036);
and U8359 (N_8359,N_7570,N_7373);
nand U8360 (N_8360,N_7873,N_6567);
or U8361 (N_8361,N_6716,N_6912);
or U8362 (N_8362,N_7809,N_7117);
nand U8363 (N_8363,N_6593,N_6481);
nand U8364 (N_8364,N_6027,N_7356);
and U8365 (N_8365,N_7991,N_6208);
nor U8366 (N_8366,N_6843,N_7898);
xor U8367 (N_8367,N_6896,N_6797);
nor U8368 (N_8368,N_6218,N_7918);
nor U8369 (N_8369,N_6354,N_6649);
nand U8370 (N_8370,N_6444,N_7916);
and U8371 (N_8371,N_6217,N_6124);
xnor U8372 (N_8372,N_6614,N_6733);
or U8373 (N_8373,N_6771,N_7133);
nor U8374 (N_8374,N_7620,N_6322);
xor U8375 (N_8375,N_7493,N_6829);
nor U8376 (N_8376,N_7952,N_7233);
xnor U8377 (N_8377,N_6211,N_7028);
xor U8378 (N_8378,N_7352,N_6694);
or U8379 (N_8379,N_7143,N_6343);
nor U8380 (N_8380,N_6181,N_6000);
nand U8381 (N_8381,N_7481,N_7635);
or U8382 (N_8382,N_6468,N_7144);
nor U8383 (N_8383,N_6998,N_6479);
and U8384 (N_8384,N_6091,N_7348);
nor U8385 (N_8385,N_6688,N_7939);
nor U8386 (N_8386,N_7657,N_7115);
xor U8387 (N_8387,N_6891,N_7756);
nor U8388 (N_8388,N_6040,N_6372);
or U8389 (N_8389,N_6695,N_6439);
nor U8390 (N_8390,N_7469,N_6870);
nand U8391 (N_8391,N_6717,N_6400);
or U8392 (N_8392,N_6431,N_7466);
xnor U8393 (N_8393,N_6382,N_7851);
nand U8394 (N_8394,N_6916,N_6135);
or U8395 (N_8395,N_6052,N_7986);
and U8396 (N_8396,N_6927,N_7767);
and U8397 (N_8397,N_6851,N_6232);
nor U8398 (N_8398,N_7345,N_7889);
nand U8399 (N_8399,N_7909,N_7792);
xor U8400 (N_8400,N_7579,N_7354);
xnor U8401 (N_8401,N_7810,N_7314);
nand U8402 (N_8402,N_6919,N_6781);
and U8403 (N_8403,N_6901,N_7259);
xnor U8404 (N_8404,N_6712,N_6117);
nor U8405 (N_8405,N_6119,N_6583);
and U8406 (N_8406,N_6418,N_6025);
nand U8407 (N_8407,N_7950,N_6110);
or U8408 (N_8408,N_6524,N_6426);
xnor U8409 (N_8409,N_7263,N_7835);
nor U8410 (N_8410,N_6580,N_6190);
or U8411 (N_8411,N_7712,N_7268);
nand U8412 (N_8412,N_6889,N_7479);
nand U8413 (N_8413,N_6459,N_6754);
nor U8414 (N_8414,N_7527,N_7171);
nand U8415 (N_8415,N_7985,N_7588);
and U8416 (N_8416,N_7404,N_6147);
or U8417 (N_8417,N_6033,N_7877);
nor U8418 (N_8418,N_7250,N_7199);
xor U8419 (N_8419,N_6629,N_7666);
nor U8420 (N_8420,N_6323,N_7329);
nor U8421 (N_8421,N_6987,N_6517);
and U8422 (N_8422,N_6955,N_7303);
and U8423 (N_8423,N_7885,N_6083);
and U8424 (N_8424,N_7630,N_6186);
nor U8425 (N_8425,N_7994,N_6172);
or U8426 (N_8426,N_6007,N_7486);
and U8427 (N_8427,N_7238,N_7934);
nor U8428 (N_8428,N_7782,N_6436);
or U8429 (N_8429,N_7580,N_6242);
or U8430 (N_8430,N_6071,N_7507);
and U8431 (N_8431,N_6951,N_6259);
and U8432 (N_8432,N_7982,N_7643);
and U8433 (N_8433,N_7484,N_6814);
nand U8434 (N_8434,N_6865,N_7105);
xnor U8435 (N_8435,N_6201,N_6933);
xor U8436 (N_8436,N_7008,N_6194);
nand U8437 (N_8437,N_7243,N_6681);
or U8438 (N_8438,N_6487,N_7393);
and U8439 (N_8439,N_6743,N_7072);
nand U8440 (N_8440,N_7455,N_7868);
nand U8441 (N_8441,N_6249,N_7220);
nand U8442 (N_8442,N_6157,N_7292);
and U8443 (N_8443,N_7628,N_6638);
or U8444 (N_8444,N_6162,N_6687);
nand U8445 (N_8445,N_6385,N_6581);
or U8446 (N_8446,N_6857,N_6586);
xor U8447 (N_8447,N_6603,N_6846);
or U8448 (N_8448,N_7473,N_6443);
nor U8449 (N_8449,N_7766,N_7843);
and U8450 (N_8450,N_7009,N_7795);
nor U8451 (N_8451,N_7956,N_6452);
or U8452 (N_8452,N_6875,N_6755);
xnor U8453 (N_8453,N_6244,N_7096);
nor U8454 (N_8454,N_7741,N_6107);
nand U8455 (N_8455,N_6028,N_6420);
nor U8456 (N_8456,N_7344,N_6778);
nor U8457 (N_8457,N_7886,N_6067);
xor U8458 (N_8458,N_6335,N_7491);
and U8459 (N_8459,N_6178,N_6527);
and U8460 (N_8460,N_6928,N_7747);
or U8461 (N_8461,N_6213,N_7623);
and U8462 (N_8462,N_7301,N_6908);
or U8463 (N_8463,N_6849,N_7495);
xnor U8464 (N_8464,N_7103,N_6170);
or U8465 (N_8465,N_6082,N_7667);
and U8466 (N_8466,N_6421,N_6662);
xor U8467 (N_8467,N_7582,N_6764);
nand U8468 (N_8468,N_7832,N_6281);
or U8469 (N_8469,N_7591,N_6167);
nor U8470 (N_8470,N_7030,N_6384);
or U8471 (N_8471,N_6985,N_7693);
nand U8472 (N_8472,N_7603,N_6516);
xor U8473 (N_8473,N_6471,N_7499);
xnor U8474 (N_8474,N_7714,N_7980);
nand U8475 (N_8475,N_7664,N_7217);
xor U8476 (N_8476,N_7604,N_6538);
xnor U8477 (N_8477,N_6961,N_7677);
xor U8478 (N_8478,N_6763,N_7661);
nor U8479 (N_8479,N_7276,N_7929);
nand U8480 (N_8480,N_6390,N_6222);
xor U8481 (N_8481,N_6541,N_7644);
nor U8482 (N_8482,N_6821,N_7039);
xnor U8483 (N_8483,N_7168,N_7074);
and U8484 (N_8484,N_6227,N_6819);
and U8485 (N_8485,N_7685,N_6277);
and U8486 (N_8486,N_6478,N_6470);
nor U8487 (N_8487,N_6048,N_7223);
nand U8488 (N_8488,N_7088,N_7463);
nor U8489 (N_8489,N_6959,N_6302);
and U8490 (N_8490,N_6461,N_7043);
nor U8491 (N_8491,N_7269,N_7252);
nor U8492 (N_8492,N_6922,N_6177);
nor U8493 (N_8493,N_6499,N_7646);
and U8494 (N_8494,N_7698,N_7574);
xor U8495 (N_8495,N_7248,N_7024);
xor U8496 (N_8496,N_7662,N_7386);
nand U8497 (N_8497,N_7020,N_7786);
and U8498 (N_8498,N_6611,N_7717);
nand U8499 (N_8499,N_6796,N_7789);
nand U8500 (N_8500,N_6554,N_7231);
xor U8501 (N_8501,N_6523,N_7050);
or U8502 (N_8502,N_6640,N_7945);
or U8503 (N_8503,N_6008,N_6512);
nand U8504 (N_8504,N_6634,N_7979);
nor U8505 (N_8505,N_7318,N_7280);
nand U8506 (N_8506,N_6948,N_7961);
or U8507 (N_8507,N_7139,N_6958);
nor U8508 (N_8508,N_6745,N_6815);
and U8509 (N_8509,N_7702,N_6954);
or U8510 (N_8510,N_6266,N_6832);
and U8511 (N_8511,N_7065,N_7110);
and U8512 (N_8512,N_6381,N_7044);
and U8513 (N_8513,N_6132,N_7421);
xor U8514 (N_8514,N_6430,N_6551);
nor U8515 (N_8515,N_6233,N_6054);
and U8516 (N_8516,N_7498,N_6329);
and U8517 (N_8517,N_7965,N_6182);
and U8518 (N_8518,N_7776,N_6880);
and U8519 (N_8519,N_6753,N_7575);
nor U8520 (N_8520,N_7830,N_7098);
and U8521 (N_8521,N_6804,N_6191);
nand U8522 (N_8522,N_7430,N_7012);
or U8523 (N_8523,N_7006,N_6863);
nand U8524 (N_8524,N_6500,N_6398);
xor U8525 (N_8525,N_6288,N_6816);
nor U8526 (N_8526,N_7572,N_7632);
nand U8527 (N_8527,N_6393,N_6666);
nor U8528 (N_8528,N_7634,N_7015);
or U8529 (N_8529,N_7343,N_7749);
or U8530 (N_8530,N_6790,N_7104);
nor U8531 (N_8531,N_6228,N_6862);
nor U8532 (N_8532,N_7215,N_6383);
xnor U8533 (N_8533,N_6435,N_7515);
xnor U8534 (N_8534,N_7759,N_6102);
and U8535 (N_8535,N_7944,N_7682);
nor U8536 (N_8536,N_7780,N_7497);
nand U8537 (N_8537,N_6650,N_7424);
or U8538 (N_8538,N_6405,N_6339);
or U8539 (N_8539,N_6051,N_6596);
nand U8540 (N_8540,N_7645,N_7378);
nor U8541 (N_8541,N_7261,N_6262);
nor U8542 (N_8542,N_6356,N_7135);
or U8543 (N_8543,N_7852,N_6457);
nor U8544 (N_8544,N_7880,N_7462);
nand U8545 (N_8545,N_6785,N_7925);
xor U8546 (N_8546,N_7278,N_7781);
nand U8547 (N_8547,N_6786,N_6126);
xor U8548 (N_8548,N_6508,N_6321);
xnor U8549 (N_8549,N_6647,N_7256);
xor U8550 (N_8550,N_6294,N_6442);
or U8551 (N_8551,N_6104,N_6109);
nand U8552 (N_8552,N_6279,N_6675);
or U8553 (N_8553,N_6388,N_6652);
and U8554 (N_8554,N_6046,N_6014);
xor U8555 (N_8555,N_7565,N_7882);
and U8556 (N_8556,N_7642,N_7325);
and U8557 (N_8557,N_7435,N_7722);
nor U8558 (N_8558,N_7867,N_6345);
and U8559 (N_8559,N_6496,N_6353);
nand U8560 (N_8560,N_7057,N_7246);
and U8561 (N_8561,N_7118,N_6010);
xnor U8562 (N_8562,N_7147,N_6497);
nand U8563 (N_8563,N_7622,N_7709);
xnor U8564 (N_8564,N_7875,N_6263);
nor U8565 (N_8565,N_7266,N_7407);
or U8566 (N_8566,N_7518,N_7905);
xnor U8567 (N_8567,N_6026,N_6902);
nor U8568 (N_8568,N_6820,N_7409);
nor U8569 (N_8569,N_6859,N_7125);
or U8570 (N_8570,N_7414,N_7920);
and U8571 (N_8571,N_6409,N_7441);
and U8572 (N_8572,N_7342,N_7533);
xnor U8573 (N_8573,N_6328,N_7336);
and U8574 (N_8574,N_7856,N_7210);
nand U8575 (N_8575,N_6498,N_7942);
and U8576 (N_8576,N_7106,N_6013);
xor U8577 (N_8577,N_6445,N_6946);
nor U8578 (N_8578,N_7029,N_6548);
nand U8579 (N_8579,N_7511,N_7804);
or U8580 (N_8580,N_7207,N_7140);
or U8581 (N_8581,N_7984,N_6114);
xor U8582 (N_8582,N_6462,N_6571);
nor U8583 (N_8583,N_7744,N_6824);
and U8584 (N_8584,N_6970,N_6252);
nor U8585 (N_8585,N_6685,N_6975);
nor U8586 (N_8586,N_7494,N_6817);
or U8587 (N_8587,N_6065,N_6853);
xor U8588 (N_8588,N_7720,N_7066);
and U8589 (N_8589,N_6412,N_6601);
nor U8590 (N_8590,N_6977,N_7154);
and U8591 (N_8591,N_6031,N_6624);
and U8592 (N_8592,N_7694,N_7175);
nand U8593 (N_8593,N_7606,N_7244);
nand U8594 (N_8594,N_7848,N_7131);
xor U8595 (N_8595,N_7836,N_6724);
nand U8596 (N_8596,N_6004,N_7734);
or U8597 (N_8597,N_6140,N_7021);
and U8598 (N_8598,N_7753,N_6488);
and U8599 (N_8599,N_6783,N_6924);
and U8600 (N_8600,N_6298,N_6112);
nand U8601 (N_8601,N_6292,N_7536);
nand U8602 (N_8602,N_7290,N_7631);
or U8603 (N_8603,N_6782,N_7775);
xnor U8604 (N_8604,N_6367,N_7999);
nand U8605 (N_8605,N_6173,N_7762);
and U8606 (N_8606,N_7313,N_6736);
or U8607 (N_8607,N_7554,N_7475);
nor U8608 (N_8608,N_7755,N_7673);
and U8609 (N_8609,N_7594,N_6732);
xnor U8610 (N_8610,N_7394,N_6850);
nor U8611 (N_8611,N_7156,N_6394);
nand U8612 (N_8612,N_6830,N_7423);
nand U8613 (N_8613,N_7438,N_6568);
xnor U8614 (N_8614,N_7940,N_6423);
nor U8615 (N_8615,N_7101,N_6894);
nor U8616 (N_8616,N_7138,N_6005);
or U8617 (N_8617,N_6690,N_6671);
and U8618 (N_8618,N_7893,N_6626);
nand U8619 (N_8619,N_6628,N_6092);
and U8620 (N_8620,N_7052,N_7371);
nor U8621 (N_8621,N_7090,N_7549);
xnor U8622 (N_8622,N_7298,N_6246);
and U8623 (N_8623,N_7460,N_6134);
nor U8624 (N_8624,N_7773,N_7718);
or U8625 (N_8625,N_6749,N_6176);
xor U8626 (N_8626,N_7737,N_6873);
xor U8627 (N_8627,N_6709,N_7813);
nand U8628 (N_8628,N_6773,N_7871);
nor U8629 (N_8629,N_6206,N_6525);
xnor U8630 (N_8630,N_6377,N_7483);
nand U8631 (N_8631,N_6812,N_6892);
or U8632 (N_8632,N_7708,N_6752);
nand U8633 (N_8633,N_6600,N_6607);
xor U8634 (N_8634,N_6654,N_7086);
nor U8635 (N_8635,N_6845,N_7976);
and U8636 (N_8636,N_6179,N_7470);
nor U8637 (N_8637,N_6837,N_7457);
nor U8638 (N_8638,N_6349,N_7617);
and U8639 (N_8639,N_7660,N_6475);
or U8640 (N_8640,N_7531,N_6136);
nor U8641 (N_8641,N_6722,N_6990);
and U8642 (N_8642,N_7937,N_6881);
xor U8643 (N_8643,N_6575,N_7200);
xnor U8644 (N_8644,N_7190,N_6608);
nor U8645 (N_8645,N_6895,N_6159);
nor U8646 (N_8646,N_7954,N_6800);
or U8647 (N_8647,N_7596,N_6240);
or U8648 (N_8648,N_7790,N_7500);
nor U8649 (N_8649,N_6682,N_7772);
xor U8650 (N_8650,N_7818,N_6131);
nor U8651 (N_8651,N_6730,N_7791);
nand U8652 (N_8652,N_6788,N_7592);
or U8653 (N_8653,N_6196,N_7209);
nand U8654 (N_8654,N_7166,N_6708);
nor U8655 (N_8655,N_6058,N_6313);
and U8656 (N_8656,N_6015,N_6974);
nor U8657 (N_8657,N_7308,N_6691);
xnor U8658 (N_8658,N_7187,N_6466);
or U8659 (N_8659,N_6631,N_6460);
nand U8660 (N_8660,N_7204,N_6949);
nand U8661 (N_8661,N_6616,N_6984);
and U8662 (N_8662,N_6257,N_6001);
and U8663 (N_8663,N_7487,N_7719);
or U8664 (N_8664,N_7211,N_7153);
nand U8665 (N_8665,N_6404,N_6373);
or U8666 (N_8666,N_7216,N_7610);
nor U8667 (N_8667,N_6312,N_7953);
nor U8668 (N_8668,N_6234,N_7196);
or U8669 (N_8669,N_7501,N_6304);
nor U8670 (N_8670,N_6703,N_7713);
nor U8671 (N_8671,N_6700,N_6203);
and U8672 (N_8672,N_7328,N_6535);
nor U8673 (N_8673,N_6963,N_6981);
nor U8674 (N_8674,N_7461,N_6757);
or U8675 (N_8675,N_7653,N_7338);
nand U8676 (N_8676,N_7045,N_6750);
nand U8677 (N_8677,N_7686,N_6680);
xor U8678 (N_8678,N_7608,N_7226);
or U8679 (N_8679,N_6950,N_7535);
and U8680 (N_8680,N_6210,N_6019);
nand U8681 (N_8681,N_7908,N_6165);
nand U8682 (N_8682,N_6598,N_6215);
or U8683 (N_8683,N_6006,N_7710);
nor U8684 (N_8684,N_6099,N_7963);
xor U8685 (N_8685,N_6472,N_7735);
nor U8686 (N_8686,N_7894,N_7315);
xor U8687 (N_8687,N_6204,N_6074);
nor U8688 (N_8688,N_7805,N_7689);
and U8689 (N_8689,N_7048,N_6224);
nor U8690 (N_8690,N_7162,N_7188);
or U8691 (N_8691,N_6396,N_6602);
or U8692 (N_8692,N_7679,N_6320);
nand U8693 (N_8693,N_7037,N_6375);
nor U8694 (N_8694,N_7778,N_7881);
and U8695 (N_8695,N_6108,N_6737);
nor U8696 (N_8696,N_6555,N_7282);
nor U8697 (N_8697,N_6146,N_6639);
xnor U8698 (N_8698,N_7614,N_7458);
or U8699 (N_8699,N_6791,N_6677);
nor U8700 (N_8700,N_7340,N_7797);
and U8701 (N_8701,N_6129,N_6806);
and U8702 (N_8702,N_6971,N_7068);
nor U8703 (N_8703,N_7611,N_7177);
nor U8704 (N_8704,N_6931,N_6645);
and U8705 (N_8705,N_6742,N_6447);
nor U8706 (N_8706,N_6149,N_7823);
nor U8707 (N_8707,N_7036,N_6930);
nand U8708 (N_8708,N_6544,N_7324);
or U8709 (N_8709,N_7784,N_7077);
or U8710 (N_8710,N_6180,N_6145);
or U8711 (N_8711,N_7729,N_6860);
nor U8712 (N_8712,N_7910,N_7284);
nor U8713 (N_8713,N_7169,N_6684);
xor U8714 (N_8714,N_7978,N_7471);
or U8715 (N_8715,N_7731,N_6374);
and U8716 (N_8716,N_7363,N_6792);
xnor U8717 (N_8717,N_6738,N_7433);
xor U8718 (N_8718,N_6477,N_7612);
and U8719 (N_8719,N_6247,N_6414);
nor U8720 (N_8720,N_6018,N_7164);
nand U8721 (N_8721,N_6842,N_6702);
nand U8722 (N_8722,N_7542,N_7069);
and U8723 (N_8723,N_6979,N_6798);
nor U8724 (N_8724,N_6609,N_6642);
nand U8725 (N_8725,N_6574,N_7388);
xnor U8726 (N_8726,N_6888,N_7697);
or U8727 (N_8727,N_6673,N_6212);
and U8728 (N_8728,N_7165,N_6362);
xor U8729 (N_8729,N_7381,N_6775);
and U8730 (N_8730,N_7425,N_7145);
or U8731 (N_8731,N_7192,N_6852);
or U8732 (N_8732,N_7422,N_6314);
nand U8733 (N_8733,N_7184,N_7108);
nand U8734 (N_8734,N_6560,N_6187);
nand U8735 (N_8735,N_7432,N_7031);
and U8736 (N_8736,N_6122,N_6123);
nor U8737 (N_8737,N_7332,N_6906);
and U8738 (N_8738,N_7532,N_6925);
xnor U8739 (N_8739,N_6833,N_7639);
nand U8740 (N_8740,N_7569,N_6992);
nand U8741 (N_8741,N_6887,N_7277);
nand U8742 (N_8742,N_7427,N_7724);
xor U8743 (N_8743,N_6050,N_7539);
nand U8744 (N_8744,N_6696,N_6868);
nor U8745 (N_8745,N_7237,N_6918);
nor U8746 (N_8746,N_6223,N_6300);
and U8747 (N_8747,N_7742,N_7884);
and U8748 (N_8748,N_7241,N_7191);
nand U8749 (N_8749,N_6276,N_6826);
nor U8750 (N_8750,N_6882,N_7562);
or U8751 (N_8751,N_7513,N_7785);
or U8752 (N_8752,N_7752,N_7738);
and U8753 (N_8753,N_7663,N_7914);
xnor U8754 (N_8754,N_6341,N_7802);
nor U8755 (N_8755,N_7063,N_7602);
and U8756 (N_8756,N_7855,N_6137);
and U8757 (N_8757,N_6886,N_6509);
nand U8758 (N_8758,N_7948,N_7157);
or U8759 (N_8759,N_7969,N_7746);
nand U8760 (N_8760,N_7478,N_6458);
and U8761 (N_8761,N_7034,N_7900);
xnor U8762 (N_8762,N_6360,N_7550);
xor U8763 (N_8763,N_6890,N_6482);
and U8764 (N_8764,N_6699,N_6258);
nand U8765 (N_8765,N_6897,N_7636);
nor U8766 (N_8766,N_6549,N_6923);
and U8767 (N_8767,N_7558,N_7806);
and U8768 (N_8768,N_7919,N_7968);
or U8769 (N_8769,N_6337,N_6143);
nor U8770 (N_8770,N_7330,N_6151);
and U8771 (N_8771,N_7563,N_6072);
and U8772 (N_8772,N_6769,N_6739);
nand U8773 (N_8773,N_7801,N_7578);
or U8774 (N_8774,N_6831,N_7228);
and U8775 (N_8775,N_7289,N_6299);
or U8776 (N_8776,N_7464,N_6562);
and U8777 (N_8777,N_7655,N_7047);
and U8778 (N_8778,N_6507,N_6269);
nand U8779 (N_8779,N_6486,N_7696);
nand U8780 (N_8780,N_7446,N_7055);
nand U8781 (N_8781,N_6327,N_7680);
nor U8782 (N_8782,N_7659,N_7265);
or U8783 (N_8783,N_7648,N_6610);
nor U8784 (N_8784,N_7136,N_6774);
and U8785 (N_8785,N_6741,N_6885);
nand U8786 (N_8786,N_6787,N_6406);
nor U8787 (N_8787,N_7076,N_7548);
nand U8788 (N_8788,N_6495,N_6802);
xor U8789 (N_8789,N_7489,N_6023);
xor U8790 (N_8790,N_7970,N_7957);
and U8791 (N_8791,N_7294,N_7989);
nor U8792 (N_8792,N_7062,N_7350);
nor U8793 (N_8793,N_6306,N_7059);
nor U8794 (N_8794,N_7764,N_7840);
nand U8795 (N_8795,N_6464,N_6225);
nand U8796 (N_8796,N_6428,N_7740);
and U8797 (N_8797,N_7932,N_7960);
xnor U8798 (N_8798,N_7520,N_6063);
xnor U8799 (N_8799,N_7078,N_7214);
xor U8800 (N_8800,N_6440,N_7866);
nor U8801 (N_8801,N_7085,N_6772);
and U8802 (N_8802,N_6840,N_6869);
xor U8803 (N_8803,N_7111,N_7800);
and U8804 (N_8804,N_6999,N_7647);
nand U8805 (N_8805,N_7456,N_6633);
nor U8806 (N_8806,N_7374,N_6605);
and U8807 (N_8807,N_6090,N_7443);
and U8808 (N_8808,N_6138,N_6956);
nor U8809 (N_8809,N_7428,N_6668);
nor U8810 (N_8810,N_7150,N_6011);
xnor U8811 (N_8811,N_7387,N_6828);
xnor U8812 (N_8812,N_7707,N_6929);
xor U8813 (N_8813,N_6518,N_6540);
and U8814 (N_8814,N_7267,N_7906);
nand U8815 (N_8815,N_7148,N_7274);
and U8816 (N_8816,N_6856,N_6827);
and U8817 (N_8817,N_7788,N_6526);
xnor U8818 (N_8818,N_6926,N_7091);
nand U8819 (N_8819,N_6438,N_6594);
nand U8820 (N_8820,N_6163,N_6453);
xor U8821 (N_8821,N_7408,N_7492);
nand U8822 (N_8822,N_6914,N_7054);
nor U8823 (N_8823,N_7240,N_6982);
or U8824 (N_8824,N_7385,N_6911);
nor U8825 (N_8825,N_6064,N_6286);
nand U8826 (N_8826,N_6876,N_7828);
and U8827 (N_8827,N_7403,N_7426);
xnor U8828 (N_8828,N_6095,N_7041);
nor U8829 (N_8829,N_6419,N_6184);
or U8830 (N_8830,N_6884,N_7262);
nor U8831 (N_8831,N_7750,N_6995);
and U8832 (N_8832,N_6759,N_6042);
and U8833 (N_8833,N_7016,N_6510);
and U8834 (N_8834,N_7857,N_7941);
or U8835 (N_8835,N_6590,N_7279);
nand U8836 (N_8836,N_7358,N_6111);
nor U8837 (N_8837,N_6205,N_7834);
and U8838 (N_8838,N_6045,N_7251);
xnor U8839 (N_8839,N_6130,N_6086);
or U8840 (N_8840,N_6424,N_7046);
and U8841 (N_8841,N_7120,N_6913);
nand U8842 (N_8842,N_6002,N_7547);
nand U8843 (N_8843,N_7459,N_6801);
or U8844 (N_8844,N_7316,N_7633);
and U8845 (N_8845,N_7727,N_7629);
nor U8846 (N_8846,N_7365,N_6326);
nand U8847 (N_8847,N_7733,N_7907);
or U8848 (N_8848,N_6579,N_6077);
xnor U8849 (N_8849,N_6660,N_6545);
nor U8850 (N_8850,N_7911,N_7253);
nand U8851 (N_8851,N_7418,N_7212);
xnor U8852 (N_8852,N_7597,N_6656);
xor U8853 (N_8853,N_7202,N_7977);
nand U8854 (N_8854,N_7506,N_6153);
or U8855 (N_8855,N_7132,N_6907);
xor U8856 (N_8856,N_6434,N_7768);
xor U8857 (N_8857,N_6577,N_6665);
nand U8858 (N_8858,N_7346,N_6089);
xor U8859 (N_8859,N_7419,N_7992);
nand U8860 (N_8860,N_7453,N_6469);
and U8861 (N_8861,N_6272,N_7413);
and U8862 (N_8862,N_7402,N_6844);
xnor U8863 (N_8863,N_6658,N_7302);
xnor U8864 (N_8864,N_6653,N_6746);
xor U8865 (N_8865,N_7027,N_7093);
nand U8866 (N_8866,N_6519,N_7014);
xor U8867 (N_8867,N_7924,N_6229);
and U8868 (N_8868,N_7361,N_6576);
or U8869 (N_8869,N_7935,N_6899);
xnor U8870 (N_8870,N_7936,N_6566);
nor U8871 (N_8871,N_7931,N_6197);
nor U8872 (N_8872,N_7305,N_7534);
or U8873 (N_8873,N_7621,N_7073);
nor U8874 (N_8874,N_7540,N_7678);
nand U8875 (N_8875,N_6055,N_6921);
nor U8876 (N_8876,N_7842,N_7839);
or U8877 (N_8877,N_6324,N_7725);
or U8878 (N_8878,N_7321,N_7794);
nor U8879 (N_8879,N_6030,N_7658);
xor U8880 (N_8880,N_7019,N_7205);
and U8881 (N_8881,N_6537,N_6032);
nor U8882 (N_8882,N_6207,N_6241);
and U8883 (N_8883,N_7808,N_6103);
or U8884 (N_8884,N_6411,N_7883);
and U8885 (N_8885,N_7189,N_7224);
xor U8886 (N_8886,N_6076,N_6762);
nor U8887 (N_8887,N_7416,N_6053);
nand U8888 (N_8888,N_7323,N_7049);
or U8889 (N_8889,N_6632,N_6714);
nor U8890 (N_8890,N_7649,N_6483);
nor U8891 (N_8891,N_6417,N_7272);
or U8892 (N_8892,N_7035,N_7369);
nor U8893 (N_8893,N_7964,N_6960);
nand U8894 (N_8894,N_6557,N_6175);
or U8895 (N_8895,N_7771,N_7509);
nand U8896 (N_8896,N_7862,N_7870);
xor U8897 (N_8897,N_6202,N_6941);
xor U8898 (N_8898,N_6158,N_7530);
nand U8899 (N_8899,N_6808,N_7601);
or U8900 (N_8900,N_6020,N_6506);
nand U8901 (N_8901,N_7665,N_7415);
nor U8902 (N_8902,N_6644,N_6389);
nor U8903 (N_8903,N_7798,N_7296);
or U8904 (N_8904,N_7736,N_6291);
nor U8905 (N_8905,N_7546,N_6253);
nand U8906 (N_8906,N_6239,N_6625);
or U8907 (N_8907,N_6667,N_7420);
xnor U8908 (N_8908,N_6410,N_7996);
nor U8909 (N_8909,N_6094,N_6017);
nand U8910 (N_8910,N_7703,N_6813);
or U8911 (N_8911,N_6770,N_7584);
xor U8912 (N_8912,N_6303,N_7641);
xnor U8913 (N_8913,N_6079,N_7320);
nand U8914 (N_8914,N_6456,N_7566);
nand U8915 (N_8915,N_7229,N_7485);
xor U8916 (N_8916,N_6041,N_6429);
nand U8917 (N_8917,N_6485,N_6463);
or U8918 (N_8918,N_6727,N_6221);
nor U8919 (N_8919,N_6515,N_7206);
nor U8920 (N_8920,N_6088,N_6166);
xor U8921 (N_8921,N_6734,N_6669);
xor U8922 (N_8922,N_7695,N_6432);
or U8923 (N_8923,N_7245,N_7180);
xnor U8924 (N_8924,N_7384,N_7892);
and U8925 (N_8925,N_6062,N_7364);
and U8926 (N_8926,N_7503,N_6592);
and U8927 (N_8927,N_6416,N_7395);
nor U8928 (N_8928,N_6012,N_6513);
or U8929 (N_8929,N_6226,N_7341);
nor U8930 (N_8930,N_6883,N_7260);
or U8931 (N_8931,N_7730,N_7195);
nor U8932 (N_8932,N_7787,N_7376);
and U8933 (N_8933,N_6265,N_6238);
or U8934 (N_8934,N_6214,N_6274);
or U8935 (N_8935,N_6623,N_6670);
nor U8936 (N_8936,N_7692,N_7758);
nand U8937 (N_8937,N_6944,N_7890);
nand U8938 (N_8938,N_7080,N_7514);
nor U8939 (N_8939,N_6080,N_6584);
nand U8940 (N_8940,N_6900,N_7599);
nor U8941 (N_8941,N_6248,N_7770);
nand U8942 (N_8942,N_6408,N_7972);
and U8943 (N_8943,N_6864,N_6993);
or U8944 (N_8944,N_7962,N_7748);
nand U8945 (N_8945,N_7058,N_7141);
nor U8946 (N_8946,N_6799,N_6595);
or U8947 (N_8947,N_7899,N_7872);
xnor U8948 (N_8948,N_6427,N_7326);
or U8949 (N_8949,N_6522,N_6243);
and U8950 (N_8950,N_7821,N_7405);
xor U8951 (N_8951,N_7587,N_6171);
nor U8952 (N_8952,N_6983,N_6338);
or U8953 (N_8953,N_6271,N_7151);
xnor U8954 (N_8954,N_6391,N_6550);
or U8955 (N_8955,N_6346,N_7236);
and U8956 (N_8956,N_7335,N_6199);
xor U8957 (N_8957,N_7928,N_6494);
or U8958 (N_8958,N_7333,N_6331);
and U8959 (N_8959,N_7181,N_6357);
or U8960 (N_8960,N_6150,N_6358);
xnor U8961 (N_8961,N_7128,N_7543);
nand U8962 (N_8962,N_7172,N_6947);
nand U8963 (N_8963,N_6936,N_7576);
nand U8964 (N_8964,N_7102,N_7845);
nand U8965 (N_8965,N_6078,N_7545);
nor U8966 (N_8966,N_6256,N_7585);
xor U8967 (N_8967,N_6059,N_7690);
or U8968 (N_8968,N_7983,N_6192);
nor U8969 (N_8969,N_7124,N_6996);
nor U8970 (N_8970,N_7538,N_6834);
or U8971 (N_8971,N_6209,N_7480);
xnor U8972 (N_8972,N_7300,N_7504);
or U8973 (N_8973,N_7955,N_6556);
and U8974 (N_8974,N_6169,N_6606);
xor U8975 (N_8975,N_7837,N_7337);
nand U8976 (N_8976,N_6976,N_7552);
nor U8977 (N_8977,N_6087,N_7951);
and U8978 (N_8978,N_7095,N_6679);
nor U8979 (N_8979,N_7264,N_7865);
nand U8980 (N_8980,N_6972,N_6280);
nor U8981 (N_8981,N_6511,N_6879);
nor U8982 (N_8982,N_7377,N_7079);
xor U8983 (N_8983,N_6342,N_6838);
nand U8984 (N_8984,N_7675,N_6836);
nand U8985 (N_8985,N_6719,N_6777);
and U8986 (N_8986,N_7902,N_6585);
or U8987 (N_8987,N_6514,N_6386);
xor U8988 (N_8988,N_6301,N_7577);
or U8989 (N_8989,N_7194,N_7221);
xor U8990 (N_8990,N_7615,N_7760);
nand U8991 (N_8991,N_7360,N_7213);
and U8992 (N_8992,N_6422,N_6043);
nor U8993 (N_8993,N_7075,N_6877);
xnor U8994 (N_8994,N_7567,N_6587);
nor U8995 (N_8995,N_7876,N_6697);
xor U8996 (N_8996,N_6097,N_7990);
nand U8997 (N_8997,N_6098,N_7042);
xnor U8998 (N_8998,N_6334,N_6133);
and U8999 (N_8999,N_6612,N_7796);
nor U9000 (N_9000,N_6541,N_6178);
xor U9001 (N_9001,N_7269,N_6925);
nand U9002 (N_9002,N_6994,N_6862);
and U9003 (N_9003,N_6833,N_7611);
nor U9004 (N_9004,N_6852,N_6872);
and U9005 (N_9005,N_7719,N_6483);
or U9006 (N_9006,N_6452,N_7191);
nand U9007 (N_9007,N_6394,N_6432);
nor U9008 (N_9008,N_7439,N_6724);
nor U9009 (N_9009,N_7624,N_7135);
nand U9010 (N_9010,N_6922,N_7080);
nor U9011 (N_9011,N_7519,N_6454);
nor U9012 (N_9012,N_7862,N_6652);
and U9013 (N_9013,N_7257,N_7732);
nand U9014 (N_9014,N_6337,N_7576);
and U9015 (N_9015,N_6726,N_7209);
or U9016 (N_9016,N_7091,N_6178);
or U9017 (N_9017,N_6637,N_6707);
or U9018 (N_9018,N_7991,N_7172);
nand U9019 (N_9019,N_6065,N_7989);
and U9020 (N_9020,N_7724,N_6985);
nand U9021 (N_9021,N_6264,N_6500);
xor U9022 (N_9022,N_6603,N_7946);
and U9023 (N_9023,N_6382,N_6957);
xor U9024 (N_9024,N_6272,N_7497);
xnor U9025 (N_9025,N_6072,N_6618);
xnor U9026 (N_9026,N_6613,N_7085);
nor U9027 (N_9027,N_6936,N_6101);
or U9028 (N_9028,N_6730,N_6171);
nand U9029 (N_9029,N_7484,N_6424);
nor U9030 (N_9030,N_7008,N_7639);
nand U9031 (N_9031,N_7872,N_7485);
nand U9032 (N_9032,N_6421,N_7364);
xor U9033 (N_9033,N_6695,N_6884);
nand U9034 (N_9034,N_6030,N_6524);
nor U9035 (N_9035,N_7778,N_7098);
nor U9036 (N_9036,N_6886,N_6358);
xor U9037 (N_9037,N_6307,N_7321);
nand U9038 (N_9038,N_7804,N_7602);
and U9039 (N_9039,N_6971,N_7103);
xnor U9040 (N_9040,N_7496,N_7195);
xnor U9041 (N_9041,N_6246,N_7241);
xnor U9042 (N_9042,N_7088,N_7696);
nor U9043 (N_9043,N_7175,N_6468);
or U9044 (N_9044,N_7845,N_7447);
nand U9045 (N_9045,N_7749,N_7034);
or U9046 (N_9046,N_6203,N_6110);
and U9047 (N_9047,N_6409,N_6964);
nor U9048 (N_9048,N_6182,N_6837);
and U9049 (N_9049,N_7192,N_7004);
or U9050 (N_9050,N_6065,N_6546);
and U9051 (N_9051,N_6440,N_6792);
or U9052 (N_9052,N_6618,N_7895);
or U9053 (N_9053,N_6923,N_7747);
nand U9054 (N_9054,N_6397,N_6861);
or U9055 (N_9055,N_7834,N_6701);
and U9056 (N_9056,N_6526,N_6174);
nand U9057 (N_9057,N_7041,N_7681);
nor U9058 (N_9058,N_7576,N_7683);
and U9059 (N_9059,N_6414,N_6202);
xnor U9060 (N_9060,N_6418,N_6427);
xnor U9061 (N_9061,N_6610,N_7953);
xor U9062 (N_9062,N_7951,N_7250);
or U9063 (N_9063,N_7226,N_6776);
and U9064 (N_9064,N_6764,N_6261);
and U9065 (N_9065,N_7184,N_7573);
nand U9066 (N_9066,N_6805,N_7758);
and U9067 (N_9067,N_6346,N_7407);
nand U9068 (N_9068,N_6040,N_6320);
or U9069 (N_9069,N_6855,N_6017);
xnor U9070 (N_9070,N_6137,N_6306);
and U9071 (N_9071,N_7810,N_7337);
xor U9072 (N_9072,N_7158,N_6556);
or U9073 (N_9073,N_7610,N_6187);
nand U9074 (N_9074,N_6066,N_6007);
nand U9075 (N_9075,N_7579,N_6298);
nor U9076 (N_9076,N_6757,N_6790);
and U9077 (N_9077,N_6480,N_6697);
xor U9078 (N_9078,N_6377,N_6418);
nor U9079 (N_9079,N_7962,N_6356);
xnor U9080 (N_9080,N_6265,N_7489);
or U9081 (N_9081,N_7430,N_6813);
nor U9082 (N_9082,N_6112,N_7032);
nand U9083 (N_9083,N_7889,N_6835);
nor U9084 (N_9084,N_7300,N_7762);
and U9085 (N_9085,N_7734,N_6992);
xnor U9086 (N_9086,N_7747,N_6303);
nor U9087 (N_9087,N_7667,N_6698);
and U9088 (N_9088,N_6979,N_6397);
nand U9089 (N_9089,N_6661,N_7325);
or U9090 (N_9090,N_6589,N_6600);
and U9091 (N_9091,N_6038,N_7529);
nand U9092 (N_9092,N_6243,N_6723);
or U9093 (N_9093,N_7492,N_7838);
and U9094 (N_9094,N_7418,N_6554);
and U9095 (N_9095,N_6776,N_6182);
xnor U9096 (N_9096,N_7663,N_7279);
nand U9097 (N_9097,N_7512,N_7264);
and U9098 (N_9098,N_6666,N_7131);
and U9099 (N_9099,N_7699,N_7706);
nand U9100 (N_9100,N_6442,N_7321);
nand U9101 (N_9101,N_6412,N_6152);
or U9102 (N_9102,N_7053,N_7623);
or U9103 (N_9103,N_7841,N_7681);
and U9104 (N_9104,N_6609,N_7220);
xor U9105 (N_9105,N_6700,N_6119);
or U9106 (N_9106,N_6841,N_6474);
xnor U9107 (N_9107,N_6098,N_7769);
xor U9108 (N_9108,N_6538,N_6436);
nand U9109 (N_9109,N_7175,N_7771);
and U9110 (N_9110,N_6020,N_6272);
and U9111 (N_9111,N_7827,N_6698);
nand U9112 (N_9112,N_7934,N_6419);
and U9113 (N_9113,N_7959,N_7718);
xnor U9114 (N_9114,N_7043,N_7130);
or U9115 (N_9115,N_6935,N_7344);
and U9116 (N_9116,N_6761,N_6051);
xnor U9117 (N_9117,N_7814,N_6463);
xor U9118 (N_9118,N_7714,N_7336);
xnor U9119 (N_9119,N_6109,N_6665);
nor U9120 (N_9120,N_6396,N_7713);
and U9121 (N_9121,N_6398,N_7761);
xnor U9122 (N_9122,N_7027,N_6993);
nand U9123 (N_9123,N_7797,N_7444);
xnor U9124 (N_9124,N_6002,N_7258);
xor U9125 (N_9125,N_6855,N_6065);
or U9126 (N_9126,N_7608,N_7017);
and U9127 (N_9127,N_6743,N_6739);
and U9128 (N_9128,N_7763,N_6749);
or U9129 (N_9129,N_6549,N_7284);
nor U9130 (N_9130,N_7958,N_7289);
nand U9131 (N_9131,N_7454,N_6172);
and U9132 (N_9132,N_7639,N_6628);
or U9133 (N_9133,N_6216,N_6135);
or U9134 (N_9134,N_7818,N_7044);
xnor U9135 (N_9135,N_6157,N_6992);
and U9136 (N_9136,N_6479,N_6369);
nor U9137 (N_9137,N_7921,N_6339);
xnor U9138 (N_9138,N_6104,N_6755);
nor U9139 (N_9139,N_7046,N_6677);
nand U9140 (N_9140,N_7684,N_6080);
xor U9141 (N_9141,N_7447,N_7015);
or U9142 (N_9142,N_6378,N_7484);
and U9143 (N_9143,N_6793,N_6392);
or U9144 (N_9144,N_6880,N_7672);
nand U9145 (N_9145,N_6494,N_7057);
nor U9146 (N_9146,N_7796,N_6933);
nand U9147 (N_9147,N_6417,N_7999);
nor U9148 (N_9148,N_7079,N_6276);
or U9149 (N_9149,N_7499,N_6117);
nand U9150 (N_9150,N_6095,N_6850);
nor U9151 (N_9151,N_6963,N_6662);
or U9152 (N_9152,N_7666,N_6540);
xor U9153 (N_9153,N_6918,N_7576);
nor U9154 (N_9154,N_7152,N_7587);
nand U9155 (N_9155,N_6966,N_6093);
or U9156 (N_9156,N_6829,N_6173);
nor U9157 (N_9157,N_6546,N_6230);
nor U9158 (N_9158,N_7312,N_7083);
or U9159 (N_9159,N_7309,N_7580);
and U9160 (N_9160,N_7986,N_6813);
xnor U9161 (N_9161,N_7747,N_7090);
nor U9162 (N_9162,N_7767,N_6026);
nand U9163 (N_9163,N_7666,N_7279);
and U9164 (N_9164,N_7637,N_6278);
nor U9165 (N_9165,N_7373,N_6130);
nand U9166 (N_9166,N_6035,N_7591);
and U9167 (N_9167,N_7908,N_6774);
and U9168 (N_9168,N_6638,N_6249);
or U9169 (N_9169,N_7327,N_7621);
or U9170 (N_9170,N_7811,N_6842);
nand U9171 (N_9171,N_7032,N_7367);
xnor U9172 (N_9172,N_7439,N_7203);
or U9173 (N_9173,N_6478,N_6823);
nand U9174 (N_9174,N_7019,N_7976);
nand U9175 (N_9175,N_6647,N_7000);
nor U9176 (N_9176,N_6423,N_6311);
and U9177 (N_9177,N_6237,N_6990);
nor U9178 (N_9178,N_7936,N_6854);
or U9179 (N_9179,N_7907,N_7621);
xnor U9180 (N_9180,N_7995,N_6442);
or U9181 (N_9181,N_6081,N_7631);
xor U9182 (N_9182,N_6962,N_7339);
xor U9183 (N_9183,N_7806,N_7715);
nor U9184 (N_9184,N_6842,N_7331);
nor U9185 (N_9185,N_6762,N_6952);
or U9186 (N_9186,N_7304,N_6756);
and U9187 (N_9187,N_7391,N_6367);
or U9188 (N_9188,N_7594,N_6072);
xnor U9189 (N_9189,N_7625,N_6561);
nand U9190 (N_9190,N_6394,N_7696);
nand U9191 (N_9191,N_6550,N_7704);
xor U9192 (N_9192,N_7648,N_7736);
nor U9193 (N_9193,N_6082,N_7153);
xnor U9194 (N_9194,N_6227,N_6248);
and U9195 (N_9195,N_6047,N_7111);
xnor U9196 (N_9196,N_7432,N_7122);
nor U9197 (N_9197,N_7260,N_6484);
nand U9198 (N_9198,N_6034,N_7055);
nand U9199 (N_9199,N_7389,N_6646);
and U9200 (N_9200,N_6376,N_7883);
or U9201 (N_9201,N_7478,N_6133);
nor U9202 (N_9202,N_6327,N_7601);
and U9203 (N_9203,N_6013,N_7839);
nor U9204 (N_9204,N_6216,N_6087);
nor U9205 (N_9205,N_7476,N_6674);
xor U9206 (N_9206,N_7369,N_7226);
nand U9207 (N_9207,N_7752,N_7188);
xnor U9208 (N_9208,N_6077,N_7843);
or U9209 (N_9209,N_6375,N_7400);
nor U9210 (N_9210,N_6170,N_6674);
nor U9211 (N_9211,N_6937,N_7295);
nand U9212 (N_9212,N_6463,N_7946);
or U9213 (N_9213,N_6669,N_6232);
and U9214 (N_9214,N_6705,N_7328);
and U9215 (N_9215,N_6103,N_7241);
and U9216 (N_9216,N_7118,N_7162);
xor U9217 (N_9217,N_7455,N_6881);
xnor U9218 (N_9218,N_7770,N_6923);
and U9219 (N_9219,N_6476,N_6228);
xor U9220 (N_9220,N_6112,N_7957);
nand U9221 (N_9221,N_6225,N_7404);
or U9222 (N_9222,N_6903,N_6469);
or U9223 (N_9223,N_7508,N_6267);
nor U9224 (N_9224,N_7932,N_6230);
and U9225 (N_9225,N_6495,N_7177);
nand U9226 (N_9226,N_7138,N_7692);
or U9227 (N_9227,N_7338,N_7997);
xnor U9228 (N_9228,N_7336,N_7306);
and U9229 (N_9229,N_6442,N_6951);
and U9230 (N_9230,N_7555,N_7282);
or U9231 (N_9231,N_7546,N_6313);
nand U9232 (N_9232,N_7666,N_7880);
or U9233 (N_9233,N_6884,N_7618);
nand U9234 (N_9234,N_6538,N_6867);
nand U9235 (N_9235,N_6144,N_7213);
and U9236 (N_9236,N_6881,N_7735);
nand U9237 (N_9237,N_6564,N_7732);
and U9238 (N_9238,N_6146,N_6754);
xor U9239 (N_9239,N_6274,N_7320);
and U9240 (N_9240,N_7477,N_7540);
nor U9241 (N_9241,N_6055,N_7806);
nand U9242 (N_9242,N_7301,N_6101);
or U9243 (N_9243,N_6064,N_6334);
nand U9244 (N_9244,N_6864,N_7785);
nor U9245 (N_9245,N_7368,N_7458);
or U9246 (N_9246,N_7362,N_7000);
xor U9247 (N_9247,N_6867,N_7708);
nor U9248 (N_9248,N_6948,N_7390);
nor U9249 (N_9249,N_6940,N_6423);
and U9250 (N_9250,N_7062,N_7701);
or U9251 (N_9251,N_7609,N_7328);
and U9252 (N_9252,N_7355,N_6034);
and U9253 (N_9253,N_6233,N_7255);
xnor U9254 (N_9254,N_6114,N_7837);
nand U9255 (N_9255,N_7677,N_7162);
and U9256 (N_9256,N_6603,N_6633);
or U9257 (N_9257,N_6869,N_6224);
nor U9258 (N_9258,N_6362,N_6320);
or U9259 (N_9259,N_6560,N_7637);
nor U9260 (N_9260,N_6758,N_7457);
and U9261 (N_9261,N_6283,N_6617);
or U9262 (N_9262,N_7941,N_6869);
or U9263 (N_9263,N_7239,N_7865);
xnor U9264 (N_9264,N_7244,N_7097);
nor U9265 (N_9265,N_6245,N_6402);
nand U9266 (N_9266,N_6187,N_7408);
xnor U9267 (N_9267,N_7013,N_7437);
xnor U9268 (N_9268,N_6871,N_7834);
and U9269 (N_9269,N_6561,N_7817);
or U9270 (N_9270,N_7768,N_6703);
nor U9271 (N_9271,N_6441,N_6024);
or U9272 (N_9272,N_6908,N_6400);
nand U9273 (N_9273,N_6884,N_7233);
and U9274 (N_9274,N_7482,N_7177);
xnor U9275 (N_9275,N_7647,N_7296);
nand U9276 (N_9276,N_7691,N_7166);
xor U9277 (N_9277,N_7116,N_7375);
and U9278 (N_9278,N_6785,N_6919);
nand U9279 (N_9279,N_7268,N_7288);
and U9280 (N_9280,N_7141,N_7087);
nand U9281 (N_9281,N_7415,N_6665);
or U9282 (N_9282,N_6355,N_7069);
or U9283 (N_9283,N_7539,N_7429);
nand U9284 (N_9284,N_7430,N_7833);
nand U9285 (N_9285,N_7403,N_6166);
nand U9286 (N_9286,N_7961,N_6987);
or U9287 (N_9287,N_6974,N_7844);
and U9288 (N_9288,N_7804,N_7690);
and U9289 (N_9289,N_7829,N_7184);
or U9290 (N_9290,N_6796,N_6513);
xor U9291 (N_9291,N_7846,N_7593);
xor U9292 (N_9292,N_7323,N_6433);
xnor U9293 (N_9293,N_6260,N_7101);
and U9294 (N_9294,N_7318,N_6600);
nor U9295 (N_9295,N_7087,N_7491);
nor U9296 (N_9296,N_7444,N_7146);
nor U9297 (N_9297,N_7147,N_6818);
nand U9298 (N_9298,N_7907,N_7161);
and U9299 (N_9299,N_6922,N_6992);
xor U9300 (N_9300,N_6599,N_6213);
nor U9301 (N_9301,N_7188,N_6941);
and U9302 (N_9302,N_6083,N_7249);
or U9303 (N_9303,N_7133,N_7501);
nand U9304 (N_9304,N_7979,N_6466);
and U9305 (N_9305,N_7734,N_6372);
and U9306 (N_9306,N_6298,N_6481);
and U9307 (N_9307,N_7967,N_6884);
nor U9308 (N_9308,N_6081,N_6565);
or U9309 (N_9309,N_6930,N_7311);
nor U9310 (N_9310,N_7357,N_7955);
and U9311 (N_9311,N_7911,N_6779);
nand U9312 (N_9312,N_7359,N_6065);
and U9313 (N_9313,N_6612,N_7742);
and U9314 (N_9314,N_7149,N_6078);
or U9315 (N_9315,N_6987,N_7288);
or U9316 (N_9316,N_7615,N_7126);
and U9317 (N_9317,N_7362,N_6607);
xor U9318 (N_9318,N_7850,N_7348);
xor U9319 (N_9319,N_6899,N_6151);
and U9320 (N_9320,N_6488,N_7134);
or U9321 (N_9321,N_7797,N_7945);
nand U9322 (N_9322,N_7039,N_6950);
or U9323 (N_9323,N_7034,N_6582);
nor U9324 (N_9324,N_6067,N_6454);
nand U9325 (N_9325,N_6355,N_7715);
nand U9326 (N_9326,N_7716,N_6150);
nor U9327 (N_9327,N_6345,N_7835);
xor U9328 (N_9328,N_7902,N_7702);
xor U9329 (N_9329,N_6019,N_6307);
nor U9330 (N_9330,N_7281,N_7720);
or U9331 (N_9331,N_7152,N_6405);
or U9332 (N_9332,N_7195,N_6360);
nand U9333 (N_9333,N_6424,N_7728);
nor U9334 (N_9334,N_6490,N_6139);
nand U9335 (N_9335,N_6670,N_7878);
xnor U9336 (N_9336,N_6808,N_7822);
nand U9337 (N_9337,N_7353,N_7617);
or U9338 (N_9338,N_6520,N_6223);
and U9339 (N_9339,N_7458,N_6931);
xnor U9340 (N_9340,N_6657,N_7060);
nand U9341 (N_9341,N_7125,N_7331);
nand U9342 (N_9342,N_7573,N_6323);
and U9343 (N_9343,N_7880,N_7595);
xnor U9344 (N_9344,N_6645,N_7786);
nand U9345 (N_9345,N_7303,N_7889);
or U9346 (N_9346,N_7031,N_7959);
xor U9347 (N_9347,N_6661,N_6972);
or U9348 (N_9348,N_7138,N_7678);
nor U9349 (N_9349,N_7677,N_6537);
or U9350 (N_9350,N_7336,N_7068);
xnor U9351 (N_9351,N_6795,N_6707);
xor U9352 (N_9352,N_6075,N_6121);
and U9353 (N_9353,N_7615,N_7948);
and U9354 (N_9354,N_6116,N_6381);
xor U9355 (N_9355,N_6883,N_6730);
xor U9356 (N_9356,N_6008,N_6852);
and U9357 (N_9357,N_7702,N_6907);
nand U9358 (N_9358,N_6282,N_7163);
nand U9359 (N_9359,N_6034,N_6669);
and U9360 (N_9360,N_6854,N_6610);
xnor U9361 (N_9361,N_7167,N_6201);
nor U9362 (N_9362,N_6739,N_7889);
nor U9363 (N_9363,N_7069,N_6316);
and U9364 (N_9364,N_7875,N_7482);
xor U9365 (N_9365,N_7883,N_7585);
nor U9366 (N_9366,N_7718,N_6245);
nor U9367 (N_9367,N_6958,N_6650);
or U9368 (N_9368,N_7392,N_6849);
or U9369 (N_9369,N_7860,N_6779);
nand U9370 (N_9370,N_7997,N_6364);
xnor U9371 (N_9371,N_6830,N_6275);
nor U9372 (N_9372,N_6762,N_6379);
xnor U9373 (N_9373,N_6914,N_7245);
and U9374 (N_9374,N_7740,N_7862);
and U9375 (N_9375,N_7661,N_6024);
nor U9376 (N_9376,N_6305,N_7298);
or U9377 (N_9377,N_7015,N_6212);
or U9378 (N_9378,N_6002,N_6071);
nand U9379 (N_9379,N_6540,N_7556);
nor U9380 (N_9380,N_7380,N_7518);
nand U9381 (N_9381,N_6863,N_7372);
and U9382 (N_9382,N_6592,N_6580);
xnor U9383 (N_9383,N_6997,N_7762);
or U9384 (N_9384,N_6312,N_7185);
and U9385 (N_9385,N_6712,N_6346);
and U9386 (N_9386,N_6351,N_7110);
nor U9387 (N_9387,N_6537,N_6285);
nand U9388 (N_9388,N_6201,N_6034);
or U9389 (N_9389,N_7063,N_6177);
or U9390 (N_9390,N_6942,N_7373);
or U9391 (N_9391,N_7601,N_6712);
nor U9392 (N_9392,N_6551,N_7343);
and U9393 (N_9393,N_6370,N_6317);
nand U9394 (N_9394,N_6851,N_7465);
or U9395 (N_9395,N_6057,N_7529);
nand U9396 (N_9396,N_7668,N_7374);
nand U9397 (N_9397,N_7817,N_7759);
xnor U9398 (N_9398,N_6112,N_7866);
nor U9399 (N_9399,N_6217,N_7549);
xnor U9400 (N_9400,N_6741,N_7974);
nand U9401 (N_9401,N_7478,N_6318);
xnor U9402 (N_9402,N_7000,N_7778);
xor U9403 (N_9403,N_6670,N_7020);
nand U9404 (N_9404,N_7885,N_7629);
xor U9405 (N_9405,N_7336,N_7490);
and U9406 (N_9406,N_6271,N_7451);
or U9407 (N_9407,N_7753,N_7542);
nor U9408 (N_9408,N_7964,N_6669);
nor U9409 (N_9409,N_7067,N_7925);
xor U9410 (N_9410,N_6714,N_6627);
xor U9411 (N_9411,N_7849,N_7961);
nor U9412 (N_9412,N_7704,N_6882);
and U9413 (N_9413,N_6467,N_6408);
or U9414 (N_9414,N_7174,N_7337);
and U9415 (N_9415,N_7359,N_7989);
or U9416 (N_9416,N_6951,N_7455);
nand U9417 (N_9417,N_7394,N_7815);
or U9418 (N_9418,N_6571,N_6934);
and U9419 (N_9419,N_7313,N_7764);
and U9420 (N_9420,N_7676,N_6636);
or U9421 (N_9421,N_7480,N_6121);
nor U9422 (N_9422,N_6637,N_7635);
and U9423 (N_9423,N_6258,N_6019);
or U9424 (N_9424,N_6709,N_6759);
or U9425 (N_9425,N_6792,N_6480);
nor U9426 (N_9426,N_6376,N_7828);
nor U9427 (N_9427,N_6610,N_7634);
and U9428 (N_9428,N_6727,N_7483);
nand U9429 (N_9429,N_6912,N_7683);
nor U9430 (N_9430,N_7931,N_7259);
nor U9431 (N_9431,N_7760,N_6282);
nand U9432 (N_9432,N_6675,N_6710);
and U9433 (N_9433,N_6407,N_6548);
nand U9434 (N_9434,N_7538,N_7595);
and U9435 (N_9435,N_7548,N_7702);
and U9436 (N_9436,N_6191,N_6719);
xnor U9437 (N_9437,N_7932,N_6358);
xor U9438 (N_9438,N_7104,N_6935);
nand U9439 (N_9439,N_7156,N_7179);
nand U9440 (N_9440,N_6398,N_6042);
nand U9441 (N_9441,N_6475,N_7529);
and U9442 (N_9442,N_6902,N_6230);
or U9443 (N_9443,N_7918,N_6918);
and U9444 (N_9444,N_6378,N_6996);
and U9445 (N_9445,N_6982,N_7156);
xor U9446 (N_9446,N_7855,N_6178);
or U9447 (N_9447,N_6897,N_6390);
and U9448 (N_9448,N_7429,N_7499);
or U9449 (N_9449,N_7195,N_7207);
or U9450 (N_9450,N_7624,N_6800);
nand U9451 (N_9451,N_6362,N_6702);
xor U9452 (N_9452,N_6107,N_7442);
or U9453 (N_9453,N_6217,N_6125);
and U9454 (N_9454,N_6589,N_7535);
nand U9455 (N_9455,N_6296,N_6796);
and U9456 (N_9456,N_6516,N_6499);
or U9457 (N_9457,N_6047,N_6234);
nand U9458 (N_9458,N_6730,N_7924);
nand U9459 (N_9459,N_6710,N_6313);
and U9460 (N_9460,N_6718,N_7790);
nor U9461 (N_9461,N_6584,N_7130);
nor U9462 (N_9462,N_6549,N_6034);
nand U9463 (N_9463,N_6343,N_7597);
and U9464 (N_9464,N_7431,N_6071);
xnor U9465 (N_9465,N_6038,N_6481);
or U9466 (N_9466,N_7088,N_6301);
or U9467 (N_9467,N_6129,N_6081);
or U9468 (N_9468,N_6934,N_6703);
nand U9469 (N_9469,N_6284,N_7007);
or U9470 (N_9470,N_6344,N_6879);
and U9471 (N_9471,N_6771,N_7912);
or U9472 (N_9472,N_6438,N_6018);
nor U9473 (N_9473,N_6386,N_7742);
or U9474 (N_9474,N_7006,N_6196);
and U9475 (N_9475,N_7853,N_7850);
and U9476 (N_9476,N_6614,N_6426);
nand U9477 (N_9477,N_6232,N_7309);
xor U9478 (N_9478,N_7177,N_7901);
or U9479 (N_9479,N_7313,N_6659);
nand U9480 (N_9480,N_6664,N_6470);
nor U9481 (N_9481,N_7509,N_7533);
and U9482 (N_9482,N_6042,N_7121);
xnor U9483 (N_9483,N_7667,N_6579);
or U9484 (N_9484,N_6214,N_7039);
xor U9485 (N_9485,N_6451,N_7712);
nand U9486 (N_9486,N_7713,N_7019);
nor U9487 (N_9487,N_7651,N_7849);
or U9488 (N_9488,N_7036,N_6144);
nor U9489 (N_9489,N_7050,N_6124);
and U9490 (N_9490,N_7513,N_7589);
and U9491 (N_9491,N_7326,N_6278);
nand U9492 (N_9492,N_7755,N_6341);
nor U9493 (N_9493,N_6565,N_6977);
or U9494 (N_9494,N_6602,N_7594);
or U9495 (N_9495,N_7028,N_7657);
or U9496 (N_9496,N_6884,N_6889);
and U9497 (N_9497,N_7674,N_7627);
nor U9498 (N_9498,N_7046,N_7236);
nand U9499 (N_9499,N_6838,N_6442);
and U9500 (N_9500,N_6945,N_6954);
xnor U9501 (N_9501,N_7111,N_7894);
and U9502 (N_9502,N_6927,N_7399);
nand U9503 (N_9503,N_7896,N_6824);
or U9504 (N_9504,N_6156,N_7547);
nand U9505 (N_9505,N_6711,N_7484);
xnor U9506 (N_9506,N_7836,N_7680);
and U9507 (N_9507,N_6977,N_6413);
nor U9508 (N_9508,N_6394,N_6644);
nor U9509 (N_9509,N_6102,N_7184);
nor U9510 (N_9510,N_6308,N_7484);
nor U9511 (N_9511,N_6841,N_7958);
nor U9512 (N_9512,N_6298,N_6901);
nand U9513 (N_9513,N_6322,N_7101);
or U9514 (N_9514,N_7802,N_7327);
or U9515 (N_9515,N_6688,N_7660);
nor U9516 (N_9516,N_7593,N_7843);
or U9517 (N_9517,N_7127,N_6306);
xor U9518 (N_9518,N_7537,N_7006);
or U9519 (N_9519,N_6746,N_6072);
xnor U9520 (N_9520,N_6622,N_6233);
nand U9521 (N_9521,N_6505,N_7255);
nand U9522 (N_9522,N_6027,N_6993);
nor U9523 (N_9523,N_6312,N_7434);
xnor U9524 (N_9524,N_7649,N_6580);
xnor U9525 (N_9525,N_6902,N_6768);
nand U9526 (N_9526,N_6157,N_7900);
nor U9527 (N_9527,N_6225,N_6457);
xor U9528 (N_9528,N_6843,N_7536);
nand U9529 (N_9529,N_7861,N_7734);
xor U9530 (N_9530,N_6914,N_7626);
nand U9531 (N_9531,N_7333,N_7496);
nand U9532 (N_9532,N_7222,N_6789);
nor U9533 (N_9533,N_6218,N_7839);
and U9534 (N_9534,N_6981,N_6086);
and U9535 (N_9535,N_7404,N_7307);
nand U9536 (N_9536,N_7681,N_6404);
xor U9537 (N_9537,N_6243,N_6834);
nand U9538 (N_9538,N_7213,N_7732);
and U9539 (N_9539,N_6400,N_6622);
nand U9540 (N_9540,N_7126,N_6667);
nor U9541 (N_9541,N_6916,N_7046);
nor U9542 (N_9542,N_6274,N_6385);
and U9543 (N_9543,N_7319,N_6166);
nor U9544 (N_9544,N_7218,N_6804);
xnor U9545 (N_9545,N_6852,N_7014);
xor U9546 (N_9546,N_6525,N_6702);
or U9547 (N_9547,N_7390,N_7832);
nor U9548 (N_9548,N_6773,N_6630);
nand U9549 (N_9549,N_6232,N_7048);
nor U9550 (N_9550,N_7736,N_7074);
nor U9551 (N_9551,N_6605,N_6977);
nor U9552 (N_9552,N_7690,N_6257);
nor U9553 (N_9553,N_7842,N_6931);
nor U9554 (N_9554,N_7703,N_7690);
nand U9555 (N_9555,N_6122,N_6252);
or U9556 (N_9556,N_6747,N_6349);
and U9557 (N_9557,N_6836,N_7810);
nor U9558 (N_9558,N_6879,N_6107);
or U9559 (N_9559,N_6887,N_7595);
or U9560 (N_9560,N_6768,N_7317);
or U9561 (N_9561,N_6177,N_6336);
or U9562 (N_9562,N_6604,N_6419);
nand U9563 (N_9563,N_6384,N_6702);
nor U9564 (N_9564,N_7382,N_7711);
nand U9565 (N_9565,N_6267,N_7877);
nor U9566 (N_9566,N_6900,N_7030);
and U9567 (N_9567,N_7186,N_7123);
nand U9568 (N_9568,N_7233,N_6813);
or U9569 (N_9569,N_6230,N_7962);
or U9570 (N_9570,N_6002,N_7371);
nor U9571 (N_9571,N_6724,N_6594);
xor U9572 (N_9572,N_7962,N_7951);
xnor U9573 (N_9573,N_7849,N_6698);
nand U9574 (N_9574,N_7920,N_7431);
nand U9575 (N_9575,N_7749,N_6925);
xnor U9576 (N_9576,N_7646,N_6096);
and U9577 (N_9577,N_6738,N_7236);
or U9578 (N_9578,N_6540,N_6453);
and U9579 (N_9579,N_6881,N_6535);
and U9580 (N_9580,N_6641,N_6953);
or U9581 (N_9581,N_6804,N_6994);
and U9582 (N_9582,N_6952,N_6049);
nand U9583 (N_9583,N_6777,N_6039);
nand U9584 (N_9584,N_7248,N_6060);
and U9585 (N_9585,N_7293,N_6554);
and U9586 (N_9586,N_7781,N_6039);
and U9587 (N_9587,N_7384,N_7649);
or U9588 (N_9588,N_6947,N_7031);
nand U9589 (N_9589,N_6175,N_7789);
and U9590 (N_9590,N_6716,N_7819);
xor U9591 (N_9591,N_7572,N_6059);
and U9592 (N_9592,N_7376,N_7427);
or U9593 (N_9593,N_7757,N_6689);
nand U9594 (N_9594,N_6743,N_6749);
xor U9595 (N_9595,N_6933,N_6635);
xor U9596 (N_9596,N_6195,N_7150);
and U9597 (N_9597,N_6567,N_6829);
nor U9598 (N_9598,N_6795,N_7192);
nand U9599 (N_9599,N_7183,N_7107);
nor U9600 (N_9600,N_7300,N_7074);
nand U9601 (N_9601,N_7703,N_6689);
and U9602 (N_9602,N_6975,N_7432);
nor U9603 (N_9603,N_6014,N_7849);
nor U9604 (N_9604,N_7147,N_6301);
nor U9605 (N_9605,N_6412,N_6999);
xnor U9606 (N_9606,N_6987,N_6730);
or U9607 (N_9607,N_6041,N_6727);
nand U9608 (N_9608,N_7339,N_6072);
nand U9609 (N_9609,N_7138,N_6860);
and U9610 (N_9610,N_6297,N_6962);
or U9611 (N_9611,N_6406,N_6732);
or U9612 (N_9612,N_6704,N_6732);
and U9613 (N_9613,N_7753,N_7133);
or U9614 (N_9614,N_7952,N_6426);
nand U9615 (N_9615,N_6440,N_6805);
nand U9616 (N_9616,N_7957,N_6709);
nand U9617 (N_9617,N_6547,N_7823);
nand U9618 (N_9618,N_6503,N_7294);
xor U9619 (N_9619,N_7642,N_6542);
nor U9620 (N_9620,N_6135,N_7109);
and U9621 (N_9621,N_7855,N_6791);
nand U9622 (N_9622,N_6990,N_6825);
or U9623 (N_9623,N_7906,N_6167);
nand U9624 (N_9624,N_7077,N_6103);
and U9625 (N_9625,N_7367,N_7905);
nor U9626 (N_9626,N_7772,N_6712);
xnor U9627 (N_9627,N_7977,N_7389);
nand U9628 (N_9628,N_7660,N_7083);
nor U9629 (N_9629,N_7580,N_7844);
and U9630 (N_9630,N_7629,N_6469);
and U9631 (N_9631,N_7130,N_6462);
or U9632 (N_9632,N_6875,N_6550);
nand U9633 (N_9633,N_6832,N_6917);
nand U9634 (N_9634,N_7473,N_7879);
nand U9635 (N_9635,N_7556,N_6092);
xnor U9636 (N_9636,N_7203,N_6930);
nand U9637 (N_9637,N_6618,N_7919);
nor U9638 (N_9638,N_6673,N_6974);
nor U9639 (N_9639,N_7329,N_6126);
xor U9640 (N_9640,N_7311,N_6624);
or U9641 (N_9641,N_7641,N_6079);
nor U9642 (N_9642,N_6779,N_7654);
or U9643 (N_9643,N_7185,N_6324);
and U9644 (N_9644,N_6339,N_7405);
nand U9645 (N_9645,N_6577,N_7023);
nor U9646 (N_9646,N_6611,N_6322);
and U9647 (N_9647,N_7749,N_7508);
nand U9648 (N_9648,N_7021,N_7542);
and U9649 (N_9649,N_6498,N_6690);
xor U9650 (N_9650,N_6738,N_6599);
nor U9651 (N_9651,N_7814,N_7872);
nor U9652 (N_9652,N_6137,N_7709);
nand U9653 (N_9653,N_7689,N_7856);
xor U9654 (N_9654,N_7410,N_6984);
nor U9655 (N_9655,N_7584,N_7394);
and U9656 (N_9656,N_6608,N_6471);
nand U9657 (N_9657,N_6195,N_6232);
or U9658 (N_9658,N_6630,N_7388);
nand U9659 (N_9659,N_6351,N_6287);
nand U9660 (N_9660,N_6664,N_6160);
nand U9661 (N_9661,N_6893,N_7556);
and U9662 (N_9662,N_6842,N_7893);
and U9663 (N_9663,N_6720,N_7874);
or U9664 (N_9664,N_6876,N_7011);
nor U9665 (N_9665,N_6797,N_7932);
or U9666 (N_9666,N_7674,N_7104);
xnor U9667 (N_9667,N_7737,N_7141);
or U9668 (N_9668,N_6866,N_6124);
nand U9669 (N_9669,N_6427,N_7933);
xor U9670 (N_9670,N_6973,N_7403);
xor U9671 (N_9671,N_6950,N_7613);
or U9672 (N_9672,N_6120,N_6566);
xor U9673 (N_9673,N_6728,N_6990);
nor U9674 (N_9674,N_6718,N_7841);
nand U9675 (N_9675,N_7991,N_6018);
nor U9676 (N_9676,N_7633,N_7991);
nor U9677 (N_9677,N_7108,N_7616);
or U9678 (N_9678,N_6133,N_6496);
nor U9679 (N_9679,N_6510,N_6709);
and U9680 (N_9680,N_6903,N_6125);
nor U9681 (N_9681,N_7488,N_6951);
xor U9682 (N_9682,N_6592,N_7424);
and U9683 (N_9683,N_6900,N_6105);
or U9684 (N_9684,N_7296,N_6680);
or U9685 (N_9685,N_6701,N_6505);
and U9686 (N_9686,N_7645,N_7327);
xor U9687 (N_9687,N_7087,N_6552);
nor U9688 (N_9688,N_6274,N_7964);
and U9689 (N_9689,N_7735,N_6815);
or U9690 (N_9690,N_6922,N_7023);
or U9691 (N_9691,N_6889,N_7210);
nand U9692 (N_9692,N_6694,N_6754);
or U9693 (N_9693,N_7464,N_6883);
xor U9694 (N_9694,N_7677,N_7855);
nor U9695 (N_9695,N_7914,N_6532);
nand U9696 (N_9696,N_7737,N_6583);
nand U9697 (N_9697,N_6849,N_7875);
nand U9698 (N_9698,N_7142,N_6004);
nor U9699 (N_9699,N_7507,N_6911);
or U9700 (N_9700,N_6477,N_7715);
or U9701 (N_9701,N_6551,N_6192);
and U9702 (N_9702,N_7964,N_6859);
and U9703 (N_9703,N_6567,N_7210);
and U9704 (N_9704,N_7894,N_6623);
nand U9705 (N_9705,N_6659,N_6140);
nor U9706 (N_9706,N_6676,N_7868);
and U9707 (N_9707,N_6644,N_7657);
nor U9708 (N_9708,N_6026,N_7789);
or U9709 (N_9709,N_7088,N_6303);
nand U9710 (N_9710,N_6904,N_6150);
nor U9711 (N_9711,N_6881,N_6366);
and U9712 (N_9712,N_7628,N_7763);
nand U9713 (N_9713,N_7810,N_7163);
xnor U9714 (N_9714,N_7657,N_6055);
xnor U9715 (N_9715,N_7804,N_6483);
nand U9716 (N_9716,N_7432,N_6647);
xor U9717 (N_9717,N_7576,N_6743);
and U9718 (N_9718,N_6212,N_6822);
nand U9719 (N_9719,N_7366,N_6862);
or U9720 (N_9720,N_7792,N_7606);
nor U9721 (N_9721,N_7700,N_6777);
or U9722 (N_9722,N_6459,N_6899);
and U9723 (N_9723,N_7593,N_6674);
and U9724 (N_9724,N_6917,N_6756);
xor U9725 (N_9725,N_7685,N_6906);
or U9726 (N_9726,N_6627,N_6970);
or U9727 (N_9727,N_7470,N_6340);
nor U9728 (N_9728,N_7402,N_7105);
and U9729 (N_9729,N_7506,N_6224);
and U9730 (N_9730,N_6771,N_7667);
and U9731 (N_9731,N_6490,N_6250);
xor U9732 (N_9732,N_6848,N_6011);
nand U9733 (N_9733,N_7302,N_6505);
xnor U9734 (N_9734,N_7576,N_6891);
nand U9735 (N_9735,N_7330,N_6472);
xnor U9736 (N_9736,N_7066,N_6816);
nor U9737 (N_9737,N_6547,N_7180);
nand U9738 (N_9738,N_6389,N_6848);
and U9739 (N_9739,N_6669,N_7098);
nand U9740 (N_9740,N_6612,N_6382);
or U9741 (N_9741,N_7202,N_7940);
or U9742 (N_9742,N_6808,N_7588);
nor U9743 (N_9743,N_6660,N_6184);
nand U9744 (N_9744,N_6661,N_6131);
xor U9745 (N_9745,N_6546,N_7999);
nor U9746 (N_9746,N_7621,N_6786);
nand U9747 (N_9747,N_6692,N_6072);
nand U9748 (N_9748,N_6380,N_6495);
xnor U9749 (N_9749,N_6830,N_7123);
nand U9750 (N_9750,N_6630,N_7066);
nor U9751 (N_9751,N_6034,N_7831);
or U9752 (N_9752,N_7954,N_7901);
xor U9753 (N_9753,N_6382,N_6840);
nand U9754 (N_9754,N_7599,N_7616);
or U9755 (N_9755,N_6427,N_6762);
or U9756 (N_9756,N_6511,N_6883);
xor U9757 (N_9757,N_6143,N_7531);
nand U9758 (N_9758,N_6399,N_7084);
xor U9759 (N_9759,N_6535,N_6983);
and U9760 (N_9760,N_7617,N_7494);
nand U9761 (N_9761,N_6954,N_6427);
nor U9762 (N_9762,N_6567,N_6215);
nor U9763 (N_9763,N_7126,N_7176);
nand U9764 (N_9764,N_6195,N_7179);
nor U9765 (N_9765,N_6339,N_6277);
and U9766 (N_9766,N_6807,N_6514);
and U9767 (N_9767,N_7378,N_7391);
nor U9768 (N_9768,N_7891,N_7918);
and U9769 (N_9769,N_7017,N_6258);
or U9770 (N_9770,N_6877,N_7344);
nor U9771 (N_9771,N_7656,N_6650);
nor U9772 (N_9772,N_6199,N_6796);
xnor U9773 (N_9773,N_6090,N_7600);
nor U9774 (N_9774,N_7307,N_6481);
nand U9775 (N_9775,N_6827,N_7445);
nor U9776 (N_9776,N_7647,N_7977);
nor U9777 (N_9777,N_7750,N_6907);
or U9778 (N_9778,N_7553,N_6190);
nand U9779 (N_9779,N_6463,N_6655);
or U9780 (N_9780,N_7159,N_6136);
nor U9781 (N_9781,N_6605,N_7471);
xnor U9782 (N_9782,N_6605,N_6087);
and U9783 (N_9783,N_7812,N_7536);
and U9784 (N_9784,N_6388,N_7677);
and U9785 (N_9785,N_6009,N_7849);
xor U9786 (N_9786,N_6360,N_6779);
nand U9787 (N_9787,N_7257,N_7336);
and U9788 (N_9788,N_6315,N_6289);
or U9789 (N_9789,N_6702,N_6715);
xor U9790 (N_9790,N_6974,N_7389);
or U9791 (N_9791,N_7774,N_6292);
and U9792 (N_9792,N_7875,N_6668);
nand U9793 (N_9793,N_7082,N_7999);
and U9794 (N_9794,N_6179,N_6029);
nor U9795 (N_9795,N_6954,N_7106);
or U9796 (N_9796,N_7005,N_7970);
nor U9797 (N_9797,N_6742,N_6968);
nand U9798 (N_9798,N_6053,N_7743);
xor U9799 (N_9799,N_7358,N_7209);
and U9800 (N_9800,N_6661,N_7009);
nand U9801 (N_9801,N_6047,N_6040);
nand U9802 (N_9802,N_6697,N_6867);
nor U9803 (N_9803,N_7806,N_7526);
nand U9804 (N_9804,N_6536,N_6668);
or U9805 (N_9805,N_7942,N_6807);
nor U9806 (N_9806,N_7189,N_7779);
and U9807 (N_9807,N_7664,N_6851);
and U9808 (N_9808,N_6640,N_7068);
and U9809 (N_9809,N_6204,N_7548);
or U9810 (N_9810,N_7882,N_6699);
or U9811 (N_9811,N_6297,N_6415);
and U9812 (N_9812,N_7039,N_7427);
nor U9813 (N_9813,N_7471,N_6167);
or U9814 (N_9814,N_7088,N_6487);
nor U9815 (N_9815,N_7251,N_7637);
and U9816 (N_9816,N_7395,N_6203);
nand U9817 (N_9817,N_7119,N_7851);
and U9818 (N_9818,N_7474,N_6744);
xor U9819 (N_9819,N_6920,N_6060);
xnor U9820 (N_9820,N_6630,N_7133);
and U9821 (N_9821,N_7232,N_7087);
nor U9822 (N_9822,N_6766,N_7785);
or U9823 (N_9823,N_6924,N_6169);
nand U9824 (N_9824,N_7352,N_7499);
or U9825 (N_9825,N_6498,N_7348);
nand U9826 (N_9826,N_7190,N_7375);
or U9827 (N_9827,N_6104,N_6719);
nand U9828 (N_9828,N_7773,N_7841);
and U9829 (N_9829,N_7399,N_6245);
nor U9830 (N_9830,N_7530,N_6925);
nand U9831 (N_9831,N_7771,N_7451);
or U9832 (N_9832,N_7668,N_6268);
nor U9833 (N_9833,N_7942,N_6453);
nand U9834 (N_9834,N_7336,N_6024);
xor U9835 (N_9835,N_7111,N_6347);
xnor U9836 (N_9836,N_7947,N_7036);
and U9837 (N_9837,N_6900,N_7056);
or U9838 (N_9838,N_7523,N_6317);
nand U9839 (N_9839,N_7080,N_6277);
xor U9840 (N_9840,N_6539,N_7612);
xor U9841 (N_9841,N_7340,N_6937);
or U9842 (N_9842,N_6203,N_7169);
xnor U9843 (N_9843,N_6951,N_6251);
nand U9844 (N_9844,N_6036,N_6465);
nand U9845 (N_9845,N_6272,N_6693);
nand U9846 (N_9846,N_6918,N_7539);
xnor U9847 (N_9847,N_7461,N_6419);
nor U9848 (N_9848,N_6375,N_6476);
and U9849 (N_9849,N_6552,N_7571);
or U9850 (N_9850,N_7268,N_7521);
and U9851 (N_9851,N_7608,N_7331);
nand U9852 (N_9852,N_6921,N_7469);
xnor U9853 (N_9853,N_6103,N_6898);
nor U9854 (N_9854,N_7607,N_7442);
or U9855 (N_9855,N_6732,N_6174);
or U9856 (N_9856,N_7810,N_6800);
and U9857 (N_9857,N_6238,N_7252);
and U9858 (N_9858,N_6182,N_7388);
nor U9859 (N_9859,N_7109,N_7213);
nor U9860 (N_9860,N_7366,N_7750);
and U9861 (N_9861,N_6551,N_6535);
nor U9862 (N_9862,N_6139,N_7307);
and U9863 (N_9863,N_7851,N_6409);
nand U9864 (N_9864,N_6087,N_7717);
nand U9865 (N_9865,N_7768,N_6094);
or U9866 (N_9866,N_6537,N_6077);
and U9867 (N_9867,N_6057,N_6218);
and U9868 (N_9868,N_6995,N_6901);
or U9869 (N_9869,N_7820,N_6340);
and U9870 (N_9870,N_7522,N_7271);
or U9871 (N_9871,N_6922,N_6960);
nor U9872 (N_9872,N_6694,N_7954);
or U9873 (N_9873,N_6642,N_7932);
nand U9874 (N_9874,N_7670,N_6697);
xor U9875 (N_9875,N_7796,N_6987);
xnor U9876 (N_9876,N_7602,N_6893);
xor U9877 (N_9877,N_6578,N_7222);
and U9878 (N_9878,N_7410,N_6167);
xnor U9879 (N_9879,N_6472,N_6241);
nor U9880 (N_9880,N_7671,N_7573);
and U9881 (N_9881,N_6947,N_7068);
xnor U9882 (N_9882,N_7418,N_6917);
or U9883 (N_9883,N_6827,N_7804);
and U9884 (N_9884,N_7173,N_6886);
and U9885 (N_9885,N_6386,N_6032);
and U9886 (N_9886,N_6957,N_6238);
xor U9887 (N_9887,N_7622,N_7376);
nor U9888 (N_9888,N_7154,N_7060);
nor U9889 (N_9889,N_6050,N_6043);
xnor U9890 (N_9890,N_6770,N_6838);
or U9891 (N_9891,N_7525,N_7707);
nor U9892 (N_9892,N_7304,N_7450);
or U9893 (N_9893,N_6598,N_6349);
and U9894 (N_9894,N_6600,N_6603);
nor U9895 (N_9895,N_6201,N_7204);
xor U9896 (N_9896,N_7217,N_6716);
nor U9897 (N_9897,N_6339,N_6434);
xor U9898 (N_9898,N_6289,N_7932);
and U9899 (N_9899,N_6343,N_6815);
xor U9900 (N_9900,N_7147,N_6244);
and U9901 (N_9901,N_7396,N_7844);
xor U9902 (N_9902,N_6247,N_6908);
or U9903 (N_9903,N_6155,N_6828);
xnor U9904 (N_9904,N_6340,N_6498);
xor U9905 (N_9905,N_6672,N_6980);
and U9906 (N_9906,N_7523,N_6522);
xnor U9907 (N_9907,N_7174,N_6510);
and U9908 (N_9908,N_7024,N_7615);
xor U9909 (N_9909,N_6191,N_6214);
and U9910 (N_9910,N_6576,N_7970);
nand U9911 (N_9911,N_6682,N_7859);
xnor U9912 (N_9912,N_6588,N_6398);
xnor U9913 (N_9913,N_6143,N_6162);
xor U9914 (N_9914,N_6199,N_6488);
nand U9915 (N_9915,N_6042,N_7463);
and U9916 (N_9916,N_7242,N_7907);
xnor U9917 (N_9917,N_7514,N_7462);
or U9918 (N_9918,N_6066,N_6183);
xnor U9919 (N_9919,N_7620,N_7180);
nand U9920 (N_9920,N_7525,N_6646);
nor U9921 (N_9921,N_7352,N_6119);
nor U9922 (N_9922,N_6855,N_7143);
nand U9923 (N_9923,N_6194,N_7051);
or U9924 (N_9924,N_7072,N_7710);
or U9925 (N_9925,N_6181,N_7196);
or U9926 (N_9926,N_7481,N_6396);
or U9927 (N_9927,N_7846,N_6520);
xor U9928 (N_9928,N_7254,N_7342);
and U9929 (N_9929,N_7286,N_7648);
and U9930 (N_9930,N_6888,N_7999);
xnor U9931 (N_9931,N_7709,N_7858);
and U9932 (N_9932,N_7962,N_7400);
nand U9933 (N_9933,N_6315,N_6431);
nor U9934 (N_9934,N_7722,N_6567);
xnor U9935 (N_9935,N_6254,N_6974);
and U9936 (N_9936,N_7192,N_6148);
nand U9937 (N_9937,N_6574,N_6198);
nor U9938 (N_9938,N_6481,N_6128);
xnor U9939 (N_9939,N_6281,N_6539);
xor U9940 (N_9940,N_7127,N_6726);
or U9941 (N_9941,N_7175,N_6835);
xnor U9942 (N_9942,N_6801,N_6986);
nand U9943 (N_9943,N_6645,N_6337);
xor U9944 (N_9944,N_7614,N_7811);
nor U9945 (N_9945,N_6872,N_7524);
xnor U9946 (N_9946,N_6620,N_7173);
nor U9947 (N_9947,N_7568,N_7011);
nor U9948 (N_9948,N_7543,N_7354);
or U9949 (N_9949,N_7722,N_7512);
and U9950 (N_9950,N_6593,N_7822);
or U9951 (N_9951,N_6051,N_6611);
or U9952 (N_9952,N_7131,N_7521);
nor U9953 (N_9953,N_7648,N_7292);
xnor U9954 (N_9954,N_7251,N_6351);
nand U9955 (N_9955,N_7810,N_6134);
nand U9956 (N_9956,N_6816,N_6106);
or U9957 (N_9957,N_7528,N_7119);
nand U9958 (N_9958,N_7414,N_7635);
xor U9959 (N_9959,N_6150,N_6469);
nor U9960 (N_9960,N_6512,N_7377);
and U9961 (N_9961,N_6978,N_6937);
and U9962 (N_9962,N_6707,N_7946);
or U9963 (N_9963,N_6700,N_6355);
and U9964 (N_9964,N_6976,N_7193);
or U9965 (N_9965,N_6008,N_6785);
xnor U9966 (N_9966,N_6574,N_6110);
or U9967 (N_9967,N_7666,N_7723);
xnor U9968 (N_9968,N_6532,N_7981);
xnor U9969 (N_9969,N_7783,N_6449);
nand U9970 (N_9970,N_7672,N_6209);
and U9971 (N_9971,N_7298,N_7581);
or U9972 (N_9972,N_6758,N_7104);
and U9973 (N_9973,N_6747,N_7151);
nor U9974 (N_9974,N_7497,N_6634);
xnor U9975 (N_9975,N_7530,N_6823);
or U9976 (N_9976,N_6596,N_7990);
and U9977 (N_9977,N_6910,N_7800);
xnor U9978 (N_9978,N_6029,N_7979);
or U9979 (N_9979,N_7218,N_6117);
xor U9980 (N_9980,N_7822,N_6096);
or U9981 (N_9981,N_7192,N_6872);
or U9982 (N_9982,N_7135,N_7187);
nand U9983 (N_9983,N_6187,N_7685);
and U9984 (N_9984,N_6097,N_7092);
xor U9985 (N_9985,N_6871,N_6365);
xnor U9986 (N_9986,N_6361,N_6947);
xnor U9987 (N_9987,N_6942,N_6265);
xor U9988 (N_9988,N_6825,N_7592);
nor U9989 (N_9989,N_7230,N_7088);
nand U9990 (N_9990,N_6128,N_7748);
or U9991 (N_9991,N_6728,N_6202);
nand U9992 (N_9992,N_7891,N_6098);
xor U9993 (N_9993,N_6879,N_7286);
nand U9994 (N_9994,N_6940,N_7848);
nand U9995 (N_9995,N_7314,N_7253);
and U9996 (N_9996,N_7465,N_6156);
xor U9997 (N_9997,N_6790,N_7101);
nor U9998 (N_9998,N_7550,N_7765);
nor U9999 (N_9999,N_6665,N_6333);
nand UO_0 (O_0,N_8284,N_8897);
or UO_1 (O_1,N_9861,N_8115);
nor UO_2 (O_2,N_9674,N_9933);
and UO_3 (O_3,N_8416,N_9431);
nor UO_4 (O_4,N_8433,N_9243);
or UO_5 (O_5,N_8578,N_8007);
and UO_6 (O_6,N_9554,N_8582);
or UO_7 (O_7,N_9626,N_9163);
or UO_8 (O_8,N_8310,N_8363);
xnor UO_9 (O_9,N_9551,N_9493);
xnor UO_10 (O_10,N_8927,N_8367);
or UO_11 (O_11,N_8583,N_9498);
and UO_12 (O_12,N_9833,N_8577);
xnor UO_13 (O_13,N_9687,N_8269);
xnor UO_14 (O_14,N_8759,N_9753);
xor UO_15 (O_15,N_8697,N_9781);
nor UO_16 (O_16,N_8459,N_9420);
or UO_17 (O_17,N_8353,N_9476);
nor UO_18 (O_18,N_8740,N_9596);
or UO_19 (O_19,N_8045,N_9682);
nor UO_20 (O_20,N_9218,N_9441);
nand UO_21 (O_21,N_8711,N_8151);
nand UO_22 (O_22,N_8898,N_8214);
or UO_23 (O_23,N_9110,N_8820);
nor UO_24 (O_24,N_8256,N_9808);
nor UO_25 (O_25,N_9726,N_8610);
nor UO_26 (O_26,N_9225,N_8388);
xnor UO_27 (O_27,N_9750,N_8192);
and UO_28 (O_28,N_9349,N_9401);
xor UO_29 (O_29,N_9516,N_9670);
nand UO_30 (O_30,N_9459,N_8602);
or UO_31 (O_31,N_8948,N_9511);
and UO_32 (O_32,N_8790,N_8035);
or UO_33 (O_33,N_9041,N_9346);
and UO_34 (O_34,N_9928,N_8975);
nor UO_35 (O_35,N_9977,N_8712);
xnor UO_36 (O_36,N_8634,N_8095);
xor UO_37 (O_37,N_8184,N_8937);
nand UO_38 (O_38,N_9767,N_9644);
nand UO_39 (O_39,N_8798,N_9173);
or UO_40 (O_40,N_9294,N_8465);
and UO_41 (O_41,N_8397,N_9117);
nor UO_42 (O_42,N_9895,N_8633);
and UO_43 (O_43,N_8562,N_9413);
nand UO_44 (O_44,N_9048,N_8042);
and UO_45 (O_45,N_9394,N_9399);
nor UO_46 (O_46,N_9318,N_8274);
or UO_47 (O_47,N_8655,N_8406);
nand UO_48 (O_48,N_8263,N_9412);
and UO_49 (O_49,N_9544,N_9744);
xnor UO_50 (O_50,N_9558,N_8296);
or UO_51 (O_51,N_9968,N_9052);
and UO_52 (O_52,N_9663,N_9321);
and UO_53 (O_53,N_9245,N_8495);
xnor UO_54 (O_54,N_9502,N_9375);
and UO_55 (O_55,N_8421,N_9652);
nor UO_56 (O_56,N_9074,N_8466);
nor UO_57 (O_57,N_9961,N_8598);
nor UO_58 (O_58,N_9365,N_8411);
nor UO_59 (O_59,N_8906,N_9216);
nor UO_60 (O_60,N_9098,N_8096);
or UO_61 (O_61,N_8036,N_9610);
nor UO_62 (O_62,N_8166,N_8858);
xnor UO_63 (O_63,N_9971,N_9746);
xnor UO_64 (O_64,N_9478,N_8793);
xor UO_65 (O_65,N_8735,N_8567);
and UO_66 (O_66,N_8765,N_9514);
nand UO_67 (O_67,N_8855,N_8227);
or UO_68 (O_68,N_9875,N_9143);
nor UO_69 (O_69,N_9784,N_8928);
xor UO_70 (O_70,N_9240,N_8805);
or UO_71 (O_71,N_9211,N_8581);
and UO_72 (O_72,N_8891,N_9629);
and UO_73 (O_73,N_8208,N_9060);
xor UO_74 (O_74,N_9927,N_8165);
nor UO_75 (O_75,N_9319,N_8448);
xor UO_76 (O_76,N_9046,N_8778);
xor UO_77 (O_77,N_9569,N_9721);
and UO_78 (O_78,N_9988,N_9757);
and UO_79 (O_79,N_8969,N_9012);
xor UO_80 (O_80,N_9035,N_8326);
nand UO_81 (O_81,N_8113,N_8400);
xor UO_82 (O_82,N_9992,N_9850);
nand UO_83 (O_83,N_8624,N_9199);
nand UO_84 (O_84,N_8369,N_9181);
nand UO_85 (O_85,N_9882,N_8625);
nand UO_86 (O_86,N_8961,N_9696);
and UO_87 (O_87,N_8370,N_8059);
or UO_88 (O_88,N_8878,N_8279);
nand UO_89 (O_89,N_9632,N_8707);
nor UO_90 (O_90,N_9135,N_9924);
and UO_91 (O_91,N_9213,N_9567);
xnor UO_92 (O_92,N_8484,N_9407);
nor UO_93 (O_93,N_8365,N_8239);
nor UO_94 (O_94,N_8360,N_8201);
and UO_95 (O_95,N_8571,N_8978);
xor UO_96 (O_96,N_9112,N_9241);
and UO_97 (O_97,N_8398,N_8687);
or UO_98 (O_98,N_8872,N_9492);
or UO_99 (O_99,N_9804,N_9150);
and UO_100 (O_100,N_8109,N_9279);
xor UO_101 (O_101,N_8882,N_8250);
or UO_102 (O_102,N_9075,N_8440);
nand UO_103 (O_103,N_9376,N_8973);
xor UO_104 (O_104,N_8290,N_9935);
and UO_105 (O_105,N_9174,N_9071);
nand UO_106 (O_106,N_9751,N_8833);
or UO_107 (O_107,N_9919,N_9536);
and UO_108 (O_108,N_8424,N_9404);
xnor UO_109 (O_109,N_9897,N_9568);
nor UO_110 (O_110,N_9099,N_9377);
or UO_111 (O_111,N_8061,N_9450);
nor UO_112 (O_112,N_8838,N_8866);
and UO_113 (O_113,N_9590,N_8220);
nor UO_114 (O_114,N_9406,N_8216);
or UO_115 (O_115,N_9288,N_9555);
nand UO_116 (O_116,N_9534,N_8880);
nor UO_117 (O_117,N_8899,N_8422);
nand UO_118 (O_118,N_8168,N_9417);
xor UO_119 (O_119,N_8609,N_9396);
xor UO_120 (O_120,N_9352,N_9649);
or UO_121 (O_121,N_9853,N_9341);
or UO_122 (O_122,N_8195,N_9540);
nand UO_123 (O_123,N_9081,N_9316);
nand UO_124 (O_124,N_8301,N_9068);
or UO_125 (O_125,N_8558,N_8563);
nand UO_126 (O_126,N_9194,N_9965);
xnor UO_127 (O_127,N_9917,N_8734);
nand UO_128 (O_128,N_8233,N_9799);
and UO_129 (O_129,N_9446,N_8011);
nor UO_130 (O_130,N_8393,N_9521);
and UO_131 (O_131,N_8314,N_9599);
and UO_132 (O_132,N_8156,N_9323);
or UO_133 (O_133,N_9116,N_9080);
nor UO_134 (O_134,N_9617,N_8447);
or UO_135 (O_135,N_8530,N_8564);
nor UO_136 (O_136,N_8514,N_8506);
xor UO_137 (O_137,N_8731,N_9711);
xnor UO_138 (O_138,N_8933,N_8328);
nand UO_139 (O_139,N_9891,N_8589);
or UO_140 (O_140,N_8922,N_9328);
and UO_141 (O_141,N_9970,N_8110);
and UO_142 (O_142,N_9641,N_8278);
xnor UO_143 (O_143,N_9628,N_8334);
nor UO_144 (O_144,N_8728,N_9087);
and UO_145 (O_145,N_9921,N_8202);
nand UO_146 (O_146,N_9039,N_9593);
or UO_147 (O_147,N_8392,N_8623);
nor UO_148 (O_148,N_8368,N_9077);
nor UO_149 (O_149,N_9154,N_9300);
nand UO_150 (O_150,N_8283,N_8148);
and UO_151 (O_151,N_8870,N_9219);
xnor UO_152 (O_152,N_9748,N_8966);
xor UO_153 (O_153,N_9095,N_8129);
nand UO_154 (O_154,N_8139,N_8854);
nor UO_155 (O_155,N_8967,N_9957);
nor UO_156 (O_156,N_9911,N_8699);
nand UO_157 (O_157,N_9723,N_8814);
nand UO_158 (O_158,N_8128,N_8942);
nor UO_159 (O_159,N_9036,N_9545);
nor UO_160 (O_160,N_9899,N_9474);
nor UO_161 (O_161,N_8458,N_8487);
or UO_162 (O_162,N_8277,N_9614);
and UO_163 (O_163,N_9572,N_8786);
nor UO_164 (O_164,N_9651,N_8690);
nand UO_165 (O_165,N_8750,N_8030);
nand UO_166 (O_166,N_9156,N_8654);
xor UO_167 (O_167,N_9477,N_8588);
xor UO_168 (O_168,N_9857,N_9597);
or UO_169 (O_169,N_8513,N_9105);
and UO_170 (O_170,N_8902,N_8819);
and UO_171 (O_171,N_8286,N_8299);
xnor UO_172 (O_172,N_8916,N_9267);
xor UO_173 (O_173,N_9463,N_9938);
or UO_174 (O_174,N_9662,N_8641);
or UO_175 (O_175,N_9955,N_9166);
nor UO_176 (O_176,N_8794,N_9761);
nand UO_177 (O_177,N_9419,N_9167);
nand UO_178 (O_178,N_8124,N_8173);
xnor UO_179 (O_179,N_9027,N_9290);
nor UO_180 (O_180,N_9981,N_8232);
xnor UO_181 (O_181,N_9089,N_8158);
or UO_182 (O_182,N_9284,N_8373);
nand UO_183 (O_183,N_9887,N_8839);
and UO_184 (O_184,N_8518,N_8442);
xor UO_185 (O_185,N_8021,N_8169);
and UO_186 (O_186,N_9920,N_8685);
or UO_187 (O_187,N_8972,N_8748);
nor UO_188 (O_188,N_9340,N_8593);
and UO_189 (O_189,N_8663,N_9265);
xnor UO_190 (O_190,N_9136,N_9625);
nand UO_191 (O_191,N_9805,N_8108);
and UO_192 (O_192,N_9313,N_8445);
nor UO_193 (O_193,N_9310,N_9846);
nand UO_194 (O_194,N_9795,N_9679);
nor UO_195 (O_195,N_8758,N_8816);
nand UO_196 (O_196,N_8517,N_9496);
and UO_197 (O_197,N_9220,N_8742);
nor UO_198 (O_198,N_9004,N_8006);
nor UO_199 (O_199,N_8535,N_9524);
nor UO_200 (O_200,N_8428,N_8215);
and UO_201 (O_201,N_9342,N_8436);
and UO_202 (O_202,N_8070,N_8954);
or UO_203 (O_203,N_9683,N_8318);
nor UO_204 (O_204,N_9792,N_8426);
nor UO_205 (O_205,N_9315,N_8483);
nor UO_206 (O_206,N_9699,N_8842);
nand UO_207 (O_207,N_8811,N_9791);
or UO_208 (O_208,N_9725,N_8821);
xnor UO_209 (O_209,N_8383,N_8651);
nand UO_210 (O_210,N_8425,N_9734);
nand UO_211 (O_211,N_8000,N_9209);
or UO_212 (O_212,N_9034,N_8417);
and UO_213 (O_213,N_8313,N_8726);
nand UO_214 (O_214,N_9661,N_9690);
or UO_215 (O_215,N_8604,N_8116);
nor UO_216 (O_216,N_9630,N_8949);
nor UO_217 (O_217,N_8481,N_9325);
nor UO_218 (O_218,N_8595,N_8437);
xnor UO_219 (O_219,N_8971,N_8812);
or UO_220 (O_220,N_9429,N_8402);
or UO_221 (O_221,N_9374,N_8378);
and UO_222 (O_222,N_8607,N_8753);
xnor UO_223 (O_223,N_8701,N_9088);
nor UO_224 (O_224,N_8456,N_8196);
nor UO_225 (O_225,N_9435,N_9364);
and UO_226 (O_226,N_8253,N_9494);
xnor UO_227 (O_227,N_9983,N_8432);
nand UO_228 (O_228,N_8941,N_8910);
and UO_229 (O_229,N_9118,N_8025);
nor UO_230 (O_230,N_8919,N_8836);
or UO_231 (O_231,N_8499,N_8903);
nor UO_232 (O_232,N_9519,N_8862);
nand UO_233 (O_233,N_8935,N_8123);
and UO_234 (O_234,N_9888,N_9353);
nand UO_235 (O_235,N_9266,N_9594);
and UO_236 (O_236,N_8665,N_8159);
nor UO_237 (O_237,N_9892,N_9874);
and UO_238 (O_238,N_9930,N_8078);
nand UO_239 (O_239,N_9100,N_8852);
xor UO_240 (O_240,N_8657,N_9103);
or UO_241 (O_241,N_9264,N_8901);
and UO_242 (O_242,N_8646,N_8469);
nor UO_243 (O_243,N_8741,N_9102);
nand UO_244 (O_244,N_8280,N_8692);
xnor UO_245 (O_245,N_9416,N_8028);
nor UO_246 (O_246,N_8700,N_8213);
nor UO_247 (O_247,N_8549,N_8174);
xnor UO_248 (O_248,N_8240,N_9769);
nor UO_249 (O_249,N_8218,N_8755);
nor UO_250 (O_250,N_8621,N_9581);
nor UO_251 (O_251,N_8292,N_9789);
xor UO_252 (O_252,N_9856,N_9454);
nand UO_253 (O_253,N_8815,N_9021);
or UO_254 (O_254,N_9849,N_8675);
or UO_255 (O_255,N_9692,N_9042);
nand UO_256 (O_256,N_8223,N_9274);
and UO_257 (O_257,N_9326,N_9573);
and UO_258 (O_258,N_8611,N_9164);
or UO_259 (O_259,N_9383,N_8323);
nor UO_260 (O_260,N_9871,N_9282);
or UO_261 (O_261,N_9738,N_9660);
and UO_262 (O_262,N_8531,N_9432);
xor UO_263 (O_263,N_9586,N_8463);
xnor UO_264 (O_264,N_9841,N_9504);
nand UO_265 (O_265,N_9385,N_8049);
or UO_266 (O_266,N_9121,N_8260);
nor UO_267 (O_267,N_8614,N_8863);
nor UO_268 (O_268,N_9691,N_8014);
nor UO_269 (O_269,N_9794,N_8211);
nor UO_270 (O_270,N_8527,N_8546);
nor UO_271 (O_271,N_9720,N_9873);
nand UO_272 (O_272,N_8023,N_9400);
nor UO_273 (O_273,N_8075,N_9025);
xnor UO_274 (O_274,N_8013,N_9905);
xor UO_275 (O_275,N_9855,N_8027);
xor UO_276 (O_276,N_9427,N_9602);
and UO_277 (O_277,N_8390,N_8552);
and UO_278 (O_278,N_8224,N_9591);
or UO_279 (O_279,N_9158,N_8565);
xnor UO_280 (O_280,N_8236,N_8321);
xnor UO_281 (O_281,N_9276,N_9996);
nand UO_282 (O_282,N_9190,N_8057);
nand UO_283 (O_283,N_8818,N_9939);
nand UO_284 (O_284,N_9575,N_9183);
or UO_285 (O_285,N_8860,N_9155);
nor UO_286 (O_286,N_8715,N_8478);
and UO_287 (O_287,N_8770,N_9522);
xor UO_288 (O_288,N_9178,N_8887);
and UO_289 (O_289,N_9775,N_9595);
nand UO_290 (O_290,N_8122,N_9329);
xnor UO_291 (O_291,N_9758,N_8405);
nand UO_292 (O_292,N_8352,N_9191);
nor UO_293 (O_293,N_8460,N_9210);
xor UO_294 (O_294,N_9999,N_8620);
xnor UO_295 (O_295,N_9906,N_9923);
or UO_296 (O_296,N_8217,N_8963);
or UO_297 (O_297,N_9169,N_9017);
nand UO_298 (O_298,N_8376,N_9640);
nor UO_299 (O_299,N_9526,N_9186);
and UO_300 (O_300,N_8317,N_9373);
nand UO_301 (O_301,N_8627,N_8990);
xnor UO_302 (O_302,N_8234,N_9562);
nand UO_303 (O_303,N_9509,N_9051);
nor UO_304 (O_304,N_9127,N_9826);
nand UO_305 (O_305,N_9161,N_9782);
nor UO_306 (O_306,N_8681,N_8039);
xnor UO_307 (O_307,N_8282,N_9543);
and UO_308 (O_308,N_8419,N_9370);
or UO_309 (O_309,N_9330,N_8067);
or UO_310 (O_310,N_9079,N_8490);
nand UO_311 (O_311,N_8024,N_9876);
nor UO_312 (O_312,N_9713,N_8658);
xnor UO_313 (O_313,N_9254,N_8890);
and UO_314 (O_314,N_8892,N_8287);
xor UO_315 (O_315,N_8394,N_9903);
and UO_316 (O_316,N_8205,N_9528);
and UO_317 (O_317,N_9234,N_9106);
nand UO_318 (O_318,N_8841,N_9836);
nand UO_319 (O_319,N_9816,N_8354);
xor UO_320 (O_320,N_8653,N_8320);
nor UO_321 (O_321,N_8356,N_8795);
xor UO_322 (O_322,N_8958,N_9842);
and UO_323 (O_323,N_9643,N_8467);
and UO_324 (O_324,N_9016,N_9650);
xnor UO_325 (O_325,N_9623,N_9913);
xnor UO_326 (O_326,N_9442,N_8180);
nor UO_327 (O_327,N_8915,N_8566);
nor UO_328 (O_328,N_9718,N_8084);
and UO_329 (O_329,N_9667,N_8612);
nor UO_330 (O_330,N_9179,N_8529);
and UO_331 (O_331,N_9580,N_8034);
nand UO_332 (O_332,N_9680,N_8785);
nand UO_333 (O_333,N_9860,N_9578);
nor UO_334 (O_334,N_8808,N_9658);
xor UO_335 (O_335,N_8064,N_8606);
xor UO_336 (O_336,N_8187,N_9987);
xor UO_337 (O_337,N_9946,N_9023);
nor UO_338 (O_338,N_9390,N_9722);
and UO_339 (O_339,N_9076,N_9908);
or UO_340 (O_340,N_8957,N_9295);
xnor UO_341 (O_341,N_8666,N_8569);
and UO_342 (O_342,N_9635,N_8893);
nand UO_343 (O_343,N_9348,N_8207);
and UO_344 (O_344,N_9986,N_8473);
and UO_345 (O_345,N_9205,N_9759);
nand UO_346 (O_346,N_8721,N_8724);
nor UO_347 (O_347,N_8077,N_9851);
and UO_348 (O_348,N_8702,N_8757);
nand UO_349 (O_349,N_9773,N_8306);
xnor UO_350 (O_350,N_9246,N_9609);
and UO_351 (O_351,N_9272,N_9426);
nand UO_352 (O_352,N_8051,N_9786);
or UO_353 (O_353,N_8349,N_8760);
nor UO_354 (O_354,N_8541,N_9015);
nand UO_355 (O_355,N_8337,N_9716);
or UO_356 (O_356,N_8270,N_8194);
nand UO_357 (O_357,N_9384,N_9501);
nor UO_358 (O_358,N_8093,N_9737);
and UO_359 (O_359,N_8097,N_9688);
nor UO_360 (O_360,N_9527,N_8576);
nor UO_361 (O_361,N_9483,N_8150);
xor UO_362 (O_362,N_9359,N_9852);
nand UO_363 (O_363,N_8829,N_9506);
nand UO_364 (O_364,N_8824,N_9393);
xnor UO_365 (O_365,N_8508,N_8912);
nand UO_366 (O_366,N_8943,N_9916);
or UO_367 (O_367,N_9508,N_9756);
and UO_368 (O_368,N_9481,N_8178);
xnor UO_369 (O_369,N_9010,N_9411);
or UO_370 (O_370,N_9584,N_8950);
nand UO_371 (O_371,N_8273,N_8964);
or UO_372 (O_372,N_9050,N_9779);
nor UO_373 (O_373,N_8082,N_8412);
or UO_374 (O_374,N_8226,N_8331);
nand UO_375 (O_375,N_9337,N_9410);
xnor UO_376 (O_376,N_9320,N_9956);
xor UO_377 (O_377,N_9133,N_9336);
or UO_378 (O_378,N_8905,N_9083);
or UO_379 (O_379,N_9520,N_9589);
nand UO_380 (O_380,N_8308,N_8081);
or UO_381 (O_381,N_9648,N_8525);
and UO_382 (O_382,N_9530,N_9712);
xnor UO_383 (O_383,N_9188,N_8026);
xor UO_384 (O_384,N_8381,N_8859);
xnor UO_385 (O_385,N_8868,N_9512);
nor UO_386 (O_386,N_9460,N_8800);
and UO_387 (O_387,N_8477,N_8198);
or UO_388 (O_388,N_9217,N_9557);
xor UO_389 (O_389,N_9303,N_8351);
and UO_390 (O_390,N_9587,N_8848);
xnor UO_391 (O_391,N_8387,N_9269);
and UO_392 (O_392,N_9745,N_8120);
or UO_393 (O_393,N_8560,N_9382);
xor UO_394 (O_394,N_8519,N_9812);
and UO_395 (O_395,N_8019,N_9838);
xor UO_396 (O_396,N_9252,N_8175);
nor UO_397 (O_397,N_9624,N_8407);
or UO_398 (O_398,N_9566,N_8145);
or UO_399 (O_399,N_9685,N_8012);
and UO_400 (O_400,N_9764,N_8341);
and UO_401 (O_401,N_8058,N_8522);
and UO_402 (O_402,N_9736,N_8930);
xor UO_403 (O_403,N_8678,N_8831);
and UO_404 (O_404,N_8118,N_8345);
or UO_405 (O_405,N_8510,N_8225);
or UO_406 (O_406,N_9162,N_8293);
xor UO_407 (O_407,N_8568,N_8585);
nand UO_408 (O_408,N_8300,N_9458);
nand UO_409 (O_409,N_9292,N_9616);
nand UO_410 (O_410,N_9697,N_9006);
or UO_411 (O_411,N_8737,N_9107);
nor UO_412 (O_412,N_8291,N_9249);
nand UO_413 (O_413,N_9433,N_8083);
nand UO_414 (O_414,N_9499,N_9468);
and UO_415 (O_415,N_9490,N_8521);
nor UO_416 (O_416,N_9031,N_9148);
xnor UO_417 (O_417,N_9084,N_9024);
xor UO_418 (O_418,N_9980,N_8777);
or UO_419 (O_419,N_9028,N_8020);
nor UO_420 (O_420,N_9994,N_8162);
nor UO_421 (O_421,N_8864,N_9467);
or UO_422 (O_422,N_8106,N_8696);
nor UO_423 (O_423,N_9627,N_8660);
nand UO_424 (O_424,N_8479,N_9991);
and UO_425 (O_425,N_8252,N_8523);
nand UO_426 (O_426,N_8616,N_9139);
and UO_427 (O_427,N_8524,N_9408);
nor UO_428 (O_428,N_9695,N_9275);
nor UO_429 (O_429,N_9440,N_9086);
or UO_430 (O_430,N_9742,N_8430);
or UO_431 (O_431,N_9090,N_8248);
nand UO_432 (O_432,N_9108,N_9176);
nand UO_433 (O_433,N_8289,N_8584);
nor UO_434 (O_434,N_9879,N_9356);
nand UO_435 (O_435,N_8114,N_9771);
and UO_436 (O_436,N_8257,N_8810);
xnor UO_437 (O_437,N_9403,N_8255);
or UO_438 (O_438,N_8925,N_9355);
and UO_439 (O_439,N_9259,N_8222);
xnor UO_440 (O_440,N_9262,N_8764);
or UO_441 (O_441,N_8404,N_8200);
or UO_442 (O_442,N_9634,N_8684);
xnor UO_443 (O_443,N_8587,N_8705);
or UO_444 (O_444,N_8126,N_9029);
xor UO_445 (O_445,N_9618,N_9487);
and UO_446 (O_446,N_8497,N_9455);
and UO_447 (O_447,N_8475,N_9807);
or UO_448 (O_448,N_8135,N_9130);
and UO_449 (O_449,N_8107,N_8883);
nand UO_450 (O_450,N_8998,N_9470);
and UO_451 (O_451,N_9867,N_9193);
xnor UO_452 (O_452,N_8063,N_9507);
nor UO_453 (O_453,N_9126,N_9308);
nand UO_454 (O_454,N_8160,N_9324);
nand UO_455 (O_455,N_8676,N_9449);
nor UO_456 (O_456,N_9009,N_9840);
and UO_457 (O_457,N_8285,N_8244);
or UO_458 (O_458,N_8254,N_9914);
nor UO_459 (O_459,N_9729,N_8913);
and UO_460 (O_460,N_8994,N_8347);
xnor UO_461 (O_461,N_8085,N_9054);
nor UO_462 (O_462,N_9960,N_8544);
nand UO_463 (O_463,N_9367,N_9546);
or UO_464 (O_464,N_9457,N_8782);
nand UO_465 (O_465,N_9157,N_8879);
xor UO_466 (O_466,N_8488,N_8867);
xor UO_467 (O_467,N_9604,N_9797);
nor UO_468 (O_468,N_8837,N_8668);
and UO_469 (O_469,N_8190,N_9395);
or UO_470 (O_470,N_9832,N_8679);
nor UO_471 (O_471,N_8851,N_9684);
or UO_472 (O_472,N_9196,N_9639);
and UO_473 (O_473,N_8149,N_9883);
nand UO_474 (O_474,N_9865,N_9366);
and UO_475 (O_475,N_8336,N_8993);
or UO_476 (O_476,N_8502,N_8276);
or UO_477 (O_477,N_8888,N_8454);
xnor UO_478 (O_478,N_9656,N_9995);
nor UO_479 (O_479,N_9304,N_8926);
nor UO_480 (O_480,N_8209,N_8018);
nor UO_481 (O_481,N_9915,N_9280);
and UO_482 (O_482,N_8505,N_8717);
nand UO_483 (O_483,N_8267,N_8686);
and UO_484 (O_484,N_9945,N_9184);
xnor UO_485 (O_485,N_8762,N_9170);
nor UO_486 (O_486,N_9984,N_9369);
nor UO_487 (O_487,N_8297,N_9621);
and UO_488 (O_488,N_8212,N_9447);
xor UO_489 (O_489,N_8143,N_9825);
and UO_490 (O_490,N_8161,N_8141);
nor UO_491 (O_491,N_8959,N_8086);
or UO_492 (O_492,N_8573,N_8545);
nor UO_493 (O_493,N_8089,N_8738);
nor UO_494 (O_494,N_9011,N_8179);
and UO_495 (O_495,N_9706,N_8896);
xnor UO_496 (O_496,N_9392,N_8340);
xnor UO_497 (O_497,N_9398,N_8048);
xnor UO_498 (O_498,N_9704,N_9032);
and UO_499 (O_499,N_8710,N_9951);
and UO_500 (O_500,N_8774,N_9338);
or UO_501 (O_501,N_8999,N_9654);
and UO_502 (O_502,N_9870,N_9822);
nor UO_503 (O_503,N_8043,N_9676);
and UO_504 (O_504,N_9475,N_9787);
and UO_505 (O_505,N_9452,N_9529);
and UO_506 (O_506,N_9577,N_9675);
and UO_507 (O_507,N_8540,N_8894);
nor UO_508 (O_508,N_9912,N_9293);
nand UO_509 (O_509,N_8929,N_9926);
nand UO_510 (O_510,N_8603,N_9270);
and UO_511 (O_511,N_8622,N_8435);
or UO_512 (O_512,N_8979,N_8840);
or UO_513 (O_513,N_8694,N_8644);
xnor UO_514 (O_514,N_9005,N_9138);
xnor UO_515 (O_515,N_8041,N_9715);
and UO_516 (O_516,N_8924,N_9045);
nand UO_517 (O_517,N_8674,N_8379);
or UO_518 (O_518,N_9619,N_8727);
and UO_519 (O_519,N_9067,N_8264);
xnor UO_520 (O_520,N_8142,N_9070);
nand UO_521 (O_521,N_8137,N_9014);
nand UO_522 (O_522,N_8427,N_9189);
nand UO_523 (O_523,N_8548,N_9443);
nor UO_524 (O_524,N_9880,N_9693);
xnor UO_525 (O_525,N_8374,N_8889);
and UO_526 (O_526,N_8471,N_9877);
and UO_527 (O_527,N_8989,N_8493);
nand UO_528 (O_528,N_9236,N_9603);
or UO_529 (O_529,N_8956,N_9372);
xnor UO_530 (O_530,N_9762,N_9525);
nor UO_531 (O_531,N_9064,N_8638);
nand UO_532 (O_532,N_8511,N_9668);
xor UO_533 (O_533,N_8673,N_9129);
xor UO_534 (O_534,N_9488,N_9985);
or UO_535 (O_535,N_9497,N_8281);
xnor UO_536 (O_536,N_9043,N_9535);
or UO_537 (O_537,N_9934,N_9612);
or UO_538 (O_538,N_8875,N_8635);
or UO_539 (O_539,N_9843,N_8102);
xnor UO_540 (O_540,N_8932,N_9776);
and UO_541 (O_541,N_9462,N_8884);
nand UO_542 (O_542,N_9778,N_8921);
or UO_543 (O_543,N_9285,N_9834);
nand UO_544 (O_544,N_9653,N_8130);
xor UO_545 (O_545,N_9113,N_9228);
and UO_546 (O_546,N_8494,N_9247);
nor UO_547 (O_547,N_9258,N_9018);
or UO_548 (O_548,N_9495,N_9149);
nor UO_549 (O_549,N_8713,N_8642);
xor UO_550 (O_550,N_8305,N_9503);
xor UO_551 (O_551,N_9765,N_9085);
nor UO_552 (O_552,N_9044,N_8050);
nand UO_553 (O_553,N_9114,N_8462);
and UO_554 (O_554,N_8303,N_9013);
nand UO_555 (O_555,N_9542,N_9571);
and UO_556 (O_556,N_8788,N_9645);
or UO_557 (O_557,N_9907,N_8617);
nor UO_558 (O_558,N_8366,N_9466);
nand UO_559 (O_559,N_9388,N_9159);
nand UO_560 (O_560,N_9901,N_9473);
or UO_561 (O_561,N_8265,N_9140);
and UO_562 (O_562,N_8453,N_8722);
or UO_563 (O_563,N_9289,N_8125);
nand UO_564 (O_564,N_8055,N_8613);
or UO_565 (O_565,N_8052,N_8556);
nor UO_566 (O_566,N_8991,N_8251);
xnor UO_567 (O_567,N_9890,N_9523);
nor UO_568 (O_568,N_8500,N_9491);
nor UO_569 (O_569,N_8934,N_8418);
nand UO_570 (O_570,N_9539,N_8672);
or UO_571 (O_571,N_9561,N_8485);
and UO_572 (O_572,N_8992,N_8714);
and UO_573 (O_573,N_8261,N_9425);
nand UO_574 (O_574,N_8662,N_9958);
xnor UO_575 (O_575,N_9471,N_8339);
xor UO_576 (O_576,N_9671,N_9096);
nand UO_577 (O_577,N_9343,N_9277);
nand UO_578 (O_578,N_9563,N_8984);
and UO_579 (O_579,N_9741,N_9302);
nand UO_580 (O_580,N_8865,N_9172);
nor UO_581 (O_581,N_8350,N_8335);
and UO_582 (O_582,N_9091,N_9197);
and UO_583 (O_583,N_9109,N_9553);
and UO_584 (O_584,N_8586,N_8316);
nand UO_585 (O_585,N_9378,N_9831);
nor UO_586 (O_586,N_9898,N_8241);
xnor UO_587 (O_587,N_9824,N_8009);
and UO_588 (O_588,N_9165,N_9312);
or UO_589 (O_589,N_8074,N_8103);
xor UO_590 (O_590,N_8420,N_9798);
nor UO_591 (O_591,N_9620,N_8974);
nor UO_592 (O_592,N_9803,N_9423);
or UO_593 (O_593,N_8791,N_8784);
and UO_594 (O_594,N_8723,N_8804);
nand UO_595 (O_595,N_9248,N_9698);
nor UO_596 (O_596,N_8689,N_9869);
xor UO_597 (O_597,N_8004,N_8329);
and UO_598 (O_598,N_8615,N_8532);
and UO_599 (O_599,N_9207,N_9864);
nand UO_600 (O_600,N_8033,N_8375);
nor UO_601 (O_601,N_8091,N_9037);
xor UO_602 (O_602,N_8008,N_9469);
and UO_603 (O_603,N_9049,N_9802);
nand UO_604 (O_604,N_9730,N_9607);
and UO_605 (O_605,N_9132,N_8749);
xor UO_606 (O_606,N_9700,N_8503);
or UO_607 (O_607,N_9301,N_9672);
and UO_608 (O_608,N_9686,N_8649);
nand UO_609 (O_609,N_9889,N_9152);
nand UO_610 (O_610,N_9200,N_8767);
or UO_611 (O_611,N_8987,N_8570);
or UO_612 (O_612,N_9942,N_9214);
or UO_613 (O_613,N_8457,N_8766);
nand UO_614 (O_614,N_8268,N_8885);
nand UO_615 (O_615,N_9192,N_9380);
xor UO_616 (O_616,N_9451,N_8719);
xor UO_617 (O_617,N_9760,N_8163);
or UO_618 (O_618,N_8533,N_8450);
nor UO_619 (O_619,N_8590,N_9436);
nand UO_620 (O_620,N_8423,N_8364);
and UO_621 (O_621,N_9421,N_9533);
xnor UO_622 (O_622,N_9783,N_9515);
and UO_623 (O_623,N_8536,N_8652);
xor UO_624 (O_624,N_9570,N_9673);
and UO_625 (O_625,N_9151,N_9097);
nand UO_626 (O_626,N_9952,N_8643);
xnor UO_627 (O_627,N_8618,N_9171);
or UO_628 (O_628,N_8154,N_8040);
nand UO_629 (O_629,N_8031,N_8140);
or UO_630 (O_630,N_9268,N_8605);
or UO_631 (O_631,N_8005,N_9309);
nand UO_632 (O_632,N_9229,N_8258);
xnor UO_633 (O_633,N_8661,N_8294);
and UO_634 (O_634,N_8189,N_9894);
nand UO_635 (O_635,N_8362,N_9754);
xnor UO_636 (O_636,N_8434,N_8324);
nor UO_637 (O_637,N_9622,N_9772);
or UO_638 (O_638,N_9859,N_8001);
nor UO_639 (O_639,N_9717,N_8080);
xnor UO_640 (O_640,N_8986,N_8144);
nand UO_641 (O_641,N_9397,N_9978);
nand UO_642 (O_642,N_8346,N_9485);
nand UO_643 (O_643,N_8703,N_9975);
nor UO_644 (O_644,N_9976,N_9752);
or UO_645 (O_645,N_8066,N_8630);
nand UO_646 (O_646,N_9047,N_9513);
and UO_647 (O_647,N_8773,N_8537);
or UO_648 (O_648,N_8157,N_9453);
nand UO_649 (O_649,N_9583,N_9973);
and UO_650 (O_650,N_8520,N_9909);
nand UO_651 (O_651,N_8608,N_8333);
or UO_652 (O_652,N_8199,N_8761);
nand UO_653 (O_653,N_9809,N_9582);
nand UO_654 (O_654,N_9344,N_8695);
and UO_655 (O_655,N_8650,N_8243);
xnor UO_656 (O_656,N_8539,N_8111);
xnor UO_657 (O_657,N_8245,N_9227);
and UO_658 (O_658,N_9424,N_8789);
nand UO_659 (O_659,N_8834,N_8626);
nor UO_660 (O_660,N_8637,N_9780);
xnor UO_661 (O_661,N_9678,N_8743);
and UO_662 (O_662,N_8708,N_8776);
or UO_663 (O_663,N_9585,N_9297);
xnor UO_664 (O_664,N_9204,N_8164);
xor UO_665 (O_665,N_9287,N_9931);
nand UO_666 (O_666,N_8147,N_8221);
or UO_667 (O_667,N_8170,N_8799);
and UO_668 (O_668,N_8206,N_9235);
xnor UO_669 (O_669,N_8688,N_9101);
nand UO_670 (O_670,N_9777,N_8988);
nor UO_671 (O_671,N_9705,N_9002);
xor UO_672 (O_672,N_9445,N_9714);
and UO_673 (O_673,N_9351,N_8002);
or UO_674 (O_674,N_9954,N_8104);
or UO_675 (O_675,N_8191,N_8572);
and UO_676 (O_676,N_9813,N_8900);
nand UO_677 (O_677,N_8003,N_8312);
xnor UO_678 (O_678,N_8797,N_8983);
nor UO_679 (O_679,N_8904,N_9422);
xnor UO_680 (O_680,N_8580,N_8629);
xnor UO_681 (O_681,N_8357,N_9038);
nor UO_682 (O_682,N_9059,N_8358);
nand UO_683 (O_683,N_9719,N_9405);
nor UO_684 (O_684,N_8718,N_9232);
and UO_685 (O_685,N_8507,N_9339);
nand UO_686 (O_686,N_9055,N_8844);
nor UO_687 (O_687,N_8874,N_9910);
or UO_688 (O_688,N_9922,N_8022);
and UO_689 (O_689,N_9637,N_9579);
nand UO_690 (O_690,N_8843,N_9918);
xnor UO_691 (O_691,N_8322,N_8302);
nor UO_692 (O_692,N_9180,N_9966);
xnor UO_693 (O_693,N_9537,N_8449);
and UO_694 (O_694,N_9886,N_8229);
xor UO_695 (O_695,N_9962,N_8596);
nand UO_696 (O_696,N_8575,N_9221);
nor UO_697 (O_697,N_9989,N_8414);
nor UO_698 (O_698,N_8574,N_8410);
or UO_699 (O_699,N_8094,N_9104);
nand UO_700 (O_700,N_8908,N_8088);
nor UO_701 (O_701,N_8677,N_8249);
and UO_702 (O_702,N_8015,N_9147);
and UO_703 (O_703,N_9438,N_8729);
and UO_704 (O_704,N_8047,N_8079);
nor UO_705 (O_705,N_9335,N_9605);
xnor UO_706 (O_706,N_9611,N_9868);
or UO_707 (O_707,N_9815,N_8807);
and UO_708 (O_708,N_9702,N_8599);
and UO_709 (O_709,N_8592,N_8468);
nor UO_710 (O_710,N_9564,N_9732);
nand UO_711 (O_711,N_8133,N_8330);
nor UO_712 (O_712,N_8600,N_9830);
and UO_713 (O_713,N_8976,N_9974);
or UO_714 (O_714,N_9820,N_8667);
nor UO_715 (O_715,N_9122,N_9418);
or UO_716 (O_716,N_9222,N_9128);
and UO_717 (O_717,N_8628,N_9260);
xor UO_718 (O_718,N_9206,N_8730);
nand UO_719 (O_719,N_8639,N_8237);
nand UO_720 (O_720,N_9368,N_9829);
nor UO_721 (O_721,N_9817,N_9314);
and UO_722 (O_722,N_8183,N_9810);
xor UO_723 (O_723,N_9636,N_8825);
and UO_724 (O_724,N_8792,N_9026);
nand UO_725 (O_725,N_9253,N_8228);
nand UO_726 (O_726,N_9936,N_8835);
nand UO_727 (O_727,N_8876,N_9361);
and UO_728 (O_728,N_8155,N_9766);
and UO_729 (O_729,N_8826,N_9866);
or UO_730 (O_730,N_9263,N_9198);
nor UO_731 (O_731,N_8172,N_9552);
nand UO_732 (O_732,N_9998,N_9053);
nand UO_733 (O_733,N_8752,N_8298);
and UO_734 (O_734,N_9517,N_8669);
nand UO_735 (O_735,N_8775,N_8551);
nand UO_736 (O_736,N_8846,N_8431);
nor UO_737 (O_737,N_9689,N_9657);
nand UO_738 (O_738,N_8733,N_8751);
nand UO_739 (O_739,N_9298,N_9331);
or UO_740 (O_740,N_8579,N_8997);
nor UO_741 (O_741,N_9940,N_9238);
xnor UO_742 (O_742,N_9230,N_9647);
xnor UO_743 (O_743,N_9884,N_9215);
and UO_744 (O_744,N_8338,N_9550);
or UO_745 (O_745,N_9990,N_9819);
nor UO_746 (O_746,N_9233,N_8985);
or UO_747 (O_747,N_8319,N_9137);
nor UO_748 (O_748,N_9703,N_9677);
and UO_749 (O_749,N_8704,N_8181);
xor UO_750 (O_750,N_8832,N_8072);
nor UO_751 (O_751,N_9022,N_8909);
nor UO_752 (O_752,N_9949,N_8136);
xnor UO_753 (O_753,N_8389,N_8698);
nor UO_754 (O_754,N_9434,N_8944);
xor UO_755 (O_755,N_8343,N_8745);
nor UO_756 (O_756,N_8796,N_8850);
nand UO_757 (O_757,N_9311,N_9033);
nand UO_758 (O_758,N_9510,N_8691);
xnor UO_759 (O_759,N_9659,N_8396);
and UO_760 (O_760,N_9997,N_9387);
and UO_761 (O_761,N_8803,N_8355);
xnor UO_762 (O_762,N_8073,N_8670);
nand UO_763 (O_763,N_9747,N_8444);
or UO_764 (O_764,N_8542,N_8955);
xnor UO_765 (O_765,N_8401,N_8640);
or UO_766 (O_766,N_8032,N_8101);
or UO_767 (O_767,N_8092,N_8732);
nor UO_768 (O_768,N_8046,N_8953);
nor UO_769 (O_769,N_9707,N_9929);
xnor UO_770 (O_770,N_8619,N_8739);
and UO_771 (O_771,N_9160,N_9291);
and UO_772 (O_772,N_8307,N_9224);
or UO_773 (O_773,N_8809,N_9724);
xnor UO_774 (O_774,N_8486,N_9900);
nand UO_775 (O_775,N_9371,N_9201);
nor UO_776 (O_776,N_9768,N_8017);
nand UO_777 (O_777,N_8636,N_9360);
nand UO_778 (O_778,N_8981,N_8996);
and UO_779 (O_779,N_8911,N_8553);
nor UO_780 (O_780,N_9120,N_9057);
xnor UO_781 (O_781,N_8482,N_8756);
nand UO_782 (O_782,N_9003,N_9278);
and UO_783 (O_783,N_9959,N_9208);
nand UO_784 (O_784,N_8895,N_8951);
nor UO_785 (O_785,N_8152,N_8725);
and UO_786 (O_786,N_9710,N_8671);
or UO_787 (O_787,N_8827,N_9142);
or UO_788 (O_788,N_9333,N_9444);
or UO_789 (O_789,N_9963,N_8461);
or UO_790 (O_790,N_8534,N_9835);
nand UO_791 (O_791,N_9242,N_9203);
and UO_792 (O_792,N_9556,N_8931);
or UO_793 (O_793,N_8038,N_9231);
nor UO_794 (O_794,N_9941,N_8385);
nor UO_795 (O_795,N_9576,N_9354);
nand UO_796 (O_796,N_9251,N_8391);
and UO_797 (O_797,N_8176,N_8559);
or UO_798 (O_798,N_9008,N_9480);
and UO_799 (O_799,N_9862,N_9598);
and UO_800 (O_800,N_8185,N_8056);
nor UO_801 (O_801,N_9063,N_8968);
xnor UO_802 (O_802,N_8087,N_9790);
xnor UO_803 (O_803,N_8439,N_9058);
xnor UO_804 (O_804,N_8403,N_9363);
and UO_805 (O_805,N_8246,N_8230);
xor UO_806 (O_806,N_9932,N_8801);
and UO_807 (O_807,N_8763,N_9548);
and UO_808 (O_808,N_9414,N_8501);
xor UO_809 (O_809,N_9559,N_8769);
and UO_810 (O_810,N_8962,N_9827);
nor UO_811 (O_811,N_9072,N_8787);
xnor UO_812 (O_812,N_8204,N_8464);
nand UO_813 (O_813,N_9872,N_8062);
nor UO_814 (O_814,N_9549,N_8492);
nand UO_815 (O_815,N_9733,N_8452);
and UO_816 (O_816,N_8693,N_8119);
or UO_817 (O_817,N_9357,N_9056);
nand UO_818 (O_818,N_8371,N_8409);
nor UO_819 (O_819,N_8780,N_9299);
nor UO_820 (O_820,N_9666,N_9237);
or UO_821 (O_821,N_8474,N_8938);
or UO_822 (O_822,N_8555,N_9273);
xnor UO_823 (O_823,N_9858,N_9642);
and UO_824 (O_824,N_8044,N_8408);
nand UO_825 (O_825,N_8395,N_8847);
xor UO_826 (O_826,N_8772,N_9327);
and UO_827 (O_827,N_8977,N_9125);
nand UO_828 (O_828,N_8631,N_9701);
or UO_829 (O_829,N_9261,N_8873);
xor UO_830 (O_830,N_9669,N_9631);
nand UO_831 (O_831,N_8188,N_8415);
or UO_832 (O_832,N_8413,N_9863);
or UO_833 (O_833,N_8550,N_8945);
xor UO_834 (O_834,N_9123,N_9801);
or UO_835 (O_835,N_9547,N_9175);
or UO_836 (O_836,N_9226,N_9811);
nor UO_837 (O_837,N_8438,N_9531);
or UO_838 (O_838,N_8231,N_8382);
and UO_839 (O_839,N_8496,N_9588);
nor UO_840 (O_840,N_8526,N_9739);
nor UO_841 (O_841,N_8262,N_9250);
xor UO_842 (O_842,N_8965,N_9681);
xnor UO_843 (O_843,N_9111,N_9950);
nand UO_844 (O_844,N_9560,N_8386);
nand UO_845 (O_845,N_8886,N_9828);
xnor UO_846 (O_846,N_8736,N_9456);
nand UO_847 (O_847,N_9428,N_8311);
nor UO_848 (O_848,N_9202,N_9893);
nor UO_849 (O_849,N_8516,N_9818);
and UO_850 (O_850,N_8380,N_9145);
or UO_851 (O_851,N_8817,N_9953);
nand UO_852 (O_852,N_9305,N_9007);
nand UO_853 (O_853,N_8554,N_8754);
nand UO_854 (O_854,N_8823,N_9541);
and UO_855 (O_855,N_9878,N_8881);
nand UO_856 (O_856,N_9461,N_8960);
and UO_857 (O_857,N_8441,N_8235);
or UO_858 (O_858,N_8342,N_8861);
nand UO_859 (O_859,N_9082,N_8127);
nor UO_860 (O_860,N_9358,N_8065);
and UO_861 (O_861,N_9073,N_9069);
xnor UO_862 (O_862,N_9430,N_8920);
xnor UO_863 (O_863,N_9785,N_8219);
nand UO_864 (O_864,N_8455,N_8443);
nor UO_865 (O_865,N_8940,N_9124);
nor UO_866 (O_866,N_8053,N_8186);
or UO_867 (O_867,N_9947,N_9532);
nor UO_868 (O_868,N_9982,N_9821);
or UO_869 (O_869,N_8069,N_8771);
xnor UO_870 (O_870,N_8632,N_8489);
and UO_871 (O_871,N_9592,N_8591);
xor UO_872 (O_872,N_9538,N_9943);
nor UO_873 (O_873,N_8429,N_8295);
and UO_874 (O_874,N_9638,N_9770);
nor UO_875 (O_875,N_8309,N_8947);
xnor UO_876 (O_876,N_9479,N_8016);
nor UO_877 (O_877,N_9141,N_9439);
and UO_878 (O_878,N_8830,N_8918);
xor UO_879 (O_879,N_9239,N_8010);
or UO_880 (O_880,N_8849,N_8682);
xor UO_881 (O_881,N_8597,N_9144);
or UO_882 (O_882,N_9472,N_8247);
nand UO_883 (O_883,N_8747,N_8182);
nand UO_884 (O_884,N_9944,N_8939);
xor UO_885 (O_885,N_9608,N_9489);
nand UO_886 (O_886,N_9964,N_9381);
and UO_887 (O_887,N_8645,N_9574);
xor UO_888 (O_888,N_8344,N_9409);
xnor UO_889 (O_889,N_8134,N_9345);
or UO_890 (O_890,N_9131,N_8683);
nand UO_891 (O_891,N_9223,N_9646);
xnor UO_892 (O_892,N_8498,N_9146);
nor UO_893 (O_893,N_9979,N_9257);
and UO_894 (O_894,N_8361,N_8813);
xnor UO_895 (O_895,N_8806,N_9185);
nor UO_896 (O_896,N_8076,N_8275);
or UO_897 (O_897,N_8822,N_9389);
xor UO_898 (O_898,N_8561,N_9800);
or UO_899 (O_899,N_9168,N_9740);
nand UO_900 (O_900,N_9065,N_9092);
nor UO_901 (O_901,N_8480,N_9814);
nand UO_902 (O_902,N_9774,N_9484);
or UO_903 (O_903,N_8068,N_9119);
nand UO_904 (O_904,N_8197,N_9904);
and UO_905 (O_905,N_8272,N_8952);
nor UO_906 (O_906,N_8543,N_8504);
nor UO_907 (O_907,N_8781,N_8647);
and UO_908 (O_908,N_8060,N_9749);
and UO_909 (O_909,N_8288,N_8071);
and UO_910 (O_910,N_9153,N_9500);
nand UO_911 (O_911,N_8105,N_9969);
and UO_912 (O_912,N_8768,N_8515);
and UO_913 (O_913,N_9837,N_8098);
nand UO_914 (O_914,N_8325,N_8491);
and UO_915 (O_915,N_8100,N_9844);
or UO_916 (O_916,N_9937,N_9793);
or UO_917 (O_917,N_8980,N_9334);
nor UO_918 (O_918,N_8648,N_9600);
xor UO_919 (O_919,N_9885,N_8664);
or UO_920 (O_920,N_9379,N_8242);
nor UO_921 (O_921,N_8470,N_9655);
nand UO_922 (O_922,N_8853,N_8472);
and UO_923 (O_923,N_8680,N_9839);
nand UO_924 (O_924,N_9482,N_9613);
xnor UO_925 (O_925,N_9465,N_9896);
xnor UO_926 (O_926,N_8720,N_9464);
or UO_927 (O_927,N_8359,N_9735);
xnor UO_928 (O_928,N_8877,N_9195);
xor UO_929 (O_929,N_9606,N_8054);
and UO_930 (O_930,N_8716,N_8132);
nor UO_931 (O_931,N_9317,N_8315);
nand UO_932 (O_932,N_8601,N_9788);
or UO_933 (O_933,N_8332,N_9845);
xnor UO_934 (O_934,N_9271,N_9727);
xnor UO_935 (O_935,N_9743,N_8266);
nand UO_936 (O_936,N_9094,N_8538);
nand UO_937 (O_937,N_9505,N_9694);
xnor UO_938 (O_938,N_8802,N_9925);
xor UO_939 (O_939,N_8138,N_9755);
and UO_940 (O_940,N_8238,N_8090);
xor UO_941 (O_941,N_9347,N_8029);
and UO_942 (O_942,N_9823,N_8153);
xnor UO_943 (O_943,N_9362,N_9062);
and UO_944 (O_944,N_8112,N_9565);
nand UO_945 (O_945,N_8656,N_9386);
and UO_946 (O_946,N_9134,N_8372);
nor UO_947 (O_947,N_9182,N_8845);
xnor UO_948 (O_948,N_8871,N_9902);
and UO_949 (O_949,N_8171,N_9763);
nand UO_950 (O_950,N_9332,N_9286);
nand UO_951 (O_951,N_9881,N_8995);
nand UO_952 (O_952,N_9307,N_9093);
or UO_953 (O_953,N_9306,N_8557);
nor UO_954 (O_954,N_8384,N_9061);
and UO_955 (O_955,N_8917,N_9615);
nand UO_956 (O_956,N_8259,N_8509);
xor UO_957 (O_957,N_9437,N_9708);
nor UO_958 (O_958,N_8037,N_9709);
and UO_959 (O_959,N_8177,N_8528);
xnor UO_960 (O_960,N_9066,N_8659);
and UO_961 (O_961,N_9115,N_8117);
nor UO_962 (O_962,N_8099,N_8982);
nand UO_963 (O_963,N_8946,N_9350);
nor UO_964 (O_964,N_9000,N_8512);
and UO_965 (O_965,N_8706,N_8377);
xor UO_966 (O_966,N_8193,N_8451);
nor UO_967 (O_967,N_9993,N_8446);
and UO_968 (O_968,N_9256,N_9001);
nor UO_969 (O_969,N_9020,N_9848);
xnor UO_970 (O_970,N_9518,N_8547);
xor UO_971 (O_971,N_9177,N_8709);
nand UO_972 (O_972,N_8970,N_8203);
or UO_973 (O_973,N_9731,N_8594);
nand UO_974 (O_974,N_8304,N_8828);
or UO_975 (O_975,N_9847,N_9078);
nand UO_976 (O_976,N_9948,N_9665);
xnor UO_977 (O_977,N_9854,N_8923);
xnor UO_978 (O_978,N_8907,N_8210);
nor UO_979 (O_979,N_8744,N_9806);
nand UO_980 (O_980,N_8167,N_9728);
xnor UO_981 (O_981,N_8856,N_8327);
and UO_982 (O_982,N_9255,N_8746);
nand UO_983 (O_983,N_9486,N_9633);
and UO_984 (O_984,N_8869,N_9296);
nor UO_985 (O_985,N_9601,N_8914);
nand UO_986 (O_986,N_8783,N_9448);
and UO_987 (O_987,N_8779,N_8936);
xor UO_988 (O_988,N_8399,N_9040);
xnor UO_989 (O_989,N_9030,N_9019);
xor UO_990 (O_990,N_9391,N_9402);
nand UO_991 (O_991,N_9322,N_9796);
nand UO_992 (O_992,N_8131,N_8476);
xnor UO_993 (O_993,N_9415,N_9664);
or UO_994 (O_994,N_8348,N_9283);
xnor UO_995 (O_995,N_9972,N_8271);
xnor UO_996 (O_996,N_8857,N_9281);
and UO_997 (O_997,N_8146,N_9967);
xnor UO_998 (O_998,N_9244,N_9212);
nand UO_999 (O_999,N_9187,N_8121);
and UO_1000 (O_1000,N_8951,N_9064);
xnor UO_1001 (O_1001,N_8782,N_9077);
or UO_1002 (O_1002,N_9999,N_9666);
xor UO_1003 (O_1003,N_9977,N_8233);
and UO_1004 (O_1004,N_8995,N_9065);
or UO_1005 (O_1005,N_9101,N_8321);
nand UO_1006 (O_1006,N_8788,N_8408);
or UO_1007 (O_1007,N_8977,N_8539);
and UO_1008 (O_1008,N_8207,N_8783);
xnor UO_1009 (O_1009,N_8506,N_8103);
nand UO_1010 (O_1010,N_8591,N_9503);
nor UO_1011 (O_1011,N_9333,N_9376);
or UO_1012 (O_1012,N_8013,N_9394);
and UO_1013 (O_1013,N_8113,N_9708);
and UO_1014 (O_1014,N_8511,N_8013);
xor UO_1015 (O_1015,N_8732,N_8741);
nor UO_1016 (O_1016,N_9471,N_8447);
nor UO_1017 (O_1017,N_9569,N_8008);
nand UO_1018 (O_1018,N_8863,N_9662);
and UO_1019 (O_1019,N_8777,N_9927);
xor UO_1020 (O_1020,N_9894,N_9085);
nor UO_1021 (O_1021,N_8960,N_8507);
nor UO_1022 (O_1022,N_8035,N_9242);
or UO_1023 (O_1023,N_8472,N_8670);
nand UO_1024 (O_1024,N_8706,N_9650);
and UO_1025 (O_1025,N_9179,N_8926);
or UO_1026 (O_1026,N_8192,N_8090);
nor UO_1027 (O_1027,N_9999,N_9026);
nand UO_1028 (O_1028,N_9389,N_8625);
nor UO_1029 (O_1029,N_8186,N_9017);
nand UO_1030 (O_1030,N_9493,N_9689);
and UO_1031 (O_1031,N_8580,N_9555);
xnor UO_1032 (O_1032,N_9858,N_8728);
xnor UO_1033 (O_1033,N_9156,N_9861);
xor UO_1034 (O_1034,N_9170,N_9877);
xor UO_1035 (O_1035,N_9050,N_9080);
or UO_1036 (O_1036,N_8149,N_9060);
or UO_1037 (O_1037,N_8558,N_8814);
nor UO_1038 (O_1038,N_8914,N_9246);
nand UO_1039 (O_1039,N_9343,N_9150);
and UO_1040 (O_1040,N_9871,N_9958);
or UO_1041 (O_1041,N_8480,N_9865);
nand UO_1042 (O_1042,N_8610,N_8493);
nand UO_1043 (O_1043,N_8839,N_8627);
xor UO_1044 (O_1044,N_9594,N_8978);
or UO_1045 (O_1045,N_8844,N_9770);
xor UO_1046 (O_1046,N_8432,N_8797);
nor UO_1047 (O_1047,N_8807,N_9680);
nor UO_1048 (O_1048,N_9633,N_9407);
and UO_1049 (O_1049,N_8686,N_9943);
nor UO_1050 (O_1050,N_9841,N_9174);
and UO_1051 (O_1051,N_8697,N_8130);
nor UO_1052 (O_1052,N_8293,N_8631);
nand UO_1053 (O_1053,N_8440,N_9141);
nor UO_1054 (O_1054,N_9954,N_8195);
and UO_1055 (O_1055,N_8122,N_9429);
nor UO_1056 (O_1056,N_8668,N_8423);
nand UO_1057 (O_1057,N_9659,N_8092);
nand UO_1058 (O_1058,N_9794,N_8787);
or UO_1059 (O_1059,N_8763,N_8928);
nor UO_1060 (O_1060,N_9684,N_9867);
xor UO_1061 (O_1061,N_8715,N_9525);
nand UO_1062 (O_1062,N_9700,N_8076);
and UO_1063 (O_1063,N_9169,N_9597);
xnor UO_1064 (O_1064,N_9763,N_8744);
and UO_1065 (O_1065,N_8083,N_8254);
and UO_1066 (O_1066,N_8493,N_8620);
nand UO_1067 (O_1067,N_8183,N_9259);
and UO_1068 (O_1068,N_9777,N_8153);
nor UO_1069 (O_1069,N_9417,N_9425);
and UO_1070 (O_1070,N_8330,N_8836);
or UO_1071 (O_1071,N_8298,N_8556);
nand UO_1072 (O_1072,N_9021,N_8019);
and UO_1073 (O_1073,N_9635,N_9640);
nand UO_1074 (O_1074,N_9550,N_8001);
and UO_1075 (O_1075,N_8554,N_9193);
and UO_1076 (O_1076,N_9345,N_9273);
or UO_1077 (O_1077,N_8932,N_9575);
xnor UO_1078 (O_1078,N_9453,N_8446);
or UO_1079 (O_1079,N_8012,N_8857);
xnor UO_1080 (O_1080,N_9309,N_8244);
or UO_1081 (O_1081,N_9147,N_9175);
nand UO_1082 (O_1082,N_9973,N_9449);
nand UO_1083 (O_1083,N_8628,N_8526);
or UO_1084 (O_1084,N_9754,N_9235);
nand UO_1085 (O_1085,N_9317,N_8763);
and UO_1086 (O_1086,N_9312,N_8058);
and UO_1087 (O_1087,N_9393,N_8107);
or UO_1088 (O_1088,N_8664,N_9706);
or UO_1089 (O_1089,N_9583,N_8689);
xor UO_1090 (O_1090,N_9631,N_8038);
nand UO_1091 (O_1091,N_8504,N_9821);
nand UO_1092 (O_1092,N_9374,N_8387);
or UO_1093 (O_1093,N_9173,N_9267);
xor UO_1094 (O_1094,N_9799,N_8120);
and UO_1095 (O_1095,N_9667,N_9863);
or UO_1096 (O_1096,N_9541,N_9986);
xor UO_1097 (O_1097,N_8722,N_8048);
nand UO_1098 (O_1098,N_9863,N_8391);
xor UO_1099 (O_1099,N_8314,N_9444);
and UO_1100 (O_1100,N_9705,N_8177);
xor UO_1101 (O_1101,N_9250,N_8737);
and UO_1102 (O_1102,N_9628,N_9057);
nor UO_1103 (O_1103,N_9339,N_9455);
xor UO_1104 (O_1104,N_9067,N_9765);
and UO_1105 (O_1105,N_8587,N_8420);
or UO_1106 (O_1106,N_8919,N_9858);
nor UO_1107 (O_1107,N_9161,N_8408);
xnor UO_1108 (O_1108,N_8510,N_8279);
nand UO_1109 (O_1109,N_9060,N_8626);
nor UO_1110 (O_1110,N_9925,N_8365);
nand UO_1111 (O_1111,N_8899,N_9166);
nor UO_1112 (O_1112,N_8339,N_9827);
xor UO_1113 (O_1113,N_9203,N_9443);
nor UO_1114 (O_1114,N_8513,N_8049);
and UO_1115 (O_1115,N_9075,N_8408);
or UO_1116 (O_1116,N_9562,N_9556);
and UO_1117 (O_1117,N_8841,N_9031);
nor UO_1118 (O_1118,N_8563,N_8566);
xor UO_1119 (O_1119,N_9903,N_9737);
and UO_1120 (O_1120,N_8398,N_9258);
or UO_1121 (O_1121,N_8235,N_8799);
and UO_1122 (O_1122,N_9140,N_9844);
nor UO_1123 (O_1123,N_8460,N_8583);
and UO_1124 (O_1124,N_8114,N_9510);
xnor UO_1125 (O_1125,N_8511,N_8422);
and UO_1126 (O_1126,N_8452,N_9828);
or UO_1127 (O_1127,N_8434,N_9796);
and UO_1128 (O_1128,N_9592,N_9254);
nand UO_1129 (O_1129,N_8043,N_9473);
xor UO_1130 (O_1130,N_9213,N_8606);
nand UO_1131 (O_1131,N_8935,N_9858);
xnor UO_1132 (O_1132,N_8189,N_8470);
and UO_1133 (O_1133,N_8326,N_9975);
and UO_1134 (O_1134,N_8895,N_9152);
nand UO_1135 (O_1135,N_8973,N_9888);
nand UO_1136 (O_1136,N_9642,N_9088);
nand UO_1137 (O_1137,N_8848,N_8634);
nor UO_1138 (O_1138,N_9418,N_9915);
or UO_1139 (O_1139,N_8705,N_8489);
and UO_1140 (O_1140,N_9340,N_9688);
nand UO_1141 (O_1141,N_9260,N_9606);
or UO_1142 (O_1142,N_8317,N_9475);
nor UO_1143 (O_1143,N_8153,N_8614);
xnor UO_1144 (O_1144,N_9523,N_9293);
nor UO_1145 (O_1145,N_9516,N_8351);
and UO_1146 (O_1146,N_9699,N_8000);
nand UO_1147 (O_1147,N_8161,N_8945);
nor UO_1148 (O_1148,N_9489,N_8882);
xnor UO_1149 (O_1149,N_8786,N_8602);
or UO_1150 (O_1150,N_9417,N_9520);
nand UO_1151 (O_1151,N_9984,N_9390);
nor UO_1152 (O_1152,N_9036,N_8815);
nor UO_1153 (O_1153,N_8341,N_9423);
nand UO_1154 (O_1154,N_9849,N_8317);
and UO_1155 (O_1155,N_8869,N_8251);
nand UO_1156 (O_1156,N_8333,N_9820);
nand UO_1157 (O_1157,N_9590,N_9697);
nand UO_1158 (O_1158,N_8136,N_9118);
and UO_1159 (O_1159,N_8327,N_8893);
xnor UO_1160 (O_1160,N_8245,N_9993);
xnor UO_1161 (O_1161,N_8663,N_9396);
nor UO_1162 (O_1162,N_8611,N_8267);
or UO_1163 (O_1163,N_9418,N_8151);
or UO_1164 (O_1164,N_9206,N_9433);
or UO_1165 (O_1165,N_8836,N_8443);
and UO_1166 (O_1166,N_8033,N_8496);
nor UO_1167 (O_1167,N_9404,N_8476);
nand UO_1168 (O_1168,N_8304,N_9282);
or UO_1169 (O_1169,N_8074,N_9452);
xnor UO_1170 (O_1170,N_8286,N_8246);
nand UO_1171 (O_1171,N_8730,N_9365);
xnor UO_1172 (O_1172,N_8190,N_9041);
or UO_1173 (O_1173,N_8547,N_8487);
and UO_1174 (O_1174,N_9886,N_9230);
or UO_1175 (O_1175,N_9104,N_8939);
xor UO_1176 (O_1176,N_8796,N_9160);
and UO_1177 (O_1177,N_9961,N_9112);
or UO_1178 (O_1178,N_8583,N_9370);
xnor UO_1179 (O_1179,N_9912,N_9671);
xor UO_1180 (O_1180,N_8923,N_9632);
and UO_1181 (O_1181,N_8390,N_9731);
nand UO_1182 (O_1182,N_9607,N_8165);
xnor UO_1183 (O_1183,N_8383,N_9576);
nand UO_1184 (O_1184,N_9885,N_8810);
or UO_1185 (O_1185,N_9764,N_9705);
nand UO_1186 (O_1186,N_8441,N_8287);
nor UO_1187 (O_1187,N_9912,N_9838);
nand UO_1188 (O_1188,N_9338,N_9987);
and UO_1189 (O_1189,N_9865,N_9996);
nand UO_1190 (O_1190,N_9217,N_8221);
nand UO_1191 (O_1191,N_9049,N_8129);
and UO_1192 (O_1192,N_8333,N_8241);
or UO_1193 (O_1193,N_9402,N_9425);
nor UO_1194 (O_1194,N_8261,N_9545);
or UO_1195 (O_1195,N_8144,N_9711);
xor UO_1196 (O_1196,N_8533,N_9226);
xnor UO_1197 (O_1197,N_8683,N_8785);
and UO_1198 (O_1198,N_9534,N_8590);
xor UO_1199 (O_1199,N_9226,N_9392);
or UO_1200 (O_1200,N_9957,N_8027);
nand UO_1201 (O_1201,N_8214,N_9996);
nor UO_1202 (O_1202,N_9549,N_8999);
xor UO_1203 (O_1203,N_8921,N_8029);
nor UO_1204 (O_1204,N_9762,N_8616);
xor UO_1205 (O_1205,N_9281,N_8661);
nand UO_1206 (O_1206,N_9628,N_8446);
nor UO_1207 (O_1207,N_8145,N_8695);
xor UO_1208 (O_1208,N_9343,N_9720);
xor UO_1209 (O_1209,N_9369,N_8387);
nand UO_1210 (O_1210,N_8913,N_8099);
and UO_1211 (O_1211,N_8986,N_9084);
nand UO_1212 (O_1212,N_9804,N_9491);
nand UO_1213 (O_1213,N_8795,N_9593);
or UO_1214 (O_1214,N_9835,N_8823);
or UO_1215 (O_1215,N_8855,N_9238);
xor UO_1216 (O_1216,N_9989,N_8748);
nor UO_1217 (O_1217,N_8797,N_8082);
nor UO_1218 (O_1218,N_8275,N_8627);
and UO_1219 (O_1219,N_8468,N_8095);
xor UO_1220 (O_1220,N_8857,N_8822);
and UO_1221 (O_1221,N_9041,N_9350);
xnor UO_1222 (O_1222,N_8743,N_9572);
xnor UO_1223 (O_1223,N_9884,N_8337);
nand UO_1224 (O_1224,N_9480,N_8220);
nand UO_1225 (O_1225,N_9323,N_8855);
xnor UO_1226 (O_1226,N_9620,N_8422);
xnor UO_1227 (O_1227,N_9511,N_8281);
xnor UO_1228 (O_1228,N_9170,N_9021);
or UO_1229 (O_1229,N_8915,N_8764);
or UO_1230 (O_1230,N_8771,N_9210);
nor UO_1231 (O_1231,N_9051,N_9351);
nand UO_1232 (O_1232,N_8399,N_9516);
xor UO_1233 (O_1233,N_9988,N_8507);
nor UO_1234 (O_1234,N_9611,N_9472);
xor UO_1235 (O_1235,N_8819,N_9860);
and UO_1236 (O_1236,N_8649,N_8143);
xor UO_1237 (O_1237,N_8272,N_8346);
nand UO_1238 (O_1238,N_9222,N_9587);
nor UO_1239 (O_1239,N_8483,N_8115);
nor UO_1240 (O_1240,N_8843,N_9735);
nor UO_1241 (O_1241,N_8144,N_8685);
nand UO_1242 (O_1242,N_9473,N_8884);
nor UO_1243 (O_1243,N_8213,N_8307);
and UO_1244 (O_1244,N_9847,N_9366);
xnor UO_1245 (O_1245,N_9625,N_8851);
nor UO_1246 (O_1246,N_8258,N_9944);
and UO_1247 (O_1247,N_8746,N_9505);
or UO_1248 (O_1248,N_8979,N_8748);
or UO_1249 (O_1249,N_8778,N_8525);
and UO_1250 (O_1250,N_9658,N_9656);
or UO_1251 (O_1251,N_8769,N_8624);
xnor UO_1252 (O_1252,N_9713,N_8968);
or UO_1253 (O_1253,N_8484,N_8817);
nor UO_1254 (O_1254,N_9706,N_9454);
or UO_1255 (O_1255,N_9584,N_9796);
or UO_1256 (O_1256,N_8486,N_8351);
or UO_1257 (O_1257,N_9332,N_8378);
nand UO_1258 (O_1258,N_8229,N_9226);
and UO_1259 (O_1259,N_8142,N_9812);
xor UO_1260 (O_1260,N_9927,N_8914);
or UO_1261 (O_1261,N_8186,N_8312);
nor UO_1262 (O_1262,N_9201,N_8382);
nand UO_1263 (O_1263,N_9961,N_9972);
or UO_1264 (O_1264,N_8704,N_8479);
and UO_1265 (O_1265,N_9228,N_8014);
and UO_1266 (O_1266,N_8332,N_9451);
or UO_1267 (O_1267,N_9998,N_8269);
nand UO_1268 (O_1268,N_8467,N_9918);
xor UO_1269 (O_1269,N_9511,N_8342);
nand UO_1270 (O_1270,N_9377,N_9603);
xor UO_1271 (O_1271,N_8497,N_8002);
nand UO_1272 (O_1272,N_8808,N_9992);
nor UO_1273 (O_1273,N_9933,N_8355);
and UO_1274 (O_1274,N_8052,N_8134);
or UO_1275 (O_1275,N_8978,N_8645);
nor UO_1276 (O_1276,N_9825,N_8025);
nand UO_1277 (O_1277,N_9586,N_8333);
nor UO_1278 (O_1278,N_9724,N_9161);
nand UO_1279 (O_1279,N_8884,N_8259);
xor UO_1280 (O_1280,N_9069,N_8980);
or UO_1281 (O_1281,N_8612,N_8842);
xor UO_1282 (O_1282,N_8027,N_8217);
nor UO_1283 (O_1283,N_9061,N_8437);
and UO_1284 (O_1284,N_9848,N_9636);
nor UO_1285 (O_1285,N_9808,N_9089);
and UO_1286 (O_1286,N_8288,N_9677);
or UO_1287 (O_1287,N_9388,N_8441);
nand UO_1288 (O_1288,N_8800,N_9325);
xor UO_1289 (O_1289,N_8679,N_8220);
nand UO_1290 (O_1290,N_9737,N_9444);
and UO_1291 (O_1291,N_9207,N_9789);
and UO_1292 (O_1292,N_9578,N_8305);
nor UO_1293 (O_1293,N_8208,N_8759);
nand UO_1294 (O_1294,N_9888,N_8363);
xnor UO_1295 (O_1295,N_9544,N_9198);
and UO_1296 (O_1296,N_9122,N_9939);
nand UO_1297 (O_1297,N_9608,N_9126);
xnor UO_1298 (O_1298,N_8445,N_9182);
nand UO_1299 (O_1299,N_8931,N_9910);
nand UO_1300 (O_1300,N_8628,N_9137);
nand UO_1301 (O_1301,N_8381,N_8478);
nor UO_1302 (O_1302,N_8076,N_8258);
nand UO_1303 (O_1303,N_8169,N_8131);
nor UO_1304 (O_1304,N_9018,N_8513);
and UO_1305 (O_1305,N_9057,N_9170);
or UO_1306 (O_1306,N_9569,N_8642);
and UO_1307 (O_1307,N_8458,N_9222);
xnor UO_1308 (O_1308,N_8509,N_8057);
and UO_1309 (O_1309,N_9988,N_9828);
nor UO_1310 (O_1310,N_9010,N_9605);
or UO_1311 (O_1311,N_9027,N_8053);
xor UO_1312 (O_1312,N_8096,N_8391);
and UO_1313 (O_1313,N_9386,N_9780);
and UO_1314 (O_1314,N_9182,N_9361);
and UO_1315 (O_1315,N_9034,N_8620);
and UO_1316 (O_1316,N_9967,N_8596);
nor UO_1317 (O_1317,N_8478,N_8567);
or UO_1318 (O_1318,N_8021,N_8451);
nand UO_1319 (O_1319,N_9095,N_8746);
or UO_1320 (O_1320,N_8984,N_8217);
xnor UO_1321 (O_1321,N_8310,N_8066);
and UO_1322 (O_1322,N_8405,N_8721);
nand UO_1323 (O_1323,N_8451,N_9550);
nor UO_1324 (O_1324,N_9402,N_8890);
and UO_1325 (O_1325,N_9382,N_9173);
nor UO_1326 (O_1326,N_8869,N_9328);
and UO_1327 (O_1327,N_8120,N_9501);
or UO_1328 (O_1328,N_9440,N_9495);
xnor UO_1329 (O_1329,N_9192,N_8044);
nor UO_1330 (O_1330,N_8369,N_8784);
xor UO_1331 (O_1331,N_9930,N_9018);
and UO_1332 (O_1332,N_9345,N_9054);
nor UO_1333 (O_1333,N_8650,N_9056);
or UO_1334 (O_1334,N_9338,N_8915);
nor UO_1335 (O_1335,N_8041,N_8275);
or UO_1336 (O_1336,N_8690,N_9615);
nand UO_1337 (O_1337,N_9917,N_8046);
nand UO_1338 (O_1338,N_8423,N_9594);
nand UO_1339 (O_1339,N_8768,N_9893);
or UO_1340 (O_1340,N_9474,N_8777);
and UO_1341 (O_1341,N_8745,N_9709);
and UO_1342 (O_1342,N_9941,N_9378);
xnor UO_1343 (O_1343,N_8855,N_8036);
nand UO_1344 (O_1344,N_9545,N_9743);
xnor UO_1345 (O_1345,N_8792,N_9493);
nor UO_1346 (O_1346,N_8495,N_8849);
and UO_1347 (O_1347,N_8816,N_8642);
nor UO_1348 (O_1348,N_9428,N_8351);
nor UO_1349 (O_1349,N_9472,N_9163);
and UO_1350 (O_1350,N_9461,N_9540);
or UO_1351 (O_1351,N_9304,N_8928);
nor UO_1352 (O_1352,N_8172,N_8654);
or UO_1353 (O_1353,N_8106,N_9553);
nor UO_1354 (O_1354,N_9608,N_9005);
xor UO_1355 (O_1355,N_9839,N_9021);
nand UO_1356 (O_1356,N_9807,N_9662);
nand UO_1357 (O_1357,N_9125,N_9270);
nand UO_1358 (O_1358,N_9829,N_8433);
or UO_1359 (O_1359,N_9564,N_8126);
nor UO_1360 (O_1360,N_9381,N_8338);
nor UO_1361 (O_1361,N_8372,N_9346);
nand UO_1362 (O_1362,N_8569,N_9005);
and UO_1363 (O_1363,N_9683,N_8977);
nand UO_1364 (O_1364,N_8580,N_9736);
nand UO_1365 (O_1365,N_9274,N_8552);
or UO_1366 (O_1366,N_9295,N_8694);
or UO_1367 (O_1367,N_9398,N_8518);
nor UO_1368 (O_1368,N_9818,N_9454);
xor UO_1369 (O_1369,N_9916,N_9590);
xor UO_1370 (O_1370,N_9320,N_8905);
xnor UO_1371 (O_1371,N_9317,N_8934);
and UO_1372 (O_1372,N_9197,N_8700);
xor UO_1373 (O_1373,N_9119,N_9485);
or UO_1374 (O_1374,N_9207,N_8238);
or UO_1375 (O_1375,N_8030,N_9417);
nand UO_1376 (O_1376,N_8841,N_9062);
nand UO_1377 (O_1377,N_9853,N_8116);
xnor UO_1378 (O_1378,N_9288,N_9258);
and UO_1379 (O_1379,N_9729,N_8030);
or UO_1380 (O_1380,N_8396,N_8581);
nor UO_1381 (O_1381,N_8757,N_8464);
or UO_1382 (O_1382,N_9405,N_8995);
xnor UO_1383 (O_1383,N_9677,N_9422);
nand UO_1384 (O_1384,N_8937,N_9562);
or UO_1385 (O_1385,N_9859,N_9278);
xor UO_1386 (O_1386,N_8207,N_8499);
xnor UO_1387 (O_1387,N_8433,N_8430);
nand UO_1388 (O_1388,N_9250,N_8034);
and UO_1389 (O_1389,N_9723,N_9145);
nand UO_1390 (O_1390,N_8252,N_9029);
xnor UO_1391 (O_1391,N_9539,N_8681);
nand UO_1392 (O_1392,N_9504,N_8187);
xor UO_1393 (O_1393,N_9954,N_9366);
and UO_1394 (O_1394,N_9851,N_9242);
nand UO_1395 (O_1395,N_9222,N_9164);
and UO_1396 (O_1396,N_8476,N_8292);
xor UO_1397 (O_1397,N_8078,N_8332);
nor UO_1398 (O_1398,N_9942,N_8604);
nor UO_1399 (O_1399,N_8713,N_8345);
nor UO_1400 (O_1400,N_9013,N_9155);
xor UO_1401 (O_1401,N_9433,N_8580);
and UO_1402 (O_1402,N_8622,N_8781);
nand UO_1403 (O_1403,N_9925,N_9134);
or UO_1404 (O_1404,N_8410,N_9320);
and UO_1405 (O_1405,N_9746,N_9781);
and UO_1406 (O_1406,N_8160,N_9299);
and UO_1407 (O_1407,N_9942,N_9622);
xor UO_1408 (O_1408,N_8266,N_9198);
nor UO_1409 (O_1409,N_8908,N_8597);
nand UO_1410 (O_1410,N_9992,N_9109);
nor UO_1411 (O_1411,N_9114,N_9222);
nand UO_1412 (O_1412,N_9185,N_8833);
and UO_1413 (O_1413,N_8935,N_8799);
nor UO_1414 (O_1414,N_9777,N_8535);
xor UO_1415 (O_1415,N_8639,N_9842);
or UO_1416 (O_1416,N_9221,N_8406);
or UO_1417 (O_1417,N_9683,N_8172);
nor UO_1418 (O_1418,N_8471,N_8536);
or UO_1419 (O_1419,N_8100,N_9246);
nand UO_1420 (O_1420,N_8300,N_9606);
nand UO_1421 (O_1421,N_8309,N_9551);
nand UO_1422 (O_1422,N_9145,N_9611);
and UO_1423 (O_1423,N_9144,N_8233);
and UO_1424 (O_1424,N_9228,N_8505);
and UO_1425 (O_1425,N_9359,N_8383);
or UO_1426 (O_1426,N_8032,N_9010);
and UO_1427 (O_1427,N_9719,N_9225);
and UO_1428 (O_1428,N_8998,N_8166);
and UO_1429 (O_1429,N_8529,N_9676);
or UO_1430 (O_1430,N_8456,N_9025);
xor UO_1431 (O_1431,N_8163,N_9353);
and UO_1432 (O_1432,N_8605,N_8560);
nand UO_1433 (O_1433,N_8500,N_8323);
or UO_1434 (O_1434,N_9102,N_9873);
nand UO_1435 (O_1435,N_8356,N_9578);
nand UO_1436 (O_1436,N_8431,N_9237);
or UO_1437 (O_1437,N_8268,N_9042);
xor UO_1438 (O_1438,N_9907,N_8760);
nand UO_1439 (O_1439,N_9773,N_8786);
or UO_1440 (O_1440,N_9582,N_8279);
and UO_1441 (O_1441,N_8051,N_8385);
and UO_1442 (O_1442,N_8276,N_8599);
xor UO_1443 (O_1443,N_9420,N_8595);
xor UO_1444 (O_1444,N_8492,N_8143);
and UO_1445 (O_1445,N_8296,N_9726);
xnor UO_1446 (O_1446,N_8604,N_8921);
nor UO_1447 (O_1447,N_8111,N_9882);
nand UO_1448 (O_1448,N_9148,N_8123);
and UO_1449 (O_1449,N_9903,N_8224);
or UO_1450 (O_1450,N_8206,N_8131);
xnor UO_1451 (O_1451,N_9002,N_8123);
and UO_1452 (O_1452,N_9423,N_8729);
nor UO_1453 (O_1453,N_9616,N_8197);
nor UO_1454 (O_1454,N_8968,N_8268);
and UO_1455 (O_1455,N_9012,N_8019);
or UO_1456 (O_1456,N_8037,N_9774);
xor UO_1457 (O_1457,N_9471,N_9767);
xnor UO_1458 (O_1458,N_8115,N_8308);
or UO_1459 (O_1459,N_8099,N_8968);
and UO_1460 (O_1460,N_9744,N_9079);
nand UO_1461 (O_1461,N_8403,N_8088);
and UO_1462 (O_1462,N_9239,N_9108);
or UO_1463 (O_1463,N_8645,N_9734);
and UO_1464 (O_1464,N_8913,N_8004);
and UO_1465 (O_1465,N_9846,N_8329);
and UO_1466 (O_1466,N_8799,N_8836);
or UO_1467 (O_1467,N_9870,N_8732);
nor UO_1468 (O_1468,N_8040,N_9073);
or UO_1469 (O_1469,N_8065,N_9580);
nor UO_1470 (O_1470,N_8760,N_8185);
nand UO_1471 (O_1471,N_8594,N_8194);
and UO_1472 (O_1472,N_9992,N_8468);
nor UO_1473 (O_1473,N_8940,N_9434);
nand UO_1474 (O_1474,N_8948,N_8462);
and UO_1475 (O_1475,N_8483,N_8784);
xnor UO_1476 (O_1476,N_8338,N_8707);
nand UO_1477 (O_1477,N_9190,N_8199);
and UO_1478 (O_1478,N_8014,N_9129);
xor UO_1479 (O_1479,N_9664,N_8297);
nand UO_1480 (O_1480,N_9588,N_9669);
xnor UO_1481 (O_1481,N_8271,N_8471);
xor UO_1482 (O_1482,N_9244,N_9692);
nand UO_1483 (O_1483,N_9511,N_9966);
and UO_1484 (O_1484,N_9844,N_8239);
nor UO_1485 (O_1485,N_8459,N_9425);
nand UO_1486 (O_1486,N_9555,N_9738);
xor UO_1487 (O_1487,N_8726,N_9272);
nand UO_1488 (O_1488,N_8018,N_9436);
or UO_1489 (O_1489,N_9706,N_8498);
nor UO_1490 (O_1490,N_8127,N_8962);
xor UO_1491 (O_1491,N_9396,N_8463);
or UO_1492 (O_1492,N_8378,N_8242);
nor UO_1493 (O_1493,N_9575,N_9050);
xor UO_1494 (O_1494,N_9814,N_8842);
nand UO_1495 (O_1495,N_9896,N_8787);
nor UO_1496 (O_1496,N_8528,N_8233);
and UO_1497 (O_1497,N_8644,N_9550);
and UO_1498 (O_1498,N_9510,N_9807);
nor UO_1499 (O_1499,N_9236,N_8996);
endmodule