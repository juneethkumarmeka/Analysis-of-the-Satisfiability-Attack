module basic_5000_50000_5000_20_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
xnor U0 (N_0,In_3805,In_3823);
xnor U1 (N_1,In_1970,In_3365);
or U2 (N_2,In_2626,In_854);
and U3 (N_3,In_2545,In_3436);
or U4 (N_4,In_2315,In_2783);
and U5 (N_5,In_36,In_1803);
or U6 (N_6,In_4213,In_2933);
nand U7 (N_7,In_79,In_1484);
nand U8 (N_8,In_1254,In_2089);
xnor U9 (N_9,In_356,In_3222);
or U10 (N_10,In_2342,In_1015);
nand U11 (N_11,In_1292,In_2820);
xnor U12 (N_12,In_2020,In_3822);
xnor U13 (N_13,In_4454,In_820);
nor U14 (N_14,In_3173,In_4099);
xnor U15 (N_15,In_376,In_3988);
nand U16 (N_16,In_2531,In_4087);
nor U17 (N_17,In_4408,In_4278);
and U18 (N_18,In_1971,In_2978);
or U19 (N_19,In_4260,In_2344);
or U20 (N_20,In_4244,In_3477);
xor U21 (N_21,In_468,In_2015);
or U22 (N_22,In_4496,In_697);
and U23 (N_23,In_4538,In_3313);
nand U24 (N_24,In_115,In_3569);
nand U25 (N_25,In_2222,In_244);
and U26 (N_26,In_4162,In_371);
nor U27 (N_27,In_3116,In_3568);
or U28 (N_28,In_3931,In_2443);
nand U29 (N_29,In_2209,In_2348);
xor U30 (N_30,In_1533,In_1024);
xnor U31 (N_31,In_2358,In_2335);
and U32 (N_32,In_2511,In_2004);
and U33 (N_33,In_4438,In_1171);
nand U34 (N_34,In_3296,In_2042);
and U35 (N_35,In_3841,In_554);
xor U36 (N_36,In_1119,In_1954);
and U37 (N_37,In_216,In_2182);
nand U38 (N_38,In_4748,In_784);
or U39 (N_39,In_4554,In_4406);
nor U40 (N_40,In_1857,In_24);
nand U41 (N_41,In_2942,In_4614);
and U42 (N_42,In_3530,In_3708);
or U43 (N_43,In_1973,In_2446);
and U44 (N_44,In_373,In_2628);
xor U45 (N_45,In_423,In_3194);
xor U46 (N_46,In_2773,In_4448);
xor U47 (N_47,In_4030,In_3687);
or U48 (N_48,In_4613,In_1231);
nand U49 (N_49,In_3926,In_1674);
and U50 (N_50,In_3873,In_1099);
nor U51 (N_51,In_299,In_1814);
nor U52 (N_52,In_785,In_257);
and U53 (N_53,In_4410,In_4733);
and U54 (N_54,In_4924,In_3730);
xor U55 (N_55,In_2457,In_2958);
and U56 (N_56,In_3628,In_907);
xnor U57 (N_57,In_4096,In_4306);
or U58 (N_58,In_4389,In_2100);
and U59 (N_59,In_4719,In_1017);
xor U60 (N_60,In_4771,In_4794);
nand U61 (N_61,In_1488,In_2075);
and U62 (N_62,In_885,In_4738);
nor U63 (N_63,In_2745,In_3681);
nand U64 (N_64,In_728,In_4744);
nor U65 (N_65,In_3242,In_1772);
and U66 (N_66,In_3092,In_2211);
nand U67 (N_67,In_381,In_2139);
nand U68 (N_68,In_4185,In_2018);
xor U69 (N_69,In_2702,In_1304);
and U70 (N_70,In_4394,In_2821);
or U71 (N_71,In_1398,In_2000);
and U72 (N_72,In_548,In_724);
nor U73 (N_73,In_4941,In_643);
and U74 (N_74,In_131,In_3740);
xnor U75 (N_75,In_3279,In_2035);
or U76 (N_76,In_1957,In_1875);
and U77 (N_77,In_3758,In_876);
xor U78 (N_78,In_734,In_3095);
nand U79 (N_79,In_1356,In_2711);
nand U80 (N_80,In_2596,In_3502);
and U81 (N_81,In_254,In_3744);
or U82 (N_82,In_2259,In_2332);
xor U83 (N_83,In_4460,In_4315);
or U84 (N_84,In_970,In_1877);
and U85 (N_85,In_2538,In_4256);
xor U86 (N_86,In_1681,In_716);
or U87 (N_87,In_936,In_1588);
nand U88 (N_88,In_2402,In_2737);
nand U89 (N_89,In_1438,In_1131);
xnor U90 (N_90,In_2126,In_1281);
nand U91 (N_91,In_2453,In_1520);
nor U92 (N_92,In_4402,In_1262);
xnor U93 (N_93,In_1215,In_3960);
nand U94 (N_94,In_1168,In_105);
or U95 (N_95,In_4223,In_1890);
or U96 (N_96,In_3013,In_471);
xor U97 (N_97,In_515,In_4634);
and U98 (N_98,In_4426,In_4240);
and U99 (N_99,In_2281,In_1183);
and U100 (N_100,In_4418,In_1998);
nor U101 (N_101,In_234,In_4204);
nor U102 (N_102,In_2649,In_2098);
nor U103 (N_103,In_4157,In_1039);
nor U104 (N_104,In_2132,In_4894);
and U105 (N_105,In_2718,In_4884);
nor U106 (N_106,In_118,In_2508);
nor U107 (N_107,In_1881,In_440);
xor U108 (N_108,In_750,In_1680);
nand U109 (N_109,In_3547,In_3494);
or U110 (N_110,In_699,In_4487);
and U111 (N_111,In_900,In_1671);
and U112 (N_112,In_2034,In_749);
nor U113 (N_113,In_4056,In_4103);
and U114 (N_114,In_82,In_3361);
or U115 (N_115,In_4999,In_4210);
xnor U116 (N_116,In_4928,In_897);
and U117 (N_117,In_2024,In_2186);
and U118 (N_118,In_1236,In_2834);
and U119 (N_119,In_2826,In_788);
or U120 (N_120,In_388,In_3803);
and U121 (N_121,In_4669,In_1936);
and U122 (N_122,In_2485,In_4022);
nor U123 (N_123,In_3150,In_3695);
nand U124 (N_124,In_4169,In_1260);
and U125 (N_125,In_455,In_1858);
or U126 (N_126,In_963,In_4447);
or U127 (N_127,In_3349,In_1736);
and U128 (N_128,In_78,In_62);
and U129 (N_129,In_4543,In_510);
nor U130 (N_130,In_3192,In_4588);
nand U131 (N_131,In_1928,In_613);
nor U132 (N_132,In_1525,In_1412);
nor U133 (N_133,In_457,In_4308);
xor U134 (N_134,In_3323,In_1620);
or U135 (N_135,In_4481,In_4398);
or U136 (N_136,In_4222,In_3937);
nand U137 (N_137,In_3972,In_4396);
xor U138 (N_138,In_3989,In_2179);
xor U139 (N_139,In_4388,In_849);
and U140 (N_140,In_3186,In_3892);
or U141 (N_141,In_4325,In_1237);
or U142 (N_142,In_1612,In_4386);
xnor U143 (N_143,In_1018,In_1933);
xor U144 (N_144,In_4996,In_1902);
or U145 (N_145,In_3123,In_4997);
xnor U146 (N_146,In_4174,In_971);
or U147 (N_147,In_2329,In_2990);
nor U148 (N_148,In_145,In_1797);
nand U149 (N_149,In_4734,In_1923);
xor U150 (N_150,In_3402,In_3451);
nor U151 (N_151,In_2982,In_3334);
nand U152 (N_152,In_4505,In_2591);
and U153 (N_153,In_4439,In_1617);
nand U154 (N_154,In_4028,In_2349);
and U155 (N_155,In_3968,In_1603);
and U156 (N_156,In_4642,In_4098);
and U157 (N_157,In_472,In_987);
and U158 (N_158,In_1251,In_3300);
nand U159 (N_159,In_924,In_523);
nor U160 (N_160,In_1668,In_3239);
xnor U161 (N_161,In_4284,In_2327);
and U162 (N_162,In_4102,In_2249);
xor U163 (N_163,In_2390,In_3827);
nor U164 (N_164,In_1110,In_2127);
nand U165 (N_165,In_4566,In_4175);
nand U166 (N_166,In_4182,In_831);
or U167 (N_167,In_2399,In_1546);
nor U168 (N_168,In_4121,In_1409);
xnor U169 (N_169,In_1032,In_1975);
xnor U170 (N_170,In_2372,In_3454);
xnor U171 (N_171,In_2612,In_4957);
and U172 (N_172,In_3995,In_3401);
xnor U173 (N_173,In_4313,In_3241);
nand U174 (N_174,In_842,In_4808);
nand U175 (N_175,In_4931,In_2665);
nor U176 (N_176,In_2487,In_1618);
nand U177 (N_177,In_3738,In_387);
and U178 (N_178,In_990,In_2570);
and U179 (N_179,In_2013,In_2924);
xnor U180 (N_180,In_939,In_222);
xnor U181 (N_181,In_1322,In_3657);
nand U182 (N_182,In_4112,In_3601);
nand U183 (N_183,In_531,In_4078);
nand U184 (N_184,In_544,In_2846);
nor U185 (N_185,In_4639,In_3286);
or U186 (N_186,In_863,In_1937);
or U187 (N_187,In_2636,In_3799);
nand U188 (N_188,In_2375,In_4785);
xor U189 (N_189,In_2685,In_3004);
or U190 (N_190,In_4369,In_4013);
or U191 (N_191,In_1165,In_1467);
xnor U192 (N_192,In_4138,In_4293);
or U193 (N_193,In_4758,In_2227);
nand U194 (N_194,In_1255,In_4883);
nand U195 (N_195,In_3206,In_1296);
or U196 (N_196,In_3309,In_843);
nand U197 (N_197,In_4827,In_311);
nor U198 (N_198,In_2960,In_1700);
nor U199 (N_199,In_1299,In_3088);
and U200 (N_200,In_3419,In_4820);
nor U201 (N_201,In_3947,In_4647);
or U202 (N_202,In_4541,In_3588);
xor U203 (N_203,In_1396,In_4423);
nor U204 (N_204,In_3749,In_2096);
xnor U205 (N_205,In_3292,In_2751);
nand U206 (N_206,In_2483,In_1275);
nand U207 (N_207,In_467,In_1946);
nor U208 (N_208,In_3754,In_3354);
nand U209 (N_209,In_413,In_3729);
or U210 (N_210,In_1784,In_2418);
xnor U211 (N_211,In_485,In_1175);
or U212 (N_212,In_4362,In_181);
nor U213 (N_213,In_4847,In_4564);
nand U214 (N_214,In_4237,In_3669);
nand U215 (N_215,In_4641,In_404);
and U216 (N_216,In_1905,In_4077);
nor U217 (N_217,In_1726,In_4462);
or U218 (N_218,In_3903,In_173);
or U219 (N_219,In_3545,In_1447);
or U220 (N_220,In_47,In_3204);
xnor U221 (N_221,In_3227,In_4401);
nand U222 (N_222,In_2285,In_2660);
nor U223 (N_223,In_220,In_3479);
or U224 (N_224,In_1074,In_1474);
and U225 (N_225,In_3128,In_137);
xnor U226 (N_226,In_2407,In_2242);
or U227 (N_227,In_2717,In_435);
and U228 (N_228,In_3544,In_3327);
nor U229 (N_229,In_3717,In_4353);
xnor U230 (N_230,In_1182,In_3442);
nand U231 (N_231,In_1143,In_4959);
nor U232 (N_232,In_3920,In_3929);
nor U233 (N_233,In_4699,In_1350);
and U234 (N_234,In_2906,In_4580);
nand U235 (N_235,In_3278,In_4788);
or U236 (N_236,In_185,In_1750);
nand U237 (N_237,In_106,In_896);
nand U238 (N_238,In_4685,In_726);
and U239 (N_239,In_911,In_2775);
or U240 (N_240,In_1127,In_2835);
or U241 (N_241,In_1712,In_2682);
and U242 (N_242,In_4472,In_2214);
nand U243 (N_243,In_1465,In_3752);
nor U244 (N_244,In_4648,In_2011);
nand U245 (N_245,In_1830,In_1118);
nand U246 (N_246,In_281,In_598);
xnor U247 (N_247,In_4630,In_2149);
xor U248 (N_248,In_1939,In_4535);
xor U249 (N_249,In_2202,In_4277);
nand U250 (N_250,In_4004,In_966);
nor U251 (N_251,In_1558,In_1103);
xor U252 (N_252,In_1195,In_3166);
nand U253 (N_253,In_286,In_2620);
nor U254 (N_254,In_469,In_1723);
xor U255 (N_255,In_258,In_1425);
and U256 (N_256,In_3289,In_498);
xnor U257 (N_257,In_1242,In_2415);
nand U258 (N_258,In_864,In_519);
nor U259 (N_259,In_4866,In_4303);
and U260 (N_260,In_985,In_213);
xnor U261 (N_261,In_1504,In_2472);
xor U262 (N_262,In_2056,In_4802);
or U263 (N_263,In_2025,In_4760);
nand U264 (N_264,In_46,In_1354);
and U265 (N_265,In_4149,In_3474);
nand U266 (N_266,In_756,In_3688);
or U267 (N_267,In_1130,In_1590);
xnor U268 (N_268,In_2610,In_1196);
or U269 (N_269,In_856,In_2171);
nor U270 (N_270,In_3865,In_1059);
or U271 (N_271,In_2684,In_3054);
nor U272 (N_272,In_3945,In_2266);
nor U273 (N_273,In_3528,In_2563);
or U274 (N_274,In_650,In_1641);
and U275 (N_275,In_4250,In_182);
nor U276 (N_276,In_3009,In_692);
and U277 (N_277,In_1573,In_2896);
nand U278 (N_278,In_3115,In_4804);
nor U279 (N_279,In_3043,In_0);
and U280 (N_280,In_1943,In_2696);
xnor U281 (N_281,In_1486,In_3584);
nand U282 (N_282,In_1966,In_2495);
nand U283 (N_283,In_2655,In_436);
nor U284 (N_284,In_304,In_1692);
xnor U285 (N_285,In_3180,In_3161);
xnor U286 (N_286,In_1194,In_3246);
or U287 (N_287,In_1310,In_54);
or U288 (N_288,In_3619,In_301);
nand U289 (N_289,In_3846,In_3218);
xor U290 (N_290,In_550,In_2290);
or U291 (N_291,In_3693,In_3498);
nand U292 (N_292,In_1748,In_979);
nor U293 (N_293,In_2355,In_2791);
nor U294 (N_294,In_4898,In_3486);
and U295 (N_295,In_1536,In_1252);
xnor U296 (N_296,In_4469,In_652);
nand U297 (N_297,In_1506,In_4867);
nand U298 (N_298,In_1731,In_3935);
and U299 (N_299,In_1704,In_2254);
and U300 (N_300,In_4814,In_3538);
nor U301 (N_301,In_3913,In_4490);
xor U302 (N_302,In_2027,In_3067);
and U303 (N_303,In_4166,In_3103);
nor U304 (N_304,In_4909,In_3720);
nand U305 (N_305,In_4524,In_4864);
nand U306 (N_306,In_2299,In_420);
xnor U307 (N_307,In_1058,In_1204);
nor U308 (N_308,In_3750,In_3443);
and U309 (N_309,In_2189,In_4990);
and U310 (N_310,In_3036,In_2746);
xor U311 (N_311,In_4938,In_4702);
nor U312 (N_312,In_562,In_585);
and U313 (N_313,In_159,In_4671);
or U314 (N_314,In_4826,In_3093);
nor U315 (N_315,In_4415,In_4739);
or U316 (N_316,In_4600,In_2287);
nor U317 (N_317,In_590,In_3760);
nor U318 (N_318,In_1046,In_156);
or U319 (N_319,In_561,In_4697);
and U320 (N_320,In_1336,In_3119);
xor U321 (N_321,In_4766,In_1375);
nor U322 (N_322,In_803,In_3121);
or U323 (N_323,In_1882,In_1656);
and U324 (N_324,In_103,In_3453);
nand U325 (N_325,In_2233,In_4368);
and U326 (N_326,In_4305,In_4993);
xor U327 (N_327,In_556,In_4672);
or U328 (N_328,In_2311,In_4217);
xor U329 (N_329,In_3397,In_4845);
nand U330 (N_330,In_2873,In_2449);
xor U331 (N_331,In_4893,In_818);
xnor U332 (N_332,In_4212,In_2919);
xor U333 (N_333,In_623,In_1141);
nand U334 (N_334,In_3175,In_4779);
nor U335 (N_335,In_3050,In_2510);
xnor U336 (N_336,In_1220,In_2267);
and U337 (N_337,In_769,In_2050);
nand U338 (N_338,In_4746,In_3065);
nand U339 (N_339,In_1448,In_1807);
and U340 (N_340,In_3434,In_2093);
xor U341 (N_341,In_4335,In_41);
nand U342 (N_342,In_190,In_2855);
and U343 (N_343,In_2221,In_4608);
nand U344 (N_344,In_2276,In_2062);
or U345 (N_345,In_4970,In_2288);
nand U346 (N_346,In_1529,In_1364);
or U347 (N_347,In_4191,In_1725);
xor U348 (N_348,In_567,In_4376);
or U349 (N_349,In_1167,In_317);
or U350 (N_350,In_2165,In_1497);
nand U351 (N_351,In_4253,In_4629);
nor U352 (N_352,In_3656,In_1264);
nor U353 (N_353,In_3312,In_2392);
nand U354 (N_354,In_1424,In_895);
xnor U355 (N_355,In_2515,In_4531);
xnor U356 (N_356,In_4687,In_3084);
xor U357 (N_357,In_931,In_4711);
or U358 (N_358,In_4323,In_745);
xor U359 (N_359,In_3651,In_3141);
nand U360 (N_360,In_2169,In_2535);
and U361 (N_361,In_2184,In_44);
and U362 (N_362,In_3345,In_3041);
xor U363 (N_363,In_3718,In_1650);
and U364 (N_364,In_4862,In_153);
nand U365 (N_365,In_432,In_327);
xor U366 (N_366,In_3655,In_1791);
nand U367 (N_367,In_4787,In_2815);
xnor U368 (N_368,In_3376,In_3645);
xnor U369 (N_369,In_2984,In_1604);
and U370 (N_370,In_2082,In_4085);
and U371 (N_371,In_4290,In_3553);
xor U372 (N_372,In_1665,In_1114);
and U373 (N_373,In_3866,In_3492);
nand U374 (N_374,In_3953,In_3371);
nor U375 (N_375,In_4186,In_504);
or U376 (N_376,In_1824,In_3868);
nor U377 (N_377,In_1147,In_1135);
xor U378 (N_378,In_1487,In_1913);
or U379 (N_379,In_2353,In_1980);
nand U380 (N_380,In_4266,In_835);
xnor U381 (N_381,In_1286,In_1948);
nor U382 (N_382,In_1117,In_4603);
or U383 (N_383,In_2832,In_3412);
nor U384 (N_384,In_3364,In_1308);
and U385 (N_385,In_976,In_3691);
nand U386 (N_386,In_2615,In_1470);
or U387 (N_387,In_4715,In_3839);
nor U388 (N_388,In_2282,In_4885);
nand U389 (N_389,In_2770,In_322);
nand U390 (N_390,In_337,In_4638);
nor U391 (N_391,In_4320,In_99);
nand U392 (N_392,In_113,In_272);
nor U393 (N_393,In_4128,In_2010);
or U394 (N_394,In_4450,In_2293);
nand U395 (N_395,In_2614,In_3415);
or U396 (N_396,In_983,In_3398);
nor U397 (N_397,In_3185,In_589);
and U398 (N_398,In_1274,In_1329);
nor U399 (N_399,In_651,In_2092);
and U400 (N_400,In_1372,In_3711);
or U401 (N_401,In_1433,In_1050);
or U402 (N_402,In_3576,In_1380);
or U403 (N_403,In_4624,In_3181);
and U404 (N_404,In_263,In_3973);
or U405 (N_405,In_2198,In_339);
and U406 (N_406,In_189,In_3163);
and U407 (N_407,In_4007,In_3460);
nand U408 (N_408,In_3350,In_3684);
nor U409 (N_409,In_2863,In_3014);
nor U410 (N_410,In_3894,In_86);
xor U411 (N_411,In_50,In_1810);
xnor U412 (N_412,In_2362,In_277);
or U413 (N_413,In_1269,In_3254);
nand U414 (N_414,In_830,In_4326);
xnor U415 (N_415,In_4264,In_2576);
and U416 (N_416,In_2695,In_1044);
nand U417 (N_417,In_1982,In_3238);
nand U418 (N_418,In_582,In_2860);
and U419 (N_419,In_1104,In_4177);
xor U420 (N_420,In_95,In_2364);
nor U421 (N_421,In_2196,In_4553);
xnor U422 (N_422,In_4843,In_2152);
and U423 (N_423,In_595,In_3082);
nand U424 (N_424,In_1592,In_3410);
nor U425 (N_425,In_3692,In_1508);
and U426 (N_426,In_4683,In_4385);
nand U427 (N_427,In_101,In_1631);
nor U428 (N_428,In_2818,In_3074);
or U429 (N_429,In_630,In_3168);
and U430 (N_430,In_4962,In_960);
nand U431 (N_431,In_111,In_3801);
nand U432 (N_432,In_3617,In_3616);
nand U433 (N_433,In_450,In_4700);
and U434 (N_434,In_4981,In_3374);
or U435 (N_435,In_1266,In_2514);
xor U436 (N_436,In_3887,In_4486);
nor U437 (N_437,In_1722,In_599);
nand U438 (N_438,In_61,In_60);
xnor U439 (N_439,In_334,In_3560);
nor U440 (N_440,In_1026,In_2819);
and U441 (N_441,In_1883,In_2484);
and U442 (N_442,In_298,In_53);
nor U443 (N_443,In_3363,In_410);
xnor U444 (N_444,In_1972,In_2580);
and U445 (N_445,In_4127,In_1895);
and U446 (N_446,In_4404,In_2031);
xor U447 (N_447,In_3336,In_2895);
and U448 (N_448,In_3814,In_4458);
and U449 (N_449,In_3796,In_3506);
nor U450 (N_450,In_1809,In_1666);
and U451 (N_451,In_3638,In_1483);
xnor U452 (N_452,In_3317,In_3137);
and U453 (N_453,In_2710,In_840);
or U454 (N_454,In_2956,In_1476);
and U455 (N_455,In_2912,In_4465);
xor U456 (N_456,In_4020,In_1009);
and U457 (N_457,In_2437,In_1755);
nand U458 (N_458,In_4784,In_1277);
or U459 (N_459,In_2579,In_1615);
or U460 (N_460,In_3941,In_1871);
or U461 (N_461,In_4592,In_3793);
nand U462 (N_462,In_3042,In_4689);
nand U463 (N_463,In_1563,In_1745);
xor U464 (N_464,In_3273,In_760);
nor U465 (N_465,In_3220,In_867);
nand U466 (N_466,In_4343,In_3176);
and U467 (N_467,In_2590,In_3936);
nand U468 (N_468,In_4065,In_1762);
or U469 (N_469,In_2882,In_2128);
or U470 (N_470,In_4132,In_682);
nand U471 (N_471,In_3196,In_1889);
nor U472 (N_472,In_2848,In_4170);
nand U473 (N_473,In_3129,In_2173);
nand U474 (N_474,In_4471,In_815);
or U475 (N_475,In_3636,In_4615);
and U476 (N_476,In_3643,In_489);
xnor U477 (N_477,In_4951,In_2121);
xnor U478 (N_478,In_2441,In_3097);
nand U479 (N_479,In_2934,In_3904);
nor U480 (N_480,In_935,In_3907);
xnor U481 (N_481,In_973,In_3783);
xor U482 (N_482,In_4095,In_4747);
or U483 (N_483,In_4610,In_419);
nand U484 (N_484,In_4932,In_3607);
and U485 (N_485,In_4913,In_1095);
and U486 (N_486,In_3831,In_316);
nor U487 (N_487,In_730,In_355);
or U488 (N_488,In_4618,In_4660);
and U489 (N_489,In_1545,In_2539);
or U490 (N_490,In_3112,In_3390);
nor U491 (N_491,In_2491,In_1786);
nor U492 (N_492,In_933,In_4100);
nor U493 (N_493,In_33,In_1644);
nor U494 (N_494,In_1100,In_1938);
nand U495 (N_495,In_2361,In_2516);
nor U496 (N_496,In_3439,In_3932);
xor U497 (N_497,In_4443,In_3027);
and U498 (N_498,In_3499,In_563);
or U499 (N_499,In_1414,In_1023);
nor U500 (N_500,In_4206,In_4530);
xor U501 (N_501,In_3403,In_537);
or U502 (N_502,In_2572,In_4344);
nand U503 (N_503,In_754,In_1327);
or U504 (N_504,In_4891,In_3063);
nor U505 (N_505,In_18,In_1553);
xnor U506 (N_506,In_3757,In_1862);
xnor U507 (N_507,In_2878,In_4791);
or U508 (N_508,In_2145,In_1222);
nand U509 (N_509,In_3427,In_952);
or U510 (N_510,In_3979,In_2509);
nand U511 (N_511,In_3413,In_3420);
or U512 (N_512,In_52,In_170);
and U513 (N_513,In_2393,In_409);
nor U514 (N_514,In_4165,In_346);
nor U515 (N_515,In_3435,In_171);
xor U516 (N_516,In_488,In_4051);
or U517 (N_517,In_486,In_4094);
xnor U518 (N_518,In_2429,In_4086);
or U519 (N_519,In_3158,In_1028);
xor U520 (N_520,In_4545,In_1609);
nor U521 (N_521,In_2651,In_3099);
and U522 (N_522,In_2807,In_2507);
and U523 (N_523,In_3114,In_1079);
or U524 (N_524,In_4332,In_1540);
or U525 (N_525,In_1090,In_883);
and U526 (N_526,In_1036,In_2460);
xnor U527 (N_527,In_1199,In_292);
xnor U528 (N_528,In_5,In_662);
nand U529 (N_529,In_2688,In_3602);
nand U530 (N_530,In_2229,In_3262);
or U531 (N_531,In_4786,In_1677);
nor U532 (N_532,In_642,In_781);
xor U533 (N_533,In_1727,In_4617);
nand U534 (N_534,In_4707,In_2271);
and U535 (N_535,In_3458,In_1811);
xnor U536 (N_536,In_177,In_1385);
xor U537 (N_537,In_3608,In_2613);
xnor U538 (N_538,In_611,In_261);
and U539 (N_539,In_1770,In_26);
nor U540 (N_540,In_1353,In_3694);
xnor U541 (N_541,In_1706,In_3117);
nand U542 (N_542,In_3627,In_3038);
nand U543 (N_543,In_2448,In_1158);
and U544 (N_544,In_3301,In_1156);
nand U545 (N_545,In_2320,In_2792);
nor U546 (N_546,In_3131,In_3030);
nor U547 (N_547,In_3049,In_4805);
or U548 (N_548,In_1343,In_116);
xnor U549 (N_549,In_3551,In_491);
nand U550 (N_550,In_641,In_3817);
xnor U551 (N_551,In_1060,In_3537);
nor U552 (N_552,In_4038,In_1326);
nor U553 (N_553,In_407,In_2892);
or U554 (N_554,In_4679,In_1960);
nor U555 (N_555,In_1211,In_4675);
nor U556 (N_556,In_290,In_1002);
nor U557 (N_557,In_74,In_114);
xor U558 (N_558,In_2286,In_1645);
or U559 (N_559,In_955,In_218);
nor U560 (N_560,In_3265,In_4842);
or U561 (N_561,In_4035,In_1218);
nor U562 (N_562,In_4176,In_1265);
or U563 (N_563,In_2482,In_3559);
and U564 (N_564,In_2757,In_947);
and U565 (N_565,In_1900,In_1829);
and U566 (N_566,In_4442,In_1587);
or U567 (N_567,In_1585,In_1756);
nand U568 (N_568,In_3348,In_367);
nor U569 (N_569,In_1405,In_2829);
nor U570 (N_570,In_1309,In_2403);
nor U571 (N_571,In_2943,In_1843);
nor U572 (N_572,In_3224,In_3216);
xor U573 (N_573,In_3039,In_1284);
and U574 (N_574,In_4706,In_4273);
and U575 (N_575,In_476,In_850);
or U576 (N_576,In_4853,In_133);
xnor U577 (N_577,In_2391,In_4552);
and U578 (N_578,In_1468,In_3126);
xor U579 (N_579,In_4214,In_2814);
and U580 (N_580,In_4161,In_2017);
and U581 (N_581,In_1225,In_758);
nand U582 (N_582,In_4520,In_2120);
and U583 (N_583,In_2084,In_3587);
or U584 (N_584,In_660,In_2822);
xor U585 (N_585,In_3683,In_1834);
nor U586 (N_586,In_812,In_2886);
xor U587 (N_587,In_1458,In_4992);
or U588 (N_588,In_2357,In_215);
and U589 (N_589,In_4888,In_1842);
and U590 (N_590,In_780,In_3096);
xnor U591 (N_591,In_1422,In_1294);
nand U592 (N_592,In_1351,In_2578);
and U593 (N_593,In_1763,In_3319);
and U594 (N_594,In_4934,In_2527);
and U595 (N_595,In_1214,In_2040);
or U596 (N_596,In_739,In_1962);
nand U597 (N_597,In_3795,In_1232);
nor U598 (N_598,In_1865,In_2643);
and U599 (N_599,In_4667,In_2987);
xor U600 (N_600,In_4045,In_237);
nand U601 (N_601,In_3476,In_1170);
or U602 (N_602,In_2537,In_4159);
nand U603 (N_603,In_1144,In_2467);
nor U604 (N_604,In_3772,In_1187);
nand U605 (N_605,In_212,In_2065);
nor U606 (N_606,In_312,In_2630);
nor U607 (N_607,In_65,In_839);
nand U608 (N_608,In_374,In_1369);
xor U609 (N_609,In_1096,In_1991);
nor U610 (N_610,In_2347,In_172);
or U611 (N_611,In_459,In_4097);
or U612 (N_612,In_2532,In_4060);
nand U613 (N_613,In_776,In_748);
nand U614 (N_614,In_3400,In_4529);
or U615 (N_615,In_194,In_2030);
xor U616 (N_616,In_1718,In_1820);
and U617 (N_617,In_1502,In_2884);
nand U618 (N_618,In_3558,In_4267);
or U619 (N_619,In_624,In_2162);
xor U620 (N_620,In_1557,In_4595);
or U621 (N_621,In_4728,In_1593);
xor U622 (N_622,In_688,In_1581);
and U623 (N_623,In_1460,In_639);
xor U624 (N_624,In_3784,In_3709);
and U625 (N_625,In_3733,In_1316);
or U626 (N_626,In_3465,In_536);
nand U627 (N_627,In_4574,In_2675);
nand U628 (N_628,In_4088,In_1776);
xor U629 (N_629,In_330,In_3395);
or U630 (N_630,In_727,In_1800);
and U631 (N_631,In_2644,In_4859);
nor U632 (N_632,In_2801,In_3127);
and U633 (N_633,In_3880,In_4765);
xnor U634 (N_634,In_4936,In_379);
nor U635 (N_635,In_1073,In_425);
and U636 (N_636,In_2966,In_3781);
or U637 (N_637,In_3102,In_3574);
and U638 (N_638,In_1087,In_4732);
nor U639 (N_639,In_4631,In_3108);
and U640 (N_640,In_2176,In_2261);
nand U641 (N_641,In_2813,In_1908);
and U642 (N_642,In_2377,In_2319);
xor U643 (N_643,In_689,In_3940);
or U644 (N_644,In_4265,In_1851);
nor U645 (N_645,In_923,In_3264);
nand U646 (N_646,In_1081,In_3324);
nor U647 (N_647,In_2726,In_4964);
nand U648 (N_648,In_3406,In_2172);
or U649 (N_649,In_3017,In_2739);
nor U650 (N_650,In_276,In_4619);
nand U651 (N_651,In_3522,In_588);
and U652 (N_652,In_3514,In_275);
xor U653 (N_653,In_1221,In_1478);
nor U654 (N_654,In_2724,In_323);
or U655 (N_655,In_4047,In_2861);
nor U656 (N_656,In_4577,In_742);
nor U657 (N_657,In_4963,In_3426);
nor U658 (N_658,In_2503,In_2870);
and U659 (N_659,In_3533,In_1201);
xor U660 (N_660,In_1891,In_2425);
and U661 (N_661,In_1703,In_4646);
and U662 (N_662,In_314,In_4757);
nor U663 (N_663,In_2812,In_2430);
xnor U664 (N_664,In_4205,In_591);
and U665 (N_665,In_3769,In_865);
nand U666 (N_666,In_1112,In_2422);
and U667 (N_667,In_1123,In_810);
or U668 (N_668,In_331,In_2883);
and U669 (N_669,In_792,In_3748);
and U670 (N_670,In_1282,In_4330);
xor U671 (N_671,In_1339,In_3230);
xnor U672 (N_672,In_2948,In_3531);
nand U673 (N_673,In_1628,In_2754);
nor U674 (N_674,In_1004,In_3835);
or U675 (N_675,In_1888,In_2842);
and U676 (N_676,In_3001,In_2663);
or U677 (N_677,In_974,In_1805);
or U678 (N_678,In_1918,In_1200);
xnor U679 (N_679,In_4737,In_846);
xnor U680 (N_680,In_3853,In_1798);
nor U681 (N_681,In_3614,In_3193);
xor U682 (N_682,In_2394,In_2917);
nand U683 (N_683,In_3942,In_723);
and U684 (N_684,In_3854,In_1694);
nor U685 (N_685,In_1055,In_1693);
nor U686 (N_686,In_3347,In_12);
and U687 (N_687,In_870,In_1556);
or U688 (N_688,In_1042,In_3734);
or U689 (N_689,In_3950,In_1052);
nand U690 (N_690,In_1289,In_1780);
nand U691 (N_691,In_3513,In_3025);
nor U692 (N_692,In_4281,In_1495);
or U693 (N_693,In_661,In_3837);
xor U694 (N_694,In_1815,In_2069);
or U695 (N_695,In_1241,In_4953);
nand U696 (N_696,In_259,In_340);
nor U697 (N_697,In_4824,In_4812);
nor U698 (N_698,In_1571,In_681);
nor U699 (N_699,In_4391,In_2256);
or U700 (N_700,In_4998,In_3763);
xor U701 (N_701,In_3613,In_2102);
xnor U702 (N_702,In_3773,In_4470);
xor U703 (N_703,In_1446,In_325);
nor U704 (N_704,In_4037,In_11);
nand U705 (N_705,In_2302,In_609);
xor U706 (N_706,In_673,In_3199);
nor U707 (N_707,In_4873,In_112);
nand U708 (N_708,In_3411,In_1614);
and U709 (N_709,In_3741,In_3228);
xnor U710 (N_710,In_4082,In_2297);
xor U711 (N_711,In_453,In_762);
nand U712 (N_712,In_4972,In_108);
and U713 (N_713,In_2387,In_3340);
nor U714 (N_714,In_4338,In_3375);
nor U715 (N_715,In_4488,In_2365);
or U716 (N_716,In_2993,In_2053);
xor U717 (N_717,In_2512,In_553);
or U718 (N_718,In_4195,In_431);
nand U719 (N_719,In_2036,In_1007);
nor U720 (N_720,In_3316,In_1528);
xor U721 (N_721,In_1802,In_1270);
and U722 (N_722,In_3804,In_4032);
nor U723 (N_723,In_1490,In_3202);
nand U724 (N_724,In_1793,In_2218);
and U725 (N_725,In_1010,In_2223);
nor U726 (N_726,In_4651,In_1159);
and U727 (N_727,In_1000,In_2006);
and U728 (N_728,In_852,In_4514);
xnor U729 (N_729,In_3834,In_4023);
nor U730 (N_730,In_207,In_4887);
nor U731 (N_731,In_2602,In_72);
nand U732 (N_732,In_1526,In_4753);
or U733 (N_733,In_2779,In_1552);
xor U734 (N_734,In_4512,In_3060);
xor U735 (N_735,In_2188,In_2977);
or U736 (N_736,In_2853,In_1926);
nor U737 (N_737,In_3353,In_4430);
or U738 (N_738,In_3652,In_3500);
or U739 (N_739,In_358,In_4995);
nor U740 (N_740,In_901,In_3970);
nor U741 (N_741,In_4314,In_4923);
nor U742 (N_742,In_4324,In_2331);
and U743 (N_743,In_2788,In_2523);
nor U744 (N_744,In_2183,In_2647);
and U745 (N_745,In_1624,In_205);
and U746 (N_746,In_4852,In_3768);
nand U747 (N_747,In_251,In_3610);
or U748 (N_748,In_2940,In_2831);
xor U749 (N_749,In_226,In_1751);
xor U750 (N_750,In_3618,In_3532);
and U751 (N_751,In_1273,In_3271);
or U752 (N_752,In_2657,In_1293);
xnor U753 (N_753,In_4790,In_2891);
xor U754 (N_754,In_368,In_581);
nor U755 (N_755,In_4361,In_3824);
and U756 (N_756,In_1136,In_2504);
and U757 (N_757,In_1463,In_1783);
nor U758 (N_758,In_695,In_1574);
xor U759 (N_759,In_3852,In_4201);
xor U760 (N_760,In_1670,In_3244);
and U761 (N_761,In_1288,In_2463);
nand U762 (N_762,In_1125,In_4494);
nand U763 (N_763,In_2235,In_2244);
nor U764 (N_764,In_1057,In_3982);
xor U765 (N_765,In_3780,In_71);
and U766 (N_766,In_1632,In_2797);
and U767 (N_767,In_2099,In_4969);
or U768 (N_768,In_2417,In_428);
nor U769 (N_769,In_2787,In_2709);
and U770 (N_770,In_4039,In_288);
xnor U771 (N_771,In_3235,In_1947);
nand U772 (N_772,In_535,In_3833);
nor U773 (N_773,In_3591,In_4724);
nand U774 (N_774,In_3006,In_4328);
or U775 (N_775,In_267,In_2061);
and U776 (N_776,In_3106,In_721);
nand U777 (N_777,In_2631,In_3697);
or U778 (N_778,In_821,In_4063);
nor U779 (N_779,In_3022,In_3702);
and U780 (N_780,In_4257,In_2719);
and U781 (N_781,In_2257,In_2925);
and U782 (N_782,In_3843,In_708);
xor U783 (N_783,In_2279,In_3061);
xor U784 (N_784,In_1942,In_4111);
nand U785 (N_785,In_4775,In_2493);
xor U786 (N_786,In_3139,In_2558);
xnor U787 (N_787,In_2314,In_1916);
nand U788 (N_788,In_3659,In_816);
nand U789 (N_789,In_1782,In_1555);
xor U790 (N_790,In_4151,In_88);
nand U791 (N_791,In_3646,In_3125);
nor U792 (N_792,In_1658,In_4919);
or U793 (N_793,In_4233,In_3787);
xor U794 (N_794,In_671,In_3182);
and U795 (N_795,In_572,In_4276);
nor U796 (N_796,In_2343,In_1663);
nor U797 (N_797,In_1034,In_2154);
or U798 (N_798,In_1013,In_3661);
xor U799 (N_799,In_4517,In_4006);
nand U800 (N_800,In_2851,In_2313);
nand U801 (N_801,In_919,In_320);
xor U802 (N_802,In_2571,In_4080);
xor U803 (N_803,In_2683,In_1822);
nor U804 (N_804,In_1072,In_2346);
xnor U805 (N_805,In_3142,In_2112);
or U806 (N_806,In_1635,In_2318);
nor U807 (N_807,In_3064,In_1539);
or U808 (N_808,In_4816,In_120);
or U809 (N_809,In_3705,In_2859);
and U810 (N_810,In_1333,In_2996);
xnor U811 (N_811,In_2686,In_3840);
and U812 (N_812,In_1056,In_3707);
nand U813 (N_813,In_3069,In_4484);
and U814 (N_814,In_694,In_3890);
nand U815 (N_815,In_2246,In_4409);
nor U816 (N_816,In_2811,In_918);
xor U817 (N_817,In_2627,In_2652);
nor U818 (N_818,In_227,In_1038);
and U819 (N_819,In_447,In_722);
nand U820 (N_820,In_4515,In_3621);
nor U821 (N_821,In_3943,In_736);
or U822 (N_822,In_1864,In_161);
and U823 (N_823,In_577,In_1338);
or U824 (N_824,In_514,In_3938);
nor U825 (N_825,In_1105,In_3654);
nor U826 (N_826,In_2486,In_1124);
nand U827 (N_827,In_2070,In_1852);
xor U828 (N_828,In_4584,In_2601);
nor U829 (N_829,In_4383,In_4501);
nand U830 (N_830,In_1575,In_2517);
xnor U831 (N_831,In_315,In_4050);
nor U832 (N_832,In_2048,In_2150);
nor U833 (N_833,In_2187,In_2103);
and U834 (N_834,In_752,In_495);
nor U835 (N_835,In_4117,In_2380);
or U836 (N_836,In_293,In_4583);
or U837 (N_837,In_487,In_4115);
and U838 (N_838,In_204,In_1092);
and U839 (N_839,In_3495,In_4763);
xor U840 (N_840,In_2324,In_797);
and U841 (N_841,In_4872,In_1250);
xnor U842 (N_842,In_825,In_909);
nand U843 (N_843,In_2194,In_2789);
and U844 (N_844,In_1192,In_4730);
xor U845 (N_845,In_3679,In_3954);
nand U846 (N_846,In_3663,In_193);
or U847 (N_847,In_4559,In_3633);
and U848 (N_848,In_4832,In_155);
xor U849 (N_849,In_2905,In_3000);
nor U850 (N_850,In_1416,In_3882);
nand U851 (N_851,In_3207,In_1256);
and U852 (N_852,In_1992,In_285);
and U853 (N_853,In_667,In_3322);
xor U854 (N_854,In_1894,In_2747);
nor U855 (N_855,In_4058,In_956);
nand U856 (N_856,In_811,In_3315);
nand U857 (N_857,In_280,In_4774);
nand U858 (N_858,In_4662,In_2914);
xor U859 (N_859,In_3358,In_268);
and U860 (N_860,In_1956,In_2317);
xnor U861 (N_861,In_3511,In_4571);
nor U862 (N_862,In_2854,In_4819);
nor U863 (N_863,In_3255,In_3861);
nor U864 (N_864,In_4300,In_4725);
or U865 (N_865,In_151,In_2777);
xnor U866 (N_866,In_3387,In_475);
nor U867 (N_867,In_2178,In_2689);
and U868 (N_868,In_142,In_4122);
nor U869 (N_869,In_3534,In_2395);
xnor U870 (N_870,In_4349,In_4150);
nand U871 (N_871,In_437,In_4770);
nor U872 (N_872,In_2489,In_3356);
xor U873 (N_873,In_3475,In_1597);
nand U874 (N_874,In_1837,In_860);
and U875 (N_875,In_2911,In_2561);
or U876 (N_876,In_307,In_512);
nand U877 (N_877,In_2248,In_1713);
xor U878 (N_878,In_759,In_4989);
xnor U879 (N_879,In_1764,In_2063);
or U880 (N_880,In_2699,In_4341);
nor U881 (N_881,In_3603,In_4317);
nand U882 (N_882,In_4828,In_2354);
and U883 (N_883,In_3379,In_3876);
nor U884 (N_884,In_3874,In_4861);
nand U885 (N_885,In_3666,In_2305);
or U886 (N_886,In_1701,In_2367);
and U887 (N_887,In_3736,In_4040);
nand U888 (N_888,In_4777,In_4637);
or U889 (N_889,In_4947,In_4991);
nor U890 (N_890,In_1667,In_3310);
and U891 (N_891,In_4381,In_774);
and U892 (N_892,In_1391,In_832);
and U893 (N_893,In_3087,In_4500);
and U894 (N_894,In_4026,In_4858);
xor U895 (N_895,In_4231,In_1016);
xnor U896 (N_896,In_1833,In_1489);
nand U897 (N_897,In_3919,In_3554);
and U898 (N_898,In_805,In_4492);
nand U899 (N_899,In_1402,In_448);
nor U900 (N_900,In_1347,In_1739);
xor U901 (N_901,In_782,In_1757);
xor U902 (N_902,In_3990,In_2157);
xor U903 (N_903,In_3747,In_4654);
xor U904 (N_904,In_3821,In_4200);
or U905 (N_905,In_3615,In_1404);
and U906 (N_906,In_3120,In_2544);
nor U907 (N_907,In_1657,In_1025);
and U908 (N_908,In_508,In_2398);
nor U909 (N_909,In_4336,In_2479);
nand U910 (N_910,In_2833,In_614);
xnor U911 (N_911,In_1983,In_4994);
or U912 (N_912,In_2066,In_2584);
xor U913 (N_913,In_3889,In_632);
or U914 (N_914,In_3152,In_1921);
and U915 (N_915,In_702,In_2181);
nand U916 (N_916,In_3107,In_1532);
and U917 (N_917,In_4557,In_1166);
xnor U918 (N_918,In_2758,In_4684);
nand U919 (N_919,In_2945,In_1394);
or U920 (N_920,In_2946,In_3790);
and U921 (N_921,In_3066,In_4966);
and U922 (N_922,In_135,In_993);
nor U923 (N_923,In_2265,In_4573);
nor U924 (N_924,In_4694,In_2119);
nand U925 (N_925,In_3225,In_621);
nand U926 (N_926,In_2658,In_3884);
and U927 (N_927,In_4511,In_3675);
and U928 (N_928,In_4158,In_3252);
xnor U929 (N_929,In_705,In_4897);
or U930 (N_930,In_2536,In_625);
and U931 (N_931,In_4502,In_2961);
nand U932 (N_932,In_2078,In_1371);
or U933 (N_933,In_3483,In_644);
xnor U934 (N_934,In_372,In_2714);
and U935 (N_935,In_2784,In_4405);
or U936 (N_936,In_1787,In_1494);
or U937 (N_937,In_1331,In_3034);
and U938 (N_938,In_3548,In_2005);
and U939 (N_939,In_4682,In_418);
xor U940 (N_940,In_1435,In_1078);
nand U941 (N_941,In_3829,In_1053);
or U942 (N_942,In_2153,In_4536);
nand U943 (N_943,In_2622,In_3939);
xnor U944 (N_944,In_3058,In_817);
nand U945 (N_945,In_3759,In_594);
and U946 (N_946,In_3704,In_3449);
xnor U947 (N_947,In_916,In_1863);
or U948 (N_948,In_1219,In_4863);
nand U949 (N_949,In_786,In_4633);
nor U950 (N_950,In_3385,In_4918);
nand U951 (N_951,In_398,In_4145);
or U952 (N_952,In_4590,In_4147);
xnor U953 (N_953,In_4283,In_492);
and U954 (N_954,In_4350,In_132);
nor U955 (N_955,In_3994,In_3916);
and U956 (N_956,In_15,In_3622);
xor U957 (N_957,In_4907,In_4378);
nor U958 (N_958,In_1958,In_2796);
and U959 (N_959,In_2049,In_4202);
or U960 (N_960,In_2312,In_1378);
nor U961 (N_961,In_3715,In_1637);
nand U962 (N_962,In_996,In_4635);
xor U963 (N_963,In_1070,In_4681);
nor U964 (N_964,In_3523,In_2918);
nor U965 (N_965,In_1276,In_3563);
or U966 (N_966,In_3135,In_1089);
nor U967 (N_967,In_3237,In_497);
nor U968 (N_968,In_1238,In_1291);
or U969 (N_969,In_2850,In_1708);
nor U970 (N_970,In_345,In_2967);
nor U971 (N_971,In_1113,In_4834);
or U972 (N_972,In_712,In_1314);
or U973 (N_973,In_321,In_873);
nand U974 (N_974,In_4575,In_887);
or U975 (N_975,In_1462,In_3580);
nor U976 (N_976,In_3766,In_691);
nor U977 (N_977,In_1720,In_380);
xnor U978 (N_978,In_4688,In_2475);
xor U979 (N_979,In_4066,In_3052);
nor U980 (N_980,In_2095,In_3983);
nor U981 (N_981,In_2621,In_4025);
nor U982 (N_982,In_1233,In_3917);
nor U983 (N_983,In_1819,In_2245);
nand U984 (N_984,In_2146,In_3589);
or U985 (N_985,In_64,In_1625);
xnor U986 (N_986,In_2459,In_2416);
or U987 (N_987,In_266,In_4445);
nor U988 (N_988,In_1929,In_4431);
and U989 (N_989,In_3630,In_211);
nand U990 (N_990,In_580,In_4935);
or U991 (N_991,In_362,In_3540);
and U992 (N_992,In_4886,In_1774);
or U993 (N_993,In_1041,In_732);
nand U994 (N_994,In_1097,In_2502);
and U995 (N_995,In_365,In_2262);
nand U996 (N_996,In_2935,In_1313);
and U997 (N_997,In_824,In_479);
nand U998 (N_998,In_3845,In_1098);
nand U999 (N_999,In_1818,In_767);
nor U1000 (N_1000,In_4239,In_2765);
and U1001 (N_1001,In_4370,In_383);
and U1002 (N_1002,In_117,In_4759);
or U1003 (N_1003,In_2490,In_2869);
xnor U1004 (N_1004,In_4245,In_335);
or U1005 (N_1005,In_1381,In_3525);
xnor U1006 (N_1006,In_1181,In_3786);
and U1007 (N_1007,In_1964,In_2793);
or U1008 (N_1008,In_4310,In_807);
xor U1009 (N_1009,In_4001,In_2426);
or U1010 (N_1010,In_725,In_3764);
and U1011 (N_1011,In_4544,In_2748);
nand U1012 (N_1012,In_3138,In_175);
xor U1013 (N_1013,In_4255,In_2750);
or U1014 (N_1014,In_604,In_283);
nand U1015 (N_1015,In_2847,In_415);
nand U1016 (N_1016,In_2866,In_4705);
and U1017 (N_1017,In_2136,In_848);
nand U1018 (N_1018,In_746,In_3585);
nor U1019 (N_1019,In_3478,In_3077);
or U1020 (N_1020,In_1914,In_3996);
nor U1021 (N_1021,In_2088,In_2573);
or U1022 (N_1022,In_2574,In_370);
and U1023 (N_1023,In_2795,In_1990);
or U1024 (N_1024,In_1021,In_1976);
and U1025 (N_1025,In_4451,In_1001);
nor U1026 (N_1026,In_1661,In_396);
nor U1027 (N_1027,In_4048,In_4288);
and U1028 (N_1028,In_2081,In_2659);
xor U1029 (N_1029,In_1441,In_890);
or U1030 (N_1030,In_4093,In_4904);
nand U1031 (N_1031,In_3519,In_2462);
nand U1032 (N_1032,In_19,In_1564);
xor U1033 (N_1033,In_1930,In_2280);
or U1034 (N_1034,In_3981,In_4640);
and U1035 (N_1035,In_2258,In_1760);
xor U1036 (N_1036,In_470,In_3261);
or U1037 (N_1037,In_3198,In_2447);
xnor U1038 (N_1038,In_3595,In_3676);
nand U1039 (N_1039,In_2901,In_3081);
xor U1040 (N_1040,In_4692,In_2474);
nand U1041 (N_1041,In_2816,In_1685);
nand U1042 (N_1042,In_3648,In_1963);
nor U1043 (N_1043,In_804,In_4243);
and U1044 (N_1044,In_4655,In_4340);
and U1045 (N_1045,In_2874,In_3029);
and U1046 (N_1046,In_147,In_402);
nor U1047 (N_1047,In_3735,In_3712);
xnor U1048 (N_1048,In_2609,In_3912);
and U1049 (N_1049,In_4522,In_14);
and U1050 (N_1050,In_4537,In_1792);
nor U1051 (N_1051,In_2992,In_2129);
nand U1052 (N_1052,In_4153,In_3143);
and U1053 (N_1053,In_1534,In_875);
nor U1054 (N_1054,In_4542,In_1457);
nand U1055 (N_1055,In_2888,In_2206);
nor U1056 (N_1056,In_353,In_1169);
nor U1057 (N_1057,In_2825,In_1247);
nand U1058 (N_1058,In_2562,In_1610);
and U1059 (N_1059,In_494,In_4419);
nor U1060 (N_1060,In_466,In_1741);
nand U1061 (N_1061,In_795,In_4348);
and U1062 (N_1062,In_2306,In_4916);
nor U1063 (N_1063,In_4769,In_3886);
nor U1064 (N_1064,In_4279,In_2131);
or U1065 (N_1065,In_2728,In_97);
nand U1066 (N_1066,In_693,In_452);
nand U1067 (N_1067,In_3251,In_4569);
xnor U1068 (N_1068,In_264,In_1999);
nor U1069 (N_1069,In_3812,In_2161);
xnor U1070 (N_1070,In_2174,In_4130);
xnor U1071 (N_1071,In_3464,In_3828);
or U1072 (N_1072,In_1740,In_3725);
and U1073 (N_1073,In_3362,In_393);
and U1074 (N_1074,In_1003,In_3229);
nand U1075 (N_1075,In_3524,In_1368);
and U1076 (N_1076,In_1855,In_704);
xor U1077 (N_1077,In_2887,In_920);
and U1078 (N_1078,In_2889,In_1801);
nor U1079 (N_1079,In_1734,In_2607);
nor U1080 (N_1080,In_1790,In_1827);
nand U1081 (N_1081,In_3650,In_3110);
nor U1082 (N_1082,In_1686,In_4713);
and U1083 (N_1083,In_3674,In_4304);
and U1084 (N_1084,In_1872,In_2400);
and U1085 (N_1085,In_2585,In_3612);
nand U1086 (N_1086,In_446,In_4424);
or U1087 (N_1087,In_2464,In_1560);
nor U1088 (N_1088,In_3965,In_3098);
xnor U1089 (N_1089,In_104,In_654);
xor U1090 (N_1090,In_603,In_3351);
nor U1091 (N_1091,In_4377,In_4876);
nand U1092 (N_1092,In_4801,In_3543);
nor U1093 (N_1093,In_1576,In_1935);
nor U1094 (N_1094,In_3899,In_3703);
nand U1095 (N_1095,In_4171,In_1);
or U1096 (N_1096,In_2690,In_4414);
nand U1097 (N_1097,In_1655,In_3807);
and U1098 (N_1098,In_4136,In_3969);
xnor U1099 (N_1099,In_3105,In_4508);
or U1100 (N_1100,In_4555,In_458);
and U1101 (N_1101,In_703,In_3211);
nand U1102 (N_1102,In_4865,In_1426);
xnor U1103 (N_1103,In_4011,In_2073);
nand U1104 (N_1104,In_2679,In_685);
and U1105 (N_1105,In_3934,In_3274);
or U1106 (N_1106,In_3047,In_683);
nor U1107 (N_1107,In_2195,In_4016);
nor U1108 (N_1108,In_4190,In_1565);
or U1109 (N_1109,In_2666,In_4673);
and U1110 (N_1110,In_4420,In_378);
and U1111 (N_1111,In_714,In_2650);
and U1112 (N_1112,In_456,In_4717);
xor U1113 (N_1113,In_4379,In_844);
nor U1114 (N_1114,In_1759,In_4363);
nand U1115 (N_1115,In_2755,In_3433);
nor U1116 (N_1116,In_3259,In_516);
xor U1117 (N_1117,In_4329,In_1767);
nand U1118 (N_1118,In_3667,In_4582);
or U1119 (N_1119,In_3101,In_2731);
nand U1120 (N_1120,In_3028,In_2542);
or U1121 (N_1121,In_2135,In_209);
nor U1122 (N_1122,In_3819,In_4123);
nand U1123 (N_1123,In_344,In_2989);
xnor U1124 (N_1124,In_1162,In_2212);
and U1125 (N_1125,In_2239,In_1907);
or U1126 (N_1126,In_2732,In_1346);
nor U1127 (N_1127,In_2160,In_3556);
nor U1128 (N_1128,In_249,In_4892);
or U1129 (N_1129,In_3438,In_3713);
or U1130 (N_1130,In_1173,In_2830);
or U1131 (N_1131,In_2269,In_3071);
or U1132 (N_1132,In_1459,In_3167);
and U1133 (N_1133,In_3634,In_3384);
and U1134 (N_1134,In_2988,In_2038);
nor U1135 (N_1135,In_629,In_2926);
nor U1136 (N_1136,In_4690,In_2564);
nor U1137 (N_1137,In_201,In_4729);
xnor U1138 (N_1138,In_4523,In_2454);
or U1139 (N_1139,In_2981,In_1374);
nand U1140 (N_1140,In_733,In_2436);
or U1141 (N_1141,In_1616,In_1388);
or U1142 (N_1142,In_1607,In_633);
xor U1143 (N_1143,In_3963,In_2519);
or U1144 (N_1144,In_1634,In_1922);
xor U1145 (N_1145,In_1403,In_4691);
nor U1146 (N_1146,In_2546,In_17);
nor U1147 (N_1147,In_3512,In_529);
xor U1148 (N_1148,In_2700,In_4207);
nor U1149 (N_1149,In_4856,In_3448);
nor U1150 (N_1150,In_354,In_4230);
and U1151 (N_1151,In_765,In_2864);
xor U1152 (N_1152,In_902,In_570);
and U1153 (N_1153,In_3794,In_422);
xor U1154 (N_1154,In_2554,In_4427);
nand U1155 (N_1155,In_58,In_1029);
xnor U1156 (N_1156,In_2963,In_1732);
xnor U1157 (N_1157,In_150,In_4143);
xnor U1158 (N_1158,In_2916,In_2106);
or U1159 (N_1159,In_2032,In_3);
nand U1160 (N_1160,In_4708,In_3314);
xor U1161 (N_1161,In_4975,In_4817);
xnor U1162 (N_1162,In_4258,In_1696);
or U1163 (N_1163,In_2238,In_525);
or U1164 (N_1164,In_2768,In_2598);
xor U1165 (N_1165,In_4879,In_2014);
and U1166 (N_1166,In_1702,In_3178);
nand U1167 (N_1167,In_871,In_3516);
and U1168 (N_1168,In_3200,In_527);
nor U1169 (N_1169,In_4179,In_1589);
xnor U1170 (N_1170,In_3189,In_3640);
nand U1171 (N_1171,In_4940,In_4437);
nand U1172 (N_1172,In_1675,In_1746);
and U1173 (N_1173,In_4319,In_4527);
nor U1174 (N_1174,In_2548,In_4645);
xor U1175 (N_1175,In_1654,In_1710);
nand U1176 (N_1176,In_3665,In_4846);
nor U1177 (N_1177,In_3428,In_2155);
xnor U1178 (N_1178,In_2908,In_3302);
nand U1179 (N_1179,In_4781,In_2890);
nor U1180 (N_1180,In_3872,In_2582);
nand U1181 (N_1181,In_445,In_30);
xor U1182 (N_1182,In_2877,In_926);
or U1183 (N_1183,In_4933,In_2974);
or U1184 (N_1184,In_2781,In_686);
nor U1185 (N_1185,In_2741,In_4821);
and U1186 (N_1186,In_246,In_3810);
and U1187 (N_1187,In_4339,In_798);
nand U1188 (N_1188,In_4952,In_2168);
and U1189 (N_1189,In_2255,In_1606);
nor U1190 (N_1190,In_4914,In_635);
nand U1191 (N_1191,In_4726,In_3728);
and U1192 (N_1192,In_2404,In_4055);
nor U1193 (N_1193,In_1643,In_4270);
and U1194 (N_1194,In_3526,In_136);
or U1195 (N_1195,In_4903,In_809);
xnor U1196 (N_1196,In_3470,In_881);
nand U1197 (N_1197,In_3706,In_127);
nand U1198 (N_1198,In_3536,In_2560);
nor U1199 (N_1199,In_2166,In_490);
nor U1200 (N_1200,In_945,In_496);
xnor U1201 (N_1201,In_927,In_915);
nor U1202 (N_1202,In_3642,In_4686);
nor U1203 (N_1203,In_2720,In_2440);
nor U1204 (N_1204,In_138,In_3719);
and U1205 (N_1205,In_134,In_1150);
xnor U1206 (N_1206,In_505,In_3360);
or U1207 (N_1207,In_4922,In_48);
xor U1208 (N_1208,In_302,In_606);
nor U1209 (N_1209,In_1133,In_70);
nor U1210 (N_1210,In_4782,In_3944);
or U1211 (N_1211,In_1912,In_3031);
nand U1212 (N_1212,In_2316,In_1869);
and U1213 (N_1213,In_3263,In_2345);
and U1214 (N_1214,In_800,In_2423);
and U1215 (N_1215,In_4282,In_1418);
and U1216 (N_1216,In_4742,In_1101);
xor U1217 (N_1217,In_700,In_3431);
xor U1218 (N_1218,In_3059,In_674);
nor U1219 (N_1219,In_3417,In_4203);
nor U1220 (N_1220,In_2307,In_1518);
xor U1221 (N_1221,In_2738,In_1493);
nand U1222 (N_1222,In_1417,In_877);
nand U1223 (N_1223,In_4567,In_579);
or U1224 (N_1224,In_4896,In_3156);
nand U1225 (N_1225,In_1687,In_3497);
and U1226 (N_1226,In_612,In_1733);
nand U1227 (N_1227,In_184,In_4937);
xor U1228 (N_1228,In_4625,In_991);
and U1229 (N_1229,In_1152,In_3213);
nor U1230 (N_1230,In_4965,In_3187);
xor U1231 (N_1231,In_1370,In_2086);
and U1232 (N_1232,In_636,In_3306);
or U1233 (N_1233,In_269,In_2427);
and U1234 (N_1234,In_2871,In_3871);
and U1235 (N_1235,In_2444,In_2969);
nor U1236 (N_1236,In_4252,In_1138);
xnor U1237 (N_1237,In_2902,In_3800);
nand U1238 (N_1238,In_1949,In_4973);
nand U1239 (N_1239,In_2016,In_4905);
nand U1240 (N_1240,In_391,In_2338);
nand U1241 (N_1241,In_4764,In_2064);
nand U1242 (N_1242,In_4678,In_4289);
nand U1243 (N_1243,In_2125,In_3100);
or U1244 (N_1244,In_3864,In_56);
nand U1245 (N_1245,In_707,In_3739);
xor U1246 (N_1246,In_148,In_3223);
xnor U1247 (N_1247,In_3774,In_3967);
xor U1248 (N_1248,In_1047,In_4345);
nor U1249 (N_1249,In_542,In_709);
and U1250 (N_1250,In_1516,In_965);
xor U1251 (N_1251,In_1319,In_4811);
or U1252 (N_1252,In_3226,In_1272);
and U1253 (N_1253,In_1845,In_822);
or U1254 (N_1254,In_3481,In_3923);
and U1255 (N_1255,In_2994,In_3172);
nor U1256 (N_1256,In_2433,In_1249);
or U1257 (N_1257,In_829,In_1320);
and U1258 (N_1258,In_3951,In_2001);
nand U1259 (N_1259,In_1006,In_2204);
xor U1260 (N_1260,In_4027,In_1359);
nand U1261 (N_1261,In_4605,In_4579);
and U1262 (N_1262,In_1994,In_1091);
nor U1263 (N_1263,In_1605,In_696);
xor U1264 (N_1264,In_3830,In_1672);
xnor U1265 (N_1265,In_4509,In_607);
xnor U1266 (N_1266,In_180,In_4428);
xnor U1267 (N_1267,In_2021,In_55);
nor U1268 (N_1268,In_4228,In_49);
nor U1269 (N_1269,In_2932,In_2124);
nor U1270 (N_1270,In_202,In_1646);
nor U1271 (N_1271,In_2191,In_4906);
or U1272 (N_1272,In_2904,In_4456);
xor U1273 (N_1273,In_2236,In_4002);
or U1274 (N_1274,In_837,In_4877);
nor U1275 (N_1275,In_1357,In_665);
xnor U1276 (N_1276,In_892,In_3503);
xnor U1277 (N_1277,In_2529,In_146);
xor U1278 (N_1278,In_513,In_4489);
nand U1279 (N_1279,In_4565,In_3699);
nand U1280 (N_1280,In_2894,In_3700);
or U1281 (N_1281,In_4133,In_4483);
and U1282 (N_1282,In_808,In_1226);
and U1283 (N_1283,In_2599,In_1813);
or U1284 (N_1284,In_2923,In_162);
or U1285 (N_1285,In_1651,In_1640);
xnor U1286 (N_1286,In_3305,In_3957);
nand U1287 (N_1287,In_1899,In_1979);
nand U1288 (N_1288,In_1649,In_2003);
and U1289 (N_1289,In_3761,In_2637);
nand U1290 (N_1290,In_4822,In_1005);
xor U1291 (N_1291,In_4663,In_930);
nor U1292 (N_1292,In_1453,In_4360);
nand U1293 (N_1293,In_1180,In_4773);
nor U1294 (N_1294,In_861,In_4269);
or U1295 (N_1295,In_819,In_1069);
xor U1296 (N_1296,In_424,In_4286);
nor U1297 (N_1297,In_3277,In_4950);
xor U1298 (N_1298,In_3696,In_1148);
nand U1299 (N_1299,In_3048,In_332);
nor U1300 (N_1300,In_2337,In_3344);
or U1301 (N_1301,In_2060,In_1543);
and U1302 (N_1302,In_1303,In_3169);
nor U1303 (N_1303,In_543,In_2167);
xnor U1304 (N_1304,In_2669,In_1115);
xor U1305 (N_1305,In_1307,In_2641);
nand U1306 (N_1306,In_4331,In_4602);
nand U1307 (N_1307,In_3891,In_1189);
nand U1308 (N_1308,In_3493,In_1586);
nand U1309 (N_1309,In_4727,In_3056);
and U1310 (N_1310,In_1094,In_3298);
or U1311 (N_1311,In_4184,In_192);
nand U1312 (N_1312,In_4144,In_3032);
or U1313 (N_1313,In_4495,In_4053);
nand U1314 (N_1314,In_2771,In_1559);
or U1315 (N_1315,In_2903,In_1917);
and U1316 (N_1316,In_3746,In_1208);
or U1317 (N_1317,In_2045,In_3008);
nand U1318 (N_1318,In_1985,In_771);
nor U1319 (N_1319,In_957,In_4956);
and U1320 (N_1320,In_1823,In_1263);
xor U1321 (N_1321,In_1202,In_2595);
and U1322 (N_1322,In_352,In_4108);
nand U1323 (N_1323,In_4072,In_167);
or U1324 (N_1324,In_4658,In_3762);
and U1325 (N_1325,In_2760,In_3270);
and U1326 (N_1326,In_3507,In_958);
nand U1327 (N_1327,In_3383,In_4587);
and U1328 (N_1328,In_2363,In_1906);
and U1329 (N_1329,In_2284,In_1271);
nor U1330 (N_1330,In_879,In_3726);
xnor U1331 (N_1331,In_541,In_775);
or U1332 (N_1332,In_3510,In_2046);
xnor U1333 (N_1333,In_3577,In_4850);
nand U1334 (N_1334,In_2565,In_3756);
xor U1335 (N_1335,In_4327,In_3971);
nor U1336 (N_1336,In_1927,In_2805);
xnor U1337 (N_1337,In_4003,In_4875);
or U1338 (N_1338,In_1045,In_2568);
and U1339 (N_1339,In_2438,In_245);
xor U1340 (N_1340,In_1995,In_4550);
nor U1341 (N_1341,In_3611,In_2321);
or U1342 (N_1342,In_2232,In_1594);
nand U1343 (N_1343,In_2586,In_2225);
and U1344 (N_1344,In_4422,In_1602);
nor U1345 (N_1345,In_3946,In_3678);
nand U1346 (N_1346,In_3598,In_4628);
or U1347 (N_1347,In_4572,In_1898);
and U1348 (N_1348,In_4870,In_3257);
xor U1349 (N_1349,In_341,In_274);
and U1350 (N_1350,In_1472,In_794);
or U1351 (N_1351,In_238,In_67);
and U1352 (N_1352,In_1399,In_3308);
nand U1353 (N_1353,In_1442,In_141);
nor U1354 (N_1354,In_2097,In_4262);
nand U1355 (N_1355,In_80,In_1305);
nor U1356 (N_1356,In_401,In_940);
xnor U1357 (N_1357,In_426,In_874);
and U1358 (N_1358,In_617,In_3629);
and U1359 (N_1359,In_2192,In_3863);
or U1360 (N_1360,In_4800,In_2039);
nor U1361 (N_1361,In_3275,In_4955);
nor U1362 (N_1362,In_4352,In_375);
or U1363 (N_1363,In_2083,In_3552);
nand U1364 (N_1364,In_1116,In_442);
nor U1365 (N_1365,In_3160,In_16);
xnor U1366 (N_1366,In_1258,In_1984);
and U1367 (N_1367,In_3902,In_1940);
xnor U1368 (N_1368,In_102,In_2804);
and U1369 (N_1369,In_3295,In_1456);
or U1370 (N_1370,In_4295,In_4601);
or U1371 (N_1371,In_2553,In_363);
and U1372 (N_1372,In_1348,In_2220);
and U1373 (N_1373,In_1566,In_3658);
nand U1374 (N_1374,In_3414,In_1887);
nor U1375 (N_1375,In_1577,In_4029);
xor U1376 (N_1376,In_2140,In_63);
nand U1377 (N_1377,In_4772,In_43);
xor U1378 (N_1378,In_1611,In_622);
and U1379 (N_1379,In_600,In_2243);
or U1380 (N_1380,In_3698,In_4291);
nand U1381 (N_1381,In_1630,In_1743);
nor U1382 (N_1382,In_4116,In_3555);
xnor U1383 (N_1383,In_1108,In_3952);
nand U1384 (N_1384,In_2492,In_1064);
xor U1385 (N_1385,In_3291,In_51);
nor U1386 (N_1386,In_1410,In_1217);
xor U1387 (N_1387,In_2340,In_3987);
and U1388 (N_1388,In_3287,In_910);
and U1389 (N_1389,In_2497,In_4292);
and U1390 (N_1390,In_2881,In_1030);
nor U1391 (N_1391,In_2687,In_3148);
nand U1392 (N_1392,In_569,In_208);
xor U1393 (N_1393,In_1901,In_1919);
or U1394 (N_1394,In_1128,In_2763);
and U1395 (N_1395,In_1145,In_3964);
xnor U1396 (N_1396,In_4249,In_1419);
nor U1397 (N_1397,In_1796,In_1477);
and U1398 (N_1398,In_3091,In_1054);
or U1399 (N_1399,In_4723,In_2301);
xor U1400 (N_1400,In_1479,In_1893);
xor U1401 (N_1401,In_76,In_4670);
and U1402 (N_1402,In_4382,In_1729);
and U1403 (N_1403,In_1360,In_4948);
nand U1404 (N_1404,In_3723,In_4882);
nand U1405 (N_1405,In_1300,In_2715);
or U1406 (N_1406,In_3978,In_1206);
nand U1407 (N_1407,In_4485,In_3565);
and U1408 (N_1408,In_2480,In_1191);
and U1409 (N_1409,In_4803,In_3641);
or U1410 (N_1410,In_1838,In_3233);
xnor U1411 (N_1411,In_2328,In_430);
nand U1412 (N_1412,In_4604,In_2413);
nand U1413 (N_1413,In_1384,In_1437);
xor U1414 (N_1414,In_3266,In_4140);
or U1415 (N_1415,In_994,In_1020);
or U1416 (N_1416,In_2533,In_2593);
nand U1417 (N_1417,In_1836,In_1728);
nand U1418 (N_1418,In_1485,In_1711);
and U1419 (N_1419,In_1245,In_2727);
nor U1420 (N_1420,In_3862,In_2057);
and U1421 (N_1421,In_4466,In_499);
and U1422 (N_1422,In_3183,In_40);
nand U1423 (N_1423,In_2836,In_2043);
or U1424 (N_1424,In_3875,In_3407);
nor U1425 (N_1425,In_3975,In_2975);
nand U1426 (N_1426,In_4154,In_4591);
nand U1427 (N_1427,In_3072,In_1062);
and U1428 (N_1428,In_3320,In_4626);
xnor U1429 (N_1429,In_2217,In_908);
xnor U1430 (N_1430,In_4754,In_2079);
and U1431 (N_1431,In_4232,In_2412);
and U1432 (N_1432,In_4322,In_1904);
and U1433 (N_1433,In_3527,In_3078);
and U1434 (N_1434,In_2704,In_1423);
nor U1435 (N_1435,In_4939,In_2774);
nor U1436 (N_1436,In_2838,In_149);
nor U1437 (N_1437,In_4434,In_287);
or U1438 (N_1438,In_3469,In_2384);
or U1439 (N_1439,In_1386,In_20);
and U1440 (N_1440,In_1235,In_1806);
or U1441 (N_1441,In_342,In_297);
or U1442 (N_1442,In_560,In_1689);
nand U1443 (N_1443,In_3055,In_2692);
xor U1444 (N_1444,In_1535,In_4211);
nor U1445 (N_1445,In_3959,In_4751);
and U1446 (N_1446,In_1444,In_1876);
xor U1447 (N_1447,In_1155,In_255);
or U1448 (N_1448,In_645,In_1503);
and U1449 (N_1449,In_2488,In_2386);
nor U1450 (N_1450,In_4860,In_2208);
or U1451 (N_1451,In_1227,In_982);
nand U1452 (N_1452,In_2646,In_3463);
nor U1453 (N_1453,In_4761,In_2414);
or U1454 (N_1454,In_571,In_1690);
xnor U1455 (N_1455,In_75,In_592);
and U1456 (N_1456,In_823,In_3958);
or U1457 (N_1457,In_1093,In_3592);
nor U1458 (N_1458,In_2893,In_3331);
or U1459 (N_1459,In_1816,In_3210);
xor U1460 (N_1460,In_1229,In_2638);
nand U1461 (N_1461,In_796,In_1014);
nand U1462 (N_1462,In_3321,In_4017);
nor U1463 (N_1463,In_1102,In_3040);
or U1464 (N_1464,In_4297,In_555);
nand U1465 (N_1465,In_199,In_1840);
and U1466 (N_1466,In_3689,In_4076);
or U1467 (N_1467,In_2694,In_2068);
xnor U1468 (N_1468,In_1491,In_4806);
nor U1469 (N_1469,In_684,In_3542);
or U1470 (N_1470,In_3355,In_640);
or U1471 (N_1471,In_2701,In_4467);
and U1472 (N_1472,In_130,In_2577);
and U1473 (N_1473,In_2876,In_1522);
nor U1474 (N_1474,In_551,In_4644);
or U1475 (N_1475,In_1688,In_1401);
and U1476 (N_1476,In_4268,In_898);
nor U1477 (N_1477,In_766,In_4351);
xnor U1478 (N_1478,In_1088,In_377);
and U1479 (N_1479,In_1547,In_1037);
and U1480 (N_1480,In_1295,In_2985);
nor U1481 (N_1481,In_4880,In_4961);
xor U1482 (N_1482,In_3432,In_2477);
nor U1483 (N_1483,In_2817,In_3020);
or U1484 (N_1484,In_4878,In_4005);
or U1485 (N_1485,In_4452,In_706);
and U1486 (N_1486,In_273,In_4196);
and U1487 (N_1487,In_389,In_4073);
nor U1488 (N_1488,In_3673,In_2680);
nor U1489 (N_1489,In_3472,In_1312);
or U1490 (N_1490,In_3778,In_4636);
nor U1491 (N_1491,In_2681,In_481);
xnor U1492 (N_1492,In_1652,In_3888);
nor U1493 (N_1493,In_2909,In_2351);
nand U1494 (N_1494,In_231,In_2411);
nor U1495 (N_1495,In_4504,In_3386);
xor U1496 (N_1496,In_4311,In_4661);
and U1497 (N_1497,In_4180,In_3284);
or U1498 (N_1498,In_2921,In_2445);
nand U1499 (N_1499,In_4823,In_2841);
nor U1500 (N_1500,In_4967,In_2104);
nor U1501 (N_1501,In_4120,In_526);
xor U1502 (N_1502,In_3582,In_4167);
nand U1503 (N_1503,In_2706,In_669);
xnor U1504 (N_1504,In_3473,In_3677);
nand U1505 (N_1505,In_4810,In_3132);
nand U1506 (N_1506,In_3366,In_1915);
nor U1507 (N_1507,In_4163,In_4131);
nor U1508 (N_1508,In_3109,In_3421);
xor U1509 (N_1509,In_4021,In_659);
or U1510 (N_1510,In_1367,In_4578);
or U1511 (N_1511,In_986,In_2141);
nand U1512 (N_1512,In_3567,In_2461);
nand U1513 (N_1513,In_953,In_2470);
nand U1514 (N_1514,In_1932,In_3389);
or U1515 (N_1515,In_666,In_4977);
nor U1516 (N_1516,In_2142,In_2733);
and U1517 (N_1517,In_1626,In_4059);
and U1518 (N_1518,In_2117,In_3346);
or U1519 (N_1519,In_294,In_1911);
nor U1520 (N_1520,In_764,In_3896);
nor U1521 (N_1521,In_1439,In_2875);
xor U1522 (N_1522,In_1063,In_2175);
or U1523 (N_1523,In_4225,In_3396);
nor U1524 (N_1524,In_4813,In_1246);
nor U1525 (N_1525,In_306,In_313);
nor U1526 (N_1526,In_4307,In_1769);
xor U1527 (N_1527,In_1738,In_740);
and U1528 (N_1528,In_4148,In_125);
nor U1529 (N_1529,In_1561,In_988);
nor U1530 (N_1530,In_42,In_3529);
nor U1531 (N_1531,In_1595,In_265);
nand U1532 (N_1532,In_3089,In_221);
xnor U1533 (N_1533,In_4316,In_3268);
nand U1534 (N_1534,In_4413,In_1449);
and U1535 (N_1535,In_270,In_3133);
or U1536 (N_1536,In_2693,In_946);
and U1537 (N_1537,In_1154,In_4740);
and U1538 (N_1538,In_4622,In_351);
and U1539 (N_1539,In_3573,In_790);
or U1540 (N_1540,In_4915,In_3037);
xor U1541 (N_1541,In_2421,In_4235);
nand U1542 (N_1542,In_2177,In_4052);
and U1543 (N_1543,In_2575,In_1109);
xor U1544 (N_1544,In_4461,In_3541);
or U1545 (N_1545,In_888,In_3294);
or U1546 (N_1546,In_474,In_29);
and U1547 (N_1547,In_4219,In_3844);
nand U1548 (N_1548,In_4224,In_69);
or U1549 (N_1549,In_557,In_4109);
nand U1550 (N_1550,In_2867,In_3885);
xnor U1551 (N_1551,In_1598,In_1977);
nor U1552 (N_1552,In_3624,In_2283);
or U1553 (N_1553,In_4756,In_1554);
xnor U1554 (N_1554,In_4374,In_4188);
nand U1555 (N_1555,In_2998,In_2110);
and U1556 (N_1556,In_4899,In_3075);
xnor U1557 (N_1557,In_3586,In_2291);
or U1558 (N_1558,In_38,In_566);
nor U1559 (N_1559,In_461,In_4221);
nand U1560 (N_1560,In_2634,In_2130);
nand U1561 (N_1561,In_3455,In_3900);
xnor U1562 (N_1562,In_4146,In_4090);
or U1563 (N_1563,In_564,In_3572);
nor U1564 (N_1564,In_3002,In_3441);
nand U1565 (N_1565,In_2275,In_2965);
nor U1566 (N_1566,In_3898,In_90);
or U1567 (N_1567,In_3631,In_2780);
nor U1568 (N_1568,In_81,In_98);
and U1569 (N_1569,In_929,In_1753);
xor U1570 (N_1570,In_2764,In_4141);
and U1571 (N_1571,In_3977,In_1340);
nand U1572 (N_1572,In_119,In_1253);
xnor U1573 (N_1573,In_2603,In_813);
nor U1574 (N_1574,In_992,In_2534);
nand U1575 (N_1575,In_2839,In_4156);
and U1576 (N_1576,In_2559,In_4581);
xor U1577 (N_1577,In_2716,In_2456);
nand U1578 (N_1578,In_2753,In_2721);
or U1579 (N_1579,In_1164,In_68);
and U1580 (N_1580,In_4152,In_2270);
and U1581 (N_1581,In_711,In_2524);
nand U1582 (N_1582,In_880,In_1321);
nor U1583 (N_1583,In_1022,In_2794);
nand U1584 (N_1584,In_4220,In_3388);
nor U1585 (N_1585,In_4710,In_1925);
nand U1586 (N_1586,In_4367,In_1754);
xor U1587 (N_1587,In_777,In_2424);
nor U1588 (N_1588,In_4449,In_3517);
nand U1589 (N_1589,In_2606,In_1071);
nor U1590 (N_1590,In_3686,In_4474);
nor U1591 (N_1591,In_1548,In_3394);
xor U1592 (N_1592,In_1012,In_2837);
nor U1593 (N_1593,In_2113,In_1986);
nor U1594 (N_1594,In_3893,In_2520);
xnor U1595 (N_1595,In_4365,In_866);
or U1596 (N_1596,In_4525,In_4568);
xnor U1597 (N_1597,In_1683,In_1850);
nand U1598 (N_1598,In_3165,In_4946);
xnor U1599 (N_1599,In_540,In_1366);
or U1600 (N_1600,In_1844,In_1302);
and U1601 (N_1601,In_303,In_3776);
or U1602 (N_1602,In_2469,In_4659);
xor U1603 (N_1603,In_1134,In_2772);
or U1604 (N_1604,In_2264,In_522);
nor U1605 (N_1605,In_203,In_941);
or U1606 (N_1606,In_3792,In_2742);
nor U1607 (N_1607,In_369,In_649);
xor U1608 (N_1608,In_3149,In_549);
and U1609 (N_1609,In_13,In_1040);
xor U1610 (N_1610,In_1301,In_2633);
and U1611 (N_1611,In_3260,In_3849);
or U1612 (N_1612,In_1077,In_4464);
xnor U1613 (N_1613,In_3258,In_1761);
or U1614 (N_1614,In_3714,In_2037);
nand U1615 (N_1615,In_3710,In_3785);
xor U1616 (N_1616,In_4346,In_546);
xnor U1617 (N_1617,In_1969,In_57);
nand U1618 (N_1618,In_2325,In_2671);
nor U1619 (N_1619,In_2158,In_1679);
or U1620 (N_1620,In_942,In_3575);
or U1621 (N_1621,In_737,In_3130);
nand U1622 (N_1622,In_509,In_2782);
or U1623 (N_1623,In_4071,In_434);
xnor U1624 (N_1624,In_3073,In_3170);
nand U1625 (N_1625,In_3682,In_3948);
nor U1626 (N_1626,In_627,In_1648);
or U1627 (N_1627,In_284,In_4046);
xor U1628 (N_1628,In_2752,In_4714);
xnor U1629 (N_1629,In_4539,In_3596);
and U1630 (N_1630,In_3399,In_647);
nand U1631 (N_1631,In_3450,In_4598);
nor U1632 (N_1632,In_2843,In_770);
nor U1633 (N_1633,In_646,In_1737);
nor U1634 (N_1634,In_1523,In_3209);
nor U1635 (N_1635,In_1892,In_443);
nand U1636 (N_1636,In_3197,In_2823);
nor U1637 (N_1637,In_2252,In_608);
and U1638 (N_1638,In_3405,In_3546);
and U1639 (N_1639,In_3928,In_2968);
nor U1640 (N_1640,In_3299,In_1768);
and U1641 (N_1641,In_4164,In_601);
and U1642 (N_1642,In_3961,In_1853);
xnor U1643 (N_1643,In_4477,In_2808);
nand U1644 (N_1644,In_4254,In_84);
and U1645 (N_1645,In_3208,In_96);
and U1646 (N_1646,In_656,In_1035);
nand U1647 (N_1647,In_4479,In_2703);
nor U1648 (N_1648,In_1139,In_1210);
and U1649 (N_1649,In_4506,In_2105);
nor U1650 (N_1650,In_2617,In_4364);
nand U1651 (N_1651,In_2215,In_1224);
nor U1652 (N_1652,In_3818,In_1856);
and U1653 (N_1653,In_4848,In_2810);
or U1654 (N_1654,In_2044,In_2705);
nand U1655 (N_1655,In_3870,In_905);
or U1656 (N_1656,In_4208,In_2698);
or U1657 (N_1657,In_3409,In_3146);
nand U1658 (N_1658,In_1397,In_2476);
nor U1659 (N_1659,In_1861,In_1527);
nor U1660 (N_1660,In_160,In_1551);
xor U1661 (N_1661,In_2303,In_975);
xnor U1662 (N_1662,In_399,In_4333);
or U1663 (N_1663,In_4432,In_1846);
or U1664 (N_1664,In_1031,In_4534);
or U1665 (N_1665,In_4926,In_995);
and U1666 (N_1666,In_4960,In_2691);
or U1667 (N_1667,In_4881,In_1622);
and U1668 (N_1668,In_3418,In_4429);
nor U1669 (N_1669,In_1735,In_4101);
nand U1670 (N_1670,In_25,In_539);
nand U1671 (N_1671,In_3007,In_1085);
nor U1672 (N_1672,In_357,In_31);
xnor U1673 (N_1673,In_1287,In_1659);
and U1674 (N_1674,In_4193,In_917);
or U1675 (N_1675,In_2274,In_4079);
nor U1676 (N_1676,In_2356,In_4570);
and U1677 (N_1677,In_1280,In_2115);
and U1678 (N_1678,In_2087,In_4275);
nor U1679 (N_1679,In_2133,In_1509);
nand U1680 (N_1680,In_501,In_3408);
or U1681 (N_1681,In_3484,In_3341);
nand U1682 (N_1682,In_4294,In_3019);
xnor U1683 (N_1683,In_2521,In_3297);
xor U1684 (N_1684,In_2498,In_1903);
nor U1685 (N_1685,In_2915,In_3035);
nand U1686 (N_1686,In_239,In_1582);
or U1687 (N_1687,In_3980,In_2373);
and U1688 (N_1688,In_2164,In_2522);
xor U1689 (N_1689,In_168,In_4173);
and U1690 (N_1690,In_793,In_483);
nor U1691 (N_1691,In_545,In_2224);
or U1692 (N_1692,In_2827,In_675);
and U1693 (N_1693,In_838,In_2910);
nor U1694 (N_1694,In_165,In_2138);
nor U1695 (N_1695,In_3325,In_2108);
and U1696 (N_1696,In_4649,In_2547);
and U1697 (N_1697,In_3010,In_35);
nor U1698 (N_1698,In_3662,In_4718);
or U1699 (N_1699,In_1352,In_2661);
nand U1700 (N_1700,In_232,In_279);
or U1701 (N_1701,In_615,In_634);
and U1702 (N_1702,In_3788,In_4187);
nand U1703 (N_1703,In_597,In_2494);
xor U1704 (N_1704,In_4049,In_3018);
nor U1705 (N_1705,In_2653,In_3549);
or U1706 (N_1706,In_4829,In_1335);
or U1707 (N_1707,In_416,In_4356);
and U1708 (N_1708,In_4216,In_2856);
or U1709 (N_1709,In_3370,In_851);
nand U1710 (N_1710,In_3487,In_3240);
nand U1711 (N_1711,In_3153,In_4134);
or U1712 (N_1712,In_158,In_2530);
xnor U1713 (N_1713,In_4558,In_129);
nand U1714 (N_1714,In_3157,In_1411);
nor U1715 (N_1715,In_3813,In_3359);
nand U1716 (N_1716,In_3644,In_889);
xor U1717 (N_1717,In_4241,In_2667);
nor U1718 (N_1718,In_2526,In_482);
xnor U1719 (N_1719,In_122,In_3378);
or U1720 (N_1720,In_2471,In_3743);
nor U1721 (N_1721,In_1669,In_3832);
nand U1722 (N_1722,In_107,In_3901);
nand U1723 (N_1723,In_4110,In_3446);
xor U1724 (N_1724,In_4435,In_1584);
or U1725 (N_1725,In_364,In_2002);
nor U1726 (N_1726,In_961,In_262);
xnor U1727 (N_1727,In_806,In_2309);
or U1728 (N_1728,In_3742,In_1873);
nor U1729 (N_1729,In_3637,In_1415);
nor U1730 (N_1730,In_1330,In_1521);
xor U1731 (N_1731,In_319,In_214);
xor U1732 (N_1732,In_493,In_3164);
xor U1733 (N_1733,In_1177,In_1968);
nand U1734 (N_1734,In_2885,In_1785);
and U1735 (N_1735,In_4178,In_862);
nand U1736 (N_1736,In_2952,In_1544);
nor U1737 (N_1737,In_670,In_2616);
nand U1738 (N_1738,In_3918,In_2054);
xnor U1739 (N_1739,In_3518,In_4809);
xnor U1740 (N_1740,In_4693,In_2428);
xnor U1741 (N_1741,In_3243,In_4246);
and U1742 (N_1742,In_2067,In_3307);
xnor U1743 (N_1743,In_943,In_4703);
or U1744 (N_1744,In_886,In_2852);
or U1745 (N_1745,In_77,In_1515);
or U1746 (N_1746,In_628,In_2879);
xor U1747 (N_1747,In_679,In_21);
or U1748 (N_1748,In_845,In_968);
or U1749 (N_1749,In_4126,In_3664);
nor U1750 (N_1750,In_230,In_2528);
and U1751 (N_1751,In_3440,In_2360);
nand U1752 (N_1752,In_4695,In_3303);
or U1753 (N_1753,In_2029,In_427);
and U1754 (N_1754,In_1323,In_1427);
or U1755 (N_1755,In_441,In_3722);
xor U1756 (N_1756,In_2936,In_4768);
and U1757 (N_1757,In_3380,In_2406);
nor U1758 (N_1758,In_4533,In_1570);
nand U1759 (N_1759,In_2639,In_2397);
and U1760 (N_1760,In_3381,In_573);
or U1761 (N_1761,In_1885,In_4607);
nand U1762 (N_1762,In_3597,In_3021);
and U1763 (N_1763,In_477,In_503);
or U1764 (N_1764,In_4929,In_507);
nand U1765 (N_1765,In_3489,In_4954);
or U1766 (N_1766,In_2629,In_1188);
and U1767 (N_1767,In_1355,In_2778);
and U1768 (N_1768,In_3485,In_1389);
xor U1769 (N_1769,In_4789,In_1390);
xor U1770 (N_1770,In_2597,In_1550);
xnor U1771 (N_1771,In_2730,In_2766);
and U1772 (N_1772,In_605,In_937);
and U1773 (N_1773,In_242,In_3466);
nor U1774 (N_1774,In_3468,In_3910);
and U1775 (N_1775,In_3515,In_1176);
xor U1776 (N_1776,In_338,In_4446);
or U1777 (N_1777,In_3124,In_2072);
or U1778 (N_1778,In_1332,In_4868);
xnor U1779 (N_1779,In_4984,In_3068);
xor U1780 (N_1780,In_3053,In_3877);
nor U1781 (N_1781,In_3520,In_3269);
or U1782 (N_1782,In_1789,In_4302);
xnor U1783 (N_1783,In_3190,In_2707);
and U1784 (N_1784,In_1664,In_4540);
xor U1785 (N_1785,In_4838,In_1341);
and U1786 (N_1786,In_972,In_869);
and U1787 (N_1787,In_1345,In_3505);
and U1788 (N_1788,In_4480,In_3159);
and U1789 (N_1789,In_1337,In_655);
or U1790 (N_1790,In_638,In_676);
nand U1791 (N_1791,In_731,In_4271);
or U1792 (N_1792,In_2734,In_1466);
nor U1793 (N_1793,In_4912,In_1662);
nor U1794 (N_1794,In_4309,In_3897);
nand U1795 (N_1795,In_857,In_3276);
and U1796 (N_1796,In_465,In_1065);
xor U1797 (N_1797,In_3281,In_1709);
and U1798 (N_1798,In_4696,In_3044);
nor U1799 (N_1799,In_4251,In_4921);
nand U1800 (N_1800,In_3836,In_2725);
or U1801 (N_1801,In_4958,In_4104);
xnor U1802 (N_1802,In_4797,In_4716);
and U1803 (N_1803,In_1440,In_1623);
and U1804 (N_1804,In_4869,In_698);
or U1805 (N_1805,In_1193,In_1804);
nand U1806 (N_1806,In_1178,In_1716);
or U1807 (N_1807,In_1344,In_2028);
xor U1808 (N_1808,In_903,In_1392);
xnor U1809 (N_1809,In_2434,In_4606);
nor U1810 (N_1810,In_3859,In_2118);
or U1811 (N_1811,In_4741,In_3457);
nand U1812 (N_1812,In_3393,In_1567);
nor U1813 (N_1813,In_3623,In_4735);
or U1814 (N_1814,In_217,In_1190);
or U1815 (N_1815,In_2295,In_484);
xnor U1816 (N_1816,In_1126,In_2107);
nand U1817 (N_1817,In_3721,In_3329);
nand U1818 (N_1818,In_2678,In_858);
or U1819 (N_1819,In_841,In_989);
and U1820 (N_1820,In_2983,In_4366);
nor U1821 (N_1821,In_747,In_1682);
nor U1822 (N_1822,In_4242,In_4057);
nand U1823 (N_1823,In_2330,In_1517);
and U1824 (N_1824,In_1395,In_3424);
nand U1825 (N_1825,In_999,In_2366);
or U1826 (N_1826,In_4459,In_2388);
or U1827 (N_1827,In_2645,In_2200);
and U1828 (N_1828,In_3765,In_34);
xnor U1829 (N_1829,In_289,In_3234);
nor U1830 (N_1830,In_4296,In_7);
xor U1831 (N_1831,In_2201,In_1542);
nor U1832 (N_1832,In_3467,In_2231);
nor U1833 (N_1833,In_3570,In_163);
nor U1834 (N_1834,In_4197,In_206);
xnor U1835 (N_1835,In_1639,In_1599);
and U1836 (N_1836,In_3051,In_4069);
xnor U1837 (N_1837,In_3283,In_1684);
xor U1838 (N_1838,In_3869,In_4510);
and U1839 (N_1839,In_1944,In_1358);
nand U1840 (N_1840,In_2159,In_4463);
or U1841 (N_1841,In_3878,In_2668);
nand U1842 (N_1842,In_4561,In_1373);
xnor U1843 (N_1843,In_2556,In_533);
and U1844 (N_1844,In_4666,In_2929);
or U1845 (N_1845,In_2743,In_39);
nand U1846 (N_1846,In_3003,In_3151);
nand U1847 (N_1847,In_1061,In_2465);
xnor U1848 (N_1848,In_3288,In_1579);
nor U1849 (N_1849,In_2583,In_3911);
nand U1850 (N_1850,In_3564,In_847);
nor U1851 (N_1851,In_3282,In_2022);
nor U1852 (N_1852,In_3745,In_3908);
or U1853 (N_1853,In_3147,In_89);
or U1854 (N_1854,In_1377,In_3343);
xor U1855 (N_1855,In_395,In_532);
xnor U1856 (N_1856,In_174,In_2928);
xor U1857 (N_1857,In_326,In_2640);
or U1858 (N_1858,In_87,In_1596);
and U1859 (N_1859,In_318,In_195);
nor U1860 (N_1860,In_1185,In_3883);
nand U1861 (N_1861,In_1660,In_417);
xor U1862 (N_1862,In_3985,In_1499);
nor U1863 (N_1863,In_4499,In_1043);
and U1864 (N_1864,In_1068,In_3578);
nor U1865 (N_1865,In_1160,In_4298);
or U1866 (N_1866,In_411,In_3820);
nor U1867 (N_1867,In_3482,In_4968);
nand U1868 (N_1868,In_997,In_980);
xnor U1869 (N_1869,In_1619,In_4974);
or U1870 (N_1870,In_2973,In_4623);
and U1871 (N_1871,In_1505,In_668);
or U1872 (N_1872,In_2148,In_4395);
or U1873 (N_1873,In_3771,In_2980);
xor U1874 (N_1874,In_791,In_4920);
or U1875 (N_1875,In_3955,In_4337);
or U1876 (N_1876,In_3561,In_4616);
or U1877 (N_1877,In_3272,In_2803);
or U1878 (N_1878,In_3162,In_3797);
and U1879 (N_1879,In_2203,In_899);
xor U1880 (N_1880,In_834,In_534);
nor U1881 (N_1881,In_2723,In_4312);
nor U1882 (N_1882,In_2007,In_2298);
nand U1883 (N_1883,In_1387,In_1839);
nand U1884 (N_1884,In_3248,In_3057);
nand U1885 (N_1885,In_1205,In_3367);
or U1886 (N_1886,In_3921,In_4889);
nand U1887 (N_1887,In_2052,In_4752);
nor U1888 (N_1888,In_4280,In_4441);
nor U1889 (N_1889,In_761,In_859);
xor U1890 (N_1890,In_2642,In_2499);
or U1891 (N_1891,In_3933,In_4019);
and U1892 (N_1892,In_2986,In_2379);
and U1893 (N_1893,In_4945,In_538);
nor U1894 (N_1894,In_2389,In_1285);
or U1895 (N_1895,In_4263,In_4259);
and U1896 (N_1896,In_743,In_1186);
nor U1897 (N_1897,In_460,In_2080);
xnor U1898 (N_1898,In_1278,In_4393);
xnor U1899 (N_1899,In_3231,In_310);
and U1900 (N_1900,In_1719,In_3445);
xor U1901 (N_1901,In_3311,In_3076);
or U1902 (N_1902,In_2625,In_2250);
nand U1903 (N_1903,In_4299,In_4980);
nor U1904 (N_1904,In_1383,In_593);
or U1905 (N_1905,In_1831,In_4183);
or U1906 (N_1906,In_1142,In_2241);
xor U1907 (N_1907,In_4160,In_4988);
nor U1908 (N_1908,In_4476,In_2971);
xnor U1909 (N_1909,In_4668,In_962);
or U1910 (N_1910,In_3490,In_3070);
xor U1911 (N_1911,In_738,In_4493);
or U1912 (N_1912,In_801,In_4857);
or U1913 (N_1913,In_1866,In_128);
or U1914 (N_1914,In_1492,In_2930);
xor U1915 (N_1915,In_412,In_1008);
nor U1916 (N_1916,In_3562,In_1613);
xnor U1917 (N_1917,In_506,In_1705);
nor U1918 (N_1918,In_2550,In_4917);
nor U1919 (N_1919,In_1408,In_3690);
and U1920 (N_1920,In_2552,In_200);
nor U1921 (N_1921,In_3625,In_1132);
xor U1922 (N_1922,In_473,In_2213);
nand U1923 (N_1923,In_4657,In_3521);
nand U1924 (N_1924,In_3808,In_2207);
and U1925 (N_1925,In_390,In_3221);
or U1926 (N_1926,In_240,In_3236);
nand U1927 (N_1927,In_2382,In_1676);
and U1928 (N_1928,In_2352,In_4033);
nor U1929 (N_1929,In_2033,In_602);
or U1930 (N_1930,In_4,In_2339);
nor U1931 (N_1931,In_400,In_3639);
nor U1932 (N_1932,In_2635,In_3357);
xnor U1933 (N_1933,In_1627,In_3851);
or U1934 (N_1934,In_2964,In_4664);
or U1935 (N_1935,In_1469,In_3501);
nand U1936 (N_1936,In_4549,In_978);
or U1937 (N_1937,In_252,In_3496);
nor U1938 (N_1938,In_3620,In_1019);
xnor U1939 (N_1939,In_4709,In_3798);
nand U1940 (N_1940,In_1867,In_4261);
xor U1941 (N_1941,In_2378,In_3155);
or U1942 (N_1942,In_3191,In_1562);
nand U1943 (N_1943,In_964,In_3716);
nand U1944 (N_1944,In_4599,In_1067);
nor U1945 (N_1945,In_1812,In_2954);
and U1946 (N_1946,In_3609,In_3879);
nor U1947 (N_1947,In_4783,In_1429);
xnor U1948 (N_1948,In_3998,In_4247);
nor U1949 (N_1949,In_1879,In_1909);
nor U1950 (N_1950,In_4105,In_4209);
nor U1951 (N_1951,In_783,In_3212);
and U1952 (N_1952,In_2900,In_4516);
nand U1953 (N_1953,In_4355,In_154);
and U1954 (N_1954,In_4215,In_2023);
or U1955 (N_1955,In_359,In_2205);
nor U1956 (N_1956,In_3062,In_687);
or U1957 (N_1957,In_680,In_1298);
and U1958 (N_1958,In_4433,In_1951);
xnor U1959 (N_1959,In_2785,In_1955);
nor U1960 (N_1960,In_4285,In_3915);
nor U1961 (N_1961,In_984,In_772);
nor U1962 (N_1962,In_2543,In_256);
nor U1963 (N_1963,In_521,In_176);
or U1964 (N_1964,In_2555,In_3491);
or U1965 (N_1965,In_37,In_4712);
nor U1966 (N_1966,In_2435,In_3685);
nor U1967 (N_1967,In_2938,In_1510);
xnor U1968 (N_1968,In_2041,In_1328);
or U1969 (N_1969,In_4192,In_143);
and U1970 (N_1970,In_3905,In_1137);
xnor U1971 (N_1971,In_3604,In_2071);
and U1972 (N_1972,In_3855,In_4839);
and U1973 (N_1973,In_720,In_4491);
and U1974 (N_1974,In_3815,In_183);
or U1975 (N_1975,In_583,In_4942);
xor U1976 (N_1976,In_3858,In_4411);
xnor U1977 (N_1977,In_4068,In_894);
nand U1978 (N_1978,In_1880,In_166);
nand U1979 (N_1979,In_2432,In_517);
or U1980 (N_1980,In_802,In_23);
xnor U1981 (N_1981,In_1480,In_1240);
nand U1982 (N_1982,In_1530,In_3806);
nand U1983 (N_1983,In_4031,In_1996);
or U1984 (N_1984,In_4835,In_1311);
or U1985 (N_1985,In_528,In_229);
nand U1986 (N_1986,In_878,In_243);
nor U1987 (N_1987,In_4799,In_828);
and U1988 (N_1988,In_3653,In_4034);
and U1989 (N_1989,In_1501,In_763);
xnor U1990 (N_1990,In_1828,In_1376);
nor U1991 (N_1991,In_1642,In_1257);
xnor U1992 (N_1992,In_3535,In_405);
or U1993 (N_1993,In_2809,In_2381);
or U1994 (N_1994,In_2541,In_2137);
and U1995 (N_1995,In_4532,In_2396);
or U1996 (N_1996,In_4620,In_3671);
nor U1997 (N_1997,In_4142,In_2419);
and U1998 (N_1998,In_4473,In_3012);
and U1999 (N_1999,In_1835,In_3847);
xor U2000 (N_2000,In_4585,In_1512);
nand U2001 (N_2001,In_32,In_3079);
nor U2002 (N_2002,In_1076,In_3782);
nor U2003 (N_2003,In_2618,In_1825);
xnor U2004 (N_2004,In_2385,In_2500);
or U2005 (N_2005,In_2294,In_3860);
or U2006 (N_2006,In_3557,In_2147);
xor U2007 (N_2007,In_2047,In_2322);
nor U2008 (N_2008,In_637,In_4750);
or U2009 (N_2009,In_2439,In_2624);
xor U2010 (N_2010,In_3701,In_1315);
nor U2011 (N_2011,In_1808,In_3456);
or U2012 (N_2012,In_4609,In_1924);
and U2013 (N_2013,In_4851,In_3177);
nor U2014 (N_2014,In_3606,In_3154);
xnor U2015 (N_2015,In_4911,In_4457);
or U2016 (N_2016,In_1870,In_188);
or U2017 (N_2017,In_2193,In_1541);
nor U2018 (N_2018,In_925,In_2505);
nor U2019 (N_2019,In_1279,In_2473);
nor U2020 (N_2020,In_4546,In_2670);
xor U2021 (N_2021,In_1580,In_2722);
and U2022 (N_2022,In_2481,In_1993);
nand U2023 (N_2023,In_1362,In_3423);
xnor U2024 (N_2024,In_4736,In_2253);
and U2025 (N_2025,In_3090,In_653);
or U2026 (N_2026,In_1324,In_3416);
or U2027 (N_2027,In_4274,In_3791);
nor U2028 (N_2028,In_2409,In_578);
xnor U2029 (N_2029,In_3670,In_178);
nand U2030 (N_2030,In_511,In_2114);
xnor U2031 (N_2031,In_690,In_4091);
nor U2032 (N_2032,In_1766,In_3430);
nor U2033 (N_2033,In_478,In_4000);
nand U2034 (N_2034,In_2557,In_729);
nand U2035 (N_2035,In_3809,In_2800);
xnor U2036 (N_2036,In_586,In_2401);
and U2037 (N_2037,In_1752,In_2844);
nand U2038 (N_2038,In_4155,In_1965);
nor U2039 (N_2039,In_959,In_552);
nand U2040 (N_2040,In_1481,In_4925);
or U2041 (N_2041,In_833,In_2009);
or U2042 (N_2042,In_1157,In_2350);
nor U2043 (N_2043,In_3480,In_210);
xnor U2044 (N_2044,In_1454,In_1198);
nor U2045 (N_2045,In_1778,In_3326);
nor U2046 (N_2046,In_2962,In_164);
nor U2047 (N_2047,In_1239,In_755);
and U2048 (N_2048,In_4397,In_2953);
xor U2049 (N_2049,In_1511,In_1436);
nand U2050 (N_2050,In_3779,In_4830);
or U2051 (N_2051,In_2260,In_3755);
and U2052 (N_2052,In_3867,In_4062);
nand U2053 (N_2053,In_2263,In_3134);
nor U2054 (N_2054,In_4497,In_949);
and U2055 (N_2055,In_1832,In_4930);
nand U2056 (N_2056,In_4831,In_1496);
and U2057 (N_2057,In_3986,In_4611);
xnor U2058 (N_2058,In_1950,In_2059);
xor U2059 (N_2059,In_4403,In_2008);
nand U2060 (N_2060,In_658,In_2513);
nand U2061 (N_2061,In_4978,In_4455);
nor U2062 (N_2062,In_324,In_4818);
or U2063 (N_2063,In_2898,In_3174);
xor U2064 (N_2064,In_2369,In_2);
xnor U2065 (N_2065,In_4236,In_664);
and U2066 (N_2066,In_2708,In_1981);
xor U2067 (N_2067,In_1715,In_502);
xor U2068 (N_2068,In_520,In_3680);
or U2069 (N_2069,In_4653,In_2156);
nor U2070 (N_2070,In_4560,In_4767);
and U2071 (N_2071,In_2941,In_1601);
or U2072 (N_2072,In_4478,In_2226);
xor U2073 (N_2073,In_2740,In_4528);
and U2074 (N_2074,In_4119,In_2697);
nor U2075 (N_2075,In_248,In_4547);
and U2076 (N_2076,In_73,In_1317);
and U2077 (N_2077,In_2648,In_751);
and U2078 (N_2078,In_1482,In_2713);
nand U2079 (N_2079,In_1075,In_715);
and U2080 (N_2080,In_2210,In_2237);
nor U2081 (N_2081,In_2308,In_3377);
or U2082 (N_2082,In_3962,In_433);
or U2083 (N_2083,In_789,In_2478);
nor U2084 (N_2084,In_2767,In_4776);
and U2085 (N_2085,In_295,In_584);
and U2086 (N_2086,In_126,In_3802);
nand U2087 (N_2087,In_1779,In_4421);
xnor U2088 (N_2088,In_3600,In_4749);
or U2089 (N_2089,In_2673,In_2026);
or U2090 (N_2090,In_1349,In_2632);
or U2091 (N_2091,In_8,In_2551);
nor U2092 (N_2092,In_3848,In_1978);
or U2093 (N_2093,In_3425,In_1334);
and U2094 (N_2094,In_4042,In_4416);
nand U2095 (N_2095,In_1961,In_4227);
nand U2096 (N_2096,In_1500,In_4498);
nand U2097 (N_2097,In_2431,In_2359);
nor U2098 (N_2098,In_2587,In_4983);
and U2099 (N_2099,In_2197,In_4387);
nand U2100 (N_2100,In_3922,In_406);
and U2101 (N_2101,In_778,In_3930);
nor U2102 (N_2102,In_1817,In_530);
xnor U2103 (N_2103,In_4807,In_4677);
or U2104 (N_2104,In_2790,In_1600);
and U2105 (N_2105,In_2951,In_3925);
nor U2106 (N_2106,In_4139,In_4198);
nand U2107 (N_2107,In_4593,In_884);
xnor U2108 (N_2108,In_169,In_397);
nor U2109 (N_2109,In_4556,In_94);
and U2110 (N_2110,In_2405,In_3974);
and U2111 (N_2111,In_1724,In_4562);
or U2112 (N_2112,In_1569,In_2085);
nor U2113 (N_2113,In_328,In_2442);
and U2114 (N_2114,In_4114,In_2858);
and U2115 (N_2115,In_2304,In_1431);
or U2116 (N_2116,In_3214,In_912);
xnor U2117 (N_2117,In_2604,In_744);
nand U2118 (N_2118,In_1826,In_1537);
nor U2119 (N_2119,In_4597,In_3767);
nand U2120 (N_2120,In_414,In_2144);
or U2121 (N_2121,In_1514,In_1297);
nand U2122 (N_2122,In_524,In_4762);
xor U2123 (N_2123,In_1591,In_4976);
nand U2124 (N_2124,In_2296,In_2664);
nand U2125 (N_2125,In_2786,In_333);
or U2126 (N_2126,In_2077,In_4971);
and U2127 (N_2127,In_1421,In_296);
and U2128 (N_2128,In_3318,In_4704);
or U2129 (N_2129,In_4092,In_124);
xor U2130 (N_2130,In_934,In_2091);
and U2131 (N_2131,In_4248,In_3737);
xnor U2132 (N_2132,In_3842,In_3338);
xnor U2133 (N_2133,In_1997,In_1967);
nor U2134 (N_2134,In_3731,In_1886);
xnor U2135 (N_2135,In_1821,In_1471);
or U2136 (N_2136,In_2326,In_198);
and U2137 (N_2137,In_4075,In_444);
nand U2138 (N_2138,In_701,In_1959);
or U2139 (N_2139,In_568,In_4849);
or U2140 (N_2140,In_4676,In_2845);
nand U2141 (N_2141,In_2828,In_3016);
nor U2142 (N_2142,In_1874,In_4043);
or U2143 (N_2143,In_2074,In_1203);
nand U2144 (N_2144,In_4334,In_768);
or U2145 (N_2145,In_3247,In_2594);
or U2146 (N_2146,In_4656,In_2058);
xnor U2147 (N_2147,In_1120,In_4392);
nand U2148 (N_2148,In_1849,In_1243);
xnor U2149 (N_2149,In_4780,In_3909);
or U2150 (N_2150,In_2300,In_4135);
xnor U2151 (N_2151,In_1653,In_3140);
nor U2152 (N_2152,In_4815,In_109);
xor U2153 (N_2153,In_191,In_1859);
nor U2154 (N_2154,In_3444,In_1678);
or U2155 (N_2155,In_3267,In_1084);
nor U2156 (N_2156,In_3789,In_3509);
nor U2157 (N_2157,In_950,In_4347);
nor U2158 (N_2158,In_22,In_4444);
nor U2159 (N_2159,In_2802,In_2450);
or U2160 (N_2160,In_4643,In_152);
nor U2161 (N_2161,In_224,In_922);
xnor U2162 (N_2162,In_140,In_4218);
xnor U2163 (N_2163,In_2111,In_1207);
or U2164 (N_2164,In_1107,In_3145);
and U2165 (N_2165,In_1027,In_1122);
nor U2166 (N_2166,In_3488,In_565);
nor U2167 (N_2167,In_3895,In_1498);
or U2168 (N_2168,In_2410,In_1524);
xnor U2169 (N_2169,In_1151,In_872);
nand U2170 (N_2170,In_4301,In_3461);
or U2171 (N_2171,In_1953,In_4650);
or U2172 (N_2172,In_4837,In_454);
nor U2173 (N_2173,In_3045,In_1197);
nand U2174 (N_2174,In_4482,In_2920);
and U2175 (N_2175,In_904,In_4010);
nor U2176 (N_2176,In_4722,In_3949);
nor U2177 (N_2177,In_2957,In_348);
xor U2178 (N_2178,In_948,In_2151);
xor U2179 (N_2179,In_928,In_4074);
or U2180 (N_2180,In_977,In_2605);
and U2181 (N_2181,In_3550,In_1744);
and U2182 (N_2182,In_620,In_1445);
xor U2183 (N_2183,In_1473,In_3422);
or U2184 (N_2184,In_913,In_2944);
nor U2185 (N_2185,In_4199,In_2370);
or U2186 (N_2186,In_1443,In_753);
nor U2187 (N_2187,In_998,In_1775);
nor U2188 (N_2188,In_2762,In_271);
xor U2189 (N_2189,In_1717,In_1080);
nor U2190 (N_2190,In_799,In_1121);
xnor U2191 (N_2191,In_1848,In_282);
or U2192 (N_2192,In_4008,In_361);
nor U2193 (N_2193,In_1048,In_575);
or U2194 (N_2194,In_3647,In_2729);
xor U2195 (N_2195,In_2180,In_1234);
nand U2196 (N_2196,In_1432,In_3583);
nand U2197 (N_2197,In_196,In_1086);
nand U2198 (N_2198,In_305,In_2336);
and U2199 (N_2199,In_1538,In_3770);
nor U2200 (N_2200,In_385,In_1400);
xnor U2201 (N_2201,In_3333,In_3217);
and U2202 (N_2202,In_3249,In_1988);
and U2203 (N_2203,In_1638,In_2333);
nor U2204 (N_2204,In_250,In_2289);
nand U2205 (N_2205,In_3471,In_773);
xnor U2206 (N_2206,In_1129,In_4652);
nor U2207 (N_2207,In_3924,In_2949);
xor U2208 (N_2208,In_3372,In_1111);
or U2209 (N_2209,In_3857,In_1379);
or U2210 (N_2210,In_4563,In_893);
nor U2211 (N_2211,In_2371,In_3991);
and U2212 (N_2212,In_300,In_2677);
nor U2213 (N_2213,In_463,In_2341);
xnor U2214 (N_2214,In_779,In_2272);
nor U2215 (N_2215,In_3136,In_713);
xnor U2216 (N_2216,In_4436,In_1699);
and U2217 (N_2217,In_4018,In_1583);
and U2218 (N_2218,In_1149,In_2383);
or U2219 (N_2219,In_3392,In_2674);
and U2220 (N_2220,In_1267,In_2134);
or U2221 (N_2221,In_4453,In_4181);
and U2222 (N_2222,In_3447,In_408);
xnor U2223 (N_2223,In_914,In_3811);
nand U2224 (N_2224,In_1549,In_4895);
xnor U2225 (N_2225,In_2588,In_2913);
nor U2226 (N_2226,In_2116,In_2950);
nor U2227 (N_2227,In_59,In_3605);
xnor U2228 (N_2228,In_4399,In_4113);
nor U2229 (N_2229,In_4129,In_3033);
nor U2230 (N_2230,In_3571,In_3080);
nor U2231 (N_2231,In_1066,In_4384);
nand U2232 (N_2232,In_2268,In_4836);
and U2233 (N_2233,In_1934,In_657);
and U2234 (N_2234,In_4796,In_421);
xnor U2235 (N_2235,In_4081,In_2251);
nor U2236 (N_2236,In_2540,In_3369);
xnor U2237 (N_2237,In_123,In_3579);
or U2238 (N_2238,In_3118,In_2323);
nand U2239 (N_2239,In_2619,In_1910);
and U2240 (N_2240,In_1268,In_4795);
xnor U2241 (N_2241,In_4987,In_1011);
xor U2242 (N_2242,In_449,In_4798);
xor U2243 (N_2243,In_717,In_187);
xor U2244 (N_2244,In_3672,In_4701);
nand U2245 (N_2245,In_2228,In_3508);
and U2246 (N_2246,In_2849,In_906);
nor U2247 (N_2247,In_2076,In_2094);
xnor U2248 (N_2248,In_350,In_2995);
nand U2249 (N_2249,In_1153,In_1083);
nand U2250 (N_2250,In_3342,In_1695);
and U2251 (N_2251,In_1209,In_3459);
or U2252 (N_2252,In_3404,In_3856);
nor U2253 (N_2253,In_3825,In_3976);
or U2254 (N_2254,In_4844,In_2662);
and U2255 (N_2255,In_2927,In_1531);
and U2256 (N_2256,In_3023,In_3256);
nand U2257 (N_2257,In_4854,In_677);
and U2258 (N_2258,In_1216,In_954);
or U2259 (N_2259,In_2334,In_1847);
or U2260 (N_2260,In_631,In_814);
and U2261 (N_2261,In_1974,In_1854);
xnor U2262 (N_2262,In_439,In_710);
nor U2263 (N_2263,In_882,In_719);
or U2264 (N_2264,In_616,In_1519);
or U2265 (N_2265,In_4358,In_3391);
xnor U2266 (N_2266,In_4036,In_2549);
xor U2267 (N_2267,In_1223,In_1691);
xor U2268 (N_2268,In_4576,In_3632);
nor U2269 (N_2269,In_547,In_253);
or U2270 (N_2270,In_3668,In_2466);
or U2271 (N_2271,In_4680,In_2185);
nor U2272 (N_2272,In_3992,In_4793);
nand U2273 (N_2273,In_1673,In_4390);
nor U2274 (N_2274,In_1788,In_1464);
nor U2275 (N_2275,In_619,In_4627);
and U2276 (N_2276,In_219,In_2931);
or U2277 (N_2277,In_1749,In_186);
xor U2278 (N_2278,In_2970,In_3304);
nand U2279 (N_2279,In_1771,In_1629);
xor U2280 (N_2280,In_4731,In_1621);
or U2281 (N_2281,In_3775,In_2862);
nor U2282 (N_2282,In_4137,In_1455);
nor U2283 (N_2283,In_1428,In_2672);
and U2284 (N_2284,In_2749,In_1230);
xnor U2285 (N_2285,In_3437,In_826);
nor U2286 (N_2286,In_4229,In_4380);
and U2287 (N_2287,In_1106,In_2216);
nand U2288 (N_2288,In_2959,In_4015);
nand U2289 (N_2289,In_2654,In_2656);
nand U2290 (N_2290,In_3046,In_4107);
nor U2291 (N_2291,In_309,In_4067);
and U2292 (N_2292,In_4902,In_2567);
or U2293 (N_2293,In_1452,In_3094);
xor U2294 (N_2294,In_1450,In_2907);
or U2295 (N_2295,In_4407,In_3332);
and U2296 (N_2296,In_2451,In_4412);
nor U2297 (N_2297,In_3144,In_233);
or U2298 (N_2298,In_741,In_3881);
xnor U2299 (N_2299,In_4632,In_2840);
and U2300 (N_2300,In_3906,In_336);
xor U2301 (N_2301,In_3085,In_3850);
or U2302 (N_2302,In_3999,In_2247);
or U2303 (N_2303,In_4551,In_1608);
and U2304 (N_2304,In_1714,In_2506);
and U2305 (N_2305,In_3184,In_1475);
nand U2306 (N_2306,In_2109,In_1325);
or U2307 (N_2307,In_1363,In_247);
nor U2308 (N_2308,In_2759,In_480);
or U2309 (N_2309,In_2277,In_139);
or U2310 (N_2310,In_3751,In_1461);
xor U2311 (N_2311,In_2999,In_4982);
and U2312 (N_2312,In_451,In_1868);
nor U2313 (N_2313,In_92,In_4943);
xor U2314 (N_2314,In_2776,In_558);
xor U2315 (N_2315,In_384,In_83);
nand U2316 (N_2316,In_4900,In_3339);
xor U2317 (N_2317,In_3293,In_1290);
xor U2318 (N_2318,In_3253,In_157);
nand U2319 (N_2319,In_4612,In_4272);
nand U2320 (N_2320,In_1860,In_2123);
xor U2321 (N_2321,In_3504,In_4901);
nor U2322 (N_2322,In_4674,In_3250);
nand U2323 (N_2323,In_4825,In_3195);
nor U2324 (N_2324,In_4234,In_2408);
and U2325 (N_2325,In_2857,In_394);
xnor U2326 (N_2326,In_308,In_4044);
nand U2327 (N_2327,In_4373,In_1213);
xnor U2328 (N_2328,In_4507,In_932);
nor U2329 (N_2329,In_626,In_1318);
xor U2330 (N_2330,In_4908,In_891);
or U2331 (N_2331,In_4089,In_1636);
xor U2332 (N_2332,In_3086,In_2501);
or U2333 (N_2333,In_10,In_969);
and U2334 (N_2334,In_1051,In_464);
nand U2335 (N_2335,In_4743,In_2240);
xor U2336 (N_2336,In_1248,In_2735);
and U2337 (N_2337,In_1773,In_4521);
or U2338 (N_2338,In_4519,In_3382);
xnor U2339 (N_2339,In_4586,In_1342);
nand U2340 (N_2340,In_3539,In_2122);
nand U2341 (N_2341,In_236,In_678);
nand U2342 (N_2342,In_1163,In_3280);
nor U2343 (N_2343,In_3914,In_4009);
xnor U2344 (N_2344,In_2525,In_2608);
xnor U2345 (N_2345,In_3777,In_921);
nand U2346 (N_2346,In_2769,In_648);
or U2347 (N_2347,In_66,In_4833);
nor U2348 (N_2348,In_4855,In_1179);
or U2349 (N_2349,In_1698,In_386);
and U2350 (N_2350,In_4014,In_1259);
nand U2351 (N_2351,In_1781,In_3956);
nand U2352 (N_2352,In_6,In_2569);
nand U2353 (N_2353,In_3203,In_4548);
nand U2354 (N_2354,In_1568,In_4596);
xnor U2355 (N_2355,In_1777,In_1361);
and U2356 (N_2356,In_3122,In_1365);
or U2357 (N_2357,In_3462,In_1306);
and U2358 (N_2358,In_2581,In_2947);
nand U2359 (N_2359,In_4594,In_944);
nor U2360 (N_2360,In_4064,In_4721);
nor U2361 (N_2361,In_4084,In_3984);
or U2362 (N_2362,In_3015,In_1799);
nand U2363 (N_2363,In_4372,In_3649);
nand U2364 (N_2364,In_2101,In_3024);
and U2365 (N_2365,In_3011,In_4518);
xor U2366 (N_2366,In_3215,In_1174);
xor U2367 (N_2367,In_2452,In_1896);
or U2368 (N_2368,In_4840,In_241);
nand U2369 (N_2369,In_179,In_735);
and U2370 (N_2370,In_1406,In_1945);
and U2371 (N_2371,In_235,In_4503);
xnor U2372 (N_2372,In_1742,In_1434);
or U2373 (N_2373,In_4321,In_3335);
nor U2374 (N_2374,In_1878,In_3179);
or U2375 (N_2375,In_1513,In_1941);
nor U2376 (N_2376,In_4041,In_1952);
or U2377 (N_2377,In_4985,In_4475);
nand U2378 (N_2378,In_3927,In_1261);
nor U2379 (N_2379,In_1382,In_2163);
or U2380 (N_2380,In_718,In_1730);
xnor U2381 (N_2381,In_618,In_2012);
or U2382 (N_2382,In_3635,In_2589);
nand U2383 (N_2383,In_2712,In_1989);
or U2384 (N_2384,In_4359,In_4755);
nor U2385 (N_2385,In_2939,In_4125);
nor U2386 (N_2386,In_2190,In_4106);
or U2387 (N_2387,In_3026,In_4226);
xor U2388 (N_2388,In_2019,In_2230);
xnor U2389 (N_2389,In_1795,In_2090);
or U2390 (N_2390,In_2991,In_2976);
or U2391 (N_2391,In_4986,In_1758);
or U2392 (N_2392,In_787,In_827);
nor U2393 (N_2393,In_2170,In_144);
xnor U2394 (N_2394,In_2880,In_2455);
xnor U2395 (N_2395,In_4172,In_559);
or U2396 (N_2396,In_3826,In_1578);
and U2397 (N_2397,In_2897,In_4665);
nand U2398 (N_2398,In_3816,In_1140);
nor U2399 (N_2399,In_45,In_110);
and U2400 (N_2400,In_4927,In_4778);
nor U2401 (N_2401,In_3753,In_3581);
xnor U2402 (N_2402,In_2872,In_4698);
nand U2403 (N_2403,In_868,In_1420);
and U2404 (N_2404,In_4425,In_610);
and U2405 (N_2405,In_28,In_4910);
and U2406 (N_2406,In_1244,In_1228);
xnor U2407 (N_2407,In_3290,In_225);
nand U2408 (N_2408,In_2374,In_3171);
and U2409 (N_2409,In_1413,In_2420);
or U2410 (N_2410,In_3626,In_4526);
xnor U2411 (N_2411,In_3005,In_2310);
xor U2412 (N_2412,In_4118,In_1697);
xor U2413 (N_2413,In_3566,In_3201);
or U2414 (N_2414,In_3111,In_1507);
and U2415 (N_2415,In_2143,In_3113);
nor U2416 (N_2416,In_2051,In_392);
and U2417 (N_2417,In_3328,In_360);
and U2418 (N_2418,In_2600,In_1884);
nor U2419 (N_2419,In_4513,In_278);
nor U2420 (N_2420,In_2972,In_4949);
and U2421 (N_2421,In_1721,In_1033);
or U2422 (N_2422,In_2055,In_4792);
nand U2423 (N_2423,In_429,In_4342);
nor U2424 (N_2424,In_2566,In_4589);
or U2425 (N_2425,In_2496,In_3285);
and U2426 (N_2426,In_228,In_382);
nor U2427 (N_2427,In_981,In_2761);
nor U2428 (N_2428,In_197,In_4070);
and U2429 (N_2429,In_3966,In_1393);
nor U2430 (N_2430,In_2937,In_3188);
and U2431 (N_2431,In_500,In_4238);
nor U2432 (N_2432,In_3838,In_1407);
nor U2433 (N_2433,In_3245,In_1841);
nand U2434 (N_2434,In_2798,In_4371);
nand U2435 (N_2435,In_1647,In_2979);
and U2436 (N_2436,In_1212,In_2744);
or U2437 (N_2437,In_1747,In_3997);
and U2438 (N_2438,In_663,In_3993);
xnor U2439 (N_2439,In_2865,In_2824);
nand U2440 (N_2440,In_3219,In_1172);
nand U2441 (N_2441,In_1451,In_1146);
nand U2442 (N_2442,In_347,In_2806);
nand U2443 (N_2443,In_3429,In_121);
and U2444 (N_2444,In_4189,In_2199);
nand U2445 (N_2445,In_2592,In_3590);
nand U2446 (N_2446,In_853,In_518);
nand U2447 (N_2447,In_403,In_3352);
nand U2448 (N_2448,In_260,In_2997);
nand U2449 (N_2449,In_2623,In_1897);
and U2450 (N_2450,In_855,In_3660);
or U2451 (N_2451,In_4061,In_1765);
nor U2452 (N_2452,In_4745,In_2273);
nand U2453 (N_2453,In_100,In_4054);
nand U2454 (N_2454,In_4375,In_2756);
or U2455 (N_2455,In_4944,In_4979);
or U2456 (N_2456,In_1794,In_3368);
xor U2457 (N_2457,In_596,In_4012);
nor U2458 (N_2458,In_1049,In_3330);
nand U2459 (N_2459,In_2468,In_85);
nor U2460 (N_2460,In_2376,In_3599);
and U2461 (N_2461,In_574,In_2518);
nor U2462 (N_2462,In_2278,In_4354);
and U2463 (N_2463,In_3452,In_1572);
and U2464 (N_2464,In_1430,In_4440);
nor U2465 (N_2465,In_4168,In_4194);
and U2466 (N_2466,In_3205,In_1283);
or U2467 (N_2467,In_4024,In_4871);
and U2468 (N_2468,In_2292,In_438);
nor U2469 (N_2469,In_4417,In_1161);
nand U2470 (N_2470,In_3337,In_2676);
nor U2471 (N_2471,In_2219,In_3104);
and U2472 (N_2472,In_3593,In_4621);
or U2473 (N_2473,In_462,In_576);
nor U2474 (N_2474,In_1082,In_3232);
or U2475 (N_2475,In_2922,In_4083);
nor U2476 (N_2476,In_4841,In_343);
or U2477 (N_2477,In_4357,In_4468);
xnor U2478 (N_2478,In_3594,In_672);
and U2479 (N_2479,In_2799,In_2234);
nor U2480 (N_2480,In_223,In_3724);
xor U2481 (N_2481,In_349,In_938);
xnor U2482 (N_2482,In_3727,In_4124);
and U2483 (N_2483,In_4720,In_1184);
nor U2484 (N_2484,In_4287,In_4890);
nand U2485 (N_2485,In_2955,In_587);
xor U2486 (N_2486,In_3083,In_27);
or U2487 (N_2487,In_1920,In_3732);
xnor U2488 (N_2488,In_2368,In_2458);
nor U2489 (N_2489,In_91,In_1633);
and U2490 (N_2490,In_291,In_2868);
xor U2491 (N_2491,In_2611,In_836);
nor U2492 (N_2492,In_4874,In_1707);
and U2493 (N_2493,In_2736,In_4318);
and U2494 (N_2494,In_9,In_4400);
nor U2495 (N_2495,In_1931,In_93);
xnor U2496 (N_2496,In_366,In_3373);
and U2497 (N_2497,In_1987,In_951);
or U2498 (N_2498,In_967,In_757);
and U2499 (N_2499,In_329,In_2899);
xor U2500 (N_2500,N_2382,N_1802);
xor U2501 (N_2501,N_1723,N_188);
xor U2502 (N_2502,N_405,N_472);
and U2503 (N_2503,N_559,N_365);
xor U2504 (N_2504,N_687,N_2373);
xnor U2505 (N_2505,N_266,N_691);
xor U2506 (N_2506,N_2459,N_1314);
nor U2507 (N_2507,N_320,N_1355);
nor U2508 (N_2508,N_1876,N_447);
and U2509 (N_2509,N_1700,N_429);
or U2510 (N_2510,N_974,N_1473);
nor U2511 (N_2511,N_428,N_1343);
or U2512 (N_2512,N_1116,N_1776);
xor U2513 (N_2513,N_1749,N_760);
or U2514 (N_2514,N_211,N_1046);
nor U2515 (N_2515,N_839,N_750);
nand U2516 (N_2516,N_1824,N_1169);
nor U2517 (N_2517,N_1195,N_1950);
nand U2518 (N_2518,N_1651,N_1159);
xnor U2519 (N_2519,N_1470,N_636);
nand U2520 (N_2520,N_1477,N_831);
nor U2521 (N_2521,N_1100,N_672);
or U2522 (N_2522,N_1007,N_1809);
nand U2523 (N_2523,N_2088,N_825);
xor U2524 (N_2524,N_761,N_1271);
nor U2525 (N_2525,N_1713,N_523);
or U2526 (N_2526,N_256,N_1660);
xor U2527 (N_2527,N_1581,N_1170);
xnor U2528 (N_2528,N_2159,N_413);
or U2529 (N_2529,N_1358,N_880);
xnor U2530 (N_2530,N_1381,N_2273);
nand U2531 (N_2531,N_240,N_1460);
nor U2532 (N_2532,N_925,N_637);
and U2533 (N_2533,N_1655,N_971);
nor U2534 (N_2534,N_2447,N_13);
nor U2535 (N_2535,N_205,N_1413);
and U2536 (N_2536,N_2328,N_2496);
nor U2537 (N_2537,N_2448,N_330);
nor U2538 (N_2538,N_276,N_1575);
or U2539 (N_2539,N_418,N_888);
nor U2540 (N_2540,N_953,N_2326);
nor U2541 (N_2541,N_2428,N_493);
and U2542 (N_2542,N_1508,N_2409);
nand U2543 (N_2543,N_1264,N_846);
and U2544 (N_2544,N_918,N_620);
xor U2545 (N_2545,N_1111,N_1792);
xnor U2546 (N_2546,N_286,N_1134);
and U2547 (N_2547,N_1813,N_1178);
nor U2548 (N_2548,N_2177,N_2263);
nor U2549 (N_2549,N_44,N_963);
and U2550 (N_2550,N_1738,N_867);
and U2551 (N_2551,N_1455,N_1610);
xnor U2552 (N_2552,N_98,N_2228);
nand U2553 (N_2553,N_967,N_1637);
xnor U2554 (N_2554,N_1871,N_1210);
nand U2555 (N_2555,N_160,N_1);
nor U2556 (N_2556,N_2345,N_424);
or U2557 (N_2557,N_690,N_46);
xnor U2558 (N_2558,N_311,N_1843);
nand U2559 (N_2559,N_545,N_2434);
and U2560 (N_2560,N_1616,N_1668);
xnor U2561 (N_2561,N_1596,N_1770);
nand U2562 (N_2562,N_673,N_2202);
nand U2563 (N_2563,N_2265,N_1020);
nand U2564 (N_2564,N_392,N_952);
nor U2565 (N_2565,N_1211,N_1274);
and U2566 (N_2566,N_986,N_1775);
or U2567 (N_2567,N_217,N_105);
xor U2568 (N_2568,N_2184,N_693);
nor U2569 (N_2569,N_1681,N_210);
nand U2570 (N_2570,N_170,N_1244);
nor U2571 (N_2571,N_1250,N_1374);
nor U2572 (N_2572,N_1853,N_201);
nor U2573 (N_2573,N_1694,N_1137);
or U2574 (N_2574,N_2309,N_546);
and U2575 (N_2575,N_536,N_2090);
nand U2576 (N_2576,N_1277,N_21);
nand U2577 (N_2577,N_2096,N_2091);
or U2578 (N_2578,N_1526,N_183);
and U2579 (N_2579,N_209,N_767);
and U2580 (N_2580,N_425,N_1024);
nor U2581 (N_2581,N_1621,N_1816);
nor U2582 (N_2582,N_602,N_1400);
nor U2583 (N_2583,N_1035,N_862);
nor U2584 (N_2584,N_2436,N_306);
xnor U2585 (N_2585,N_1688,N_2267);
nor U2586 (N_2586,N_1428,N_650);
and U2587 (N_2587,N_1014,N_2457);
nand U2588 (N_2588,N_1615,N_1942);
nand U2589 (N_2589,N_101,N_258);
and U2590 (N_2590,N_560,N_1851);
nor U2591 (N_2591,N_2283,N_384);
nor U2592 (N_2592,N_2187,N_1260);
and U2593 (N_2593,N_2498,N_1349);
and U2594 (N_2594,N_1612,N_1590);
xnor U2595 (N_2595,N_965,N_1377);
nor U2596 (N_2596,N_689,N_784);
nand U2597 (N_2597,N_937,N_208);
nor U2598 (N_2598,N_510,N_2218);
or U2599 (N_2599,N_2020,N_2418);
or U2600 (N_2600,N_1263,N_2161);
nand U2601 (N_2601,N_207,N_1897);
or U2602 (N_2602,N_2480,N_909);
nor U2603 (N_2603,N_2348,N_464);
nand U2604 (N_2604,N_2433,N_1893);
nand U2605 (N_2605,N_1439,N_193);
xnor U2606 (N_2606,N_165,N_1577);
xor U2607 (N_2607,N_487,N_1078);
or U2608 (N_2608,N_2139,N_2086);
or U2609 (N_2609,N_94,N_1513);
nand U2610 (N_2610,N_896,N_728);
and U2611 (N_2611,N_1790,N_337);
xnor U2612 (N_2612,N_334,N_914);
and U2613 (N_2613,N_1567,N_1835);
nand U2614 (N_2614,N_87,N_1762);
nor U2615 (N_2615,N_619,N_412);
xnor U2616 (N_2616,N_1782,N_2035);
and U2617 (N_2617,N_25,N_2341);
and U2618 (N_2618,N_865,N_1949);
xor U2619 (N_2619,N_549,N_1807);
nand U2620 (N_2620,N_1002,N_448);
and U2621 (N_2621,N_268,N_1429);
nor U2622 (N_2622,N_2259,N_528);
nand U2623 (N_2623,N_265,N_519);
nand U2624 (N_2624,N_1874,N_1784);
xnor U2625 (N_2625,N_289,N_1204);
nand U2626 (N_2626,N_1885,N_2232);
or U2627 (N_2627,N_1704,N_1487);
xor U2628 (N_2628,N_819,N_2122);
and U2629 (N_2629,N_2393,N_2287);
or U2630 (N_2630,N_647,N_195);
nor U2631 (N_2631,N_924,N_1080);
nor U2632 (N_2632,N_1026,N_1437);
xnor U2633 (N_2633,N_938,N_1001);
nand U2634 (N_2634,N_2493,N_45);
nor U2635 (N_2635,N_2237,N_247);
and U2636 (N_2636,N_768,N_2201);
nand U2637 (N_2637,N_227,N_1654);
and U2638 (N_2638,N_2340,N_216);
and U2639 (N_2639,N_90,N_1129);
xnor U2640 (N_2640,N_2484,N_1541);
nor U2641 (N_2641,N_14,N_2145);
or U2642 (N_2642,N_754,N_1452);
and U2643 (N_2643,N_494,N_2198);
xnor U2644 (N_2644,N_39,N_1417);
nand U2645 (N_2645,N_395,N_993);
nor U2646 (N_2646,N_212,N_1741);
nand U2647 (N_2647,N_1328,N_2281);
or U2648 (N_2648,N_1918,N_1372);
or U2649 (N_2649,N_485,N_747);
xor U2650 (N_2650,N_2467,N_1607);
nor U2651 (N_2651,N_1865,N_575);
xor U2652 (N_2652,N_2374,N_1225);
or U2653 (N_2653,N_81,N_854);
xnor U2654 (N_2654,N_1407,N_1861);
or U2655 (N_2655,N_1150,N_1863);
nor U2656 (N_2656,N_2238,N_2185);
nor U2657 (N_2657,N_177,N_1088);
nand U2658 (N_2658,N_15,N_1803);
or U2659 (N_2659,N_2193,N_1383);
nor U2660 (N_2660,N_692,N_206);
or U2661 (N_2661,N_855,N_53);
and U2662 (N_2662,N_1102,N_980);
and U2663 (N_2663,N_1650,N_1633);
xor U2664 (N_2664,N_1983,N_452);
or U2665 (N_2665,N_2044,N_73);
and U2666 (N_2666,N_1198,N_460);
xor U2667 (N_2667,N_1773,N_390);
or U2668 (N_2668,N_1933,N_934);
xnor U2669 (N_2669,N_280,N_1342);
and U2670 (N_2670,N_2065,N_1181);
or U2671 (N_2671,N_2495,N_1265);
or U2672 (N_2672,N_1889,N_1245);
xor U2673 (N_2673,N_368,N_1005);
or U2674 (N_2674,N_155,N_778);
xor U2675 (N_2675,N_2454,N_350);
or U2676 (N_2676,N_1719,N_1724);
nand U2677 (N_2677,N_1311,N_696);
or U2678 (N_2678,N_2427,N_1795);
xor U2679 (N_2679,N_645,N_2449);
nor U2680 (N_2680,N_1391,N_336);
nor U2681 (N_2681,N_853,N_2053);
and U2682 (N_2682,N_594,N_961);
and U2683 (N_2683,N_2379,N_592);
nor U2684 (N_2684,N_940,N_158);
xnor U2685 (N_2685,N_997,N_32);
nand U2686 (N_2686,N_1368,N_710);
nor U2687 (N_2687,N_878,N_1533);
or U2688 (N_2688,N_327,N_2258);
xnor U2689 (N_2689,N_623,N_490);
xor U2690 (N_2690,N_2231,N_1016);
nor U2691 (N_2691,N_125,N_1187);
xor U2692 (N_2692,N_251,N_462);
or U2693 (N_2693,N_1869,N_2017);
and U2694 (N_2694,N_2097,N_532);
nor U2695 (N_2695,N_495,N_716);
and U2696 (N_2696,N_1769,N_2112);
and U2697 (N_2697,N_1721,N_659);
xor U2698 (N_2698,N_8,N_176);
xor U2699 (N_2699,N_474,N_1891);
xor U2700 (N_2700,N_866,N_588);
xnor U2701 (N_2701,N_926,N_2026);
and U2702 (N_2702,N_2067,N_1435);
or U2703 (N_2703,N_1718,N_254);
or U2704 (N_2704,N_2197,N_34);
nor U2705 (N_2705,N_2012,N_300);
xor U2706 (N_2706,N_1309,N_426);
and U2707 (N_2707,N_1303,N_1284);
and U2708 (N_2708,N_2465,N_1173);
nand U2709 (N_2709,N_64,N_2170);
and U2710 (N_2710,N_62,N_634);
nand U2711 (N_2711,N_2421,N_391);
xnor U2712 (N_2712,N_1798,N_543);
or U2713 (N_2713,N_2420,N_2289);
nor U2714 (N_2714,N_982,N_168);
and U2715 (N_2715,N_2183,N_1067);
nor U2716 (N_2716,N_1631,N_1947);
nor U2717 (N_2717,N_1747,N_1494);
nand U2718 (N_2718,N_998,N_1378);
or U2719 (N_2719,N_2068,N_2299);
xnor U2720 (N_2720,N_790,N_2473);
nand U2721 (N_2721,N_1862,N_2370);
nand U2722 (N_2722,N_1249,N_369);
or U2723 (N_2723,N_2194,N_2356);
or U2724 (N_2724,N_1845,N_1711);
and U2725 (N_2725,N_1691,N_1850);
or U2726 (N_2726,N_1171,N_1604);
nand U2727 (N_2727,N_2288,N_496);
or U2728 (N_2728,N_38,N_1739);
or U2729 (N_2729,N_1043,N_2404);
nand U2730 (N_2730,N_1986,N_2414);
nand U2731 (N_2731,N_126,N_2352);
or U2732 (N_2732,N_1971,N_916);
and U2733 (N_2733,N_644,N_367);
nor U2734 (N_2734,N_2027,N_1566);
xor U2735 (N_2735,N_2431,N_145);
xor U2736 (N_2736,N_1337,N_1888);
nand U2737 (N_2737,N_427,N_869);
nor U2738 (N_2738,N_705,N_617);
or U2739 (N_2739,N_2349,N_1825);
nand U2740 (N_2740,N_80,N_1414);
nand U2741 (N_2741,N_497,N_756);
nand U2742 (N_2742,N_1628,N_553);
and U2743 (N_2743,N_2158,N_456);
or U2744 (N_2744,N_1786,N_2461);
nor U2745 (N_2745,N_128,N_2372);
nand U2746 (N_2746,N_957,N_2142);
nor U2747 (N_2747,N_291,N_2062);
and U2748 (N_2748,N_1517,N_1144);
and U2749 (N_2749,N_759,N_1138);
xor U2750 (N_2750,N_2134,N_59);
nor U2751 (N_2751,N_2257,N_2042);
and U2752 (N_2752,N_739,N_1695);
or U2753 (N_2753,N_135,N_197);
nor U2754 (N_2754,N_2430,N_2308);
or U2755 (N_2755,N_1670,N_58);
nand U2756 (N_2756,N_518,N_1488);
and U2757 (N_2757,N_455,N_33);
or U2758 (N_2758,N_252,N_2074);
nand U2759 (N_2759,N_410,N_131);
xor U2760 (N_2760,N_1332,N_1029);
xnor U2761 (N_2761,N_2305,N_93);
and U2762 (N_2762,N_1938,N_298);
and U2763 (N_2763,N_1287,N_380);
xnor U2764 (N_2764,N_1013,N_2019);
xnor U2765 (N_2765,N_983,N_586);
or U2766 (N_2766,N_148,N_364);
xnor U2767 (N_2767,N_1962,N_1838);
nor U2768 (N_2768,N_2103,N_1913);
xor U2769 (N_2769,N_1787,N_2350);
or U2770 (N_2770,N_1620,N_255);
and U2771 (N_2771,N_2261,N_2329);
nand U2772 (N_2772,N_565,N_738);
and U2773 (N_2773,N_2123,N_360);
xor U2774 (N_2774,N_1205,N_1267);
nand U2775 (N_2775,N_1890,N_1857);
xnor U2776 (N_2776,N_232,N_1237);
nor U2777 (N_2777,N_1426,N_1502);
xor U2778 (N_2778,N_723,N_2140);
or U2779 (N_2779,N_121,N_357);
xor U2780 (N_2780,N_12,N_627);
and U2781 (N_2781,N_1136,N_674);
nand U2782 (N_2782,N_1594,N_861);
nor U2783 (N_2783,N_2060,N_1406);
nand U2784 (N_2784,N_2082,N_292);
or U2785 (N_2785,N_318,N_1597);
and U2786 (N_2786,N_449,N_1228);
xor U2787 (N_2787,N_48,N_713);
nand U2788 (N_2788,N_1860,N_347);
nor U2789 (N_2789,N_1832,N_2162);
nor U2790 (N_2790,N_2113,N_1877);
and U2791 (N_2791,N_582,N_1980);
nor U2792 (N_2792,N_167,N_1906);
and U2793 (N_2793,N_649,N_304);
or U2794 (N_2794,N_844,N_1968);
and U2795 (N_2795,N_2176,N_1427);
xnor U2796 (N_2796,N_222,N_2336);
nor U2797 (N_2797,N_264,N_178);
nand U2798 (N_2798,N_1251,N_51);
xor U2799 (N_2799,N_1050,N_2233);
or U2800 (N_2800,N_871,N_1261);
and U2801 (N_2801,N_1586,N_1475);
nand U2802 (N_2802,N_224,N_230);
or U2803 (N_2803,N_1164,N_2313);
xnor U2804 (N_2804,N_1810,N_1659);
xor U2805 (N_2805,N_1232,N_781);
and U2806 (N_2806,N_801,N_1096);
and U2807 (N_2807,N_840,N_338);
nor U2808 (N_2808,N_1397,N_615);
nor U2809 (N_2809,N_1120,N_873);
or U2810 (N_2810,N_420,N_2410);
and U2811 (N_2811,N_1532,N_1565);
xor U2812 (N_2812,N_438,N_226);
nor U2813 (N_2813,N_1037,N_1822);
nor U2814 (N_2814,N_1834,N_1085);
nor U2815 (N_2815,N_2485,N_2392);
nand U2816 (N_2816,N_1320,N_1006);
xnor U2817 (N_2817,N_960,N_1990);
nand U2818 (N_2818,N_1965,N_1525);
nor U2819 (N_2819,N_1736,N_1305);
nor U2820 (N_2820,N_1151,N_590);
nand U2821 (N_2821,N_134,N_1730);
or U2822 (N_2822,N_421,N_1583);
nor U2823 (N_2823,N_1931,N_1767);
and U2824 (N_2824,N_1558,N_2018);
xor U2825 (N_2825,N_544,N_908);
and U2826 (N_2826,N_2051,N_803);
or U2827 (N_2827,N_301,N_2422);
nor U2828 (N_2828,N_2456,N_1732);
nand U2829 (N_2829,N_2400,N_1247);
nand U2830 (N_2830,N_881,N_2272);
and U2831 (N_2831,N_2056,N_1665);
nand U2832 (N_2832,N_1077,N_731);
and U2833 (N_2833,N_1573,N_706);
nor U2834 (N_2834,N_1471,N_1817);
nand U2835 (N_2835,N_221,N_1412);
or U2836 (N_2836,N_775,N_1568);
nand U2837 (N_2837,N_1093,N_2115);
nand U2838 (N_2838,N_1672,N_1466);
xor U2839 (N_2839,N_1369,N_1584);
nand U2840 (N_2840,N_2411,N_1595);
nand U2841 (N_2841,N_618,N_2151);
or U2842 (N_2842,N_915,N_54);
nor U2843 (N_2843,N_1048,N_1639);
or U2844 (N_2844,N_2247,N_837);
and U2845 (N_2845,N_2337,N_2174);
xor U2846 (N_2846,N_2081,N_1556);
nor U2847 (N_2847,N_535,N_707);
nor U2848 (N_2848,N_1549,N_2204);
nor U2849 (N_2849,N_797,N_807);
nor U2850 (N_2850,N_1319,N_595);
or U2851 (N_2851,N_1056,N_987);
nand U2852 (N_2852,N_2104,N_1168);
nor U2853 (N_2853,N_1800,N_1109);
xnor U2854 (N_2854,N_2355,N_599);
or U2855 (N_2855,N_1658,N_275);
and U2856 (N_2856,N_2052,N_505);
nor U2857 (N_2857,N_1622,N_2253);
and U2858 (N_2858,N_945,N_612);
xor U2859 (N_2859,N_753,N_736);
nand U2860 (N_2860,N_274,N_1047);
and U2861 (N_2861,N_1061,N_944);
and U2862 (N_2862,N_1486,N_1291);
nor U2863 (N_2863,N_1106,N_2450);
xor U2864 (N_2864,N_2029,N_529);
nand U2865 (N_2865,N_382,N_1161);
nor U2866 (N_2866,N_2451,N_1399);
and U2867 (N_2867,N_1018,N_151);
nor U2868 (N_2868,N_2458,N_2063);
nor U2869 (N_2869,N_583,N_715);
xor U2870 (N_2870,N_859,N_407);
or U2871 (N_2871,N_2129,N_2001);
or U2872 (N_2872,N_1602,N_2280);
and U2873 (N_2873,N_1587,N_1032);
or U2874 (N_2874,N_1632,N_669);
or U2875 (N_2875,N_1829,N_2083);
nand U2876 (N_2876,N_648,N_2266);
or U2877 (N_2877,N_1425,N_1553);
xnor U2878 (N_2878,N_563,N_1112);
or U2879 (N_2879,N_2284,N_1640);
nand U2880 (N_2880,N_2487,N_1742);
nand U2881 (N_2881,N_42,N_933);
xor U2882 (N_2882,N_851,N_2127);
xnor U2883 (N_2883,N_451,N_1939);
and U2884 (N_2884,N_1201,N_2069);
nor U2885 (N_2885,N_638,N_1347);
and U2886 (N_2886,N_555,N_657);
and U2887 (N_2887,N_776,N_1371);
nor U2888 (N_2888,N_2072,N_1031);
nand U2889 (N_2889,N_770,N_1952);
xnor U2890 (N_2890,N_872,N_484);
xor U2891 (N_2891,N_1392,N_1367);
and U2892 (N_2892,N_1300,N_444);
xnor U2893 (N_2893,N_959,N_1868);
and U2894 (N_2894,N_1076,N_1310);
or U2895 (N_2895,N_1192,N_2242);
xor U2896 (N_2896,N_370,N_1768);
nor U2897 (N_2897,N_2039,N_2107);
nand U2898 (N_2898,N_198,N_1126);
and U2899 (N_2899,N_1238,N_661);
nand U2900 (N_2900,N_717,N_1656);
and U2901 (N_2901,N_968,N_1131);
nor U2902 (N_2902,N_2130,N_522);
nand U2903 (N_2903,N_1440,N_1820);
nor U2904 (N_2904,N_1248,N_2028);
nand U2905 (N_2905,N_1197,N_2189);
nand U2906 (N_2906,N_1924,N_1463);
or U2907 (N_2907,N_43,N_2398);
and U2908 (N_2908,N_18,N_901);
nand U2909 (N_2909,N_2339,N_65);
and U2910 (N_2910,N_2312,N_1958);
and U2911 (N_2911,N_1752,N_1712);
xnor U2912 (N_2912,N_498,N_83);
or U2913 (N_2913,N_2375,N_132);
or U2914 (N_2914,N_406,N_2116);
or U2915 (N_2915,N_319,N_1348);
and U2916 (N_2916,N_1149,N_23);
xnor U2917 (N_2917,N_215,N_2364);
xor U2918 (N_2918,N_718,N_624);
nor U2919 (N_2919,N_2160,N_2150);
xor U2920 (N_2920,N_29,N_1548);
and U2921 (N_2921,N_1570,N_1403);
nand U2922 (N_2922,N_589,N_762);
and U2923 (N_2923,N_2025,N_2325);
and U2924 (N_2924,N_294,N_2225);
and U2925 (N_2925,N_450,N_1789);
and U2926 (N_2926,N_703,N_1432);
nor U2927 (N_2927,N_1456,N_1881);
and U2928 (N_2928,N_2285,N_1550);
nand U2929 (N_2929,N_999,N_1702);
nor U2930 (N_2930,N_780,N_1158);
xor U2931 (N_2931,N_1411,N_1256);
xor U2932 (N_2932,N_1922,N_681);
nand U2933 (N_2933,N_662,N_1282);
nor U2934 (N_2934,N_1199,N_1469);
or U2935 (N_2935,N_1344,N_157);
nand U2936 (N_2936,N_2076,N_295);
nand U2937 (N_2937,N_1734,N_1783);
and U2938 (N_2938,N_1837,N_1454);
xnor U2939 (N_2939,N_743,N_830);
nand U2940 (N_2940,N_966,N_469);
nand U2941 (N_2941,N_2327,N_1200);
xor U2942 (N_2942,N_1049,N_1230);
and U2943 (N_2943,N_566,N_895);
xnor U2944 (N_2944,N_114,N_515);
xor U2945 (N_2945,N_1357,N_1193);
and U2946 (N_2946,N_2108,N_1107);
and U2947 (N_2947,N_682,N_343);
nor U2948 (N_2948,N_379,N_142);
nand U2949 (N_2949,N_2383,N_2157);
nand U2950 (N_2950,N_1686,N_1777);
or U2951 (N_2951,N_1805,N_1993);
and U2952 (N_2952,N_698,N_1735);
nor U2953 (N_2953,N_2260,N_2306);
and U2954 (N_2954,N_2058,N_2221);
xnor U2955 (N_2955,N_1353,N_992);
or U2956 (N_2956,N_1313,N_223);
xnor U2957 (N_2957,N_1935,N_1053);
nor U2958 (N_2958,N_2008,N_1366);
nand U2959 (N_2959,N_607,N_1467);
nand U2960 (N_2960,N_2136,N_538);
or U2961 (N_2961,N_810,N_900);
xnor U2962 (N_2962,N_1509,N_626);
or U2963 (N_2963,N_2424,N_1917);
nand U2964 (N_2964,N_86,N_2262);
or U2965 (N_2965,N_1443,N_233);
nand U2966 (N_2966,N_1666,N_958);
and U2967 (N_2967,N_943,N_1104);
or U2968 (N_2968,N_939,N_1981);
and U2969 (N_2969,N_2222,N_1393);
nand U2970 (N_2970,N_1864,N_1852);
or U2971 (N_2971,N_1405,N_796);
and U2972 (N_2972,N_1506,N_1995);
xor U2973 (N_2973,N_414,N_1269);
nor U2974 (N_2974,N_2054,N_931);
nand U2975 (N_2975,N_2464,N_1543);
or U2976 (N_2976,N_2094,N_111);
nor U2977 (N_2977,N_1523,N_746);
and U2978 (N_2978,N_2439,N_501);
and U2979 (N_2979,N_2126,N_430);
xnor U2980 (N_2980,N_376,N_1716);
nor U2981 (N_2981,N_2316,N_622);
nor U2982 (N_2982,N_541,N_2200);
nand U2983 (N_2983,N_1040,N_61);
nand U2984 (N_2984,N_1304,N_153);
nand U2985 (N_2985,N_1335,N_1395);
and U2986 (N_2986,N_2073,N_2359);
or U2987 (N_2987,N_1177,N_1234);
nand U2988 (N_2988,N_2169,N_2011);
or U2989 (N_2989,N_667,N_1979);
or U2990 (N_2990,N_1207,N_1012);
nand U2991 (N_2991,N_1507,N_2138);
and U2992 (N_2992,N_817,N_1647);
nor U2993 (N_2993,N_2460,N_2417);
and U2994 (N_2994,N_1848,N_1840);
and U2995 (N_2995,N_1341,N_2210);
nor U2996 (N_2996,N_1290,N_400);
nor U2997 (N_2997,N_398,N_680);
xnor U2998 (N_2998,N_113,N_632);
nand U2999 (N_2999,N_2271,N_1683);
and U3000 (N_3000,N_729,N_678);
or U3001 (N_3001,N_323,N_603);
or U3002 (N_3002,N_1329,N_1415);
or U3003 (N_3003,N_506,N_990);
nor U3004 (N_3004,N_1272,N_1756);
or U3005 (N_3005,N_362,N_1294);
nand U3006 (N_3006,N_1438,N_100);
xnor U3007 (N_3007,N_187,N_1559);
and U3008 (N_3008,N_2371,N_1608);
nand U3009 (N_3009,N_601,N_2021);
and U3010 (N_3010,N_1521,N_1926);
and U3011 (N_3011,N_832,N_1472);
or U3012 (N_3012,N_655,N_863);
and U3013 (N_3013,N_2226,N_2438);
nand U3014 (N_3014,N_2037,N_2114);
nor U3015 (N_3015,N_1288,N_1243);
or U3016 (N_3016,N_112,N_2041);
nor U3017 (N_3017,N_598,N_1844);
nand U3018 (N_3018,N_639,N_2478);
nor U3019 (N_3019,N_2085,N_1614);
or U3020 (N_3020,N_2230,N_1125);
nand U3021 (N_3021,N_2207,N_246);
and U3022 (N_3022,N_1160,N_1360);
and U3023 (N_3023,N_1669,N_175);
and U3024 (N_3024,N_1582,N_277);
or U3025 (N_3025,N_771,N_1649);
xnor U3026 (N_3026,N_573,N_972);
or U3027 (N_3027,N_244,N_235);
nand U3028 (N_3028,N_184,N_66);
and U3029 (N_3029,N_2220,N_1791);
nand U3030 (N_3030,N_2124,N_2307);
nand U3031 (N_3031,N_630,N_1017);
xor U3032 (N_3032,N_1699,N_1912);
nand U3033 (N_3033,N_1387,N_795);
xor U3034 (N_3034,N_1379,N_2335);
nand U3035 (N_3035,N_1388,N_2203);
and U3036 (N_3036,N_2486,N_1424);
nand U3037 (N_3037,N_1492,N_1461);
and U3038 (N_3038,N_514,N_2396);
or U3039 (N_3039,N_1645,N_1957);
xnor U3040 (N_3040,N_1644,N_1330);
or U3041 (N_3041,N_699,N_733);
nand U3042 (N_3042,N_702,N_2215);
and U3043 (N_3043,N_1948,N_561);
nor U3044 (N_3044,N_1866,N_1833);
xor U3045 (N_3045,N_970,N_1626);
and U3046 (N_3046,N_1879,N_242);
xor U3047 (N_3047,N_847,N_1978);
nor U3048 (N_3048,N_1538,N_1398);
nor U3049 (N_3049,N_572,N_231);
and U3050 (N_3050,N_1765,N_2455);
and U3051 (N_3051,N_2049,N_1618);
nor U3052 (N_3052,N_203,N_1384);
nand U3053 (N_3053,N_1780,N_1110);
and U3054 (N_3054,N_278,N_1709);
and U3055 (N_3055,N_1396,N_1380);
and U3056 (N_3056,N_1592,N_902);
nor U3057 (N_3057,N_110,N_1153);
nand U3058 (N_3058,N_2282,N_2077);
xor U3059 (N_3059,N_419,N_82);
and U3060 (N_3060,N_471,N_1674);
xor U3061 (N_3061,N_371,N_826);
and U3062 (N_3062,N_2346,N_2223);
or U3063 (N_3063,N_580,N_1450);
xor U3064 (N_3064,N_1292,N_969);
xor U3065 (N_3065,N_989,N_179);
nand U3066 (N_3066,N_1841,N_2133);
xnor U3067 (N_3067,N_1015,N_1004);
xnor U3068 (N_3068,N_339,N_791);
and U3069 (N_3069,N_303,N_608);
nand U3070 (N_3070,N_1870,N_36);
nor U3071 (N_3071,N_660,N_1057);
or U3072 (N_3072,N_149,N_1814);
xnor U3073 (N_3073,N_503,N_633);
nand U3074 (N_3074,N_2293,N_454);
nor U3075 (N_3075,N_2038,N_1598);
and U3076 (N_3076,N_954,N_1190);
nand U3077 (N_3077,N_1629,N_1551);
nor U3078 (N_3078,N_1726,N_431);
xor U3079 (N_3079,N_950,N_467);
or U3080 (N_3080,N_1318,N_883);
and U3081 (N_3081,N_377,N_1821);
xnor U3082 (N_3082,N_1087,N_2239);
nor U3083 (N_3083,N_834,N_508);
and U3084 (N_3084,N_806,N_1748);
nor U3085 (N_3085,N_1194,N_857);
nor U3086 (N_3086,N_2241,N_2463);
or U3087 (N_3087,N_554,N_7);
nand U3088 (N_3088,N_2472,N_1707);
nand U3089 (N_3089,N_1994,N_287);
or U3090 (N_3090,N_1281,N_181);
nand U3091 (N_3091,N_978,N_1246);
and U3092 (N_3092,N_164,N_1321);
xnor U3093 (N_3093,N_1402,N_1206);
nor U3094 (N_3094,N_1060,N_375);
nand U3095 (N_3095,N_1054,N_1066);
xnor U3096 (N_3096,N_1905,N_2391);
nand U3097 (N_3097,N_1761,N_2055);
xnor U3098 (N_3098,N_2084,N_272);
and U3099 (N_3099,N_2442,N_913);
nand U3100 (N_3100,N_1720,N_587);
xnor U3101 (N_3101,N_2032,N_499);
xnor U3102 (N_3102,N_27,N_885);
nand U3103 (N_3103,N_2483,N_625);
nand U3104 (N_3104,N_2059,N_1630);
and U3105 (N_3105,N_481,N_1627);
and U3106 (N_3106,N_1166,N_1363);
nand U3107 (N_3107,N_2432,N_1090);
nand U3108 (N_3108,N_1359,N_1479);
nor U3109 (N_3109,N_1324,N_2407);
nor U3110 (N_3110,N_1385,N_1172);
or U3111 (N_3111,N_1685,N_1510);
xnor U3112 (N_3112,N_726,N_838);
nor U3113 (N_3113,N_2030,N_1836);
xor U3114 (N_3114,N_141,N_1514);
or U3115 (N_3115,N_1585,N_2435);
or U3116 (N_3116,N_1481,N_159);
and U3117 (N_3117,N_973,N_1985);
nand U3118 (N_3118,N_685,N_1336);
nand U3119 (N_3119,N_1572,N_1804);
or U3120 (N_3120,N_841,N_1216);
xor U3121 (N_3121,N_1420,N_2180);
or U3122 (N_3122,N_1401,N_1536);
or U3123 (N_3123,N_1914,N_76);
xnor U3124 (N_3124,N_26,N_1323);
nand U3125 (N_3125,N_1916,N_2499);
nand U3126 (N_3126,N_22,N_10);
xor U3127 (N_3127,N_457,N_1408);
and U3128 (N_3128,N_1953,N_2279);
nor U3129 (N_3129,N_2323,N_905);
and U3130 (N_3130,N_2022,N_1280);
or U3131 (N_3131,N_279,N_1934);
and U3132 (N_3132,N_1921,N_1223);
nand U3133 (N_3133,N_1867,N_1667);
nand U3134 (N_3134,N_1527,N_314);
and U3135 (N_3135,N_182,N_2154);
or U3136 (N_3136,N_1788,N_346);
xnor U3137 (N_3137,N_1710,N_1708);
or U3138 (N_3138,N_1972,N_1653);
or U3139 (N_3139,N_1316,N_1546);
nor U3140 (N_3140,N_1498,N_2212);
nor U3141 (N_3141,N_2118,N_635);
nand U3142 (N_3142,N_290,N_397);
and U3143 (N_3143,N_1588,N_2111);
nor U3144 (N_3144,N_892,N_1763);
nor U3145 (N_3145,N_2098,N_1932);
or U3146 (N_3146,N_2469,N_0);
xor U3147 (N_3147,N_1184,N_1799);
xor U3148 (N_3148,N_764,N_1697);
nand U3149 (N_3149,N_663,N_2095);
or U3150 (N_3150,N_297,N_1725);
and U3151 (N_3151,N_1603,N_440);
nor U3152 (N_3152,N_354,N_2368);
or U3153 (N_3153,N_248,N_1530);
nand U3154 (N_3154,N_1350,N_374);
and U3155 (N_3155,N_409,N_1143);
xor U3156 (N_3156,N_238,N_2331);
or U3157 (N_3157,N_1499,N_856);
xnor U3158 (N_3158,N_1998,N_1505);
or U3159 (N_3159,N_530,N_628);
or U3160 (N_3160,N_2064,N_2235);
or U3161 (N_3161,N_2099,N_788);
or U3162 (N_3162,N_237,N_793);
or U3163 (N_3163,N_2195,N_1208);
xor U3164 (N_3164,N_2321,N_394);
nand U3165 (N_3165,N_827,N_2132);
or U3166 (N_3166,N_1661,N_568);
xnor U3167 (N_3167,N_2402,N_1278);
and U3168 (N_3168,N_1312,N_1489);
nand U3169 (N_3169,N_363,N_898);
nor U3170 (N_3170,N_1196,N_1375);
xor U3171 (N_3171,N_1065,N_1089);
nand U3172 (N_3172,N_714,N_2490);
xor U3173 (N_3173,N_829,N_876);
or U3174 (N_3174,N_2466,N_1929);
nor U3175 (N_3175,N_2304,N_1646);
xnor U3176 (N_3176,N_1919,N_1000);
nor U3177 (N_3177,N_1528,N_2256);
nor U3178 (N_3178,N_1854,N_443);
nand U3179 (N_3179,N_366,N_2286);
xor U3180 (N_3180,N_2381,N_2013);
nor U3181 (N_3181,N_701,N_194);
and U3182 (N_3182,N_604,N_1019);
xnor U3183 (N_3183,N_166,N_2249);
xor U3184 (N_3184,N_828,N_2416);
nand U3185 (N_3185,N_2387,N_1235);
and U3186 (N_3186,N_1760,N_127);
nand U3187 (N_3187,N_2246,N_77);
or U3188 (N_3188,N_1547,N_1887);
and U3189 (N_3189,N_2093,N_404);
or U3190 (N_3190,N_1673,N_2143);
nor U3191 (N_3191,N_1976,N_677);
or U3192 (N_3192,N_842,N_932);
xnor U3193 (N_3193,N_326,N_2369);
nor U3194 (N_3194,N_2300,N_270);
and U3195 (N_3195,N_2191,N_2110);
nand U3196 (N_3196,N_875,N_2390);
or U3197 (N_3197,N_1678,N_889);
xnor U3198 (N_3198,N_1812,N_2405);
nand U3199 (N_3199,N_1447,N_1535);
nor U3200 (N_3200,N_136,N_1657);
nor U3201 (N_3201,N_1458,N_118);
or U3202 (N_3202,N_1944,N_1222);
nand U3203 (N_3203,N_2179,N_109);
xor U3204 (N_3204,N_137,N_2208);
or U3205 (N_3205,N_1283,N_2453);
xnor U3206 (N_3206,N_283,N_631);
nand U3207 (N_3207,N_1878,N_752);
nor U3208 (N_3208,N_1955,N_814);
nand U3209 (N_3209,N_185,N_2100);
nand U3210 (N_3210,N_1418,N_2292);
nor U3211 (N_3211,N_611,N_820);
nand U3212 (N_3212,N_1152,N_1345);
xnor U3213 (N_3213,N_1524,N_2276);
xor U3214 (N_3214,N_96,N_527);
xnor U3215 (N_3215,N_1097,N_1262);
xnor U3216 (N_3216,N_1842,N_964);
nor U3217 (N_3217,N_789,N_1186);
and U3218 (N_3218,N_1797,N_1930);
nand U3219 (N_3219,N_316,N_1818);
or U3220 (N_3220,N_904,N_422);
or U3221 (N_3221,N_2403,N_1448);
or U3222 (N_3222,N_1883,N_156);
or U3223 (N_3223,N_2164,N_245);
and U3224 (N_3224,N_24,N_2357);
or U3225 (N_3225,N_1082,N_16);
xor U3226 (N_3226,N_228,N_629);
nor U3227 (N_3227,N_1634,N_281);
nor U3228 (N_3228,N_2213,N_2188);
nor U3229 (N_3229,N_1593,N_122);
nor U3230 (N_3230,N_1623,N_191);
nand U3231 (N_3231,N_2057,N_2290);
nand U3232 (N_3232,N_2010,N_340);
nand U3233 (N_3233,N_858,N_725);
or U3234 (N_3234,N_1920,N_2317);
or U3235 (N_3235,N_1044,N_2007);
and U3236 (N_3236,N_666,N_2178);
or U3237 (N_3237,N_1296,N_1285);
nor U3238 (N_3238,N_309,N_1516);
nand U3239 (N_3239,N_1218,N_1010);
or U3240 (N_3240,N_2149,N_769);
or U3241 (N_3241,N_610,N_928);
or U3242 (N_3242,N_267,N_688);
or U3243 (N_3243,N_2014,N_1959);
nor U3244 (N_3244,N_605,N_2386);
or U3245 (N_3245,N_2089,N_1563);
and U3246 (N_3246,N_984,N_991);
nor U3247 (N_3247,N_1943,N_1600);
nand U3248 (N_3248,N_1531,N_1179);
or U3249 (N_3249,N_1449,N_2033);
xnor U3250 (N_3250,N_1182,N_1706);
and U3251 (N_3251,N_335,N_200);
nand U3252 (N_3252,N_2397,N_199);
xor U3253 (N_3253,N_897,N_1317);
nor U3254 (N_3254,N_2385,N_1520);
or U3255 (N_3255,N_437,N_1497);
xnor U3256 (N_3256,N_2445,N_1501);
nand U3257 (N_3257,N_910,N_1468);
or U3258 (N_3258,N_1055,N_1690);
and U3259 (N_3259,N_1365,N_1286);
or U3260 (N_3260,N_1858,N_652);
or U3261 (N_3261,N_124,N_1113);
xor U3262 (N_3262,N_1175,N_2399);
and U3263 (N_3263,N_174,N_1638);
or U3264 (N_3264,N_385,N_1241);
xor U3265 (N_3265,N_1275,N_1202);
nor U3266 (N_3266,N_1295,N_930);
or U3267 (N_3267,N_1431,N_315);
xor U3268 (N_3268,N_1880,N_571);
nand U3269 (N_3269,N_1167,N_2181);
nor U3270 (N_3270,N_2268,N_2471);
xor U3271 (N_3271,N_656,N_2347);
nor U3272 (N_3272,N_1778,N_683);
nor U3273 (N_3273,N_1519,N_2389);
xor U3274 (N_3274,N_2000,N_882);
or U3275 (N_3275,N_2318,N_730);
nor U3276 (N_3276,N_749,N_988);
xnor U3277 (N_3277,N_1457,N_1619);
and U3278 (N_3278,N_1951,N_2102);
or U3279 (N_3279,N_1534,N_1253);
xnor U3280 (N_3280,N_1676,N_2314);
nand U3281 (N_3281,N_792,N_1999);
nor U3282 (N_3282,N_31,N_172);
xor U3283 (N_3283,N_225,N_2024);
nand U3284 (N_3284,N_57,N_1609);
or U3285 (N_3285,N_2360,N_2141);
xor U3286 (N_3286,N_1483,N_28);
or U3287 (N_3287,N_737,N_351);
xnor U3288 (N_3288,N_1491,N_1064);
nor U3289 (N_3289,N_441,N_482);
or U3290 (N_3290,N_2234,N_1404);
nor U3291 (N_3291,N_609,N_1185);
nor U3292 (N_3292,N_679,N_1970);
and U3293 (N_3293,N_2437,N_1105);
or U3294 (N_3294,N_2109,N_324);
xnor U3295 (N_3295,N_1569,N_709);
nor U3296 (N_3296,N_884,N_2277);
nor U3297 (N_3297,N_860,N_823);
and U3298 (N_3298,N_2489,N_317);
nand U3299 (N_3299,N_2366,N_864);
nor U3300 (N_3300,N_1485,N_818);
xnor U3301 (N_3301,N_2196,N_1500);
or U3302 (N_3302,N_1240,N_517);
and U3303 (N_3303,N_2048,N_1662);
xor U3304 (N_3304,N_1872,N_1338);
and U3305 (N_3305,N_836,N_1909);
and U3306 (N_3306,N_1083,N_1028);
xnor U3307 (N_3307,N_92,N_654);
nand U3308 (N_3308,N_249,N_402);
and U3309 (N_3309,N_2137,N_552);
and U3310 (N_3310,N_719,N_79);
xnor U3311 (N_3311,N_1859,N_1680);
nor U3312 (N_3312,N_1465,N_435);
and U3313 (N_3313,N_2087,N_1898);
xor U3314 (N_3314,N_1785,N_55);
and U3315 (N_3315,N_919,N_2);
xnor U3316 (N_3316,N_1239,N_389);
and U3317 (N_3317,N_1522,N_1663);
nand U3318 (N_3318,N_651,N_332);
and U3319 (N_3319,N_2245,N_477);
nor U3320 (N_3320,N_1030,N_1462);
nor U3321 (N_3321,N_2482,N_218);
or U3322 (N_3322,N_2351,N_525);
and U3323 (N_3323,N_2075,N_2298);
and U3324 (N_3324,N_1960,N_1423);
and U3325 (N_3325,N_341,N_381);
or U3326 (N_3326,N_1781,N_1099);
xnor U3327 (N_3327,N_1301,N_107);
nand U3328 (N_3328,N_1062,N_946);
nand U3329 (N_3329,N_2443,N_824);
nand U3330 (N_3330,N_670,N_1315);
xor U3331 (N_3331,N_1356,N_1259);
nand U3332 (N_3332,N_1636,N_1793);
xor U3333 (N_3333,N_47,N_1503);
nor U3334 (N_3334,N_1504,N_1894);
or U3335 (N_3335,N_2080,N_550);
xnor U3336 (N_3336,N_584,N_640);
nand U3337 (N_3337,N_1599,N_2358);
or U3338 (N_3338,N_329,N_1370);
or U3339 (N_3339,N_1969,N_1904);
or U3340 (N_3340,N_2002,N_123);
or U3341 (N_3341,N_1459,N_1213);
or U3342 (N_3342,N_1334,N_1091);
nand U3343 (N_3343,N_154,N_1146);
or U3344 (N_3344,N_735,N_312);
and U3345 (N_3345,N_1148,N_2217);
nor U3346 (N_3346,N_1495,N_899);
or U3347 (N_3347,N_1557,N_516);
and U3348 (N_3348,N_2199,N_616);
nor U3349 (N_3349,N_539,N_1191);
or U3350 (N_3350,N_1611,N_483);
and U3351 (N_3351,N_56,N_296);
nor U3352 (N_3352,N_773,N_1717);
nand U3353 (N_3353,N_1941,N_1911);
or U3354 (N_3354,N_1846,N_2380);
or U3355 (N_3355,N_711,N_985);
nor U3356 (N_3356,N_1826,N_1892);
and U3357 (N_3357,N_173,N_1340);
and U3358 (N_3358,N_1529,N_1737);
nand U3359 (N_3359,N_63,N_1220);
or U3360 (N_3360,N_84,N_1692);
nor U3361 (N_3361,N_542,N_261);
and U3362 (N_3362,N_877,N_2023);
xor U3363 (N_3363,N_2378,N_313);
or U3364 (N_3364,N_2440,N_1434);
and U3365 (N_3365,N_1578,N_812);
nand U3366 (N_3366,N_1308,N_1490);
nor U3367 (N_3367,N_772,N_2406);
and U3368 (N_3368,N_2423,N_2121);
or U3369 (N_3369,N_1176,N_2163);
nand U3370 (N_3370,N_1991,N_642);
and U3371 (N_3371,N_204,N_1464);
or U3372 (N_3372,N_2408,N_1731);
or U3373 (N_3373,N_1759,N_2206);
or U3374 (N_3374,N_2236,N_1693);
or U3375 (N_3375,N_2315,N_1022);
xnor U3376 (N_3376,N_1772,N_906);
nand U3377 (N_3377,N_1988,N_911);
nand U3378 (N_3378,N_331,N_234);
nor U3379 (N_3379,N_220,N_2168);
and U3380 (N_3380,N_1242,N_887);
or U3381 (N_3381,N_1419,N_41);
xor U3382 (N_3382,N_352,N_2243);
xor U3383 (N_3383,N_432,N_551);
and U3384 (N_3384,N_947,N_2446);
or U3385 (N_3385,N_740,N_1188);
xor U3386 (N_3386,N_1174,N_1127);
nor U3387 (N_3387,N_17,N_446);
and U3388 (N_3388,N_434,N_1696);
nand U3389 (N_3389,N_138,N_1794);
or U3390 (N_3390,N_1069,N_108);
nor U3391 (N_3391,N_1189,N_1900);
xnor U3392 (N_3392,N_786,N_2192);
nand U3393 (N_3393,N_463,N_171);
nor U3394 (N_3394,N_815,N_102);
xnor U3395 (N_3395,N_2252,N_2342);
or U3396 (N_3396,N_1299,N_2240);
xnor U3397 (N_3397,N_613,N_1364);
nor U3398 (N_3398,N_1122,N_1394);
nor U3399 (N_3399,N_567,N_461);
or U3400 (N_3400,N_163,N_1937);
or U3401 (N_3401,N_1236,N_1997);
nand U3402 (N_3402,N_2003,N_358);
xnor U3403 (N_3403,N_2319,N_1945);
or U3404 (N_3404,N_783,N_700);
and U3405 (N_3405,N_2148,N_1333);
and U3406 (N_3406,N_2412,N_2415);
or U3407 (N_3407,N_1624,N_1808);
xor U3408 (N_3408,N_1297,N_843);
nand U3409 (N_3409,N_2452,N_569);
and U3410 (N_3410,N_1307,N_2106);
and U3411 (N_3411,N_1936,N_2152);
or U3412 (N_3412,N_1442,N_1118);
xor U3413 (N_3413,N_2146,N_2264);
xnor U3414 (N_3414,N_196,N_229);
or U3415 (N_3415,N_2050,N_1745);
and U3416 (N_3416,N_475,N_282);
nor U3417 (N_3417,N_1270,N_1875);
or U3418 (N_3418,N_724,N_1928);
nand U3419 (N_3419,N_2441,N_1361);
nor U3420 (N_3420,N_1907,N_401);
or U3421 (N_3421,N_1051,N_799);
or U3422 (N_3422,N_1042,N_500);
nor U3423 (N_3423,N_470,N_1386);
nor U3424 (N_3424,N_1766,N_507);
nand U3425 (N_3425,N_1641,N_579);
or U3426 (N_3426,N_1555,N_879);
or U3427 (N_3427,N_1966,N_1101);
or U3428 (N_3428,N_2334,N_1758);
xnor U3429 (N_3429,N_2310,N_1084);
xnor U3430 (N_3430,N_2250,N_981);
and U3431 (N_3431,N_2036,N_1542);
xor U3432 (N_3432,N_1480,N_1902);
nor U3433 (N_3433,N_1512,N_2333);
nand U3434 (N_3434,N_1072,N_2477);
and U3435 (N_3435,N_116,N_403);
or U3436 (N_3436,N_593,N_1698);
or U3437 (N_3437,N_1989,N_2005);
nor U3438 (N_3438,N_1157,N_2302);
nor U3439 (N_3439,N_2070,N_1705);
xor U3440 (N_3440,N_1279,N_2474);
nor U3441 (N_3441,N_328,N_935);
nand U3442 (N_3442,N_373,N_1648);
nand U3443 (N_3443,N_540,N_1819);
xnor U3444 (N_3444,N_956,N_845);
xor U3445 (N_3445,N_712,N_2303);
nor U3446 (N_3446,N_1045,N_1849);
xor U3447 (N_3447,N_996,N_1940);
nor U3448 (N_3448,N_1923,N_433);
nand U3449 (N_3449,N_1254,N_537);
or U3450 (N_3450,N_1038,N_513);
or U3451 (N_3451,N_721,N_907);
xnor U3452 (N_3452,N_299,N_359);
nand U3453 (N_3453,N_75,N_2047);
nand U3454 (N_3454,N_445,N_1613);
nand U3455 (N_3455,N_40,N_798);
nand U3456 (N_3456,N_288,N_1119);
and U3457 (N_3457,N_1021,N_765);
nor U3458 (N_3458,N_597,N_162);
and U3459 (N_3459,N_2425,N_72);
nand U3460 (N_3460,N_1139,N_262);
xnor U3461 (N_3461,N_106,N_1132);
or U3462 (N_3462,N_1422,N_1373);
nor U3463 (N_3463,N_621,N_727);
nor U3464 (N_3464,N_694,N_2479);
xor U3465 (N_3465,N_704,N_833);
nand U3466 (N_3466,N_1231,N_606);
or U3467 (N_3467,N_2255,N_751);
and U3468 (N_3468,N_941,N_2294);
or U3469 (N_3469,N_1293,N_2344);
nand U3470 (N_3470,N_744,N_2488);
xnor U3471 (N_3471,N_2016,N_1352);
xor U3472 (N_3472,N_97,N_2429);
or U3473 (N_3473,N_653,N_1095);
and U3474 (N_3474,N_1011,N_800);
and U3475 (N_3475,N_2491,N_1895);
and U3476 (N_3476,N_1727,N_2361);
nand U3477 (N_3477,N_2395,N_1801);
xor U3478 (N_3478,N_473,N_2254);
or U3479 (N_3479,N_2167,N_129);
nor U3480 (N_3480,N_1103,N_822);
and U3481 (N_3481,N_994,N_1576);
and U3482 (N_3482,N_2105,N_491);
nor U3483 (N_3483,N_675,N_805);
nand U3484 (N_3484,N_2043,N_1071);
and U3485 (N_3485,N_949,N_891);
nor U3486 (N_3486,N_2354,N_1003);
nand U3487 (N_3487,N_2278,N_720);
nand U3488 (N_3488,N_777,N_1714);
xor U3489 (N_3489,N_2468,N_2071);
nor U3490 (N_3490,N_52,N_293);
and U3491 (N_3491,N_1561,N_1436);
nand U3492 (N_3492,N_4,N_259);
nor U3493 (N_3493,N_1073,N_349);
nor U3494 (N_3494,N_236,N_250);
and U3495 (N_3495,N_11,N_1823);
nor U3496 (N_3496,N_1684,N_2426);
or U3497 (N_3497,N_1474,N_2497);
nor U3498 (N_3498,N_202,N_557);
or U3499 (N_3499,N_779,N_758);
xor U3500 (N_3500,N_570,N_868);
xnor U3501 (N_3501,N_49,N_2009);
xnor U3502 (N_3502,N_436,N_1899);
nor U3503 (N_3503,N_2462,N_1975);
and U3504 (N_3504,N_578,N_91);
or U3505 (N_3505,N_2125,N_886);
nand U3506 (N_3506,N_50,N_1910);
or U3507 (N_3507,N_192,N_802);
nor U3508 (N_3508,N_948,N_2384);
and U3509 (N_3509,N_1430,N_1226);
or U3510 (N_3510,N_849,N_1155);
xnor U3511 (N_3511,N_835,N_585);
nand U3512 (N_3512,N_591,N_120);
or U3513 (N_3513,N_89,N_74);
nand U3514 (N_3514,N_686,N_923);
nor U3515 (N_3515,N_2131,N_1729);
nand U3516 (N_3516,N_466,N_1740);
and U3517 (N_3517,N_1771,N_1268);
nand U3518 (N_3518,N_1142,N_1075);
and U3519 (N_3519,N_1537,N_2353);
xor U3520 (N_3520,N_975,N_1289);
nor U3521 (N_3521,N_977,N_492);
and U3522 (N_3522,N_1896,N_2153);
nand U3523 (N_3523,N_665,N_104);
nor U3524 (N_3524,N_2274,N_1255);
or U3525 (N_3525,N_504,N_1233);
xor U3526 (N_3526,N_356,N_1227);
and U3527 (N_3527,N_912,N_19);
or U3528 (N_3528,N_348,N_2295);
nor U3529 (N_3529,N_1229,N_920);
nor U3530 (N_3530,N_671,N_556);
nand U3531 (N_3531,N_852,N_774);
xor U3532 (N_3532,N_2297,N_1257);
nor U3533 (N_3533,N_1036,N_1518);
nand U3534 (N_3534,N_1266,N_423);
xor U3535 (N_3535,N_1302,N_1108);
xor U3536 (N_3536,N_2171,N_2046);
or U3537 (N_3537,N_1703,N_1114);
or U3538 (N_3538,N_416,N_321);
xnor U3539 (N_3539,N_88,N_2166);
xnor U3540 (N_3540,N_1544,N_2120);
xor U3541 (N_3541,N_1165,N_458);
nand U3542 (N_3542,N_1963,N_78);
nand U3543 (N_3543,N_2079,N_2248);
or U3544 (N_3544,N_1416,N_1130);
and U3545 (N_3545,N_305,N_468);
xor U3546 (N_3546,N_870,N_2388);
xnor U3547 (N_3547,N_1306,N_1446);
or U3548 (N_3548,N_787,N_2244);
or U3549 (N_3549,N_378,N_2061);
nand U3550 (N_3550,N_1643,N_763);
or U3551 (N_3551,N_1733,N_658);
xnor U3552 (N_3552,N_186,N_2211);
xnor U3553 (N_3553,N_676,N_60);
and U3554 (N_3554,N_600,N_1679);
nor U3555 (N_3555,N_486,N_1540);
and U3556 (N_3556,N_1224,N_929);
and U3557 (N_3557,N_2006,N_372);
nand U3558 (N_3558,N_1092,N_1410);
and U3559 (N_3559,N_1390,N_1973);
xor U3560 (N_3560,N_558,N_2135);
or U3561 (N_3561,N_307,N_804);
nand U3562 (N_3562,N_995,N_2144);
nand U3563 (N_3563,N_1856,N_1074);
or U3564 (N_3564,N_146,N_6);
nand U3565 (N_3565,N_808,N_386);
nor U3566 (N_3566,N_521,N_1562);
nor U3567 (N_3567,N_894,N_344);
nor U3568 (N_3568,N_614,N_1276);
or U3569 (N_3569,N_2338,N_189);
or U3570 (N_3570,N_1560,N_1855);
nor U3571 (N_3571,N_417,N_2362);
nor U3572 (N_3572,N_1484,N_1008);
or U3573 (N_3573,N_263,N_1162);
nand U3574 (N_3574,N_564,N_2296);
xor U3575 (N_3575,N_1133,N_512);
or U3576 (N_3576,N_2275,N_1221);
nand U3577 (N_3577,N_1984,N_1755);
nand U3578 (N_3578,N_2494,N_180);
and U3579 (N_3579,N_1389,N_1815);
nor U3580 (N_3580,N_271,N_708);
xor U3581 (N_3581,N_962,N_213);
nand U3582 (N_3582,N_2147,N_1605);
or U3583 (N_3583,N_1954,N_1215);
and U3584 (N_3584,N_1039,N_30);
nor U3585 (N_3585,N_1154,N_596);
and U3586 (N_3586,N_388,N_1750);
or U3587 (N_3587,N_1034,N_1180);
xor U3588 (N_3588,N_1496,N_643);
xnor U3589 (N_3589,N_664,N_1376);
and U3590 (N_3590,N_2269,N_3);
xnor U3591 (N_3591,N_2190,N_757);
or U3592 (N_3592,N_1574,N_741);
or U3593 (N_3593,N_2045,N_745);
xor U3594 (N_3594,N_1140,N_1033);
or U3595 (N_3595,N_1183,N_2031);
xnor U3596 (N_3596,N_2101,N_1147);
nor U3597 (N_3597,N_2119,N_342);
xor U3598 (N_3598,N_1325,N_1258);
xor U3599 (N_3599,N_1493,N_67);
nor U3600 (N_3600,N_755,N_476);
and U3601 (N_3601,N_2330,N_2481);
xnor U3602 (N_3602,N_1982,N_85);
xor U3603 (N_3603,N_1086,N_697);
and U3604 (N_3604,N_35,N_1552);
nor U3605 (N_3605,N_1675,N_1121);
xor U3606 (N_3606,N_465,N_821);
and U3607 (N_3607,N_874,N_2172);
nand U3608 (N_3608,N_562,N_922);
nand U3609 (N_3609,N_442,N_1946);
or U3610 (N_3610,N_1617,N_1124);
and U3611 (N_3611,N_2175,N_816);
xor U3612 (N_3612,N_1796,N_2186);
and U3613 (N_3613,N_2078,N_748);
xor U3614 (N_3614,N_241,N_1830);
xor U3615 (N_3615,N_2332,N_214);
or U3616 (N_3616,N_1212,N_5);
nand U3617 (N_3617,N_1539,N_453);
nor U3618 (N_3618,N_273,N_1476);
or U3619 (N_3619,N_1421,N_2401);
xor U3620 (N_3620,N_1362,N_285);
and U3621 (N_3621,N_2034,N_130);
or U3622 (N_3622,N_1094,N_68);
nor U3623 (N_3623,N_143,N_2128);
and U3624 (N_3624,N_1041,N_480);
nor U3625 (N_3625,N_1515,N_1956);
nor U3626 (N_3626,N_150,N_2419);
or U3627 (N_3627,N_1839,N_2219);
nor U3628 (N_3628,N_2040,N_2476);
xnor U3629 (N_3629,N_581,N_1063);
and U3630 (N_3630,N_1882,N_520);
nor U3631 (N_3631,N_1764,N_1652);
and U3632 (N_3632,N_411,N_383);
nor U3633 (N_3633,N_1903,N_646);
xor U3634 (N_3634,N_1482,N_2301);
nor U3635 (N_3635,N_1806,N_782);
or U3636 (N_3636,N_794,N_139);
or U3637 (N_3637,N_2209,N_2322);
xnor U3638 (N_3638,N_1682,N_239);
or U3639 (N_3639,N_1564,N_1642);
and U3640 (N_3640,N_103,N_1884);
nand U3641 (N_3641,N_361,N_1135);
nor U3642 (N_3642,N_399,N_117);
xnor U3643 (N_3643,N_531,N_2363);
and U3644 (N_3644,N_478,N_893);
nand U3645 (N_3645,N_1701,N_1511);
and U3646 (N_3646,N_684,N_1441);
and U3647 (N_3647,N_1117,N_2270);
nand U3648 (N_3648,N_576,N_526);
or U3649 (N_3649,N_408,N_890);
xnor U3650 (N_3650,N_1252,N_2444);
or U3651 (N_3651,N_1580,N_95);
or U3652 (N_3652,N_1331,N_2475);
and U3653 (N_3653,N_459,N_2320);
and U3654 (N_3654,N_2155,N_734);
nand U3655 (N_3655,N_2413,N_936);
or U3656 (N_3656,N_1757,N_811);
and U3657 (N_3657,N_1098,N_548);
nand U3658 (N_3658,N_2224,N_1992);
or U3659 (N_3659,N_1589,N_1451);
nand U3660 (N_3660,N_1987,N_161);
nand U3661 (N_3661,N_533,N_2394);
nor U3662 (N_3662,N_1751,N_1339);
nand U3663 (N_3663,N_439,N_190);
or U3664 (N_3664,N_509,N_20);
or U3665 (N_3665,N_2324,N_1115);
and U3666 (N_3666,N_1908,N_813);
and U3667 (N_3667,N_1025,N_1915);
or U3668 (N_3668,N_1977,N_1925);
and U3669 (N_3669,N_2343,N_1744);
xnor U3670 (N_3670,N_1996,N_942);
and U3671 (N_3671,N_850,N_345);
xnor U3672 (N_3672,N_260,N_1409);
xor U3673 (N_3673,N_133,N_976);
or U3674 (N_3674,N_1831,N_2173);
nor U3675 (N_3675,N_119,N_695);
and U3676 (N_3676,N_1163,N_479);
or U3677 (N_3677,N_1591,N_1774);
xnor U3678 (N_3678,N_1974,N_1058);
and U3679 (N_3679,N_903,N_1059);
xnor U3680 (N_3680,N_1219,N_1722);
nor U3681 (N_3681,N_1811,N_766);
nor U3682 (N_3682,N_848,N_284);
or U3683 (N_3683,N_574,N_152);
xnor U3684 (N_3684,N_547,N_2214);
and U3685 (N_3685,N_2066,N_732);
nand U3686 (N_3686,N_502,N_2156);
and U3687 (N_3687,N_1689,N_921);
and U3688 (N_3688,N_2311,N_668);
or U3689 (N_3689,N_1827,N_1664);
nor U3690 (N_3690,N_1753,N_809);
or U3691 (N_3691,N_1728,N_722);
or U3692 (N_3692,N_1445,N_2229);
nor U3693 (N_3693,N_1298,N_1023);
and U3694 (N_3694,N_1635,N_2165);
xor U3695 (N_3695,N_415,N_387);
or U3696 (N_3696,N_1886,N_1779);
xnor U3697 (N_3697,N_1606,N_1351);
nand U3698 (N_3698,N_1052,N_2205);
or U3699 (N_3699,N_144,N_2492);
nor U3700 (N_3700,N_534,N_1847);
xnor U3701 (N_3701,N_1901,N_927);
xor U3702 (N_3702,N_489,N_1671);
nor U3703 (N_3703,N_1964,N_269);
xor U3704 (N_3704,N_577,N_1123);
xnor U3705 (N_3705,N_955,N_71);
nor U3706 (N_3706,N_1128,N_524);
nor U3707 (N_3707,N_1273,N_1079);
nand U3708 (N_3708,N_2227,N_1382);
and U3709 (N_3709,N_99,N_2470);
nand U3710 (N_3710,N_333,N_2365);
and U3711 (N_3711,N_2251,N_2182);
or U3712 (N_3712,N_1141,N_70);
or U3713 (N_3713,N_9,N_1873);
or U3714 (N_3714,N_785,N_169);
or U3715 (N_3715,N_2367,N_302);
xor U3716 (N_3716,N_396,N_1677);
nor U3717 (N_3717,N_69,N_2004);
nand U3718 (N_3718,N_488,N_1326);
nor U3719 (N_3719,N_1217,N_1209);
xor U3720 (N_3720,N_353,N_1214);
nand U3721 (N_3721,N_511,N_308);
nor U3722 (N_3722,N_951,N_2291);
or U3723 (N_3723,N_979,N_1009);
nand U3724 (N_3724,N_243,N_1156);
nand U3725 (N_3725,N_1327,N_1828);
nor U3726 (N_3726,N_1743,N_147);
nor U3727 (N_3727,N_1081,N_1070);
nor U3728 (N_3728,N_742,N_1478);
xor U3729 (N_3729,N_1927,N_140);
or U3730 (N_3730,N_1687,N_1625);
xnor U3731 (N_3731,N_1433,N_1967);
and U3732 (N_3732,N_1444,N_1145);
nand U3733 (N_3733,N_37,N_1961);
nand U3734 (N_3734,N_1068,N_2216);
and U3735 (N_3735,N_1754,N_1027);
xnor U3736 (N_3736,N_253,N_1715);
or U3737 (N_3737,N_115,N_1545);
nor U3738 (N_3738,N_917,N_641);
xnor U3739 (N_3739,N_2376,N_322);
xnor U3740 (N_3740,N_2377,N_1322);
and U3741 (N_3741,N_1554,N_2092);
and U3742 (N_3742,N_219,N_393);
or U3743 (N_3743,N_1571,N_325);
or U3744 (N_3744,N_310,N_1354);
and U3745 (N_3745,N_1203,N_1579);
and U3746 (N_3746,N_1346,N_1453);
xnor U3747 (N_3747,N_2117,N_257);
and U3748 (N_3748,N_2015,N_1601);
xnor U3749 (N_3749,N_355,N_1746);
nor U3750 (N_3750,N_924,N_2134);
or U3751 (N_3751,N_369,N_1497);
xor U3752 (N_3752,N_2151,N_1406);
xnor U3753 (N_3753,N_336,N_609);
and U3754 (N_3754,N_1780,N_1212);
xor U3755 (N_3755,N_365,N_709);
or U3756 (N_3756,N_1662,N_1313);
or U3757 (N_3757,N_2038,N_575);
and U3758 (N_3758,N_522,N_385);
xnor U3759 (N_3759,N_1248,N_2100);
xnor U3760 (N_3760,N_2150,N_857);
nand U3761 (N_3761,N_1335,N_1759);
nor U3762 (N_3762,N_1650,N_2136);
and U3763 (N_3763,N_1213,N_1456);
xor U3764 (N_3764,N_30,N_634);
nand U3765 (N_3765,N_378,N_1953);
or U3766 (N_3766,N_472,N_642);
and U3767 (N_3767,N_2039,N_2232);
xnor U3768 (N_3768,N_1399,N_1836);
nand U3769 (N_3769,N_1432,N_1470);
nor U3770 (N_3770,N_287,N_679);
or U3771 (N_3771,N_1047,N_440);
nand U3772 (N_3772,N_756,N_2037);
xor U3773 (N_3773,N_1819,N_620);
nand U3774 (N_3774,N_2226,N_966);
or U3775 (N_3775,N_121,N_389);
nand U3776 (N_3776,N_2489,N_2116);
or U3777 (N_3777,N_341,N_210);
nor U3778 (N_3778,N_1214,N_1296);
and U3779 (N_3779,N_987,N_324);
or U3780 (N_3780,N_2367,N_938);
nor U3781 (N_3781,N_909,N_195);
and U3782 (N_3782,N_1671,N_2034);
nor U3783 (N_3783,N_325,N_2209);
nor U3784 (N_3784,N_1455,N_2140);
and U3785 (N_3785,N_2391,N_1645);
and U3786 (N_3786,N_962,N_2222);
xnor U3787 (N_3787,N_374,N_2051);
nand U3788 (N_3788,N_1278,N_934);
nand U3789 (N_3789,N_1768,N_1866);
nand U3790 (N_3790,N_1560,N_2490);
xnor U3791 (N_3791,N_1442,N_64);
nand U3792 (N_3792,N_1727,N_856);
nand U3793 (N_3793,N_651,N_972);
xor U3794 (N_3794,N_1039,N_1375);
nand U3795 (N_3795,N_2213,N_1418);
and U3796 (N_3796,N_1173,N_2351);
nor U3797 (N_3797,N_1825,N_1100);
xnor U3798 (N_3798,N_1297,N_821);
and U3799 (N_3799,N_557,N_490);
and U3800 (N_3800,N_1976,N_1525);
nand U3801 (N_3801,N_1017,N_2249);
or U3802 (N_3802,N_1849,N_515);
or U3803 (N_3803,N_598,N_2358);
xor U3804 (N_3804,N_1605,N_645);
and U3805 (N_3805,N_1113,N_1074);
nand U3806 (N_3806,N_371,N_250);
and U3807 (N_3807,N_1078,N_2438);
or U3808 (N_3808,N_1885,N_1270);
or U3809 (N_3809,N_262,N_388);
and U3810 (N_3810,N_1656,N_1786);
or U3811 (N_3811,N_1356,N_2031);
xnor U3812 (N_3812,N_1713,N_2349);
nor U3813 (N_3813,N_690,N_884);
xor U3814 (N_3814,N_2200,N_113);
or U3815 (N_3815,N_1333,N_1604);
or U3816 (N_3816,N_400,N_1417);
nand U3817 (N_3817,N_732,N_579);
and U3818 (N_3818,N_539,N_2342);
or U3819 (N_3819,N_1518,N_2103);
xnor U3820 (N_3820,N_805,N_1030);
xor U3821 (N_3821,N_2314,N_2153);
or U3822 (N_3822,N_1063,N_2409);
and U3823 (N_3823,N_1133,N_1750);
nand U3824 (N_3824,N_1648,N_31);
nand U3825 (N_3825,N_2406,N_1898);
nor U3826 (N_3826,N_1680,N_1671);
or U3827 (N_3827,N_1269,N_652);
and U3828 (N_3828,N_738,N_1286);
and U3829 (N_3829,N_1534,N_2484);
xnor U3830 (N_3830,N_494,N_1552);
xnor U3831 (N_3831,N_120,N_1299);
xor U3832 (N_3832,N_60,N_1740);
nor U3833 (N_3833,N_903,N_1328);
xor U3834 (N_3834,N_1311,N_1469);
xnor U3835 (N_3835,N_1723,N_1329);
xor U3836 (N_3836,N_1815,N_1949);
and U3837 (N_3837,N_1904,N_44);
nor U3838 (N_3838,N_1985,N_400);
or U3839 (N_3839,N_930,N_1368);
or U3840 (N_3840,N_2407,N_412);
xnor U3841 (N_3841,N_441,N_343);
or U3842 (N_3842,N_908,N_1813);
nor U3843 (N_3843,N_1718,N_2393);
and U3844 (N_3844,N_2123,N_740);
nor U3845 (N_3845,N_1204,N_1931);
or U3846 (N_3846,N_388,N_1457);
or U3847 (N_3847,N_2129,N_396);
nor U3848 (N_3848,N_2225,N_2075);
xnor U3849 (N_3849,N_437,N_195);
or U3850 (N_3850,N_1282,N_2495);
or U3851 (N_3851,N_2392,N_463);
or U3852 (N_3852,N_2115,N_1492);
nand U3853 (N_3853,N_2483,N_1710);
or U3854 (N_3854,N_2325,N_681);
or U3855 (N_3855,N_2137,N_1800);
or U3856 (N_3856,N_1773,N_1992);
or U3857 (N_3857,N_1573,N_1485);
nand U3858 (N_3858,N_203,N_1852);
or U3859 (N_3859,N_2381,N_1743);
nand U3860 (N_3860,N_1829,N_2182);
nand U3861 (N_3861,N_1010,N_2359);
or U3862 (N_3862,N_1047,N_1632);
nand U3863 (N_3863,N_1577,N_59);
nor U3864 (N_3864,N_1338,N_322);
nand U3865 (N_3865,N_1161,N_312);
nand U3866 (N_3866,N_2392,N_1200);
nor U3867 (N_3867,N_837,N_1623);
nand U3868 (N_3868,N_754,N_1513);
nor U3869 (N_3869,N_420,N_704);
or U3870 (N_3870,N_2365,N_181);
xor U3871 (N_3871,N_1955,N_38);
nand U3872 (N_3872,N_163,N_292);
and U3873 (N_3873,N_664,N_579);
and U3874 (N_3874,N_464,N_355);
nand U3875 (N_3875,N_225,N_502);
nor U3876 (N_3876,N_1587,N_2187);
xor U3877 (N_3877,N_953,N_681);
nand U3878 (N_3878,N_1433,N_2175);
nand U3879 (N_3879,N_305,N_2024);
and U3880 (N_3880,N_391,N_368);
xor U3881 (N_3881,N_2019,N_27);
or U3882 (N_3882,N_466,N_586);
xnor U3883 (N_3883,N_2255,N_1014);
and U3884 (N_3884,N_2083,N_1805);
and U3885 (N_3885,N_1639,N_1385);
nand U3886 (N_3886,N_513,N_668);
nand U3887 (N_3887,N_1892,N_1838);
and U3888 (N_3888,N_1374,N_1313);
xor U3889 (N_3889,N_307,N_2067);
xor U3890 (N_3890,N_129,N_2140);
xor U3891 (N_3891,N_674,N_1695);
nor U3892 (N_3892,N_448,N_2274);
and U3893 (N_3893,N_2054,N_234);
xor U3894 (N_3894,N_1153,N_1772);
or U3895 (N_3895,N_1205,N_1518);
xnor U3896 (N_3896,N_46,N_2336);
xnor U3897 (N_3897,N_446,N_1187);
nand U3898 (N_3898,N_1324,N_488);
and U3899 (N_3899,N_1714,N_1399);
and U3900 (N_3900,N_594,N_1140);
xnor U3901 (N_3901,N_202,N_1925);
and U3902 (N_3902,N_39,N_233);
nand U3903 (N_3903,N_2305,N_1696);
nor U3904 (N_3904,N_144,N_1631);
xnor U3905 (N_3905,N_319,N_1472);
nand U3906 (N_3906,N_1304,N_1229);
nor U3907 (N_3907,N_904,N_1906);
or U3908 (N_3908,N_410,N_52);
and U3909 (N_3909,N_722,N_750);
nor U3910 (N_3910,N_909,N_1583);
xnor U3911 (N_3911,N_2129,N_522);
and U3912 (N_3912,N_1132,N_595);
xor U3913 (N_3913,N_486,N_2105);
nand U3914 (N_3914,N_2272,N_2340);
xor U3915 (N_3915,N_1086,N_1576);
xnor U3916 (N_3916,N_652,N_959);
nand U3917 (N_3917,N_1279,N_426);
and U3918 (N_3918,N_665,N_810);
xnor U3919 (N_3919,N_139,N_2285);
xor U3920 (N_3920,N_1379,N_1349);
and U3921 (N_3921,N_1410,N_208);
nor U3922 (N_3922,N_1570,N_2023);
xnor U3923 (N_3923,N_1076,N_2381);
or U3924 (N_3924,N_124,N_359);
and U3925 (N_3925,N_729,N_1805);
and U3926 (N_3926,N_223,N_1849);
and U3927 (N_3927,N_2264,N_1933);
and U3928 (N_3928,N_216,N_2422);
and U3929 (N_3929,N_2419,N_2105);
or U3930 (N_3930,N_622,N_71);
xnor U3931 (N_3931,N_177,N_823);
or U3932 (N_3932,N_2050,N_373);
and U3933 (N_3933,N_551,N_1482);
xnor U3934 (N_3934,N_292,N_2249);
nand U3935 (N_3935,N_208,N_1057);
nor U3936 (N_3936,N_2077,N_2400);
nor U3937 (N_3937,N_1901,N_2426);
xnor U3938 (N_3938,N_871,N_1005);
nor U3939 (N_3939,N_2364,N_340);
nand U3940 (N_3940,N_328,N_1237);
nor U3941 (N_3941,N_613,N_1729);
xor U3942 (N_3942,N_674,N_2082);
and U3943 (N_3943,N_818,N_1584);
and U3944 (N_3944,N_710,N_1989);
and U3945 (N_3945,N_567,N_1869);
xor U3946 (N_3946,N_270,N_1344);
nor U3947 (N_3947,N_1189,N_1844);
nand U3948 (N_3948,N_937,N_974);
or U3949 (N_3949,N_986,N_840);
and U3950 (N_3950,N_2343,N_1600);
or U3951 (N_3951,N_543,N_617);
nor U3952 (N_3952,N_47,N_1252);
nand U3953 (N_3953,N_801,N_1026);
nor U3954 (N_3954,N_1561,N_267);
or U3955 (N_3955,N_981,N_723);
and U3956 (N_3956,N_1641,N_2101);
xnor U3957 (N_3957,N_1016,N_1913);
and U3958 (N_3958,N_789,N_2060);
and U3959 (N_3959,N_1900,N_2008);
and U3960 (N_3960,N_1051,N_533);
or U3961 (N_3961,N_2450,N_1555);
nand U3962 (N_3962,N_802,N_2337);
or U3963 (N_3963,N_1827,N_1056);
and U3964 (N_3964,N_880,N_1280);
and U3965 (N_3965,N_1691,N_2402);
or U3966 (N_3966,N_2284,N_2193);
or U3967 (N_3967,N_1288,N_1581);
or U3968 (N_3968,N_78,N_1431);
xor U3969 (N_3969,N_240,N_1773);
nand U3970 (N_3970,N_1206,N_247);
xor U3971 (N_3971,N_2441,N_534);
and U3972 (N_3972,N_213,N_1477);
or U3973 (N_3973,N_335,N_1122);
xor U3974 (N_3974,N_1428,N_779);
and U3975 (N_3975,N_0,N_2449);
xor U3976 (N_3976,N_2449,N_601);
or U3977 (N_3977,N_1196,N_2448);
or U3978 (N_3978,N_1792,N_65);
nand U3979 (N_3979,N_398,N_470);
or U3980 (N_3980,N_1384,N_721);
nand U3981 (N_3981,N_210,N_2061);
nor U3982 (N_3982,N_436,N_2111);
nand U3983 (N_3983,N_1078,N_2220);
or U3984 (N_3984,N_2286,N_597);
nand U3985 (N_3985,N_851,N_478);
nor U3986 (N_3986,N_39,N_182);
and U3987 (N_3987,N_1755,N_961);
and U3988 (N_3988,N_1735,N_1367);
and U3989 (N_3989,N_707,N_1764);
xor U3990 (N_3990,N_558,N_112);
or U3991 (N_3991,N_1531,N_1378);
or U3992 (N_3992,N_938,N_1710);
nor U3993 (N_3993,N_1713,N_1499);
or U3994 (N_3994,N_126,N_1736);
nand U3995 (N_3995,N_381,N_404);
xor U3996 (N_3996,N_2205,N_112);
nand U3997 (N_3997,N_2051,N_1828);
and U3998 (N_3998,N_2284,N_1972);
nor U3999 (N_3999,N_2028,N_353);
nor U4000 (N_4000,N_1381,N_2378);
nor U4001 (N_4001,N_1768,N_968);
and U4002 (N_4002,N_1230,N_2235);
nor U4003 (N_4003,N_139,N_2117);
or U4004 (N_4004,N_2121,N_666);
nor U4005 (N_4005,N_199,N_1577);
and U4006 (N_4006,N_1867,N_1433);
nor U4007 (N_4007,N_2430,N_792);
nor U4008 (N_4008,N_1821,N_1508);
and U4009 (N_4009,N_249,N_108);
and U4010 (N_4010,N_1070,N_239);
xnor U4011 (N_4011,N_491,N_482);
nor U4012 (N_4012,N_837,N_2098);
or U4013 (N_4013,N_814,N_1809);
nor U4014 (N_4014,N_675,N_2073);
nor U4015 (N_4015,N_816,N_1281);
xor U4016 (N_4016,N_1795,N_2167);
xor U4017 (N_4017,N_1211,N_172);
or U4018 (N_4018,N_1196,N_2270);
nand U4019 (N_4019,N_1878,N_257);
nor U4020 (N_4020,N_2260,N_220);
nor U4021 (N_4021,N_201,N_265);
nor U4022 (N_4022,N_2472,N_2172);
or U4023 (N_4023,N_1025,N_2110);
nand U4024 (N_4024,N_1269,N_1418);
or U4025 (N_4025,N_2324,N_1383);
xor U4026 (N_4026,N_125,N_1424);
xor U4027 (N_4027,N_2065,N_592);
nand U4028 (N_4028,N_678,N_1977);
nor U4029 (N_4029,N_638,N_717);
nor U4030 (N_4030,N_1303,N_1981);
xnor U4031 (N_4031,N_588,N_45);
and U4032 (N_4032,N_1303,N_885);
nor U4033 (N_4033,N_318,N_432);
and U4034 (N_4034,N_484,N_2189);
xnor U4035 (N_4035,N_466,N_385);
xnor U4036 (N_4036,N_2082,N_377);
nor U4037 (N_4037,N_2295,N_466);
and U4038 (N_4038,N_595,N_2139);
nor U4039 (N_4039,N_815,N_2290);
nand U4040 (N_4040,N_1798,N_346);
nand U4041 (N_4041,N_716,N_646);
or U4042 (N_4042,N_2354,N_1992);
or U4043 (N_4043,N_2275,N_824);
and U4044 (N_4044,N_2268,N_1843);
nand U4045 (N_4045,N_2173,N_1423);
and U4046 (N_4046,N_553,N_2415);
nor U4047 (N_4047,N_2377,N_2476);
or U4048 (N_4048,N_227,N_997);
or U4049 (N_4049,N_874,N_1415);
or U4050 (N_4050,N_1796,N_739);
and U4051 (N_4051,N_1002,N_1468);
nor U4052 (N_4052,N_1122,N_826);
nand U4053 (N_4053,N_2031,N_1448);
and U4054 (N_4054,N_1087,N_2026);
xor U4055 (N_4055,N_736,N_2403);
nor U4056 (N_4056,N_2305,N_1278);
nand U4057 (N_4057,N_265,N_1041);
and U4058 (N_4058,N_1837,N_1805);
xnor U4059 (N_4059,N_1884,N_2359);
nand U4060 (N_4060,N_400,N_1785);
xnor U4061 (N_4061,N_1506,N_173);
nand U4062 (N_4062,N_2019,N_895);
nand U4063 (N_4063,N_1162,N_1793);
nand U4064 (N_4064,N_801,N_633);
and U4065 (N_4065,N_331,N_3);
nand U4066 (N_4066,N_779,N_2445);
nor U4067 (N_4067,N_2478,N_2139);
nand U4068 (N_4068,N_611,N_1234);
or U4069 (N_4069,N_194,N_1422);
xnor U4070 (N_4070,N_329,N_323);
nand U4071 (N_4071,N_1547,N_1281);
and U4072 (N_4072,N_1266,N_22);
or U4073 (N_4073,N_107,N_2269);
and U4074 (N_4074,N_1252,N_2306);
nand U4075 (N_4075,N_1674,N_361);
or U4076 (N_4076,N_1566,N_2320);
nor U4077 (N_4077,N_945,N_2068);
and U4078 (N_4078,N_1044,N_599);
or U4079 (N_4079,N_1471,N_620);
nand U4080 (N_4080,N_535,N_881);
nor U4081 (N_4081,N_564,N_1812);
nand U4082 (N_4082,N_1661,N_1522);
xor U4083 (N_4083,N_2041,N_2308);
nand U4084 (N_4084,N_575,N_2345);
xnor U4085 (N_4085,N_2092,N_1614);
nand U4086 (N_4086,N_791,N_1197);
nand U4087 (N_4087,N_1469,N_1870);
nand U4088 (N_4088,N_631,N_626);
and U4089 (N_4089,N_1316,N_1375);
nand U4090 (N_4090,N_2199,N_370);
nand U4091 (N_4091,N_1425,N_1673);
and U4092 (N_4092,N_1532,N_392);
nand U4093 (N_4093,N_361,N_2491);
or U4094 (N_4094,N_699,N_1548);
nand U4095 (N_4095,N_1491,N_67);
and U4096 (N_4096,N_192,N_469);
or U4097 (N_4097,N_2034,N_2366);
or U4098 (N_4098,N_2277,N_1290);
or U4099 (N_4099,N_197,N_333);
nor U4100 (N_4100,N_1315,N_88);
nor U4101 (N_4101,N_2034,N_556);
xor U4102 (N_4102,N_1523,N_272);
nand U4103 (N_4103,N_1910,N_2125);
xnor U4104 (N_4104,N_918,N_544);
and U4105 (N_4105,N_250,N_2016);
or U4106 (N_4106,N_469,N_139);
or U4107 (N_4107,N_123,N_1606);
nor U4108 (N_4108,N_1475,N_1137);
or U4109 (N_4109,N_1388,N_1462);
and U4110 (N_4110,N_507,N_1636);
xor U4111 (N_4111,N_429,N_1966);
nand U4112 (N_4112,N_977,N_1416);
xor U4113 (N_4113,N_1836,N_1722);
xor U4114 (N_4114,N_1756,N_1386);
nor U4115 (N_4115,N_829,N_325);
nand U4116 (N_4116,N_532,N_1433);
nand U4117 (N_4117,N_2191,N_2101);
nand U4118 (N_4118,N_1010,N_1224);
xnor U4119 (N_4119,N_1562,N_2300);
nand U4120 (N_4120,N_1197,N_1614);
nor U4121 (N_4121,N_1236,N_2179);
xor U4122 (N_4122,N_1853,N_2140);
nor U4123 (N_4123,N_987,N_605);
nor U4124 (N_4124,N_531,N_2048);
xnor U4125 (N_4125,N_2378,N_153);
xor U4126 (N_4126,N_2113,N_1394);
and U4127 (N_4127,N_2093,N_2481);
or U4128 (N_4128,N_2491,N_2159);
nor U4129 (N_4129,N_189,N_2236);
nor U4130 (N_4130,N_2388,N_1948);
or U4131 (N_4131,N_983,N_2071);
and U4132 (N_4132,N_1323,N_73);
nand U4133 (N_4133,N_1998,N_454);
xnor U4134 (N_4134,N_1581,N_797);
or U4135 (N_4135,N_867,N_1785);
xor U4136 (N_4136,N_1053,N_668);
nand U4137 (N_4137,N_2261,N_192);
and U4138 (N_4138,N_2018,N_1235);
nand U4139 (N_4139,N_25,N_2385);
xnor U4140 (N_4140,N_1379,N_2497);
and U4141 (N_4141,N_1155,N_1542);
xor U4142 (N_4142,N_1132,N_2361);
nand U4143 (N_4143,N_933,N_712);
nand U4144 (N_4144,N_2498,N_778);
nor U4145 (N_4145,N_2031,N_1425);
nor U4146 (N_4146,N_1256,N_493);
or U4147 (N_4147,N_542,N_246);
xor U4148 (N_4148,N_1390,N_109);
or U4149 (N_4149,N_1838,N_1078);
xnor U4150 (N_4150,N_324,N_1580);
or U4151 (N_4151,N_1525,N_2045);
and U4152 (N_4152,N_862,N_1961);
nor U4153 (N_4153,N_2428,N_1083);
and U4154 (N_4154,N_1354,N_1701);
nand U4155 (N_4155,N_233,N_1315);
and U4156 (N_4156,N_2359,N_2232);
xnor U4157 (N_4157,N_536,N_202);
and U4158 (N_4158,N_233,N_175);
nand U4159 (N_4159,N_1192,N_1220);
nand U4160 (N_4160,N_2349,N_766);
or U4161 (N_4161,N_648,N_1132);
nand U4162 (N_4162,N_987,N_947);
or U4163 (N_4163,N_808,N_2418);
nor U4164 (N_4164,N_529,N_825);
and U4165 (N_4165,N_1549,N_970);
nand U4166 (N_4166,N_996,N_325);
nand U4167 (N_4167,N_2214,N_1323);
xor U4168 (N_4168,N_2082,N_1744);
and U4169 (N_4169,N_1004,N_367);
nor U4170 (N_4170,N_1445,N_896);
xor U4171 (N_4171,N_2033,N_1485);
and U4172 (N_4172,N_1178,N_2265);
xor U4173 (N_4173,N_1502,N_2338);
and U4174 (N_4174,N_2384,N_516);
or U4175 (N_4175,N_2005,N_711);
and U4176 (N_4176,N_585,N_589);
and U4177 (N_4177,N_151,N_2252);
nor U4178 (N_4178,N_2278,N_10);
nor U4179 (N_4179,N_30,N_2101);
xnor U4180 (N_4180,N_2112,N_172);
nor U4181 (N_4181,N_359,N_837);
nand U4182 (N_4182,N_1444,N_536);
xor U4183 (N_4183,N_1553,N_2336);
nand U4184 (N_4184,N_1236,N_170);
nor U4185 (N_4185,N_547,N_269);
nor U4186 (N_4186,N_1802,N_1070);
xor U4187 (N_4187,N_1234,N_188);
xnor U4188 (N_4188,N_1294,N_1473);
xor U4189 (N_4189,N_2472,N_1519);
or U4190 (N_4190,N_2247,N_287);
and U4191 (N_4191,N_693,N_1956);
and U4192 (N_4192,N_1602,N_980);
nand U4193 (N_4193,N_2337,N_598);
nand U4194 (N_4194,N_2073,N_2099);
and U4195 (N_4195,N_56,N_674);
nor U4196 (N_4196,N_1507,N_187);
and U4197 (N_4197,N_2295,N_1254);
xor U4198 (N_4198,N_246,N_979);
nand U4199 (N_4199,N_1637,N_1405);
or U4200 (N_4200,N_1745,N_2481);
xnor U4201 (N_4201,N_2264,N_2440);
and U4202 (N_4202,N_709,N_1634);
nor U4203 (N_4203,N_2363,N_44);
xnor U4204 (N_4204,N_2158,N_704);
and U4205 (N_4205,N_2103,N_1933);
nand U4206 (N_4206,N_797,N_2106);
and U4207 (N_4207,N_1811,N_1369);
xnor U4208 (N_4208,N_1655,N_1019);
nor U4209 (N_4209,N_1723,N_352);
nor U4210 (N_4210,N_339,N_1494);
xnor U4211 (N_4211,N_2412,N_876);
nor U4212 (N_4212,N_300,N_861);
xor U4213 (N_4213,N_1757,N_2023);
or U4214 (N_4214,N_274,N_108);
xor U4215 (N_4215,N_1128,N_615);
and U4216 (N_4216,N_1117,N_1091);
xor U4217 (N_4217,N_2349,N_562);
xnor U4218 (N_4218,N_2024,N_2334);
nor U4219 (N_4219,N_2160,N_937);
xor U4220 (N_4220,N_1452,N_1524);
nand U4221 (N_4221,N_1732,N_2465);
nor U4222 (N_4222,N_1422,N_332);
xor U4223 (N_4223,N_1544,N_2004);
or U4224 (N_4224,N_406,N_1268);
or U4225 (N_4225,N_2382,N_1624);
nor U4226 (N_4226,N_2224,N_1475);
nand U4227 (N_4227,N_1045,N_1282);
or U4228 (N_4228,N_124,N_474);
and U4229 (N_4229,N_469,N_959);
nand U4230 (N_4230,N_671,N_38);
and U4231 (N_4231,N_446,N_1540);
or U4232 (N_4232,N_322,N_140);
and U4233 (N_4233,N_587,N_265);
and U4234 (N_4234,N_1486,N_346);
xor U4235 (N_4235,N_669,N_1000);
nor U4236 (N_4236,N_2462,N_868);
nand U4237 (N_4237,N_867,N_2400);
nor U4238 (N_4238,N_1561,N_1260);
and U4239 (N_4239,N_809,N_651);
and U4240 (N_4240,N_1861,N_1526);
nor U4241 (N_4241,N_2142,N_2349);
and U4242 (N_4242,N_549,N_2315);
xnor U4243 (N_4243,N_2359,N_23);
or U4244 (N_4244,N_1817,N_1358);
or U4245 (N_4245,N_1711,N_792);
and U4246 (N_4246,N_2295,N_1623);
or U4247 (N_4247,N_2401,N_906);
nand U4248 (N_4248,N_98,N_2090);
xnor U4249 (N_4249,N_608,N_1943);
and U4250 (N_4250,N_1789,N_2216);
xor U4251 (N_4251,N_37,N_1341);
nor U4252 (N_4252,N_1290,N_857);
xnor U4253 (N_4253,N_835,N_2026);
and U4254 (N_4254,N_957,N_337);
or U4255 (N_4255,N_1436,N_850);
xnor U4256 (N_4256,N_981,N_805);
nand U4257 (N_4257,N_317,N_1605);
and U4258 (N_4258,N_763,N_664);
nor U4259 (N_4259,N_699,N_333);
or U4260 (N_4260,N_545,N_1143);
or U4261 (N_4261,N_299,N_27);
and U4262 (N_4262,N_2382,N_1410);
nor U4263 (N_4263,N_1246,N_278);
or U4264 (N_4264,N_809,N_774);
and U4265 (N_4265,N_2386,N_1991);
xor U4266 (N_4266,N_1550,N_1572);
nor U4267 (N_4267,N_1246,N_798);
xnor U4268 (N_4268,N_2304,N_355);
or U4269 (N_4269,N_809,N_615);
nand U4270 (N_4270,N_853,N_834);
xnor U4271 (N_4271,N_1058,N_1525);
nor U4272 (N_4272,N_476,N_2020);
xnor U4273 (N_4273,N_1524,N_317);
or U4274 (N_4274,N_2274,N_2365);
nor U4275 (N_4275,N_1513,N_1694);
and U4276 (N_4276,N_1637,N_1635);
or U4277 (N_4277,N_2301,N_1416);
or U4278 (N_4278,N_662,N_763);
nor U4279 (N_4279,N_1943,N_2269);
or U4280 (N_4280,N_1019,N_51);
or U4281 (N_4281,N_481,N_1847);
and U4282 (N_4282,N_2362,N_2278);
and U4283 (N_4283,N_2499,N_1547);
nand U4284 (N_4284,N_521,N_1787);
nor U4285 (N_4285,N_2258,N_2414);
nand U4286 (N_4286,N_1550,N_1903);
nand U4287 (N_4287,N_2148,N_1851);
xor U4288 (N_4288,N_1000,N_2034);
and U4289 (N_4289,N_1618,N_411);
nor U4290 (N_4290,N_802,N_1543);
xor U4291 (N_4291,N_1232,N_1165);
or U4292 (N_4292,N_76,N_570);
and U4293 (N_4293,N_1025,N_1663);
and U4294 (N_4294,N_205,N_1358);
nor U4295 (N_4295,N_1863,N_770);
nand U4296 (N_4296,N_470,N_164);
nor U4297 (N_4297,N_2388,N_626);
xor U4298 (N_4298,N_2164,N_2338);
xor U4299 (N_4299,N_2132,N_362);
nand U4300 (N_4300,N_1799,N_2453);
nor U4301 (N_4301,N_189,N_2216);
xnor U4302 (N_4302,N_232,N_2496);
and U4303 (N_4303,N_2378,N_875);
nor U4304 (N_4304,N_775,N_1944);
nand U4305 (N_4305,N_373,N_215);
and U4306 (N_4306,N_235,N_993);
nor U4307 (N_4307,N_2087,N_493);
xor U4308 (N_4308,N_59,N_953);
xnor U4309 (N_4309,N_2211,N_130);
or U4310 (N_4310,N_651,N_1733);
and U4311 (N_4311,N_2324,N_1499);
nand U4312 (N_4312,N_1631,N_1446);
xnor U4313 (N_4313,N_1913,N_2214);
nor U4314 (N_4314,N_1791,N_842);
or U4315 (N_4315,N_819,N_424);
and U4316 (N_4316,N_1142,N_1120);
nor U4317 (N_4317,N_2382,N_1039);
nor U4318 (N_4318,N_20,N_697);
xnor U4319 (N_4319,N_1448,N_1);
nand U4320 (N_4320,N_1377,N_1779);
nor U4321 (N_4321,N_952,N_1050);
and U4322 (N_4322,N_276,N_1545);
or U4323 (N_4323,N_466,N_705);
nand U4324 (N_4324,N_741,N_1622);
and U4325 (N_4325,N_1837,N_596);
nor U4326 (N_4326,N_35,N_2283);
or U4327 (N_4327,N_659,N_514);
and U4328 (N_4328,N_898,N_51);
and U4329 (N_4329,N_2367,N_1908);
or U4330 (N_4330,N_1918,N_2031);
nor U4331 (N_4331,N_93,N_1371);
xor U4332 (N_4332,N_1243,N_856);
nand U4333 (N_4333,N_477,N_402);
xor U4334 (N_4334,N_796,N_976);
nand U4335 (N_4335,N_564,N_1982);
and U4336 (N_4336,N_1665,N_1633);
nand U4337 (N_4337,N_1052,N_1092);
nand U4338 (N_4338,N_2339,N_2422);
xor U4339 (N_4339,N_671,N_1188);
xnor U4340 (N_4340,N_994,N_1557);
nor U4341 (N_4341,N_1033,N_950);
nor U4342 (N_4342,N_193,N_2017);
nand U4343 (N_4343,N_1074,N_1988);
or U4344 (N_4344,N_1587,N_552);
or U4345 (N_4345,N_1156,N_148);
nor U4346 (N_4346,N_62,N_1);
xor U4347 (N_4347,N_1253,N_2220);
xor U4348 (N_4348,N_593,N_1839);
nand U4349 (N_4349,N_2170,N_741);
and U4350 (N_4350,N_1204,N_302);
or U4351 (N_4351,N_496,N_1500);
nor U4352 (N_4352,N_1453,N_1030);
nor U4353 (N_4353,N_1313,N_137);
nor U4354 (N_4354,N_1054,N_1848);
or U4355 (N_4355,N_197,N_593);
nand U4356 (N_4356,N_752,N_2329);
and U4357 (N_4357,N_1569,N_1860);
or U4358 (N_4358,N_82,N_160);
or U4359 (N_4359,N_2139,N_1214);
and U4360 (N_4360,N_2012,N_837);
xor U4361 (N_4361,N_1020,N_2033);
nand U4362 (N_4362,N_48,N_1310);
xor U4363 (N_4363,N_2004,N_1745);
nor U4364 (N_4364,N_708,N_1502);
xor U4365 (N_4365,N_2181,N_371);
nand U4366 (N_4366,N_146,N_2422);
nor U4367 (N_4367,N_1069,N_2322);
xor U4368 (N_4368,N_1710,N_1608);
or U4369 (N_4369,N_376,N_574);
nand U4370 (N_4370,N_1790,N_1943);
nor U4371 (N_4371,N_1273,N_1860);
nand U4372 (N_4372,N_1896,N_894);
and U4373 (N_4373,N_2090,N_1758);
nand U4374 (N_4374,N_239,N_210);
xor U4375 (N_4375,N_1398,N_721);
or U4376 (N_4376,N_1608,N_129);
nand U4377 (N_4377,N_1456,N_2336);
xnor U4378 (N_4378,N_1895,N_1844);
and U4379 (N_4379,N_635,N_145);
xor U4380 (N_4380,N_282,N_1678);
or U4381 (N_4381,N_2366,N_758);
nand U4382 (N_4382,N_1620,N_1062);
or U4383 (N_4383,N_1843,N_917);
nand U4384 (N_4384,N_1408,N_1534);
and U4385 (N_4385,N_1185,N_1473);
or U4386 (N_4386,N_2438,N_233);
xnor U4387 (N_4387,N_844,N_1245);
or U4388 (N_4388,N_837,N_266);
xnor U4389 (N_4389,N_701,N_2135);
and U4390 (N_4390,N_210,N_1939);
and U4391 (N_4391,N_1217,N_2214);
nor U4392 (N_4392,N_260,N_1405);
and U4393 (N_4393,N_340,N_127);
and U4394 (N_4394,N_71,N_1278);
and U4395 (N_4395,N_722,N_1992);
or U4396 (N_4396,N_2308,N_1183);
xor U4397 (N_4397,N_1544,N_1119);
and U4398 (N_4398,N_1357,N_1707);
and U4399 (N_4399,N_816,N_2186);
and U4400 (N_4400,N_519,N_1952);
nand U4401 (N_4401,N_706,N_1289);
xnor U4402 (N_4402,N_1718,N_2127);
xnor U4403 (N_4403,N_2028,N_1596);
or U4404 (N_4404,N_613,N_1758);
nand U4405 (N_4405,N_1358,N_180);
nor U4406 (N_4406,N_2308,N_1919);
xor U4407 (N_4407,N_981,N_1426);
nor U4408 (N_4408,N_1570,N_1730);
nor U4409 (N_4409,N_2356,N_2012);
nor U4410 (N_4410,N_1488,N_1368);
and U4411 (N_4411,N_2392,N_2227);
xnor U4412 (N_4412,N_2004,N_2420);
xnor U4413 (N_4413,N_1088,N_701);
and U4414 (N_4414,N_1931,N_2243);
or U4415 (N_4415,N_536,N_1973);
nor U4416 (N_4416,N_17,N_63);
or U4417 (N_4417,N_218,N_2072);
or U4418 (N_4418,N_1483,N_1690);
nor U4419 (N_4419,N_2107,N_1351);
or U4420 (N_4420,N_2004,N_1159);
nand U4421 (N_4421,N_2365,N_1498);
xor U4422 (N_4422,N_806,N_1056);
xor U4423 (N_4423,N_1464,N_1633);
or U4424 (N_4424,N_1281,N_2403);
nand U4425 (N_4425,N_2410,N_1949);
nand U4426 (N_4426,N_1055,N_499);
and U4427 (N_4427,N_1677,N_657);
nor U4428 (N_4428,N_795,N_1542);
or U4429 (N_4429,N_783,N_1109);
nand U4430 (N_4430,N_982,N_2435);
nor U4431 (N_4431,N_1659,N_2124);
or U4432 (N_4432,N_1732,N_725);
and U4433 (N_4433,N_179,N_1209);
or U4434 (N_4434,N_427,N_1287);
xor U4435 (N_4435,N_2426,N_850);
nor U4436 (N_4436,N_754,N_1278);
nand U4437 (N_4437,N_73,N_882);
xor U4438 (N_4438,N_928,N_846);
nand U4439 (N_4439,N_354,N_2292);
nor U4440 (N_4440,N_1002,N_2441);
or U4441 (N_4441,N_744,N_706);
xor U4442 (N_4442,N_2050,N_2385);
nor U4443 (N_4443,N_309,N_360);
and U4444 (N_4444,N_1642,N_1610);
and U4445 (N_4445,N_122,N_1891);
nand U4446 (N_4446,N_724,N_636);
or U4447 (N_4447,N_1224,N_1563);
xor U4448 (N_4448,N_669,N_1808);
or U4449 (N_4449,N_1653,N_907);
and U4450 (N_4450,N_1480,N_483);
xnor U4451 (N_4451,N_1263,N_1759);
nor U4452 (N_4452,N_1967,N_2316);
and U4453 (N_4453,N_2108,N_1816);
and U4454 (N_4454,N_1169,N_2027);
or U4455 (N_4455,N_1934,N_2499);
nor U4456 (N_4456,N_1892,N_1306);
nor U4457 (N_4457,N_540,N_669);
and U4458 (N_4458,N_914,N_1683);
or U4459 (N_4459,N_1203,N_871);
and U4460 (N_4460,N_1175,N_534);
nand U4461 (N_4461,N_1999,N_842);
or U4462 (N_4462,N_359,N_83);
or U4463 (N_4463,N_1271,N_1452);
nand U4464 (N_4464,N_2417,N_675);
xnor U4465 (N_4465,N_741,N_408);
nor U4466 (N_4466,N_231,N_559);
or U4467 (N_4467,N_1401,N_2087);
or U4468 (N_4468,N_1480,N_1726);
nand U4469 (N_4469,N_1686,N_1454);
or U4470 (N_4470,N_1088,N_735);
or U4471 (N_4471,N_1763,N_1200);
nand U4472 (N_4472,N_562,N_1302);
xor U4473 (N_4473,N_6,N_46);
and U4474 (N_4474,N_1677,N_2208);
nor U4475 (N_4475,N_1541,N_1996);
and U4476 (N_4476,N_1073,N_1159);
nor U4477 (N_4477,N_269,N_345);
xnor U4478 (N_4478,N_2320,N_300);
xor U4479 (N_4479,N_2431,N_1379);
xor U4480 (N_4480,N_422,N_1762);
and U4481 (N_4481,N_498,N_570);
nor U4482 (N_4482,N_1253,N_463);
nand U4483 (N_4483,N_1749,N_2106);
nand U4484 (N_4484,N_210,N_1844);
xor U4485 (N_4485,N_1503,N_453);
nor U4486 (N_4486,N_2223,N_735);
and U4487 (N_4487,N_662,N_1351);
xnor U4488 (N_4488,N_1535,N_1487);
xnor U4489 (N_4489,N_922,N_2350);
nor U4490 (N_4490,N_2043,N_940);
nand U4491 (N_4491,N_113,N_1029);
nand U4492 (N_4492,N_618,N_660);
or U4493 (N_4493,N_828,N_1233);
nor U4494 (N_4494,N_145,N_2322);
or U4495 (N_4495,N_1408,N_2213);
and U4496 (N_4496,N_1731,N_2059);
xnor U4497 (N_4497,N_1448,N_2441);
or U4498 (N_4498,N_693,N_1081);
or U4499 (N_4499,N_572,N_1840);
nand U4500 (N_4500,N_1632,N_1245);
or U4501 (N_4501,N_626,N_1571);
or U4502 (N_4502,N_228,N_1071);
nand U4503 (N_4503,N_2184,N_2335);
nand U4504 (N_4504,N_1572,N_32);
and U4505 (N_4505,N_1925,N_1361);
nand U4506 (N_4506,N_842,N_417);
xnor U4507 (N_4507,N_1674,N_860);
or U4508 (N_4508,N_2341,N_711);
or U4509 (N_4509,N_1419,N_2366);
nor U4510 (N_4510,N_320,N_1635);
nand U4511 (N_4511,N_1292,N_447);
or U4512 (N_4512,N_1794,N_328);
nand U4513 (N_4513,N_1639,N_2346);
nor U4514 (N_4514,N_355,N_539);
or U4515 (N_4515,N_2152,N_2279);
nor U4516 (N_4516,N_1445,N_1261);
xor U4517 (N_4517,N_1605,N_144);
xor U4518 (N_4518,N_1704,N_1163);
nand U4519 (N_4519,N_2282,N_579);
nand U4520 (N_4520,N_1568,N_2250);
nor U4521 (N_4521,N_2266,N_1498);
and U4522 (N_4522,N_932,N_2455);
nor U4523 (N_4523,N_2015,N_511);
nor U4524 (N_4524,N_2444,N_592);
or U4525 (N_4525,N_1050,N_1249);
and U4526 (N_4526,N_962,N_380);
xnor U4527 (N_4527,N_338,N_927);
or U4528 (N_4528,N_1920,N_2446);
nor U4529 (N_4529,N_203,N_2359);
and U4530 (N_4530,N_2139,N_1430);
xnor U4531 (N_4531,N_717,N_1059);
xor U4532 (N_4532,N_1570,N_374);
nand U4533 (N_4533,N_2134,N_313);
nand U4534 (N_4534,N_1260,N_2129);
xnor U4535 (N_4535,N_2410,N_2377);
and U4536 (N_4536,N_394,N_148);
nor U4537 (N_4537,N_1471,N_363);
nand U4538 (N_4538,N_499,N_2209);
xnor U4539 (N_4539,N_1951,N_2456);
or U4540 (N_4540,N_2419,N_335);
or U4541 (N_4541,N_588,N_1305);
xnor U4542 (N_4542,N_1924,N_1535);
nor U4543 (N_4543,N_802,N_1915);
nand U4544 (N_4544,N_1878,N_1842);
nor U4545 (N_4545,N_504,N_183);
and U4546 (N_4546,N_1754,N_1039);
nor U4547 (N_4547,N_2313,N_1658);
and U4548 (N_4548,N_1740,N_1151);
xnor U4549 (N_4549,N_1427,N_523);
and U4550 (N_4550,N_1643,N_406);
or U4551 (N_4551,N_1223,N_137);
nand U4552 (N_4552,N_1520,N_2364);
xnor U4553 (N_4553,N_1691,N_2461);
or U4554 (N_4554,N_307,N_1144);
nor U4555 (N_4555,N_1390,N_2116);
and U4556 (N_4556,N_1574,N_1805);
xnor U4557 (N_4557,N_1676,N_2403);
or U4558 (N_4558,N_1974,N_283);
nand U4559 (N_4559,N_1969,N_157);
or U4560 (N_4560,N_2183,N_115);
nor U4561 (N_4561,N_2010,N_2176);
or U4562 (N_4562,N_1354,N_822);
nor U4563 (N_4563,N_1683,N_1237);
and U4564 (N_4564,N_1536,N_1397);
nor U4565 (N_4565,N_1799,N_1888);
nor U4566 (N_4566,N_59,N_1902);
or U4567 (N_4567,N_1711,N_842);
xnor U4568 (N_4568,N_2127,N_247);
or U4569 (N_4569,N_2238,N_1626);
xor U4570 (N_4570,N_169,N_540);
and U4571 (N_4571,N_550,N_1852);
nand U4572 (N_4572,N_1517,N_143);
or U4573 (N_4573,N_913,N_1198);
nand U4574 (N_4574,N_2407,N_1763);
nor U4575 (N_4575,N_962,N_1524);
and U4576 (N_4576,N_623,N_649);
nor U4577 (N_4577,N_2012,N_1457);
xnor U4578 (N_4578,N_1261,N_339);
nor U4579 (N_4579,N_1196,N_1899);
nor U4580 (N_4580,N_2472,N_1804);
xor U4581 (N_4581,N_374,N_2350);
or U4582 (N_4582,N_1945,N_452);
or U4583 (N_4583,N_563,N_2073);
nor U4584 (N_4584,N_1868,N_2093);
xor U4585 (N_4585,N_232,N_1879);
or U4586 (N_4586,N_1548,N_262);
nand U4587 (N_4587,N_30,N_1041);
and U4588 (N_4588,N_2114,N_2016);
and U4589 (N_4589,N_2337,N_403);
nand U4590 (N_4590,N_1358,N_995);
nor U4591 (N_4591,N_350,N_1429);
xnor U4592 (N_4592,N_124,N_837);
nor U4593 (N_4593,N_1233,N_484);
nand U4594 (N_4594,N_277,N_1803);
and U4595 (N_4595,N_577,N_2032);
nor U4596 (N_4596,N_220,N_2080);
nor U4597 (N_4597,N_1386,N_172);
nand U4598 (N_4598,N_662,N_497);
nor U4599 (N_4599,N_1032,N_137);
and U4600 (N_4600,N_1416,N_186);
or U4601 (N_4601,N_1645,N_1178);
nand U4602 (N_4602,N_1267,N_924);
nor U4603 (N_4603,N_715,N_1039);
xnor U4604 (N_4604,N_86,N_822);
nand U4605 (N_4605,N_2258,N_2474);
nand U4606 (N_4606,N_36,N_2059);
nand U4607 (N_4607,N_325,N_1254);
nand U4608 (N_4608,N_1581,N_1898);
xnor U4609 (N_4609,N_2392,N_2031);
nor U4610 (N_4610,N_1135,N_1485);
or U4611 (N_4611,N_2355,N_1);
nand U4612 (N_4612,N_2084,N_788);
nor U4613 (N_4613,N_833,N_346);
and U4614 (N_4614,N_631,N_2036);
and U4615 (N_4615,N_1998,N_2226);
nor U4616 (N_4616,N_326,N_1414);
nand U4617 (N_4617,N_259,N_1493);
or U4618 (N_4618,N_2073,N_2427);
or U4619 (N_4619,N_497,N_1903);
and U4620 (N_4620,N_351,N_1775);
nand U4621 (N_4621,N_2478,N_1131);
and U4622 (N_4622,N_1011,N_1159);
nor U4623 (N_4623,N_209,N_1183);
nor U4624 (N_4624,N_1443,N_1976);
nand U4625 (N_4625,N_1003,N_1662);
nand U4626 (N_4626,N_2260,N_1039);
nand U4627 (N_4627,N_1890,N_101);
or U4628 (N_4628,N_1310,N_679);
xor U4629 (N_4629,N_846,N_1954);
and U4630 (N_4630,N_642,N_2276);
nand U4631 (N_4631,N_1229,N_1884);
and U4632 (N_4632,N_346,N_1512);
and U4633 (N_4633,N_1534,N_807);
or U4634 (N_4634,N_290,N_2162);
nor U4635 (N_4635,N_2344,N_580);
xor U4636 (N_4636,N_118,N_480);
nor U4637 (N_4637,N_777,N_2378);
xor U4638 (N_4638,N_372,N_1112);
and U4639 (N_4639,N_785,N_341);
or U4640 (N_4640,N_1212,N_11);
nor U4641 (N_4641,N_744,N_634);
nand U4642 (N_4642,N_1840,N_2165);
nand U4643 (N_4643,N_1819,N_878);
and U4644 (N_4644,N_1927,N_1241);
nor U4645 (N_4645,N_377,N_1996);
or U4646 (N_4646,N_1726,N_2450);
or U4647 (N_4647,N_1572,N_1512);
or U4648 (N_4648,N_388,N_2338);
and U4649 (N_4649,N_1807,N_1404);
xor U4650 (N_4650,N_748,N_1658);
or U4651 (N_4651,N_197,N_94);
and U4652 (N_4652,N_0,N_994);
nor U4653 (N_4653,N_1245,N_475);
and U4654 (N_4654,N_971,N_1072);
or U4655 (N_4655,N_1142,N_2020);
nand U4656 (N_4656,N_841,N_1204);
xnor U4657 (N_4657,N_152,N_1791);
nor U4658 (N_4658,N_1758,N_232);
or U4659 (N_4659,N_2475,N_1432);
nand U4660 (N_4660,N_729,N_1166);
or U4661 (N_4661,N_781,N_1953);
and U4662 (N_4662,N_1020,N_821);
or U4663 (N_4663,N_695,N_2162);
nand U4664 (N_4664,N_576,N_1409);
and U4665 (N_4665,N_1949,N_115);
and U4666 (N_4666,N_2393,N_1743);
xor U4667 (N_4667,N_2475,N_136);
and U4668 (N_4668,N_201,N_1763);
xnor U4669 (N_4669,N_1813,N_360);
and U4670 (N_4670,N_1156,N_1867);
xnor U4671 (N_4671,N_932,N_1696);
nor U4672 (N_4672,N_633,N_1542);
xor U4673 (N_4673,N_3,N_1424);
nand U4674 (N_4674,N_1298,N_242);
or U4675 (N_4675,N_1696,N_348);
nor U4676 (N_4676,N_546,N_1529);
or U4677 (N_4677,N_2100,N_1715);
or U4678 (N_4678,N_567,N_1945);
nand U4679 (N_4679,N_812,N_2261);
xnor U4680 (N_4680,N_1624,N_2438);
and U4681 (N_4681,N_1016,N_919);
nor U4682 (N_4682,N_2389,N_1482);
xor U4683 (N_4683,N_150,N_2144);
or U4684 (N_4684,N_405,N_652);
xnor U4685 (N_4685,N_826,N_1327);
or U4686 (N_4686,N_1006,N_2077);
nand U4687 (N_4687,N_987,N_949);
and U4688 (N_4688,N_1340,N_1776);
and U4689 (N_4689,N_908,N_2226);
xnor U4690 (N_4690,N_1111,N_1589);
nor U4691 (N_4691,N_1923,N_1739);
and U4692 (N_4692,N_847,N_1820);
and U4693 (N_4693,N_1691,N_273);
xnor U4694 (N_4694,N_2351,N_2439);
xor U4695 (N_4695,N_218,N_2044);
nor U4696 (N_4696,N_2103,N_2428);
nor U4697 (N_4697,N_2268,N_2313);
nand U4698 (N_4698,N_1771,N_2118);
and U4699 (N_4699,N_987,N_1109);
and U4700 (N_4700,N_2140,N_1415);
and U4701 (N_4701,N_1666,N_920);
nor U4702 (N_4702,N_811,N_401);
and U4703 (N_4703,N_1685,N_1506);
and U4704 (N_4704,N_284,N_55);
nand U4705 (N_4705,N_24,N_388);
and U4706 (N_4706,N_1671,N_1481);
nand U4707 (N_4707,N_2419,N_587);
nor U4708 (N_4708,N_433,N_1377);
and U4709 (N_4709,N_1699,N_1617);
nand U4710 (N_4710,N_978,N_320);
or U4711 (N_4711,N_312,N_1417);
xor U4712 (N_4712,N_1383,N_420);
or U4713 (N_4713,N_2391,N_1306);
and U4714 (N_4714,N_1195,N_376);
and U4715 (N_4715,N_1937,N_1725);
nand U4716 (N_4716,N_1783,N_2297);
and U4717 (N_4717,N_648,N_417);
or U4718 (N_4718,N_247,N_1213);
nand U4719 (N_4719,N_1630,N_1842);
or U4720 (N_4720,N_897,N_788);
nand U4721 (N_4721,N_291,N_332);
nor U4722 (N_4722,N_1893,N_2034);
or U4723 (N_4723,N_2155,N_300);
xnor U4724 (N_4724,N_2269,N_758);
xor U4725 (N_4725,N_822,N_1720);
xor U4726 (N_4726,N_434,N_990);
nor U4727 (N_4727,N_561,N_1405);
xnor U4728 (N_4728,N_800,N_620);
nor U4729 (N_4729,N_1167,N_1139);
nor U4730 (N_4730,N_1978,N_376);
nor U4731 (N_4731,N_1298,N_1925);
xor U4732 (N_4732,N_2172,N_1448);
xnor U4733 (N_4733,N_2036,N_2397);
and U4734 (N_4734,N_782,N_802);
and U4735 (N_4735,N_565,N_857);
nor U4736 (N_4736,N_289,N_1553);
xor U4737 (N_4737,N_1460,N_2327);
xor U4738 (N_4738,N_1765,N_962);
or U4739 (N_4739,N_797,N_232);
or U4740 (N_4740,N_870,N_1999);
xnor U4741 (N_4741,N_602,N_1188);
or U4742 (N_4742,N_644,N_653);
or U4743 (N_4743,N_2468,N_1670);
or U4744 (N_4744,N_1455,N_1371);
nand U4745 (N_4745,N_712,N_315);
nor U4746 (N_4746,N_1037,N_1881);
xnor U4747 (N_4747,N_2309,N_2227);
and U4748 (N_4748,N_1137,N_2098);
or U4749 (N_4749,N_300,N_955);
or U4750 (N_4750,N_558,N_1632);
nand U4751 (N_4751,N_142,N_1472);
nand U4752 (N_4752,N_1870,N_459);
nand U4753 (N_4753,N_1395,N_991);
nor U4754 (N_4754,N_2052,N_2007);
xor U4755 (N_4755,N_1917,N_1871);
xor U4756 (N_4756,N_1643,N_519);
xor U4757 (N_4757,N_1225,N_620);
and U4758 (N_4758,N_1391,N_605);
xnor U4759 (N_4759,N_2424,N_1908);
and U4760 (N_4760,N_189,N_1773);
and U4761 (N_4761,N_401,N_250);
nor U4762 (N_4762,N_593,N_1251);
xor U4763 (N_4763,N_1497,N_1631);
nor U4764 (N_4764,N_247,N_1094);
or U4765 (N_4765,N_619,N_132);
nand U4766 (N_4766,N_2374,N_311);
xnor U4767 (N_4767,N_274,N_1488);
xor U4768 (N_4768,N_1780,N_1447);
or U4769 (N_4769,N_2367,N_674);
nand U4770 (N_4770,N_2420,N_37);
nand U4771 (N_4771,N_1320,N_1220);
xnor U4772 (N_4772,N_1709,N_873);
or U4773 (N_4773,N_1770,N_884);
and U4774 (N_4774,N_2405,N_1853);
xor U4775 (N_4775,N_1391,N_51);
nor U4776 (N_4776,N_9,N_1677);
or U4777 (N_4777,N_289,N_1165);
nor U4778 (N_4778,N_1532,N_1243);
nor U4779 (N_4779,N_1912,N_787);
nand U4780 (N_4780,N_1269,N_896);
nand U4781 (N_4781,N_1629,N_1857);
xnor U4782 (N_4782,N_1756,N_2485);
nand U4783 (N_4783,N_1193,N_681);
nor U4784 (N_4784,N_232,N_1768);
and U4785 (N_4785,N_2197,N_600);
nor U4786 (N_4786,N_2143,N_485);
nor U4787 (N_4787,N_1465,N_538);
xnor U4788 (N_4788,N_2460,N_2301);
xnor U4789 (N_4789,N_1824,N_682);
nand U4790 (N_4790,N_1289,N_2428);
and U4791 (N_4791,N_213,N_1342);
nand U4792 (N_4792,N_1151,N_1241);
or U4793 (N_4793,N_2165,N_118);
or U4794 (N_4794,N_2215,N_551);
nor U4795 (N_4795,N_1220,N_1929);
or U4796 (N_4796,N_210,N_668);
and U4797 (N_4797,N_1425,N_553);
or U4798 (N_4798,N_1660,N_1443);
and U4799 (N_4799,N_1812,N_2198);
nand U4800 (N_4800,N_1162,N_16);
or U4801 (N_4801,N_1226,N_204);
or U4802 (N_4802,N_1802,N_2236);
and U4803 (N_4803,N_386,N_1191);
nor U4804 (N_4804,N_705,N_337);
nor U4805 (N_4805,N_588,N_2072);
xor U4806 (N_4806,N_457,N_822);
and U4807 (N_4807,N_437,N_1345);
nand U4808 (N_4808,N_158,N_171);
xnor U4809 (N_4809,N_425,N_1010);
nand U4810 (N_4810,N_1482,N_489);
and U4811 (N_4811,N_1017,N_160);
and U4812 (N_4812,N_416,N_713);
xnor U4813 (N_4813,N_1890,N_281);
nand U4814 (N_4814,N_2289,N_1417);
xnor U4815 (N_4815,N_506,N_2293);
nand U4816 (N_4816,N_1296,N_2396);
nor U4817 (N_4817,N_184,N_2351);
xnor U4818 (N_4818,N_372,N_1255);
or U4819 (N_4819,N_2012,N_808);
nand U4820 (N_4820,N_681,N_1266);
and U4821 (N_4821,N_1198,N_1057);
nor U4822 (N_4822,N_1411,N_1050);
nor U4823 (N_4823,N_16,N_2498);
xnor U4824 (N_4824,N_1613,N_884);
xnor U4825 (N_4825,N_1235,N_170);
nand U4826 (N_4826,N_122,N_1365);
xnor U4827 (N_4827,N_1566,N_2268);
or U4828 (N_4828,N_27,N_988);
xnor U4829 (N_4829,N_1115,N_1530);
nor U4830 (N_4830,N_742,N_1965);
nor U4831 (N_4831,N_318,N_1490);
xnor U4832 (N_4832,N_1605,N_1943);
xnor U4833 (N_4833,N_1658,N_1557);
xnor U4834 (N_4834,N_1055,N_2120);
and U4835 (N_4835,N_839,N_718);
nor U4836 (N_4836,N_430,N_96);
or U4837 (N_4837,N_145,N_1505);
nor U4838 (N_4838,N_1228,N_2345);
xor U4839 (N_4839,N_1247,N_2413);
or U4840 (N_4840,N_1248,N_1972);
and U4841 (N_4841,N_819,N_153);
nand U4842 (N_4842,N_929,N_1375);
or U4843 (N_4843,N_2469,N_2208);
xor U4844 (N_4844,N_372,N_1396);
and U4845 (N_4845,N_1510,N_1535);
nor U4846 (N_4846,N_1931,N_1268);
xnor U4847 (N_4847,N_2339,N_2117);
and U4848 (N_4848,N_368,N_561);
nor U4849 (N_4849,N_1671,N_198);
or U4850 (N_4850,N_2071,N_51);
and U4851 (N_4851,N_1877,N_1822);
nand U4852 (N_4852,N_1999,N_1722);
nand U4853 (N_4853,N_2019,N_2032);
xor U4854 (N_4854,N_1581,N_1108);
nor U4855 (N_4855,N_1341,N_710);
xor U4856 (N_4856,N_882,N_1424);
or U4857 (N_4857,N_818,N_801);
and U4858 (N_4858,N_1181,N_690);
and U4859 (N_4859,N_277,N_666);
nand U4860 (N_4860,N_868,N_335);
nand U4861 (N_4861,N_1163,N_492);
or U4862 (N_4862,N_2176,N_1934);
nor U4863 (N_4863,N_492,N_709);
xor U4864 (N_4864,N_1749,N_1550);
nand U4865 (N_4865,N_1658,N_314);
and U4866 (N_4866,N_1359,N_1793);
nand U4867 (N_4867,N_1276,N_1960);
or U4868 (N_4868,N_2214,N_212);
nor U4869 (N_4869,N_284,N_2272);
nor U4870 (N_4870,N_179,N_1380);
or U4871 (N_4871,N_1238,N_1039);
and U4872 (N_4872,N_21,N_1252);
nand U4873 (N_4873,N_28,N_1488);
xnor U4874 (N_4874,N_2002,N_1264);
and U4875 (N_4875,N_543,N_235);
nand U4876 (N_4876,N_1742,N_941);
nand U4877 (N_4877,N_825,N_1280);
and U4878 (N_4878,N_402,N_2139);
and U4879 (N_4879,N_657,N_1170);
nor U4880 (N_4880,N_740,N_958);
and U4881 (N_4881,N_832,N_1894);
nor U4882 (N_4882,N_1458,N_977);
nor U4883 (N_4883,N_173,N_2160);
or U4884 (N_4884,N_32,N_1826);
nor U4885 (N_4885,N_979,N_211);
xor U4886 (N_4886,N_328,N_2374);
nand U4887 (N_4887,N_1055,N_795);
or U4888 (N_4888,N_2344,N_444);
and U4889 (N_4889,N_2378,N_1670);
and U4890 (N_4890,N_1428,N_1472);
nor U4891 (N_4891,N_2008,N_2224);
nor U4892 (N_4892,N_1209,N_1788);
or U4893 (N_4893,N_456,N_1733);
and U4894 (N_4894,N_1235,N_2496);
nand U4895 (N_4895,N_2497,N_1426);
nor U4896 (N_4896,N_1099,N_1536);
xnor U4897 (N_4897,N_379,N_74);
or U4898 (N_4898,N_1208,N_569);
and U4899 (N_4899,N_1765,N_1471);
and U4900 (N_4900,N_2072,N_180);
and U4901 (N_4901,N_982,N_1512);
or U4902 (N_4902,N_1341,N_1772);
nor U4903 (N_4903,N_386,N_421);
nand U4904 (N_4904,N_125,N_1603);
nor U4905 (N_4905,N_152,N_1230);
or U4906 (N_4906,N_2288,N_980);
or U4907 (N_4907,N_214,N_1457);
nor U4908 (N_4908,N_300,N_1236);
or U4909 (N_4909,N_919,N_2207);
xor U4910 (N_4910,N_996,N_420);
or U4911 (N_4911,N_1107,N_774);
xnor U4912 (N_4912,N_726,N_1475);
nand U4913 (N_4913,N_181,N_1486);
nor U4914 (N_4914,N_1372,N_1808);
nor U4915 (N_4915,N_1360,N_1981);
nand U4916 (N_4916,N_995,N_335);
xor U4917 (N_4917,N_787,N_2466);
xnor U4918 (N_4918,N_970,N_363);
or U4919 (N_4919,N_1473,N_56);
xor U4920 (N_4920,N_1387,N_2392);
nor U4921 (N_4921,N_1957,N_2314);
xor U4922 (N_4922,N_155,N_1280);
nand U4923 (N_4923,N_1426,N_947);
nor U4924 (N_4924,N_1910,N_145);
or U4925 (N_4925,N_2495,N_1739);
or U4926 (N_4926,N_2484,N_1401);
or U4927 (N_4927,N_1100,N_295);
nand U4928 (N_4928,N_2308,N_624);
and U4929 (N_4929,N_2247,N_1383);
and U4930 (N_4930,N_942,N_56);
nand U4931 (N_4931,N_2139,N_231);
nor U4932 (N_4932,N_1183,N_1033);
nor U4933 (N_4933,N_2065,N_2217);
xnor U4934 (N_4934,N_866,N_2161);
and U4935 (N_4935,N_729,N_1975);
or U4936 (N_4936,N_2046,N_329);
nor U4937 (N_4937,N_720,N_2197);
nand U4938 (N_4938,N_1064,N_2378);
nor U4939 (N_4939,N_1207,N_613);
or U4940 (N_4940,N_585,N_907);
xnor U4941 (N_4941,N_101,N_350);
or U4942 (N_4942,N_807,N_958);
nand U4943 (N_4943,N_601,N_2279);
nor U4944 (N_4944,N_1437,N_463);
nor U4945 (N_4945,N_976,N_1071);
xor U4946 (N_4946,N_905,N_1234);
nand U4947 (N_4947,N_1508,N_271);
or U4948 (N_4948,N_1294,N_262);
nor U4949 (N_4949,N_2180,N_1400);
nand U4950 (N_4950,N_1098,N_2355);
xor U4951 (N_4951,N_227,N_1373);
and U4952 (N_4952,N_833,N_155);
and U4953 (N_4953,N_1959,N_508);
nand U4954 (N_4954,N_1275,N_1248);
xor U4955 (N_4955,N_738,N_1510);
or U4956 (N_4956,N_22,N_2143);
xor U4957 (N_4957,N_1367,N_1797);
nand U4958 (N_4958,N_998,N_1731);
xor U4959 (N_4959,N_889,N_1757);
xnor U4960 (N_4960,N_915,N_2242);
nand U4961 (N_4961,N_1348,N_89);
or U4962 (N_4962,N_918,N_1147);
xor U4963 (N_4963,N_863,N_1276);
or U4964 (N_4964,N_20,N_2349);
nor U4965 (N_4965,N_44,N_1797);
or U4966 (N_4966,N_2351,N_1333);
or U4967 (N_4967,N_1629,N_659);
xnor U4968 (N_4968,N_1520,N_752);
xor U4969 (N_4969,N_1218,N_1164);
nor U4970 (N_4970,N_1236,N_6);
nor U4971 (N_4971,N_2494,N_817);
nor U4972 (N_4972,N_972,N_2410);
xor U4973 (N_4973,N_2108,N_1702);
nor U4974 (N_4974,N_580,N_2014);
nor U4975 (N_4975,N_2257,N_1028);
or U4976 (N_4976,N_445,N_1153);
xnor U4977 (N_4977,N_234,N_1495);
or U4978 (N_4978,N_1740,N_1575);
or U4979 (N_4979,N_264,N_459);
and U4980 (N_4980,N_1803,N_2271);
nor U4981 (N_4981,N_260,N_1194);
xnor U4982 (N_4982,N_393,N_2280);
nor U4983 (N_4983,N_1694,N_294);
and U4984 (N_4984,N_1875,N_705);
nand U4985 (N_4985,N_167,N_788);
xnor U4986 (N_4986,N_328,N_2230);
and U4987 (N_4987,N_1055,N_146);
nor U4988 (N_4988,N_1982,N_2334);
nand U4989 (N_4989,N_1176,N_862);
nand U4990 (N_4990,N_56,N_985);
nor U4991 (N_4991,N_936,N_1904);
nand U4992 (N_4992,N_1832,N_781);
xor U4993 (N_4993,N_2362,N_689);
nor U4994 (N_4994,N_1626,N_943);
or U4995 (N_4995,N_2145,N_1633);
and U4996 (N_4996,N_152,N_1000);
nor U4997 (N_4997,N_880,N_1192);
and U4998 (N_4998,N_936,N_698);
nand U4999 (N_4999,N_1835,N_1396);
or U5000 (N_5000,N_4055,N_4191);
or U5001 (N_5001,N_3489,N_4910);
xor U5002 (N_5002,N_2989,N_4435);
xnor U5003 (N_5003,N_4460,N_3031);
nor U5004 (N_5004,N_2773,N_2797);
nand U5005 (N_5005,N_2829,N_3310);
nand U5006 (N_5006,N_3472,N_4316);
nand U5007 (N_5007,N_3320,N_2738);
xnor U5008 (N_5008,N_4373,N_3191);
xor U5009 (N_5009,N_3155,N_3890);
nand U5010 (N_5010,N_3332,N_3734);
and U5011 (N_5011,N_3801,N_2867);
nand U5012 (N_5012,N_4178,N_3099);
nand U5013 (N_5013,N_4858,N_4992);
and U5014 (N_5014,N_4146,N_4400);
nand U5015 (N_5015,N_3073,N_3604);
or U5016 (N_5016,N_4260,N_4063);
and U5017 (N_5017,N_3770,N_2525);
nand U5018 (N_5018,N_4788,N_2912);
or U5019 (N_5019,N_3828,N_3863);
nand U5020 (N_5020,N_2849,N_4136);
xnor U5021 (N_5021,N_2613,N_2670);
nand U5022 (N_5022,N_4167,N_2999);
and U5023 (N_5023,N_4831,N_2536);
nor U5024 (N_5024,N_4701,N_4439);
or U5025 (N_5025,N_3351,N_4590);
xnor U5026 (N_5026,N_2633,N_3212);
nand U5027 (N_5027,N_3291,N_4344);
or U5028 (N_5028,N_4547,N_3426);
nor U5029 (N_5029,N_4044,N_2991);
xnor U5030 (N_5030,N_4479,N_3660);
nor U5031 (N_5031,N_4397,N_3941);
nor U5032 (N_5032,N_4770,N_2658);
nand U5033 (N_5033,N_3597,N_3199);
and U5034 (N_5034,N_4718,N_4293);
xnor U5035 (N_5035,N_4060,N_4140);
xnor U5036 (N_5036,N_4527,N_2638);
nor U5037 (N_5037,N_4036,N_4698);
nand U5038 (N_5038,N_4394,N_2614);
or U5039 (N_5039,N_4990,N_4923);
nor U5040 (N_5040,N_3123,N_2714);
nand U5041 (N_5041,N_3282,N_2951);
nand U5042 (N_5042,N_3668,N_2655);
and U5043 (N_5043,N_4068,N_4607);
and U5044 (N_5044,N_2676,N_3717);
or U5045 (N_5045,N_2672,N_3701);
nand U5046 (N_5046,N_3072,N_2982);
nor U5047 (N_5047,N_3578,N_4895);
nand U5048 (N_5048,N_4972,N_4970);
nor U5049 (N_5049,N_2767,N_3859);
xnor U5050 (N_5050,N_2842,N_2623);
or U5051 (N_5051,N_3672,N_4314);
and U5052 (N_5052,N_4517,N_4180);
nand U5053 (N_5053,N_4671,N_2504);
nand U5054 (N_5054,N_3030,N_3807);
xnor U5055 (N_5055,N_3362,N_3877);
and U5056 (N_5056,N_4300,N_4742);
xnor U5057 (N_5057,N_4282,N_4752);
and U5058 (N_5058,N_4776,N_3816);
nor U5059 (N_5059,N_4598,N_4372);
and U5060 (N_5060,N_4550,N_2922);
nand U5061 (N_5061,N_4451,N_4796);
nor U5062 (N_5062,N_4716,N_4334);
nor U5063 (N_5063,N_3341,N_4454);
and U5064 (N_5064,N_3224,N_3736);
and U5065 (N_5065,N_4464,N_3560);
nand U5066 (N_5066,N_4892,N_3152);
nor U5067 (N_5067,N_4386,N_2921);
nor U5068 (N_5068,N_2752,N_2503);
or U5069 (N_5069,N_4213,N_3933);
nor U5070 (N_5070,N_2656,N_3068);
or U5071 (N_5071,N_2558,N_2539);
and U5072 (N_5072,N_4336,N_4309);
and U5073 (N_5073,N_4093,N_3994);
and U5074 (N_5074,N_3242,N_2863);
or U5075 (N_5075,N_3886,N_3596);
nand U5076 (N_5076,N_2875,N_2839);
or U5077 (N_5077,N_4872,N_4944);
xnor U5078 (N_5078,N_4906,N_4905);
nand U5079 (N_5079,N_2846,N_2807);
and U5080 (N_5080,N_4769,N_4891);
and U5081 (N_5081,N_3730,N_2641);
or U5082 (N_5082,N_2800,N_2566);
nor U5083 (N_5083,N_2749,N_3891);
nor U5084 (N_5084,N_4071,N_2704);
nor U5085 (N_5085,N_4247,N_4926);
nor U5086 (N_5086,N_3234,N_4047);
or U5087 (N_5087,N_3096,N_2903);
xor U5088 (N_5088,N_4930,N_4982);
nand U5089 (N_5089,N_2682,N_4080);
xnor U5090 (N_5090,N_3461,N_3391);
or U5091 (N_5091,N_4353,N_3448);
and U5092 (N_5092,N_2854,N_4288);
or U5093 (N_5093,N_3616,N_3769);
and U5094 (N_5094,N_2733,N_4586);
xnor U5095 (N_5095,N_3586,N_3685);
xor U5096 (N_5096,N_4898,N_2601);
and U5097 (N_5097,N_3283,N_3095);
nand U5098 (N_5098,N_4131,N_4409);
nand U5099 (N_5099,N_4790,N_4508);
nor U5100 (N_5100,N_2644,N_4363);
and U5101 (N_5101,N_2571,N_4816);
xnor U5102 (N_5102,N_4406,N_2699);
or U5103 (N_5103,N_4122,N_4579);
nor U5104 (N_5104,N_3460,N_4775);
nand U5105 (N_5105,N_4385,N_2684);
or U5106 (N_5106,N_4856,N_3402);
nand U5107 (N_5107,N_3164,N_4161);
and U5108 (N_5108,N_3075,N_2642);
nor U5109 (N_5109,N_3427,N_3343);
or U5110 (N_5110,N_2980,N_3371);
xnor U5111 (N_5111,N_3547,N_3327);
and U5112 (N_5112,N_4472,N_4149);
nand U5113 (N_5113,N_3177,N_4393);
or U5114 (N_5114,N_2883,N_2817);
or U5115 (N_5115,N_3554,N_4367);
or U5116 (N_5116,N_3404,N_3467);
nor U5117 (N_5117,N_2877,N_4268);
and U5118 (N_5118,N_4621,N_3374);
xnor U5119 (N_5119,N_2500,N_3186);
nand U5120 (N_5120,N_3057,N_4578);
nand U5121 (N_5121,N_2998,N_4396);
xnor U5122 (N_5122,N_4021,N_2560);
and U5123 (N_5123,N_2988,N_2565);
or U5124 (N_5124,N_3579,N_2852);
xor U5125 (N_5125,N_4571,N_2774);
xor U5126 (N_5126,N_3087,N_2652);
or U5127 (N_5127,N_4203,N_3696);
nand U5128 (N_5128,N_2981,N_4381);
and U5129 (N_5129,N_3926,N_3934);
nand U5130 (N_5130,N_4274,N_3998);
or U5131 (N_5131,N_3516,N_3936);
or U5132 (N_5132,N_4325,N_3708);
or U5133 (N_5133,N_3179,N_4050);
nor U5134 (N_5134,N_3773,N_2730);
nand U5135 (N_5135,N_4988,N_3421);
xor U5136 (N_5136,N_2803,N_3102);
or U5137 (N_5137,N_4295,N_4227);
or U5138 (N_5138,N_3496,N_4430);
xor U5139 (N_5139,N_4211,N_3814);
xor U5140 (N_5140,N_4675,N_3325);
nor U5141 (N_5141,N_4588,N_2971);
nor U5142 (N_5142,N_4214,N_4876);
nand U5143 (N_5143,N_2758,N_4998);
xnor U5144 (N_5144,N_4807,N_2847);
nor U5145 (N_5145,N_3002,N_2820);
nand U5146 (N_5146,N_3157,N_3272);
nor U5147 (N_5147,N_3248,N_4572);
and U5148 (N_5148,N_4182,N_4552);
nor U5149 (N_5149,N_2516,N_4429);
nor U5150 (N_5150,N_3757,N_4436);
or U5151 (N_5151,N_3085,N_3832);
nand U5152 (N_5152,N_3630,N_4190);
xor U5153 (N_5153,N_2794,N_4916);
and U5154 (N_5154,N_3469,N_3942);
and U5155 (N_5155,N_4101,N_4835);
or U5156 (N_5156,N_4783,N_4737);
nor U5157 (N_5157,N_3409,N_2519);
and U5158 (N_5158,N_3714,N_4426);
nor U5159 (N_5159,N_2943,N_3084);
or U5160 (N_5160,N_4407,N_4064);
or U5161 (N_5161,N_3023,N_3308);
nor U5162 (N_5162,N_3670,N_3928);
or U5163 (N_5163,N_4541,N_4584);
nand U5164 (N_5164,N_3275,N_4967);
nand U5165 (N_5165,N_3722,N_2799);
xnor U5166 (N_5166,N_4948,N_3357);
and U5167 (N_5167,N_2972,N_4975);
or U5168 (N_5168,N_3870,N_4069);
nand U5169 (N_5169,N_4627,N_3788);
nand U5170 (N_5170,N_4756,N_2635);
nand U5171 (N_5171,N_3278,N_3497);
nand U5172 (N_5172,N_4630,N_4315);
nand U5173 (N_5173,N_2984,N_4357);
and U5174 (N_5174,N_2535,N_2890);
xor U5175 (N_5175,N_4270,N_4431);
nand U5176 (N_5176,N_3008,N_4803);
nand U5177 (N_5177,N_4734,N_3463);
or U5178 (N_5178,N_2961,N_4567);
and U5179 (N_5179,N_2569,N_4777);
nor U5180 (N_5180,N_3988,N_3216);
or U5181 (N_5181,N_3262,N_3546);
and U5182 (N_5182,N_3603,N_3168);
nor U5183 (N_5183,N_4039,N_3778);
or U5184 (N_5184,N_2592,N_2743);
nor U5185 (N_5185,N_4951,N_3522);
nor U5186 (N_5186,N_3055,N_4465);
xor U5187 (N_5187,N_4506,N_2994);
nand U5188 (N_5188,N_4204,N_2750);
and U5189 (N_5189,N_3957,N_4434);
nand U5190 (N_5190,N_4414,N_4925);
nand U5191 (N_5191,N_3313,N_4907);
or U5192 (N_5192,N_4001,N_3836);
nand U5193 (N_5193,N_3798,N_4185);
nand U5194 (N_5194,N_3440,N_3297);
nor U5195 (N_5195,N_4338,N_4448);
nand U5196 (N_5196,N_2593,N_4249);
nand U5197 (N_5197,N_4020,N_3160);
xor U5198 (N_5198,N_2748,N_3751);
nand U5199 (N_5199,N_2792,N_4450);
or U5200 (N_5200,N_2995,N_3260);
and U5201 (N_5201,N_4751,N_3299);
xnor U5202 (N_5202,N_3004,N_3150);
nand U5203 (N_5203,N_3366,N_3447);
nor U5204 (N_5204,N_4619,N_3114);
nand U5205 (N_5205,N_3764,N_4401);
and U5206 (N_5206,N_4674,N_3611);
xnor U5207 (N_5207,N_2705,N_3478);
or U5208 (N_5208,N_2555,N_3290);
nor U5209 (N_5209,N_3569,N_3585);
nand U5210 (N_5210,N_3333,N_4974);
xor U5211 (N_5211,N_4613,N_2896);
nand U5212 (N_5212,N_3386,N_3678);
nand U5213 (N_5213,N_3052,N_4291);
or U5214 (N_5214,N_4244,N_4484);
or U5215 (N_5215,N_3720,N_3459);
nor U5216 (N_5216,N_2722,N_4252);
xnor U5217 (N_5217,N_2657,N_3881);
nor U5218 (N_5218,N_4921,N_4124);
nand U5219 (N_5219,N_2606,N_2956);
xor U5220 (N_5220,N_4085,N_3698);
or U5221 (N_5221,N_2531,N_3382);
and U5222 (N_5222,N_3927,N_4786);
or U5223 (N_5223,N_4943,N_3767);
or U5224 (N_5224,N_3132,N_3515);
nor U5225 (N_5225,N_3491,N_2802);
nand U5226 (N_5226,N_4509,N_4861);
and U5227 (N_5227,N_3935,N_2939);
or U5228 (N_5228,N_3744,N_4228);
nor U5229 (N_5229,N_2880,N_4838);
and U5230 (N_5230,N_4684,N_3873);
nand U5231 (N_5231,N_4649,N_2919);
or U5232 (N_5232,N_2729,N_2851);
xor U5233 (N_5233,N_3951,N_2583);
nor U5234 (N_5234,N_3705,N_4323);
and U5235 (N_5235,N_3026,N_4886);
and U5236 (N_5236,N_3316,N_3652);
nand U5237 (N_5237,N_3692,N_4792);
and U5238 (N_5238,N_4466,N_4486);
and U5239 (N_5239,N_3917,N_2709);
and U5240 (N_5240,N_3434,N_3221);
xnor U5241 (N_5241,N_3561,N_4714);
xnor U5242 (N_5242,N_4241,N_3484);
nor U5243 (N_5243,N_3388,N_4004);
xnor U5244 (N_5244,N_3317,N_2879);
nand U5245 (N_5245,N_4117,N_4947);
nor U5246 (N_5246,N_4965,N_3563);
and U5247 (N_5247,N_3488,N_2791);
nand U5248 (N_5248,N_2731,N_2804);
nand U5249 (N_5249,N_2881,N_4958);
xor U5250 (N_5250,N_4404,N_4804);
nand U5251 (N_5251,N_2837,N_3745);
nand U5252 (N_5252,N_2823,N_4232);
nand U5253 (N_5253,N_2955,N_4853);
nand U5254 (N_5254,N_3479,N_4492);
and U5255 (N_5255,N_4519,N_4938);
and U5256 (N_5256,N_2764,N_4868);
nand U5257 (N_5257,N_4841,N_3449);
nor U5258 (N_5258,N_4797,N_4881);
nor U5259 (N_5259,N_2910,N_3194);
nand U5260 (N_5260,N_4153,N_4410);
nor U5261 (N_5261,N_3575,N_4257);
nor U5262 (N_5262,N_4801,N_3509);
and U5263 (N_5263,N_4529,N_4667);
nand U5264 (N_5264,N_4016,N_3700);
or U5265 (N_5265,N_2987,N_4896);
or U5266 (N_5266,N_4639,N_4349);
and U5267 (N_5267,N_2680,N_2685);
nor U5268 (N_5268,N_3746,N_3158);
nand U5269 (N_5269,N_3978,N_4570);
or U5270 (N_5270,N_4577,N_2702);
or U5271 (N_5271,N_3664,N_4894);
nor U5272 (N_5272,N_2825,N_3043);
nand U5273 (N_5273,N_4904,N_4711);
and U5274 (N_5274,N_4462,N_2781);
or U5275 (N_5275,N_2600,N_3804);
xor U5276 (N_5276,N_3053,N_2882);
or U5277 (N_5277,N_2806,N_3949);
or U5278 (N_5278,N_4311,N_2788);
nor U5279 (N_5279,N_4278,N_2537);
or U5280 (N_5280,N_4163,N_4764);
nor U5281 (N_5281,N_3127,N_2591);
nor U5282 (N_5282,N_4605,N_2515);
nand U5283 (N_5283,N_4638,N_3711);
nand U5284 (N_5284,N_4864,N_3028);
and U5285 (N_5285,N_3851,N_2885);
nand U5286 (N_5286,N_3422,N_3955);
nor U5287 (N_5287,N_3056,N_4237);
or U5288 (N_5288,N_4280,N_2717);
and U5289 (N_5289,N_2665,N_2900);
nand U5290 (N_5290,N_4545,N_2628);
or U5291 (N_5291,N_3962,N_3149);
nand U5292 (N_5292,N_3372,N_3480);
xnor U5293 (N_5293,N_4978,N_3618);
nor U5294 (N_5294,N_3334,N_4507);
or U5295 (N_5295,N_2771,N_4743);
and U5296 (N_5296,N_3166,N_3898);
and U5297 (N_5297,N_3347,N_3116);
nor U5298 (N_5298,N_3286,N_3187);
nand U5299 (N_5299,N_4903,N_2857);
and U5300 (N_5300,N_2726,N_4745);
nor U5301 (N_5301,N_3661,N_3256);
or U5302 (N_5302,N_3277,N_2718);
nor U5303 (N_5303,N_4837,N_4231);
xor U5304 (N_5304,N_2514,N_3694);
and U5305 (N_5305,N_3328,N_4172);
and U5306 (N_5306,N_3727,N_3458);
nand U5307 (N_5307,N_4310,N_3601);
nand U5308 (N_5308,N_4780,N_3889);
nor U5309 (N_5309,N_3531,N_4986);
nor U5310 (N_5310,N_3502,N_2521);
xnor U5311 (N_5311,N_2858,N_3133);
and U5312 (N_5312,N_4164,N_2732);
nand U5313 (N_5313,N_3580,N_4233);
nor U5314 (N_5314,N_2831,N_3592);
nor U5315 (N_5315,N_4806,N_4676);
and U5316 (N_5316,N_2697,N_3355);
and U5317 (N_5317,N_3475,N_4901);
nor U5318 (N_5318,N_4973,N_3445);
xnor U5319 (N_5319,N_3182,N_4361);
xor U5320 (N_5320,N_4432,N_2627);
nor U5321 (N_5321,N_3444,N_4695);
nor U5322 (N_5322,N_3946,N_4289);
nand U5323 (N_5323,N_3573,N_4932);
nand U5324 (N_5324,N_4284,N_3633);
xor U5325 (N_5325,N_3017,N_2549);
nor U5326 (N_5326,N_3198,N_2878);
or U5327 (N_5327,N_3035,N_3691);
nand U5328 (N_5328,N_4443,N_2992);
or U5329 (N_5329,N_4006,N_4489);
nor U5330 (N_5330,N_4785,N_3874);
or U5331 (N_5331,N_4113,N_3925);
xnor U5332 (N_5332,N_4319,N_4771);
nand U5333 (N_5333,N_4165,N_3724);
nand U5334 (N_5334,N_4893,N_2666);
nor U5335 (N_5335,N_4834,N_3178);
nand U5336 (N_5336,N_4819,N_3987);
nor U5337 (N_5337,N_3039,N_4035);
and U5338 (N_5338,N_3864,N_3803);
nand U5339 (N_5339,N_4915,N_3003);
nor U5340 (N_5340,N_3113,N_4647);
nor U5341 (N_5341,N_4285,N_4616);
or U5342 (N_5342,N_4350,N_4503);
nor U5343 (N_5343,N_4618,N_4246);
nor U5344 (N_5344,N_3315,N_3209);
nor U5345 (N_5345,N_2827,N_2946);
and U5346 (N_5346,N_2808,N_4437);
and U5347 (N_5347,N_4902,N_3014);
nor U5348 (N_5348,N_4042,N_4345);
and U5349 (N_5349,N_4679,N_4713);
nand U5350 (N_5350,N_3094,N_3457);
or U5351 (N_5351,N_4840,N_4920);
and U5352 (N_5352,N_3074,N_3012);
xor U5353 (N_5353,N_4263,N_4582);
xor U5354 (N_5354,N_4624,N_4481);
nor U5355 (N_5355,N_4909,N_4245);
nor U5356 (N_5356,N_3654,N_2643);
and U5357 (N_5357,N_4480,N_4427);
and U5358 (N_5358,N_4087,N_3368);
nand U5359 (N_5359,N_3681,N_3914);
or U5360 (N_5360,N_4761,N_3674);
nand U5361 (N_5361,N_3818,N_2511);
and U5362 (N_5362,N_2734,N_4885);
xnor U5363 (N_5363,N_3011,N_4599);
or U5364 (N_5364,N_4558,N_2720);
or U5365 (N_5365,N_3302,N_4302);
xor U5366 (N_5366,N_4748,N_2548);
nor U5367 (N_5367,N_4625,N_3270);
xor U5368 (N_5368,N_4542,N_4936);
and U5369 (N_5369,N_2577,N_3019);
or U5370 (N_5370,N_4176,N_4534);
and U5371 (N_5371,N_3274,N_3703);
xnor U5372 (N_5372,N_2559,N_4854);
and U5373 (N_5373,N_2612,N_2715);
and U5374 (N_5374,N_3184,N_2969);
and U5375 (N_5375,N_4195,N_2621);
nand U5376 (N_5376,N_2891,N_4694);
nor U5377 (N_5377,N_4942,N_3916);
nand U5378 (N_5378,N_3101,N_4878);
xor U5379 (N_5379,N_4828,N_3909);
nand U5380 (N_5380,N_3806,N_3977);
nor U5381 (N_5381,N_3837,N_3206);
and U5382 (N_5382,N_2901,N_2864);
or U5383 (N_5383,N_3380,N_3415);
nand U5384 (N_5384,N_3849,N_2966);
nor U5385 (N_5385,N_4095,N_4850);
and U5386 (N_5386,N_2974,N_3662);
and U5387 (N_5387,N_4557,N_3229);
nor U5388 (N_5388,N_3431,N_3367);
xnor U5389 (N_5389,N_3675,N_3862);
nand U5390 (N_5390,N_2605,N_2540);
xnor U5391 (N_5391,N_3439,N_4849);
or U5392 (N_5392,N_3776,N_4056);
nor U5393 (N_5393,N_3495,N_3059);
nor U5394 (N_5394,N_2907,N_2742);
nand U5395 (N_5395,N_2532,N_3524);
nor U5396 (N_5396,N_3839,N_4715);
and U5397 (N_5397,N_4415,N_3846);
nor U5398 (N_5398,N_3303,N_3944);
or U5399 (N_5399,N_3841,N_3128);
or U5400 (N_5400,N_3385,N_2761);
xnor U5401 (N_5401,N_3600,N_4335);
nand U5402 (N_5402,N_2664,N_3456);
nand U5403 (N_5403,N_3240,N_4660);
nor U5404 (N_5404,N_2787,N_4145);
or U5405 (N_5405,N_3226,N_4461);
nor U5406 (N_5406,N_4238,N_3840);
nand U5407 (N_5407,N_3474,N_4591);
xnor U5408 (N_5408,N_2712,N_4495);
nor U5409 (N_5409,N_3397,N_4908);
nor U5410 (N_5410,N_4683,N_4762);
nor U5411 (N_5411,N_2942,N_4672);
nor U5412 (N_5412,N_4049,N_3103);
nor U5413 (N_5413,N_3399,N_2597);
xor U5414 (N_5414,N_4815,N_3289);
or U5415 (N_5415,N_3759,N_4077);
xor U5416 (N_5416,N_4691,N_4287);
xor U5417 (N_5417,N_4078,N_3477);
xor U5418 (N_5418,N_4096,N_4147);
nor U5419 (N_5419,N_4387,N_4626);
xnor U5420 (N_5420,N_2609,N_4569);
or U5421 (N_5421,N_2648,N_4061);
nand U5422 (N_5422,N_4248,N_4845);
nand U5423 (N_5423,N_2816,N_3970);
xor U5424 (N_5424,N_3301,N_2790);
xnor U5425 (N_5425,N_3353,N_3823);
nand U5426 (N_5426,N_3518,N_3381);
and U5427 (N_5427,N_4979,N_4433);
nor U5428 (N_5428,N_2745,N_3659);
or U5429 (N_5429,N_4193,N_3610);
nor U5430 (N_5430,N_2967,N_3716);
and U5431 (N_5431,N_3799,N_3843);
nor U5432 (N_5432,N_4076,N_2945);
and U5433 (N_5433,N_3067,N_3507);
nor U5434 (N_5434,N_2868,N_4470);
xnor U5435 (N_5435,N_3490,N_3911);
nand U5436 (N_5436,N_4987,N_3238);
xnor U5437 (N_5437,N_4239,N_3822);
nand U5438 (N_5438,N_2746,N_4086);
nand U5439 (N_5439,N_3393,N_4208);
nand U5440 (N_5440,N_4888,N_3631);
nand U5441 (N_5441,N_4833,N_3728);
and U5442 (N_5442,N_3394,N_3305);
nor U5443 (N_5443,N_4262,N_4912);
xor U5444 (N_5444,N_3510,N_4732);
nand U5445 (N_5445,N_3151,N_4928);
nor U5446 (N_5446,N_3271,N_4601);
nand U5447 (N_5447,N_4202,N_4121);
and U5448 (N_5448,N_3860,N_2626);
nand U5449 (N_5449,N_4360,N_4189);
nand U5450 (N_5450,N_4216,N_4829);
and U5451 (N_5451,N_4298,N_3188);
nand U5452 (N_5452,N_4286,N_3855);
xnor U5453 (N_5453,N_3342,N_2833);
nand U5454 (N_5454,N_3958,N_4469);
or U5455 (N_5455,N_3782,N_3642);
xnor U5456 (N_5456,N_3687,N_3765);
and U5457 (N_5457,N_4041,N_4995);
or U5458 (N_5458,N_4155,N_4874);
xor U5459 (N_5459,N_4900,N_4559);
nor U5460 (N_5460,N_3774,N_2985);
or U5461 (N_5461,N_3693,N_3587);
nand U5462 (N_5462,N_3538,N_4817);
and U5463 (N_5463,N_4179,N_3145);
xnor U5464 (N_5464,N_3257,N_3192);
or U5465 (N_5465,N_3626,N_3219);
or U5466 (N_5466,N_3591,N_3755);
xnor U5467 (N_5467,N_4941,N_4418);
nor U5468 (N_5468,N_4610,N_3710);
nor U5469 (N_5469,N_4159,N_3280);
xnor U5470 (N_5470,N_4617,N_4151);
or U5471 (N_5471,N_4802,N_3779);
xor U5472 (N_5472,N_4120,N_3365);
xor U5473 (N_5473,N_2893,N_3910);
nand U5474 (N_5474,N_3329,N_4370);
or U5475 (N_5475,N_3247,N_4824);
or U5476 (N_5476,N_2568,N_4961);
and U5477 (N_5477,N_3293,N_3231);
nor U5478 (N_5478,N_2646,N_2810);
nor U5479 (N_5479,N_4346,N_3953);
xor U5480 (N_5480,N_4632,N_4725);
or U5481 (N_5481,N_4391,N_3134);
and U5482 (N_5482,N_4953,N_2843);
xor U5483 (N_5483,N_2552,N_3009);
and U5484 (N_5484,N_3689,N_4499);
and U5485 (N_5485,N_3433,N_3125);
nor U5486 (N_5486,N_2584,N_3852);
or U5487 (N_5487,N_3140,N_4482);
or U5488 (N_5488,N_4264,N_4494);
nand U5489 (N_5489,N_3220,N_2551);
or U5490 (N_5490,N_2929,N_3967);
nand U5491 (N_5491,N_3867,N_2894);
nor U5492 (N_5492,N_3702,N_4911);
xor U5493 (N_5493,N_4075,N_3752);
and U5494 (N_5494,N_2735,N_4065);
xor U5495 (N_5495,N_3679,N_3665);
and U5496 (N_5496,N_3676,N_3786);
nor U5497 (N_5497,N_2869,N_3153);
nand U5498 (N_5498,N_4668,N_2904);
or U5499 (N_5499,N_4651,N_3838);
xnor U5500 (N_5500,N_4100,N_2990);
xnor U5501 (N_5501,N_3135,N_4197);
or U5502 (N_5502,N_4132,N_3793);
xnor U5503 (N_5503,N_2975,N_2688);
or U5504 (N_5504,N_4791,N_4997);
nand U5505 (N_5505,N_4051,N_2824);
or U5506 (N_5506,N_3078,N_3241);
xor U5507 (N_5507,N_4846,N_2836);
or U5508 (N_5508,N_3339,N_4883);
nor U5509 (N_5509,N_4091,N_4511);
and U5510 (N_5510,N_3468,N_4554);
xnor U5511 (N_5511,N_3943,N_3655);
nor U5512 (N_5512,N_2622,N_4747);
xor U5513 (N_5513,N_2917,N_2741);
and U5514 (N_5514,N_3647,N_4689);
nor U5515 (N_5515,N_3628,N_3139);
nand U5516 (N_5516,N_3945,N_4983);
xnor U5517 (N_5517,N_2844,N_4186);
or U5518 (N_5518,N_4899,N_4832);
xnor U5519 (N_5519,N_4304,N_3753);
and U5520 (N_5520,N_3537,N_4646);
nand U5521 (N_5521,N_3016,N_3922);
nand U5522 (N_5522,N_2724,N_3820);
nor U5523 (N_5523,N_3425,N_4536);
and U5524 (N_5524,N_3718,N_2865);
and U5525 (N_5525,N_3737,N_3285);
and U5526 (N_5526,N_4991,N_4730);
nand U5527 (N_5527,N_4692,N_2862);
nor U5528 (N_5528,N_4157,N_4798);
xnor U5529 (N_5529,N_2651,N_4820);
nand U5530 (N_5530,N_3775,N_3006);
nor U5531 (N_5531,N_4533,N_2509);
or U5532 (N_5532,N_2703,N_2747);
or U5533 (N_5533,N_3193,N_3549);
and U5534 (N_5534,N_3331,N_4099);
nand U5535 (N_5535,N_3632,N_3264);
or U5536 (N_5536,N_3536,N_3713);
nand U5537 (N_5537,N_4512,N_4267);
or U5538 (N_5538,N_4158,N_2895);
xor U5539 (N_5539,N_4518,N_2629);
and U5540 (N_5540,N_4420,N_3956);
nand U5541 (N_5541,N_3966,N_2780);
and U5542 (N_5542,N_3097,N_2822);
nor U5543 (N_5543,N_3930,N_2779);
and U5544 (N_5544,N_4666,N_4556);
nor U5545 (N_5545,N_4389,N_3483);
nand U5546 (N_5546,N_4028,N_3784);
nand U5547 (N_5547,N_2898,N_4793);
nor U5548 (N_5548,N_2782,N_3845);
nand U5549 (N_5549,N_4709,N_4971);
and U5550 (N_5550,N_4474,N_3739);
and U5551 (N_5551,N_3252,N_2654);
nand U5552 (N_5552,N_2667,N_3412);
or U5553 (N_5553,N_3237,N_2693);
xnor U5554 (N_5554,N_2700,N_2830);
nor U5555 (N_5555,N_3120,N_3871);
or U5556 (N_5556,N_4359,N_4890);
and U5557 (N_5557,N_3454,N_3041);
nand U5558 (N_5558,N_3999,N_4364);
and U5559 (N_5559,N_3232,N_2866);
and U5560 (N_5560,N_2660,N_3663);
xor U5561 (N_5561,N_4581,N_4879);
or U5562 (N_5562,N_3947,N_2826);
nand U5563 (N_5563,N_4989,N_2813);
xnor U5564 (N_5564,N_4171,N_4813);
and U5565 (N_5565,N_2772,N_3373);
nand U5566 (N_5566,N_2708,N_3932);
nor U5567 (N_5567,N_2534,N_3584);
or U5568 (N_5568,N_4369,N_3356);
nand U5569 (N_5569,N_2501,N_4177);
or U5570 (N_5570,N_3124,N_3980);
xnor U5571 (N_5571,N_3529,N_4636);
xor U5572 (N_5572,N_3562,N_3344);
nand U5573 (N_5573,N_4867,N_2953);
and U5574 (N_5574,N_4693,N_4956);
or U5575 (N_5575,N_3599,N_4059);
xor U5576 (N_5576,N_4889,N_2793);
or U5577 (N_5577,N_2959,N_3527);
nand U5578 (N_5578,N_3204,N_3697);
xor U5579 (N_5579,N_4825,N_4946);
nor U5580 (N_5580,N_3138,N_4219);
nand U5581 (N_5581,N_3117,N_3887);
nor U5582 (N_5582,N_3077,N_4648);
and U5583 (N_5583,N_3062,N_3589);
xor U5584 (N_5584,N_4468,N_4229);
or U5585 (N_5585,N_4768,N_3858);
and U5586 (N_5586,N_3519,N_3222);
nand U5587 (N_5587,N_3406,N_4875);
nor U5588 (N_5588,N_2909,N_2637);
nor U5589 (N_5589,N_2923,N_4321);
or U5590 (N_5590,N_2986,N_3583);
and U5591 (N_5591,N_2711,N_4478);
xor U5592 (N_5592,N_3666,N_3423);
nor U5593 (N_5593,N_3805,N_4521);
nor U5594 (N_5594,N_2529,N_2850);
nand U5595 (N_5595,N_4614,N_3992);
nor U5596 (N_5596,N_2860,N_3107);
and U5597 (N_5597,N_2544,N_3005);
nor U5598 (N_5598,N_4859,N_3273);
xnor U5599 (N_5599,N_2542,N_2587);
nand U5600 (N_5600,N_2550,N_4968);
xor U5601 (N_5601,N_3088,N_2589);
or U5602 (N_5602,N_4993,N_2798);
and U5603 (N_5603,N_4013,N_4269);
and U5604 (N_5604,N_2751,N_2595);
and U5605 (N_5605,N_2763,N_4757);
nand U5606 (N_5606,N_3025,N_3122);
nor U5607 (N_5607,N_3080,N_2968);
and U5608 (N_5608,N_2562,N_3492);
xor U5609 (N_5609,N_2706,N_2567);
nor U5610 (N_5610,N_4573,N_4150);
and U5611 (N_5611,N_3990,N_4568);
nor U5612 (N_5612,N_4329,N_4224);
or U5613 (N_5613,N_3338,N_2815);
nand U5614 (N_5614,N_3712,N_3740);
and U5615 (N_5615,N_4629,N_2777);
nor U5616 (N_5616,N_3109,N_4724);
nor U5617 (N_5617,N_4955,N_3438);
and U5618 (N_5618,N_3539,N_3211);
xnor U5619 (N_5619,N_4810,N_4438);
or U5620 (N_5620,N_4072,N_3130);
or U5621 (N_5621,N_3621,N_3392);
nand U5622 (N_5622,N_3236,N_3500);
xnor U5623 (N_5623,N_4594,N_4773);
and U5624 (N_5624,N_4812,N_3403);
xnor U5625 (N_5625,N_4640,N_2546);
and U5626 (N_5626,N_3559,N_3446);
xor U5627 (N_5627,N_4729,N_3263);
and U5628 (N_5628,N_3215,N_4272);
xnor U5629 (N_5629,N_3643,N_3471);
and U5630 (N_5630,N_4116,N_3535);
xor U5631 (N_5631,N_2934,N_2675);
xor U5632 (N_5632,N_3255,N_3170);
and U5633 (N_5633,N_4187,N_3210);
nand U5634 (N_5634,N_3481,N_2821);
nor U5635 (N_5635,N_2778,N_2828);
and U5636 (N_5636,N_3856,N_4175);
or U5637 (N_5637,N_4183,N_4827);
nor U5638 (N_5638,N_2845,N_4753);
and U5639 (N_5639,N_4653,N_3108);
nand U5640 (N_5640,N_4976,N_3817);
xnor U5641 (N_5641,N_3985,N_4657);
xnor U5642 (N_5642,N_3369,N_3743);
xor U5643 (N_5643,N_4682,N_3214);
xnor U5644 (N_5644,N_2937,N_4294);
nand U5645 (N_5645,N_4645,N_4862);
nand U5646 (N_5646,N_2818,N_2809);
xnor U5647 (N_5647,N_3815,N_3564);
and U5648 (N_5648,N_3868,N_2617);
nor U5649 (N_5649,N_3809,N_2561);
or U5650 (N_5650,N_2812,N_3246);
and U5651 (N_5651,N_4070,N_3395);
or U5652 (N_5652,N_3045,N_4148);
nor U5653 (N_5653,N_3148,N_3424);
nor U5654 (N_5654,N_4778,N_3390);
nand U5655 (N_5655,N_3854,N_3079);
nor U5656 (N_5656,N_3861,N_4243);
xnor U5657 (N_5657,N_4421,N_4048);
or U5658 (N_5658,N_4317,N_3185);
and U5659 (N_5659,N_2756,N_4090);
nand U5660 (N_5660,N_4741,N_4408);
nor U5661 (N_5661,N_2768,N_3629);
and U5662 (N_5662,N_3119,N_3882);
nand U5663 (N_5663,N_2938,N_3842);
nand U5664 (N_5664,N_4412,N_2970);
or U5665 (N_5665,N_4440,N_4697);
and U5666 (N_5666,N_3007,N_4760);
nor U5667 (N_5667,N_4548,N_4027);
nor U5668 (N_5668,N_4331,N_3251);
nand U5669 (N_5669,N_3964,N_3173);
nand U5670 (N_5670,N_4937,N_4996);
nand U5671 (N_5671,N_2888,N_3878);
nand U5672 (N_5672,N_4253,N_2727);
nand U5673 (N_5673,N_2636,N_3646);
nand U5674 (N_5674,N_4608,N_3022);
or U5675 (N_5675,N_4222,N_2578);
or U5676 (N_5676,N_2625,N_3401);
xnor U5677 (N_5677,N_3590,N_2572);
or U5678 (N_5678,N_2775,N_3254);
nor U5679 (N_5679,N_4207,N_3027);
and U5680 (N_5680,N_2710,N_3893);
and U5681 (N_5681,N_4144,N_4209);
and U5682 (N_5682,N_4330,N_4623);
nand U5683 (N_5683,N_4656,N_3337);
and U5684 (N_5684,N_4098,N_4458);
nand U5685 (N_5685,N_3189,N_4818);
and U5686 (N_5686,N_4563,N_4375);
nor U5687 (N_5687,N_3810,N_4597);
xnor U5688 (N_5688,N_2608,N_3276);
or U5689 (N_5689,N_3482,N_3742);
xor U5690 (N_5690,N_2526,N_3938);
xnor U5691 (N_5691,N_3081,N_4054);
xnor U5692 (N_5692,N_4115,N_3090);
nor U5693 (N_5693,N_2543,N_3295);
nor U5694 (N_5694,N_4215,N_3976);
nor U5695 (N_5695,N_4513,N_4669);
nand U5696 (N_5696,N_2962,N_3112);
nor U5697 (N_5697,N_3307,N_4731);
nand U5698 (N_5698,N_4673,N_3499);
xor U5699 (N_5699,N_4585,N_4067);
nand U5700 (N_5700,N_3892,N_3682);
or U5701 (N_5701,N_2785,N_4690);
and U5702 (N_5702,N_3615,N_2884);
and U5703 (N_5703,N_2997,N_3533);
or U5704 (N_5704,N_3551,N_3069);
nor U5705 (N_5705,N_4014,N_3322);
and U5706 (N_5706,N_3975,N_3915);
nand U5707 (N_5707,N_4152,N_3635);
nor U5708 (N_5708,N_4073,N_3258);
and U5709 (N_5709,N_4107,N_3576);
nand U5710 (N_5710,N_4281,N_4583);
xnor U5711 (N_5711,N_3648,N_3378);
nand U5712 (N_5712,N_4168,N_3800);
or U5713 (N_5713,N_3826,N_3010);
xor U5714 (N_5714,N_3568,N_2683);
or U5715 (N_5715,N_4746,N_4772);
and U5716 (N_5716,N_2873,N_3176);
nand U5717 (N_5717,N_4303,N_4024);
or U5718 (N_5718,N_4687,N_3673);
or U5719 (N_5719,N_2795,N_2686);
xnor U5720 (N_5720,N_4650,N_2585);
and U5721 (N_5721,N_2570,N_3831);
or U5722 (N_5722,N_3418,N_4799);
or U5723 (N_5723,N_3544,N_4327);
and U5724 (N_5724,N_4154,N_3669);
nor U5725 (N_5725,N_4954,N_3619);
xnor U5726 (N_5726,N_4576,N_4685);
or U5727 (N_5727,N_2957,N_4296);
or U5728 (N_5728,N_4395,N_4089);
nand U5729 (N_5729,N_3645,N_2530);
and U5730 (N_5730,N_3105,N_4417);
nand U5731 (N_5731,N_3924,N_2759);
nand U5732 (N_5732,N_4143,N_4789);
nand U5733 (N_5733,N_4952,N_4516);
nand U5734 (N_5734,N_2721,N_4251);
nand U5735 (N_5735,N_4220,N_3653);
nor U5736 (N_5736,N_3617,N_4062);
nand U5737 (N_5737,N_4445,N_2649);
and U5738 (N_5738,N_4723,N_4538);
xnor U5739 (N_5739,N_4927,N_3634);
xor U5740 (N_5740,N_4455,N_4104);
nand U5741 (N_5741,N_4037,N_3314);
nor U5742 (N_5742,N_4471,N_3345);
nand U5743 (N_5743,N_4739,N_4960);
and U5744 (N_5744,N_3143,N_4265);
xor U5745 (N_5745,N_3897,N_2596);
xor U5746 (N_5746,N_4324,N_4081);
nor U5747 (N_5747,N_3000,N_3950);
nor U5748 (N_5748,N_3443,N_3118);
and U5749 (N_5749,N_4088,N_4704);
nand U5750 (N_5750,N_3121,N_3208);
xnor U5751 (N_5751,N_3487,N_3265);
xnor U5752 (N_5752,N_4949,N_4306);
and U5753 (N_5753,N_3046,N_4959);
xor U5754 (N_5754,N_2573,N_3044);
nand U5755 (N_5755,N_3726,N_4416);
and U5756 (N_5756,N_3638,N_4749);
nand U5757 (N_5757,N_3350,N_2739);
nand U5758 (N_5758,N_3233,N_4212);
nor U5759 (N_5759,N_2933,N_3594);
nor U5760 (N_5760,N_4663,N_3644);
or U5761 (N_5761,N_3811,N_2650);
nand U5762 (N_5762,N_4863,N_3605);
and U5763 (N_5763,N_3570,N_2647);
xnor U5764 (N_5764,N_4196,N_3572);
or U5765 (N_5765,N_3725,N_3723);
or U5766 (N_5766,N_4774,N_3508);
nand U5767 (N_5767,N_2872,N_3699);
and U5768 (N_5768,N_3606,N_3971);
or U5769 (N_5769,N_4539,N_3249);
and U5770 (N_5770,N_3354,N_4275);
or U5771 (N_5771,N_2563,N_2590);
xnor U5772 (N_5772,N_3250,N_3131);
or U5773 (N_5773,N_3142,N_4223);
nor U5774 (N_5774,N_4382,N_4917);
xnor U5775 (N_5775,N_4322,N_4531);
or U5776 (N_5776,N_3311,N_2716);
nor U5777 (N_5777,N_2978,N_4194);
or U5778 (N_5778,N_3268,N_3181);
xor U5779 (N_5779,N_2575,N_2805);
nor U5780 (N_5780,N_3651,N_3530);
xnor U5781 (N_5781,N_4950,N_2668);
and U5782 (N_5782,N_3671,N_3464);
or U5783 (N_5783,N_3335,N_3895);
or U5784 (N_5784,N_3542,N_2925);
nor U5785 (N_5785,N_4514,N_4504);
xnor U5786 (N_5786,N_3989,N_3034);
and U5787 (N_5787,N_3906,N_3485);
nand U5788 (N_5788,N_2848,N_3253);
and U5789 (N_5789,N_3894,N_4301);
nor U5790 (N_5790,N_2915,N_4009);
xnor U5791 (N_5791,N_4842,N_2930);
xnor U5792 (N_5792,N_4299,N_2553);
or U5793 (N_5793,N_4611,N_2517);
xnor U5794 (N_5794,N_4622,N_2838);
nor U5795 (N_5795,N_2602,N_4276);
nor U5796 (N_5796,N_3396,N_2973);
and U5797 (N_5797,N_4188,N_4358);
nand U5798 (N_5798,N_4596,N_2958);
or U5799 (N_5799,N_3995,N_4717);
or U5800 (N_5800,N_3389,N_3921);
nand U5801 (N_5801,N_3162,N_4053);
nor U5802 (N_5802,N_3190,N_4017);
xor U5803 (N_5803,N_2728,N_3450);
nand U5804 (N_5804,N_4112,N_4273);
or U5805 (N_5805,N_3318,N_4643);
or U5806 (N_5806,N_3639,N_3419);
or U5807 (N_5807,N_4722,N_4852);
and U5808 (N_5808,N_3306,N_3526);
xnor U5809 (N_5809,N_3292,N_3183);
nand U5810 (N_5810,N_4376,N_4082);
nand U5811 (N_5811,N_3540,N_3558);
nand U5812 (N_5812,N_3038,N_2678);
xnor U5813 (N_5813,N_2744,N_3235);
nand U5814 (N_5814,N_3574,N_3735);
or U5815 (N_5815,N_4703,N_3106);
or U5816 (N_5816,N_4106,N_3174);
or U5817 (N_5817,N_3912,N_4337);
nor U5818 (N_5818,N_3352,N_3110);
nor U5819 (N_5819,N_3521,N_2796);
xor U5820 (N_5820,N_3959,N_3683);
nand U5821 (N_5821,N_3430,N_4641);
xor U5822 (N_5822,N_2964,N_3309);
nor U5823 (N_5823,N_4399,N_3900);
and U5824 (N_5824,N_2935,N_3416);
or U5825 (N_5825,N_3049,N_4800);
and U5826 (N_5826,N_4705,N_3783);
or U5827 (N_5827,N_4138,N_4546);
or U5828 (N_5828,N_4377,N_2786);
xnor U5829 (N_5829,N_4794,N_4130);
xnor U5830 (N_5830,N_4442,N_3567);
nand U5831 (N_5831,N_4326,N_3375);
xor U5832 (N_5832,N_4957,N_4005);
and U5833 (N_5833,N_3001,N_3029);
or U5834 (N_5834,N_2835,N_4873);
and U5835 (N_5835,N_4939,N_3296);
or U5836 (N_5836,N_4700,N_2918);
xnor U5837 (N_5837,N_4332,N_3470);
or U5838 (N_5838,N_2887,N_3504);
nand U5839 (N_5839,N_4870,N_3163);
nand U5840 (N_5840,N_2677,N_3623);
and U5841 (N_5841,N_4019,N_4210);
and U5842 (N_5842,N_4530,N_3888);
nor U5843 (N_5843,N_2681,N_4447);
and U5844 (N_5844,N_4493,N_3607);
nand U5845 (N_5845,N_3901,N_2694);
and U5846 (N_5846,N_3506,N_2819);
and U5847 (N_5847,N_3089,N_3239);
nand U5848 (N_5848,N_4940,N_3048);
and U5849 (N_5849,N_3802,N_3965);
and U5850 (N_5850,N_4642,N_4766);
or U5851 (N_5851,N_4292,N_4765);
xnor U5852 (N_5852,N_2506,N_2811);
xnor U5853 (N_5853,N_3098,N_3545);
xor U5854 (N_5854,N_4114,N_4999);
and U5855 (N_5855,N_4452,N_2671);
xnor U5856 (N_5856,N_4030,N_4354);
nor U5857 (N_5857,N_2645,N_3750);
nand U5858 (N_5858,N_4283,N_3920);
or U5859 (N_5859,N_2586,N_4234);
xor U5860 (N_5860,N_4686,N_2950);
and U5861 (N_5861,N_4033,N_2619);
xnor U5862 (N_5862,N_3923,N_4279);
and U5863 (N_5863,N_3902,N_3829);
and U5864 (N_5864,N_4348,N_2692);
or U5865 (N_5865,N_4575,N_3690);
and U5866 (N_5866,N_4102,N_3608);
xnor U5867 (N_5867,N_2653,N_4994);
or U5868 (N_5868,N_3532,N_3083);
and U5869 (N_5869,N_3960,N_4092);
and U5870 (N_5870,N_3795,N_4365);
nand U5871 (N_5871,N_3721,N_4083);
nor U5872 (N_5872,N_2576,N_4045);
xor U5873 (N_5873,N_3825,N_3261);
xnor U5874 (N_5874,N_3400,N_3453);
or U5875 (N_5875,N_3284,N_3768);
nor U5876 (N_5876,N_4500,N_2502);
or U5877 (N_5877,N_3834,N_3797);
and U5878 (N_5878,N_2631,N_3566);
or U5879 (N_5879,N_4865,N_3169);
or U5880 (N_5880,N_3050,N_4966);
xnor U5881 (N_5881,N_3517,N_3281);
xnor U5882 (N_5882,N_3384,N_4199);
and U5883 (N_5883,N_4537,N_2620);
nor U5884 (N_5884,N_4929,N_4384);
xor U5885 (N_5885,N_4544,N_4388);
nor U5886 (N_5886,N_3195,N_4670);
nand U5887 (N_5887,N_2947,N_4561);
xnor U5888 (N_5888,N_2783,N_3156);
xnor U5889 (N_5889,N_3872,N_3503);
xnor U5890 (N_5890,N_2776,N_2524);
and U5891 (N_5891,N_3808,N_3407);
nand U5892 (N_5892,N_2936,N_4659);
xnor U5893 (N_5893,N_4977,N_4490);
nand U5894 (N_5894,N_2765,N_4884);
nand U5895 (N_5895,N_3144,N_4740);
nor U5896 (N_5896,N_4985,N_2618);
xor U5897 (N_5897,N_2599,N_2762);
xnor U5898 (N_5898,N_4720,N_4141);
and U5899 (N_5899,N_4129,N_4913);
or U5900 (N_5900,N_3707,N_2941);
or U5901 (N_5901,N_2906,N_4535);
and U5902 (N_5902,N_3213,N_3218);
nor U5903 (N_5903,N_4423,N_4633);
nand U5904 (N_5904,N_2801,N_4712);
and U5905 (N_5905,N_4236,N_4356);
and U5906 (N_5906,N_3111,N_3847);
or U5907 (N_5907,N_3437,N_3885);
and U5908 (N_5908,N_3376,N_4964);
nor U5909 (N_5909,N_3649,N_4532);
nor U5910 (N_5910,N_2928,N_3441);
xnor U5911 (N_5911,N_4441,N_4551);
nor U5912 (N_5912,N_3054,N_3066);
or U5913 (N_5913,N_2960,N_3154);
nand U5914 (N_5914,N_2736,N_2507);
nor U5915 (N_5915,N_3771,N_3780);
or U5916 (N_5916,N_3748,N_2870);
nand U5917 (N_5917,N_4398,N_4137);
nor U5918 (N_5918,N_3919,N_4453);
and U5919 (N_5919,N_3787,N_3432);
and U5920 (N_5920,N_3245,N_3493);
nor U5921 (N_5921,N_4887,N_3512);
nor U5922 (N_5922,N_3319,N_4328);
or U5923 (N_5923,N_3398,N_4710);
xor U5924 (N_5924,N_4339,N_3324);
xor U5925 (N_5925,N_2662,N_3042);
xor U5926 (N_5926,N_3819,N_2554);
nor U5927 (N_5927,N_4528,N_2948);
nor U5928 (N_5928,N_4609,N_2582);
nor U5929 (N_5929,N_4008,N_2977);
or U5930 (N_5930,N_3760,N_3650);
xnor U5931 (N_5931,N_4011,N_4736);
or U5932 (N_5932,N_3047,N_3205);
nor U5933 (N_5933,N_3129,N_4606);
nor U5934 (N_5934,N_4342,N_3541);
xor U5935 (N_5935,N_4424,N_3904);
nor U5936 (N_5936,N_4413,N_4066);
and U5937 (N_5937,N_4644,N_3167);
nand U5938 (N_5938,N_4708,N_4847);
or U5939 (N_5939,N_4380,N_4411);
or U5940 (N_5940,N_3076,N_3146);
nand U5941 (N_5941,N_4549,N_4520);
nor U5942 (N_5942,N_3907,N_4522);
nand U5943 (N_5943,N_2689,N_4543);
or U5944 (N_5944,N_3534,N_4706);
nand U5945 (N_5945,N_3228,N_4498);
nand U5946 (N_5946,N_3982,N_3323);
xnor U5947 (N_5947,N_4023,N_2949);
or U5948 (N_5948,N_3528,N_2663);
or U5949 (N_5949,N_4079,N_3058);
or U5950 (N_5950,N_3033,N_3018);
xnor U5951 (N_5951,N_3880,N_4733);
xor U5952 (N_5952,N_4963,N_4758);
nor U5953 (N_5953,N_3879,N_4135);
nor U5954 (N_5954,N_4105,N_4661);
or U5955 (N_5955,N_4945,N_2512);
or U5956 (N_5956,N_4604,N_2996);
nand U5957 (N_5957,N_4826,N_3414);
nand U5958 (N_5958,N_4012,N_4225);
nor U5959 (N_5959,N_3498,N_3243);
and U5960 (N_5960,N_3684,N_3411);
nand U5961 (N_5961,N_4271,N_4560);
or U5962 (N_5962,N_4266,N_4110);
xor U5963 (N_5963,N_3571,N_3715);
xor U5964 (N_5964,N_3595,N_2541);
nor U5965 (N_5965,N_3092,N_2841);
nor U5966 (N_5966,N_4491,N_4457);
or U5967 (N_5967,N_2701,N_2856);
and U5968 (N_5968,N_3321,N_3223);
or U5969 (N_5969,N_4392,N_4040);
nor U5970 (N_5970,N_4759,N_4379);
xor U5971 (N_5971,N_4031,N_2634);
xor U5972 (N_5972,N_2740,N_4043);
nand U5973 (N_5973,N_4419,N_2610);
nor U5974 (N_5974,N_2615,N_2520);
or U5975 (N_5975,N_4217,N_2924);
or U5976 (N_5976,N_2920,N_3040);
nor U5977 (N_5977,N_3180,N_4403);
or U5978 (N_5978,N_3557,N_4133);
nand U5979 (N_5979,N_3070,N_4719);
or U5980 (N_5980,N_3588,N_4726);
and U5981 (N_5981,N_4351,N_4603);
nand U5982 (N_5982,N_3695,N_4018);
and U5983 (N_5983,N_3511,N_3688);
nor U5984 (N_5984,N_3348,N_3225);
xnor U5985 (N_5985,N_2876,N_4744);
nand U5986 (N_5986,N_3363,N_3361);
and U5987 (N_5987,N_4654,N_3171);
and U5988 (N_5988,N_3071,N_4782);
or U5989 (N_5989,N_4111,N_4052);
and U5990 (N_5990,N_4242,N_2690);
nor U5991 (N_5991,N_4980,N_4565);
nand U5992 (N_5992,N_4767,N_2737);
nor U5993 (N_5993,N_4205,N_4664);
nand U5994 (N_5994,N_4378,N_4277);
nor U5995 (N_5995,N_2871,N_4127);
and U5996 (N_5996,N_4821,N_4808);
nand U5997 (N_5997,N_4297,N_3543);
and U5998 (N_5998,N_2581,N_4313);
and U5999 (N_5999,N_2913,N_4446);
xnor U6000 (N_6000,N_4477,N_3869);
nor U6001 (N_6001,N_4355,N_3636);
or U6002 (N_6002,N_3777,N_2931);
nand U6003 (N_6003,N_4347,N_2669);
nand U6004 (N_6004,N_4254,N_4428);
nand U6005 (N_6005,N_4123,N_3550);
or U6006 (N_6006,N_3954,N_3657);
nor U6007 (N_6007,N_4094,N_3161);
or U6008 (N_6008,N_3844,N_4735);
nor U6009 (N_6009,N_4118,N_3796);
or U6010 (N_6010,N_3230,N_4058);
xor U6011 (N_6011,N_3974,N_2673);
or U6012 (N_6012,N_4497,N_3624);
xnor U6013 (N_6013,N_3704,N_3513);
xor U6014 (N_6014,N_3383,N_4162);
or U6015 (N_6015,N_4206,N_4218);
or U6016 (N_6016,N_2698,N_4526);
nor U6017 (N_6017,N_3963,N_4857);
nor U6018 (N_6018,N_4312,N_4057);
xnor U6019 (N_6019,N_2965,N_2528);
or U6020 (N_6020,N_3598,N_3622);
xor U6021 (N_6021,N_4160,N_3435);
nand U6022 (N_6022,N_2707,N_4727);
nor U6023 (N_6023,N_4795,N_3709);
and U6024 (N_6024,N_2659,N_3785);
nand U6025 (N_6025,N_2630,N_3364);
nand U6026 (N_6026,N_3465,N_4589);
nor U6027 (N_6027,N_4620,N_3520);
nand U6028 (N_6028,N_4969,N_4602);
or U6029 (N_6029,N_4502,N_3706);
or U6030 (N_6030,N_2579,N_4483);
and U6031 (N_6031,N_4505,N_3991);
xnor U6032 (N_6032,N_3899,N_4877);
or U6033 (N_6033,N_3207,N_2687);
or U6034 (N_6034,N_4866,N_2753);
and U6035 (N_6035,N_3609,N_3812);
nand U6036 (N_6036,N_4255,N_3593);
xor U6037 (N_6037,N_4170,N_4201);
or U6038 (N_6038,N_3741,N_3853);
or U6039 (N_6039,N_3227,N_3336);
and U6040 (N_6040,N_3581,N_4046);
or U6041 (N_6041,N_3060,N_4580);
nor U6042 (N_6042,N_3905,N_3577);
or U6043 (N_6043,N_3505,N_4261);
nor U6044 (N_6044,N_4677,N_2574);
or U6045 (N_6045,N_4169,N_2993);
xnor U6046 (N_6046,N_4240,N_2639);
nand U6047 (N_6047,N_4628,N_3883);
nand U6048 (N_6048,N_3613,N_4383);
or U6049 (N_6049,N_3555,N_3203);
nor U6050 (N_6050,N_3514,N_2832);
xnor U6051 (N_6051,N_3939,N_3762);
nand U6052 (N_6052,N_4880,N_2691);
or U6053 (N_6053,N_2616,N_2510);
and U6054 (N_6054,N_4173,N_4352);
or U6055 (N_6055,N_3136,N_3556);
xnor U6056 (N_6056,N_3937,N_4678);
and U6057 (N_6057,N_4156,N_3346);
nor U6058 (N_6058,N_3525,N_3377);
nand U6059 (N_6059,N_4984,N_4487);
nand U6060 (N_6060,N_4456,N_2674);
and U6061 (N_6061,N_2611,N_4318);
nand U6062 (N_6062,N_4839,N_2908);
nor U6063 (N_6063,N_3857,N_4564);
nand U6064 (N_6064,N_4250,N_4843);
nor U6065 (N_6065,N_4830,N_4463);
nand U6066 (N_6066,N_4871,N_3417);
xor U6067 (N_6067,N_3326,N_2892);
or U6068 (N_6068,N_4631,N_3175);
and U6069 (N_6069,N_4524,N_4034);
or U6070 (N_6070,N_2725,N_3172);
nor U6071 (N_6071,N_3833,N_3761);
or U6072 (N_6072,N_3979,N_3789);
nand U6073 (N_6073,N_3387,N_4184);
xnor U6074 (N_6074,N_3115,N_4814);
and U6075 (N_6075,N_2564,N_2695);
nor U6076 (N_6076,N_3428,N_3061);
nand U6077 (N_6077,N_3137,N_4390);
xnor U6078 (N_6078,N_4449,N_4362);
and U6079 (N_6079,N_3637,N_2983);
nor U6080 (N_6080,N_4897,N_4696);
nand U6081 (N_6081,N_3200,N_3763);
nor U6082 (N_6082,N_4103,N_4007);
nand U6083 (N_6083,N_2927,N_3827);
nor U6084 (N_6084,N_2580,N_3973);
and U6085 (N_6085,N_3288,N_4553);
nand U6086 (N_6086,N_4174,N_3452);
nor U6087 (N_6087,N_4781,N_3756);
xnor U6088 (N_6088,N_3486,N_2861);
and U6089 (N_6089,N_4707,N_3625);
and U6090 (N_6090,N_3733,N_3969);
xnor U6091 (N_6091,N_3738,N_2547);
nand U6092 (N_6092,N_3686,N_4754);
xnor U6093 (N_6093,N_4922,N_4750);
nand U6094 (N_6094,N_4755,N_3036);
or U6095 (N_6095,N_4931,N_2640);
nand U6096 (N_6096,N_3093,N_4475);
nor U6097 (N_6097,N_4662,N_3442);
nor U6098 (N_6098,N_2770,N_3996);
nand U6099 (N_6099,N_3781,N_3790);
and U6100 (N_6100,N_3436,N_4119);
nor U6101 (N_6101,N_2533,N_4763);
or U6102 (N_6102,N_3279,N_3147);
or U6103 (N_6103,N_2944,N_4574);
xor U6104 (N_6104,N_4142,N_2723);
nor U6105 (N_6105,N_3754,N_3159);
xnor U6106 (N_6106,N_3758,N_2814);
nor U6107 (N_6107,N_3656,N_4333);
nand U6108 (N_6108,N_4010,N_4555);
and U6109 (N_6109,N_2757,N_2952);
nand U6110 (N_6110,N_3747,N_3918);
or U6111 (N_6111,N_4181,N_2598);
xor U6112 (N_6112,N_2522,N_4015);
nand U6113 (N_6113,N_3948,N_4402);
xnor U6114 (N_6114,N_2696,N_4688);
xor U6115 (N_6115,N_4366,N_3165);
or U6116 (N_6116,N_2624,N_3813);
xnor U6117 (N_6117,N_2902,N_2932);
xor U6118 (N_6118,N_4473,N_2954);
or U6119 (N_6119,N_4540,N_3791);
xnor U6120 (N_6120,N_2523,N_2755);
or U6121 (N_6121,N_4307,N_2769);
nand U6122 (N_6122,N_2518,N_3298);
and U6123 (N_6123,N_2889,N_3473);
xnor U6124 (N_6124,N_4851,N_2545);
nor U6125 (N_6125,N_3476,N_4200);
nor U6126 (N_6126,N_4981,N_4340);
nand U6127 (N_6127,N_3929,N_3015);
and U6128 (N_6128,N_2886,N_3972);
nor U6129 (N_6129,N_2632,N_4655);
nand U6130 (N_6130,N_3913,N_3259);
nor U6131 (N_6131,N_2899,N_4025);
nand U6132 (N_6132,N_3082,N_3349);
nor U6133 (N_6133,N_4029,N_4405);
nand U6134 (N_6134,N_2905,N_3680);
or U6135 (N_6135,N_2789,N_4074);
xor U6136 (N_6136,N_2527,N_4226);
and U6137 (N_6137,N_4652,N_4425);
or U6138 (N_6138,N_3340,N_4256);
and U6139 (N_6139,N_4869,N_2853);
or U6140 (N_6140,N_4935,N_3908);
xor U6141 (N_6141,N_3100,N_4566);
or U6142 (N_6142,N_3620,N_4592);
xnor U6143 (N_6143,N_4467,N_2897);
and U6144 (N_6144,N_4235,N_3896);
nor U6145 (N_6145,N_4855,N_3749);
or U6146 (N_6146,N_3358,N_3197);
nor U6147 (N_6147,N_4166,N_3548);
nor U6148 (N_6148,N_4126,N_4918);
or U6149 (N_6149,N_3244,N_3940);
and U6150 (N_6150,N_3865,N_4003);
nor U6151 (N_6151,N_3086,N_3051);
or U6152 (N_6152,N_4305,N_4128);
nand U6153 (N_6153,N_4882,N_3494);
nor U6154 (N_6154,N_3202,N_3370);
xnor U6155 (N_6155,N_4844,N_4488);
or U6156 (N_6156,N_4525,N_3766);
and U6157 (N_6157,N_3772,N_4665);
nand U6158 (N_6158,N_2588,N_3466);
or U6159 (N_6159,N_4595,N_4962);
and U6160 (N_6160,N_3294,N_4787);
xor U6161 (N_6161,N_3984,N_2556);
nor U6162 (N_6162,N_4108,N_4615);
xor U6163 (N_6163,N_4699,N_3104);
nand U6164 (N_6164,N_4259,N_3552);
nand U6165 (N_6165,N_3983,N_2754);
and U6166 (N_6166,N_4811,N_2607);
nand U6167 (N_6167,N_3287,N_4919);
nor U6168 (N_6168,N_4721,N_2840);
or U6169 (N_6169,N_3420,N_3379);
and U6170 (N_6170,N_4459,N_4515);
nor U6171 (N_6171,N_2874,N_2557);
xnor U6172 (N_6172,N_3065,N_3304);
nand U6173 (N_6173,N_2916,N_3201);
xnor U6174 (N_6174,N_4290,N_4933);
and U6175 (N_6175,N_3196,N_4635);
or U6176 (N_6176,N_3037,N_2513);
or U6177 (N_6177,N_4681,N_2760);
and U6178 (N_6178,N_3677,N_2603);
nor U6179 (N_6179,N_4026,N_3565);
nand U6180 (N_6180,N_3993,N_3360);
or U6181 (N_6181,N_2505,N_2926);
xnor U6182 (N_6182,N_3032,N_4097);
nor U6183 (N_6183,N_2859,N_4368);
nor U6184 (N_6184,N_3719,N_4109);
or U6185 (N_6185,N_3952,N_3627);
nand U6186 (N_6186,N_4822,N_3021);
nand U6187 (N_6187,N_3523,N_4320);
or U6188 (N_6188,N_3903,N_4032);
or U6189 (N_6189,N_3217,N_2911);
nand U6190 (N_6190,N_3884,N_4258);
or U6191 (N_6191,N_4371,N_3850);
or U6192 (N_6192,N_2538,N_4738);
nand U6193 (N_6193,N_4000,N_4308);
nand U6194 (N_6194,N_3876,N_2719);
and U6195 (N_6195,N_3359,N_4924);
nand U6196 (N_6196,N_4784,N_3300);
nand U6197 (N_6197,N_2979,N_3931);
and U6198 (N_6198,N_3024,N_3875);
xnor U6199 (N_6199,N_4221,N_2976);
nand U6200 (N_6200,N_4779,N_4084);
or U6201 (N_6201,N_3866,N_2834);
or U6202 (N_6202,N_3835,N_4809);
or U6203 (N_6203,N_3410,N_3455);
nand U6204 (N_6204,N_3792,N_4343);
nand U6205 (N_6205,N_4658,N_4914);
nor U6206 (N_6206,N_3986,N_3020);
or U6207 (N_6207,N_4134,N_4587);
nor U6208 (N_6208,N_4728,N_3640);
nor U6209 (N_6209,N_4496,N_4805);
nor U6210 (N_6210,N_3830,N_2855);
xor U6211 (N_6211,N_3602,N_3312);
nand U6212 (N_6212,N_3997,N_4038);
and U6213 (N_6213,N_2784,N_3267);
and U6214 (N_6214,N_3821,N_3824);
xnor U6215 (N_6215,N_2679,N_2661);
or U6216 (N_6216,N_3266,N_3501);
nand U6217 (N_6217,N_4022,N_2713);
xnor U6218 (N_6218,N_3848,N_3408);
or U6219 (N_6219,N_3794,N_4444);
xor U6220 (N_6220,N_4341,N_4836);
or U6221 (N_6221,N_4476,N_4002);
or U6222 (N_6222,N_4125,N_4198);
and U6223 (N_6223,N_3731,N_3429);
nand U6224 (N_6224,N_4139,N_3064);
and U6225 (N_6225,N_3553,N_4848);
xnor U6226 (N_6226,N_2940,N_4612);
xor U6227 (N_6227,N_3405,N_4823);
and U6228 (N_6228,N_3658,N_3269);
or U6229 (N_6229,N_3614,N_4702);
xor U6230 (N_6230,N_3330,N_2914);
or U6231 (N_6231,N_3582,N_3981);
nor U6232 (N_6232,N_3729,N_3126);
nand U6233 (N_6233,N_4593,N_3063);
and U6234 (N_6234,N_4422,N_2508);
nor U6235 (N_6235,N_3732,N_2963);
or U6236 (N_6236,N_4637,N_3968);
nor U6237 (N_6237,N_4192,N_4485);
xor U6238 (N_6238,N_4374,N_3451);
or U6239 (N_6239,N_4934,N_2604);
and U6240 (N_6240,N_2766,N_3667);
nor U6241 (N_6241,N_4562,N_4860);
nand U6242 (N_6242,N_4523,N_3462);
nor U6243 (N_6243,N_3612,N_4634);
or U6244 (N_6244,N_3091,N_4230);
nand U6245 (N_6245,N_3013,N_3141);
and U6246 (N_6246,N_4510,N_4680);
xnor U6247 (N_6247,N_4600,N_3641);
nor U6248 (N_6248,N_4501,N_3413);
or U6249 (N_6249,N_2594,N_3961);
or U6250 (N_6250,N_2885,N_4447);
or U6251 (N_6251,N_4692,N_3817);
nand U6252 (N_6252,N_2873,N_3689);
xnor U6253 (N_6253,N_3754,N_4021);
xnor U6254 (N_6254,N_3298,N_4169);
or U6255 (N_6255,N_4203,N_3459);
nor U6256 (N_6256,N_3643,N_3272);
xnor U6257 (N_6257,N_3716,N_4007);
nor U6258 (N_6258,N_3541,N_4887);
and U6259 (N_6259,N_3492,N_3317);
nand U6260 (N_6260,N_4399,N_3986);
and U6261 (N_6261,N_4484,N_4287);
nor U6262 (N_6262,N_4879,N_3371);
nor U6263 (N_6263,N_4191,N_2845);
xnor U6264 (N_6264,N_4757,N_4307);
and U6265 (N_6265,N_4843,N_3529);
xor U6266 (N_6266,N_3312,N_3108);
or U6267 (N_6267,N_3170,N_4701);
and U6268 (N_6268,N_4395,N_4752);
nor U6269 (N_6269,N_4571,N_2553);
and U6270 (N_6270,N_3671,N_2908);
or U6271 (N_6271,N_2758,N_4887);
xnor U6272 (N_6272,N_4930,N_2597);
nand U6273 (N_6273,N_3786,N_4369);
xnor U6274 (N_6274,N_4756,N_3605);
nand U6275 (N_6275,N_2934,N_3988);
or U6276 (N_6276,N_3430,N_4341);
nand U6277 (N_6277,N_3469,N_2701);
and U6278 (N_6278,N_4597,N_3227);
nor U6279 (N_6279,N_3042,N_3388);
nor U6280 (N_6280,N_4681,N_4240);
xor U6281 (N_6281,N_4610,N_2574);
xor U6282 (N_6282,N_2921,N_3100);
nor U6283 (N_6283,N_4111,N_2606);
or U6284 (N_6284,N_3466,N_4467);
and U6285 (N_6285,N_3565,N_2811);
nor U6286 (N_6286,N_3833,N_2972);
and U6287 (N_6287,N_3051,N_3835);
xor U6288 (N_6288,N_2593,N_3896);
or U6289 (N_6289,N_4229,N_2737);
xor U6290 (N_6290,N_3826,N_4499);
or U6291 (N_6291,N_3316,N_3845);
xnor U6292 (N_6292,N_3958,N_2900);
and U6293 (N_6293,N_4716,N_2601);
nor U6294 (N_6294,N_4494,N_4837);
or U6295 (N_6295,N_2717,N_3943);
nor U6296 (N_6296,N_2830,N_4225);
nand U6297 (N_6297,N_4051,N_2530);
and U6298 (N_6298,N_3622,N_2576);
and U6299 (N_6299,N_4377,N_3073);
nor U6300 (N_6300,N_2771,N_4004);
nand U6301 (N_6301,N_3329,N_4120);
or U6302 (N_6302,N_4591,N_4145);
xnor U6303 (N_6303,N_3102,N_2630);
and U6304 (N_6304,N_4480,N_3800);
or U6305 (N_6305,N_2807,N_4381);
xor U6306 (N_6306,N_2910,N_4260);
or U6307 (N_6307,N_3373,N_3101);
xor U6308 (N_6308,N_4056,N_3883);
or U6309 (N_6309,N_4705,N_4016);
nor U6310 (N_6310,N_4017,N_4302);
or U6311 (N_6311,N_3724,N_2842);
and U6312 (N_6312,N_2612,N_4533);
nor U6313 (N_6313,N_4585,N_4534);
or U6314 (N_6314,N_4964,N_3556);
and U6315 (N_6315,N_3047,N_4771);
nor U6316 (N_6316,N_4924,N_3957);
nand U6317 (N_6317,N_3527,N_4172);
nor U6318 (N_6318,N_4423,N_4679);
nor U6319 (N_6319,N_4967,N_3771);
nor U6320 (N_6320,N_4892,N_3772);
xor U6321 (N_6321,N_3862,N_4693);
nor U6322 (N_6322,N_4687,N_3042);
and U6323 (N_6323,N_3521,N_2798);
nor U6324 (N_6324,N_3463,N_4076);
nor U6325 (N_6325,N_3011,N_4491);
and U6326 (N_6326,N_3332,N_4001);
nor U6327 (N_6327,N_4325,N_4567);
nor U6328 (N_6328,N_4558,N_4336);
and U6329 (N_6329,N_2717,N_4282);
xnor U6330 (N_6330,N_3374,N_3797);
nand U6331 (N_6331,N_4657,N_4850);
nor U6332 (N_6332,N_4843,N_2811);
or U6333 (N_6333,N_2940,N_4913);
nor U6334 (N_6334,N_3759,N_4888);
or U6335 (N_6335,N_4057,N_4476);
nand U6336 (N_6336,N_4721,N_4102);
nor U6337 (N_6337,N_3339,N_3563);
or U6338 (N_6338,N_3168,N_3086);
or U6339 (N_6339,N_4162,N_3007);
or U6340 (N_6340,N_4435,N_4599);
and U6341 (N_6341,N_2743,N_4239);
nand U6342 (N_6342,N_4987,N_3479);
nor U6343 (N_6343,N_2727,N_4230);
or U6344 (N_6344,N_4419,N_2799);
xnor U6345 (N_6345,N_4738,N_4162);
nand U6346 (N_6346,N_3810,N_4532);
and U6347 (N_6347,N_3575,N_4091);
or U6348 (N_6348,N_4994,N_4090);
or U6349 (N_6349,N_4941,N_3358);
nand U6350 (N_6350,N_3381,N_4375);
xor U6351 (N_6351,N_3586,N_4550);
nor U6352 (N_6352,N_3377,N_3038);
xnor U6353 (N_6353,N_3278,N_3042);
and U6354 (N_6354,N_4343,N_2815);
nand U6355 (N_6355,N_3606,N_3372);
xnor U6356 (N_6356,N_3630,N_2925);
nor U6357 (N_6357,N_4473,N_4395);
nand U6358 (N_6358,N_3426,N_4667);
nor U6359 (N_6359,N_3483,N_2983);
xnor U6360 (N_6360,N_3758,N_2525);
nor U6361 (N_6361,N_3516,N_3895);
xnor U6362 (N_6362,N_2703,N_3842);
nor U6363 (N_6363,N_2964,N_4832);
nand U6364 (N_6364,N_4054,N_4371);
or U6365 (N_6365,N_4455,N_4243);
nor U6366 (N_6366,N_3950,N_4030);
or U6367 (N_6367,N_3493,N_4005);
nand U6368 (N_6368,N_2761,N_3528);
nand U6369 (N_6369,N_3076,N_3809);
nor U6370 (N_6370,N_2552,N_3023);
nor U6371 (N_6371,N_3328,N_3775);
nor U6372 (N_6372,N_4876,N_3838);
nor U6373 (N_6373,N_4653,N_4026);
nor U6374 (N_6374,N_2618,N_3094);
or U6375 (N_6375,N_4892,N_4740);
nand U6376 (N_6376,N_3847,N_2978);
nor U6377 (N_6377,N_3248,N_4243);
and U6378 (N_6378,N_3115,N_3368);
xor U6379 (N_6379,N_3826,N_4356);
nor U6380 (N_6380,N_2822,N_4757);
and U6381 (N_6381,N_4879,N_4620);
and U6382 (N_6382,N_3605,N_2925);
nor U6383 (N_6383,N_2786,N_3040);
or U6384 (N_6384,N_3966,N_3411);
and U6385 (N_6385,N_2678,N_2742);
nand U6386 (N_6386,N_3350,N_2882);
and U6387 (N_6387,N_4154,N_2520);
nand U6388 (N_6388,N_3043,N_4407);
nand U6389 (N_6389,N_3464,N_4714);
xnor U6390 (N_6390,N_4061,N_3593);
and U6391 (N_6391,N_2564,N_3293);
nor U6392 (N_6392,N_2526,N_4902);
or U6393 (N_6393,N_4109,N_2668);
xnor U6394 (N_6394,N_2787,N_3056);
or U6395 (N_6395,N_3494,N_4761);
xor U6396 (N_6396,N_4727,N_3000);
or U6397 (N_6397,N_2620,N_3139);
xor U6398 (N_6398,N_2791,N_4149);
or U6399 (N_6399,N_3951,N_3709);
and U6400 (N_6400,N_2734,N_3544);
xor U6401 (N_6401,N_2668,N_4356);
nor U6402 (N_6402,N_2573,N_3372);
nand U6403 (N_6403,N_4875,N_4127);
and U6404 (N_6404,N_3438,N_3942);
nor U6405 (N_6405,N_2642,N_2690);
xnor U6406 (N_6406,N_3377,N_4514);
xor U6407 (N_6407,N_2646,N_4223);
or U6408 (N_6408,N_4551,N_3160);
xor U6409 (N_6409,N_2962,N_4287);
xor U6410 (N_6410,N_4660,N_4513);
nand U6411 (N_6411,N_3984,N_2918);
nand U6412 (N_6412,N_2532,N_2878);
or U6413 (N_6413,N_4674,N_3732);
and U6414 (N_6414,N_4311,N_4441);
and U6415 (N_6415,N_2770,N_4464);
xnor U6416 (N_6416,N_2604,N_4508);
xnor U6417 (N_6417,N_4630,N_2968);
nand U6418 (N_6418,N_4211,N_4950);
nor U6419 (N_6419,N_4008,N_4016);
nand U6420 (N_6420,N_2525,N_2745);
xor U6421 (N_6421,N_4278,N_4613);
nand U6422 (N_6422,N_3694,N_3376);
and U6423 (N_6423,N_4158,N_2958);
xnor U6424 (N_6424,N_4651,N_4283);
nand U6425 (N_6425,N_3342,N_4258);
xnor U6426 (N_6426,N_2657,N_2830);
or U6427 (N_6427,N_3176,N_4974);
and U6428 (N_6428,N_4312,N_3462);
or U6429 (N_6429,N_3619,N_4306);
or U6430 (N_6430,N_4487,N_4728);
or U6431 (N_6431,N_2587,N_3163);
and U6432 (N_6432,N_4226,N_3061);
and U6433 (N_6433,N_4994,N_3706);
and U6434 (N_6434,N_3426,N_3892);
xor U6435 (N_6435,N_2943,N_4488);
nor U6436 (N_6436,N_2918,N_3472);
nor U6437 (N_6437,N_4798,N_2876);
and U6438 (N_6438,N_3853,N_4812);
nor U6439 (N_6439,N_3490,N_2871);
and U6440 (N_6440,N_2954,N_4441);
nor U6441 (N_6441,N_2634,N_3133);
xnor U6442 (N_6442,N_3291,N_3821);
or U6443 (N_6443,N_4517,N_4885);
or U6444 (N_6444,N_2657,N_4657);
or U6445 (N_6445,N_2865,N_3393);
xor U6446 (N_6446,N_4046,N_2792);
nor U6447 (N_6447,N_3110,N_4012);
xor U6448 (N_6448,N_3916,N_2989);
nor U6449 (N_6449,N_3097,N_4761);
nor U6450 (N_6450,N_4503,N_4696);
nand U6451 (N_6451,N_4823,N_4686);
nor U6452 (N_6452,N_4111,N_3954);
or U6453 (N_6453,N_4483,N_4260);
xor U6454 (N_6454,N_4177,N_4355);
or U6455 (N_6455,N_3599,N_4883);
xor U6456 (N_6456,N_3938,N_2828);
xnor U6457 (N_6457,N_2628,N_4300);
and U6458 (N_6458,N_4460,N_2582);
nor U6459 (N_6459,N_3596,N_3894);
xor U6460 (N_6460,N_2780,N_2888);
nor U6461 (N_6461,N_3268,N_4131);
and U6462 (N_6462,N_4775,N_4520);
xnor U6463 (N_6463,N_3286,N_3122);
nand U6464 (N_6464,N_2519,N_4552);
xor U6465 (N_6465,N_3080,N_3337);
nand U6466 (N_6466,N_2950,N_2931);
xnor U6467 (N_6467,N_3361,N_3349);
nand U6468 (N_6468,N_4201,N_3388);
and U6469 (N_6469,N_2926,N_3093);
nand U6470 (N_6470,N_3474,N_4098);
nor U6471 (N_6471,N_4545,N_2868);
or U6472 (N_6472,N_4354,N_3488);
and U6473 (N_6473,N_3056,N_2513);
xnor U6474 (N_6474,N_4076,N_4948);
nor U6475 (N_6475,N_3398,N_4317);
xor U6476 (N_6476,N_3248,N_3383);
nor U6477 (N_6477,N_4990,N_4211);
or U6478 (N_6478,N_3191,N_4947);
or U6479 (N_6479,N_4382,N_4180);
nand U6480 (N_6480,N_3747,N_2742);
xor U6481 (N_6481,N_3599,N_4205);
nand U6482 (N_6482,N_4025,N_3388);
nor U6483 (N_6483,N_3460,N_3907);
nand U6484 (N_6484,N_4691,N_4001);
or U6485 (N_6485,N_4781,N_4587);
and U6486 (N_6486,N_2892,N_3162);
or U6487 (N_6487,N_4302,N_4438);
nor U6488 (N_6488,N_4382,N_3122);
and U6489 (N_6489,N_3018,N_3236);
nand U6490 (N_6490,N_4796,N_3087);
and U6491 (N_6491,N_3884,N_3589);
and U6492 (N_6492,N_4373,N_3460);
xnor U6493 (N_6493,N_3146,N_4548);
and U6494 (N_6494,N_4569,N_4982);
nand U6495 (N_6495,N_4369,N_3362);
nand U6496 (N_6496,N_4109,N_4395);
xnor U6497 (N_6497,N_3896,N_4253);
nand U6498 (N_6498,N_3277,N_2693);
and U6499 (N_6499,N_4529,N_3527);
or U6500 (N_6500,N_3680,N_4217);
xor U6501 (N_6501,N_4116,N_4385);
and U6502 (N_6502,N_3392,N_2510);
and U6503 (N_6503,N_4634,N_3206);
nor U6504 (N_6504,N_4000,N_4240);
nand U6505 (N_6505,N_4793,N_4984);
nand U6506 (N_6506,N_3633,N_4656);
nand U6507 (N_6507,N_3969,N_3288);
or U6508 (N_6508,N_3373,N_4506);
or U6509 (N_6509,N_3483,N_3533);
xnor U6510 (N_6510,N_2752,N_4984);
nor U6511 (N_6511,N_4764,N_3246);
xor U6512 (N_6512,N_4260,N_4595);
and U6513 (N_6513,N_3852,N_3935);
or U6514 (N_6514,N_4073,N_4719);
nor U6515 (N_6515,N_4726,N_3226);
nor U6516 (N_6516,N_2991,N_2690);
or U6517 (N_6517,N_4969,N_4504);
nand U6518 (N_6518,N_2712,N_3981);
nor U6519 (N_6519,N_4239,N_4031);
or U6520 (N_6520,N_4288,N_4203);
nand U6521 (N_6521,N_3175,N_3404);
nand U6522 (N_6522,N_3020,N_2584);
and U6523 (N_6523,N_4344,N_2771);
xnor U6524 (N_6524,N_2864,N_4927);
nor U6525 (N_6525,N_4166,N_4122);
nor U6526 (N_6526,N_4530,N_4231);
nor U6527 (N_6527,N_2725,N_2772);
nor U6528 (N_6528,N_3135,N_4625);
and U6529 (N_6529,N_3866,N_2628);
nor U6530 (N_6530,N_2752,N_3158);
and U6531 (N_6531,N_3634,N_4154);
or U6532 (N_6532,N_4840,N_4589);
or U6533 (N_6533,N_3551,N_3530);
nand U6534 (N_6534,N_3834,N_3300);
or U6535 (N_6535,N_2809,N_3189);
nor U6536 (N_6536,N_3789,N_4197);
or U6537 (N_6537,N_4774,N_4625);
and U6538 (N_6538,N_3211,N_3713);
nand U6539 (N_6539,N_3453,N_4940);
xor U6540 (N_6540,N_3087,N_3389);
xor U6541 (N_6541,N_3932,N_3269);
xor U6542 (N_6542,N_4261,N_4820);
nor U6543 (N_6543,N_3451,N_4278);
or U6544 (N_6544,N_3877,N_2555);
nand U6545 (N_6545,N_2923,N_4000);
nor U6546 (N_6546,N_4174,N_4863);
xor U6547 (N_6547,N_2596,N_4233);
or U6548 (N_6548,N_4769,N_4866);
nand U6549 (N_6549,N_2794,N_3816);
or U6550 (N_6550,N_3908,N_4193);
nor U6551 (N_6551,N_2604,N_4453);
nor U6552 (N_6552,N_4125,N_4305);
nor U6553 (N_6553,N_3267,N_4096);
xor U6554 (N_6554,N_4270,N_3163);
and U6555 (N_6555,N_2688,N_3337);
and U6556 (N_6556,N_4964,N_3713);
xor U6557 (N_6557,N_4403,N_3177);
nor U6558 (N_6558,N_3474,N_3119);
nor U6559 (N_6559,N_2854,N_4027);
xor U6560 (N_6560,N_2947,N_3967);
or U6561 (N_6561,N_2938,N_4424);
nor U6562 (N_6562,N_4400,N_2968);
and U6563 (N_6563,N_4645,N_2828);
nand U6564 (N_6564,N_3842,N_3814);
and U6565 (N_6565,N_4418,N_4638);
nor U6566 (N_6566,N_2671,N_4832);
and U6567 (N_6567,N_3289,N_2882);
nand U6568 (N_6568,N_4472,N_2904);
or U6569 (N_6569,N_4636,N_3585);
nor U6570 (N_6570,N_4528,N_4554);
or U6571 (N_6571,N_4690,N_3218);
nor U6572 (N_6572,N_4650,N_4105);
nand U6573 (N_6573,N_4121,N_4857);
xnor U6574 (N_6574,N_3640,N_2858);
or U6575 (N_6575,N_3912,N_4773);
and U6576 (N_6576,N_4684,N_4520);
xor U6577 (N_6577,N_4965,N_3702);
and U6578 (N_6578,N_4217,N_4280);
nand U6579 (N_6579,N_2682,N_2784);
nor U6580 (N_6580,N_3789,N_2761);
or U6581 (N_6581,N_4793,N_4751);
nor U6582 (N_6582,N_2683,N_3437);
or U6583 (N_6583,N_3994,N_4742);
xor U6584 (N_6584,N_4806,N_4674);
xor U6585 (N_6585,N_4598,N_4550);
nor U6586 (N_6586,N_2968,N_2685);
or U6587 (N_6587,N_3835,N_3091);
nor U6588 (N_6588,N_4414,N_2998);
and U6589 (N_6589,N_3621,N_3184);
and U6590 (N_6590,N_3194,N_3130);
nand U6591 (N_6591,N_4319,N_4409);
and U6592 (N_6592,N_3762,N_4839);
xor U6593 (N_6593,N_2700,N_4642);
xnor U6594 (N_6594,N_4715,N_2541);
xnor U6595 (N_6595,N_4972,N_3903);
and U6596 (N_6596,N_3415,N_3815);
xnor U6597 (N_6597,N_4865,N_3697);
and U6598 (N_6598,N_4999,N_3845);
or U6599 (N_6599,N_4428,N_4682);
nand U6600 (N_6600,N_3302,N_2945);
nor U6601 (N_6601,N_4149,N_3969);
xor U6602 (N_6602,N_4328,N_3248);
or U6603 (N_6603,N_4199,N_2518);
xnor U6604 (N_6604,N_2783,N_3332);
or U6605 (N_6605,N_2894,N_2962);
and U6606 (N_6606,N_2558,N_4694);
nand U6607 (N_6607,N_3909,N_3595);
xnor U6608 (N_6608,N_4655,N_3106);
and U6609 (N_6609,N_4561,N_4923);
and U6610 (N_6610,N_3538,N_3733);
xnor U6611 (N_6611,N_4598,N_3706);
nor U6612 (N_6612,N_3629,N_4266);
nand U6613 (N_6613,N_3574,N_3826);
or U6614 (N_6614,N_3328,N_4886);
or U6615 (N_6615,N_4419,N_3652);
nand U6616 (N_6616,N_2657,N_4165);
nor U6617 (N_6617,N_2850,N_4717);
xnor U6618 (N_6618,N_3066,N_2723);
nor U6619 (N_6619,N_4728,N_3911);
xor U6620 (N_6620,N_3121,N_2894);
xor U6621 (N_6621,N_4691,N_2900);
xor U6622 (N_6622,N_4345,N_4098);
and U6623 (N_6623,N_4270,N_4825);
or U6624 (N_6624,N_4386,N_4054);
nand U6625 (N_6625,N_4459,N_4625);
nor U6626 (N_6626,N_4429,N_3818);
or U6627 (N_6627,N_2576,N_4016);
nor U6628 (N_6628,N_4584,N_2692);
nand U6629 (N_6629,N_4224,N_4671);
and U6630 (N_6630,N_3502,N_4952);
and U6631 (N_6631,N_4919,N_2664);
or U6632 (N_6632,N_2924,N_4026);
and U6633 (N_6633,N_4500,N_2889);
and U6634 (N_6634,N_2554,N_3583);
xnor U6635 (N_6635,N_3198,N_2927);
xnor U6636 (N_6636,N_3474,N_2827);
xor U6637 (N_6637,N_3308,N_3413);
nand U6638 (N_6638,N_4260,N_4571);
nor U6639 (N_6639,N_4253,N_4878);
or U6640 (N_6640,N_4421,N_3047);
nand U6641 (N_6641,N_3152,N_3599);
or U6642 (N_6642,N_2941,N_3595);
nor U6643 (N_6643,N_4716,N_4739);
nand U6644 (N_6644,N_2993,N_4882);
or U6645 (N_6645,N_3960,N_2891);
nand U6646 (N_6646,N_2832,N_4744);
nand U6647 (N_6647,N_4305,N_2915);
and U6648 (N_6648,N_2577,N_2667);
or U6649 (N_6649,N_4706,N_3479);
xor U6650 (N_6650,N_4330,N_2709);
and U6651 (N_6651,N_4073,N_2922);
or U6652 (N_6652,N_2698,N_2611);
xor U6653 (N_6653,N_4118,N_2748);
and U6654 (N_6654,N_3518,N_4024);
or U6655 (N_6655,N_4305,N_2598);
xnor U6656 (N_6656,N_3005,N_3640);
and U6657 (N_6657,N_4666,N_3326);
nand U6658 (N_6658,N_3881,N_4215);
nor U6659 (N_6659,N_3728,N_3122);
nor U6660 (N_6660,N_3189,N_3337);
nor U6661 (N_6661,N_3651,N_4831);
or U6662 (N_6662,N_2851,N_4246);
nor U6663 (N_6663,N_4153,N_3682);
nor U6664 (N_6664,N_4208,N_4882);
or U6665 (N_6665,N_2588,N_4112);
and U6666 (N_6666,N_4131,N_3969);
and U6667 (N_6667,N_2902,N_4248);
xnor U6668 (N_6668,N_4852,N_3546);
nand U6669 (N_6669,N_3093,N_3682);
nor U6670 (N_6670,N_3299,N_3794);
nor U6671 (N_6671,N_2958,N_4635);
xnor U6672 (N_6672,N_3062,N_3153);
nand U6673 (N_6673,N_2880,N_2729);
nor U6674 (N_6674,N_3095,N_3631);
or U6675 (N_6675,N_4907,N_3987);
xnor U6676 (N_6676,N_3971,N_3070);
xor U6677 (N_6677,N_3961,N_4986);
nor U6678 (N_6678,N_3117,N_4105);
nand U6679 (N_6679,N_3166,N_3603);
nand U6680 (N_6680,N_2524,N_4656);
xnor U6681 (N_6681,N_3165,N_4302);
xnor U6682 (N_6682,N_4183,N_3269);
and U6683 (N_6683,N_2843,N_3425);
nand U6684 (N_6684,N_4550,N_4496);
or U6685 (N_6685,N_4665,N_4200);
xnor U6686 (N_6686,N_3003,N_4093);
nand U6687 (N_6687,N_3674,N_4856);
and U6688 (N_6688,N_4346,N_3634);
or U6689 (N_6689,N_2925,N_4503);
nor U6690 (N_6690,N_4315,N_2799);
or U6691 (N_6691,N_2595,N_2874);
or U6692 (N_6692,N_3137,N_2691);
nand U6693 (N_6693,N_3782,N_2710);
nor U6694 (N_6694,N_4054,N_2595);
and U6695 (N_6695,N_4760,N_3587);
nand U6696 (N_6696,N_3185,N_2878);
and U6697 (N_6697,N_4472,N_3601);
nand U6698 (N_6698,N_3528,N_4068);
nand U6699 (N_6699,N_4668,N_3163);
nor U6700 (N_6700,N_2715,N_3192);
and U6701 (N_6701,N_3722,N_3872);
nor U6702 (N_6702,N_3950,N_3728);
nor U6703 (N_6703,N_4500,N_2517);
and U6704 (N_6704,N_3794,N_4719);
xor U6705 (N_6705,N_3303,N_3823);
nor U6706 (N_6706,N_2780,N_3885);
and U6707 (N_6707,N_2986,N_2980);
nor U6708 (N_6708,N_3296,N_3627);
and U6709 (N_6709,N_2539,N_4304);
xnor U6710 (N_6710,N_4507,N_4514);
nand U6711 (N_6711,N_3363,N_3703);
and U6712 (N_6712,N_4243,N_3809);
nand U6713 (N_6713,N_4838,N_4711);
or U6714 (N_6714,N_2649,N_4983);
or U6715 (N_6715,N_4021,N_4702);
and U6716 (N_6716,N_3601,N_4645);
xor U6717 (N_6717,N_3672,N_3607);
xor U6718 (N_6718,N_2623,N_3031);
nand U6719 (N_6719,N_3007,N_2860);
nand U6720 (N_6720,N_4604,N_2662);
or U6721 (N_6721,N_4661,N_3297);
nor U6722 (N_6722,N_4120,N_2961);
or U6723 (N_6723,N_4538,N_2915);
nand U6724 (N_6724,N_2925,N_3939);
nand U6725 (N_6725,N_2512,N_3107);
nor U6726 (N_6726,N_2970,N_3579);
nand U6727 (N_6727,N_3054,N_3631);
nor U6728 (N_6728,N_2625,N_3322);
and U6729 (N_6729,N_4528,N_3995);
and U6730 (N_6730,N_4150,N_2610);
nor U6731 (N_6731,N_4776,N_3623);
or U6732 (N_6732,N_4297,N_4257);
xnor U6733 (N_6733,N_3540,N_4403);
nand U6734 (N_6734,N_3056,N_2612);
and U6735 (N_6735,N_4461,N_4546);
and U6736 (N_6736,N_3047,N_4018);
and U6737 (N_6737,N_3128,N_2761);
nor U6738 (N_6738,N_4903,N_3208);
nand U6739 (N_6739,N_4979,N_2982);
xor U6740 (N_6740,N_2918,N_2825);
and U6741 (N_6741,N_2581,N_3298);
or U6742 (N_6742,N_4987,N_3884);
or U6743 (N_6743,N_3357,N_4736);
nor U6744 (N_6744,N_4098,N_3443);
and U6745 (N_6745,N_2556,N_2542);
or U6746 (N_6746,N_4213,N_4230);
or U6747 (N_6747,N_3317,N_3144);
nand U6748 (N_6748,N_4309,N_3685);
and U6749 (N_6749,N_3185,N_3432);
or U6750 (N_6750,N_4117,N_4827);
xnor U6751 (N_6751,N_2587,N_3272);
xnor U6752 (N_6752,N_2671,N_2659);
nor U6753 (N_6753,N_3423,N_4796);
nor U6754 (N_6754,N_4207,N_3932);
nand U6755 (N_6755,N_4853,N_3216);
xor U6756 (N_6756,N_4004,N_3775);
nand U6757 (N_6757,N_4185,N_3116);
or U6758 (N_6758,N_2542,N_3024);
nand U6759 (N_6759,N_3192,N_4658);
nor U6760 (N_6760,N_2816,N_4670);
nor U6761 (N_6761,N_3872,N_2962);
nand U6762 (N_6762,N_3615,N_3206);
nor U6763 (N_6763,N_3448,N_2702);
or U6764 (N_6764,N_3550,N_2922);
or U6765 (N_6765,N_4886,N_4056);
xnor U6766 (N_6766,N_3093,N_3943);
nor U6767 (N_6767,N_4620,N_2853);
nor U6768 (N_6768,N_4877,N_4559);
or U6769 (N_6769,N_3971,N_4120);
or U6770 (N_6770,N_4960,N_4023);
nand U6771 (N_6771,N_3237,N_4725);
or U6772 (N_6772,N_4042,N_3904);
or U6773 (N_6773,N_4168,N_3809);
or U6774 (N_6774,N_2580,N_4811);
xnor U6775 (N_6775,N_3096,N_4899);
or U6776 (N_6776,N_4380,N_3242);
nor U6777 (N_6777,N_2674,N_3782);
nor U6778 (N_6778,N_3725,N_4712);
and U6779 (N_6779,N_4088,N_4696);
and U6780 (N_6780,N_3961,N_2873);
nand U6781 (N_6781,N_2731,N_3567);
nor U6782 (N_6782,N_3983,N_4024);
or U6783 (N_6783,N_4694,N_3609);
nor U6784 (N_6784,N_2938,N_2922);
nand U6785 (N_6785,N_4341,N_3291);
nand U6786 (N_6786,N_4363,N_4802);
nand U6787 (N_6787,N_2723,N_2806);
xor U6788 (N_6788,N_3549,N_2739);
nand U6789 (N_6789,N_4123,N_4779);
nor U6790 (N_6790,N_2787,N_4322);
xnor U6791 (N_6791,N_2528,N_4277);
nand U6792 (N_6792,N_2999,N_4506);
nand U6793 (N_6793,N_2532,N_4832);
nand U6794 (N_6794,N_4900,N_4664);
xnor U6795 (N_6795,N_3268,N_4134);
nand U6796 (N_6796,N_3613,N_4796);
nor U6797 (N_6797,N_3222,N_2905);
and U6798 (N_6798,N_4425,N_4329);
nand U6799 (N_6799,N_4899,N_3471);
xor U6800 (N_6800,N_3663,N_2695);
nand U6801 (N_6801,N_4103,N_3693);
xnor U6802 (N_6802,N_3916,N_2895);
nand U6803 (N_6803,N_3086,N_4589);
nand U6804 (N_6804,N_2904,N_4293);
and U6805 (N_6805,N_2854,N_4715);
xor U6806 (N_6806,N_3249,N_3055);
xnor U6807 (N_6807,N_4198,N_4177);
nor U6808 (N_6808,N_4293,N_4006);
and U6809 (N_6809,N_2689,N_2741);
nor U6810 (N_6810,N_4456,N_4608);
nor U6811 (N_6811,N_3733,N_4632);
nor U6812 (N_6812,N_4211,N_4371);
xor U6813 (N_6813,N_3614,N_3585);
or U6814 (N_6814,N_4894,N_3983);
nor U6815 (N_6815,N_3669,N_2802);
xor U6816 (N_6816,N_4343,N_2554);
and U6817 (N_6817,N_3506,N_2612);
nand U6818 (N_6818,N_4211,N_4393);
xor U6819 (N_6819,N_3979,N_4891);
nor U6820 (N_6820,N_2536,N_4775);
nor U6821 (N_6821,N_3017,N_3539);
and U6822 (N_6822,N_4747,N_4153);
nor U6823 (N_6823,N_4484,N_3084);
nor U6824 (N_6824,N_3038,N_3681);
nor U6825 (N_6825,N_3652,N_3729);
and U6826 (N_6826,N_3700,N_3161);
and U6827 (N_6827,N_4957,N_3282);
xnor U6828 (N_6828,N_3624,N_4066);
xor U6829 (N_6829,N_4109,N_3957);
and U6830 (N_6830,N_4870,N_4637);
and U6831 (N_6831,N_2631,N_4512);
nor U6832 (N_6832,N_4235,N_4153);
and U6833 (N_6833,N_4958,N_3124);
xnor U6834 (N_6834,N_2508,N_4621);
nor U6835 (N_6835,N_3565,N_3309);
nand U6836 (N_6836,N_4020,N_3152);
nand U6837 (N_6837,N_4835,N_3069);
xnor U6838 (N_6838,N_3107,N_4900);
or U6839 (N_6839,N_3302,N_3520);
and U6840 (N_6840,N_4375,N_4193);
nand U6841 (N_6841,N_2605,N_4541);
nand U6842 (N_6842,N_4946,N_4341);
nor U6843 (N_6843,N_4984,N_3576);
nor U6844 (N_6844,N_3884,N_4091);
or U6845 (N_6845,N_4227,N_4365);
nor U6846 (N_6846,N_3103,N_2965);
nor U6847 (N_6847,N_4392,N_2505);
nor U6848 (N_6848,N_3836,N_3724);
or U6849 (N_6849,N_3386,N_3904);
and U6850 (N_6850,N_3617,N_3810);
nand U6851 (N_6851,N_3682,N_4733);
or U6852 (N_6852,N_3854,N_3090);
or U6853 (N_6853,N_2516,N_3603);
or U6854 (N_6854,N_3744,N_3679);
and U6855 (N_6855,N_2592,N_3848);
xnor U6856 (N_6856,N_4857,N_3738);
or U6857 (N_6857,N_3130,N_3200);
or U6858 (N_6858,N_3102,N_4969);
xor U6859 (N_6859,N_3665,N_4553);
xnor U6860 (N_6860,N_4954,N_2789);
nor U6861 (N_6861,N_3092,N_4940);
nand U6862 (N_6862,N_2904,N_2944);
nor U6863 (N_6863,N_4358,N_2934);
or U6864 (N_6864,N_2961,N_4680);
xnor U6865 (N_6865,N_4567,N_3781);
nor U6866 (N_6866,N_4059,N_4544);
nand U6867 (N_6867,N_4587,N_2643);
or U6868 (N_6868,N_2548,N_3606);
xor U6869 (N_6869,N_3857,N_3406);
and U6870 (N_6870,N_4637,N_3349);
xnor U6871 (N_6871,N_4758,N_3386);
or U6872 (N_6872,N_4026,N_3454);
or U6873 (N_6873,N_3727,N_4687);
nor U6874 (N_6874,N_4986,N_3940);
nand U6875 (N_6875,N_2882,N_2628);
nor U6876 (N_6876,N_3634,N_4729);
and U6877 (N_6877,N_2868,N_3753);
or U6878 (N_6878,N_4305,N_3942);
and U6879 (N_6879,N_3221,N_3100);
and U6880 (N_6880,N_2506,N_4801);
or U6881 (N_6881,N_3416,N_4079);
or U6882 (N_6882,N_4567,N_4394);
nor U6883 (N_6883,N_3328,N_3788);
nand U6884 (N_6884,N_2601,N_2513);
xnor U6885 (N_6885,N_3276,N_2614);
or U6886 (N_6886,N_2864,N_3109);
nor U6887 (N_6887,N_4360,N_4344);
xor U6888 (N_6888,N_4832,N_4889);
nor U6889 (N_6889,N_3371,N_2856);
and U6890 (N_6890,N_4998,N_3871);
and U6891 (N_6891,N_3397,N_2934);
and U6892 (N_6892,N_4249,N_2586);
or U6893 (N_6893,N_4485,N_3456);
xor U6894 (N_6894,N_4284,N_3188);
and U6895 (N_6895,N_4048,N_4876);
nor U6896 (N_6896,N_2526,N_2862);
nand U6897 (N_6897,N_4408,N_2746);
or U6898 (N_6898,N_2952,N_4514);
nor U6899 (N_6899,N_2647,N_2639);
nand U6900 (N_6900,N_4259,N_4599);
xnor U6901 (N_6901,N_4995,N_3076);
nor U6902 (N_6902,N_2731,N_4338);
and U6903 (N_6903,N_2842,N_4102);
nand U6904 (N_6904,N_4897,N_3074);
or U6905 (N_6905,N_3193,N_3209);
or U6906 (N_6906,N_4842,N_2866);
xnor U6907 (N_6907,N_4961,N_3807);
or U6908 (N_6908,N_3890,N_2833);
xor U6909 (N_6909,N_4320,N_3367);
nor U6910 (N_6910,N_4807,N_3673);
or U6911 (N_6911,N_2576,N_4845);
and U6912 (N_6912,N_3070,N_3710);
and U6913 (N_6913,N_3284,N_4648);
nor U6914 (N_6914,N_2916,N_4257);
nor U6915 (N_6915,N_3507,N_2901);
nor U6916 (N_6916,N_2692,N_4764);
nand U6917 (N_6917,N_3448,N_2835);
and U6918 (N_6918,N_4130,N_3386);
nand U6919 (N_6919,N_4807,N_3194);
xnor U6920 (N_6920,N_4025,N_4371);
nand U6921 (N_6921,N_3306,N_4426);
and U6922 (N_6922,N_2974,N_4939);
and U6923 (N_6923,N_3592,N_4684);
xor U6924 (N_6924,N_3636,N_3255);
or U6925 (N_6925,N_4853,N_4217);
or U6926 (N_6926,N_3829,N_3691);
or U6927 (N_6927,N_3317,N_2802);
or U6928 (N_6928,N_3860,N_4201);
and U6929 (N_6929,N_4038,N_3867);
nor U6930 (N_6930,N_4579,N_4865);
and U6931 (N_6931,N_3278,N_3054);
and U6932 (N_6932,N_4318,N_4771);
and U6933 (N_6933,N_3326,N_3949);
nor U6934 (N_6934,N_3573,N_2601);
and U6935 (N_6935,N_2597,N_2875);
and U6936 (N_6936,N_2773,N_3249);
or U6937 (N_6937,N_3088,N_3243);
nand U6938 (N_6938,N_4355,N_2798);
nor U6939 (N_6939,N_3887,N_4302);
nor U6940 (N_6940,N_4822,N_3516);
xnor U6941 (N_6941,N_4652,N_3027);
xnor U6942 (N_6942,N_4246,N_3382);
xor U6943 (N_6943,N_4143,N_4314);
and U6944 (N_6944,N_4143,N_3638);
or U6945 (N_6945,N_2723,N_2772);
xor U6946 (N_6946,N_3225,N_4849);
or U6947 (N_6947,N_4280,N_3704);
nor U6948 (N_6948,N_3591,N_3863);
xnor U6949 (N_6949,N_3227,N_4178);
and U6950 (N_6950,N_2890,N_3741);
nor U6951 (N_6951,N_4435,N_3745);
xnor U6952 (N_6952,N_3569,N_3449);
or U6953 (N_6953,N_4746,N_2766);
nor U6954 (N_6954,N_3773,N_4108);
xor U6955 (N_6955,N_2576,N_3556);
nor U6956 (N_6956,N_3510,N_2605);
or U6957 (N_6957,N_2890,N_2611);
nand U6958 (N_6958,N_4773,N_2582);
xor U6959 (N_6959,N_2677,N_3002);
nand U6960 (N_6960,N_4959,N_4740);
xnor U6961 (N_6961,N_3430,N_4159);
and U6962 (N_6962,N_2842,N_3709);
nor U6963 (N_6963,N_2936,N_4233);
xor U6964 (N_6964,N_4830,N_4631);
nor U6965 (N_6965,N_4391,N_4110);
and U6966 (N_6966,N_3164,N_3751);
or U6967 (N_6967,N_3777,N_3876);
and U6968 (N_6968,N_4928,N_4620);
xnor U6969 (N_6969,N_3331,N_3782);
nand U6970 (N_6970,N_3198,N_4514);
xor U6971 (N_6971,N_4061,N_3400);
xor U6972 (N_6972,N_4992,N_4591);
nand U6973 (N_6973,N_3203,N_3970);
nand U6974 (N_6974,N_4494,N_3463);
and U6975 (N_6975,N_3863,N_4530);
xor U6976 (N_6976,N_4777,N_4397);
xnor U6977 (N_6977,N_4157,N_3931);
nand U6978 (N_6978,N_3176,N_3513);
and U6979 (N_6979,N_3777,N_2811);
and U6980 (N_6980,N_3285,N_3774);
or U6981 (N_6981,N_3062,N_4099);
xor U6982 (N_6982,N_2843,N_3626);
and U6983 (N_6983,N_4915,N_3018);
nand U6984 (N_6984,N_4101,N_2656);
and U6985 (N_6985,N_3058,N_4640);
xor U6986 (N_6986,N_3474,N_2958);
xor U6987 (N_6987,N_3164,N_4694);
nand U6988 (N_6988,N_3055,N_3476);
xnor U6989 (N_6989,N_4791,N_4052);
or U6990 (N_6990,N_4838,N_3744);
and U6991 (N_6991,N_3356,N_4650);
nand U6992 (N_6992,N_4506,N_2689);
nor U6993 (N_6993,N_3872,N_4447);
and U6994 (N_6994,N_3904,N_4637);
or U6995 (N_6995,N_3353,N_2766);
nor U6996 (N_6996,N_3185,N_3775);
xor U6997 (N_6997,N_2972,N_2861);
xor U6998 (N_6998,N_3656,N_4904);
or U6999 (N_6999,N_4157,N_3017);
nor U7000 (N_7000,N_2773,N_4565);
nor U7001 (N_7001,N_2963,N_2529);
nor U7002 (N_7002,N_3011,N_2742);
nand U7003 (N_7003,N_3586,N_3025);
xor U7004 (N_7004,N_3501,N_3688);
or U7005 (N_7005,N_2800,N_4448);
nor U7006 (N_7006,N_3928,N_3711);
and U7007 (N_7007,N_4765,N_4047);
and U7008 (N_7008,N_3225,N_4717);
nand U7009 (N_7009,N_3276,N_4311);
nand U7010 (N_7010,N_3769,N_4733);
nand U7011 (N_7011,N_2662,N_4242);
and U7012 (N_7012,N_2783,N_3232);
nor U7013 (N_7013,N_3887,N_3285);
nor U7014 (N_7014,N_3022,N_3427);
xor U7015 (N_7015,N_4146,N_4224);
nor U7016 (N_7016,N_3224,N_4377);
xor U7017 (N_7017,N_3687,N_4060);
nor U7018 (N_7018,N_2947,N_4690);
nor U7019 (N_7019,N_2990,N_2970);
or U7020 (N_7020,N_4475,N_2721);
and U7021 (N_7021,N_4613,N_3009);
xnor U7022 (N_7022,N_3487,N_3532);
nand U7023 (N_7023,N_4492,N_2809);
xor U7024 (N_7024,N_2973,N_3446);
nor U7025 (N_7025,N_4788,N_2684);
or U7026 (N_7026,N_3040,N_4005);
nor U7027 (N_7027,N_3110,N_3108);
nor U7028 (N_7028,N_4025,N_3591);
or U7029 (N_7029,N_4116,N_3223);
xor U7030 (N_7030,N_4657,N_4561);
nor U7031 (N_7031,N_2553,N_4274);
and U7032 (N_7032,N_3803,N_4466);
nor U7033 (N_7033,N_4497,N_3286);
or U7034 (N_7034,N_4725,N_2955);
xor U7035 (N_7035,N_4873,N_3768);
nor U7036 (N_7036,N_4505,N_2920);
xor U7037 (N_7037,N_4872,N_3847);
nand U7038 (N_7038,N_3683,N_3422);
and U7039 (N_7039,N_3887,N_4584);
nand U7040 (N_7040,N_3681,N_3551);
nor U7041 (N_7041,N_4458,N_3477);
xor U7042 (N_7042,N_2877,N_4143);
nand U7043 (N_7043,N_4344,N_3180);
or U7044 (N_7044,N_3262,N_4344);
xnor U7045 (N_7045,N_2708,N_4305);
xnor U7046 (N_7046,N_3859,N_4614);
nand U7047 (N_7047,N_4419,N_3278);
and U7048 (N_7048,N_3534,N_3719);
nand U7049 (N_7049,N_4773,N_4850);
nand U7050 (N_7050,N_3150,N_4617);
xor U7051 (N_7051,N_3843,N_3062);
or U7052 (N_7052,N_3244,N_2749);
xnor U7053 (N_7053,N_2683,N_3793);
and U7054 (N_7054,N_4173,N_3649);
and U7055 (N_7055,N_4714,N_2753);
and U7056 (N_7056,N_3053,N_2919);
nand U7057 (N_7057,N_3675,N_3574);
xor U7058 (N_7058,N_3487,N_3235);
xnor U7059 (N_7059,N_3908,N_3549);
nor U7060 (N_7060,N_3742,N_3010);
xnor U7061 (N_7061,N_4426,N_3167);
and U7062 (N_7062,N_2916,N_3326);
and U7063 (N_7063,N_2863,N_2509);
or U7064 (N_7064,N_4370,N_4974);
nand U7065 (N_7065,N_3669,N_2669);
nor U7066 (N_7066,N_3233,N_4918);
nor U7067 (N_7067,N_3016,N_2737);
and U7068 (N_7068,N_2984,N_2604);
or U7069 (N_7069,N_2654,N_4536);
nor U7070 (N_7070,N_3577,N_4511);
and U7071 (N_7071,N_3000,N_3187);
nand U7072 (N_7072,N_4942,N_4386);
xnor U7073 (N_7073,N_3347,N_3291);
or U7074 (N_7074,N_4187,N_4397);
and U7075 (N_7075,N_4105,N_3908);
xor U7076 (N_7076,N_4743,N_2887);
xor U7077 (N_7077,N_4049,N_3858);
nand U7078 (N_7078,N_4948,N_3023);
nor U7079 (N_7079,N_4135,N_4338);
or U7080 (N_7080,N_2895,N_4529);
xnor U7081 (N_7081,N_4120,N_3429);
nor U7082 (N_7082,N_2610,N_3267);
nand U7083 (N_7083,N_3581,N_2729);
or U7084 (N_7084,N_2728,N_3064);
and U7085 (N_7085,N_3531,N_4506);
xnor U7086 (N_7086,N_2724,N_4976);
nor U7087 (N_7087,N_4844,N_3901);
and U7088 (N_7088,N_4316,N_4961);
nand U7089 (N_7089,N_4934,N_4384);
or U7090 (N_7090,N_3503,N_3960);
or U7091 (N_7091,N_4641,N_3950);
nand U7092 (N_7092,N_4014,N_3769);
nand U7093 (N_7093,N_3976,N_4072);
nand U7094 (N_7094,N_3596,N_3683);
nor U7095 (N_7095,N_3098,N_3238);
or U7096 (N_7096,N_4629,N_2980);
nand U7097 (N_7097,N_2986,N_2580);
or U7098 (N_7098,N_2571,N_3264);
and U7099 (N_7099,N_4992,N_3986);
nand U7100 (N_7100,N_3346,N_4515);
or U7101 (N_7101,N_2963,N_4141);
xnor U7102 (N_7102,N_4430,N_4477);
xnor U7103 (N_7103,N_3979,N_4032);
nand U7104 (N_7104,N_3651,N_4430);
or U7105 (N_7105,N_3172,N_4737);
and U7106 (N_7106,N_4132,N_3382);
and U7107 (N_7107,N_4395,N_4851);
nand U7108 (N_7108,N_2505,N_2807);
nor U7109 (N_7109,N_4573,N_4482);
and U7110 (N_7110,N_2557,N_4194);
nand U7111 (N_7111,N_3014,N_3438);
nand U7112 (N_7112,N_4173,N_2657);
xor U7113 (N_7113,N_4894,N_3593);
nand U7114 (N_7114,N_4977,N_4507);
nand U7115 (N_7115,N_3468,N_2953);
xnor U7116 (N_7116,N_2777,N_2735);
xor U7117 (N_7117,N_3645,N_3996);
xnor U7118 (N_7118,N_2756,N_3023);
nor U7119 (N_7119,N_3609,N_2917);
or U7120 (N_7120,N_3174,N_2599);
and U7121 (N_7121,N_4148,N_3572);
and U7122 (N_7122,N_2907,N_3093);
and U7123 (N_7123,N_4351,N_4525);
nor U7124 (N_7124,N_3428,N_3608);
xor U7125 (N_7125,N_4910,N_2863);
nand U7126 (N_7126,N_3862,N_4131);
xor U7127 (N_7127,N_4604,N_4183);
nor U7128 (N_7128,N_3576,N_3058);
or U7129 (N_7129,N_3997,N_4673);
nand U7130 (N_7130,N_4603,N_3415);
or U7131 (N_7131,N_4035,N_3902);
or U7132 (N_7132,N_3511,N_3599);
or U7133 (N_7133,N_2555,N_4609);
xnor U7134 (N_7134,N_2642,N_4852);
nor U7135 (N_7135,N_2915,N_3858);
or U7136 (N_7136,N_4143,N_4334);
xor U7137 (N_7137,N_4055,N_3792);
nor U7138 (N_7138,N_3765,N_3839);
nor U7139 (N_7139,N_4924,N_2827);
and U7140 (N_7140,N_4692,N_2963);
and U7141 (N_7141,N_2532,N_4309);
nand U7142 (N_7142,N_4569,N_3122);
nor U7143 (N_7143,N_4501,N_4596);
and U7144 (N_7144,N_4652,N_3028);
or U7145 (N_7145,N_4785,N_3947);
or U7146 (N_7146,N_4848,N_4867);
nor U7147 (N_7147,N_4691,N_3715);
nand U7148 (N_7148,N_3399,N_3769);
nand U7149 (N_7149,N_4814,N_2647);
or U7150 (N_7150,N_3745,N_3176);
or U7151 (N_7151,N_3654,N_4871);
nand U7152 (N_7152,N_3130,N_3016);
xor U7153 (N_7153,N_4342,N_3410);
and U7154 (N_7154,N_4551,N_3990);
or U7155 (N_7155,N_3020,N_3574);
nand U7156 (N_7156,N_2854,N_4784);
xor U7157 (N_7157,N_4799,N_2560);
and U7158 (N_7158,N_4493,N_4156);
xnor U7159 (N_7159,N_4414,N_2605);
or U7160 (N_7160,N_4017,N_2767);
and U7161 (N_7161,N_4020,N_3400);
nand U7162 (N_7162,N_3024,N_4118);
and U7163 (N_7163,N_4697,N_4552);
xnor U7164 (N_7164,N_3183,N_4827);
xnor U7165 (N_7165,N_2963,N_3879);
nor U7166 (N_7166,N_4223,N_4018);
nand U7167 (N_7167,N_3588,N_3650);
and U7168 (N_7168,N_2542,N_4108);
nor U7169 (N_7169,N_4638,N_4022);
xor U7170 (N_7170,N_3060,N_3886);
and U7171 (N_7171,N_4326,N_3349);
xnor U7172 (N_7172,N_4733,N_4275);
and U7173 (N_7173,N_4919,N_3859);
and U7174 (N_7174,N_2994,N_4771);
nor U7175 (N_7175,N_4704,N_3162);
nor U7176 (N_7176,N_3203,N_4806);
nor U7177 (N_7177,N_3275,N_2707);
and U7178 (N_7178,N_3159,N_3956);
or U7179 (N_7179,N_3809,N_3852);
nand U7180 (N_7180,N_3322,N_4576);
and U7181 (N_7181,N_4198,N_3747);
or U7182 (N_7182,N_4975,N_3240);
nor U7183 (N_7183,N_4718,N_4489);
nand U7184 (N_7184,N_4950,N_3903);
xor U7185 (N_7185,N_3448,N_3963);
xor U7186 (N_7186,N_3348,N_3327);
nor U7187 (N_7187,N_4525,N_4360);
nand U7188 (N_7188,N_2937,N_3156);
nor U7189 (N_7189,N_4420,N_4887);
xor U7190 (N_7190,N_4407,N_4502);
or U7191 (N_7191,N_4094,N_4883);
or U7192 (N_7192,N_3412,N_3163);
nor U7193 (N_7193,N_4932,N_4406);
and U7194 (N_7194,N_4430,N_4037);
or U7195 (N_7195,N_2984,N_2525);
nand U7196 (N_7196,N_3512,N_3905);
and U7197 (N_7197,N_3682,N_4269);
xor U7198 (N_7198,N_3621,N_2751);
xnor U7199 (N_7199,N_3957,N_2886);
or U7200 (N_7200,N_4855,N_3703);
nand U7201 (N_7201,N_4675,N_2968);
nand U7202 (N_7202,N_3225,N_4508);
nand U7203 (N_7203,N_2649,N_3111);
and U7204 (N_7204,N_3134,N_4400);
or U7205 (N_7205,N_3133,N_4981);
nand U7206 (N_7206,N_3687,N_4571);
nand U7207 (N_7207,N_3069,N_2860);
nand U7208 (N_7208,N_4808,N_2740);
nand U7209 (N_7209,N_4546,N_4136);
nand U7210 (N_7210,N_4683,N_4561);
nor U7211 (N_7211,N_4708,N_3210);
xnor U7212 (N_7212,N_3424,N_4685);
nor U7213 (N_7213,N_2659,N_3362);
and U7214 (N_7214,N_3753,N_4916);
or U7215 (N_7215,N_2654,N_4796);
xor U7216 (N_7216,N_4879,N_4101);
nand U7217 (N_7217,N_4467,N_4925);
nand U7218 (N_7218,N_2666,N_3595);
nor U7219 (N_7219,N_3960,N_4052);
nand U7220 (N_7220,N_3404,N_4944);
nand U7221 (N_7221,N_4413,N_4125);
and U7222 (N_7222,N_4594,N_3723);
or U7223 (N_7223,N_3052,N_4030);
or U7224 (N_7224,N_3438,N_3377);
or U7225 (N_7225,N_4175,N_4364);
nand U7226 (N_7226,N_3469,N_4471);
or U7227 (N_7227,N_2568,N_4221);
or U7228 (N_7228,N_3319,N_3434);
xor U7229 (N_7229,N_4673,N_2856);
nor U7230 (N_7230,N_3054,N_3533);
xnor U7231 (N_7231,N_4613,N_3594);
or U7232 (N_7232,N_4326,N_3628);
nand U7233 (N_7233,N_2806,N_3924);
and U7234 (N_7234,N_3795,N_3506);
nand U7235 (N_7235,N_4722,N_3374);
or U7236 (N_7236,N_4038,N_3285);
or U7237 (N_7237,N_2588,N_4964);
and U7238 (N_7238,N_2846,N_2853);
xnor U7239 (N_7239,N_4097,N_3925);
xnor U7240 (N_7240,N_2870,N_3866);
xnor U7241 (N_7241,N_2809,N_4067);
nor U7242 (N_7242,N_3741,N_3519);
xor U7243 (N_7243,N_4000,N_2577);
or U7244 (N_7244,N_3508,N_3975);
and U7245 (N_7245,N_4021,N_3711);
or U7246 (N_7246,N_4412,N_4359);
nand U7247 (N_7247,N_4078,N_3794);
nand U7248 (N_7248,N_2790,N_3929);
and U7249 (N_7249,N_4639,N_3626);
nand U7250 (N_7250,N_3519,N_3767);
xor U7251 (N_7251,N_2554,N_3491);
xor U7252 (N_7252,N_4053,N_3482);
xor U7253 (N_7253,N_4305,N_4499);
or U7254 (N_7254,N_2914,N_3820);
nor U7255 (N_7255,N_3931,N_4540);
nor U7256 (N_7256,N_2887,N_3975);
and U7257 (N_7257,N_2613,N_2716);
xor U7258 (N_7258,N_4828,N_3008);
xor U7259 (N_7259,N_3349,N_2900);
nor U7260 (N_7260,N_4073,N_4003);
and U7261 (N_7261,N_4929,N_4087);
xnor U7262 (N_7262,N_3541,N_4267);
nand U7263 (N_7263,N_3055,N_4955);
nor U7264 (N_7264,N_4225,N_3684);
or U7265 (N_7265,N_3540,N_3206);
or U7266 (N_7266,N_4016,N_2504);
or U7267 (N_7267,N_2965,N_4619);
nor U7268 (N_7268,N_3253,N_3927);
nand U7269 (N_7269,N_3721,N_4759);
xnor U7270 (N_7270,N_4181,N_4474);
nor U7271 (N_7271,N_2604,N_4041);
or U7272 (N_7272,N_3515,N_4673);
or U7273 (N_7273,N_2546,N_3479);
and U7274 (N_7274,N_2719,N_3100);
nor U7275 (N_7275,N_2692,N_3714);
or U7276 (N_7276,N_3804,N_4038);
xnor U7277 (N_7277,N_4592,N_3843);
or U7278 (N_7278,N_4886,N_2950);
nand U7279 (N_7279,N_3905,N_3499);
nor U7280 (N_7280,N_3624,N_3260);
nand U7281 (N_7281,N_3839,N_3520);
xnor U7282 (N_7282,N_4689,N_3053);
or U7283 (N_7283,N_4669,N_4456);
nor U7284 (N_7284,N_3394,N_3316);
or U7285 (N_7285,N_4483,N_3210);
nand U7286 (N_7286,N_2781,N_3334);
or U7287 (N_7287,N_2885,N_2796);
nand U7288 (N_7288,N_3369,N_4877);
or U7289 (N_7289,N_3495,N_4508);
and U7290 (N_7290,N_2658,N_3555);
or U7291 (N_7291,N_4389,N_4044);
or U7292 (N_7292,N_3613,N_4194);
xnor U7293 (N_7293,N_2976,N_3329);
nor U7294 (N_7294,N_2909,N_4599);
nor U7295 (N_7295,N_3737,N_4879);
nor U7296 (N_7296,N_3783,N_2611);
nand U7297 (N_7297,N_3113,N_4353);
and U7298 (N_7298,N_4028,N_3392);
nand U7299 (N_7299,N_3442,N_3312);
xnor U7300 (N_7300,N_3061,N_2803);
and U7301 (N_7301,N_3942,N_3863);
xor U7302 (N_7302,N_3045,N_2888);
and U7303 (N_7303,N_3488,N_3572);
nand U7304 (N_7304,N_3089,N_3670);
or U7305 (N_7305,N_2723,N_4744);
and U7306 (N_7306,N_4081,N_3176);
xor U7307 (N_7307,N_3547,N_3583);
nor U7308 (N_7308,N_3160,N_2670);
nand U7309 (N_7309,N_4514,N_4547);
nand U7310 (N_7310,N_4603,N_3368);
or U7311 (N_7311,N_4268,N_3692);
xor U7312 (N_7312,N_4840,N_2810);
xnor U7313 (N_7313,N_3819,N_3737);
nor U7314 (N_7314,N_2755,N_3302);
and U7315 (N_7315,N_4597,N_4655);
or U7316 (N_7316,N_3402,N_4814);
or U7317 (N_7317,N_3898,N_2557);
nor U7318 (N_7318,N_4008,N_4275);
nand U7319 (N_7319,N_3176,N_3640);
and U7320 (N_7320,N_2620,N_4952);
nor U7321 (N_7321,N_4823,N_3372);
nor U7322 (N_7322,N_3040,N_3441);
or U7323 (N_7323,N_4531,N_3128);
xnor U7324 (N_7324,N_2607,N_3840);
xor U7325 (N_7325,N_3511,N_4872);
nand U7326 (N_7326,N_4084,N_2906);
and U7327 (N_7327,N_3388,N_2685);
or U7328 (N_7328,N_3289,N_2626);
nand U7329 (N_7329,N_4016,N_4848);
and U7330 (N_7330,N_4733,N_3357);
or U7331 (N_7331,N_2896,N_4558);
or U7332 (N_7332,N_4307,N_2553);
nand U7333 (N_7333,N_3640,N_2764);
nand U7334 (N_7334,N_4979,N_3612);
or U7335 (N_7335,N_3969,N_4076);
nand U7336 (N_7336,N_2929,N_3187);
nand U7337 (N_7337,N_3457,N_4049);
and U7338 (N_7338,N_4054,N_4248);
xnor U7339 (N_7339,N_2778,N_3050);
and U7340 (N_7340,N_4928,N_2574);
nand U7341 (N_7341,N_2829,N_2993);
nor U7342 (N_7342,N_3181,N_4405);
xnor U7343 (N_7343,N_3874,N_3561);
and U7344 (N_7344,N_4123,N_3421);
nand U7345 (N_7345,N_3102,N_3334);
and U7346 (N_7346,N_4077,N_4007);
nand U7347 (N_7347,N_3004,N_4290);
nor U7348 (N_7348,N_4450,N_2944);
nand U7349 (N_7349,N_4965,N_2698);
or U7350 (N_7350,N_3211,N_4422);
nand U7351 (N_7351,N_4813,N_4092);
nor U7352 (N_7352,N_3742,N_4960);
nand U7353 (N_7353,N_2568,N_4062);
and U7354 (N_7354,N_3002,N_4513);
or U7355 (N_7355,N_3283,N_3431);
nand U7356 (N_7356,N_3816,N_2810);
or U7357 (N_7357,N_3493,N_3114);
or U7358 (N_7358,N_4471,N_4668);
and U7359 (N_7359,N_4675,N_2534);
and U7360 (N_7360,N_2908,N_4866);
nor U7361 (N_7361,N_4501,N_3645);
nor U7362 (N_7362,N_3383,N_4443);
nor U7363 (N_7363,N_3953,N_4830);
and U7364 (N_7364,N_4972,N_3488);
or U7365 (N_7365,N_4549,N_2569);
nor U7366 (N_7366,N_4725,N_2545);
xor U7367 (N_7367,N_2669,N_2747);
and U7368 (N_7368,N_2793,N_3505);
and U7369 (N_7369,N_4397,N_3049);
and U7370 (N_7370,N_4030,N_4700);
xnor U7371 (N_7371,N_4763,N_2839);
nand U7372 (N_7372,N_4575,N_3475);
and U7373 (N_7373,N_3996,N_4156);
and U7374 (N_7374,N_4333,N_4208);
nor U7375 (N_7375,N_3346,N_2809);
or U7376 (N_7376,N_3812,N_4102);
xor U7377 (N_7377,N_3978,N_2719);
nor U7378 (N_7378,N_3316,N_4670);
xnor U7379 (N_7379,N_3630,N_3368);
and U7380 (N_7380,N_2987,N_2712);
or U7381 (N_7381,N_4891,N_2541);
xor U7382 (N_7382,N_3985,N_2634);
and U7383 (N_7383,N_3978,N_3824);
xnor U7384 (N_7384,N_3454,N_3141);
nor U7385 (N_7385,N_2987,N_4793);
nor U7386 (N_7386,N_3556,N_4499);
nand U7387 (N_7387,N_3375,N_4584);
nand U7388 (N_7388,N_3015,N_4870);
nor U7389 (N_7389,N_2529,N_4903);
and U7390 (N_7390,N_3795,N_4160);
nor U7391 (N_7391,N_4589,N_3182);
nor U7392 (N_7392,N_3116,N_3183);
nor U7393 (N_7393,N_2680,N_4867);
nand U7394 (N_7394,N_2798,N_3433);
or U7395 (N_7395,N_4490,N_4768);
nand U7396 (N_7396,N_3805,N_4597);
or U7397 (N_7397,N_2941,N_4008);
or U7398 (N_7398,N_2804,N_4238);
or U7399 (N_7399,N_3944,N_3371);
or U7400 (N_7400,N_3117,N_4650);
and U7401 (N_7401,N_4466,N_2982);
and U7402 (N_7402,N_4949,N_3738);
or U7403 (N_7403,N_4590,N_2944);
nor U7404 (N_7404,N_3498,N_3789);
and U7405 (N_7405,N_2618,N_3274);
nor U7406 (N_7406,N_3203,N_2979);
xnor U7407 (N_7407,N_3486,N_3548);
and U7408 (N_7408,N_2818,N_4280);
nor U7409 (N_7409,N_3940,N_3961);
and U7410 (N_7410,N_3676,N_4447);
and U7411 (N_7411,N_3255,N_4514);
nor U7412 (N_7412,N_2575,N_4113);
or U7413 (N_7413,N_3832,N_3744);
or U7414 (N_7414,N_4734,N_4700);
nand U7415 (N_7415,N_4778,N_4256);
or U7416 (N_7416,N_3287,N_2836);
nor U7417 (N_7417,N_2758,N_4268);
or U7418 (N_7418,N_4813,N_3870);
or U7419 (N_7419,N_2868,N_4416);
nor U7420 (N_7420,N_2808,N_4371);
and U7421 (N_7421,N_4205,N_3847);
nand U7422 (N_7422,N_4926,N_3302);
and U7423 (N_7423,N_4417,N_3668);
or U7424 (N_7424,N_3038,N_4712);
xor U7425 (N_7425,N_2804,N_4741);
or U7426 (N_7426,N_3388,N_3666);
nor U7427 (N_7427,N_4210,N_3612);
nand U7428 (N_7428,N_4080,N_3966);
and U7429 (N_7429,N_4244,N_4541);
xnor U7430 (N_7430,N_2714,N_3958);
xor U7431 (N_7431,N_3993,N_4069);
and U7432 (N_7432,N_2690,N_3608);
or U7433 (N_7433,N_4836,N_4027);
nor U7434 (N_7434,N_4842,N_4733);
or U7435 (N_7435,N_4605,N_3719);
nand U7436 (N_7436,N_2759,N_4708);
or U7437 (N_7437,N_2794,N_3080);
and U7438 (N_7438,N_3182,N_3983);
xnor U7439 (N_7439,N_3053,N_4257);
xor U7440 (N_7440,N_3733,N_4009);
and U7441 (N_7441,N_4819,N_3047);
or U7442 (N_7442,N_2903,N_3177);
or U7443 (N_7443,N_4959,N_4090);
nor U7444 (N_7444,N_3752,N_3836);
or U7445 (N_7445,N_4444,N_4182);
nor U7446 (N_7446,N_2861,N_3238);
nor U7447 (N_7447,N_2819,N_4868);
nor U7448 (N_7448,N_4694,N_2799);
and U7449 (N_7449,N_2599,N_3122);
and U7450 (N_7450,N_2910,N_4358);
nor U7451 (N_7451,N_3152,N_3362);
nand U7452 (N_7452,N_2589,N_3870);
and U7453 (N_7453,N_3880,N_3885);
nor U7454 (N_7454,N_3107,N_3816);
nor U7455 (N_7455,N_4829,N_4416);
nand U7456 (N_7456,N_4828,N_2945);
nand U7457 (N_7457,N_3969,N_3096);
and U7458 (N_7458,N_2836,N_3529);
or U7459 (N_7459,N_4326,N_4562);
or U7460 (N_7460,N_2922,N_4413);
and U7461 (N_7461,N_4063,N_3942);
or U7462 (N_7462,N_2754,N_3338);
and U7463 (N_7463,N_4734,N_3863);
nand U7464 (N_7464,N_4795,N_2656);
and U7465 (N_7465,N_2556,N_3498);
or U7466 (N_7466,N_4992,N_3104);
nor U7467 (N_7467,N_3446,N_3363);
xnor U7468 (N_7468,N_3068,N_3724);
nand U7469 (N_7469,N_2914,N_2646);
or U7470 (N_7470,N_2930,N_4411);
or U7471 (N_7471,N_3498,N_3146);
or U7472 (N_7472,N_4582,N_2868);
nor U7473 (N_7473,N_4921,N_4691);
and U7474 (N_7474,N_3158,N_4429);
or U7475 (N_7475,N_3765,N_3588);
nor U7476 (N_7476,N_2767,N_3837);
and U7477 (N_7477,N_4385,N_4261);
xnor U7478 (N_7478,N_2914,N_3286);
nand U7479 (N_7479,N_2708,N_2729);
nor U7480 (N_7480,N_4957,N_2758);
nor U7481 (N_7481,N_3329,N_4928);
xor U7482 (N_7482,N_3737,N_3430);
or U7483 (N_7483,N_3034,N_3639);
nor U7484 (N_7484,N_3072,N_3895);
or U7485 (N_7485,N_3951,N_2879);
nand U7486 (N_7486,N_4250,N_4603);
nand U7487 (N_7487,N_3427,N_4165);
or U7488 (N_7488,N_3509,N_3174);
xnor U7489 (N_7489,N_2717,N_3964);
and U7490 (N_7490,N_4930,N_2603);
nor U7491 (N_7491,N_3067,N_3092);
nand U7492 (N_7492,N_4194,N_4433);
nor U7493 (N_7493,N_3036,N_3428);
nand U7494 (N_7494,N_4394,N_3443);
nand U7495 (N_7495,N_3840,N_3548);
or U7496 (N_7496,N_2891,N_4495);
nand U7497 (N_7497,N_3625,N_3842);
and U7498 (N_7498,N_2864,N_3761);
xor U7499 (N_7499,N_4070,N_3909);
xor U7500 (N_7500,N_7339,N_6957);
or U7501 (N_7501,N_6911,N_5418);
nor U7502 (N_7502,N_5527,N_5386);
or U7503 (N_7503,N_5822,N_7095);
and U7504 (N_7504,N_6536,N_6150);
or U7505 (N_7505,N_6787,N_5765);
or U7506 (N_7506,N_5035,N_5372);
nor U7507 (N_7507,N_6280,N_5284);
nor U7508 (N_7508,N_5040,N_5764);
and U7509 (N_7509,N_6522,N_6267);
xor U7510 (N_7510,N_7357,N_7069);
nor U7511 (N_7511,N_7465,N_5147);
or U7512 (N_7512,N_5006,N_5621);
xnor U7513 (N_7513,N_7403,N_7021);
xor U7514 (N_7514,N_5201,N_7077);
nor U7515 (N_7515,N_6240,N_6465);
nand U7516 (N_7516,N_6358,N_5573);
and U7517 (N_7517,N_6793,N_5547);
nor U7518 (N_7518,N_5519,N_6934);
nand U7519 (N_7519,N_6459,N_6158);
xnor U7520 (N_7520,N_6310,N_6112);
and U7521 (N_7521,N_7059,N_5458);
or U7522 (N_7522,N_6775,N_6281);
nor U7523 (N_7523,N_5802,N_6606);
or U7524 (N_7524,N_5106,N_5430);
nor U7525 (N_7525,N_7096,N_7409);
nor U7526 (N_7526,N_6173,N_7183);
nand U7527 (N_7527,N_6423,N_7483);
nand U7528 (N_7528,N_6469,N_7002);
nor U7529 (N_7529,N_7005,N_7224);
or U7530 (N_7530,N_6406,N_5989);
xor U7531 (N_7531,N_5339,N_5716);
or U7532 (N_7532,N_6984,N_7177);
nor U7533 (N_7533,N_6737,N_5560);
nand U7534 (N_7534,N_6869,N_5775);
nand U7535 (N_7535,N_6088,N_5363);
and U7536 (N_7536,N_6422,N_5615);
nand U7537 (N_7537,N_6391,N_6917);
or U7538 (N_7538,N_6786,N_7394);
nor U7539 (N_7539,N_5266,N_6343);
nand U7540 (N_7540,N_6962,N_5829);
nor U7541 (N_7541,N_7046,N_5361);
nand U7542 (N_7542,N_6543,N_7227);
nand U7543 (N_7543,N_6419,N_6026);
and U7544 (N_7544,N_6683,N_7105);
xor U7545 (N_7545,N_5279,N_5606);
and U7546 (N_7546,N_5323,N_5794);
or U7547 (N_7547,N_7340,N_5807);
or U7548 (N_7548,N_6130,N_5774);
nand U7549 (N_7549,N_5565,N_7225);
nand U7550 (N_7550,N_5821,N_7040);
xnor U7551 (N_7551,N_7487,N_7057);
nand U7552 (N_7552,N_6379,N_6621);
and U7553 (N_7553,N_5378,N_6724);
nor U7554 (N_7554,N_7335,N_5541);
nand U7555 (N_7555,N_6361,N_5157);
xnor U7556 (N_7556,N_5081,N_6043);
xnor U7557 (N_7557,N_6409,N_7391);
xor U7558 (N_7558,N_5028,N_6372);
and U7559 (N_7559,N_6766,N_5785);
nor U7560 (N_7560,N_5950,N_7172);
or U7561 (N_7561,N_6063,N_5089);
xor U7562 (N_7562,N_5653,N_7133);
or U7563 (N_7563,N_5311,N_6972);
and U7564 (N_7564,N_5970,N_5274);
or U7565 (N_7565,N_5000,N_7416);
nor U7566 (N_7566,N_7395,N_5701);
nor U7567 (N_7567,N_6930,N_6985);
nor U7568 (N_7568,N_7404,N_7139);
nand U7569 (N_7569,N_6609,N_6738);
nor U7570 (N_7570,N_5292,N_7384);
or U7571 (N_7571,N_6178,N_5150);
nor U7572 (N_7572,N_6181,N_7106);
or U7573 (N_7573,N_5195,N_7049);
and U7574 (N_7574,N_5796,N_7498);
nand U7575 (N_7575,N_6703,N_5733);
and U7576 (N_7576,N_6380,N_6908);
xor U7577 (N_7577,N_6124,N_5041);
xor U7578 (N_7578,N_6952,N_5884);
nor U7579 (N_7579,N_5877,N_5272);
nor U7580 (N_7580,N_5403,N_5443);
nor U7581 (N_7581,N_6454,N_6504);
xor U7582 (N_7582,N_5362,N_5095);
nand U7583 (N_7583,N_7157,N_5711);
xor U7584 (N_7584,N_5235,N_5026);
xnor U7585 (N_7585,N_6219,N_7162);
xor U7586 (N_7586,N_5102,N_6821);
or U7587 (N_7587,N_6212,N_6996);
and U7588 (N_7588,N_6861,N_5551);
nor U7589 (N_7589,N_6463,N_7109);
xnor U7590 (N_7590,N_6878,N_6691);
nor U7591 (N_7591,N_6264,N_7300);
and U7592 (N_7592,N_5782,N_5481);
nor U7593 (N_7593,N_6154,N_7126);
xnor U7594 (N_7594,N_6097,N_7292);
nand U7595 (N_7595,N_5897,N_7197);
and U7596 (N_7596,N_5426,N_7481);
nand U7597 (N_7597,N_7492,N_6300);
nand U7598 (N_7598,N_5015,N_6477);
xor U7599 (N_7599,N_5413,N_5182);
and U7600 (N_7600,N_7243,N_5841);
nand U7601 (N_7601,N_5024,N_6834);
and U7602 (N_7602,N_5538,N_5126);
nor U7603 (N_7603,N_5607,N_5114);
xnor U7604 (N_7604,N_6116,N_6244);
and U7605 (N_7605,N_7097,N_7150);
or U7606 (N_7606,N_5965,N_5952);
nor U7607 (N_7607,N_6374,N_5770);
xnor U7608 (N_7608,N_5159,N_6323);
nand U7609 (N_7609,N_6944,N_5183);
xor U7610 (N_7610,N_5524,N_6881);
nand U7611 (N_7611,N_5894,N_6656);
nand U7612 (N_7612,N_7050,N_6732);
and U7613 (N_7613,N_7115,N_6639);
or U7614 (N_7614,N_5377,N_7036);
nand U7615 (N_7615,N_6571,N_5668);
nor U7616 (N_7616,N_6809,N_6981);
nand U7617 (N_7617,N_7200,N_6798);
xor U7618 (N_7618,N_6049,N_6432);
or U7619 (N_7619,N_6791,N_5437);
nor U7620 (N_7620,N_5947,N_7155);
and U7621 (N_7621,N_5713,N_7202);
nand U7622 (N_7622,N_5127,N_5011);
nand U7623 (N_7623,N_7156,N_6236);
xnor U7624 (N_7624,N_5288,N_5973);
nand U7625 (N_7625,N_5188,N_5726);
nand U7626 (N_7626,N_6449,N_5872);
xnor U7627 (N_7627,N_6533,N_5725);
xnor U7628 (N_7628,N_6591,N_5493);
or U7629 (N_7629,N_6989,N_6964);
or U7630 (N_7630,N_6385,N_5883);
nor U7631 (N_7631,N_5083,N_6935);
or U7632 (N_7632,N_6000,N_6873);
nor U7633 (N_7633,N_5972,N_5073);
nand U7634 (N_7634,N_5500,N_6257);
and U7635 (N_7635,N_7470,N_7102);
nand U7636 (N_7636,N_7027,N_6252);
or U7637 (N_7637,N_5124,N_6362);
xor U7638 (N_7638,N_6176,N_5755);
and U7639 (N_7639,N_6393,N_5555);
or U7640 (N_7640,N_6092,N_5971);
or U7641 (N_7641,N_5482,N_5463);
xor U7642 (N_7642,N_6013,N_7039);
nand U7643 (N_7643,N_5173,N_5871);
nand U7644 (N_7644,N_5999,N_6851);
or U7645 (N_7645,N_6828,N_5979);
nor U7646 (N_7646,N_5345,N_6489);
or U7647 (N_7647,N_5036,N_6760);
nor U7648 (N_7648,N_5756,N_5044);
and U7649 (N_7649,N_5091,N_7163);
nor U7650 (N_7650,N_5938,N_7438);
nand U7651 (N_7651,N_6237,N_5140);
nor U7652 (N_7652,N_6666,N_5557);
nor U7653 (N_7653,N_7192,N_6995);
nand U7654 (N_7654,N_5179,N_7426);
nor U7655 (N_7655,N_5684,N_7071);
xnor U7656 (N_7656,N_5290,N_6965);
or U7657 (N_7657,N_5255,N_6673);
xnor U7658 (N_7658,N_7314,N_6705);
xnor U7659 (N_7659,N_6781,N_6942);
nor U7660 (N_7660,N_5594,N_5833);
xnor U7661 (N_7661,N_6839,N_7186);
or U7662 (N_7662,N_6577,N_6762);
nand U7663 (N_7663,N_6476,N_5241);
or U7664 (N_7664,N_6058,N_5793);
or U7665 (N_7665,N_7052,N_6331);
nor U7666 (N_7666,N_5869,N_5856);
nand U7667 (N_7667,N_5162,N_5257);
and U7668 (N_7668,N_5795,N_5452);
and U7669 (N_7669,N_5889,N_6761);
nor U7670 (N_7670,N_5580,N_7299);
and U7671 (N_7671,N_6458,N_7078);
and U7672 (N_7672,N_6527,N_6549);
or U7673 (N_7673,N_6135,N_5222);
nand U7674 (N_7674,N_5983,N_5561);
or U7675 (N_7675,N_6330,N_7390);
nand U7676 (N_7676,N_5310,N_6700);
nand U7677 (N_7677,N_6214,N_6569);
nor U7678 (N_7678,N_6084,N_6546);
nand U7679 (N_7679,N_7354,N_6484);
nor U7680 (N_7680,N_5549,N_6344);
nor U7681 (N_7681,N_6905,N_6923);
or U7682 (N_7682,N_7334,N_6731);
nand U7683 (N_7683,N_5881,N_6417);
xnor U7684 (N_7684,N_5910,N_7067);
or U7685 (N_7685,N_7215,N_6986);
xor U7686 (N_7686,N_5401,N_6364);
nand U7687 (N_7687,N_7003,N_7325);
nand U7688 (N_7688,N_7258,N_5819);
nand U7689 (N_7689,N_7331,N_5808);
or U7690 (N_7690,N_5639,N_6452);
and U7691 (N_7691,N_5342,N_5154);
and U7692 (N_7692,N_5583,N_6435);
xor U7693 (N_7693,N_5516,N_5596);
nor U7694 (N_7694,N_6799,N_7278);
xnor U7695 (N_7695,N_6065,N_6031);
and U7696 (N_7696,N_5766,N_7283);
nor U7697 (N_7697,N_6570,N_5824);
nor U7698 (N_7698,N_6721,N_5338);
or U7699 (N_7699,N_6959,N_6871);
or U7700 (N_7700,N_7297,N_5669);
and U7701 (N_7701,N_7124,N_5674);
xnor U7702 (N_7702,N_5364,N_7143);
or U7703 (N_7703,N_6014,N_7399);
and U7704 (N_7704,N_7076,N_6702);
and U7705 (N_7705,N_5525,N_5130);
xor U7706 (N_7706,N_5034,N_6366);
or U7707 (N_7707,N_6810,N_6245);
or U7708 (N_7708,N_6963,N_7087);
xor U7709 (N_7709,N_6061,N_6636);
xnor U7710 (N_7710,N_5908,N_7479);
nand U7711 (N_7711,N_5699,N_5744);
and U7712 (N_7712,N_5904,N_6638);
nor U7713 (N_7713,N_5077,N_5567);
nand U7714 (N_7714,N_5008,N_7495);
and U7715 (N_7715,N_7427,N_5681);
xor U7716 (N_7716,N_7301,N_5178);
or U7717 (N_7717,N_7337,N_7045);
xnor U7718 (N_7718,N_7174,N_6122);
or U7719 (N_7719,N_5597,N_5400);
nand U7720 (N_7720,N_7104,N_5902);
nor U7721 (N_7721,N_6497,N_5368);
xor U7722 (N_7722,N_6537,N_5906);
and U7723 (N_7723,N_5320,N_6982);
and U7724 (N_7724,N_6302,N_6101);
nor U7725 (N_7725,N_5104,N_5806);
nor U7726 (N_7726,N_5848,N_7457);
or U7727 (N_7727,N_7121,N_7132);
nand U7728 (N_7728,N_5205,N_5286);
or U7729 (N_7729,N_6168,N_7201);
and U7730 (N_7730,N_7113,N_5566);
and U7731 (N_7731,N_6988,N_5501);
or U7732 (N_7732,N_5319,N_6661);
nor U7733 (N_7733,N_5390,N_6282);
xnor U7734 (N_7734,N_6003,N_6676);
nand U7735 (N_7735,N_5704,N_6439);
or U7736 (N_7736,N_5369,N_7084);
and U7737 (N_7737,N_7273,N_6593);
xnor U7738 (N_7738,N_6770,N_7233);
nand U7739 (N_7739,N_6596,N_6508);
or U7740 (N_7740,N_6688,N_6747);
or U7741 (N_7741,N_6650,N_5995);
or U7742 (N_7742,N_7413,N_6410);
or U7743 (N_7743,N_7220,N_5540);
or U7744 (N_7744,N_5087,N_7148);
or U7745 (N_7745,N_7327,N_6713);
nand U7746 (N_7746,N_5991,N_5510);
xor U7747 (N_7747,N_7173,N_5629);
or U7748 (N_7748,N_7171,N_7305);
and U7749 (N_7749,N_5422,N_6309);
and U7750 (N_7750,N_6462,N_5259);
or U7751 (N_7751,N_6644,N_6874);
xor U7752 (N_7752,N_7100,N_5861);
nor U7753 (N_7753,N_5899,N_6826);
or U7754 (N_7754,N_5048,N_5291);
or U7755 (N_7755,N_6074,N_5090);
nand U7756 (N_7756,N_6495,N_6266);
and U7757 (N_7757,N_5414,N_7241);
nor U7758 (N_7758,N_7356,N_6017);
xnor U7759 (N_7759,N_6394,N_5903);
or U7760 (N_7760,N_5990,N_6233);
and U7761 (N_7761,N_7128,N_5027);
nor U7762 (N_7762,N_6011,N_5522);
or U7763 (N_7763,N_5085,N_6110);
or U7764 (N_7764,N_7452,N_7499);
nor U7765 (N_7765,N_5850,N_6890);
nor U7766 (N_7766,N_6475,N_6759);
nand U7767 (N_7767,N_5544,N_7254);
xor U7768 (N_7768,N_5843,N_5101);
xor U7769 (N_7769,N_5293,N_5626);
nand U7770 (N_7770,N_5062,N_5212);
nor U7771 (N_7771,N_5859,N_5504);
nand U7772 (N_7772,N_7017,N_5105);
nand U7773 (N_7773,N_6161,N_6649);
nor U7774 (N_7774,N_5542,N_7477);
and U7775 (N_7775,N_6304,N_6598);
nand U7776 (N_7776,N_5190,N_6792);
nor U7777 (N_7777,N_5691,N_5953);
and U7778 (N_7778,N_6451,N_5053);
or U7779 (N_7779,N_7070,N_6322);
or U7780 (N_7780,N_6044,N_6064);
nand U7781 (N_7781,N_6186,N_5732);
xnor U7782 (N_7782,N_5880,N_5010);
nand U7783 (N_7783,N_5218,N_6426);
xnor U7784 (N_7784,N_5853,N_5700);
or U7785 (N_7785,N_5449,N_6938);
nand U7786 (N_7786,N_5250,N_7206);
and U7787 (N_7787,N_6496,N_6633);
or U7788 (N_7788,N_5204,N_5605);
and U7789 (N_7789,N_5767,N_5845);
nand U7790 (N_7790,N_6992,N_7072);
and U7791 (N_7791,N_6107,N_7043);
nor U7792 (N_7792,N_6886,N_6371);
or U7793 (N_7793,N_6262,N_6892);
and U7794 (N_7794,N_6696,N_5247);
or U7795 (N_7795,N_7154,N_6473);
or U7796 (N_7796,N_6744,N_6728);
and U7797 (N_7797,N_6128,N_5627);
xor U7798 (N_7798,N_5748,N_6670);
and U7799 (N_7799,N_5060,N_5409);
nor U7800 (N_7800,N_7445,N_5484);
nand U7801 (N_7801,N_5340,N_5228);
and U7802 (N_7802,N_6194,N_6316);
nor U7803 (N_7803,N_6255,N_6751);
xor U7804 (N_7804,N_5118,N_6535);
or U7805 (N_7805,N_6788,N_6453);
nand U7806 (N_7806,N_7440,N_7336);
or U7807 (N_7807,N_5064,N_6815);
nor U7808 (N_7808,N_6845,N_7193);
nor U7809 (N_7809,N_5683,N_5349);
xnor U7810 (N_7810,N_7439,N_5391);
and U7811 (N_7811,N_6669,N_5882);
xor U7812 (N_7812,N_5509,N_6610);
nor U7813 (N_7813,N_7015,N_7242);
or U7814 (N_7814,N_6286,N_6009);
nor U7815 (N_7815,N_6727,N_5963);
nand U7816 (N_7816,N_6018,N_6875);
xnor U7817 (N_7817,N_5780,N_6270);
nand U7818 (N_7818,N_5745,N_6398);
nand U7819 (N_7819,N_5037,N_6937);
xor U7820 (N_7820,N_5968,N_6032);
and U7821 (N_7821,N_6632,N_5434);
nor U7822 (N_7822,N_5588,N_5838);
nand U7823 (N_7823,N_6405,N_5002);
xor U7824 (N_7824,N_7443,N_6441);
or U7825 (N_7825,N_6138,N_5453);
or U7826 (N_7826,N_5539,N_5176);
and U7827 (N_7827,N_6619,N_7235);
nand U7828 (N_7828,N_6408,N_6831);
xor U7829 (N_7829,N_5021,N_5811);
nor U7830 (N_7830,N_6540,N_5030);
xnor U7831 (N_7831,N_5718,N_6485);
and U7832 (N_7832,N_6162,N_5280);
or U7833 (N_7833,N_6929,N_5328);
nor U7834 (N_7834,N_6196,N_5165);
nand U7835 (N_7835,N_5086,N_6748);
and U7836 (N_7836,N_5689,N_5752);
and U7837 (N_7837,N_7451,N_5631);
nor U7838 (N_7838,N_7112,N_7246);
nor U7839 (N_7839,N_5348,N_5445);
xor U7840 (N_7840,N_6295,N_6040);
nor U7841 (N_7841,N_5231,N_5798);
nor U7842 (N_7842,N_5773,N_5728);
or U7843 (N_7843,N_5855,N_5758);
xnor U7844 (N_7844,N_7471,N_7135);
nand U7845 (N_7845,N_5265,N_6675);
or U7846 (N_7846,N_6631,N_7222);
nand U7847 (N_7847,N_5543,N_6444);
xnor U7848 (N_7848,N_5813,N_7152);
or U7849 (N_7849,N_7453,N_5474);
and U7850 (N_7850,N_7011,N_6824);
and U7851 (N_7851,N_5270,N_5107);
or U7852 (N_7852,N_6434,N_5723);
and U7853 (N_7853,N_5016,N_5506);
or U7854 (N_7854,N_6599,N_7127);
nand U7855 (N_7855,N_7031,N_5136);
or U7856 (N_7856,N_5680,N_6618);
nand U7857 (N_7857,N_5628,N_7294);
xnor U7858 (N_7858,N_5405,N_5554);
or U7859 (N_7859,N_6265,N_6884);
nor U7860 (N_7860,N_6857,N_6805);
or U7861 (N_7861,N_6657,N_5558);
xnor U7862 (N_7862,N_5407,N_7265);
and U7863 (N_7863,N_6318,N_6447);
xnor U7864 (N_7864,N_6115,N_5071);
xnor U7865 (N_7865,N_7355,N_6012);
nor U7866 (N_7866,N_6250,N_5520);
and U7867 (N_7867,N_5526,N_6397);
nand U7868 (N_7868,N_7238,N_6248);
nand U7869 (N_7869,N_6498,N_5170);
xor U7870 (N_7870,N_5616,N_7352);
nor U7871 (N_7871,N_5960,N_5185);
nor U7872 (N_7872,N_5302,N_7181);
or U7873 (N_7873,N_6321,N_5110);
xnor U7874 (N_7874,N_5214,N_6575);
and U7875 (N_7875,N_6922,N_6967);
and U7876 (N_7876,N_6741,N_6224);
or U7877 (N_7877,N_5641,N_6600);
and U7878 (N_7878,N_5447,N_5707);
nand U7879 (N_7879,N_6420,N_5221);
and U7880 (N_7880,N_5797,N_6464);
and U7881 (N_7881,N_6089,N_7080);
or U7882 (N_7882,N_7144,N_6622);
nand U7883 (N_7883,N_6943,N_5617);
nand U7884 (N_7884,N_7288,N_6174);
or U7885 (N_7885,N_6842,N_5951);
nand U7886 (N_7886,N_5982,N_5134);
nor U7887 (N_7887,N_6156,N_6139);
xnor U7888 (N_7888,N_7016,N_5371);
xnor U7889 (N_7889,N_6818,N_6830);
and U7890 (N_7890,N_6594,N_6348);
or U7891 (N_7891,N_5262,N_5005);
xnor U7892 (N_7892,N_6991,N_6927);
nand U7893 (N_7893,N_5876,N_6332);
nand U7894 (N_7894,N_6872,N_5624);
xnor U7895 (N_7895,N_6777,N_6865);
xnor U7896 (N_7896,N_5387,N_5258);
xor U7897 (N_7897,N_7211,N_5942);
nor U7898 (N_7898,N_7311,N_6079);
nand U7899 (N_7899,N_7410,N_6580);
xnor U7900 (N_7900,N_5158,N_6977);
nor U7901 (N_7901,N_5977,N_6141);
or U7902 (N_7902,N_7063,N_5113);
nand U7903 (N_7903,N_6529,N_6234);
nor U7904 (N_7904,N_7038,N_5849);
nor U7905 (N_7905,N_6076,N_5578);
xor U7906 (N_7906,N_5503,N_7260);
xnor U7907 (N_7907,N_6137,N_6376);
nand U7908 (N_7908,N_6823,N_7262);
or U7909 (N_7909,N_6293,N_5264);
xor U7910 (N_7910,N_5657,N_6229);
xnor U7911 (N_7911,N_6785,N_6333);
xnor U7912 (N_7912,N_5237,N_5393);
xor U7913 (N_7913,N_5847,N_6514);
or U7914 (N_7914,N_5936,N_7058);
nand U7915 (N_7915,N_5532,N_5827);
and U7916 (N_7916,N_7175,N_6171);
and U7917 (N_7917,N_6634,N_7091);
nand U7918 (N_7918,N_7359,N_6701);
nor U7919 (N_7919,N_5357,N_7368);
and U7920 (N_7920,N_5436,N_5772);
or U7921 (N_7921,N_6072,N_6756);
and U7922 (N_7922,N_5779,N_6307);
nand U7923 (N_7923,N_5103,N_7079);
and U7924 (N_7924,N_5433,N_6932);
nand U7925 (N_7925,N_5329,N_5866);
and U7926 (N_7926,N_5751,N_5945);
or U7927 (N_7927,N_5455,N_5491);
or U7928 (N_7928,N_7264,N_6687);
and U7929 (N_7929,N_7217,N_6170);
nor U7930 (N_7930,N_7460,N_7130);
nor U7931 (N_7931,N_7195,N_5314);
nand U7932 (N_7932,N_6651,N_6941);
xnor U7933 (N_7933,N_5595,N_5946);
nand U7934 (N_7934,N_5664,N_6544);
or U7935 (N_7935,N_6354,N_5603);
xnor U7936 (N_7936,N_7051,N_7406);
and U7937 (N_7937,N_6471,N_7034);
nor U7938 (N_7938,N_5384,N_6149);
xnor U7939 (N_7939,N_6764,N_6263);
nor U7940 (N_7940,N_7248,N_5408);
and U7941 (N_7941,N_5613,N_7494);
xnor U7942 (N_7942,N_7309,N_7270);
xnor U7943 (N_7943,N_5740,N_5069);
nand U7944 (N_7944,N_7145,N_6203);
xnor U7945 (N_7945,N_6512,N_5287);
xnor U7946 (N_7946,N_7044,N_6743);
xnor U7947 (N_7947,N_6502,N_6613);
nor U7948 (N_7948,N_5789,N_5692);
xnor U7949 (N_7949,N_6069,N_5269);
xor U7950 (N_7950,N_7207,N_5198);
or U7951 (N_7951,N_6381,N_5275);
and U7952 (N_7952,N_6518,N_6106);
nand U7953 (N_7953,N_7298,N_6384);
nand U7954 (N_7954,N_6734,N_5225);
nor U7955 (N_7955,N_6730,N_7179);
nand U7956 (N_7956,N_6841,N_6152);
nor U7957 (N_7957,N_7407,N_6166);
nand U7958 (N_7958,N_6146,N_6838);
nand U7959 (N_7959,N_6228,N_6284);
nand U7960 (N_7960,N_6733,N_5985);
nor U7961 (N_7961,N_6660,N_7255);
and U7962 (N_7962,N_5410,N_6225);
and U7963 (N_7963,N_7366,N_5515);
or U7964 (N_7964,N_5251,N_6635);
or U7965 (N_7965,N_7023,N_7324);
nor U7966 (N_7966,N_7424,N_5213);
or U7967 (N_7967,N_6442,N_6885);
nor U7968 (N_7968,N_6617,N_5380);
and U7969 (N_7969,N_5809,N_7414);
nand U7970 (N_7970,N_6902,N_6652);
and U7971 (N_7971,N_6576,N_6859);
xnor U7972 (N_7972,N_6772,N_5754);
or U7973 (N_7973,N_7019,N_7188);
nor U7974 (N_7974,N_6356,N_5875);
or U7975 (N_7975,N_6913,N_5318);
or U7976 (N_7976,N_6033,N_6668);
nand U7977 (N_7977,N_5623,N_7054);
nand U7978 (N_7978,N_7386,N_5042);
or U7979 (N_7979,N_5887,N_6388);
or U7980 (N_7980,N_5720,N_6352);
and U7981 (N_7981,N_7437,N_7330);
xor U7982 (N_7982,N_7475,N_5858);
and U7983 (N_7983,N_7371,N_7468);
or U7984 (N_7984,N_5163,N_7376);
or U7985 (N_7985,N_5283,N_6445);
xnor U7986 (N_7986,N_6093,N_7486);
nand U7987 (N_7987,N_6239,N_6840);
and U7988 (N_7988,N_6648,N_7007);
nand U7989 (N_7989,N_6221,N_7401);
nand U7990 (N_7990,N_6412,N_5457);
nor U7991 (N_7991,N_7285,N_5343);
and U7992 (N_7992,N_5020,N_6305);
or U7993 (N_7993,N_5781,N_5486);
nand U7994 (N_7994,N_6769,N_6456);
xnor U7995 (N_7995,N_7377,N_6200);
nor U7996 (N_7996,N_6707,N_5468);
or U7997 (N_7997,N_5098,N_6062);
xor U7998 (N_7998,N_5898,N_5996);
or U7999 (N_7999,N_6578,N_5708);
or U8000 (N_8000,N_5659,N_6287);
nor U8001 (N_8001,N_6720,N_6742);
xnor U8002 (N_8002,N_5135,N_6400);
nand U8003 (N_8003,N_5216,N_5976);
or U8004 (N_8004,N_5529,N_6005);
or U8005 (N_8005,N_6862,N_6500);
and U8006 (N_8006,N_7397,N_5890);
nor U8007 (N_8007,N_6446,N_6365);
and U8008 (N_8008,N_5675,N_6901);
and U8009 (N_8009,N_6187,N_6349);
or U8010 (N_8010,N_6164,N_7466);
nor U8011 (N_8011,N_5927,N_5874);
or U8012 (N_8012,N_7062,N_5645);
xnor U8013 (N_8013,N_6247,N_6133);
and U8014 (N_8014,N_6948,N_6794);
nor U8015 (N_8015,N_5734,N_7431);
or U8016 (N_8016,N_6218,N_5572);
and U8017 (N_8017,N_6946,N_5075);
and U8018 (N_8018,N_6411,N_6931);
or U8019 (N_8019,N_5686,N_6836);
or U8020 (N_8020,N_6641,N_6290);
nand U8021 (N_8021,N_6757,N_5050);
or U8022 (N_8022,N_6746,N_7214);
nand U8023 (N_8023,N_6867,N_5909);
and U8024 (N_8024,N_7293,N_6501);
nor U8025 (N_8025,N_7061,N_5488);
and U8026 (N_8026,N_6887,N_5394);
or U8027 (N_8027,N_7166,N_5496);
nand U8028 (N_8028,N_5419,N_6177);
nor U8029 (N_8029,N_5648,N_6515);
nand U8030 (N_8030,N_5305,N_6564);
and U8031 (N_8031,N_5167,N_7275);
nand U8032 (N_8032,N_5724,N_5007);
xnor U8033 (N_8033,N_5495,N_6087);
nor U8034 (N_8034,N_5148,N_6679);
xor U8035 (N_8035,N_6197,N_5633);
xor U8036 (N_8036,N_6396,N_5814);
and U8037 (N_8037,N_6383,N_5844);
nand U8038 (N_8038,N_6987,N_6753);
and U8039 (N_8039,N_7244,N_5592);
nand U8040 (N_8040,N_7488,N_6157);
xor U8041 (N_8041,N_5851,N_7204);
nor U8042 (N_8042,N_6480,N_6847);
and U8043 (N_8043,N_6370,N_5416);
xnor U8044 (N_8044,N_6118,N_5642);
nor U8045 (N_8045,N_5132,N_6472);
or U8046 (N_8046,N_5579,N_6949);
nor U8047 (N_8047,N_6517,N_6466);
nor U8048 (N_8048,N_6123,N_6363);
nand U8049 (N_8049,N_5261,N_7239);
nand U8050 (N_8050,N_5835,N_6888);
xnor U8051 (N_8051,N_6373,N_5825);
and U8052 (N_8052,N_6883,N_5052);
and U8053 (N_8053,N_5959,N_5489);
nor U8054 (N_8054,N_5878,N_7212);
and U8055 (N_8055,N_5556,N_6401);
and U8056 (N_8056,N_5072,N_5230);
nor U8057 (N_8057,N_6994,N_6910);
nor U8058 (N_8058,N_5029,N_7205);
and U8059 (N_8059,N_5476,N_6208);
nand U8060 (N_8060,N_7075,N_5873);
nor U8061 (N_8061,N_6776,N_5444);
or U8062 (N_8062,N_5256,N_6783);
xnor U8063 (N_8063,N_6595,N_5316);
nor U8064 (N_8064,N_6531,N_6275);
or U8065 (N_8065,N_5161,N_7229);
nor U8066 (N_8066,N_6022,N_5354);
and U8067 (N_8067,N_6210,N_6928);
xor U8068 (N_8068,N_6042,N_5771);
nand U8069 (N_8069,N_5575,N_5964);
nand U8070 (N_8070,N_7253,N_5593);
nand U8071 (N_8071,N_5171,N_5079);
nor U8072 (N_8072,N_5406,N_5992);
or U8073 (N_8073,N_6201,N_6329);
nor U8074 (N_8074,N_6804,N_5145);
or U8075 (N_8075,N_5988,N_6202);
xnor U8076 (N_8076,N_6592,N_7348);
nor U8077 (N_8077,N_7456,N_5905);
or U8078 (N_8078,N_7194,N_7251);
xor U8079 (N_8079,N_6519,N_5344);
and U8080 (N_8080,N_6626,N_6440);
nor U8081 (N_8081,N_6966,N_5223);
or U8082 (N_8082,N_6722,N_7421);
and U8083 (N_8083,N_6429,N_6037);
or U8084 (N_8084,N_5385,N_7108);
nor U8085 (N_8085,N_6739,N_5581);
and U8086 (N_8086,N_6460,N_5059);
and U8087 (N_8087,N_6817,N_5321);
or U8088 (N_8088,N_7074,N_6803);
and U8089 (N_8089,N_5012,N_6029);
or U8090 (N_8090,N_5512,N_6630);
nand U8091 (N_8091,N_6481,N_5969);
or U8092 (N_8092,N_5207,N_5402);
xnor U8093 (N_8093,N_7497,N_6856);
xnor U8094 (N_8094,N_5099,N_5049);
nor U8095 (N_8095,N_7322,N_5168);
or U8096 (N_8096,N_7482,N_5017);
or U8097 (N_8097,N_6876,N_6357);
xor U8098 (N_8098,N_7382,N_5987);
and U8099 (N_8099,N_6800,N_5762);
and U8100 (N_8100,N_5424,N_6308);
or U8101 (N_8101,N_5638,N_7372);
and U8102 (N_8102,N_5472,N_6893);
nor U8103 (N_8103,N_5651,N_5826);
nand U8104 (N_8104,N_7138,N_6709);
xnor U8105 (N_8105,N_6552,N_5559);
xnor U8106 (N_8106,N_7240,N_7169);
or U8107 (N_8107,N_6132,N_5398);
xnor U8108 (N_8108,N_7442,N_5252);
or U8109 (N_8109,N_7053,N_5867);
or U8110 (N_8110,N_7218,N_6023);
xnor U8111 (N_8111,N_6136,N_6808);
nand U8112 (N_8112,N_6706,N_7389);
xnor U8113 (N_8113,N_5285,N_6736);
xor U8114 (N_8114,N_5295,N_6021);
nor U8115 (N_8115,N_5388,N_5730);
nand U8116 (N_8116,N_6665,N_5562);
or U8117 (N_8117,N_5018,N_6274);
or U8118 (N_8118,N_5705,N_7103);
or U8119 (N_8119,N_5854,N_5661);
and U8120 (N_8120,N_5932,N_6833);
nand U8121 (N_8121,N_6520,N_6227);
and U8122 (N_8122,N_6814,N_6377);
nor U8123 (N_8123,N_6620,N_6353);
xor U8124 (N_8124,N_6507,N_5397);
nand U8125 (N_8125,N_6159,N_5092);
nor U8126 (N_8126,N_6616,N_5485);
nand U8127 (N_8127,N_6041,N_6754);
nand U8128 (N_8128,N_6970,N_6277);
nand U8129 (N_8129,N_7158,N_6582);
nand U8130 (N_8130,N_6853,N_5141);
nand U8131 (N_8131,N_5076,N_6085);
or U8132 (N_8132,N_6147,N_6470);
and U8133 (N_8133,N_6796,N_6850);
nand U8134 (N_8134,N_7117,N_5533);
nor U8135 (N_8135,N_5706,N_5537);
or U8136 (N_8136,N_7234,N_5656);
nand U8137 (N_8137,N_5840,N_7493);
nand U8138 (N_8138,N_5703,N_5548);
or U8139 (N_8139,N_7259,N_7333);
xor U8140 (N_8140,N_6933,N_7055);
nor U8141 (N_8141,N_5260,N_6723);
nor U8142 (N_8142,N_6016,N_6712);
xnor U8143 (N_8143,N_7013,N_6539);
nand U8144 (N_8144,N_7435,N_5379);
and U8145 (N_8145,N_6692,N_5784);
nor U8146 (N_8146,N_7307,N_6837);
nand U8147 (N_8147,N_6950,N_5837);
or U8148 (N_8148,N_7026,N_5690);
and U8149 (N_8149,N_7373,N_5175);
or U8150 (N_8150,N_6051,N_7170);
and U8151 (N_8151,N_5004,N_7245);
and U8152 (N_8152,N_6193,N_5722);
xor U8153 (N_8153,N_6068,N_5038);
or U8154 (N_8154,N_6572,N_6898);
and U8155 (N_8155,N_7073,N_6002);
and U8156 (N_8156,N_7092,N_5925);
nor U8157 (N_8157,N_7000,N_5186);
nor U8158 (N_8158,N_5478,N_6778);
nor U8159 (N_8159,N_6414,N_6672);
or U8160 (N_8160,N_5498,N_5879);
nand U8161 (N_8161,N_7393,N_6345);
nand U8162 (N_8162,N_7164,N_5142);
nand U8163 (N_8163,N_5067,N_6030);
nor U8164 (N_8164,N_7107,N_5777);
xor U8165 (N_8165,N_6958,N_6378);
or U8166 (N_8166,N_5741,N_6153);
and U8167 (N_8167,N_5993,N_6513);
xnor U8168 (N_8168,N_6008,N_5299);
or U8169 (N_8169,N_7455,N_5660);
nor U8170 (N_8170,N_5523,N_6235);
xor U8171 (N_8171,N_5521,N_7088);
xor U8172 (N_8172,N_7037,N_5846);
nor U8173 (N_8173,N_7361,N_5227);
nor U8174 (N_8174,N_5460,N_7447);
or U8175 (N_8175,N_6046,N_6455);
nor U8176 (N_8176,N_5296,N_6057);
nand U8177 (N_8177,N_6647,N_7210);
nor U8178 (N_8178,N_6690,N_5045);
nand U8179 (N_8179,N_7196,N_5914);
xor U8180 (N_8180,N_5490,N_5475);
nor U8181 (N_8181,N_7304,N_6954);
xor U8182 (N_8182,N_6603,N_5749);
nor U8183 (N_8183,N_5614,N_6827);
or U8184 (N_8184,N_5330,N_5715);
and U8185 (N_8185,N_5350,N_5803);
xnor U8186 (N_8186,N_6269,N_5451);
nand U8187 (N_8187,N_5696,N_5374);
xor U8188 (N_8188,N_5376,N_7125);
xnor U8189 (N_8189,N_7370,N_6565);
xnor U8190 (N_8190,N_6169,N_7484);
and U8191 (N_8191,N_5483,N_6198);
xor U8192 (N_8192,N_7449,N_5612);
nand U8193 (N_8193,N_7462,N_5602);
and U8194 (N_8194,N_6749,N_5276);
or U8195 (N_8195,N_6907,N_5820);
nand U8196 (N_8196,N_5074,N_5719);
nand U8197 (N_8197,N_6983,N_5600);
xor U8198 (N_8198,N_6278,N_5934);
and U8199 (N_8199,N_6294,N_6433);
nand U8200 (N_8200,N_6524,N_6541);
or U8201 (N_8201,N_6961,N_5980);
nand U8202 (N_8202,N_5676,N_5438);
or U8203 (N_8203,N_7478,N_6007);
and U8204 (N_8204,N_5115,N_7185);
xnor U8205 (N_8205,N_5601,N_7180);
xnor U8206 (N_8206,N_6750,N_5459);
xnor U8207 (N_8207,N_6849,N_5944);
nand U8208 (N_8208,N_6896,N_7141);
and U8209 (N_8209,N_6425,N_5816);
or U8210 (N_8210,N_5189,N_6211);
nor U8211 (N_8211,N_5571,N_7398);
nand U8212 (N_8212,N_5063,N_5435);
nor U8213 (N_8213,N_6735,N_5263);
and U8214 (N_8214,N_6367,N_6492);
and U8215 (N_8215,N_5078,N_6682);
nand U8216 (N_8216,N_6254,N_5439);
or U8217 (N_8217,N_6226,N_5324);
nand U8218 (N_8218,N_6758,N_6297);
and U8219 (N_8219,N_5334,N_6605);
and U8220 (N_8220,N_5149,N_6067);
and U8221 (N_8221,N_5193,N_5267);
and U8222 (N_8222,N_6131,N_6960);
xnor U8223 (N_8223,N_6327,N_6075);
nand U8224 (N_8224,N_7068,N_5180);
or U8225 (N_8225,N_6677,N_6468);
and U8226 (N_8226,N_6109,N_5432);
or U8227 (N_8227,N_6587,N_5800);
and U8228 (N_8228,N_6574,N_5497);
nor U8229 (N_8229,N_6590,N_6926);
nor U8230 (N_8230,N_5832,N_5986);
or U8231 (N_8231,N_5761,N_6844);
nor U8232 (N_8232,N_5836,N_5392);
nor U8233 (N_8233,N_7380,N_5598);
nand U8234 (N_8234,N_7433,N_5860);
xor U8235 (N_8235,N_5308,N_6479);
nor U8236 (N_8236,N_7146,N_6010);
and U8237 (N_8237,N_5033,N_6253);
xor U8238 (N_8238,N_6272,N_5121);
and U8239 (N_8239,N_5300,N_5957);
or U8240 (N_8240,N_5919,N_6404);
nand U8241 (N_8241,N_6779,N_6506);
nand U8242 (N_8242,N_6711,N_6190);
or U8243 (N_8243,N_7085,N_7230);
nand U8244 (N_8244,N_6978,N_6335);
xnor U8245 (N_8245,N_6209,N_5961);
xor U8246 (N_8246,N_7441,N_6082);
or U8247 (N_8247,N_5799,N_6407);
and U8248 (N_8248,N_6102,N_7346);
and U8249 (N_8249,N_5610,N_5673);
or U8250 (N_8250,N_7110,N_5151);
or U8251 (N_8251,N_6006,N_7247);
or U8252 (N_8252,N_6117,N_7066);
xnor U8253 (N_8253,N_7415,N_5446);
nand U8254 (N_8254,N_6768,N_5922);
or U8255 (N_8255,N_6241,N_6914);
nand U8256 (N_8256,N_6588,N_6563);
nor U8257 (N_8257,N_6585,N_5536);
xor U8258 (N_8258,N_5238,N_6001);
nand U8259 (N_8259,N_5070,N_7279);
or U8260 (N_8260,N_5479,N_5590);
nand U8261 (N_8261,N_7033,N_6581);
or U8262 (N_8262,N_6607,N_5834);
xor U8263 (N_8263,N_5412,N_5923);
xnor U8264 (N_8264,N_7228,N_6103);
and U8265 (N_8265,N_6100,N_7317);
xor U8266 (N_8266,N_5643,N_5298);
xnor U8267 (N_8267,N_6567,N_6184);
nor U8268 (N_8268,N_5939,N_5146);
nor U8269 (N_8269,N_6078,N_7290);
xor U8270 (N_8270,N_5688,N_7250);
and U8271 (N_8271,N_6795,N_5665);
and U8272 (N_8272,N_6387,N_5322);
nand U8273 (N_8273,N_6431,N_5892);
or U8274 (N_8274,N_5122,N_6763);
xor U8275 (N_8275,N_5842,N_5695);
xor U8276 (N_8276,N_6806,N_5552);
nand U8277 (N_8277,N_6077,N_5649);
nand U8278 (N_8278,N_7216,N_7014);
or U8279 (N_8279,N_5710,N_6645);
nor U8280 (N_8280,N_5156,N_6860);
nand U8281 (N_8281,N_5619,N_5599);
and U8282 (N_8282,N_6719,N_7009);
nand U8283 (N_8283,N_5046,N_5172);
and U8284 (N_8284,N_5367,N_5918);
xnor U8285 (N_8285,N_6276,N_6579);
xor U8286 (N_8286,N_7412,N_7360);
or U8287 (N_8287,N_6443,N_5355);
and U8288 (N_8288,N_6879,N_5513);
xor U8289 (N_8289,N_5309,N_6491);
nor U8290 (N_8290,N_5065,N_5634);
nand U8291 (N_8291,N_6899,N_6525);
nor U8292 (N_8292,N_6053,N_6654);
and U8293 (N_8293,N_6637,N_7149);
and U8294 (N_8294,N_7098,N_6698);
and U8295 (N_8295,N_5191,N_5428);
nand U8296 (N_8296,N_6843,N_5791);
or U8297 (N_8297,N_5546,N_7090);
and U8298 (N_8298,N_7010,N_5924);
xor U8299 (N_8299,N_5219,N_5911);
and U8300 (N_8300,N_7190,N_7184);
or U8301 (N_8301,N_5112,N_7168);
xnor U8302 (N_8302,N_7161,N_5211);
xor U8303 (N_8303,N_7295,N_6142);
and U8304 (N_8304,N_7364,N_6125);
xor U8305 (N_8305,N_5307,N_7089);
nand U8306 (N_8306,N_5857,N_7064);
xnor U8307 (N_8307,N_6615,N_6625);
and U8308 (N_8308,N_5194,N_6306);
or U8309 (N_8309,N_5125,N_5032);
nor U8310 (N_8310,N_5014,N_6428);
and U8311 (N_8311,N_5731,N_5531);
and U8312 (N_8312,N_6399,N_7029);
and U8313 (N_8313,N_5133,N_5404);
xnor U8314 (N_8314,N_6882,N_5013);
nand U8315 (N_8315,N_5082,N_6035);
nand U8316 (N_8316,N_5277,N_6919);
nor U8317 (N_8317,N_7223,N_5312);
or U8318 (N_8318,N_6185,N_5094);
or U8319 (N_8319,N_6557,N_7056);
or U8320 (N_8320,N_5088,N_5577);
or U8321 (N_8321,N_7136,N_7402);
nor U8322 (N_8322,N_6643,N_5757);
and U8323 (N_8323,N_5815,N_6897);
or U8324 (N_8324,N_7342,N_6059);
xor U8325 (N_8325,N_5123,N_5518);
nor U8326 (N_8326,N_6558,N_6217);
xnor U8327 (N_8327,N_6313,N_6182);
and U8328 (N_8328,N_5553,N_5574);
or U8329 (N_8329,N_6510,N_6490);
xnor U8330 (N_8330,N_6347,N_7400);
and U8331 (N_8331,N_5019,N_6646);
xor U8332 (N_8332,N_6993,N_7282);
xnor U8333 (N_8333,N_6191,N_7329);
nand U8334 (N_8334,N_6261,N_7365);
or U8335 (N_8335,N_7199,N_5177);
or U8336 (N_8336,N_7022,N_6355);
and U8337 (N_8337,N_5215,N_5271);
nand U8338 (N_8338,N_5442,N_5862);
xnor U8339 (N_8339,N_5181,N_5931);
and U8340 (N_8340,N_5584,N_5786);
xor U8341 (N_8341,N_7159,N_6099);
and U8342 (N_8342,N_7319,N_5470);
nor U8343 (N_8343,N_6979,N_7035);
or U8344 (N_8344,N_6945,N_5679);
or U8345 (N_8345,N_5166,N_6108);
nor U8346 (N_8346,N_6568,N_6258);
nor U8347 (N_8347,N_6566,N_6390);
xor U8348 (N_8348,N_5499,N_5739);
or U8349 (N_8349,N_6807,N_7142);
xnor U8350 (N_8350,N_7047,N_6678);
and U8351 (N_8351,N_5534,N_6608);
or U8352 (N_8352,N_6601,N_5507);
nor U8353 (N_8353,N_6526,N_7418);
nor U8354 (N_8354,N_6482,N_6105);
and U8355 (N_8355,N_6395,N_6542);
or U8356 (N_8356,N_5929,N_5916);
xnor U8357 (N_8357,N_6767,N_6725);
nand U8358 (N_8358,N_7464,N_6314);
and U8359 (N_8359,N_5431,N_5196);
and U8360 (N_8360,N_5100,N_7392);
or U8361 (N_8361,N_5801,N_5254);
and U8362 (N_8362,N_6315,N_6789);
and U8363 (N_8363,N_6642,N_6812);
nand U8364 (N_8364,N_5888,N_7048);
nor U8365 (N_8365,N_6392,N_7165);
or U8366 (N_8366,N_7266,N_6811);
and U8367 (N_8367,N_7160,N_5365);
nand U8368 (N_8368,N_5128,N_5356);
nand U8369 (N_8369,N_7151,N_7345);
or U8370 (N_8370,N_7018,N_5545);
nand U8371 (N_8371,N_5672,N_5440);
xor U8372 (N_8372,N_6998,N_5473);
and U8373 (N_8373,N_6004,N_7208);
nand U8374 (N_8374,N_7344,N_6195);
and U8375 (N_8375,N_7463,N_5487);
nor U8376 (N_8376,N_5640,N_6303);
or U8377 (N_8377,N_6402,N_6288);
or U8378 (N_8378,N_5303,N_7476);
nand U8379 (N_8379,N_6699,N_5187);
xnor U8380 (N_8380,N_5921,N_7320);
and U8381 (N_8381,N_6337,N_7182);
nor U8382 (N_8382,N_6726,N_6095);
or U8383 (N_8383,N_5327,N_7323);
or U8384 (N_8384,N_5997,N_6755);
and U8385 (N_8385,N_6413,N_6326);
xor U8386 (N_8386,N_5423,N_5721);
nand U8387 (N_8387,N_7042,N_6094);
and U8388 (N_8388,N_5662,N_6659);
and U8389 (N_8389,N_6311,N_7396);
nand U8390 (N_8390,N_7385,N_5717);
nor U8391 (N_8391,N_5753,N_7276);
xnor U8392 (N_8392,N_6183,N_5735);
nand U8393 (N_8393,N_6612,N_5978);
xor U8394 (N_8394,N_5589,N_7419);
xor U8395 (N_8395,N_6350,N_7198);
xor U8396 (N_8396,N_6478,N_7284);
and U8397 (N_8397,N_7458,N_5505);
or U8398 (N_8398,N_6697,N_6340);
nor U8399 (N_8399,N_6080,N_7237);
or U8400 (N_8400,N_6167,N_5347);
nor U8401 (N_8401,N_5625,N_5511);
nand U8402 (N_8402,N_6155,N_5817);
and U8403 (N_8403,N_5783,N_5940);
or U8404 (N_8404,N_6283,N_7351);
nand U8405 (N_8405,N_7219,N_5702);
or U8406 (N_8406,N_5025,N_6825);
nand U8407 (N_8407,N_7411,N_5608);
nor U8408 (N_8408,N_7353,N_7381);
nor U8409 (N_8409,N_5517,N_5729);
nor U8410 (N_8410,N_7375,N_7347);
nor U8411 (N_8411,N_5568,N_5332);
and U8412 (N_8412,N_6488,N_7189);
or U8413 (N_8413,N_5341,N_5427);
xnor U8414 (N_8414,N_5353,N_5788);
nand U8415 (N_8415,N_7428,N_6714);
nand U8416 (N_8416,N_6773,N_6915);
and U8417 (N_8417,N_7408,N_7296);
xor U8418 (N_8418,N_6695,N_6921);
or U8419 (N_8419,N_5441,N_5926);
and U8420 (N_8420,N_5974,N_5569);
and U8421 (N_8421,N_7137,N_7232);
nor U8422 (N_8422,N_5224,N_7272);
nor U8423 (N_8423,N_5576,N_6114);
nand U8424 (N_8424,N_6260,N_5210);
or U8425 (N_8425,N_7332,N_6143);
nand U8426 (N_8426,N_6583,N_5138);
nand U8427 (N_8427,N_7349,N_5326);
or U8428 (N_8428,N_5051,N_6627);
nor U8429 (N_8429,N_5246,N_5047);
and U8430 (N_8430,N_7041,N_6483);
nor U8431 (N_8431,N_6215,N_6819);
nor U8432 (N_8432,N_5143,N_6039);
or U8433 (N_8433,N_5535,N_7489);
xor U8434 (N_8434,N_6145,N_6689);
xnor U8435 (N_8435,N_6204,N_6866);
xnor U8436 (N_8436,N_5563,N_5611);
and U8437 (N_8437,N_5209,N_5197);
nand U8438 (N_8438,N_5206,N_5351);
xor U8439 (N_8439,N_5208,N_5650);
xor U8440 (N_8440,N_6782,N_7191);
xnor U8441 (N_8441,N_6457,N_5769);
or U8442 (N_8442,N_7316,N_5480);
nor U8443 (N_8443,N_5915,N_6207);
nor U8444 (N_8444,N_5622,N_7131);
and U8445 (N_8445,N_6916,N_5586);
xnor U8446 (N_8446,N_6797,N_5448);
nand U8447 (N_8447,N_6467,N_7083);
nand U8448 (N_8448,N_6346,N_6752);
and U8449 (N_8449,N_5346,N_6336);
and U8450 (N_8450,N_5137,N_7030);
nor U8451 (N_8451,N_6165,N_7310);
nand U8452 (N_8452,N_5084,N_5055);
xor U8453 (N_8453,N_6999,N_7280);
nor U8454 (N_8454,N_5864,N_6230);
and U8455 (N_8455,N_5530,N_7281);
nand U8456 (N_8456,N_6437,N_7081);
xnor U8457 (N_8457,N_5336,N_5389);
or U8458 (N_8458,N_5759,N_6129);
or U8459 (N_8459,N_6055,N_7231);
or U8460 (N_8460,N_5636,N_6342);
nand U8461 (N_8461,N_5635,N_6231);
nor U8462 (N_8462,N_5184,N_5839);
xor U8463 (N_8463,N_6538,N_7422);
or U8464 (N_8464,N_6312,N_6771);
and U8465 (N_8465,N_6487,N_6486);
or U8466 (N_8466,N_5297,N_5528);
or U8467 (N_8467,N_5383,N_5737);
nand U8468 (N_8468,N_6956,N_5031);
nand U8469 (N_8469,N_6704,N_5097);
nand U8470 (N_8470,N_6573,N_6918);
xor U8471 (N_8471,N_6903,N_6382);
or U8472 (N_8472,N_5492,N_6813);
and U8473 (N_8473,N_7417,N_5462);
nor U8474 (N_8474,N_6784,N_7432);
nor U8475 (N_8475,N_6338,N_6179);
xor U8476 (N_8476,N_5750,N_7491);
nand U8477 (N_8477,N_5169,N_5429);
nor U8478 (N_8478,N_6098,N_6685);
and U8479 (N_8479,N_6205,N_5738);
and U8480 (N_8480,N_5747,N_5787);
and U8481 (N_8481,N_5317,N_6940);
nand U8482 (N_8482,N_7094,N_5550);
or U8483 (N_8483,N_6291,N_7326);
nand U8484 (N_8484,N_5697,N_6556);
nor U8485 (N_8485,N_6545,N_5352);
nand U8486 (N_8486,N_5863,N_5694);
or U8487 (N_8487,N_5678,N_5948);
or U8488 (N_8488,N_7469,N_7363);
and U8489 (N_8489,N_7472,N_6555);
and U8490 (N_8490,N_7459,N_6249);
nor U8491 (N_8491,N_6019,N_5289);
nand U8492 (N_8492,N_6997,N_7012);
and U8493 (N_8493,N_5454,N_6020);
nand U8494 (N_8494,N_5667,N_6436);
or U8495 (N_8495,N_7271,N_5001);
or U8496 (N_8496,N_6299,N_5943);
or U8497 (N_8497,N_6671,N_6126);
nand U8498 (N_8498,N_6765,N_7004);
xnor U8499 (N_8499,N_7178,N_5975);
nand U8500 (N_8500,N_6584,N_5117);
nand U8501 (N_8501,N_5080,N_7480);
nand U8502 (N_8502,N_5373,N_6904);
and U8503 (N_8503,N_6547,N_7328);
nand U8504 (N_8504,N_7060,N_6325);
xnor U8505 (N_8505,N_5411,N_5885);
and U8506 (N_8506,N_7436,N_7153);
nor U8507 (N_8507,N_6511,N_7454);
and U8508 (N_8508,N_7420,N_6450);
nand U8509 (N_8509,N_7008,N_7187);
nor U8510 (N_8510,N_6955,N_5935);
nand U8511 (N_8511,N_5239,N_7020);
xnor U8512 (N_8512,N_6855,N_5232);
or U8513 (N_8513,N_7111,N_5056);
nand U8514 (N_8514,N_7496,N_6066);
xnor U8515 (N_8515,N_7321,N_7490);
and U8516 (N_8516,N_7123,N_5958);
xnor U8517 (N_8517,N_5366,N_6816);
xor U8518 (N_8518,N_6474,N_5061);
nor U8519 (N_8519,N_6416,N_7221);
or U8520 (N_8520,N_6268,N_6220);
and U8521 (N_8521,N_6909,N_7448);
and U8522 (N_8522,N_5116,N_6829);
nor U8523 (N_8523,N_6560,N_5736);
xor U8524 (N_8524,N_6976,N_7450);
nor U8525 (N_8525,N_5966,N_5742);
or U8526 (N_8526,N_6036,N_5956);
and U8527 (N_8527,N_6774,N_6589);
and U8528 (N_8528,N_5994,N_5066);
nand U8529 (N_8529,N_7167,N_6801);
nor U8530 (N_8530,N_6056,N_5096);
nor U8531 (N_8531,N_6298,N_5248);
and U8532 (N_8532,N_5282,N_6553);
nand U8533 (N_8533,N_6140,N_5912);
and U8534 (N_8534,N_6389,N_6864);
nor U8535 (N_8535,N_5399,N_5202);
or U8536 (N_8536,N_6920,N_5790);
and U8537 (N_8537,N_6604,N_5192);
xnor U8538 (N_8538,N_6924,N_5570);
nor U8539 (N_8539,N_5630,N_6189);
and U8540 (N_8540,N_7338,N_6045);
nand U8541 (N_8541,N_6048,N_7423);
or U8542 (N_8542,N_6292,N_6403);
nor U8543 (N_8543,N_6640,N_7289);
and U8544 (N_8544,N_5415,N_5281);
nor U8545 (N_8545,N_5930,N_6674);
and U8546 (N_8546,N_7378,N_5058);
nor U8547 (N_8547,N_6163,N_5823);
xor U8548 (N_8548,N_6054,N_6317);
or U8549 (N_8549,N_6554,N_6351);
nand U8550 (N_8550,N_5591,N_6655);
xor U8551 (N_8551,N_7256,N_6532);
and U8552 (N_8552,N_7226,N_5831);
or U8553 (N_8553,N_7430,N_7383);
and U8554 (N_8554,N_6438,N_5417);
nor U8555 (N_8555,N_6243,N_6360);
nand U8556 (N_8556,N_6493,N_6083);
nand U8557 (N_8557,N_7099,N_6662);
nand U8558 (N_8558,N_6894,N_6369);
and U8559 (N_8559,N_6729,N_6222);
xnor U8560 (N_8560,N_6852,N_6969);
nand U8561 (N_8561,N_5609,N_6104);
or U8562 (N_8562,N_6900,N_5294);
nor U8563 (N_8563,N_7116,N_7203);
or U8564 (N_8564,N_5109,N_7315);
and U8565 (N_8565,N_5477,N_6499);
and U8566 (N_8566,N_5714,N_7387);
nand U8567 (N_8567,N_6971,N_5370);
xnor U8568 (N_8568,N_6664,N_5620);
nand U8569 (N_8569,N_6597,N_6848);
and U8570 (N_8570,N_7236,N_5949);
or U8571 (N_8571,N_6521,N_5654);
nor U8572 (N_8572,N_6718,N_5335);
nor U8573 (N_8573,N_5039,N_5768);
xor U8574 (N_8574,N_6868,N_7263);
nand U8575 (N_8575,N_7341,N_7024);
and U8576 (N_8576,N_6024,N_6681);
and U8577 (N_8577,N_6242,N_6375);
xnor U8578 (N_8578,N_6854,N_5891);
xnor U8579 (N_8579,N_5685,N_7006);
or U8580 (N_8580,N_5009,N_6070);
nor U8581 (N_8581,N_5954,N_7379);
nand U8582 (N_8582,N_6663,N_5618);
nand U8583 (N_8583,N_5981,N_7122);
nor U8584 (N_8584,N_6127,N_5111);
nand U8585 (N_8585,N_6745,N_6559);
nor U8586 (N_8586,N_6121,N_5155);
or U8587 (N_8587,N_5693,N_5325);
nand U8588 (N_8588,N_7120,N_5465);
nand U8589 (N_8589,N_6175,N_6038);
and U8590 (N_8590,N_5054,N_7374);
and U8591 (N_8591,N_7429,N_6025);
nor U8592 (N_8592,N_6693,N_6223);
or U8593 (N_8593,N_5760,N_5587);
xor U8594 (N_8594,N_5709,N_5652);
and U8595 (N_8595,N_6386,N_5941);
nand U8596 (N_8596,N_5129,N_7093);
or U8597 (N_8597,N_7065,N_7343);
and U8598 (N_8598,N_5727,N_6430);
and U8599 (N_8599,N_6418,N_6858);
nor U8600 (N_8600,N_7434,N_5249);
xnor U8601 (N_8601,N_5464,N_5139);
xnor U8602 (N_8602,N_7446,N_5582);
nand U8603 (N_8603,N_5933,N_6285);
xnor U8604 (N_8604,N_5253,N_6034);
xor U8605 (N_8605,N_6832,N_6246);
or U8606 (N_8606,N_5313,N_6715);
or U8607 (N_8607,N_6974,N_7129);
and U8608 (N_8608,N_6740,N_6925);
xor U8609 (N_8609,N_7134,N_7444);
nand U8610 (N_8610,N_7209,N_5203);
nand U8611 (N_8611,N_6339,N_5743);
nand U8612 (N_8612,N_6694,N_6680);
and U8613 (N_8613,N_5637,N_6717);
xor U8614 (N_8614,N_5425,N_6551);
nand U8615 (N_8615,N_5467,N_5870);
xor U8616 (N_8616,N_5395,N_6047);
and U8617 (N_8617,N_7369,N_6090);
or U8618 (N_8618,N_5043,N_6629);
and U8619 (N_8619,N_6628,N_5955);
nand U8620 (N_8620,N_5998,N_6494);
nor U8621 (N_8621,N_5792,N_5907);
or U8622 (N_8622,N_6368,N_6134);
nand U8623 (N_8623,N_5682,N_6523);
nor U8624 (N_8624,N_5160,N_7025);
nand U8625 (N_8625,N_6050,N_5375);
nor U8626 (N_8626,N_5663,N_5917);
nand U8627 (N_8627,N_6192,N_6550);
and U8628 (N_8628,N_6216,N_6561);
xor U8629 (N_8629,N_7485,N_6320);
nand U8630 (N_8630,N_6686,N_5306);
and U8631 (N_8631,N_7119,N_5828);
nand U8632 (N_8632,N_5804,N_6936);
and U8633 (N_8633,N_5358,N_6119);
nand U8634 (N_8634,N_5331,N_5119);
and U8635 (N_8635,N_5450,N_5852);
xor U8636 (N_8636,N_6624,N_6889);
and U8637 (N_8637,N_5469,N_6951);
or U8638 (N_8638,N_6328,N_5895);
or U8639 (N_8639,N_6953,N_5396);
nor U8640 (N_8640,N_5068,N_7101);
nor U8641 (N_8641,N_5144,N_7269);
or U8642 (N_8642,N_7032,N_6160);
xnor U8643 (N_8643,N_5120,N_5502);
or U8644 (N_8644,N_5268,N_5655);
xor U8645 (N_8645,N_6939,N_5920);
or U8646 (N_8646,N_5243,N_6148);
and U8647 (N_8647,N_5646,N_5962);
or U8648 (N_8648,N_5278,N_7268);
xnor U8649 (N_8649,N_5763,N_7086);
nor U8650 (N_8650,N_5220,N_5564);
nand U8651 (N_8651,N_7350,N_5301);
xor U8652 (N_8652,N_5670,N_6180);
or U8653 (N_8653,N_6296,N_5712);
nand U8654 (N_8654,N_5244,N_6780);
and U8655 (N_8655,N_5514,N_6790);
xor U8656 (N_8656,N_6822,N_7213);
nand U8657 (N_8657,N_5830,N_7176);
nor U8658 (N_8658,N_6324,N_5273);
or U8659 (N_8659,N_5420,N_7358);
nor U8660 (N_8660,N_5234,N_6427);
or U8661 (N_8661,N_6334,N_5174);
and U8662 (N_8662,N_7405,N_5805);
xnor U8663 (N_8663,N_5778,N_6206);
xnor U8664 (N_8664,N_7318,N_6912);
xor U8665 (N_8665,N_5200,N_7308);
and U8666 (N_8666,N_5421,N_5928);
or U8667 (N_8667,N_5164,N_6091);
nand U8668 (N_8668,N_6947,N_6877);
and U8669 (N_8669,N_7287,N_7277);
nand U8670 (N_8670,N_5913,N_5242);
xor U8671 (N_8671,N_6111,N_6289);
nor U8672 (N_8672,N_6990,N_5233);
nand U8673 (N_8673,N_5229,N_6509);
xnor U8674 (N_8674,N_6667,N_5671);
and U8675 (N_8675,N_7118,N_7147);
or U8676 (N_8676,N_5585,N_6238);
or U8677 (N_8677,N_6259,N_5304);
nand U8678 (N_8678,N_5896,N_5886);
and U8679 (N_8679,N_6027,N_5644);
xnor U8680 (N_8680,N_7028,N_5677);
and U8681 (N_8681,N_6256,N_7140);
or U8682 (N_8682,N_5022,N_7362);
or U8683 (N_8683,N_5131,N_6975);
and U8684 (N_8684,N_5776,N_6880);
nand U8685 (N_8685,N_6232,N_7286);
and U8686 (N_8686,N_6505,N_6980);
and U8687 (N_8687,N_6359,N_5658);
and U8688 (N_8688,N_6802,N_6716);
or U8689 (N_8689,N_6846,N_6052);
xnor U8690 (N_8690,N_6895,N_7291);
xor U8691 (N_8691,N_6710,N_6870);
or U8692 (N_8692,N_6273,N_5456);
or U8693 (N_8693,N_6614,N_6015);
xor U8694 (N_8694,N_6503,N_6528);
nand U8695 (N_8695,N_5461,N_6081);
nor U8696 (N_8696,N_6144,N_6341);
nor U8697 (N_8697,N_7114,N_6073);
nand U8698 (N_8698,N_7261,N_7467);
xor U8699 (N_8699,N_6891,N_6835);
and U8700 (N_8700,N_7425,N_7461);
nand U8701 (N_8701,N_5199,N_7249);
nand U8702 (N_8702,N_6060,N_7252);
nor U8703 (N_8703,N_6279,N_6172);
and U8704 (N_8704,N_7306,N_7388);
and U8705 (N_8705,N_5698,N_5666);
nor U8706 (N_8706,N_5466,N_7473);
xnor U8707 (N_8707,N_5984,N_6028);
xor U8708 (N_8708,N_5217,N_6199);
and U8709 (N_8709,N_6906,N_6534);
and U8710 (N_8710,N_6968,N_5900);
xor U8711 (N_8711,N_6602,N_5471);
nand U8712 (N_8712,N_6120,N_6461);
nand U8713 (N_8713,N_6586,N_6516);
nor U8714 (N_8714,N_6213,N_5967);
xnor U8715 (N_8715,N_7474,N_5093);
nand U8716 (N_8716,N_5152,N_5632);
or U8717 (N_8717,N_5687,N_7001);
and U8718 (N_8718,N_6448,N_6424);
and U8719 (N_8719,N_5226,N_7267);
nor U8720 (N_8720,N_7312,N_5337);
nor U8721 (N_8721,N_5865,N_6548);
or U8722 (N_8722,N_7303,N_5240);
nand U8723 (N_8723,N_6611,N_5810);
or U8724 (N_8724,N_6863,N_5381);
or U8725 (N_8725,N_7274,N_6658);
nand U8726 (N_8726,N_6684,N_6271);
xnor U8727 (N_8727,N_7367,N_5604);
nand U8728 (N_8728,N_7257,N_5868);
nand U8729 (N_8729,N_5360,N_6086);
and U8730 (N_8730,N_5108,N_5746);
nor U8731 (N_8731,N_6623,N_5153);
and U8732 (N_8732,N_5057,N_6301);
xor U8733 (N_8733,N_6530,N_6415);
and U8734 (N_8734,N_5382,N_7313);
nor U8735 (N_8735,N_6653,N_6319);
nor U8736 (N_8736,N_5236,N_5003);
or U8737 (N_8737,N_6708,N_5494);
nand U8738 (N_8738,N_6071,N_5333);
nand U8739 (N_8739,N_7082,N_5245);
and U8740 (N_8740,N_6151,N_6251);
nand U8741 (N_8741,N_6973,N_6562);
nor U8742 (N_8742,N_5937,N_5023);
or U8743 (N_8743,N_6421,N_5901);
or U8744 (N_8744,N_7302,N_5508);
nor U8745 (N_8745,N_6096,N_5359);
and U8746 (N_8746,N_6820,N_5647);
xnor U8747 (N_8747,N_5818,N_6188);
nor U8748 (N_8748,N_5893,N_6113);
nor U8749 (N_8749,N_5315,N_5812);
nor U8750 (N_8750,N_5632,N_5284);
nand U8751 (N_8751,N_5383,N_5758);
or U8752 (N_8752,N_6377,N_5707);
nand U8753 (N_8753,N_7198,N_5443);
xor U8754 (N_8754,N_5280,N_6690);
nor U8755 (N_8755,N_5043,N_6070);
xor U8756 (N_8756,N_5943,N_7249);
and U8757 (N_8757,N_5195,N_5558);
and U8758 (N_8758,N_5902,N_5378);
xnor U8759 (N_8759,N_6581,N_7179);
or U8760 (N_8760,N_6919,N_6116);
xor U8761 (N_8761,N_6358,N_7188);
nor U8762 (N_8762,N_6850,N_5269);
or U8763 (N_8763,N_6047,N_7458);
nand U8764 (N_8764,N_6072,N_5449);
xor U8765 (N_8765,N_7042,N_7374);
xnor U8766 (N_8766,N_5031,N_5338);
or U8767 (N_8767,N_6219,N_6102);
and U8768 (N_8768,N_6893,N_5047);
or U8769 (N_8769,N_5964,N_5890);
or U8770 (N_8770,N_6959,N_6047);
and U8771 (N_8771,N_6069,N_6419);
nand U8772 (N_8772,N_6500,N_6251);
and U8773 (N_8773,N_5074,N_6669);
xor U8774 (N_8774,N_5511,N_5386);
or U8775 (N_8775,N_6569,N_7340);
and U8776 (N_8776,N_6911,N_5778);
xnor U8777 (N_8777,N_7113,N_5339);
and U8778 (N_8778,N_5297,N_6030);
or U8779 (N_8779,N_5631,N_6022);
and U8780 (N_8780,N_7399,N_7201);
and U8781 (N_8781,N_5523,N_7002);
nand U8782 (N_8782,N_5840,N_5714);
and U8783 (N_8783,N_7130,N_5683);
and U8784 (N_8784,N_6040,N_6780);
nand U8785 (N_8785,N_5669,N_5375);
xor U8786 (N_8786,N_5693,N_6551);
nor U8787 (N_8787,N_7325,N_5820);
and U8788 (N_8788,N_6009,N_7214);
nand U8789 (N_8789,N_5158,N_6750);
xor U8790 (N_8790,N_5356,N_6152);
nor U8791 (N_8791,N_5296,N_6716);
nor U8792 (N_8792,N_6564,N_7106);
nor U8793 (N_8793,N_7282,N_5376);
xor U8794 (N_8794,N_7075,N_5755);
nand U8795 (N_8795,N_6281,N_6493);
nand U8796 (N_8796,N_5884,N_7471);
or U8797 (N_8797,N_5491,N_7365);
xnor U8798 (N_8798,N_6458,N_7071);
nand U8799 (N_8799,N_5309,N_5385);
or U8800 (N_8800,N_7005,N_5168);
or U8801 (N_8801,N_5164,N_6495);
and U8802 (N_8802,N_6948,N_6660);
xor U8803 (N_8803,N_5084,N_6697);
xor U8804 (N_8804,N_6269,N_5324);
or U8805 (N_8805,N_5633,N_5822);
and U8806 (N_8806,N_6749,N_5945);
nand U8807 (N_8807,N_6156,N_6339);
xnor U8808 (N_8808,N_6534,N_6703);
xor U8809 (N_8809,N_6113,N_6230);
xnor U8810 (N_8810,N_6114,N_7412);
nand U8811 (N_8811,N_5225,N_6200);
or U8812 (N_8812,N_6505,N_7219);
nor U8813 (N_8813,N_6987,N_5805);
xor U8814 (N_8814,N_7422,N_6862);
nor U8815 (N_8815,N_5202,N_5456);
nand U8816 (N_8816,N_6743,N_5538);
xor U8817 (N_8817,N_5463,N_6811);
nand U8818 (N_8818,N_5629,N_5239);
and U8819 (N_8819,N_7234,N_6659);
and U8820 (N_8820,N_5146,N_5574);
xnor U8821 (N_8821,N_6705,N_5156);
and U8822 (N_8822,N_6394,N_5570);
nor U8823 (N_8823,N_7250,N_6715);
nor U8824 (N_8824,N_5527,N_5217);
nand U8825 (N_8825,N_7027,N_5004);
and U8826 (N_8826,N_5657,N_7205);
nand U8827 (N_8827,N_6484,N_6845);
nand U8828 (N_8828,N_5777,N_5873);
xor U8829 (N_8829,N_6735,N_6573);
nand U8830 (N_8830,N_5594,N_5868);
nor U8831 (N_8831,N_5169,N_6068);
nand U8832 (N_8832,N_5427,N_7358);
or U8833 (N_8833,N_6398,N_5113);
or U8834 (N_8834,N_6080,N_7259);
xor U8835 (N_8835,N_5712,N_5433);
or U8836 (N_8836,N_7196,N_6122);
and U8837 (N_8837,N_5691,N_5510);
xor U8838 (N_8838,N_5814,N_6452);
nor U8839 (N_8839,N_5693,N_7083);
nand U8840 (N_8840,N_7477,N_5015);
or U8841 (N_8841,N_6763,N_7439);
nor U8842 (N_8842,N_5163,N_5009);
nand U8843 (N_8843,N_7221,N_6437);
and U8844 (N_8844,N_6722,N_5658);
nor U8845 (N_8845,N_5110,N_5063);
xor U8846 (N_8846,N_6806,N_5641);
nor U8847 (N_8847,N_5744,N_6909);
nor U8848 (N_8848,N_6480,N_7064);
xnor U8849 (N_8849,N_6578,N_7439);
nand U8850 (N_8850,N_5208,N_6054);
or U8851 (N_8851,N_5542,N_7174);
or U8852 (N_8852,N_7492,N_5213);
xor U8853 (N_8853,N_7046,N_7107);
nand U8854 (N_8854,N_6970,N_7302);
or U8855 (N_8855,N_5088,N_5510);
or U8856 (N_8856,N_7106,N_6964);
nor U8857 (N_8857,N_5411,N_7424);
or U8858 (N_8858,N_7405,N_7212);
nor U8859 (N_8859,N_6562,N_7359);
xnor U8860 (N_8860,N_7305,N_7277);
nor U8861 (N_8861,N_5090,N_5134);
or U8862 (N_8862,N_5082,N_5761);
xor U8863 (N_8863,N_6333,N_5333);
and U8864 (N_8864,N_5310,N_5035);
nand U8865 (N_8865,N_6976,N_5919);
or U8866 (N_8866,N_5716,N_6060);
and U8867 (N_8867,N_6891,N_7149);
and U8868 (N_8868,N_5904,N_5188);
and U8869 (N_8869,N_5348,N_5938);
nor U8870 (N_8870,N_6201,N_6324);
xnor U8871 (N_8871,N_6804,N_7065);
xnor U8872 (N_8872,N_5029,N_5081);
or U8873 (N_8873,N_5846,N_6909);
and U8874 (N_8874,N_5736,N_6473);
and U8875 (N_8875,N_7362,N_6840);
and U8876 (N_8876,N_5354,N_6972);
or U8877 (N_8877,N_7138,N_5919);
and U8878 (N_8878,N_6983,N_6158);
nand U8879 (N_8879,N_5114,N_5602);
and U8880 (N_8880,N_6939,N_6151);
or U8881 (N_8881,N_5096,N_6692);
nor U8882 (N_8882,N_5431,N_5346);
nand U8883 (N_8883,N_5801,N_5770);
nor U8884 (N_8884,N_5723,N_5796);
and U8885 (N_8885,N_6320,N_5246);
xnor U8886 (N_8886,N_6517,N_6044);
xnor U8887 (N_8887,N_5802,N_7079);
nor U8888 (N_8888,N_5482,N_7499);
nor U8889 (N_8889,N_7045,N_7176);
or U8890 (N_8890,N_5486,N_5077);
nand U8891 (N_8891,N_7195,N_5078);
nand U8892 (N_8892,N_5607,N_5228);
or U8893 (N_8893,N_6003,N_6493);
xnor U8894 (N_8894,N_5680,N_5877);
xnor U8895 (N_8895,N_6270,N_5929);
nand U8896 (N_8896,N_6225,N_6342);
nand U8897 (N_8897,N_5246,N_5065);
nor U8898 (N_8898,N_7198,N_6678);
xor U8899 (N_8899,N_5990,N_6120);
or U8900 (N_8900,N_5553,N_6857);
xor U8901 (N_8901,N_6991,N_7146);
or U8902 (N_8902,N_7483,N_5181);
and U8903 (N_8903,N_7145,N_6194);
nor U8904 (N_8904,N_7107,N_6341);
xnor U8905 (N_8905,N_6063,N_5532);
nand U8906 (N_8906,N_5052,N_5993);
or U8907 (N_8907,N_5993,N_6629);
xor U8908 (N_8908,N_5790,N_6588);
nor U8909 (N_8909,N_5799,N_5855);
or U8910 (N_8910,N_5935,N_5252);
or U8911 (N_8911,N_5541,N_5676);
nand U8912 (N_8912,N_6548,N_7067);
xor U8913 (N_8913,N_6841,N_5424);
xor U8914 (N_8914,N_5980,N_6679);
nand U8915 (N_8915,N_6984,N_5139);
and U8916 (N_8916,N_5005,N_6626);
nor U8917 (N_8917,N_5305,N_5665);
and U8918 (N_8918,N_5554,N_5070);
and U8919 (N_8919,N_5627,N_5589);
and U8920 (N_8920,N_6760,N_6031);
or U8921 (N_8921,N_6666,N_6618);
nand U8922 (N_8922,N_6744,N_6678);
or U8923 (N_8923,N_6670,N_6612);
or U8924 (N_8924,N_7359,N_6285);
xnor U8925 (N_8925,N_7015,N_6040);
nand U8926 (N_8926,N_5522,N_5806);
nand U8927 (N_8927,N_7475,N_6788);
or U8928 (N_8928,N_5965,N_6834);
xor U8929 (N_8929,N_6884,N_6100);
nand U8930 (N_8930,N_5533,N_5479);
nor U8931 (N_8931,N_7063,N_7007);
nor U8932 (N_8932,N_5869,N_6661);
xor U8933 (N_8933,N_6627,N_5948);
nand U8934 (N_8934,N_5054,N_5298);
nor U8935 (N_8935,N_5160,N_5917);
and U8936 (N_8936,N_6760,N_5920);
nor U8937 (N_8937,N_5080,N_6223);
xnor U8938 (N_8938,N_6522,N_5064);
or U8939 (N_8939,N_7213,N_6976);
or U8940 (N_8940,N_7153,N_6815);
or U8941 (N_8941,N_6352,N_5529);
nand U8942 (N_8942,N_5565,N_6673);
and U8943 (N_8943,N_6922,N_6592);
xnor U8944 (N_8944,N_6278,N_6601);
or U8945 (N_8945,N_5328,N_5931);
nand U8946 (N_8946,N_6762,N_5321);
and U8947 (N_8947,N_6756,N_7161);
xnor U8948 (N_8948,N_6341,N_6434);
nand U8949 (N_8949,N_6021,N_5455);
and U8950 (N_8950,N_6893,N_7310);
and U8951 (N_8951,N_6511,N_7286);
and U8952 (N_8952,N_6010,N_6406);
and U8953 (N_8953,N_5572,N_6761);
nor U8954 (N_8954,N_5229,N_7443);
nand U8955 (N_8955,N_5747,N_6676);
nor U8956 (N_8956,N_5183,N_6791);
or U8957 (N_8957,N_5147,N_5943);
xor U8958 (N_8958,N_6501,N_6913);
and U8959 (N_8959,N_5273,N_6585);
nand U8960 (N_8960,N_7138,N_5684);
nand U8961 (N_8961,N_5949,N_6458);
or U8962 (N_8962,N_5916,N_6385);
nor U8963 (N_8963,N_5704,N_7384);
nand U8964 (N_8964,N_6519,N_6798);
xnor U8965 (N_8965,N_5713,N_5110);
or U8966 (N_8966,N_6854,N_6695);
nand U8967 (N_8967,N_5726,N_6490);
nor U8968 (N_8968,N_6200,N_6747);
nand U8969 (N_8969,N_6750,N_6567);
or U8970 (N_8970,N_6811,N_5737);
or U8971 (N_8971,N_6218,N_5157);
nor U8972 (N_8972,N_5524,N_6695);
nand U8973 (N_8973,N_7198,N_5801);
xor U8974 (N_8974,N_6157,N_6090);
and U8975 (N_8975,N_7330,N_6800);
nand U8976 (N_8976,N_5254,N_6821);
or U8977 (N_8977,N_5007,N_6731);
nand U8978 (N_8978,N_5125,N_7459);
or U8979 (N_8979,N_5514,N_6775);
nor U8980 (N_8980,N_5878,N_6895);
nand U8981 (N_8981,N_6721,N_7119);
nor U8982 (N_8982,N_7240,N_6352);
nor U8983 (N_8983,N_6994,N_5280);
nand U8984 (N_8984,N_6093,N_6799);
and U8985 (N_8985,N_6119,N_7385);
xor U8986 (N_8986,N_6274,N_6114);
nand U8987 (N_8987,N_5868,N_6716);
and U8988 (N_8988,N_6221,N_6924);
nor U8989 (N_8989,N_7219,N_6322);
nor U8990 (N_8990,N_6686,N_7319);
or U8991 (N_8991,N_7044,N_6900);
and U8992 (N_8992,N_5394,N_7267);
xor U8993 (N_8993,N_6414,N_7426);
or U8994 (N_8994,N_5421,N_7331);
and U8995 (N_8995,N_6120,N_5369);
nand U8996 (N_8996,N_6780,N_6157);
or U8997 (N_8997,N_5237,N_6535);
or U8998 (N_8998,N_7419,N_6757);
or U8999 (N_8999,N_6228,N_6412);
or U9000 (N_9000,N_6069,N_6941);
xor U9001 (N_9001,N_5455,N_6630);
nand U9002 (N_9002,N_6582,N_6503);
nor U9003 (N_9003,N_6358,N_7218);
nand U9004 (N_9004,N_5239,N_5566);
xnor U9005 (N_9005,N_6578,N_7158);
and U9006 (N_9006,N_7065,N_5935);
or U9007 (N_9007,N_6065,N_5795);
xor U9008 (N_9008,N_6717,N_6193);
or U9009 (N_9009,N_6365,N_6229);
and U9010 (N_9010,N_7107,N_6026);
and U9011 (N_9011,N_6667,N_6682);
nor U9012 (N_9012,N_7215,N_7391);
xnor U9013 (N_9013,N_5883,N_6293);
or U9014 (N_9014,N_7313,N_6178);
xor U9015 (N_9015,N_6981,N_6688);
and U9016 (N_9016,N_6868,N_5816);
or U9017 (N_9017,N_7358,N_5184);
or U9018 (N_9018,N_5705,N_5793);
or U9019 (N_9019,N_5801,N_6223);
xor U9020 (N_9020,N_7327,N_6257);
or U9021 (N_9021,N_6494,N_7291);
xnor U9022 (N_9022,N_5003,N_5361);
and U9023 (N_9023,N_7348,N_6475);
and U9024 (N_9024,N_5352,N_7341);
nor U9025 (N_9025,N_5657,N_7374);
nor U9026 (N_9026,N_6208,N_5694);
nand U9027 (N_9027,N_5622,N_5044);
xor U9028 (N_9028,N_7123,N_5483);
and U9029 (N_9029,N_6297,N_6441);
and U9030 (N_9030,N_6269,N_5464);
xor U9031 (N_9031,N_6140,N_6426);
and U9032 (N_9032,N_5865,N_5736);
nand U9033 (N_9033,N_5851,N_7203);
nand U9034 (N_9034,N_5268,N_5581);
nor U9035 (N_9035,N_7011,N_6407);
nor U9036 (N_9036,N_7089,N_5180);
and U9037 (N_9037,N_6732,N_7394);
or U9038 (N_9038,N_6556,N_6807);
xor U9039 (N_9039,N_6152,N_6537);
nand U9040 (N_9040,N_5662,N_6596);
or U9041 (N_9041,N_5706,N_7355);
or U9042 (N_9042,N_5876,N_6479);
and U9043 (N_9043,N_7325,N_5512);
or U9044 (N_9044,N_5077,N_5039);
nand U9045 (N_9045,N_6940,N_7296);
xnor U9046 (N_9046,N_6401,N_5080);
and U9047 (N_9047,N_5206,N_7034);
nand U9048 (N_9048,N_7131,N_5647);
nand U9049 (N_9049,N_7380,N_5152);
nand U9050 (N_9050,N_6115,N_6920);
nand U9051 (N_9051,N_5818,N_7469);
or U9052 (N_9052,N_5506,N_6953);
nand U9053 (N_9053,N_6980,N_5381);
nand U9054 (N_9054,N_5825,N_5841);
and U9055 (N_9055,N_6805,N_7374);
nand U9056 (N_9056,N_6997,N_5145);
and U9057 (N_9057,N_7158,N_6113);
or U9058 (N_9058,N_6651,N_5976);
nand U9059 (N_9059,N_5249,N_6288);
nor U9060 (N_9060,N_5693,N_7098);
nor U9061 (N_9061,N_6303,N_6013);
nand U9062 (N_9062,N_6793,N_7329);
or U9063 (N_9063,N_7007,N_7133);
or U9064 (N_9064,N_6686,N_6838);
nand U9065 (N_9065,N_5815,N_6355);
and U9066 (N_9066,N_5588,N_5114);
nand U9067 (N_9067,N_5612,N_6398);
and U9068 (N_9068,N_7131,N_5233);
and U9069 (N_9069,N_5214,N_7319);
nand U9070 (N_9070,N_5443,N_5922);
xnor U9071 (N_9071,N_6761,N_5142);
or U9072 (N_9072,N_7291,N_7486);
nor U9073 (N_9073,N_6321,N_5405);
or U9074 (N_9074,N_6611,N_5590);
nor U9075 (N_9075,N_7390,N_6959);
nand U9076 (N_9076,N_7155,N_5898);
xor U9077 (N_9077,N_5471,N_6928);
or U9078 (N_9078,N_7480,N_5165);
nand U9079 (N_9079,N_5774,N_7035);
xor U9080 (N_9080,N_6679,N_7281);
nor U9081 (N_9081,N_5489,N_5420);
or U9082 (N_9082,N_6468,N_7417);
or U9083 (N_9083,N_6676,N_6866);
or U9084 (N_9084,N_6042,N_5544);
and U9085 (N_9085,N_7329,N_6641);
nand U9086 (N_9086,N_5319,N_5295);
nand U9087 (N_9087,N_6959,N_6253);
and U9088 (N_9088,N_7409,N_7074);
or U9089 (N_9089,N_5671,N_5868);
xnor U9090 (N_9090,N_7229,N_6808);
nor U9091 (N_9091,N_5196,N_7291);
xor U9092 (N_9092,N_7049,N_6135);
and U9093 (N_9093,N_7491,N_6627);
xor U9094 (N_9094,N_7493,N_6302);
nand U9095 (N_9095,N_5833,N_6438);
nor U9096 (N_9096,N_5224,N_7089);
nor U9097 (N_9097,N_7029,N_5164);
nand U9098 (N_9098,N_6837,N_7288);
nand U9099 (N_9099,N_6073,N_6204);
and U9100 (N_9100,N_5302,N_6043);
nand U9101 (N_9101,N_6488,N_5432);
nand U9102 (N_9102,N_7328,N_6252);
xnor U9103 (N_9103,N_5495,N_7254);
and U9104 (N_9104,N_5962,N_5410);
or U9105 (N_9105,N_5906,N_7468);
nand U9106 (N_9106,N_5944,N_5619);
or U9107 (N_9107,N_5003,N_5970);
nor U9108 (N_9108,N_5091,N_6669);
xnor U9109 (N_9109,N_5651,N_5607);
xor U9110 (N_9110,N_6502,N_5927);
nor U9111 (N_9111,N_6037,N_6198);
and U9112 (N_9112,N_5945,N_5001);
xor U9113 (N_9113,N_5561,N_7091);
or U9114 (N_9114,N_5778,N_6954);
nand U9115 (N_9115,N_5617,N_6904);
or U9116 (N_9116,N_6322,N_7279);
nor U9117 (N_9117,N_5949,N_7471);
xnor U9118 (N_9118,N_5839,N_7397);
or U9119 (N_9119,N_7419,N_5540);
nor U9120 (N_9120,N_7154,N_5266);
xnor U9121 (N_9121,N_7065,N_6734);
and U9122 (N_9122,N_5225,N_7227);
nand U9123 (N_9123,N_7133,N_7413);
and U9124 (N_9124,N_7180,N_5437);
nor U9125 (N_9125,N_7488,N_7207);
nor U9126 (N_9126,N_7430,N_5569);
or U9127 (N_9127,N_6764,N_5854);
nor U9128 (N_9128,N_5724,N_5287);
xnor U9129 (N_9129,N_5324,N_7427);
nor U9130 (N_9130,N_5307,N_6949);
or U9131 (N_9131,N_6400,N_5806);
or U9132 (N_9132,N_5049,N_5011);
xnor U9133 (N_9133,N_5962,N_6494);
nand U9134 (N_9134,N_5612,N_5602);
nand U9135 (N_9135,N_6908,N_6289);
xor U9136 (N_9136,N_6885,N_6234);
nor U9137 (N_9137,N_7362,N_6441);
or U9138 (N_9138,N_5197,N_7131);
or U9139 (N_9139,N_6123,N_5603);
and U9140 (N_9140,N_6998,N_6048);
xor U9141 (N_9141,N_5179,N_7240);
or U9142 (N_9142,N_6207,N_6153);
nor U9143 (N_9143,N_6425,N_6989);
xor U9144 (N_9144,N_5804,N_6053);
nor U9145 (N_9145,N_6680,N_7175);
or U9146 (N_9146,N_6883,N_5904);
or U9147 (N_9147,N_6780,N_7120);
xnor U9148 (N_9148,N_7278,N_5531);
nor U9149 (N_9149,N_5562,N_5420);
xor U9150 (N_9150,N_6098,N_7377);
and U9151 (N_9151,N_6960,N_5701);
and U9152 (N_9152,N_7406,N_6343);
xor U9153 (N_9153,N_7076,N_7071);
and U9154 (N_9154,N_6318,N_5406);
nand U9155 (N_9155,N_5910,N_5950);
or U9156 (N_9156,N_5872,N_6072);
xnor U9157 (N_9157,N_5289,N_6304);
or U9158 (N_9158,N_5285,N_6920);
and U9159 (N_9159,N_7169,N_7105);
or U9160 (N_9160,N_5517,N_5750);
nor U9161 (N_9161,N_6195,N_6635);
or U9162 (N_9162,N_6851,N_5391);
and U9163 (N_9163,N_6101,N_7324);
nor U9164 (N_9164,N_5167,N_6747);
nor U9165 (N_9165,N_6580,N_5770);
nor U9166 (N_9166,N_6666,N_5403);
nand U9167 (N_9167,N_7388,N_6391);
xnor U9168 (N_9168,N_6178,N_5377);
xnor U9169 (N_9169,N_7317,N_6480);
xor U9170 (N_9170,N_6790,N_5851);
xor U9171 (N_9171,N_6671,N_5782);
or U9172 (N_9172,N_6913,N_6713);
nand U9173 (N_9173,N_5254,N_7261);
xnor U9174 (N_9174,N_6666,N_6005);
nand U9175 (N_9175,N_7360,N_7134);
nand U9176 (N_9176,N_7083,N_6879);
xnor U9177 (N_9177,N_6055,N_5412);
and U9178 (N_9178,N_6143,N_6977);
or U9179 (N_9179,N_5858,N_7016);
xnor U9180 (N_9180,N_5233,N_7165);
and U9181 (N_9181,N_6515,N_5067);
nor U9182 (N_9182,N_6478,N_5464);
and U9183 (N_9183,N_6404,N_7080);
or U9184 (N_9184,N_6607,N_7060);
xnor U9185 (N_9185,N_5694,N_7306);
nor U9186 (N_9186,N_7051,N_6047);
and U9187 (N_9187,N_7191,N_5974);
and U9188 (N_9188,N_7334,N_5727);
or U9189 (N_9189,N_7110,N_7109);
or U9190 (N_9190,N_6956,N_7443);
nor U9191 (N_9191,N_6609,N_5254);
nand U9192 (N_9192,N_5079,N_5884);
and U9193 (N_9193,N_5119,N_5358);
and U9194 (N_9194,N_5223,N_6902);
or U9195 (N_9195,N_6243,N_6266);
xor U9196 (N_9196,N_7498,N_5163);
nand U9197 (N_9197,N_5850,N_6228);
nor U9198 (N_9198,N_6356,N_7499);
nand U9199 (N_9199,N_5096,N_5422);
xnor U9200 (N_9200,N_6658,N_7323);
nand U9201 (N_9201,N_5496,N_5745);
nand U9202 (N_9202,N_6350,N_7241);
nand U9203 (N_9203,N_6768,N_6754);
and U9204 (N_9204,N_5917,N_6905);
and U9205 (N_9205,N_7432,N_5612);
nor U9206 (N_9206,N_7105,N_6226);
xor U9207 (N_9207,N_7371,N_5447);
nand U9208 (N_9208,N_6274,N_5261);
nor U9209 (N_9209,N_6171,N_7228);
xnor U9210 (N_9210,N_5809,N_5122);
and U9211 (N_9211,N_5310,N_7174);
xor U9212 (N_9212,N_6387,N_5087);
xor U9213 (N_9213,N_7061,N_7189);
nand U9214 (N_9214,N_5019,N_5729);
xnor U9215 (N_9215,N_6341,N_5006);
xnor U9216 (N_9216,N_6060,N_6398);
xor U9217 (N_9217,N_7105,N_6919);
nand U9218 (N_9218,N_5955,N_7031);
xnor U9219 (N_9219,N_5453,N_6777);
nand U9220 (N_9220,N_7442,N_5669);
nand U9221 (N_9221,N_6182,N_6424);
nor U9222 (N_9222,N_5985,N_6351);
or U9223 (N_9223,N_7350,N_6505);
and U9224 (N_9224,N_7055,N_7370);
nor U9225 (N_9225,N_7047,N_7283);
and U9226 (N_9226,N_5484,N_7395);
xor U9227 (N_9227,N_5258,N_5292);
and U9228 (N_9228,N_7035,N_6874);
and U9229 (N_9229,N_5072,N_5251);
nor U9230 (N_9230,N_7219,N_5503);
or U9231 (N_9231,N_6163,N_5403);
nor U9232 (N_9232,N_6243,N_5443);
and U9233 (N_9233,N_5707,N_5974);
nand U9234 (N_9234,N_5793,N_7053);
nor U9235 (N_9235,N_5871,N_5663);
nand U9236 (N_9236,N_5090,N_5625);
nand U9237 (N_9237,N_6680,N_5343);
nor U9238 (N_9238,N_6841,N_7070);
nor U9239 (N_9239,N_6194,N_6590);
xnor U9240 (N_9240,N_5272,N_6709);
nand U9241 (N_9241,N_5580,N_7135);
or U9242 (N_9242,N_6978,N_5463);
or U9243 (N_9243,N_6014,N_6391);
or U9244 (N_9244,N_6713,N_5007);
xor U9245 (N_9245,N_6523,N_5152);
xor U9246 (N_9246,N_5168,N_5964);
nor U9247 (N_9247,N_5254,N_5197);
and U9248 (N_9248,N_6842,N_5112);
nand U9249 (N_9249,N_5332,N_6868);
and U9250 (N_9250,N_5093,N_6441);
or U9251 (N_9251,N_6658,N_6049);
or U9252 (N_9252,N_6897,N_6490);
xnor U9253 (N_9253,N_6277,N_6159);
nand U9254 (N_9254,N_7183,N_7019);
and U9255 (N_9255,N_5476,N_5977);
or U9256 (N_9256,N_7098,N_7435);
and U9257 (N_9257,N_6515,N_5084);
or U9258 (N_9258,N_6801,N_5614);
nor U9259 (N_9259,N_6683,N_7308);
and U9260 (N_9260,N_6731,N_5574);
xnor U9261 (N_9261,N_6288,N_5424);
nand U9262 (N_9262,N_7409,N_5429);
and U9263 (N_9263,N_5819,N_5854);
nand U9264 (N_9264,N_7230,N_5039);
and U9265 (N_9265,N_7047,N_5154);
nor U9266 (N_9266,N_6788,N_6161);
nor U9267 (N_9267,N_6849,N_5647);
nand U9268 (N_9268,N_7143,N_5280);
xor U9269 (N_9269,N_5802,N_6409);
and U9270 (N_9270,N_7437,N_7024);
or U9271 (N_9271,N_5154,N_7101);
nand U9272 (N_9272,N_5117,N_5152);
and U9273 (N_9273,N_6294,N_6358);
and U9274 (N_9274,N_6900,N_6697);
and U9275 (N_9275,N_7147,N_7144);
nor U9276 (N_9276,N_6615,N_6613);
or U9277 (N_9277,N_5414,N_6164);
nand U9278 (N_9278,N_5743,N_7103);
xor U9279 (N_9279,N_5468,N_5806);
and U9280 (N_9280,N_5937,N_7339);
or U9281 (N_9281,N_5508,N_6887);
and U9282 (N_9282,N_5990,N_7455);
nor U9283 (N_9283,N_7331,N_6901);
nand U9284 (N_9284,N_5524,N_5027);
xor U9285 (N_9285,N_5303,N_6920);
or U9286 (N_9286,N_5914,N_6161);
and U9287 (N_9287,N_5343,N_6008);
nand U9288 (N_9288,N_6016,N_6577);
nor U9289 (N_9289,N_6458,N_7103);
nand U9290 (N_9290,N_6192,N_6858);
xnor U9291 (N_9291,N_6467,N_5485);
nor U9292 (N_9292,N_6275,N_5526);
or U9293 (N_9293,N_6648,N_6362);
xnor U9294 (N_9294,N_5399,N_6648);
nand U9295 (N_9295,N_6175,N_6217);
and U9296 (N_9296,N_5168,N_6963);
nor U9297 (N_9297,N_6767,N_5469);
nor U9298 (N_9298,N_7012,N_6393);
nor U9299 (N_9299,N_5266,N_5489);
nand U9300 (N_9300,N_6720,N_6088);
xor U9301 (N_9301,N_7046,N_6150);
nand U9302 (N_9302,N_6603,N_6740);
nor U9303 (N_9303,N_6498,N_5757);
xor U9304 (N_9304,N_5229,N_7285);
nand U9305 (N_9305,N_6480,N_5612);
xor U9306 (N_9306,N_5319,N_5159);
nand U9307 (N_9307,N_6296,N_5589);
xor U9308 (N_9308,N_6305,N_7493);
xor U9309 (N_9309,N_5495,N_5007);
or U9310 (N_9310,N_6099,N_7049);
or U9311 (N_9311,N_5832,N_6472);
nor U9312 (N_9312,N_5017,N_7495);
nand U9313 (N_9313,N_6104,N_7326);
nor U9314 (N_9314,N_7266,N_6574);
nand U9315 (N_9315,N_5822,N_7361);
nand U9316 (N_9316,N_6999,N_6091);
nor U9317 (N_9317,N_5523,N_6643);
nor U9318 (N_9318,N_5488,N_6262);
nor U9319 (N_9319,N_7134,N_5896);
nand U9320 (N_9320,N_7127,N_6522);
nor U9321 (N_9321,N_6283,N_7250);
nand U9322 (N_9322,N_6462,N_7413);
nand U9323 (N_9323,N_5948,N_5699);
xnor U9324 (N_9324,N_7341,N_7496);
xor U9325 (N_9325,N_6732,N_5442);
nand U9326 (N_9326,N_5512,N_7192);
xor U9327 (N_9327,N_6283,N_6876);
or U9328 (N_9328,N_5278,N_7081);
xor U9329 (N_9329,N_6426,N_5727);
nor U9330 (N_9330,N_6669,N_7075);
and U9331 (N_9331,N_5336,N_7017);
nand U9332 (N_9332,N_5486,N_6643);
nor U9333 (N_9333,N_6774,N_5264);
and U9334 (N_9334,N_6169,N_6946);
xnor U9335 (N_9335,N_5333,N_6936);
and U9336 (N_9336,N_6435,N_5968);
nor U9337 (N_9337,N_7061,N_6449);
or U9338 (N_9338,N_6049,N_7407);
nand U9339 (N_9339,N_6092,N_6395);
nor U9340 (N_9340,N_7064,N_6001);
or U9341 (N_9341,N_6958,N_5496);
nor U9342 (N_9342,N_6863,N_5125);
xnor U9343 (N_9343,N_5487,N_6764);
and U9344 (N_9344,N_5461,N_5287);
nand U9345 (N_9345,N_5378,N_7130);
or U9346 (N_9346,N_7102,N_5151);
or U9347 (N_9347,N_5883,N_6257);
or U9348 (N_9348,N_6763,N_5986);
and U9349 (N_9349,N_6208,N_5583);
nor U9350 (N_9350,N_5215,N_7353);
or U9351 (N_9351,N_6526,N_7074);
xnor U9352 (N_9352,N_5759,N_6862);
and U9353 (N_9353,N_6051,N_6810);
or U9354 (N_9354,N_6904,N_6202);
nand U9355 (N_9355,N_6230,N_5915);
or U9356 (N_9356,N_6722,N_6319);
xnor U9357 (N_9357,N_6296,N_5241);
nor U9358 (N_9358,N_7015,N_5629);
and U9359 (N_9359,N_5575,N_6969);
nor U9360 (N_9360,N_6394,N_7446);
and U9361 (N_9361,N_7320,N_6311);
xor U9362 (N_9362,N_7253,N_6777);
and U9363 (N_9363,N_6058,N_7414);
nand U9364 (N_9364,N_5911,N_5746);
or U9365 (N_9365,N_6009,N_5409);
nor U9366 (N_9366,N_5916,N_5040);
or U9367 (N_9367,N_6976,N_6161);
and U9368 (N_9368,N_6670,N_6201);
or U9369 (N_9369,N_7127,N_7280);
nor U9370 (N_9370,N_5808,N_6255);
and U9371 (N_9371,N_6276,N_6450);
or U9372 (N_9372,N_7201,N_5611);
xor U9373 (N_9373,N_6258,N_7116);
nand U9374 (N_9374,N_5163,N_5895);
nand U9375 (N_9375,N_6855,N_5588);
or U9376 (N_9376,N_5083,N_5895);
and U9377 (N_9377,N_5171,N_7033);
and U9378 (N_9378,N_5782,N_6703);
nand U9379 (N_9379,N_5202,N_6809);
or U9380 (N_9380,N_5353,N_6162);
xnor U9381 (N_9381,N_5352,N_7138);
and U9382 (N_9382,N_5214,N_6372);
nand U9383 (N_9383,N_5280,N_5463);
and U9384 (N_9384,N_6977,N_5393);
nand U9385 (N_9385,N_6438,N_6893);
and U9386 (N_9386,N_7126,N_7364);
nor U9387 (N_9387,N_6388,N_5884);
nor U9388 (N_9388,N_6197,N_6450);
nand U9389 (N_9389,N_5018,N_6139);
or U9390 (N_9390,N_6088,N_5908);
or U9391 (N_9391,N_6466,N_7010);
nand U9392 (N_9392,N_6943,N_6748);
nand U9393 (N_9393,N_6040,N_5972);
and U9394 (N_9394,N_7014,N_7266);
nand U9395 (N_9395,N_6242,N_7310);
or U9396 (N_9396,N_7383,N_7241);
and U9397 (N_9397,N_6266,N_5107);
and U9398 (N_9398,N_7346,N_6721);
or U9399 (N_9399,N_6455,N_5248);
and U9400 (N_9400,N_5221,N_5746);
xor U9401 (N_9401,N_5145,N_6507);
and U9402 (N_9402,N_6653,N_6092);
and U9403 (N_9403,N_5651,N_6687);
or U9404 (N_9404,N_5980,N_5627);
nand U9405 (N_9405,N_5394,N_5992);
nand U9406 (N_9406,N_6767,N_6308);
xor U9407 (N_9407,N_5770,N_6935);
xor U9408 (N_9408,N_5513,N_7482);
nand U9409 (N_9409,N_6877,N_6741);
and U9410 (N_9410,N_5457,N_6977);
xor U9411 (N_9411,N_5512,N_7039);
and U9412 (N_9412,N_6842,N_7387);
or U9413 (N_9413,N_6886,N_5210);
or U9414 (N_9414,N_6790,N_5628);
or U9415 (N_9415,N_7298,N_6033);
xnor U9416 (N_9416,N_5839,N_6919);
xor U9417 (N_9417,N_6718,N_6124);
xnor U9418 (N_9418,N_7069,N_5923);
and U9419 (N_9419,N_5939,N_6352);
nor U9420 (N_9420,N_6872,N_7125);
xnor U9421 (N_9421,N_5243,N_6263);
nor U9422 (N_9422,N_5247,N_6790);
and U9423 (N_9423,N_6030,N_7471);
or U9424 (N_9424,N_6002,N_5344);
and U9425 (N_9425,N_7271,N_6552);
nor U9426 (N_9426,N_7283,N_5492);
xor U9427 (N_9427,N_5313,N_6229);
nor U9428 (N_9428,N_5110,N_6626);
nor U9429 (N_9429,N_6573,N_5997);
nand U9430 (N_9430,N_6053,N_5713);
nor U9431 (N_9431,N_5209,N_7405);
nor U9432 (N_9432,N_7322,N_5611);
and U9433 (N_9433,N_6036,N_6143);
nand U9434 (N_9434,N_7408,N_5243);
and U9435 (N_9435,N_6383,N_5269);
nor U9436 (N_9436,N_7235,N_6291);
and U9437 (N_9437,N_5526,N_5817);
nor U9438 (N_9438,N_7375,N_5734);
nand U9439 (N_9439,N_6868,N_5688);
nand U9440 (N_9440,N_5433,N_5528);
xor U9441 (N_9441,N_5406,N_5380);
nor U9442 (N_9442,N_6774,N_5235);
or U9443 (N_9443,N_7213,N_5269);
or U9444 (N_9444,N_6072,N_6113);
xnor U9445 (N_9445,N_5475,N_5991);
and U9446 (N_9446,N_6804,N_5474);
nor U9447 (N_9447,N_6156,N_6250);
nand U9448 (N_9448,N_6393,N_6140);
nand U9449 (N_9449,N_5073,N_6334);
xnor U9450 (N_9450,N_5720,N_7321);
xnor U9451 (N_9451,N_6711,N_7338);
and U9452 (N_9452,N_7000,N_6253);
nor U9453 (N_9453,N_6023,N_5238);
xor U9454 (N_9454,N_5001,N_5776);
nand U9455 (N_9455,N_6903,N_6767);
nor U9456 (N_9456,N_6122,N_6936);
nor U9457 (N_9457,N_6939,N_6161);
nor U9458 (N_9458,N_7397,N_6671);
and U9459 (N_9459,N_7119,N_5049);
xor U9460 (N_9460,N_5461,N_6763);
or U9461 (N_9461,N_6849,N_6386);
nand U9462 (N_9462,N_6797,N_5892);
and U9463 (N_9463,N_7437,N_6979);
nor U9464 (N_9464,N_6296,N_7017);
xor U9465 (N_9465,N_7272,N_5343);
nor U9466 (N_9466,N_6254,N_5565);
nor U9467 (N_9467,N_6311,N_5122);
nand U9468 (N_9468,N_6439,N_7133);
and U9469 (N_9469,N_5378,N_5249);
nand U9470 (N_9470,N_5774,N_5021);
nor U9471 (N_9471,N_7255,N_5625);
xor U9472 (N_9472,N_7158,N_7357);
and U9473 (N_9473,N_7236,N_5817);
xor U9474 (N_9474,N_7364,N_6311);
nor U9475 (N_9475,N_5091,N_6336);
and U9476 (N_9476,N_5518,N_6777);
nor U9477 (N_9477,N_5384,N_5255);
nor U9478 (N_9478,N_6098,N_6307);
nand U9479 (N_9479,N_5872,N_7097);
nand U9480 (N_9480,N_5944,N_6604);
nor U9481 (N_9481,N_6166,N_5279);
xor U9482 (N_9482,N_7397,N_7381);
nor U9483 (N_9483,N_5390,N_5204);
or U9484 (N_9484,N_7057,N_6583);
xnor U9485 (N_9485,N_7079,N_6737);
nor U9486 (N_9486,N_7434,N_6335);
and U9487 (N_9487,N_7464,N_7268);
nand U9488 (N_9488,N_6684,N_5541);
and U9489 (N_9489,N_7291,N_6176);
nor U9490 (N_9490,N_7487,N_5348);
and U9491 (N_9491,N_6035,N_6545);
and U9492 (N_9492,N_6782,N_5764);
nand U9493 (N_9493,N_6288,N_6368);
xnor U9494 (N_9494,N_7198,N_6968);
xnor U9495 (N_9495,N_5627,N_7128);
nand U9496 (N_9496,N_6518,N_6615);
nor U9497 (N_9497,N_6465,N_6333);
xnor U9498 (N_9498,N_7328,N_6326);
nor U9499 (N_9499,N_6944,N_5673);
or U9500 (N_9500,N_7433,N_7460);
xnor U9501 (N_9501,N_5472,N_5492);
or U9502 (N_9502,N_6754,N_5380);
xor U9503 (N_9503,N_5820,N_5204);
xor U9504 (N_9504,N_7439,N_6121);
nand U9505 (N_9505,N_6070,N_5027);
xor U9506 (N_9506,N_7356,N_6327);
or U9507 (N_9507,N_5332,N_7350);
and U9508 (N_9508,N_6649,N_7229);
and U9509 (N_9509,N_5254,N_7273);
and U9510 (N_9510,N_6793,N_6772);
xnor U9511 (N_9511,N_5101,N_6660);
xor U9512 (N_9512,N_5023,N_5632);
nor U9513 (N_9513,N_7267,N_5605);
nor U9514 (N_9514,N_7008,N_6446);
or U9515 (N_9515,N_6618,N_5564);
and U9516 (N_9516,N_5581,N_5276);
and U9517 (N_9517,N_5256,N_5942);
nand U9518 (N_9518,N_6283,N_5105);
nor U9519 (N_9519,N_6570,N_6520);
or U9520 (N_9520,N_5347,N_6074);
or U9521 (N_9521,N_6673,N_6288);
and U9522 (N_9522,N_6118,N_5197);
nand U9523 (N_9523,N_5601,N_5027);
or U9524 (N_9524,N_6370,N_5970);
nor U9525 (N_9525,N_5023,N_6980);
and U9526 (N_9526,N_6240,N_7410);
and U9527 (N_9527,N_6270,N_5107);
nand U9528 (N_9528,N_5063,N_6585);
and U9529 (N_9529,N_7280,N_6328);
or U9530 (N_9530,N_6085,N_6185);
xor U9531 (N_9531,N_5083,N_6667);
and U9532 (N_9532,N_5334,N_6218);
xor U9533 (N_9533,N_5733,N_6635);
or U9534 (N_9534,N_6273,N_6686);
or U9535 (N_9535,N_6984,N_6411);
or U9536 (N_9536,N_5267,N_7011);
nand U9537 (N_9537,N_7030,N_7190);
and U9538 (N_9538,N_7183,N_7472);
xor U9539 (N_9539,N_5697,N_6332);
nand U9540 (N_9540,N_5467,N_5919);
or U9541 (N_9541,N_6804,N_5057);
nand U9542 (N_9542,N_5197,N_5150);
and U9543 (N_9543,N_5868,N_6547);
nor U9544 (N_9544,N_7219,N_7076);
xnor U9545 (N_9545,N_5867,N_5498);
nor U9546 (N_9546,N_6486,N_5360);
xor U9547 (N_9547,N_5837,N_5177);
nor U9548 (N_9548,N_5254,N_5508);
xnor U9549 (N_9549,N_6952,N_7121);
nor U9550 (N_9550,N_7159,N_5594);
and U9551 (N_9551,N_7032,N_5478);
nand U9552 (N_9552,N_6375,N_6882);
xnor U9553 (N_9553,N_6261,N_5428);
and U9554 (N_9554,N_5342,N_5255);
nand U9555 (N_9555,N_5911,N_5500);
nor U9556 (N_9556,N_5942,N_5811);
xor U9557 (N_9557,N_5983,N_5068);
nor U9558 (N_9558,N_6995,N_7009);
and U9559 (N_9559,N_5369,N_5338);
nand U9560 (N_9560,N_5271,N_6973);
and U9561 (N_9561,N_6490,N_5778);
nand U9562 (N_9562,N_6665,N_6414);
and U9563 (N_9563,N_6222,N_6774);
or U9564 (N_9564,N_6030,N_7246);
or U9565 (N_9565,N_6256,N_5009);
xor U9566 (N_9566,N_5522,N_5375);
xor U9567 (N_9567,N_5715,N_6369);
nand U9568 (N_9568,N_7155,N_6498);
or U9569 (N_9569,N_5950,N_5648);
nand U9570 (N_9570,N_6774,N_6264);
or U9571 (N_9571,N_6397,N_7059);
nor U9572 (N_9572,N_5040,N_7499);
nor U9573 (N_9573,N_6099,N_7374);
or U9574 (N_9574,N_6869,N_5136);
or U9575 (N_9575,N_6944,N_5127);
xor U9576 (N_9576,N_6156,N_6187);
xor U9577 (N_9577,N_5339,N_6964);
nor U9578 (N_9578,N_5598,N_6256);
and U9579 (N_9579,N_7136,N_5465);
xnor U9580 (N_9580,N_5836,N_5760);
and U9581 (N_9581,N_6861,N_5239);
nor U9582 (N_9582,N_6929,N_5584);
nor U9583 (N_9583,N_7086,N_6886);
nor U9584 (N_9584,N_5295,N_7066);
nand U9585 (N_9585,N_6202,N_5666);
or U9586 (N_9586,N_6830,N_5011);
nor U9587 (N_9587,N_7424,N_5192);
nand U9588 (N_9588,N_5379,N_7172);
and U9589 (N_9589,N_6157,N_5103);
or U9590 (N_9590,N_5398,N_5786);
or U9591 (N_9591,N_7392,N_7382);
nand U9592 (N_9592,N_5158,N_6244);
nor U9593 (N_9593,N_6007,N_6440);
xnor U9594 (N_9594,N_6899,N_6462);
xor U9595 (N_9595,N_5779,N_5467);
or U9596 (N_9596,N_7180,N_5510);
xnor U9597 (N_9597,N_6167,N_5549);
or U9598 (N_9598,N_5921,N_6928);
nand U9599 (N_9599,N_6989,N_6482);
nor U9600 (N_9600,N_7323,N_6339);
xnor U9601 (N_9601,N_6034,N_6741);
xor U9602 (N_9602,N_6798,N_6109);
xor U9603 (N_9603,N_6397,N_6174);
nor U9604 (N_9604,N_6655,N_6759);
nor U9605 (N_9605,N_5459,N_6980);
or U9606 (N_9606,N_6600,N_6033);
or U9607 (N_9607,N_6316,N_5663);
nand U9608 (N_9608,N_5331,N_6455);
or U9609 (N_9609,N_6628,N_7016);
nor U9610 (N_9610,N_7208,N_6231);
xor U9611 (N_9611,N_5310,N_6815);
nor U9612 (N_9612,N_5396,N_5649);
nor U9613 (N_9613,N_7089,N_6072);
nand U9614 (N_9614,N_5568,N_6649);
nor U9615 (N_9615,N_6046,N_5387);
nand U9616 (N_9616,N_6989,N_5034);
nand U9617 (N_9617,N_6486,N_5128);
or U9618 (N_9618,N_5184,N_6931);
xnor U9619 (N_9619,N_5369,N_6997);
xor U9620 (N_9620,N_5364,N_6214);
xnor U9621 (N_9621,N_6134,N_5613);
or U9622 (N_9622,N_5667,N_6702);
and U9623 (N_9623,N_6798,N_5355);
xor U9624 (N_9624,N_5068,N_6476);
nor U9625 (N_9625,N_5015,N_6160);
nor U9626 (N_9626,N_6019,N_7145);
or U9627 (N_9627,N_6765,N_7210);
xnor U9628 (N_9628,N_5634,N_5640);
nand U9629 (N_9629,N_5514,N_7435);
xnor U9630 (N_9630,N_6322,N_6757);
and U9631 (N_9631,N_6299,N_7134);
nor U9632 (N_9632,N_5850,N_5078);
and U9633 (N_9633,N_6752,N_5838);
nor U9634 (N_9634,N_5750,N_5823);
and U9635 (N_9635,N_5602,N_7370);
or U9636 (N_9636,N_5292,N_7048);
and U9637 (N_9637,N_5139,N_6890);
nor U9638 (N_9638,N_6110,N_6457);
or U9639 (N_9639,N_6244,N_6624);
nand U9640 (N_9640,N_5335,N_5843);
and U9641 (N_9641,N_5723,N_6042);
or U9642 (N_9642,N_6047,N_5515);
nor U9643 (N_9643,N_7237,N_5994);
or U9644 (N_9644,N_6110,N_5608);
nor U9645 (N_9645,N_6203,N_6219);
xor U9646 (N_9646,N_6578,N_5931);
or U9647 (N_9647,N_5825,N_7031);
nand U9648 (N_9648,N_5153,N_6711);
nand U9649 (N_9649,N_5129,N_6700);
nor U9650 (N_9650,N_5327,N_5777);
nor U9651 (N_9651,N_7216,N_5211);
xnor U9652 (N_9652,N_6266,N_5138);
xor U9653 (N_9653,N_5738,N_5805);
or U9654 (N_9654,N_5078,N_5791);
nor U9655 (N_9655,N_5320,N_7247);
xor U9656 (N_9656,N_6056,N_5684);
xnor U9657 (N_9657,N_7396,N_5325);
nor U9658 (N_9658,N_6595,N_7330);
or U9659 (N_9659,N_5487,N_6039);
nand U9660 (N_9660,N_6296,N_5834);
and U9661 (N_9661,N_5111,N_7190);
nor U9662 (N_9662,N_7301,N_7066);
xor U9663 (N_9663,N_5988,N_6374);
and U9664 (N_9664,N_7348,N_5730);
nand U9665 (N_9665,N_5766,N_5060);
or U9666 (N_9666,N_6914,N_6686);
or U9667 (N_9667,N_6056,N_5600);
xnor U9668 (N_9668,N_6587,N_7432);
nand U9669 (N_9669,N_6876,N_5002);
and U9670 (N_9670,N_7496,N_5619);
xnor U9671 (N_9671,N_7314,N_6696);
nand U9672 (N_9672,N_7089,N_6001);
nand U9673 (N_9673,N_6615,N_5333);
or U9674 (N_9674,N_5691,N_5555);
nand U9675 (N_9675,N_6898,N_6834);
nand U9676 (N_9676,N_5867,N_5987);
and U9677 (N_9677,N_5000,N_5878);
nor U9678 (N_9678,N_7270,N_6340);
and U9679 (N_9679,N_5597,N_7425);
nand U9680 (N_9680,N_6821,N_5063);
nor U9681 (N_9681,N_6813,N_5573);
or U9682 (N_9682,N_7351,N_6750);
and U9683 (N_9683,N_5748,N_5492);
nand U9684 (N_9684,N_7082,N_5007);
nor U9685 (N_9685,N_5099,N_6508);
nand U9686 (N_9686,N_5226,N_6733);
xnor U9687 (N_9687,N_7437,N_6323);
and U9688 (N_9688,N_7175,N_7279);
nor U9689 (N_9689,N_6992,N_7415);
or U9690 (N_9690,N_6797,N_6043);
xnor U9691 (N_9691,N_7129,N_6153);
xnor U9692 (N_9692,N_6608,N_7493);
nand U9693 (N_9693,N_5388,N_5842);
nor U9694 (N_9694,N_5338,N_5061);
and U9695 (N_9695,N_7476,N_7453);
and U9696 (N_9696,N_7095,N_5356);
nand U9697 (N_9697,N_7286,N_6966);
and U9698 (N_9698,N_7077,N_7057);
nor U9699 (N_9699,N_6676,N_5285);
or U9700 (N_9700,N_6434,N_6075);
and U9701 (N_9701,N_5851,N_6528);
xor U9702 (N_9702,N_7418,N_5553);
or U9703 (N_9703,N_5724,N_5641);
nor U9704 (N_9704,N_7137,N_5587);
xor U9705 (N_9705,N_6292,N_5944);
and U9706 (N_9706,N_7149,N_7025);
nand U9707 (N_9707,N_6623,N_7241);
nand U9708 (N_9708,N_6936,N_5080);
or U9709 (N_9709,N_5787,N_6920);
nand U9710 (N_9710,N_6357,N_7026);
or U9711 (N_9711,N_6606,N_6483);
or U9712 (N_9712,N_6903,N_6653);
nor U9713 (N_9713,N_6052,N_5437);
nor U9714 (N_9714,N_7197,N_6740);
xor U9715 (N_9715,N_7217,N_5497);
nor U9716 (N_9716,N_5270,N_7126);
and U9717 (N_9717,N_5168,N_6649);
xor U9718 (N_9718,N_5520,N_6416);
and U9719 (N_9719,N_5912,N_6539);
xnor U9720 (N_9720,N_6714,N_7299);
and U9721 (N_9721,N_6561,N_6438);
nand U9722 (N_9722,N_6279,N_5364);
nor U9723 (N_9723,N_6952,N_5614);
nand U9724 (N_9724,N_6544,N_5343);
xor U9725 (N_9725,N_6731,N_5535);
and U9726 (N_9726,N_7463,N_6884);
and U9727 (N_9727,N_6740,N_6386);
or U9728 (N_9728,N_6905,N_7400);
and U9729 (N_9729,N_7422,N_6180);
nand U9730 (N_9730,N_7153,N_5152);
nand U9731 (N_9731,N_5587,N_5127);
or U9732 (N_9732,N_6519,N_7242);
nor U9733 (N_9733,N_7035,N_5439);
or U9734 (N_9734,N_6273,N_6586);
nor U9735 (N_9735,N_5720,N_6616);
nor U9736 (N_9736,N_7472,N_5574);
and U9737 (N_9737,N_6211,N_5611);
xor U9738 (N_9738,N_7412,N_5103);
nand U9739 (N_9739,N_6943,N_7308);
and U9740 (N_9740,N_5260,N_7412);
xor U9741 (N_9741,N_7130,N_5517);
or U9742 (N_9742,N_5552,N_6313);
and U9743 (N_9743,N_6700,N_5867);
and U9744 (N_9744,N_5483,N_5997);
or U9745 (N_9745,N_6363,N_5822);
and U9746 (N_9746,N_7452,N_6559);
and U9747 (N_9747,N_7461,N_5262);
nand U9748 (N_9748,N_5750,N_6353);
or U9749 (N_9749,N_7454,N_6747);
nor U9750 (N_9750,N_6315,N_6899);
and U9751 (N_9751,N_5965,N_5953);
xor U9752 (N_9752,N_7256,N_6585);
nor U9753 (N_9753,N_6708,N_5966);
nor U9754 (N_9754,N_6141,N_5404);
or U9755 (N_9755,N_6005,N_6275);
nand U9756 (N_9756,N_5967,N_5431);
and U9757 (N_9757,N_6388,N_5343);
nor U9758 (N_9758,N_6076,N_5286);
nor U9759 (N_9759,N_7455,N_6526);
nand U9760 (N_9760,N_7304,N_5972);
nor U9761 (N_9761,N_5881,N_6686);
nand U9762 (N_9762,N_6121,N_6935);
xnor U9763 (N_9763,N_6355,N_5585);
xor U9764 (N_9764,N_6317,N_6896);
nand U9765 (N_9765,N_6455,N_6343);
nor U9766 (N_9766,N_7454,N_5974);
and U9767 (N_9767,N_6537,N_5095);
or U9768 (N_9768,N_5786,N_6933);
nor U9769 (N_9769,N_7190,N_5419);
nand U9770 (N_9770,N_7369,N_5353);
nand U9771 (N_9771,N_6473,N_6558);
and U9772 (N_9772,N_6984,N_7427);
nor U9773 (N_9773,N_7404,N_6770);
and U9774 (N_9774,N_5337,N_5872);
nor U9775 (N_9775,N_5210,N_5571);
xnor U9776 (N_9776,N_5169,N_5946);
nor U9777 (N_9777,N_5374,N_5535);
nor U9778 (N_9778,N_7047,N_6514);
or U9779 (N_9779,N_5458,N_5664);
or U9780 (N_9780,N_6876,N_7276);
or U9781 (N_9781,N_5629,N_6953);
xnor U9782 (N_9782,N_7149,N_5770);
or U9783 (N_9783,N_7418,N_6455);
nor U9784 (N_9784,N_6827,N_6037);
nand U9785 (N_9785,N_5384,N_5799);
nor U9786 (N_9786,N_5688,N_7000);
or U9787 (N_9787,N_6992,N_5487);
nand U9788 (N_9788,N_5557,N_5567);
nor U9789 (N_9789,N_5332,N_5552);
xnor U9790 (N_9790,N_5568,N_6229);
nand U9791 (N_9791,N_5568,N_6044);
nand U9792 (N_9792,N_6918,N_7018);
nor U9793 (N_9793,N_5895,N_6105);
nor U9794 (N_9794,N_5255,N_5851);
xor U9795 (N_9795,N_6562,N_6645);
xor U9796 (N_9796,N_6709,N_5557);
and U9797 (N_9797,N_5632,N_5754);
or U9798 (N_9798,N_5587,N_6768);
and U9799 (N_9799,N_5741,N_7397);
nand U9800 (N_9800,N_7297,N_7441);
nor U9801 (N_9801,N_5639,N_6066);
nand U9802 (N_9802,N_6865,N_6638);
xnor U9803 (N_9803,N_5376,N_5109);
or U9804 (N_9804,N_5650,N_7211);
or U9805 (N_9805,N_5207,N_5789);
or U9806 (N_9806,N_5217,N_5307);
and U9807 (N_9807,N_5228,N_5144);
xor U9808 (N_9808,N_5328,N_7077);
xnor U9809 (N_9809,N_5806,N_5991);
nand U9810 (N_9810,N_6432,N_6241);
xor U9811 (N_9811,N_5085,N_6901);
xor U9812 (N_9812,N_7342,N_6611);
or U9813 (N_9813,N_5384,N_6350);
nor U9814 (N_9814,N_7238,N_6831);
nor U9815 (N_9815,N_6363,N_5104);
xor U9816 (N_9816,N_7155,N_5709);
and U9817 (N_9817,N_7312,N_6367);
nor U9818 (N_9818,N_5723,N_6834);
nand U9819 (N_9819,N_5602,N_5926);
nand U9820 (N_9820,N_6742,N_7147);
nor U9821 (N_9821,N_5158,N_7331);
nand U9822 (N_9822,N_6480,N_6013);
or U9823 (N_9823,N_5432,N_6455);
xor U9824 (N_9824,N_7396,N_5223);
or U9825 (N_9825,N_6338,N_6311);
nand U9826 (N_9826,N_5908,N_6537);
and U9827 (N_9827,N_6002,N_5749);
or U9828 (N_9828,N_7259,N_5164);
or U9829 (N_9829,N_5141,N_7443);
nor U9830 (N_9830,N_5300,N_5295);
xnor U9831 (N_9831,N_7095,N_5594);
and U9832 (N_9832,N_7496,N_5087);
or U9833 (N_9833,N_7123,N_6090);
nor U9834 (N_9834,N_5862,N_5137);
nor U9835 (N_9835,N_7198,N_5113);
nor U9836 (N_9836,N_5664,N_6731);
xor U9837 (N_9837,N_5550,N_6015);
or U9838 (N_9838,N_5134,N_6601);
and U9839 (N_9839,N_6249,N_5154);
and U9840 (N_9840,N_5617,N_6150);
or U9841 (N_9841,N_6337,N_6226);
xor U9842 (N_9842,N_5755,N_5802);
nor U9843 (N_9843,N_5869,N_7186);
nand U9844 (N_9844,N_5346,N_6265);
nor U9845 (N_9845,N_7115,N_5003);
xor U9846 (N_9846,N_6415,N_7081);
xor U9847 (N_9847,N_5873,N_5427);
nand U9848 (N_9848,N_5543,N_5637);
and U9849 (N_9849,N_6323,N_7157);
xnor U9850 (N_9850,N_5696,N_5526);
nor U9851 (N_9851,N_7099,N_6638);
xnor U9852 (N_9852,N_7204,N_6378);
xnor U9853 (N_9853,N_6680,N_5643);
nor U9854 (N_9854,N_7031,N_6939);
or U9855 (N_9855,N_7286,N_6655);
nor U9856 (N_9856,N_7189,N_5724);
and U9857 (N_9857,N_6106,N_5588);
nor U9858 (N_9858,N_5719,N_5732);
or U9859 (N_9859,N_6609,N_7109);
nor U9860 (N_9860,N_6762,N_6189);
nand U9861 (N_9861,N_5098,N_6180);
nand U9862 (N_9862,N_5510,N_6233);
nor U9863 (N_9863,N_7284,N_7010);
nor U9864 (N_9864,N_7186,N_6936);
and U9865 (N_9865,N_7376,N_6176);
and U9866 (N_9866,N_6602,N_6796);
nand U9867 (N_9867,N_5420,N_7467);
or U9868 (N_9868,N_7491,N_7104);
nand U9869 (N_9869,N_5982,N_6617);
nand U9870 (N_9870,N_5835,N_6349);
nor U9871 (N_9871,N_6675,N_5284);
xnor U9872 (N_9872,N_6310,N_6843);
nor U9873 (N_9873,N_6922,N_5435);
xnor U9874 (N_9874,N_5925,N_5498);
nor U9875 (N_9875,N_7247,N_6169);
nor U9876 (N_9876,N_7087,N_7337);
nand U9877 (N_9877,N_6144,N_5348);
and U9878 (N_9878,N_7128,N_6144);
nand U9879 (N_9879,N_5479,N_7208);
and U9880 (N_9880,N_6318,N_5747);
xnor U9881 (N_9881,N_7003,N_7156);
and U9882 (N_9882,N_6203,N_7138);
nand U9883 (N_9883,N_6722,N_5645);
and U9884 (N_9884,N_6326,N_7346);
and U9885 (N_9885,N_6796,N_5793);
or U9886 (N_9886,N_6659,N_5683);
and U9887 (N_9887,N_7227,N_5650);
nor U9888 (N_9888,N_6642,N_6864);
or U9889 (N_9889,N_6272,N_6680);
xnor U9890 (N_9890,N_5508,N_5073);
and U9891 (N_9891,N_5457,N_7346);
nor U9892 (N_9892,N_7414,N_5507);
and U9893 (N_9893,N_5737,N_5870);
and U9894 (N_9894,N_7049,N_5456);
nor U9895 (N_9895,N_5048,N_6725);
and U9896 (N_9896,N_6855,N_6550);
or U9897 (N_9897,N_7473,N_6504);
xor U9898 (N_9898,N_5451,N_7153);
and U9899 (N_9899,N_6580,N_5792);
xnor U9900 (N_9900,N_6680,N_5421);
nor U9901 (N_9901,N_6082,N_6397);
nand U9902 (N_9902,N_7268,N_6239);
nand U9903 (N_9903,N_6898,N_6230);
nor U9904 (N_9904,N_7154,N_6178);
or U9905 (N_9905,N_6153,N_5500);
nand U9906 (N_9906,N_6764,N_7161);
and U9907 (N_9907,N_5508,N_5238);
xnor U9908 (N_9908,N_6234,N_6912);
and U9909 (N_9909,N_6895,N_5180);
xnor U9910 (N_9910,N_5627,N_6100);
and U9911 (N_9911,N_6820,N_6216);
nand U9912 (N_9912,N_6407,N_7253);
nand U9913 (N_9913,N_6681,N_5215);
nor U9914 (N_9914,N_5348,N_7249);
or U9915 (N_9915,N_6795,N_7179);
nor U9916 (N_9916,N_5200,N_5169);
nand U9917 (N_9917,N_5076,N_6309);
nand U9918 (N_9918,N_6500,N_5614);
nor U9919 (N_9919,N_5209,N_5646);
nor U9920 (N_9920,N_6245,N_5430);
xor U9921 (N_9921,N_5226,N_5618);
nand U9922 (N_9922,N_5771,N_5802);
nor U9923 (N_9923,N_5852,N_6173);
or U9924 (N_9924,N_5436,N_5298);
xor U9925 (N_9925,N_6441,N_5521);
and U9926 (N_9926,N_5002,N_6804);
nor U9927 (N_9927,N_5136,N_7293);
xnor U9928 (N_9928,N_6483,N_6970);
nand U9929 (N_9929,N_6814,N_6839);
or U9930 (N_9930,N_6654,N_7001);
or U9931 (N_9931,N_7276,N_5621);
and U9932 (N_9932,N_7243,N_5651);
and U9933 (N_9933,N_6403,N_6634);
nor U9934 (N_9934,N_6557,N_6703);
and U9935 (N_9935,N_5067,N_6928);
and U9936 (N_9936,N_7099,N_6816);
nor U9937 (N_9937,N_5300,N_7174);
xor U9938 (N_9938,N_7183,N_5140);
or U9939 (N_9939,N_6096,N_6026);
nor U9940 (N_9940,N_6157,N_6358);
nor U9941 (N_9941,N_7231,N_5354);
nand U9942 (N_9942,N_6261,N_6014);
nor U9943 (N_9943,N_6408,N_5377);
xnor U9944 (N_9944,N_5485,N_5787);
or U9945 (N_9945,N_6612,N_6282);
xnor U9946 (N_9946,N_7067,N_6424);
xnor U9947 (N_9947,N_5151,N_7238);
and U9948 (N_9948,N_6486,N_5484);
and U9949 (N_9949,N_5776,N_5899);
xor U9950 (N_9950,N_7174,N_5151);
or U9951 (N_9951,N_5942,N_5750);
xnor U9952 (N_9952,N_5285,N_6926);
nand U9953 (N_9953,N_7496,N_5545);
xnor U9954 (N_9954,N_5442,N_5797);
nand U9955 (N_9955,N_6396,N_5418);
and U9956 (N_9956,N_5123,N_6163);
and U9957 (N_9957,N_7135,N_7083);
nor U9958 (N_9958,N_5270,N_6509);
nor U9959 (N_9959,N_7362,N_6409);
nand U9960 (N_9960,N_7036,N_7299);
and U9961 (N_9961,N_6062,N_5497);
nand U9962 (N_9962,N_5057,N_6416);
and U9963 (N_9963,N_5071,N_5672);
or U9964 (N_9964,N_7478,N_5641);
xor U9965 (N_9965,N_5553,N_5373);
or U9966 (N_9966,N_6130,N_5772);
xnor U9967 (N_9967,N_5713,N_6305);
and U9968 (N_9968,N_6025,N_6990);
nand U9969 (N_9969,N_5281,N_7069);
nand U9970 (N_9970,N_6269,N_5939);
or U9971 (N_9971,N_6517,N_5018);
nor U9972 (N_9972,N_6426,N_7228);
nor U9973 (N_9973,N_7193,N_6345);
nor U9974 (N_9974,N_7006,N_6793);
xor U9975 (N_9975,N_6900,N_5790);
xnor U9976 (N_9976,N_7072,N_5514);
xnor U9977 (N_9977,N_6512,N_6223);
or U9978 (N_9978,N_6323,N_5700);
xor U9979 (N_9979,N_6769,N_6674);
nand U9980 (N_9980,N_6398,N_5296);
xor U9981 (N_9981,N_6394,N_5519);
and U9982 (N_9982,N_6586,N_6303);
nor U9983 (N_9983,N_6673,N_5562);
or U9984 (N_9984,N_7222,N_7449);
nor U9985 (N_9985,N_5247,N_5625);
or U9986 (N_9986,N_7153,N_5123);
xnor U9987 (N_9987,N_5881,N_5445);
nor U9988 (N_9988,N_5151,N_5577);
xor U9989 (N_9989,N_5317,N_7077);
xor U9990 (N_9990,N_6411,N_6800);
xor U9991 (N_9991,N_6835,N_6574);
or U9992 (N_9992,N_6833,N_5596);
nor U9993 (N_9993,N_5380,N_7406);
xnor U9994 (N_9994,N_5064,N_5427);
nand U9995 (N_9995,N_5582,N_6506);
or U9996 (N_9996,N_5442,N_7051);
xnor U9997 (N_9997,N_5935,N_5314);
nor U9998 (N_9998,N_6608,N_6038);
and U9999 (N_9999,N_5881,N_7404);
or U10000 (N_10000,N_9130,N_9720);
nor U10001 (N_10001,N_9005,N_9873);
nand U10002 (N_10002,N_8896,N_8025);
and U10003 (N_10003,N_8076,N_8712);
nand U10004 (N_10004,N_8840,N_9132);
or U10005 (N_10005,N_9957,N_9613);
or U10006 (N_10006,N_9315,N_9670);
nand U10007 (N_10007,N_7845,N_9323);
and U10008 (N_10008,N_7865,N_8623);
or U10009 (N_10009,N_9594,N_8189);
nand U10010 (N_10010,N_8647,N_9235);
and U10011 (N_10011,N_9621,N_9673);
xnor U10012 (N_10012,N_9208,N_7938);
xnor U10013 (N_10013,N_9691,N_8724);
and U10014 (N_10014,N_8820,N_8531);
or U10015 (N_10015,N_9635,N_8907);
nand U10016 (N_10016,N_8219,N_8023);
or U10017 (N_10017,N_9164,N_8019);
nand U10018 (N_10018,N_8425,N_9852);
nor U10019 (N_10019,N_7599,N_7579);
xnor U10020 (N_10020,N_8818,N_9129);
or U10021 (N_10021,N_7621,N_8373);
and U10022 (N_10022,N_9772,N_9950);
nand U10023 (N_10023,N_8194,N_8063);
nand U10024 (N_10024,N_9379,N_9253);
nor U10025 (N_10025,N_8708,N_7541);
nand U10026 (N_10026,N_7742,N_7616);
or U10027 (N_10027,N_7716,N_9926);
xor U10028 (N_10028,N_7650,N_9896);
and U10029 (N_10029,N_8749,N_9361);
and U10030 (N_10030,N_9462,N_7870);
xor U10031 (N_10031,N_8031,N_9649);
or U10032 (N_10032,N_9223,N_9427);
and U10033 (N_10033,N_8001,N_7757);
nand U10034 (N_10034,N_9019,N_8123);
xnor U10035 (N_10035,N_9133,N_8944);
xor U10036 (N_10036,N_8847,N_8095);
and U10037 (N_10037,N_9862,N_8470);
xnor U10038 (N_10038,N_9698,N_9537);
nor U10039 (N_10039,N_9603,N_8554);
xor U10040 (N_10040,N_9480,N_9123);
nor U10041 (N_10041,N_9230,N_7908);
and U10042 (N_10042,N_8550,N_9241);
and U10043 (N_10043,N_8282,N_7726);
nand U10044 (N_10044,N_9316,N_9712);
nor U10045 (N_10045,N_9804,N_9461);
and U10046 (N_10046,N_7822,N_8347);
xnor U10047 (N_10047,N_9411,N_8904);
nand U10048 (N_10048,N_9442,N_7888);
nor U10049 (N_10049,N_7792,N_9261);
and U10050 (N_10050,N_8655,N_8590);
and U10051 (N_10051,N_9474,N_7591);
nor U10052 (N_10052,N_8134,N_9710);
xnor U10053 (N_10053,N_8015,N_8371);
and U10054 (N_10054,N_7975,N_9451);
and U10055 (N_10055,N_8374,N_7996);
xnor U10056 (N_10056,N_7572,N_9909);
and U10057 (N_10057,N_7887,N_7948);
nand U10058 (N_10058,N_9066,N_9262);
xnor U10059 (N_10059,N_7871,N_8264);
nor U10060 (N_10060,N_8585,N_9620);
nor U10061 (N_10061,N_9373,N_8254);
or U10062 (N_10062,N_9582,N_8483);
xnor U10063 (N_10063,N_8789,N_7625);
nor U10064 (N_10064,N_9886,N_9408);
nand U10065 (N_10065,N_9291,N_9935);
or U10066 (N_10066,N_9367,N_9246);
nor U10067 (N_10067,N_8223,N_9760);
nor U10068 (N_10068,N_9871,N_9080);
and U10069 (N_10069,N_9335,N_8301);
and U10070 (N_10070,N_7668,N_9521);
or U10071 (N_10071,N_9992,N_7786);
nor U10072 (N_10072,N_7550,N_8563);
xnor U10073 (N_10073,N_9687,N_7793);
xor U10074 (N_10074,N_7943,N_7573);
nand U10075 (N_10075,N_9380,N_8143);
nand U10076 (N_10076,N_9467,N_8115);
xnor U10077 (N_10077,N_9423,N_9045);
or U10078 (N_10078,N_8379,N_9283);
nand U10079 (N_10079,N_7779,N_9440);
and U10080 (N_10080,N_7527,N_8378);
xor U10081 (N_10081,N_8258,N_9509);
xnor U10082 (N_10082,N_8584,N_9538);
or U10083 (N_10083,N_9511,N_8398);
and U10084 (N_10084,N_8049,N_9643);
nand U10085 (N_10085,N_9978,N_8948);
nor U10086 (N_10086,N_7811,N_8888);
nand U10087 (N_10087,N_7724,N_8202);
xnor U10088 (N_10088,N_9683,N_9515);
xor U10089 (N_10089,N_7615,N_7761);
nor U10090 (N_10090,N_9344,N_9659);
and U10091 (N_10091,N_9333,N_9788);
nand U10092 (N_10092,N_8089,N_7817);
xnor U10093 (N_10093,N_8499,N_7578);
or U10094 (N_10094,N_9212,N_9136);
nand U10095 (N_10095,N_7660,N_8558);
or U10096 (N_10096,N_8694,N_9924);
and U10097 (N_10097,N_8916,N_9415);
xnor U10098 (N_10098,N_8341,N_7720);
xor U10099 (N_10099,N_7755,N_9371);
nor U10100 (N_10100,N_9186,N_9662);
xnor U10101 (N_10101,N_9108,N_9434);
xor U10102 (N_10102,N_9897,N_9175);
nand U10103 (N_10103,N_7998,N_9732);
and U10104 (N_10104,N_9723,N_8087);
xor U10105 (N_10105,N_8669,N_8784);
nor U10106 (N_10106,N_9914,N_9287);
and U10107 (N_10107,N_8476,N_8777);
and U10108 (N_10108,N_8292,N_9485);
or U10109 (N_10109,N_8980,N_9225);
xnor U10110 (N_10110,N_9071,N_9457);
nor U10111 (N_10111,N_8057,N_9868);
xnor U10112 (N_10112,N_8327,N_9417);
nor U10113 (N_10113,N_9386,N_9849);
nor U10114 (N_10114,N_8949,N_9044);
xor U10115 (N_10115,N_9587,N_9820);
xnor U10116 (N_10116,N_8257,N_9837);
xor U10117 (N_10117,N_9048,N_8626);
nand U10118 (N_10118,N_9989,N_8385);
xnor U10119 (N_10119,N_7986,N_8757);
nand U10120 (N_10120,N_9233,N_8416);
nor U10121 (N_10121,N_8882,N_9701);
nand U10122 (N_10122,N_8562,N_9403);
or U10123 (N_10123,N_7713,N_8376);
nand U10124 (N_10124,N_9599,N_8879);
xor U10125 (N_10125,N_9448,N_8658);
nor U10126 (N_10126,N_8042,N_7740);
xor U10127 (N_10127,N_8690,N_9634);
nor U10128 (N_10128,N_8083,N_9733);
and U10129 (N_10129,N_8839,N_7896);
xnor U10130 (N_10130,N_9792,N_8981);
nor U10131 (N_10131,N_8932,N_8866);
xor U10132 (N_10132,N_7984,N_9383);
and U10133 (N_10133,N_9960,N_9646);
nor U10134 (N_10134,N_8136,N_7837);
nand U10135 (N_10135,N_9674,N_7892);
nand U10136 (N_10136,N_8737,N_9624);
nor U10137 (N_10137,N_8106,N_8894);
nand U10138 (N_10138,N_7899,N_8364);
nor U10139 (N_10139,N_9699,N_7647);
xor U10140 (N_10140,N_9679,N_8812);
nor U10141 (N_10141,N_8768,N_9381);
nor U10142 (N_10142,N_7514,N_9310);
xnor U10143 (N_10143,N_7708,N_8165);
or U10144 (N_10144,N_8578,N_9811);
xnor U10145 (N_10145,N_8762,N_9042);
or U10146 (N_10146,N_7500,N_8598);
or U10147 (N_10147,N_9540,N_9738);
or U10148 (N_10148,N_8711,N_8174);
nor U10149 (N_10149,N_8300,N_8654);
nor U10150 (N_10150,N_7507,N_8119);
and U10151 (N_10151,N_8148,N_8765);
or U10152 (N_10152,N_8573,N_8832);
and U10153 (N_10153,N_9161,N_9226);
nor U10154 (N_10154,N_8722,N_9706);
nor U10155 (N_10155,N_7747,N_8328);
nand U10156 (N_10156,N_9481,N_8910);
nor U10157 (N_10157,N_9013,N_9671);
nand U10158 (N_10158,N_9753,N_8231);
and U10159 (N_10159,N_7947,N_8748);
or U10160 (N_10160,N_9356,N_7831);
xor U10161 (N_10161,N_9139,N_7727);
and U10162 (N_10162,N_8852,N_8160);
nor U10163 (N_10163,N_7818,N_9334);
or U10164 (N_10164,N_8725,N_7622);
and U10165 (N_10165,N_7506,N_8715);
or U10166 (N_10166,N_9818,N_9776);
nor U10167 (N_10167,N_9784,N_7776);
xnor U10168 (N_10168,N_8054,N_9399);
or U10169 (N_10169,N_9773,N_9484);
and U10170 (N_10170,N_8596,N_8983);
nor U10171 (N_10171,N_8686,N_9990);
or U10172 (N_10172,N_9830,N_9400);
and U10173 (N_10173,N_9708,N_9860);
xor U10174 (N_10174,N_8849,N_8893);
xnor U10175 (N_10175,N_9134,N_8186);
or U10176 (N_10176,N_8291,N_9827);
nand U10177 (N_10177,N_9516,N_9554);
nor U10178 (N_10178,N_8519,N_7981);
nand U10179 (N_10179,N_8955,N_9833);
xnor U10180 (N_10180,N_9496,N_9996);
nor U10181 (N_10181,N_8078,N_8071);
xor U10182 (N_10182,N_9200,N_8897);
or U10183 (N_10183,N_8286,N_9247);
or U10184 (N_10184,N_9024,N_8609);
and U10185 (N_10185,N_9345,N_8595);
nor U10186 (N_10186,N_7575,N_8681);
xor U10187 (N_10187,N_9363,N_8520);
xnor U10188 (N_10188,N_7777,N_9444);
xor U10189 (N_10189,N_8413,N_8269);
nand U10190 (N_10190,N_8296,N_9102);
nor U10191 (N_10191,N_9799,N_9843);
or U10192 (N_10192,N_8318,N_8493);
xor U10193 (N_10193,N_8842,N_9869);
xor U10194 (N_10194,N_9105,N_8682);
or U10195 (N_10195,N_8815,N_9838);
nor U10196 (N_10196,N_8339,N_9154);
xor U10197 (N_10197,N_7582,N_8576);
nand U10198 (N_10198,N_9320,N_9985);
nand U10199 (N_10199,N_9000,N_7681);
nand U10200 (N_10200,N_8249,N_7836);
nand U10201 (N_10201,N_9302,N_9141);
or U10202 (N_10202,N_9464,N_9207);
nand U10203 (N_10203,N_7741,N_8439);
and U10204 (N_10204,N_8334,N_9368);
nor U10205 (N_10205,N_8235,N_9091);
xnor U10206 (N_10206,N_9700,N_8788);
and U10207 (N_10207,N_9801,N_8800);
and U10208 (N_10208,N_8816,N_8614);
nand U10209 (N_10209,N_7930,N_8926);
xor U10210 (N_10210,N_7942,N_8838);
and U10211 (N_10211,N_8758,N_8858);
nand U10212 (N_10212,N_8941,N_9490);
nor U10213 (N_10213,N_9277,N_9202);
nor U10214 (N_10214,N_8353,N_9745);
nor U10215 (N_10215,N_9864,N_8774);
xnor U10216 (N_10216,N_8028,N_7710);
nor U10217 (N_10217,N_7847,N_8271);
and U10218 (N_10218,N_8319,N_7587);
nor U10219 (N_10219,N_9647,N_7661);
nand U10220 (N_10220,N_8630,N_8723);
and U10221 (N_10221,N_9270,N_7510);
nand U10222 (N_10222,N_8173,N_9475);
or U10223 (N_10223,N_9436,N_9942);
nor U10224 (N_10224,N_9471,N_7982);
and U10225 (N_10225,N_7702,N_9210);
or U10226 (N_10226,N_8092,N_8208);
nor U10227 (N_10227,N_8683,N_8463);
nor U10228 (N_10228,N_8418,N_8135);
or U10229 (N_10229,N_8674,N_7788);
nor U10230 (N_10230,N_8782,N_8138);
or U10231 (N_10231,N_7964,N_7979);
xor U10232 (N_10232,N_9961,N_8921);
nand U10233 (N_10233,N_9558,N_8097);
xor U10234 (N_10234,N_9709,N_8407);
or U10235 (N_10235,N_9718,N_9279);
or U10236 (N_10236,N_9198,N_9692);
nand U10237 (N_10237,N_8600,N_8687);
nand U10238 (N_10238,N_8995,N_9583);
nor U10239 (N_10239,N_8133,N_8744);
nand U10240 (N_10240,N_8278,N_9499);
nand U10241 (N_10241,N_9842,N_9131);
and U10242 (N_10242,N_8033,N_8697);
and U10243 (N_10243,N_7540,N_9529);
nor U10244 (N_10244,N_8833,N_8330);
or U10245 (N_10245,N_9329,N_8359);
nor U10246 (N_10246,N_8671,N_8521);
or U10247 (N_10247,N_7537,N_9598);
or U10248 (N_10248,N_9993,N_9374);
or U10249 (N_10249,N_8157,N_8660);
or U10250 (N_10250,N_8113,N_8244);
xor U10251 (N_10251,N_9932,N_7645);
and U10252 (N_10252,N_9677,N_8024);
or U10253 (N_10253,N_9215,N_7770);
or U10254 (N_10254,N_9128,N_9592);
or U10255 (N_10255,N_7869,N_9174);
nor U10256 (N_10256,N_7627,N_9308);
nand U10257 (N_10257,N_8272,N_9685);
or U10258 (N_10258,N_8635,N_9314);
nor U10259 (N_10259,N_7806,N_9568);
nor U10260 (N_10260,N_9309,N_9376);
and U10261 (N_10261,N_7751,N_8781);
xor U10262 (N_10262,N_7680,N_9187);
xnor U10263 (N_10263,N_7985,N_9238);
nand U10264 (N_10264,N_9234,N_7750);
xor U10265 (N_10265,N_8314,N_9812);
nand U10266 (N_10266,N_7674,N_9878);
and U10267 (N_10267,N_8443,N_9196);
nor U10268 (N_10268,N_8766,N_8928);
or U10269 (N_10269,N_7808,N_9877);
nand U10270 (N_10270,N_8954,N_7919);
nand U10271 (N_10271,N_7790,N_8427);
nor U10272 (N_10272,N_9681,N_9626);
nand U10273 (N_10273,N_9845,N_7653);
nor U10274 (N_10274,N_8699,N_7614);
nor U10275 (N_10275,N_8207,N_8153);
or U10276 (N_10276,N_9815,N_9616);
nand U10277 (N_10277,N_8696,N_7608);
xor U10278 (N_10278,N_7688,N_7866);
xor U10279 (N_10279,N_8661,N_7538);
or U10280 (N_10280,N_9081,N_9739);
and U10281 (N_10281,N_8883,N_9636);
nand U10282 (N_10282,N_9204,N_7917);
nor U10283 (N_10283,N_9149,N_7800);
xnor U10284 (N_10284,N_9027,N_7933);
or U10285 (N_10285,N_7875,N_9747);
nand U10286 (N_10286,N_8583,N_8891);
or U10287 (N_10287,N_9967,N_9527);
nand U10288 (N_10288,N_9968,N_8402);
nor U10289 (N_10289,N_8011,N_9562);
nor U10290 (N_10290,N_9572,N_7915);
xor U10291 (N_10291,N_8363,N_8064);
or U10292 (N_10292,N_9781,N_9824);
or U10293 (N_10293,N_8603,N_7576);
or U10294 (N_10294,N_9660,N_9099);
nor U10295 (N_10295,N_8523,N_9460);
and U10296 (N_10296,N_9243,N_9742);
and U10297 (N_10297,N_8246,N_7701);
and U10298 (N_10298,N_8046,N_9790);
nand U10299 (N_10299,N_9891,N_7787);
nand U10300 (N_10300,N_7771,N_8511);
xor U10301 (N_10301,N_9525,N_9982);
or U10302 (N_10302,N_8344,N_9504);
and U10303 (N_10303,N_7585,N_7611);
and U10304 (N_10304,N_8027,N_8982);
and U10305 (N_10305,N_9795,N_7949);
xnor U10306 (N_10306,N_7501,N_9669);
nand U10307 (N_10307,N_8253,N_9519);
or U10308 (N_10308,N_9576,N_8759);
nand U10309 (N_10309,N_9893,N_9724);
xor U10310 (N_10310,N_9533,N_8565);
xnor U10311 (N_10311,N_9666,N_8146);
nand U10312 (N_10312,N_9337,N_8400);
and U10313 (N_10313,N_9392,N_9328);
nor U10314 (N_10314,N_7598,N_9292);
nand U10315 (N_10315,N_9506,N_8646);
or U10316 (N_10316,N_7853,N_8273);
and U10317 (N_10317,N_7816,N_8529);
nand U10318 (N_10318,N_7738,N_9899);
nor U10319 (N_10319,N_8404,N_9514);
or U10320 (N_10320,N_9232,N_9855);
nand U10321 (N_10321,N_8985,N_7935);
and U10322 (N_10322,N_8061,N_7901);
nor U10323 (N_10323,N_8617,N_7843);
xor U10324 (N_10324,N_8640,N_8912);
or U10325 (N_10325,N_8032,N_7665);
and U10326 (N_10326,N_8915,N_9419);
and U10327 (N_10327,N_9737,N_7781);
nor U10328 (N_10328,N_7618,N_7974);
nor U10329 (N_10329,N_9548,N_8787);
and U10330 (N_10330,N_8485,N_8191);
nand U10331 (N_10331,N_8716,N_9874);
nand U10332 (N_10332,N_9642,N_7858);
nor U10333 (N_10333,N_9413,N_9401);
or U10334 (N_10334,N_9872,N_9654);
and U10335 (N_10335,N_7851,N_8216);
nor U10336 (N_10336,N_7562,N_8796);
or U10337 (N_10337,N_7705,N_8266);
xnor U10338 (N_10338,N_9237,N_7512);
nor U10339 (N_10339,N_8739,N_7610);
nand U10340 (N_10340,N_8961,N_7523);
nand U10341 (N_10341,N_8807,N_8120);
or U10342 (N_10342,N_9991,N_8966);
nand U10343 (N_10343,N_8863,N_8856);
xor U10344 (N_10344,N_9766,N_8229);
nand U10345 (N_10345,N_8307,N_8546);
xnor U10346 (N_10346,N_8978,N_9078);
nand U10347 (N_10347,N_8785,N_9127);
nand U10348 (N_10348,N_9306,N_9284);
and U10349 (N_10349,N_9412,N_8468);
nor U10350 (N_10350,N_9491,N_7687);
nand U10351 (N_10351,N_9549,N_9920);
nand U10352 (N_10352,N_8923,N_9623);
nand U10353 (N_10353,N_8874,N_9676);
nand U10354 (N_10354,N_7569,N_8752);
xnor U10355 (N_10355,N_7605,N_9435);
and U10356 (N_10356,N_8622,N_8791);
nor U10357 (N_10357,N_9832,N_8346);
nor U10358 (N_10358,N_9173,N_9577);
nor U10359 (N_10359,N_9638,N_7881);
or U10360 (N_10360,N_7978,N_8110);
nor U10361 (N_10361,N_7544,N_8964);
nor U10362 (N_10362,N_9093,N_9547);
and U10363 (N_10363,N_9523,N_9251);
nor U10364 (N_10364,N_9902,N_9166);
nand U10365 (N_10365,N_9851,N_8551);
xor U10366 (N_10366,N_8730,N_8804);
nor U10367 (N_10367,N_9163,N_8343);
xor U10368 (N_10368,N_8467,N_8889);
or U10369 (N_10369,N_7667,N_7659);
and U10370 (N_10370,N_9492,N_9744);
nor U10371 (N_10371,N_9263,N_9295);
nand U10372 (N_10372,N_8618,N_7743);
or U10373 (N_10373,N_9998,N_9505);
and U10374 (N_10374,N_9398,N_8652);
xor U10375 (N_10375,N_8579,N_7796);
nand U10376 (N_10376,N_8719,N_9183);
nand U10377 (N_10377,N_8776,N_8677);
or U10378 (N_10378,N_9256,N_8703);
nand U10379 (N_10379,N_8536,N_8643);
nor U10380 (N_10380,N_9500,N_7838);
and U10381 (N_10381,N_8688,N_8155);
nor U10382 (N_10382,N_7977,N_7589);
nand U10383 (N_10383,N_7997,N_9217);
and U10384 (N_10384,N_8226,N_8594);
or U10385 (N_10385,N_8158,N_9915);
nor U10386 (N_10386,N_9938,N_9955);
and U10387 (N_10387,N_9227,N_8692);
or U10388 (N_10388,N_9755,N_9126);
and U10389 (N_10389,N_8974,N_7530);
or U10390 (N_10390,N_8518,N_9876);
and U10391 (N_10391,N_9336,N_8577);
and U10392 (N_10392,N_7868,N_9775);
nand U10393 (N_10393,N_9866,N_8827);
nor U10394 (N_10394,N_8215,N_9817);
or U10395 (N_10395,N_7898,N_9770);
xnor U10396 (N_10396,N_8178,N_9531);
and U10397 (N_10397,N_7723,N_7924);
and U10398 (N_10398,N_8114,N_9049);
nor U10399 (N_10399,N_7557,N_8680);
or U10400 (N_10400,N_9552,N_9796);
nand U10401 (N_10401,N_7783,N_8913);
and U10402 (N_10402,N_8919,N_9269);
nand U10403 (N_10403,N_9656,N_9486);
or U10404 (N_10404,N_7539,N_9446);
xor U10405 (N_10405,N_9189,N_9016);
and U10406 (N_10406,N_9972,N_9157);
and U10407 (N_10407,N_7696,N_9918);
nand U10408 (N_10408,N_8636,N_9581);
and U10409 (N_10409,N_7798,N_8422);
nand U10410 (N_10410,N_9047,N_9821);
and U10411 (N_10411,N_8515,N_8805);
nor U10412 (N_10412,N_8294,N_7860);
nand U10413 (N_10413,N_8547,N_9933);
nand U10414 (N_10414,N_8184,N_9258);
and U10415 (N_10415,N_8320,N_8755);
nand U10416 (N_10416,N_9736,N_8369);
xor U10417 (N_10417,N_9648,N_7878);
nor U10418 (N_10418,N_8192,N_9476);
and U10419 (N_10419,N_9199,N_9242);
or U10420 (N_10420,N_8706,N_9503);
and U10421 (N_10421,N_9420,N_7736);
nor U10422 (N_10422,N_7840,N_8731);
or U10423 (N_10423,N_8629,N_9205);
and U10424 (N_10424,N_7918,N_7521);
nor U10425 (N_10425,N_8009,N_8747);
and U10426 (N_10426,N_9567,N_8624);
and U10427 (N_10427,N_8977,N_9593);
or U10428 (N_10428,N_9853,N_8234);
nand U10429 (N_10429,N_9303,N_9304);
or U10430 (N_10430,N_8336,N_9578);
or U10431 (N_10431,N_9342,N_8675);
xor U10432 (N_10432,N_8568,N_8093);
xnor U10433 (N_10433,N_9079,N_8862);
nor U10434 (N_10434,N_8642,N_7684);
nor U10435 (N_10435,N_8446,N_8797);
nor U10436 (N_10436,N_9120,N_9319);
xor U10437 (N_10437,N_8649,N_8567);
or U10438 (N_10438,N_8736,N_8825);
or U10439 (N_10439,N_9370,N_9816);
and U10440 (N_10440,N_8122,N_8965);
xnor U10441 (N_10441,N_9348,N_7556);
nand U10442 (N_10442,N_8245,N_9997);
and U10443 (N_10443,N_9759,N_8099);
nor U10444 (N_10444,N_8612,N_9966);
or U10445 (N_10445,N_7577,N_9167);
and U10446 (N_10446,N_7960,N_8458);
or U10447 (N_10447,N_9741,N_8767);
and U10448 (N_10448,N_9143,N_9887);
or U10449 (N_10449,N_8695,N_8901);
nor U10450 (N_10450,N_9655,N_9443);
xnor U10451 (N_10451,N_9014,N_9777);
nor U10452 (N_10452,N_8062,N_9349);
nor U10453 (N_10453,N_8950,N_8287);
nor U10454 (N_10454,N_7852,N_8355);
nor U10455 (N_10455,N_8222,N_7991);
or U10456 (N_10456,N_8329,N_9501);
nand U10457 (N_10457,N_9919,N_9007);
nand U10458 (N_10458,N_8070,N_9758);
or U10459 (N_10459,N_9596,N_9299);
nor U10460 (N_10460,N_9495,N_9353);
or U10461 (N_10461,N_7749,N_8022);
xnor U10462 (N_10462,N_9271,N_7628);
nor U10463 (N_10463,N_8854,N_9168);
or U10464 (N_10464,N_7756,N_9979);
nor U10465 (N_10465,N_8338,N_8508);
nand U10466 (N_10466,N_9250,N_9439);
and U10467 (N_10467,N_8494,N_7672);
nor U10468 (N_10468,N_9021,N_9273);
nor U10469 (N_10469,N_9209,N_9389);
nand U10470 (N_10470,N_8382,N_8415);
nand U10471 (N_10471,N_8615,N_8081);
nand U10472 (N_10472,N_9793,N_8108);
xnor U10473 (N_10473,N_7597,N_8345);
or U10474 (N_10474,N_7649,N_9715);
xor U10475 (N_10475,N_8710,N_8745);
nand U10476 (N_10476,N_9663,N_8952);
nor U10477 (N_10477,N_8769,N_9289);
nand U10478 (N_10478,N_9095,N_7634);
xnor U10479 (N_10479,N_7731,N_8817);
and U10480 (N_10480,N_7504,N_9953);
xnor U10481 (N_10481,N_9559,N_9761);
xnor U10482 (N_10482,N_9946,N_8721);
nor U10483 (N_10483,N_8048,N_9780);
or U10484 (N_10484,N_8885,N_8666);
nand U10485 (N_10485,N_8572,N_9927);
xnor U10486 (N_10486,N_8899,N_9055);
or U10487 (N_10487,N_7956,N_8943);
xnor U10488 (N_10488,N_8029,N_7910);
and U10489 (N_10489,N_9840,N_7886);
nand U10490 (N_10490,N_9934,N_7821);
nand U10491 (N_10491,N_8491,N_8420);
nor U10492 (N_10492,N_7911,N_9393);
nand U10493 (N_10493,N_7666,N_8405);
and U10494 (N_10494,N_9075,N_8263);
nand U10495 (N_10495,N_9228,N_9863);
nor U10496 (N_10496,N_7546,N_8410);
or U10497 (N_10497,N_8473,N_8689);
xnor U10498 (N_10498,N_9661,N_8530);
xnor U10499 (N_10499,N_8237,N_9825);
xnor U10500 (N_10500,N_7602,N_9008);
or U10501 (N_10501,N_9541,N_7561);
nor U10502 (N_10502,N_9146,N_9274);
and U10503 (N_10503,N_8069,N_7832);
nor U10504 (N_10504,N_8218,N_8305);
or U10505 (N_10505,N_9879,N_7636);
and U10506 (N_10506,N_7580,N_9359);
and U10507 (N_10507,N_9321,N_9881);
or U10508 (N_10508,N_9033,N_9740);
and U10509 (N_10509,N_7584,N_8331);
or U10510 (N_10510,N_8538,N_7564);
and U10511 (N_10511,N_9473,N_8199);
and U10512 (N_10512,N_7891,N_8311);
nand U10513 (N_10513,N_8627,N_9062);
nor U10514 (N_10514,N_7762,N_9026);
nand U10515 (N_10515,N_9429,N_9407);
nand U10516 (N_10516,N_9728,N_7526);
xnor U10517 (N_10517,N_8945,N_8931);
nor U10518 (N_10518,N_7630,N_9936);
and U10519 (N_10519,N_9857,N_8111);
or U10520 (N_10520,N_9557,N_8662);
xnor U10521 (N_10521,N_8786,N_7678);
nor U10522 (N_10522,N_9151,N_8059);
nor U10523 (N_10523,N_8783,N_8734);
and U10524 (N_10524,N_8720,N_9458);
or U10525 (N_10525,N_9022,N_9422);
nand U10526 (N_10526,N_8096,N_9117);
or U10527 (N_10527,N_8668,N_8250);
nor U10528 (N_10528,N_8128,N_8741);
nand U10529 (N_10529,N_8464,N_8599);
and U10530 (N_10530,N_7529,N_9252);
nand U10531 (N_10531,N_8159,N_8243);
nand U10532 (N_10532,N_8566,N_9889);
nand U10533 (N_10533,N_9591,N_8052);
and U10534 (N_10534,N_7675,N_9059);
or U10535 (N_10535,N_8605,N_8993);
and U10536 (N_10536,N_9923,N_8471);
nor U10537 (N_10537,N_7931,N_9888);
or U10538 (N_10538,N_9901,N_8559);
nor U10539 (N_10539,N_9324,N_7690);
xor U10540 (N_10540,N_8238,N_8121);
nand U10541 (N_10541,N_7846,N_8150);
nor U10542 (N_10542,N_8790,N_7679);
nor U10543 (N_10543,N_7797,N_9870);
nand U10544 (N_10544,N_8200,N_9794);
nor U10545 (N_10545,N_9607,N_8406);
xor U10546 (N_10546,N_8560,N_7966);
nor U10547 (N_10547,N_8525,N_8526);
nand U10548 (N_10548,N_9883,N_7664);
and U10549 (N_10549,N_8726,N_8203);
or U10550 (N_10550,N_9756,N_9841);
nor U10551 (N_10551,N_9455,N_9023);
nor U10552 (N_10552,N_7677,N_9937);
nor U10553 (N_10553,N_9153,N_8457);
and U10554 (N_10554,N_9268,N_8366);
or U10555 (N_10555,N_9900,N_8853);
nand U10556 (N_10556,N_9083,N_7789);
nor U10557 (N_10557,N_8772,N_8809);
xor U10558 (N_10558,N_8350,N_7859);
nand U10559 (N_10559,N_7893,N_9907);
and U10560 (N_10560,N_8484,N_7842);
xor U10561 (N_10561,N_9074,N_9905);
and U10562 (N_10562,N_7658,N_8169);
xnor U10563 (N_10563,N_9201,N_9908);
and U10564 (N_10564,N_9265,N_9248);
nor U10565 (N_10565,N_8431,N_8267);
xor U10566 (N_10566,N_8665,N_9518);
or U10567 (N_10567,N_8077,N_9913);
nand U10568 (N_10568,N_8332,N_7631);
xor U10569 (N_10569,N_9895,N_9331);
nand U10570 (N_10570,N_9430,N_8997);
and U10571 (N_10571,N_8495,N_7563);
nand U10572 (N_10572,N_9088,N_8428);
nor U10573 (N_10573,N_8544,N_8756);
nor U10574 (N_10574,N_9631,N_8044);
xnor U10575 (N_10575,N_9285,N_8377);
and U10576 (N_10576,N_9601,N_9617);
xnor U10577 (N_10577,N_7697,N_7903);
and U10578 (N_10578,N_8403,N_9406);
or U10579 (N_10579,N_8474,N_9169);
and U10580 (N_10580,N_9155,N_8593);
or U10581 (N_10581,N_8824,N_7925);
and U10582 (N_10582,N_8442,N_8035);
xor U10583 (N_10583,N_8129,N_7570);
or U10584 (N_10584,N_8262,N_8969);
and U10585 (N_10585,N_9865,N_7729);
and U10586 (N_10586,N_9949,N_8079);
xnor U10587 (N_10587,N_8482,N_9916);
xnor U10588 (N_10588,N_7952,N_8268);
and U10589 (N_10589,N_9428,N_7509);
xor U10590 (N_10590,N_7912,N_7791);
nand U10591 (N_10591,N_8259,N_8588);
xnor U10592 (N_10592,N_9823,N_7999);
and U10593 (N_10593,N_7683,N_8118);
or U10594 (N_10594,N_9478,N_8388);
nor U10595 (N_10595,N_9260,N_9751);
and U10596 (N_10596,N_9693,N_7715);
nand U10597 (N_10597,N_8434,N_9765);
nor U10598 (N_10598,N_8808,N_9213);
or U10599 (N_10599,N_7983,N_8828);
nand U10600 (N_10600,N_9829,N_9553);
nand U10601 (N_10601,N_7613,N_9983);
nor U10602 (N_10602,N_9276,N_8342);
and U10603 (N_10603,N_8448,N_8650);
or U10604 (N_10604,N_8831,N_7958);
xor U10605 (N_10605,N_9532,N_9203);
xnor U10606 (N_10606,N_8038,N_7549);
or U10607 (N_10607,N_7990,N_9752);
and U10608 (N_10608,N_8444,N_8214);
nand U10609 (N_10609,N_8170,N_8227);
nor U10610 (N_10610,N_8900,N_8604);
nor U10611 (N_10611,N_8340,N_8241);
nand U10612 (N_10612,N_8979,N_9958);
and U10613 (N_10613,N_9650,N_8591);
nor U10614 (N_10614,N_9657,N_9360);
nand U10615 (N_10615,N_8274,N_8580);
nand U10616 (N_10616,N_8260,N_8771);
nor U10617 (N_10617,N_9479,N_9714);
or U10618 (N_10618,N_8356,N_9020);
nor U10619 (N_10619,N_7753,N_7909);
nand U10620 (N_10620,N_7739,N_8152);
or U10621 (N_10621,N_8962,N_9193);
nand U10622 (N_10622,N_7657,N_8998);
xnor U10623 (N_10623,N_9573,N_8505);
xnor U10624 (N_10624,N_8514,N_8351);
nor U10625 (N_10625,N_7673,N_9142);
nor U10626 (N_10626,N_9488,N_8003);
nand U10627 (N_10627,N_7854,N_8527);
xnor U10628 (N_10628,N_8613,N_7543);
nor U10629 (N_10629,N_8653,N_7944);
nand U10630 (N_10630,N_9574,N_8488);
or U10631 (N_10631,N_9686,N_9589);
nand U10632 (N_10632,N_8645,N_9312);
nand U10633 (N_10633,N_7953,N_8779);
nor U10634 (N_10634,N_9922,N_9456);
xnor U10635 (N_10635,N_9762,N_9011);
nand U10636 (N_10636,N_8875,N_9364);
or U10637 (N_10637,N_7725,N_8360);
nand U10638 (N_10638,N_8709,N_8424);
nand U10639 (N_10639,N_8441,N_8433);
nand U10640 (N_10640,N_7642,N_8392);
nor U10641 (N_10641,N_9219,N_8887);
and U10642 (N_10642,N_9318,N_8497);
nand U10643 (N_10643,N_8290,N_8080);
or U10644 (N_10644,N_9629,N_9178);
and U10645 (N_10645,N_9771,N_9550);
or U10646 (N_10646,N_9384,N_7810);
or U10647 (N_10647,N_9910,N_8168);
or U10648 (N_10648,N_9730,N_8224);
nor U10649 (N_10649,N_9051,N_8284);
nand U10650 (N_10650,N_8091,N_9716);
xnor U10651 (N_10651,N_8145,N_9140);
or U10652 (N_10652,N_9939,N_9986);
and U10653 (N_10653,N_9090,N_7955);
xor U10654 (N_10654,N_7773,N_9534);
xor U10655 (N_10655,N_9653,N_9658);
and U10656 (N_10656,N_9884,N_9338);
or U10657 (N_10657,N_7795,N_7764);
and U10658 (N_10658,N_7959,N_9690);
and U10659 (N_10659,N_8409,N_8354);
or U10660 (N_10660,N_7848,N_7559);
nand U10661 (N_10661,N_9707,N_9929);
xor U10662 (N_10662,N_8701,N_8892);
nor U10663 (N_10663,N_8084,N_9307);
xor U10664 (N_10664,N_7867,N_8834);
and U10665 (N_10665,N_8039,N_9418);
and U10666 (N_10666,N_9705,N_9885);
xor U10667 (N_10667,N_9245,N_9466);
xnor U10668 (N_10668,N_8971,N_7763);
nor U10669 (N_10669,N_9339,N_7721);
and U10670 (N_10670,N_8616,N_9101);
nor U10671 (N_10671,N_8116,N_7815);
nor U10672 (N_10672,N_9586,N_7581);
nor U10673 (N_10673,N_9987,N_9704);
or U10674 (N_10674,N_7775,N_8996);
nand U10675 (N_10675,N_8679,N_8251);
nor U10676 (N_10676,N_9177,N_7515);
nand U10677 (N_10677,N_8987,N_7531);
nor U10678 (N_10678,N_9086,N_8903);
nand U10679 (N_10679,N_8792,N_9543);
nand U10680 (N_10680,N_9684,N_7670);
nand U10681 (N_10681,N_7617,N_7922);
and U10682 (N_10682,N_9025,N_8764);
and U10683 (N_10683,N_9195,N_8067);
nand U10684 (N_10684,N_8236,N_8045);
and U10685 (N_10685,N_8691,N_9846);
nand U10686 (N_10686,N_7784,N_9396);
and U10687 (N_10687,N_8391,N_7954);
nand U10688 (N_10688,N_9769,N_7542);
xor U10689 (N_10689,N_9286,N_7603);
nor U10690 (N_10690,N_8435,N_9165);
and U10691 (N_10691,N_9787,N_9236);
or U10692 (N_10692,N_8179,N_7883);
xnor U10693 (N_10693,N_7694,N_9001);
or U10694 (N_10694,N_9280,N_9388);
and U10695 (N_10695,N_8871,N_9524);
xnor U10696 (N_10696,N_8942,N_9721);
or U10697 (N_10697,N_8066,N_7600);
xor U10698 (N_10698,N_8308,N_8309);
nand U10699 (N_10699,N_7857,N_9114);
nor U10700 (N_10700,N_8557,N_9317);
or U10701 (N_10701,N_9298,N_7593);
or U10702 (N_10702,N_8139,N_8466);
xor U10703 (N_10703,N_9867,N_7826);
nor U10704 (N_10704,N_8182,N_9848);
nor U10705 (N_10705,N_8280,N_8935);
or U10706 (N_10706,N_9702,N_9063);
or U10707 (N_10707,N_8705,N_9414);
or U10708 (N_10708,N_9627,N_7719);
xor U10709 (N_10709,N_7967,N_8124);
xor U10710 (N_10710,N_7717,N_8844);
nand U10711 (N_10711,N_9622,N_9341);
nor U10712 (N_10712,N_9182,N_7748);
nand U10713 (N_10713,N_7760,N_7813);
nor U10714 (N_10714,N_7946,N_8773);
xnor U10715 (N_10715,N_9281,N_9948);
nand U10716 (N_10716,N_7676,N_8112);
or U10717 (N_10717,N_8362,N_9152);
nor U10718 (N_10718,N_9469,N_7754);
xor U10719 (N_10719,N_9465,N_8187);
xnor U10720 (N_10720,N_9301,N_9410);
nor U10721 (N_10721,N_8857,N_7620);
or U10722 (N_10722,N_8306,N_9037);
or U10723 (N_10723,N_7767,N_7703);
or U10724 (N_10724,N_8397,N_9350);
nand U10725 (N_10725,N_8581,N_7707);
and U10726 (N_10726,N_8555,N_8247);
xnor U10727 (N_10727,N_9425,N_9767);
or U10728 (N_10728,N_8386,N_8050);
nand U10729 (N_10729,N_9806,N_9858);
nor U10730 (N_10730,N_9327,N_9483);
and U10731 (N_10731,N_9240,N_8976);
and U10732 (N_10732,N_9148,N_8127);
xnor U10733 (N_10733,N_8698,N_8589);
or U10734 (N_10734,N_7553,N_9639);
nand U10735 (N_10735,N_8198,N_7534);
xnor U10736 (N_10736,N_8212,N_9619);
xnor U10737 (N_10737,N_8535,N_7849);
and U10738 (N_10738,N_8628,N_9502);
nand U10739 (N_10739,N_9665,N_9678);
xor U10740 (N_10740,N_8498,N_9254);
and U10741 (N_10741,N_8432,N_9542);
xnor U10742 (N_10742,N_7897,N_8513);
nand U10743 (N_10743,N_9512,N_9110);
or U10744 (N_10744,N_8984,N_9510);
nand U10745 (N_10745,N_9995,N_8632);
nor U10746 (N_10746,N_8727,N_8753);
or U10747 (N_10747,N_9789,N_9778);
nor U10748 (N_10748,N_9206,N_7945);
or U10749 (N_10749,N_7560,N_7927);
and U10750 (N_10750,N_8196,N_7988);
and U10751 (N_10751,N_7873,N_8751);
and U10752 (N_10752,N_8685,N_8934);
xor U10753 (N_10753,N_8606,N_7583);
nand U10754 (N_10754,N_7812,N_8502);
and U10755 (N_10755,N_8582,N_8922);
or U10756 (N_10756,N_8507,N_9734);
nor U10757 (N_10757,N_8872,N_8678);
nor U10758 (N_10758,N_9424,N_8147);
and U10759 (N_10759,N_9584,N_7937);
nor U10760 (N_10760,N_9641,N_7785);
or U10761 (N_10761,N_7864,N_7828);
nand U10762 (N_10762,N_7803,N_9015);
and U10763 (N_10763,N_8117,N_8543);
or U10764 (N_10764,N_7994,N_8587);
nand U10765 (N_10765,N_8380,N_8283);
or U10766 (N_10766,N_8197,N_7619);
xnor U10767 (N_10767,N_8506,N_7566);
nor U10768 (N_10768,N_9945,N_7939);
xor U10769 (N_10769,N_7704,N_9035);
xnor U10770 (N_10770,N_9615,N_7932);
nor U10771 (N_10771,N_8423,N_9711);
and U10772 (N_10772,N_8929,N_9798);
nand U10773 (N_10773,N_9009,N_8221);
and U10774 (N_10774,N_7592,N_9107);
xor U10775 (N_10775,N_9218,N_7746);
nor U10776 (N_10776,N_9903,N_9729);
xnor U10777 (N_10777,N_8693,N_7652);
nand U10778 (N_10778,N_9965,N_8733);
nand U10779 (N_10779,N_9917,N_7934);
nand U10780 (N_10780,N_8846,N_7662);
and U10781 (N_10781,N_9597,N_8012);
xnor U10782 (N_10782,N_8085,N_9689);
and U10783 (N_10783,N_9847,N_7882);
nor U10784 (N_10784,N_9229,N_7732);
nor U10785 (N_10785,N_8738,N_8349);
nor U10786 (N_10786,N_7980,N_9859);
and U10787 (N_10787,N_9179,N_9038);
or U10788 (N_10788,N_9947,N_9144);
or U10789 (N_10789,N_7926,N_8323);
nor U10790 (N_10790,N_7567,N_9928);
and U10791 (N_10791,N_9118,N_8171);
xor U10792 (N_10792,N_9058,N_8970);
or U10793 (N_10793,N_8637,N_8743);
nand U10794 (N_10794,N_9974,N_9156);
nor U10795 (N_10795,N_8075,N_9046);
xnor U10796 (N_10796,N_9637,N_9355);
nand U10797 (N_10797,N_8137,N_9606);
xnor U10798 (N_10798,N_7646,N_7801);
nor U10799 (N_10799,N_9190,N_8837);
or U10800 (N_10800,N_9831,N_9018);
or U10801 (N_10801,N_8924,N_8281);
nor U10802 (N_10802,N_8304,N_8389);
and U10803 (N_10803,N_8638,N_9805);
xor U10804 (N_10804,N_7921,N_9437);
nor U10805 (N_10805,N_9070,N_7517);
or U10806 (N_10806,N_8860,N_8459);
nand U10807 (N_10807,N_9056,N_9882);
nand U10808 (N_10808,N_8242,N_9453);
or U10809 (N_10809,N_9294,N_7889);
xnor U10810 (N_10810,N_9575,N_9172);
and U10811 (N_10811,N_7730,N_7629);
xor U10812 (N_10812,N_9695,N_9171);
and U10813 (N_10813,N_8545,N_8303);
and U10814 (N_10814,N_8492,N_8861);
and U10815 (N_10815,N_9220,N_9508);
nand U10816 (N_10816,N_9943,N_8569);
and U10817 (N_10817,N_9836,N_7936);
or U10818 (N_10818,N_8641,N_8859);
xnor U10819 (N_10819,N_8592,N_8657);
xnor U10820 (N_10820,N_8884,N_9441);
or U10821 (N_10821,N_8986,N_8073);
nor U10822 (N_10822,N_7968,N_9255);
nand U10823 (N_10823,N_9912,N_8326);
nand U10824 (N_10824,N_9180,N_8105);
xor U10825 (N_10825,N_8088,N_9391);
xor U10826 (N_10826,N_8659,N_9526);
nor U10827 (N_10827,N_7880,N_8802);
or U10828 (N_10828,N_8205,N_7914);
nand U10829 (N_10829,N_8564,N_8429);
or U10830 (N_10830,N_7626,N_8436);
nor U10831 (N_10831,N_8851,N_8556);
xnor U10832 (N_10832,N_8456,N_9346);
nand U10833 (N_10833,N_8101,N_9098);
nor U10834 (N_10834,N_9890,N_9731);
and U10835 (N_10835,N_9100,N_8939);
nand U10836 (N_10836,N_9963,N_8799);
and U10837 (N_10837,N_7601,N_9111);
nor U10838 (N_10838,N_8620,N_8297);
or U10839 (N_10839,N_8509,N_8481);
xnor U10840 (N_10840,N_7752,N_7535);
or U10841 (N_10841,N_7640,N_8164);
nor U10842 (N_10842,N_8225,N_8288);
nand U10843 (N_10843,N_9808,N_9366);
xnor U10844 (N_10844,N_9802,N_7555);
nand U10845 (N_10845,N_8611,N_9609);
and U10846 (N_10846,N_8142,N_7525);
xnor U10847 (N_10847,N_8548,N_8322);
or U10848 (N_10848,N_7586,N_8517);
nor U10849 (N_10849,N_9158,N_7802);
nor U10850 (N_10850,N_9030,N_7895);
xor U10851 (N_10851,N_9138,N_8845);
xnor U10852 (N_10852,N_9191,N_9856);
or U10853 (N_10853,N_8419,N_8930);
and U10854 (N_10854,N_9244,N_7904);
and U10855 (N_10855,N_7907,N_9611);
nand U10856 (N_10856,N_8625,N_8016);
and U10857 (N_10857,N_8902,N_8006);
or U10858 (N_10858,N_8104,N_7596);
and U10859 (N_10859,N_9898,N_9362);
and U10860 (N_10860,N_8324,N_9112);
nor U10861 (N_10861,N_7671,N_7595);
nand U10862 (N_10862,N_9528,N_8007);
xnor U10863 (N_10863,N_8453,N_8261);
nand U10864 (N_10864,N_8714,N_7841);
or U10865 (N_10865,N_9999,N_7519);
or U10866 (N_10866,N_8383,N_8956);
xor U10867 (N_10867,N_8213,N_9850);
nor U10868 (N_10868,N_9043,N_8717);
xnor U10869 (N_10869,N_8561,N_9828);
or U10870 (N_10870,N_9216,N_8395);
xnor U10871 (N_10871,N_9125,N_7765);
nor U10872 (N_10872,N_7685,N_9468);
nand U10873 (N_10873,N_9925,N_7735);
and U10874 (N_10874,N_7693,N_9875);
and U10875 (N_10875,N_9387,N_7711);
or U10876 (N_10876,N_8454,N_8058);
xor U10877 (N_10877,N_8878,N_8430);
nor U10878 (N_10878,N_7565,N_9039);
or U10879 (N_10879,N_9735,N_7825);
or U10880 (N_10880,N_7609,N_9977);
nand U10881 (N_10881,N_9072,N_9618);
or U10882 (N_10882,N_8438,N_8586);
nand U10883 (N_10883,N_8412,N_9894);
nor U10884 (N_10884,N_9688,N_9426);
xor U10885 (N_10885,N_8830,N_8317);
nor U10886 (N_10886,N_9906,N_8906);
xor U10887 (N_10887,N_9313,N_9150);
and U10888 (N_10888,N_9822,N_9004);
or U10889 (N_10889,N_8056,N_9768);
nand U10890 (N_10890,N_8375,N_8487);
nand U10891 (N_10891,N_7588,N_8648);
nand U10892 (N_10892,N_9600,N_9785);
and U10893 (N_10893,N_9482,N_8302);
nor U10894 (N_10894,N_7689,N_7695);
nand U10895 (N_10895,N_8094,N_7656);
xnor U10896 (N_10896,N_9445,N_7839);
nor U10897 (N_10897,N_9951,N_8387);
or U10898 (N_10898,N_9904,N_9696);
nand U10899 (N_10899,N_9272,N_8975);
and U10900 (N_10900,N_7830,N_8181);
nor U10901 (N_10901,N_7590,N_9746);
or U10902 (N_10902,N_8574,N_8794);
xor U10903 (N_10903,N_8408,N_9065);
and U10904 (N_10904,N_8047,N_9077);
nor U10905 (N_10905,N_9782,N_7823);
or U10906 (N_10906,N_8132,N_8384);
nor U10907 (N_10907,N_8811,N_7758);
and U10908 (N_10908,N_8144,N_8008);
nand U10909 (N_10909,N_8130,N_7872);
or U10910 (N_10910,N_8041,N_9160);
and U10911 (N_10911,N_8644,N_8209);
nor U10912 (N_10912,N_9703,N_9743);
nand U10913 (N_10913,N_9211,N_8803);
or U10914 (N_10914,N_8575,N_8707);
and U10915 (N_10915,N_7780,N_7820);
or U10916 (N_10916,N_9404,N_8829);
and U10917 (N_10917,N_9290,N_9322);
or U10918 (N_10918,N_8255,N_7992);
or U10919 (N_10919,N_8034,N_8051);
nor U10920 (N_10920,N_9305,N_8451);
xnor U10921 (N_10921,N_8528,N_9854);
nor U10922 (N_10922,N_8489,N_8065);
nand U10923 (N_10923,N_9347,N_8013);
xor U10924 (N_10924,N_9113,N_8201);
nor U10925 (N_10925,N_8713,N_8651);
or U10926 (N_10926,N_7906,N_7554);
or U10927 (N_10927,N_9472,N_8855);
nor U10928 (N_10928,N_9498,N_9092);
nand U10929 (N_10929,N_8299,N_9297);
nand U10930 (N_10930,N_7722,N_8925);
xnor U10931 (N_10931,N_8933,N_7508);
nand U10932 (N_10932,N_8469,N_9954);
and U10933 (N_10933,N_8445,N_8275);
or U10934 (N_10934,N_9249,N_9585);
nand U10935 (N_10935,N_9807,N_8909);
nand U10936 (N_10936,N_8795,N_8055);
nand U10937 (N_10937,N_9002,N_9085);
xor U10938 (N_10938,N_9188,N_9754);
nor U10939 (N_10939,N_7916,N_8746);
and U10940 (N_10940,N_8399,N_9192);
nor U10941 (N_10941,N_9814,N_9668);
xnor U10942 (N_10942,N_7700,N_8335);
xor U10943 (N_10943,N_8486,N_8729);
nand U10944 (N_10944,N_9941,N_8994);
nand U10945 (N_10945,N_9628,N_9839);
xor U10946 (N_10946,N_8125,N_9975);
nand U10947 (N_10947,N_7844,N_9032);
and U10948 (N_10948,N_8239,N_8021);
or U10949 (N_10949,N_8176,N_9231);
and U10950 (N_10950,N_8673,N_9973);
xor U10951 (N_10951,N_8352,N_7971);
and U10952 (N_10952,N_7612,N_9259);
and U10953 (N_10953,N_9800,N_7804);
and U10954 (N_10954,N_9563,N_9539);
xnor U10955 (N_10955,N_9357,N_9980);
and U10956 (N_10956,N_9006,N_9145);
xor U10957 (N_10957,N_7923,N_8333);
or U10958 (N_10958,N_9545,N_7833);
nand U10959 (N_10959,N_7772,N_9311);
nor U10960 (N_10960,N_9053,N_8040);
nor U10961 (N_10961,N_8367,N_9351);
xnor U10962 (N_10962,N_7737,N_8881);
nand U10963 (N_10963,N_8895,N_8289);
xnor U10964 (N_10964,N_9197,N_7928);
or U10965 (N_10965,N_8841,N_8960);
xor U10966 (N_10966,N_9050,N_8472);
xnor U10967 (N_10967,N_8740,N_8014);
nor U10968 (N_10968,N_8020,N_7699);
and U10969 (N_10969,N_8188,N_8947);
xor U10970 (N_10970,N_7827,N_8542);
or U10971 (N_10971,N_7987,N_8877);
or U10972 (N_10972,N_8718,N_9810);
or U10973 (N_10973,N_7970,N_8664);
xor U10974 (N_10974,N_7639,N_8285);
nor U10975 (N_10975,N_8252,N_8770);
or U10976 (N_10976,N_8370,N_9984);
nand U10977 (N_10977,N_9962,N_7632);
or U10978 (N_10978,N_9546,N_7768);
and U10979 (N_10979,N_8917,N_8914);
xor U10980 (N_10980,N_9300,N_8656);
xnor U10981 (N_10981,N_9614,N_8516);
nor U10982 (N_10982,N_8920,N_9170);
xor U10983 (N_10983,N_9352,N_9082);
xor U10984 (N_10984,N_9109,N_9667);
nand U10985 (N_10985,N_9610,N_8848);
xor U10986 (N_10986,N_9569,N_9750);
or U10987 (N_10987,N_8763,N_9224);
xor U10988 (N_10988,N_9017,N_8541);
nor U10989 (N_10989,N_9288,N_9664);
nor U10990 (N_10990,N_8043,N_9375);
nor U10991 (N_10991,N_8990,N_9727);
or U10992 (N_10992,N_9520,N_8946);
or U10993 (N_10993,N_7965,N_8193);
xor U10994 (N_10994,N_8775,N_9604);
nand U10995 (N_10995,N_8102,N_7876);
nor U10996 (N_10996,N_7951,N_7778);
and U10997 (N_10997,N_7884,N_9682);
nand U10998 (N_10998,N_9293,N_7759);
nand U10999 (N_10999,N_7877,N_9416);
nor U11000 (N_11000,N_7769,N_7606);
xor U11001 (N_11001,N_9507,N_8672);
and U11002 (N_11002,N_9330,N_7663);
xnor U11003 (N_11003,N_9470,N_7941);
nor U11004 (N_11004,N_7568,N_8814);
xor U11005 (N_11005,N_9748,N_8819);
nor U11006 (N_11006,N_7814,N_7805);
or U11007 (N_11007,N_9651,N_9068);
nand U11008 (N_11008,N_9076,N_8450);
or U11009 (N_11009,N_8172,N_7637);
xnor U11010 (N_11010,N_7989,N_9409);
or U11011 (N_11011,N_9571,N_8533);
nand U11012 (N_11012,N_7635,N_9264);
xor U11013 (N_11013,N_9421,N_8490);
nor U11014 (N_11014,N_8836,N_8886);
and U11015 (N_11015,N_7733,N_9450);
xor U11016 (N_11016,N_7961,N_9725);
or U11017 (N_11017,N_9588,N_7574);
or U11018 (N_11018,N_8107,N_9786);
xnor U11019 (N_11019,N_8460,N_7856);
xor U11020 (N_11020,N_8141,N_8793);
and U11021 (N_11021,N_7520,N_8018);
nand U11022 (N_11022,N_9372,N_8321);
nor U11023 (N_11023,N_7782,N_8185);
or U11024 (N_11024,N_7905,N_8417);
or U11025 (N_11025,N_7728,N_9555);
or U11026 (N_11026,N_7712,N_7654);
or U11027 (N_11027,N_8957,N_8313);
nor U11028 (N_11028,N_7809,N_7962);
and U11029 (N_11029,N_9517,N_8394);
xor U11030 (N_11030,N_7855,N_9239);
nor U11031 (N_11031,N_9103,N_9332);
nor U11032 (N_11032,N_8810,N_8728);
xor U11033 (N_11033,N_8801,N_9640);
or U11034 (N_11034,N_9390,N_8732);
or U11035 (N_11035,N_9477,N_8503);
nor U11036 (N_11036,N_9797,N_9003);
and U11037 (N_11037,N_8004,N_7807);
and U11038 (N_11038,N_8190,N_7623);
and U11039 (N_11039,N_8393,N_8449);
nand U11040 (N_11040,N_7532,N_9084);
nor U11041 (N_11041,N_8676,N_8826);
xor U11042 (N_11042,N_8639,N_7900);
xnor U11043 (N_11043,N_9556,N_9454);
and U11044 (N_11044,N_9097,N_7879);
or U11045 (N_11045,N_8850,N_9433);
and U11046 (N_11046,N_8510,N_9162);
and U11047 (N_11047,N_9970,N_8512);
nor U11048 (N_11048,N_8634,N_7547);
nor U11049 (N_11049,N_8608,N_8702);
xnor U11050 (N_11050,N_8806,N_8276);
nor U11051 (N_11051,N_8462,N_9447);
nand U11052 (N_11052,N_7993,N_8534);
nor U11053 (N_11053,N_9459,N_7528);
nand U11054 (N_11054,N_8005,N_9267);
and U11055 (N_11055,N_9580,N_9719);
xor U11056 (N_11056,N_7920,N_9073);
nand U11057 (N_11057,N_7894,N_8390);
and U11058 (N_11058,N_8156,N_9976);
nand U11059 (N_11059,N_8455,N_9122);
and U11060 (N_11060,N_7548,N_9041);
and U11061 (N_11061,N_8938,N_7698);
xnor U11062 (N_11062,N_8240,N_9774);
nor U11063 (N_11063,N_9358,N_8700);
nor U11064 (N_11064,N_9680,N_9672);
xnor U11065 (N_11065,N_9722,N_9325);
xnor U11066 (N_11066,N_8315,N_7950);
xor U11067 (N_11067,N_9135,N_9214);
nor U11068 (N_11068,N_8798,N_9612);
or U11069 (N_11069,N_8154,N_8149);
nor U11070 (N_11070,N_9981,N_8537);
nor U11071 (N_11071,N_8911,N_9834);
xnor U11072 (N_11072,N_9394,N_8937);
xnor U11073 (N_11073,N_9115,N_8540);
and U11074 (N_11074,N_8312,N_8601);
nand U11075 (N_11075,N_8500,N_8210);
nor U11076 (N_11076,N_9779,N_9257);
and U11077 (N_11077,N_7571,N_8864);
xnor U11078 (N_11078,N_8973,N_8060);
nor U11079 (N_11079,N_9625,N_7913);
and U11080 (N_11080,N_7552,N_9094);
or U11081 (N_11081,N_7648,N_7686);
nand U11082 (N_11082,N_8414,N_8999);
nand U11083 (N_11083,N_8908,N_8968);
or U11084 (N_11084,N_7963,N_8163);
and U11085 (N_11085,N_9432,N_8265);
xnor U11086 (N_11086,N_9159,N_9764);
xor U11087 (N_11087,N_8248,N_9494);
or U11088 (N_11088,N_8670,N_9438);
or U11089 (N_11089,N_8131,N_8953);
xnor U11090 (N_11090,N_8026,N_9726);
xnor U11091 (N_11091,N_8277,N_9675);
xnor U11092 (N_11092,N_9266,N_9844);
or U11093 (N_11093,N_7545,N_8421);
nor U11094 (N_11094,N_9489,N_7644);
nand U11095 (N_11095,N_7516,N_9826);
nand U11096 (N_11096,N_9405,N_9431);
xnor U11097 (N_11097,N_7929,N_8958);
or U11098 (N_11098,N_8256,N_7957);
nor U11099 (N_11099,N_8684,N_8524);
or U11100 (N_11100,N_7774,N_9395);
and U11101 (N_11101,N_8539,N_8074);
nor U11102 (N_11102,N_8270,N_7890);
nor U11103 (N_11103,N_7624,N_8017);
xor U11104 (N_11104,N_7604,N_9181);
xor U11105 (N_11105,N_7511,N_9835);
nor U11106 (N_11106,N_8140,N_7862);
nand U11107 (N_11107,N_9031,N_8821);
nor U11108 (N_11108,N_9377,N_9930);
nor U11109 (N_11109,N_7834,N_8876);
or U11110 (N_11110,N_7706,N_8602);
nor U11111 (N_11111,N_9061,N_9176);
nor U11112 (N_11112,N_8310,N_9340);
nand U11113 (N_11113,N_9921,N_9535);
xnor U11114 (N_11114,N_7533,N_8233);
nor U11115 (N_11115,N_9296,N_9931);
xor U11116 (N_11116,N_9034,N_9969);
or U11117 (N_11117,N_9185,N_8396);
or U11118 (N_11118,N_9278,N_9365);
xor U11119 (N_11119,N_9449,N_9089);
nor U11120 (N_11120,N_8298,N_8504);
or U11121 (N_11121,N_8072,N_7594);
nand U11122 (N_11122,N_7558,N_8633);
nand U11123 (N_11123,N_8036,N_9282);
nand U11124 (N_11124,N_8868,N_8992);
xor U11125 (N_11125,N_8368,N_7850);
xor U11126 (N_11126,N_7835,N_8735);
xnor U11127 (N_11127,N_8760,N_8963);
nand U11128 (N_11128,N_8780,N_8607);
nand U11129 (N_11129,N_8750,N_9570);
nand U11130 (N_11130,N_8440,N_8667);
and U11131 (N_11131,N_8480,N_9060);
xnor U11132 (N_11132,N_8823,N_7643);
or U11133 (N_11133,N_9952,N_7861);
and U11134 (N_11134,N_8951,N_9861);
or U11135 (N_11135,N_7607,N_7718);
and U11136 (N_11136,N_9369,N_8126);
xor U11137 (N_11137,N_9012,N_9595);
nor U11138 (N_11138,N_9106,N_9028);
xor U11139 (N_11139,N_8109,N_8337);
nor U11140 (N_11140,N_9551,N_8162);
nor U11141 (N_11141,N_9880,N_8631);
nand U11142 (N_11142,N_9275,N_8167);
nand U11143 (N_11143,N_7536,N_9096);
nor U11144 (N_11144,N_8890,N_9964);
and U11145 (N_11145,N_8358,N_8204);
xnor U11146 (N_11146,N_9397,N_8478);
and U11147 (N_11147,N_7972,N_7995);
nor U11148 (N_11148,N_8357,N_8880);
xnor U11149 (N_11149,N_7709,N_8754);
or U11150 (N_11150,N_9343,N_9608);
nand U11151 (N_11151,N_8228,N_8597);
and U11152 (N_11152,N_9354,N_9892);
nor U11153 (N_11153,N_8279,N_8465);
and U11154 (N_11154,N_7973,N_8870);
and U11155 (N_11155,N_8621,N_9116);
and U11156 (N_11156,N_8610,N_8663);
and U11157 (N_11157,N_9956,N_8532);
xnor U11158 (N_11158,N_9378,N_7518);
and U11159 (N_11159,N_9052,N_8742);
xor U11160 (N_11160,N_9911,N_8988);
and U11161 (N_11161,N_8037,N_9561);
nand U11162 (N_11162,N_8549,N_9137);
and U11163 (N_11163,N_9630,N_9385);
nand U11164 (N_11164,N_9452,N_9402);
nor U11165 (N_11165,N_9713,N_7522);
xnor U11166 (N_11166,N_7502,N_9087);
nand U11167 (N_11167,N_8991,N_9119);
and U11168 (N_11168,N_8501,N_8230);
and U11169 (N_11169,N_8898,N_8325);
nor U11170 (N_11170,N_9544,N_9463);
and U11171 (N_11171,N_8479,N_8082);
or U11172 (N_11172,N_9994,N_9988);
or U11173 (N_11173,N_8869,N_8761);
nor U11174 (N_11174,N_9644,N_8220);
nor U11175 (N_11175,N_9971,N_9104);
and U11176 (N_11176,N_7734,N_9749);
xor U11177 (N_11177,N_8452,N_7638);
and U11178 (N_11178,N_8086,N_8959);
nor U11179 (N_11179,N_9944,N_8411);
or U11180 (N_11180,N_8447,N_9590);
or U11181 (N_11181,N_8778,N_9602);
nor U11182 (N_11182,N_7745,N_7885);
and U11183 (N_11183,N_8401,N_9803);
xnor U11184 (N_11184,N_9645,N_9326);
nor U11185 (N_11185,N_9697,N_9717);
nand U11186 (N_11186,N_7863,N_7655);
and U11187 (N_11187,N_7969,N_9652);
and U11188 (N_11188,N_9565,N_8972);
or U11189 (N_11189,N_9067,N_9809);
nand U11190 (N_11190,N_8100,N_9579);
and U11191 (N_11191,N_9222,N_8835);
nor U11192 (N_11192,N_8704,N_9783);
xnor U11193 (N_11193,N_8316,N_8000);
nor U11194 (N_11194,N_9757,N_8361);
nand U11195 (N_11195,N_9493,N_8206);
nand U11196 (N_11196,N_7505,N_9566);
nand U11197 (N_11197,N_7682,N_8843);
or U11198 (N_11198,N_9382,N_8936);
xnor U11199 (N_11199,N_8177,N_7744);
xor U11200 (N_11200,N_7524,N_8927);
xor U11201 (N_11201,N_8183,N_8867);
xnor U11202 (N_11202,N_9054,N_9791);
nor U11203 (N_11203,N_8967,N_9194);
nand U11204 (N_11204,N_9940,N_8195);
nand U11205 (N_11205,N_8372,N_9605);
or U11206 (N_11206,N_9064,N_9522);
nor U11207 (N_11207,N_8348,N_7824);
nand U11208 (N_11208,N_8381,N_8822);
nand U11209 (N_11209,N_9560,N_9536);
nand U11210 (N_11210,N_8865,N_8180);
xnor U11211 (N_11211,N_8010,N_7794);
nand U11212 (N_11212,N_9959,N_8053);
nand U11213 (N_11213,N_8098,N_9184);
nand U11214 (N_11214,N_7651,N_8905);
and U11215 (N_11215,N_9513,N_8232);
or U11216 (N_11216,N_8166,N_8552);
xor U11217 (N_11217,N_8940,N_7641);
or U11218 (N_11218,N_8002,N_8151);
and U11219 (N_11219,N_7551,N_8068);
nand U11220 (N_11220,N_9057,N_8103);
nor U11221 (N_11221,N_8295,N_8496);
xnor U11222 (N_11222,N_7669,N_7819);
or U11223 (N_11223,N_7503,N_8161);
and U11224 (N_11224,N_7633,N_7799);
and U11225 (N_11225,N_9147,N_8175);
nand U11226 (N_11226,N_8477,N_7692);
or U11227 (N_11227,N_8873,N_9763);
nand U11228 (N_11228,N_9564,N_8365);
or U11229 (N_11229,N_9813,N_8426);
or U11230 (N_11230,N_7829,N_9010);
xor U11231 (N_11231,N_7874,N_9633);
xnor U11232 (N_11232,N_8571,N_9530);
xnor U11233 (N_11233,N_8813,N_8030);
nand U11234 (N_11234,N_9121,N_9694);
or U11235 (N_11235,N_7940,N_7766);
nand U11236 (N_11236,N_8211,N_8461);
and U11237 (N_11237,N_9036,N_8217);
nand U11238 (N_11238,N_8522,N_8989);
nand U11239 (N_11239,N_8570,N_9819);
and U11240 (N_11240,N_9040,N_7976);
nor U11241 (N_11241,N_9029,N_7691);
nand U11242 (N_11242,N_8619,N_9124);
and U11243 (N_11243,N_9487,N_8553);
nand U11244 (N_11244,N_8437,N_9069);
or U11245 (N_11245,N_8293,N_9632);
nand U11246 (N_11246,N_7902,N_7513);
xor U11247 (N_11247,N_8090,N_8918);
nand U11248 (N_11248,N_8475,N_9497);
and U11249 (N_11249,N_7714,N_9221);
or U11250 (N_11250,N_9973,N_9401);
and U11251 (N_11251,N_8117,N_8941);
nor U11252 (N_11252,N_8980,N_7596);
nor U11253 (N_11253,N_8508,N_9408);
nand U11254 (N_11254,N_8560,N_7522);
nor U11255 (N_11255,N_8789,N_7701);
nor U11256 (N_11256,N_8641,N_7916);
xnor U11257 (N_11257,N_9523,N_9149);
nand U11258 (N_11258,N_9128,N_9229);
xor U11259 (N_11259,N_8733,N_9439);
and U11260 (N_11260,N_9809,N_8625);
and U11261 (N_11261,N_9598,N_8197);
nand U11262 (N_11262,N_8536,N_9727);
and U11263 (N_11263,N_9666,N_8015);
nor U11264 (N_11264,N_9494,N_9297);
nand U11265 (N_11265,N_8284,N_7858);
and U11266 (N_11266,N_7625,N_9608);
nor U11267 (N_11267,N_9885,N_8458);
nor U11268 (N_11268,N_7625,N_9530);
nor U11269 (N_11269,N_8223,N_8864);
and U11270 (N_11270,N_7520,N_9099);
nand U11271 (N_11271,N_9782,N_9832);
nand U11272 (N_11272,N_7776,N_9014);
nand U11273 (N_11273,N_9697,N_8507);
or U11274 (N_11274,N_8188,N_9422);
or U11275 (N_11275,N_8985,N_8871);
xnor U11276 (N_11276,N_7776,N_7719);
nor U11277 (N_11277,N_9219,N_8965);
nand U11278 (N_11278,N_8786,N_7696);
and U11279 (N_11279,N_8897,N_7545);
or U11280 (N_11280,N_9181,N_7730);
xor U11281 (N_11281,N_8274,N_8285);
nand U11282 (N_11282,N_9117,N_8587);
nand U11283 (N_11283,N_9873,N_7700);
or U11284 (N_11284,N_8706,N_7839);
xor U11285 (N_11285,N_7817,N_8607);
nor U11286 (N_11286,N_9429,N_9829);
and U11287 (N_11287,N_8649,N_8550);
nor U11288 (N_11288,N_8513,N_8882);
nand U11289 (N_11289,N_8182,N_7593);
or U11290 (N_11290,N_8973,N_7755);
and U11291 (N_11291,N_9099,N_7938);
nor U11292 (N_11292,N_8562,N_7772);
nand U11293 (N_11293,N_8950,N_9894);
and U11294 (N_11294,N_9002,N_8758);
nor U11295 (N_11295,N_9159,N_8263);
or U11296 (N_11296,N_8664,N_8014);
nand U11297 (N_11297,N_9284,N_9462);
or U11298 (N_11298,N_9672,N_8768);
xnor U11299 (N_11299,N_8707,N_7797);
and U11300 (N_11300,N_8605,N_9640);
nor U11301 (N_11301,N_8850,N_8665);
nor U11302 (N_11302,N_7724,N_9861);
nor U11303 (N_11303,N_8784,N_8715);
nor U11304 (N_11304,N_7907,N_9455);
and U11305 (N_11305,N_8533,N_9356);
and U11306 (N_11306,N_7805,N_7622);
xnor U11307 (N_11307,N_8501,N_9530);
nor U11308 (N_11308,N_9959,N_7724);
and U11309 (N_11309,N_7539,N_9730);
xnor U11310 (N_11310,N_8374,N_8432);
nand U11311 (N_11311,N_8837,N_8377);
xor U11312 (N_11312,N_8630,N_8221);
nand U11313 (N_11313,N_8493,N_9697);
xor U11314 (N_11314,N_8176,N_8386);
or U11315 (N_11315,N_7681,N_8785);
xnor U11316 (N_11316,N_9686,N_9821);
xor U11317 (N_11317,N_9238,N_8547);
nor U11318 (N_11318,N_7922,N_8156);
and U11319 (N_11319,N_8021,N_8632);
nand U11320 (N_11320,N_9231,N_7981);
nor U11321 (N_11321,N_9766,N_9405);
nand U11322 (N_11322,N_9577,N_8718);
nand U11323 (N_11323,N_9638,N_8929);
nand U11324 (N_11324,N_9583,N_8930);
nand U11325 (N_11325,N_8732,N_7819);
and U11326 (N_11326,N_8279,N_8593);
or U11327 (N_11327,N_8025,N_9446);
nor U11328 (N_11328,N_8488,N_8877);
nand U11329 (N_11329,N_9378,N_9031);
and U11330 (N_11330,N_9631,N_9851);
xor U11331 (N_11331,N_7910,N_8400);
xnor U11332 (N_11332,N_7731,N_7591);
xor U11333 (N_11333,N_8869,N_9518);
or U11334 (N_11334,N_7646,N_7906);
xnor U11335 (N_11335,N_8918,N_8472);
or U11336 (N_11336,N_7732,N_9947);
nor U11337 (N_11337,N_9621,N_9347);
nor U11338 (N_11338,N_9061,N_8107);
or U11339 (N_11339,N_8199,N_9968);
nor U11340 (N_11340,N_9669,N_7879);
nand U11341 (N_11341,N_9618,N_8000);
xor U11342 (N_11342,N_8949,N_8524);
xor U11343 (N_11343,N_9815,N_8103);
nand U11344 (N_11344,N_7965,N_9701);
xnor U11345 (N_11345,N_9743,N_9231);
nor U11346 (N_11346,N_7836,N_8490);
xnor U11347 (N_11347,N_8498,N_7951);
and U11348 (N_11348,N_8705,N_8937);
or U11349 (N_11349,N_8862,N_9594);
xor U11350 (N_11350,N_9389,N_9280);
and U11351 (N_11351,N_7916,N_7951);
or U11352 (N_11352,N_7571,N_7804);
or U11353 (N_11353,N_9695,N_9612);
xnor U11354 (N_11354,N_9304,N_9893);
and U11355 (N_11355,N_8040,N_9074);
nor U11356 (N_11356,N_9469,N_7970);
nor U11357 (N_11357,N_8355,N_9050);
nand U11358 (N_11358,N_7686,N_8103);
xnor U11359 (N_11359,N_9683,N_8810);
nor U11360 (N_11360,N_7991,N_7961);
nor U11361 (N_11361,N_9966,N_8532);
xnor U11362 (N_11362,N_8910,N_8257);
and U11363 (N_11363,N_8518,N_7656);
nand U11364 (N_11364,N_7840,N_9539);
and U11365 (N_11365,N_8209,N_9458);
nor U11366 (N_11366,N_9041,N_9141);
nor U11367 (N_11367,N_7834,N_8647);
or U11368 (N_11368,N_9384,N_9256);
xor U11369 (N_11369,N_8006,N_9009);
or U11370 (N_11370,N_7508,N_9671);
or U11371 (N_11371,N_9040,N_8587);
and U11372 (N_11372,N_7842,N_7668);
and U11373 (N_11373,N_9942,N_8927);
xnor U11374 (N_11374,N_9350,N_9417);
nor U11375 (N_11375,N_9478,N_9861);
xor U11376 (N_11376,N_9789,N_9144);
or U11377 (N_11377,N_8812,N_8123);
nand U11378 (N_11378,N_9639,N_9721);
nor U11379 (N_11379,N_8901,N_8405);
or U11380 (N_11380,N_9527,N_9205);
xnor U11381 (N_11381,N_8332,N_7628);
nor U11382 (N_11382,N_9876,N_8373);
nor U11383 (N_11383,N_7641,N_8130);
and U11384 (N_11384,N_9636,N_9393);
nor U11385 (N_11385,N_9109,N_8211);
xnor U11386 (N_11386,N_9511,N_8857);
and U11387 (N_11387,N_8814,N_8539);
nand U11388 (N_11388,N_9881,N_8892);
xor U11389 (N_11389,N_8101,N_9635);
or U11390 (N_11390,N_9449,N_9025);
nand U11391 (N_11391,N_9736,N_7768);
nand U11392 (N_11392,N_8030,N_8384);
nor U11393 (N_11393,N_9473,N_9940);
and U11394 (N_11394,N_9661,N_9658);
nor U11395 (N_11395,N_8304,N_9495);
or U11396 (N_11396,N_9771,N_9514);
and U11397 (N_11397,N_9211,N_7651);
nand U11398 (N_11398,N_7795,N_8630);
nor U11399 (N_11399,N_8873,N_9356);
nand U11400 (N_11400,N_8533,N_9052);
and U11401 (N_11401,N_8771,N_8548);
nor U11402 (N_11402,N_9824,N_8148);
and U11403 (N_11403,N_7851,N_7750);
nand U11404 (N_11404,N_7557,N_8622);
nor U11405 (N_11405,N_9710,N_9823);
or U11406 (N_11406,N_7670,N_9332);
and U11407 (N_11407,N_8274,N_7760);
nor U11408 (N_11408,N_8728,N_7549);
xor U11409 (N_11409,N_9533,N_8980);
xnor U11410 (N_11410,N_9729,N_8714);
nand U11411 (N_11411,N_8250,N_9772);
and U11412 (N_11412,N_7834,N_8278);
nor U11413 (N_11413,N_8439,N_9803);
nand U11414 (N_11414,N_8401,N_8026);
and U11415 (N_11415,N_9917,N_9409);
xnor U11416 (N_11416,N_9148,N_9935);
nor U11417 (N_11417,N_7535,N_9026);
xor U11418 (N_11418,N_9407,N_9647);
xnor U11419 (N_11419,N_9846,N_8657);
nor U11420 (N_11420,N_7994,N_8949);
nor U11421 (N_11421,N_7591,N_7821);
xnor U11422 (N_11422,N_8872,N_8576);
nand U11423 (N_11423,N_9670,N_8139);
nor U11424 (N_11424,N_9621,N_9265);
xnor U11425 (N_11425,N_7990,N_9383);
or U11426 (N_11426,N_7629,N_8556);
or U11427 (N_11427,N_7690,N_9529);
or U11428 (N_11428,N_9223,N_8102);
xnor U11429 (N_11429,N_8502,N_9667);
nor U11430 (N_11430,N_9902,N_8652);
and U11431 (N_11431,N_9776,N_9568);
nand U11432 (N_11432,N_8786,N_9032);
xnor U11433 (N_11433,N_8809,N_7717);
nand U11434 (N_11434,N_8939,N_7565);
xnor U11435 (N_11435,N_9292,N_9501);
nor U11436 (N_11436,N_8043,N_9004);
or U11437 (N_11437,N_7756,N_8317);
or U11438 (N_11438,N_9674,N_7619);
nor U11439 (N_11439,N_9978,N_9062);
xor U11440 (N_11440,N_9759,N_8404);
xnor U11441 (N_11441,N_9430,N_8917);
nor U11442 (N_11442,N_8046,N_9218);
nor U11443 (N_11443,N_9554,N_8572);
nand U11444 (N_11444,N_9661,N_9489);
or U11445 (N_11445,N_7865,N_8102);
nor U11446 (N_11446,N_7963,N_8938);
or U11447 (N_11447,N_7841,N_7628);
xnor U11448 (N_11448,N_9498,N_8183);
nand U11449 (N_11449,N_8674,N_7980);
xor U11450 (N_11450,N_9102,N_8198);
xor U11451 (N_11451,N_7690,N_9372);
nor U11452 (N_11452,N_9457,N_9630);
nor U11453 (N_11453,N_9421,N_7996);
nor U11454 (N_11454,N_9111,N_8186);
xnor U11455 (N_11455,N_8854,N_8761);
and U11456 (N_11456,N_8788,N_9856);
or U11457 (N_11457,N_9021,N_7977);
and U11458 (N_11458,N_7766,N_9977);
xnor U11459 (N_11459,N_8184,N_8704);
and U11460 (N_11460,N_7566,N_7994);
xnor U11461 (N_11461,N_9172,N_9525);
nor U11462 (N_11462,N_9803,N_9800);
nor U11463 (N_11463,N_9614,N_8817);
nand U11464 (N_11464,N_8870,N_8804);
nor U11465 (N_11465,N_9449,N_7892);
and U11466 (N_11466,N_7936,N_8312);
or U11467 (N_11467,N_8964,N_7747);
and U11468 (N_11468,N_8857,N_9668);
and U11469 (N_11469,N_8637,N_9679);
nand U11470 (N_11470,N_9370,N_9606);
nor U11471 (N_11471,N_7860,N_9785);
and U11472 (N_11472,N_9079,N_8652);
xnor U11473 (N_11473,N_8977,N_8837);
nor U11474 (N_11474,N_9314,N_8883);
or U11475 (N_11475,N_9732,N_8172);
and U11476 (N_11476,N_9378,N_9024);
xnor U11477 (N_11477,N_7804,N_8670);
xnor U11478 (N_11478,N_9176,N_9396);
or U11479 (N_11479,N_7543,N_7593);
or U11480 (N_11480,N_9828,N_8951);
or U11481 (N_11481,N_9438,N_8895);
and U11482 (N_11482,N_7927,N_7537);
or U11483 (N_11483,N_9525,N_8444);
and U11484 (N_11484,N_8074,N_9685);
xor U11485 (N_11485,N_9864,N_9256);
nand U11486 (N_11486,N_7584,N_8335);
nor U11487 (N_11487,N_8252,N_9139);
nand U11488 (N_11488,N_8028,N_8700);
nor U11489 (N_11489,N_9816,N_8028);
and U11490 (N_11490,N_9599,N_8420);
and U11491 (N_11491,N_9450,N_8462);
or U11492 (N_11492,N_7563,N_8278);
nor U11493 (N_11493,N_9457,N_8302);
nor U11494 (N_11494,N_7792,N_9746);
or U11495 (N_11495,N_9450,N_9791);
or U11496 (N_11496,N_9500,N_7854);
and U11497 (N_11497,N_7741,N_7538);
nor U11498 (N_11498,N_9647,N_9350);
xnor U11499 (N_11499,N_8237,N_8344);
nand U11500 (N_11500,N_9827,N_8379);
and U11501 (N_11501,N_8767,N_8500);
and U11502 (N_11502,N_9700,N_8359);
xnor U11503 (N_11503,N_9471,N_7804);
nor U11504 (N_11504,N_7562,N_7520);
nand U11505 (N_11505,N_8008,N_8551);
and U11506 (N_11506,N_8563,N_9811);
and U11507 (N_11507,N_7880,N_9355);
or U11508 (N_11508,N_8588,N_9392);
xor U11509 (N_11509,N_7778,N_8335);
xnor U11510 (N_11510,N_9448,N_8000);
or U11511 (N_11511,N_9785,N_7901);
and U11512 (N_11512,N_7941,N_8275);
nor U11513 (N_11513,N_9360,N_9699);
nand U11514 (N_11514,N_9118,N_9397);
xor U11515 (N_11515,N_7502,N_9646);
or U11516 (N_11516,N_7744,N_8113);
xnor U11517 (N_11517,N_8437,N_9327);
or U11518 (N_11518,N_8080,N_9828);
or U11519 (N_11519,N_7563,N_8007);
nand U11520 (N_11520,N_9678,N_8072);
nand U11521 (N_11521,N_8049,N_8276);
nor U11522 (N_11522,N_7767,N_8470);
xnor U11523 (N_11523,N_8049,N_9574);
nand U11524 (N_11524,N_9407,N_7665);
nand U11525 (N_11525,N_9434,N_8358);
and U11526 (N_11526,N_7727,N_7995);
nand U11527 (N_11527,N_8467,N_8100);
or U11528 (N_11528,N_8816,N_8465);
and U11529 (N_11529,N_9250,N_9308);
nand U11530 (N_11530,N_8203,N_9809);
xnor U11531 (N_11531,N_8263,N_9583);
nor U11532 (N_11532,N_9480,N_8562);
xor U11533 (N_11533,N_9510,N_9837);
or U11534 (N_11534,N_9532,N_9910);
nand U11535 (N_11535,N_8812,N_9449);
or U11536 (N_11536,N_8384,N_8290);
nand U11537 (N_11537,N_9831,N_7507);
nor U11538 (N_11538,N_8772,N_9328);
or U11539 (N_11539,N_9324,N_9937);
and U11540 (N_11540,N_7533,N_8730);
nand U11541 (N_11541,N_8995,N_7722);
and U11542 (N_11542,N_9306,N_9205);
xnor U11543 (N_11543,N_8527,N_8832);
xnor U11544 (N_11544,N_8964,N_7672);
xor U11545 (N_11545,N_8680,N_8826);
or U11546 (N_11546,N_9669,N_7719);
xnor U11547 (N_11547,N_7786,N_9336);
and U11548 (N_11548,N_8039,N_9325);
and U11549 (N_11549,N_9435,N_9171);
nor U11550 (N_11550,N_8863,N_7635);
or U11551 (N_11551,N_9473,N_8506);
and U11552 (N_11552,N_7614,N_9675);
nor U11553 (N_11553,N_8738,N_7966);
and U11554 (N_11554,N_9669,N_7549);
nand U11555 (N_11555,N_8224,N_7722);
and U11556 (N_11556,N_9738,N_7720);
and U11557 (N_11557,N_8683,N_8296);
nand U11558 (N_11558,N_8270,N_9338);
and U11559 (N_11559,N_9140,N_9511);
and U11560 (N_11560,N_7716,N_8078);
or U11561 (N_11561,N_8985,N_9165);
or U11562 (N_11562,N_9857,N_7903);
nand U11563 (N_11563,N_9471,N_9230);
nand U11564 (N_11564,N_7739,N_8856);
or U11565 (N_11565,N_8384,N_8455);
and U11566 (N_11566,N_9665,N_8786);
or U11567 (N_11567,N_7895,N_9335);
nand U11568 (N_11568,N_9754,N_8065);
nor U11569 (N_11569,N_9372,N_9454);
xnor U11570 (N_11570,N_8795,N_9518);
or U11571 (N_11571,N_7917,N_9080);
nor U11572 (N_11572,N_8909,N_9190);
or U11573 (N_11573,N_9832,N_9510);
and U11574 (N_11574,N_8500,N_9360);
nor U11575 (N_11575,N_9165,N_8889);
or U11576 (N_11576,N_8786,N_9234);
and U11577 (N_11577,N_7729,N_9206);
or U11578 (N_11578,N_9348,N_8092);
nand U11579 (N_11579,N_8403,N_9841);
or U11580 (N_11580,N_8171,N_8826);
nand U11581 (N_11581,N_8773,N_9886);
or U11582 (N_11582,N_7690,N_8778);
or U11583 (N_11583,N_9835,N_9929);
nor U11584 (N_11584,N_7563,N_7551);
and U11585 (N_11585,N_7696,N_8602);
nor U11586 (N_11586,N_7588,N_8348);
and U11587 (N_11587,N_9270,N_8564);
or U11588 (N_11588,N_8334,N_8928);
nand U11589 (N_11589,N_9042,N_9331);
nand U11590 (N_11590,N_8125,N_8854);
xor U11591 (N_11591,N_8575,N_8027);
and U11592 (N_11592,N_9111,N_9353);
and U11593 (N_11593,N_9624,N_7962);
nor U11594 (N_11594,N_9422,N_8784);
nor U11595 (N_11595,N_9058,N_8888);
and U11596 (N_11596,N_7521,N_9132);
and U11597 (N_11597,N_7733,N_9979);
or U11598 (N_11598,N_7959,N_9276);
or U11599 (N_11599,N_8391,N_8583);
or U11600 (N_11600,N_9740,N_7859);
or U11601 (N_11601,N_8123,N_8796);
nand U11602 (N_11602,N_9505,N_8549);
and U11603 (N_11603,N_8087,N_9217);
xor U11604 (N_11604,N_9273,N_8582);
xor U11605 (N_11605,N_9198,N_7992);
xnor U11606 (N_11606,N_8658,N_8946);
and U11607 (N_11607,N_9350,N_9125);
xnor U11608 (N_11608,N_8399,N_8307);
nor U11609 (N_11609,N_9175,N_8941);
xor U11610 (N_11610,N_7519,N_8190);
or U11611 (N_11611,N_9998,N_8450);
and U11612 (N_11612,N_9660,N_9174);
nand U11613 (N_11613,N_8773,N_8129);
nor U11614 (N_11614,N_9664,N_7968);
and U11615 (N_11615,N_9959,N_8604);
nand U11616 (N_11616,N_7827,N_9207);
or U11617 (N_11617,N_8673,N_7654);
or U11618 (N_11618,N_8141,N_7628);
nand U11619 (N_11619,N_8600,N_7739);
and U11620 (N_11620,N_9529,N_9459);
nand U11621 (N_11621,N_9915,N_8882);
nor U11622 (N_11622,N_7514,N_9929);
nand U11623 (N_11623,N_9717,N_8082);
nor U11624 (N_11624,N_7890,N_8039);
nor U11625 (N_11625,N_8214,N_9555);
xnor U11626 (N_11626,N_9587,N_8750);
xnor U11627 (N_11627,N_8968,N_9616);
or U11628 (N_11628,N_9379,N_9421);
and U11629 (N_11629,N_8092,N_8088);
xor U11630 (N_11630,N_9473,N_9028);
nand U11631 (N_11631,N_9803,N_8651);
nor U11632 (N_11632,N_9247,N_9236);
nand U11633 (N_11633,N_9498,N_9210);
nand U11634 (N_11634,N_7548,N_9240);
xor U11635 (N_11635,N_7508,N_7626);
xnor U11636 (N_11636,N_8275,N_9676);
or U11637 (N_11637,N_9410,N_7603);
or U11638 (N_11638,N_8178,N_9459);
or U11639 (N_11639,N_9044,N_8574);
nand U11640 (N_11640,N_9693,N_9533);
and U11641 (N_11641,N_9741,N_7724);
xor U11642 (N_11642,N_7991,N_8043);
or U11643 (N_11643,N_8905,N_8827);
nor U11644 (N_11644,N_9844,N_9294);
or U11645 (N_11645,N_8181,N_9657);
or U11646 (N_11646,N_8674,N_9111);
and U11647 (N_11647,N_9307,N_8332);
nand U11648 (N_11648,N_8622,N_9435);
nand U11649 (N_11649,N_9802,N_9918);
and U11650 (N_11650,N_9306,N_9279);
and U11651 (N_11651,N_7788,N_8614);
and U11652 (N_11652,N_7527,N_9875);
and U11653 (N_11653,N_9768,N_9706);
xnor U11654 (N_11654,N_8215,N_8920);
nand U11655 (N_11655,N_8121,N_8109);
nor U11656 (N_11656,N_8936,N_9415);
nor U11657 (N_11657,N_7740,N_9099);
xor U11658 (N_11658,N_9716,N_8771);
or U11659 (N_11659,N_9772,N_9135);
nand U11660 (N_11660,N_7900,N_9298);
xnor U11661 (N_11661,N_9247,N_8067);
or U11662 (N_11662,N_8044,N_9956);
nand U11663 (N_11663,N_7597,N_9687);
xnor U11664 (N_11664,N_9041,N_7900);
and U11665 (N_11665,N_8966,N_9130);
or U11666 (N_11666,N_8740,N_9311);
and U11667 (N_11667,N_9282,N_9132);
or U11668 (N_11668,N_8636,N_9329);
nor U11669 (N_11669,N_9279,N_9636);
xnor U11670 (N_11670,N_9922,N_7969);
nor U11671 (N_11671,N_9710,N_7714);
xor U11672 (N_11672,N_8108,N_9265);
nor U11673 (N_11673,N_8593,N_8432);
and U11674 (N_11674,N_9015,N_8765);
xnor U11675 (N_11675,N_8020,N_8316);
nand U11676 (N_11676,N_9163,N_8851);
and U11677 (N_11677,N_9808,N_9227);
or U11678 (N_11678,N_8197,N_8816);
xor U11679 (N_11679,N_9571,N_8102);
xnor U11680 (N_11680,N_8271,N_9245);
nor U11681 (N_11681,N_8342,N_8641);
and U11682 (N_11682,N_7715,N_8071);
nor U11683 (N_11683,N_7781,N_8254);
nor U11684 (N_11684,N_9550,N_7714);
xnor U11685 (N_11685,N_9408,N_9296);
or U11686 (N_11686,N_7855,N_9283);
or U11687 (N_11687,N_9853,N_8770);
or U11688 (N_11688,N_9502,N_8081);
or U11689 (N_11689,N_7653,N_9800);
nor U11690 (N_11690,N_8071,N_9029);
or U11691 (N_11691,N_7993,N_9068);
xnor U11692 (N_11692,N_7948,N_7622);
or U11693 (N_11693,N_9086,N_8410);
or U11694 (N_11694,N_9797,N_9816);
nor U11695 (N_11695,N_7643,N_9063);
nor U11696 (N_11696,N_8517,N_8809);
nor U11697 (N_11697,N_9922,N_7600);
nor U11698 (N_11698,N_9305,N_9520);
xnor U11699 (N_11699,N_7624,N_9979);
nor U11700 (N_11700,N_7738,N_9762);
nor U11701 (N_11701,N_8814,N_9282);
nor U11702 (N_11702,N_8060,N_8084);
nor U11703 (N_11703,N_7550,N_7599);
xnor U11704 (N_11704,N_9806,N_8137);
nand U11705 (N_11705,N_7501,N_8218);
nor U11706 (N_11706,N_8214,N_9344);
xor U11707 (N_11707,N_8160,N_8529);
xor U11708 (N_11708,N_8763,N_9495);
nor U11709 (N_11709,N_8086,N_9442);
or U11710 (N_11710,N_9908,N_8100);
and U11711 (N_11711,N_9032,N_8850);
xnor U11712 (N_11712,N_8194,N_8002);
and U11713 (N_11713,N_9290,N_8648);
nand U11714 (N_11714,N_8874,N_8186);
nor U11715 (N_11715,N_8804,N_7756);
xnor U11716 (N_11716,N_8028,N_8434);
nor U11717 (N_11717,N_9451,N_9880);
nand U11718 (N_11718,N_9226,N_7809);
nor U11719 (N_11719,N_9987,N_9496);
or U11720 (N_11720,N_7971,N_8504);
xnor U11721 (N_11721,N_9808,N_8726);
xnor U11722 (N_11722,N_8108,N_9216);
nor U11723 (N_11723,N_7574,N_8324);
nor U11724 (N_11724,N_7858,N_8916);
nand U11725 (N_11725,N_9972,N_9084);
and U11726 (N_11726,N_9235,N_8646);
or U11727 (N_11727,N_9899,N_8194);
xor U11728 (N_11728,N_8866,N_8239);
nand U11729 (N_11729,N_9272,N_7989);
or U11730 (N_11730,N_9312,N_8832);
or U11731 (N_11731,N_8008,N_9295);
xor U11732 (N_11732,N_9747,N_9945);
nor U11733 (N_11733,N_8178,N_8355);
nand U11734 (N_11734,N_8479,N_9423);
and U11735 (N_11735,N_8116,N_9032);
nand U11736 (N_11736,N_9793,N_9752);
xnor U11737 (N_11737,N_7922,N_9844);
and U11738 (N_11738,N_7681,N_8446);
xnor U11739 (N_11739,N_7660,N_9191);
nor U11740 (N_11740,N_7609,N_8062);
xor U11741 (N_11741,N_9551,N_9742);
xor U11742 (N_11742,N_8641,N_9664);
nand U11743 (N_11743,N_8689,N_7516);
nand U11744 (N_11744,N_9128,N_9631);
nor U11745 (N_11745,N_9322,N_7582);
or U11746 (N_11746,N_7986,N_9595);
or U11747 (N_11747,N_8536,N_8334);
and U11748 (N_11748,N_9798,N_8004);
xor U11749 (N_11749,N_9109,N_9308);
nor U11750 (N_11750,N_7615,N_8297);
xor U11751 (N_11751,N_9346,N_9378);
xnor U11752 (N_11752,N_7744,N_9926);
and U11753 (N_11753,N_7761,N_7977);
nand U11754 (N_11754,N_9465,N_9192);
nand U11755 (N_11755,N_9940,N_9906);
or U11756 (N_11756,N_7594,N_9467);
nor U11757 (N_11757,N_8148,N_9698);
nor U11758 (N_11758,N_8286,N_9133);
and U11759 (N_11759,N_7932,N_9963);
nand U11760 (N_11760,N_7893,N_7627);
or U11761 (N_11761,N_8902,N_9552);
nand U11762 (N_11762,N_7621,N_9438);
or U11763 (N_11763,N_8363,N_7538);
nand U11764 (N_11764,N_9420,N_9543);
nor U11765 (N_11765,N_9706,N_8433);
and U11766 (N_11766,N_9668,N_8078);
and U11767 (N_11767,N_8215,N_8981);
nand U11768 (N_11768,N_9103,N_9439);
xor U11769 (N_11769,N_9940,N_9201);
or U11770 (N_11770,N_9359,N_9808);
nand U11771 (N_11771,N_8531,N_9450);
and U11772 (N_11772,N_9037,N_7580);
nand U11773 (N_11773,N_9399,N_9292);
xor U11774 (N_11774,N_8467,N_9156);
nand U11775 (N_11775,N_7602,N_8027);
and U11776 (N_11776,N_8259,N_8069);
and U11777 (N_11777,N_7874,N_9910);
xor U11778 (N_11778,N_8430,N_9162);
nor U11779 (N_11779,N_9798,N_9820);
and U11780 (N_11780,N_9079,N_8806);
xnor U11781 (N_11781,N_8612,N_8870);
and U11782 (N_11782,N_7652,N_9197);
and U11783 (N_11783,N_9250,N_7542);
nand U11784 (N_11784,N_8215,N_7873);
and U11785 (N_11785,N_8560,N_9322);
xor U11786 (N_11786,N_9460,N_9292);
nand U11787 (N_11787,N_7556,N_7772);
and U11788 (N_11788,N_8138,N_8179);
nor U11789 (N_11789,N_8505,N_8330);
and U11790 (N_11790,N_9552,N_8288);
nor U11791 (N_11791,N_8546,N_8800);
xor U11792 (N_11792,N_8533,N_7654);
and U11793 (N_11793,N_7691,N_8997);
or U11794 (N_11794,N_9138,N_8680);
and U11795 (N_11795,N_8285,N_8192);
nand U11796 (N_11796,N_8625,N_8286);
nand U11797 (N_11797,N_7563,N_9766);
nor U11798 (N_11798,N_9640,N_8441);
nand U11799 (N_11799,N_9040,N_8267);
nor U11800 (N_11800,N_7812,N_9014);
xor U11801 (N_11801,N_7867,N_7978);
nor U11802 (N_11802,N_8695,N_9719);
nand U11803 (N_11803,N_8414,N_7876);
and U11804 (N_11804,N_8094,N_8340);
nor U11805 (N_11805,N_9336,N_9669);
nand U11806 (N_11806,N_8053,N_7881);
nand U11807 (N_11807,N_9366,N_9823);
nand U11808 (N_11808,N_9545,N_7552);
nand U11809 (N_11809,N_8426,N_8352);
nand U11810 (N_11810,N_9773,N_8502);
or U11811 (N_11811,N_8796,N_8206);
or U11812 (N_11812,N_9296,N_7673);
and U11813 (N_11813,N_8656,N_9439);
nand U11814 (N_11814,N_8480,N_9486);
nor U11815 (N_11815,N_8403,N_9123);
nand U11816 (N_11816,N_8915,N_8176);
xor U11817 (N_11817,N_8732,N_9762);
nor U11818 (N_11818,N_7690,N_9923);
nor U11819 (N_11819,N_7769,N_9862);
or U11820 (N_11820,N_8869,N_8074);
or U11821 (N_11821,N_7840,N_9902);
nand U11822 (N_11822,N_9814,N_8045);
and U11823 (N_11823,N_7844,N_8092);
and U11824 (N_11824,N_9645,N_9202);
nor U11825 (N_11825,N_9892,N_8748);
or U11826 (N_11826,N_8334,N_7899);
nor U11827 (N_11827,N_7933,N_9224);
nor U11828 (N_11828,N_9538,N_8427);
or U11829 (N_11829,N_9456,N_7627);
and U11830 (N_11830,N_7500,N_8255);
and U11831 (N_11831,N_9376,N_8592);
nand U11832 (N_11832,N_7621,N_9533);
nor U11833 (N_11833,N_8632,N_8035);
or U11834 (N_11834,N_9668,N_9583);
nand U11835 (N_11835,N_9813,N_8008);
and U11836 (N_11836,N_7870,N_9634);
xor U11837 (N_11837,N_9064,N_7538);
or U11838 (N_11838,N_9450,N_8196);
or U11839 (N_11839,N_9044,N_9149);
nor U11840 (N_11840,N_8594,N_9855);
and U11841 (N_11841,N_9266,N_8562);
nand U11842 (N_11842,N_9237,N_8549);
and U11843 (N_11843,N_8612,N_9179);
and U11844 (N_11844,N_9452,N_8710);
nor U11845 (N_11845,N_7817,N_8098);
or U11846 (N_11846,N_8077,N_8828);
and U11847 (N_11847,N_8455,N_8202);
xnor U11848 (N_11848,N_9481,N_8760);
xnor U11849 (N_11849,N_9927,N_8679);
xnor U11850 (N_11850,N_9474,N_9190);
xnor U11851 (N_11851,N_8419,N_8007);
xor U11852 (N_11852,N_7989,N_8075);
xnor U11853 (N_11853,N_9218,N_8578);
xnor U11854 (N_11854,N_9918,N_9011);
or U11855 (N_11855,N_8581,N_9832);
xnor U11856 (N_11856,N_9669,N_8393);
nand U11857 (N_11857,N_7878,N_8494);
and U11858 (N_11858,N_8659,N_9273);
or U11859 (N_11859,N_9413,N_9373);
xnor U11860 (N_11860,N_8902,N_7520);
nor U11861 (N_11861,N_8351,N_9344);
xor U11862 (N_11862,N_8438,N_7982);
xor U11863 (N_11863,N_9059,N_9413);
xor U11864 (N_11864,N_9163,N_8154);
or U11865 (N_11865,N_8199,N_9528);
xor U11866 (N_11866,N_9787,N_8455);
xnor U11867 (N_11867,N_9571,N_9869);
nor U11868 (N_11868,N_8747,N_9743);
or U11869 (N_11869,N_8302,N_8747);
and U11870 (N_11870,N_9213,N_9834);
or U11871 (N_11871,N_8483,N_9477);
and U11872 (N_11872,N_7756,N_8632);
nand U11873 (N_11873,N_7656,N_9576);
or U11874 (N_11874,N_9258,N_7709);
nor U11875 (N_11875,N_9435,N_8738);
nor U11876 (N_11876,N_8554,N_7814);
nor U11877 (N_11877,N_7923,N_8496);
nor U11878 (N_11878,N_9810,N_8725);
and U11879 (N_11879,N_9099,N_9384);
or U11880 (N_11880,N_9007,N_8918);
and U11881 (N_11881,N_9803,N_9234);
or U11882 (N_11882,N_9574,N_8135);
xnor U11883 (N_11883,N_7616,N_9092);
and U11884 (N_11884,N_9182,N_9691);
nand U11885 (N_11885,N_8696,N_8183);
and U11886 (N_11886,N_9107,N_7805);
nor U11887 (N_11887,N_8708,N_8903);
xor U11888 (N_11888,N_9888,N_7722);
xor U11889 (N_11889,N_9802,N_9861);
xnor U11890 (N_11890,N_9961,N_9696);
nor U11891 (N_11891,N_8455,N_9974);
nor U11892 (N_11892,N_7559,N_7720);
xor U11893 (N_11893,N_8221,N_8391);
nand U11894 (N_11894,N_9046,N_7735);
nor U11895 (N_11895,N_9301,N_8738);
xor U11896 (N_11896,N_8892,N_9233);
and U11897 (N_11897,N_7516,N_9425);
nand U11898 (N_11898,N_8531,N_8167);
nand U11899 (N_11899,N_9833,N_9452);
nor U11900 (N_11900,N_7675,N_9678);
or U11901 (N_11901,N_9329,N_9172);
or U11902 (N_11902,N_9254,N_7544);
nor U11903 (N_11903,N_9926,N_7569);
and U11904 (N_11904,N_9891,N_8280);
or U11905 (N_11905,N_8137,N_8082);
nor U11906 (N_11906,N_9271,N_7615);
xnor U11907 (N_11907,N_9486,N_8076);
nor U11908 (N_11908,N_9922,N_9439);
or U11909 (N_11909,N_8882,N_8010);
and U11910 (N_11910,N_7994,N_8598);
nor U11911 (N_11911,N_8380,N_9166);
nand U11912 (N_11912,N_8204,N_8568);
xnor U11913 (N_11913,N_8600,N_7794);
or U11914 (N_11914,N_8080,N_8872);
and U11915 (N_11915,N_7596,N_9724);
and U11916 (N_11916,N_7731,N_8032);
and U11917 (N_11917,N_9532,N_9201);
nor U11918 (N_11918,N_8209,N_8982);
and U11919 (N_11919,N_9610,N_7669);
or U11920 (N_11920,N_9623,N_8258);
and U11921 (N_11921,N_9287,N_9844);
nor U11922 (N_11922,N_7506,N_9300);
and U11923 (N_11923,N_9607,N_8996);
and U11924 (N_11924,N_7518,N_8678);
xnor U11925 (N_11925,N_8292,N_8029);
xor U11926 (N_11926,N_8330,N_7641);
nor U11927 (N_11927,N_9133,N_9279);
and U11928 (N_11928,N_7604,N_9750);
nor U11929 (N_11929,N_9709,N_8749);
or U11930 (N_11930,N_9464,N_9047);
xor U11931 (N_11931,N_7903,N_7737);
nor U11932 (N_11932,N_9372,N_9044);
xnor U11933 (N_11933,N_7683,N_9154);
nor U11934 (N_11934,N_8546,N_7658);
or U11935 (N_11935,N_8121,N_9931);
nand U11936 (N_11936,N_9440,N_9662);
nor U11937 (N_11937,N_8436,N_8137);
nand U11938 (N_11938,N_9508,N_8063);
nand U11939 (N_11939,N_8624,N_9874);
and U11940 (N_11940,N_7790,N_8116);
and U11941 (N_11941,N_8774,N_9537);
or U11942 (N_11942,N_7759,N_9123);
nand U11943 (N_11943,N_9447,N_9492);
xnor U11944 (N_11944,N_8157,N_9791);
nand U11945 (N_11945,N_9289,N_9398);
nand U11946 (N_11946,N_8841,N_7871);
and U11947 (N_11947,N_9952,N_9397);
nor U11948 (N_11948,N_9302,N_9030);
nor U11949 (N_11949,N_9861,N_7796);
or U11950 (N_11950,N_8767,N_8114);
xor U11951 (N_11951,N_9640,N_9087);
xor U11952 (N_11952,N_8650,N_9456);
and U11953 (N_11953,N_8815,N_7613);
and U11954 (N_11954,N_9188,N_7850);
xnor U11955 (N_11955,N_9038,N_8581);
nand U11956 (N_11956,N_8213,N_9390);
or U11957 (N_11957,N_8494,N_8338);
xnor U11958 (N_11958,N_8122,N_8808);
nand U11959 (N_11959,N_7745,N_8650);
nand U11960 (N_11960,N_8176,N_8571);
and U11961 (N_11961,N_9726,N_8908);
xnor U11962 (N_11962,N_8146,N_7871);
nor U11963 (N_11963,N_9967,N_9352);
nand U11964 (N_11964,N_8466,N_9188);
xor U11965 (N_11965,N_9909,N_9111);
and U11966 (N_11966,N_7889,N_9931);
and U11967 (N_11967,N_9788,N_7854);
nand U11968 (N_11968,N_9217,N_9308);
xnor U11969 (N_11969,N_7597,N_8879);
nor U11970 (N_11970,N_7532,N_9629);
and U11971 (N_11971,N_9851,N_8084);
nand U11972 (N_11972,N_7712,N_8935);
nor U11973 (N_11973,N_9987,N_7946);
nor U11974 (N_11974,N_9502,N_7692);
nand U11975 (N_11975,N_9917,N_9721);
nand U11976 (N_11976,N_8975,N_9914);
nand U11977 (N_11977,N_8100,N_8150);
xnor U11978 (N_11978,N_9065,N_7715);
nand U11979 (N_11979,N_8287,N_8445);
xor U11980 (N_11980,N_8631,N_7608);
xor U11981 (N_11981,N_8890,N_8003);
nand U11982 (N_11982,N_8083,N_9855);
nor U11983 (N_11983,N_8094,N_8898);
xnor U11984 (N_11984,N_9620,N_7526);
nor U11985 (N_11985,N_9870,N_9046);
xor U11986 (N_11986,N_9811,N_8709);
and U11987 (N_11987,N_9052,N_9005);
or U11988 (N_11988,N_8951,N_8233);
nand U11989 (N_11989,N_8130,N_9368);
or U11990 (N_11990,N_8107,N_9847);
nor U11991 (N_11991,N_9028,N_8508);
xnor U11992 (N_11992,N_9663,N_9939);
xor U11993 (N_11993,N_9349,N_9141);
xnor U11994 (N_11994,N_8613,N_9983);
nand U11995 (N_11995,N_7707,N_9590);
nand U11996 (N_11996,N_7519,N_9959);
nor U11997 (N_11997,N_7517,N_8482);
and U11998 (N_11998,N_9929,N_8425);
xnor U11999 (N_11999,N_8457,N_7759);
and U12000 (N_12000,N_7722,N_8294);
or U12001 (N_12001,N_9024,N_9690);
or U12002 (N_12002,N_9060,N_8892);
or U12003 (N_12003,N_9907,N_9533);
xor U12004 (N_12004,N_9117,N_9384);
nand U12005 (N_12005,N_7782,N_7565);
nand U12006 (N_12006,N_8698,N_7719);
xor U12007 (N_12007,N_7584,N_7737);
xor U12008 (N_12008,N_9470,N_9826);
nand U12009 (N_12009,N_9828,N_8111);
or U12010 (N_12010,N_7500,N_8877);
or U12011 (N_12011,N_8805,N_7950);
and U12012 (N_12012,N_8732,N_7985);
xnor U12013 (N_12013,N_8696,N_9965);
and U12014 (N_12014,N_9084,N_9668);
or U12015 (N_12015,N_9761,N_9168);
xor U12016 (N_12016,N_9411,N_9012);
xnor U12017 (N_12017,N_8451,N_8610);
nand U12018 (N_12018,N_8356,N_8940);
xnor U12019 (N_12019,N_9681,N_9148);
xnor U12020 (N_12020,N_7500,N_8427);
xnor U12021 (N_12021,N_7537,N_7867);
nand U12022 (N_12022,N_9633,N_9562);
xor U12023 (N_12023,N_9256,N_8146);
and U12024 (N_12024,N_9032,N_9502);
xor U12025 (N_12025,N_8160,N_8784);
or U12026 (N_12026,N_9276,N_9062);
nor U12027 (N_12027,N_8759,N_7649);
or U12028 (N_12028,N_9987,N_8943);
xor U12029 (N_12029,N_9418,N_8486);
or U12030 (N_12030,N_8311,N_7730);
and U12031 (N_12031,N_9365,N_9142);
xnor U12032 (N_12032,N_8108,N_7502);
nor U12033 (N_12033,N_9741,N_8063);
or U12034 (N_12034,N_9331,N_8430);
xor U12035 (N_12035,N_8198,N_8894);
nor U12036 (N_12036,N_7912,N_9760);
nor U12037 (N_12037,N_8225,N_8189);
nor U12038 (N_12038,N_9120,N_9604);
nor U12039 (N_12039,N_8005,N_8174);
nand U12040 (N_12040,N_8592,N_9640);
nor U12041 (N_12041,N_7636,N_7785);
or U12042 (N_12042,N_9526,N_9521);
and U12043 (N_12043,N_8953,N_7672);
nor U12044 (N_12044,N_9431,N_8544);
nor U12045 (N_12045,N_8228,N_9332);
nor U12046 (N_12046,N_9977,N_9545);
and U12047 (N_12047,N_8301,N_9672);
or U12048 (N_12048,N_9031,N_8077);
xnor U12049 (N_12049,N_7856,N_9451);
nand U12050 (N_12050,N_8330,N_8770);
nand U12051 (N_12051,N_8063,N_9677);
xor U12052 (N_12052,N_8272,N_9844);
or U12053 (N_12053,N_9856,N_8966);
nand U12054 (N_12054,N_8644,N_7848);
or U12055 (N_12055,N_7973,N_9368);
nor U12056 (N_12056,N_8774,N_8805);
nand U12057 (N_12057,N_9732,N_9927);
xor U12058 (N_12058,N_9464,N_9847);
xnor U12059 (N_12059,N_8298,N_9607);
xor U12060 (N_12060,N_9805,N_9938);
nand U12061 (N_12061,N_9795,N_8699);
nor U12062 (N_12062,N_7900,N_7956);
or U12063 (N_12063,N_8177,N_8183);
xnor U12064 (N_12064,N_7911,N_8094);
and U12065 (N_12065,N_9032,N_9000);
nor U12066 (N_12066,N_7652,N_8318);
nor U12067 (N_12067,N_9485,N_9323);
and U12068 (N_12068,N_8862,N_8715);
xor U12069 (N_12069,N_9010,N_9433);
nor U12070 (N_12070,N_8003,N_7529);
nor U12071 (N_12071,N_7972,N_8947);
nand U12072 (N_12072,N_8808,N_9332);
nor U12073 (N_12073,N_9955,N_8287);
xnor U12074 (N_12074,N_8058,N_9074);
xor U12075 (N_12075,N_9892,N_7593);
nor U12076 (N_12076,N_8124,N_9284);
or U12077 (N_12077,N_8397,N_7816);
xnor U12078 (N_12078,N_9124,N_9153);
and U12079 (N_12079,N_9599,N_9979);
or U12080 (N_12080,N_7518,N_8423);
nor U12081 (N_12081,N_8331,N_9677);
or U12082 (N_12082,N_9283,N_8102);
xor U12083 (N_12083,N_8528,N_8603);
xnor U12084 (N_12084,N_8330,N_9052);
or U12085 (N_12085,N_7974,N_8927);
nor U12086 (N_12086,N_9653,N_8640);
xor U12087 (N_12087,N_8778,N_7681);
nand U12088 (N_12088,N_9687,N_8606);
and U12089 (N_12089,N_9634,N_8897);
nand U12090 (N_12090,N_9121,N_9308);
xor U12091 (N_12091,N_9466,N_9459);
and U12092 (N_12092,N_9371,N_7658);
nand U12093 (N_12093,N_7869,N_9649);
nand U12094 (N_12094,N_7648,N_9399);
or U12095 (N_12095,N_8198,N_8796);
and U12096 (N_12096,N_8019,N_9607);
or U12097 (N_12097,N_9456,N_8222);
nand U12098 (N_12098,N_9595,N_8029);
nand U12099 (N_12099,N_9673,N_8922);
nand U12100 (N_12100,N_9817,N_7995);
xor U12101 (N_12101,N_7820,N_9353);
nor U12102 (N_12102,N_7942,N_8736);
xnor U12103 (N_12103,N_7999,N_9367);
or U12104 (N_12104,N_9950,N_9420);
nor U12105 (N_12105,N_8003,N_9122);
nor U12106 (N_12106,N_8699,N_8927);
xor U12107 (N_12107,N_8962,N_7992);
and U12108 (N_12108,N_8013,N_8853);
and U12109 (N_12109,N_7793,N_7821);
xnor U12110 (N_12110,N_9465,N_9187);
nor U12111 (N_12111,N_9105,N_8391);
nor U12112 (N_12112,N_7791,N_8956);
xnor U12113 (N_12113,N_8990,N_9014);
nor U12114 (N_12114,N_9654,N_9859);
and U12115 (N_12115,N_9849,N_8178);
and U12116 (N_12116,N_8358,N_8579);
nor U12117 (N_12117,N_7804,N_9904);
and U12118 (N_12118,N_7817,N_7516);
or U12119 (N_12119,N_7739,N_9255);
or U12120 (N_12120,N_9578,N_7781);
and U12121 (N_12121,N_9439,N_9078);
nand U12122 (N_12122,N_8202,N_9532);
nor U12123 (N_12123,N_8861,N_9662);
nor U12124 (N_12124,N_8295,N_9092);
xnor U12125 (N_12125,N_8104,N_8494);
nor U12126 (N_12126,N_8299,N_7789);
nor U12127 (N_12127,N_9935,N_8906);
xor U12128 (N_12128,N_8267,N_8645);
or U12129 (N_12129,N_9770,N_9601);
and U12130 (N_12130,N_8935,N_9244);
and U12131 (N_12131,N_7844,N_7578);
or U12132 (N_12132,N_9274,N_9775);
nand U12133 (N_12133,N_8953,N_7722);
nor U12134 (N_12134,N_8215,N_8993);
or U12135 (N_12135,N_9625,N_8756);
nor U12136 (N_12136,N_9719,N_9107);
or U12137 (N_12137,N_9161,N_9674);
nor U12138 (N_12138,N_9997,N_9216);
nor U12139 (N_12139,N_8397,N_8727);
nor U12140 (N_12140,N_8751,N_9523);
nand U12141 (N_12141,N_9552,N_7842);
nor U12142 (N_12142,N_9834,N_9182);
nand U12143 (N_12143,N_9882,N_7556);
nor U12144 (N_12144,N_7979,N_8763);
nor U12145 (N_12145,N_7975,N_9984);
or U12146 (N_12146,N_8302,N_8984);
nor U12147 (N_12147,N_7871,N_8944);
nor U12148 (N_12148,N_7550,N_8333);
or U12149 (N_12149,N_9698,N_9787);
and U12150 (N_12150,N_9322,N_8200);
nor U12151 (N_12151,N_8020,N_9328);
nand U12152 (N_12152,N_9380,N_9221);
nor U12153 (N_12153,N_9828,N_8555);
and U12154 (N_12154,N_9128,N_9692);
or U12155 (N_12155,N_7740,N_9869);
and U12156 (N_12156,N_9183,N_9561);
or U12157 (N_12157,N_8876,N_8106);
nand U12158 (N_12158,N_8733,N_9763);
xnor U12159 (N_12159,N_8918,N_9085);
xor U12160 (N_12160,N_8270,N_7921);
xnor U12161 (N_12161,N_9952,N_8914);
nor U12162 (N_12162,N_9838,N_8028);
nand U12163 (N_12163,N_8329,N_8915);
xnor U12164 (N_12164,N_9613,N_8093);
nor U12165 (N_12165,N_9714,N_9455);
xnor U12166 (N_12166,N_8916,N_8344);
xor U12167 (N_12167,N_8768,N_7642);
or U12168 (N_12168,N_9247,N_9200);
xnor U12169 (N_12169,N_9140,N_9565);
xnor U12170 (N_12170,N_9616,N_9738);
and U12171 (N_12171,N_8699,N_8033);
and U12172 (N_12172,N_8475,N_8626);
or U12173 (N_12173,N_8444,N_7725);
nand U12174 (N_12174,N_8911,N_9724);
or U12175 (N_12175,N_7595,N_9096);
nor U12176 (N_12176,N_7908,N_9652);
nor U12177 (N_12177,N_7907,N_8218);
and U12178 (N_12178,N_9780,N_9091);
and U12179 (N_12179,N_8692,N_9398);
nand U12180 (N_12180,N_7572,N_9986);
nor U12181 (N_12181,N_8170,N_8949);
nand U12182 (N_12182,N_8391,N_9069);
xor U12183 (N_12183,N_9303,N_8692);
xnor U12184 (N_12184,N_8202,N_9221);
xor U12185 (N_12185,N_9164,N_9902);
and U12186 (N_12186,N_7827,N_7628);
xnor U12187 (N_12187,N_9392,N_9510);
nor U12188 (N_12188,N_9611,N_9750);
or U12189 (N_12189,N_9224,N_8586);
and U12190 (N_12190,N_9454,N_7521);
and U12191 (N_12191,N_9116,N_9192);
or U12192 (N_12192,N_8844,N_9422);
or U12193 (N_12193,N_9935,N_9045);
nand U12194 (N_12194,N_8769,N_9228);
nor U12195 (N_12195,N_8204,N_9484);
nand U12196 (N_12196,N_8778,N_8883);
nor U12197 (N_12197,N_7917,N_9599);
or U12198 (N_12198,N_8128,N_8653);
and U12199 (N_12199,N_9914,N_8546);
or U12200 (N_12200,N_9377,N_8220);
nand U12201 (N_12201,N_8539,N_7776);
xnor U12202 (N_12202,N_9483,N_7668);
nor U12203 (N_12203,N_8540,N_8191);
or U12204 (N_12204,N_9726,N_8835);
nor U12205 (N_12205,N_8843,N_8785);
and U12206 (N_12206,N_7534,N_8958);
or U12207 (N_12207,N_8089,N_7529);
and U12208 (N_12208,N_8023,N_9853);
nor U12209 (N_12209,N_7986,N_8265);
or U12210 (N_12210,N_8824,N_8290);
nor U12211 (N_12211,N_9225,N_9898);
or U12212 (N_12212,N_9450,N_9788);
nand U12213 (N_12213,N_8219,N_9284);
and U12214 (N_12214,N_9429,N_8288);
and U12215 (N_12215,N_9125,N_8881);
nand U12216 (N_12216,N_8888,N_8799);
and U12217 (N_12217,N_8521,N_7662);
and U12218 (N_12218,N_9444,N_8268);
or U12219 (N_12219,N_8591,N_9059);
nand U12220 (N_12220,N_8257,N_8174);
xnor U12221 (N_12221,N_9415,N_9727);
nand U12222 (N_12222,N_7713,N_9094);
xor U12223 (N_12223,N_8350,N_8368);
nor U12224 (N_12224,N_8419,N_9600);
nand U12225 (N_12225,N_8468,N_8247);
xor U12226 (N_12226,N_8881,N_7710);
and U12227 (N_12227,N_7556,N_7710);
xnor U12228 (N_12228,N_8351,N_9782);
nand U12229 (N_12229,N_8318,N_8217);
or U12230 (N_12230,N_9366,N_9471);
or U12231 (N_12231,N_7988,N_8168);
or U12232 (N_12232,N_8020,N_8449);
nor U12233 (N_12233,N_8972,N_9239);
or U12234 (N_12234,N_7779,N_7816);
nand U12235 (N_12235,N_7533,N_8996);
nand U12236 (N_12236,N_7756,N_7899);
and U12237 (N_12237,N_8640,N_8477);
nor U12238 (N_12238,N_9918,N_8225);
or U12239 (N_12239,N_9200,N_7638);
and U12240 (N_12240,N_9842,N_9263);
xor U12241 (N_12241,N_7523,N_9629);
and U12242 (N_12242,N_8070,N_9462);
xor U12243 (N_12243,N_8532,N_7503);
and U12244 (N_12244,N_9236,N_8001);
nand U12245 (N_12245,N_9501,N_8417);
nor U12246 (N_12246,N_8507,N_8915);
and U12247 (N_12247,N_9236,N_8779);
xor U12248 (N_12248,N_9496,N_9304);
nand U12249 (N_12249,N_8843,N_9254);
nor U12250 (N_12250,N_8880,N_8380);
or U12251 (N_12251,N_9190,N_8983);
nand U12252 (N_12252,N_9673,N_9188);
or U12253 (N_12253,N_8313,N_8937);
xor U12254 (N_12254,N_9301,N_9497);
and U12255 (N_12255,N_7760,N_7797);
nand U12256 (N_12256,N_9886,N_8117);
nand U12257 (N_12257,N_7908,N_9994);
or U12258 (N_12258,N_9898,N_8256);
and U12259 (N_12259,N_8157,N_9639);
nand U12260 (N_12260,N_9915,N_7899);
or U12261 (N_12261,N_9021,N_7672);
and U12262 (N_12262,N_8839,N_8152);
xor U12263 (N_12263,N_8946,N_8229);
or U12264 (N_12264,N_9145,N_7960);
nor U12265 (N_12265,N_9762,N_8714);
xnor U12266 (N_12266,N_8767,N_7737);
xnor U12267 (N_12267,N_9681,N_7849);
xnor U12268 (N_12268,N_8819,N_8168);
nor U12269 (N_12269,N_7841,N_8937);
nand U12270 (N_12270,N_9095,N_8104);
nand U12271 (N_12271,N_8924,N_7833);
xnor U12272 (N_12272,N_8865,N_9314);
or U12273 (N_12273,N_8963,N_8461);
xor U12274 (N_12274,N_7773,N_8321);
or U12275 (N_12275,N_8157,N_8814);
xor U12276 (N_12276,N_7966,N_9726);
and U12277 (N_12277,N_8424,N_8344);
and U12278 (N_12278,N_7639,N_8725);
nor U12279 (N_12279,N_7633,N_7704);
nor U12280 (N_12280,N_7593,N_8746);
nor U12281 (N_12281,N_9493,N_8236);
or U12282 (N_12282,N_9279,N_8919);
nor U12283 (N_12283,N_9439,N_8275);
or U12284 (N_12284,N_9138,N_8585);
nor U12285 (N_12285,N_9353,N_8017);
and U12286 (N_12286,N_9171,N_9998);
nor U12287 (N_12287,N_7688,N_9047);
xnor U12288 (N_12288,N_7845,N_7611);
xor U12289 (N_12289,N_7738,N_9172);
nor U12290 (N_12290,N_9500,N_8242);
and U12291 (N_12291,N_9799,N_8226);
nor U12292 (N_12292,N_9339,N_9819);
nand U12293 (N_12293,N_7938,N_8619);
xor U12294 (N_12294,N_9316,N_8708);
and U12295 (N_12295,N_8365,N_8030);
xor U12296 (N_12296,N_8158,N_9748);
nor U12297 (N_12297,N_9554,N_9255);
or U12298 (N_12298,N_9415,N_7625);
and U12299 (N_12299,N_8379,N_8953);
nor U12300 (N_12300,N_8952,N_8607);
and U12301 (N_12301,N_8858,N_8140);
nand U12302 (N_12302,N_9718,N_8827);
and U12303 (N_12303,N_8637,N_8931);
xor U12304 (N_12304,N_9303,N_9697);
or U12305 (N_12305,N_9773,N_8962);
xnor U12306 (N_12306,N_8652,N_8315);
or U12307 (N_12307,N_9708,N_9634);
or U12308 (N_12308,N_7628,N_8893);
or U12309 (N_12309,N_9369,N_9531);
nor U12310 (N_12310,N_7702,N_9714);
or U12311 (N_12311,N_7949,N_9610);
or U12312 (N_12312,N_8660,N_7845);
and U12313 (N_12313,N_8198,N_8244);
xnor U12314 (N_12314,N_8424,N_9964);
xnor U12315 (N_12315,N_8959,N_7577);
nor U12316 (N_12316,N_9468,N_9510);
or U12317 (N_12317,N_9298,N_7865);
xnor U12318 (N_12318,N_9671,N_9720);
nand U12319 (N_12319,N_7586,N_7570);
xnor U12320 (N_12320,N_9934,N_8836);
xor U12321 (N_12321,N_7569,N_7829);
and U12322 (N_12322,N_7879,N_7546);
nand U12323 (N_12323,N_8298,N_8156);
nor U12324 (N_12324,N_8861,N_8420);
and U12325 (N_12325,N_8070,N_9485);
or U12326 (N_12326,N_9686,N_9299);
and U12327 (N_12327,N_9910,N_7720);
and U12328 (N_12328,N_9820,N_7745);
xor U12329 (N_12329,N_7714,N_8777);
xnor U12330 (N_12330,N_8114,N_8622);
nand U12331 (N_12331,N_8359,N_8304);
or U12332 (N_12332,N_9386,N_9979);
or U12333 (N_12333,N_9535,N_9657);
nand U12334 (N_12334,N_8302,N_7762);
nand U12335 (N_12335,N_9243,N_9386);
xor U12336 (N_12336,N_9018,N_7622);
xnor U12337 (N_12337,N_7703,N_8910);
and U12338 (N_12338,N_8565,N_7978);
xor U12339 (N_12339,N_9598,N_7939);
nand U12340 (N_12340,N_7880,N_8312);
and U12341 (N_12341,N_7784,N_9842);
and U12342 (N_12342,N_9746,N_9944);
and U12343 (N_12343,N_7777,N_9812);
xor U12344 (N_12344,N_8075,N_9731);
or U12345 (N_12345,N_7912,N_8717);
and U12346 (N_12346,N_8830,N_9182);
nand U12347 (N_12347,N_8193,N_7656);
nand U12348 (N_12348,N_9539,N_8799);
nor U12349 (N_12349,N_8290,N_8695);
xor U12350 (N_12350,N_8671,N_8648);
or U12351 (N_12351,N_7870,N_9827);
nand U12352 (N_12352,N_8504,N_9030);
nor U12353 (N_12353,N_8604,N_7952);
xor U12354 (N_12354,N_9615,N_8937);
nand U12355 (N_12355,N_8239,N_7620);
nand U12356 (N_12356,N_9400,N_7599);
and U12357 (N_12357,N_7567,N_9323);
nand U12358 (N_12358,N_8430,N_9709);
xnor U12359 (N_12359,N_8962,N_9590);
and U12360 (N_12360,N_9415,N_9057);
and U12361 (N_12361,N_9427,N_9076);
nand U12362 (N_12362,N_8194,N_9634);
nand U12363 (N_12363,N_9132,N_8631);
or U12364 (N_12364,N_7511,N_8765);
nand U12365 (N_12365,N_9687,N_8920);
nand U12366 (N_12366,N_9245,N_8008);
or U12367 (N_12367,N_9876,N_8712);
nand U12368 (N_12368,N_8136,N_8285);
xor U12369 (N_12369,N_7902,N_7592);
or U12370 (N_12370,N_9828,N_9830);
nor U12371 (N_12371,N_7904,N_8522);
xnor U12372 (N_12372,N_8420,N_9949);
nor U12373 (N_12373,N_7586,N_8522);
or U12374 (N_12374,N_8007,N_9668);
or U12375 (N_12375,N_7843,N_8718);
xor U12376 (N_12376,N_8602,N_9991);
or U12377 (N_12377,N_8245,N_7935);
xnor U12378 (N_12378,N_9640,N_9716);
xor U12379 (N_12379,N_8069,N_9035);
nor U12380 (N_12380,N_7883,N_8912);
nand U12381 (N_12381,N_9858,N_7554);
nor U12382 (N_12382,N_7537,N_7786);
nor U12383 (N_12383,N_8543,N_8370);
and U12384 (N_12384,N_8480,N_7543);
or U12385 (N_12385,N_8763,N_7659);
nand U12386 (N_12386,N_8253,N_8739);
or U12387 (N_12387,N_9726,N_7596);
or U12388 (N_12388,N_9581,N_9313);
nor U12389 (N_12389,N_7858,N_8518);
and U12390 (N_12390,N_8857,N_8183);
nor U12391 (N_12391,N_9632,N_7587);
or U12392 (N_12392,N_8557,N_8958);
or U12393 (N_12393,N_8858,N_8653);
xnor U12394 (N_12394,N_9358,N_8731);
nand U12395 (N_12395,N_8072,N_7581);
nor U12396 (N_12396,N_7729,N_9166);
or U12397 (N_12397,N_8679,N_8540);
and U12398 (N_12398,N_9859,N_9269);
nand U12399 (N_12399,N_9489,N_9378);
nand U12400 (N_12400,N_9086,N_8290);
and U12401 (N_12401,N_9488,N_8977);
and U12402 (N_12402,N_9344,N_8466);
nand U12403 (N_12403,N_9689,N_9574);
nand U12404 (N_12404,N_8759,N_9429);
nor U12405 (N_12405,N_7981,N_8972);
and U12406 (N_12406,N_8203,N_9335);
xnor U12407 (N_12407,N_8728,N_7813);
nand U12408 (N_12408,N_8921,N_8487);
or U12409 (N_12409,N_8924,N_7810);
xor U12410 (N_12410,N_9506,N_7559);
or U12411 (N_12411,N_9961,N_7987);
or U12412 (N_12412,N_9604,N_9847);
xor U12413 (N_12413,N_9573,N_8990);
and U12414 (N_12414,N_9613,N_8579);
xor U12415 (N_12415,N_7806,N_8025);
or U12416 (N_12416,N_8552,N_9511);
xor U12417 (N_12417,N_9129,N_9328);
and U12418 (N_12418,N_9419,N_8532);
and U12419 (N_12419,N_9259,N_9308);
nor U12420 (N_12420,N_8175,N_9733);
and U12421 (N_12421,N_9492,N_7855);
or U12422 (N_12422,N_8146,N_8777);
nand U12423 (N_12423,N_9669,N_8132);
nor U12424 (N_12424,N_8359,N_7771);
xnor U12425 (N_12425,N_8765,N_8406);
nand U12426 (N_12426,N_8586,N_8643);
and U12427 (N_12427,N_9684,N_7889);
nand U12428 (N_12428,N_9122,N_7721);
or U12429 (N_12429,N_9836,N_8404);
and U12430 (N_12430,N_7916,N_7753);
and U12431 (N_12431,N_9966,N_7683);
and U12432 (N_12432,N_8022,N_9446);
nor U12433 (N_12433,N_9001,N_8714);
xnor U12434 (N_12434,N_9170,N_9997);
or U12435 (N_12435,N_8444,N_9473);
or U12436 (N_12436,N_8167,N_9305);
xor U12437 (N_12437,N_8360,N_8261);
and U12438 (N_12438,N_9944,N_8728);
nor U12439 (N_12439,N_7997,N_9907);
nor U12440 (N_12440,N_9306,N_7806);
xnor U12441 (N_12441,N_8241,N_8539);
nor U12442 (N_12442,N_9176,N_9852);
xnor U12443 (N_12443,N_9879,N_7839);
and U12444 (N_12444,N_8271,N_9109);
and U12445 (N_12445,N_8045,N_9231);
and U12446 (N_12446,N_8340,N_9913);
or U12447 (N_12447,N_8058,N_8305);
or U12448 (N_12448,N_9455,N_8065);
and U12449 (N_12449,N_7673,N_9834);
nand U12450 (N_12450,N_8348,N_7743);
nand U12451 (N_12451,N_8867,N_8476);
nor U12452 (N_12452,N_8086,N_9747);
and U12453 (N_12453,N_9488,N_9450);
and U12454 (N_12454,N_8044,N_8019);
and U12455 (N_12455,N_9049,N_9622);
nor U12456 (N_12456,N_7711,N_8168);
nor U12457 (N_12457,N_8567,N_8791);
nand U12458 (N_12458,N_7736,N_8042);
xor U12459 (N_12459,N_8429,N_9656);
nor U12460 (N_12460,N_9139,N_8838);
and U12461 (N_12461,N_7728,N_8361);
nor U12462 (N_12462,N_8139,N_7569);
nor U12463 (N_12463,N_8212,N_9453);
nand U12464 (N_12464,N_9586,N_9739);
xnor U12465 (N_12465,N_9558,N_9295);
or U12466 (N_12466,N_9730,N_9560);
nand U12467 (N_12467,N_9205,N_8820);
xnor U12468 (N_12468,N_8187,N_8697);
nor U12469 (N_12469,N_7617,N_8456);
nor U12470 (N_12470,N_9756,N_9057);
xnor U12471 (N_12471,N_8216,N_9424);
nor U12472 (N_12472,N_9963,N_9995);
nand U12473 (N_12473,N_9212,N_7532);
and U12474 (N_12474,N_8037,N_9375);
xor U12475 (N_12475,N_8271,N_8726);
xor U12476 (N_12476,N_8547,N_7731);
or U12477 (N_12477,N_8525,N_9919);
nand U12478 (N_12478,N_8652,N_8995);
or U12479 (N_12479,N_7523,N_7722);
nand U12480 (N_12480,N_9374,N_8870);
or U12481 (N_12481,N_9829,N_9024);
or U12482 (N_12482,N_8213,N_7539);
xnor U12483 (N_12483,N_8264,N_8058);
or U12484 (N_12484,N_8619,N_8888);
nand U12485 (N_12485,N_9456,N_9179);
nor U12486 (N_12486,N_9392,N_8752);
xnor U12487 (N_12487,N_8911,N_9873);
nand U12488 (N_12488,N_8760,N_7810);
nor U12489 (N_12489,N_8669,N_7744);
nor U12490 (N_12490,N_9419,N_7554);
nor U12491 (N_12491,N_9488,N_7773);
nand U12492 (N_12492,N_9677,N_8563);
or U12493 (N_12493,N_7579,N_7966);
and U12494 (N_12494,N_8192,N_8515);
nand U12495 (N_12495,N_8192,N_9803);
or U12496 (N_12496,N_7799,N_8729);
nor U12497 (N_12497,N_8248,N_9633);
nand U12498 (N_12498,N_9086,N_8262);
or U12499 (N_12499,N_9179,N_9846);
and U12500 (N_12500,N_10445,N_11388);
or U12501 (N_12501,N_11768,N_11377);
xor U12502 (N_12502,N_11033,N_11571);
nand U12503 (N_12503,N_11090,N_10761);
and U12504 (N_12504,N_11469,N_11390);
nor U12505 (N_12505,N_10493,N_11427);
nor U12506 (N_12506,N_10471,N_12075);
xor U12507 (N_12507,N_12316,N_11275);
nor U12508 (N_12508,N_10121,N_12200);
or U12509 (N_12509,N_10741,N_11185);
nand U12510 (N_12510,N_12305,N_10838);
and U12511 (N_12511,N_11245,N_12159);
nand U12512 (N_12512,N_11880,N_11343);
xor U12513 (N_12513,N_11927,N_10459);
nor U12514 (N_12514,N_12274,N_11872);
xor U12515 (N_12515,N_10823,N_10605);
and U12516 (N_12516,N_11817,N_11823);
or U12517 (N_12517,N_12044,N_12164);
and U12518 (N_12518,N_11827,N_12267);
or U12519 (N_12519,N_11970,N_10654);
or U12520 (N_12520,N_11975,N_10461);
or U12521 (N_12521,N_12109,N_11402);
and U12522 (N_12522,N_12165,N_10062);
or U12523 (N_12523,N_10875,N_11917);
nor U12524 (N_12524,N_10725,N_10154);
nor U12525 (N_12525,N_10960,N_10424);
xnor U12526 (N_12526,N_12321,N_11789);
nand U12527 (N_12527,N_11997,N_12488);
xor U12528 (N_12528,N_10120,N_12262);
xor U12529 (N_12529,N_10063,N_10084);
or U12530 (N_12530,N_11224,N_11664);
nor U12531 (N_12531,N_10742,N_11401);
or U12532 (N_12532,N_10298,N_10150);
or U12533 (N_12533,N_11287,N_10856);
and U12534 (N_12534,N_11329,N_10125);
nor U12535 (N_12535,N_11058,N_10697);
and U12536 (N_12536,N_10480,N_10879);
nand U12537 (N_12537,N_12252,N_11755);
nand U12538 (N_12538,N_10730,N_10969);
or U12539 (N_12539,N_11238,N_11841);
or U12540 (N_12540,N_12461,N_11362);
and U12541 (N_12541,N_11910,N_11727);
xor U12542 (N_12542,N_10239,N_11658);
and U12543 (N_12543,N_10865,N_10132);
xor U12544 (N_12544,N_11251,N_10234);
or U12545 (N_12545,N_10232,N_10346);
nor U12546 (N_12546,N_11921,N_11060);
or U12547 (N_12547,N_10801,N_11095);
and U12548 (N_12548,N_10876,N_10408);
or U12549 (N_12549,N_11115,N_10770);
nand U12550 (N_12550,N_11996,N_10517);
and U12551 (N_12551,N_11121,N_12242);
and U12552 (N_12552,N_12275,N_12160);
and U12553 (N_12553,N_11886,N_11053);
xor U12554 (N_12554,N_11017,N_11083);
xor U12555 (N_12555,N_11334,N_11369);
or U12556 (N_12556,N_11415,N_11739);
nand U12557 (N_12557,N_10197,N_10092);
xnor U12558 (N_12558,N_11254,N_10256);
xnor U12559 (N_12559,N_11803,N_10302);
and U12560 (N_12560,N_10415,N_12436);
and U12561 (N_12561,N_10972,N_10262);
and U12562 (N_12562,N_10138,N_11724);
nor U12563 (N_12563,N_12009,N_10936);
or U12564 (N_12564,N_11365,N_10732);
xor U12565 (N_12565,N_12329,N_11235);
nand U12566 (N_12566,N_10859,N_10812);
and U12567 (N_12567,N_10866,N_11567);
nor U12568 (N_12568,N_12104,N_10858);
and U12569 (N_12569,N_11828,N_11111);
or U12570 (N_12570,N_10665,N_10830);
or U12571 (N_12571,N_11820,N_11485);
nand U12572 (N_12572,N_10826,N_10588);
and U12573 (N_12573,N_12096,N_10520);
nand U12574 (N_12574,N_11558,N_10990);
or U12575 (N_12575,N_11197,N_12272);
nor U12576 (N_12576,N_11067,N_11443);
or U12577 (N_12577,N_11852,N_11107);
xor U12578 (N_12578,N_10645,N_10082);
and U12579 (N_12579,N_12062,N_12086);
nand U12580 (N_12580,N_12048,N_10474);
xor U12581 (N_12581,N_11175,N_10388);
nor U12582 (N_12582,N_12209,N_10845);
and U12583 (N_12583,N_10612,N_11373);
nand U12584 (N_12584,N_11504,N_12173);
and U12585 (N_12585,N_11529,N_10235);
nand U12586 (N_12586,N_11954,N_10624);
nor U12587 (N_12587,N_11361,N_11766);
and U12588 (N_12588,N_11486,N_12391);
nand U12589 (N_12589,N_10978,N_12015);
nor U12590 (N_12590,N_12479,N_11453);
xor U12591 (N_12591,N_11769,N_11376);
xnor U12592 (N_12592,N_10921,N_11913);
nor U12593 (N_12593,N_11720,N_10935);
or U12594 (N_12594,N_11648,N_10579);
and U12595 (N_12595,N_11289,N_10486);
nand U12596 (N_12596,N_11237,N_12154);
or U12597 (N_12597,N_12487,N_11007);
xor U12598 (N_12598,N_12248,N_12481);
nand U12599 (N_12599,N_11605,N_10464);
nand U12600 (N_12600,N_11753,N_10818);
and U12601 (N_12601,N_11864,N_11578);
nor U12602 (N_12602,N_10572,N_10407);
or U12603 (N_12603,N_10767,N_11074);
nand U12604 (N_12604,N_11920,N_10429);
nand U12605 (N_12605,N_10829,N_10175);
and U12606 (N_12606,N_11048,N_11157);
nor U12607 (N_12607,N_10567,N_11773);
nor U12608 (N_12608,N_10432,N_11673);
nand U12609 (N_12609,N_10208,N_10957);
xnor U12610 (N_12610,N_11561,N_10338);
or U12611 (N_12611,N_10729,N_11831);
xor U12612 (N_12612,N_11932,N_11772);
and U12613 (N_12613,N_11903,N_10403);
or U12614 (N_12614,N_11778,N_10778);
and U12615 (N_12615,N_10023,N_10014);
xor U12616 (N_12616,N_11211,N_12230);
nor U12617 (N_12617,N_10526,N_10776);
or U12618 (N_12618,N_10350,N_11381);
nand U12619 (N_12619,N_11548,N_11608);
or U12620 (N_12620,N_10358,N_10669);
and U12621 (N_12621,N_10602,N_11981);
and U12622 (N_12622,N_11079,N_12040);
nand U12623 (N_12623,N_10056,N_10247);
nor U12624 (N_12624,N_10723,N_10805);
nor U12625 (N_12625,N_11492,N_12189);
or U12626 (N_12626,N_11893,N_11464);
nor U12627 (N_12627,N_11968,N_11716);
nor U12628 (N_12628,N_10793,N_12187);
and U12629 (N_12629,N_12083,N_12198);
nand U12630 (N_12630,N_10995,N_11835);
nor U12631 (N_12631,N_10817,N_11278);
nor U12632 (N_12632,N_10038,N_11266);
or U12633 (N_12633,N_11596,N_11318);
nor U12634 (N_12634,N_11389,N_12442);
xnor U12635 (N_12635,N_10748,N_10989);
nand U12636 (N_12636,N_12184,N_10945);
nor U12637 (N_12637,N_10837,N_11368);
or U12638 (N_12638,N_10048,N_11692);
and U12639 (N_12639,N_11512,N_11992);
and U12640 (N_12640,N_11801,N_10484);
and U12641 (N_12641,N_12234,N_12337);
or U12642 (N_12642,N_10953,N_10584);
xnor U12643 (N_12643,N_10258,N_11171);
nand U12644 (N_12644,N_11173,N_10738);
nor U12645 (N_12645,N_10981,N_11788);
nand U12646 (N_12646,N_11544,N_12494);
nand U12647 (N_12647,N_11925,N_11679);
and U12648 (N_12648,N_10068,N_11719);
and U12649 (N_12649,N_11680,N_12012);
and U12650 (N_12650,N_10521,N_12112);
and U12651 (N_12651,N_10781,N_11256);
nor U12652 (N_12652,N_12217,N_11281);
or U12653 (N_12653,N_10218,N_11301);
or U12654 (N_12654,N_12340,N_11135);
nand U12655 (N_12655,N_11723,N_10760);
nand U12656 (N_12656,N_12417,N_10582);
nor U12657 (N_12657,N_10238,N_12101);
and U12658 (N_12658,N_11645,N_10246);
xor U12659 (N_12659,N_12170,N_10965);
xor U12660 (N_12660,N_11011,N_11885);
nand U12661 (N_12661,N_10558,N_10516);
xnor U12662 (N_12662,N_10032,N_12484);
nand U12663 (N_12663,N_10337,N_10542);
nand U12664 (N_12664,N_10207,N_11814);
xnor U12665 (N_12665,N_10914,N_12413);
or U12666 (N_12666,N_10754,N_11526);
nand U12667 (N_12667,N_11955,N_11428);
and U12668 (N_12668,N_10257,N_10631);
nor U12669 (N_12669,N_11468,N_11677);
nand U12670 (N_12670,N_11220,N_12277);
and U12671 (N_12671,N_11259,N_11756);
or U12672 (N_12672,N_11454,N_11620);
nand U12673 (N_12673,N_10877,N_11812);
nor U12674 (N_12674,N_11505,N_10019);
xor U12675 (N_12675,N_11424,N_12357);
and U12676 (N_12676,N_10359,N_10052);
or U12677 (N_12677,N_10682,N_11093);
xnor U12678 (N_12678,N_12310,N_10438);
nand U12679 (N_12679,N_10946,N_11952);
and U12680 (N_12680,N_11805,N_11019);
nor U12681 (N_12681,N_11702,N_11530);
nand U12682 (N_12682,N_11044,N_12422);
and U12683 (N_12683,N_11179,N_11649);
and U12684 (N_12684,N_10304,N_11637);
and U12685 (N_12685,N_10353,N_10451);
and U12686 (N_12686,N_12314,N_10269);
nor U12687 (N_12687,N_10312,N_11566);
nor U12688 (N_12688,N_12288,N_12476);
nor U12689 (N_12689,N_12285,N_11031);
or U12690 (N_12690,N_10880,N_11589);
nand U12691 (N_12691,N_10080,N_10940);
nor U12692 (N_12692,N_11158,N_10755);
nand U12693 (N_12693,N_10814,N_10692);
nor U12694 (N_12694,N_12077,N_10255);
nand U12695 (N_12695,N_12051,N_12460);
xor U12696 (N_12696,N_11335,N_12379);
xor U12697 (N_12697,N_10721,N_11502);
and U12698 (N_12698,N_11517,N_11707);
nand U12699 (N_12699,N_11073,N_12356);
nand U12700 (N_12700,N_11172,N_12374);
or U12701 (N_12701,N_10615,N_10959);
xnor U12702 (N_12702,N_12309,N_10402);
or U12703 (N_12703,N_12097,N_10890);
nand U12704 (N_12704,N_10827,N_10580);
nor U12705 (N_12705,N_12468,N_11891);
xnor U12706 (N_12706,N_10882,N_12418);
xor U12707 (N_12707,N_11697,N_10263);
or U12708 (N_12708,N_10621,N_10822);
nand U12709 (N_12709,N_11795,N_10625);
and U12710 (N_12710,N_12081,N_12496);
nor U12711 (N_12711,N_10901,N_12495);
or U12712 (N_12712,N_10731,N_12058);
xnor U12713 (N_12713,N_10545,N_10894);
xnor U12714 (N_12714,N_12289,N_10757);
xor U12715 (N_12715,N_11202,N_11507);
and U12716 (N_12716,N_12064,N_11915);
nor U12717 (N_12717,N_11728,N_12183);
or U12718 (N_12718,N_12393,N_10927);
and U12719 (N_12719,N_10381,N_10334);
nand U12720 (N_12720,N_11935,N_10639);
nor U12721 (N_12721,N_10112,N_11693);
nor U12722 (N_12722,N_12404,N_11822);
or U12723 (N_12723,N_11824,N_10096);
nand U12724 (N_12724,N_10999,N_10368);
and U12725 (N_12725,N_11227,N_12136);
and U12726 (N_12726,N_12485,N_11042);
and U12727 (N_12727,N_10983,N_10036);
and U12728 (N_12728,N_11993,N_12045);
nor U12729 (N_12729,N_10864,N_10297);
nor U12730 (N_12730,N_11612,N_10344);
nor U12731 (N_12731,N_11447,N_12228);
nor U12732 (N_12732,N_11091,N_10076);
or U12733 (N_12733,N_11130,N_11951);
xnor U12734 (N_12734,N_10272,N_12022);
or U12735 (N_12735,N_10434,N_10657);
or U12736 (N_12736,N_12470,N_11481);
or U12737 (N_12737,N_11884,N_11367);
nand U12738 (N_12738,N_11889,N_11116);
xnor U12739 (N_12739,N_11101,N_10210);
or U12740 (N_12740,N_10984,N_10724);
and U12741 (N_12741,N_12107,N_11705);
nand U12742 (N_12742,N_10413,N_11793);
and U12743 (N_12743,N_11636,N_11830);
or U12744 (N_12744,N_10543,N_11597);
xnor U12745 (N_12745,N_10660,N_12052);
nand U12746 (N_12746,N_11644,N_10790);
nor U12747 (N_12747,N_12042,N_11147);
or U12748 (N_12748,N_10749,N_10825);
and U12749 (N_12749,N_12158,N_10792);
or U12750 (N_12750,N_11640,N_11174);
xor U12751 (N_12751,N_11592,N_10863);
nand U12752 (N_12752,N_12156,N_11523);
xor U12753 (N_12753,N_10284,N_12126);
nor U12754 (N_12754,N_10675,N_10406);
nor U12755 (N_12755,N_10676,N_12123);
nand U12756 (N_12756,N_12298,N_11770);
and U12757 (N_12757,N_10926,N_11919);
or U12758 (N_12758,N_10212,N_10930);
nor U12759 (N_12759,N_11406,N_10454);
xor U12760 (N_12760,N_12482,N_11326);
or U12761 (N_12761,N_12445,N_10924);
xnor U12762 (N_12762,N_11767,N_11375);
nor U12763 (N_12763,N_11267,N_10204);
xor U12764 (N_12764,N_10928,N_11141);
nor U12765 (N_12765,N_10411,N_10022);
and U12766 (N_12766,N_10819,N_12144);
nor U12767 (N_12767,N_11930,N_10236);
nor U12768 (N_12768,N_11718,N_11156);
and U12769 (N_12769,N_10417,N_11014);
or U12770 (N_12770,N_11626,N_10017);
nand U12771 (N_12771,N_10569,N_12318);
or U12772 (N_12772,N_11837,N_10378);
xnor U12773 (N_12773,N_10362,N_12213);
xor U12774 (N_12774,N_12348,N_10202);
nand U12775 (N_12775,N_10385,N_10189);
xor U12776 (N_12776,N_11440,N_10994);
or U12777 (N_12777,N_10922,N_12497);
or U12778 (N_12778,N_10536,N_10668);
nand U12779 (N_12779,N_12181,N_11150);
xor U12780 (N_12780,N_10634,N_11139);
nand U12781 (N_12781,N_10007,N_11686);
nand U12782 (N_12782,N_11187,N_12021);
and U12783 (N_12783,N_12134,N_12443);
xor U12784 (N_12784,N_12023,N_11004);
nand U12785 (N_12785,N_10141,N_11344);
or U12786 (N_12786,N_10209,N_10170);
xnor U12787 (N_12787,N_10511,N_11422);
xnor U12788 (N_12788,N_11153,N_10364);
or U12789 (N_12789,N_12477,N_10640);
nand U12790 (N_12790,N_10951,N_10490);
nand U12791 (N_12791,N_11409,N_10685);
xnor U12792 (N_12792,N_10199,N_11054);
or U12793 (N_12793,N_10974,N_12459);
or U12794 (N_12794,N_10977,N_10574);
xor U12795 (N_12795,N_10098,N_12448);
and U12796 (N_12796,N_11451,N_10559);
nor U12797 (N_12797,N_11871,N_11675);
xor U12798 (N_12798,N_10093,N_11874);
xnor U12799 (N_12799,N_11937,N_11869);
nand U12800 (N_12800,N_12392,N_12210);
and U12801 (N_12801,N_12306,N_11056);
and U12802 (N_12802,N_12328,N_12095);
or U12803 (N_12803,N_12268,N_11378);
xnor U12804 (N_12804,N_10041,N_12419);
or U12805 (N_12805,N_11327,N_10505);
nand U12806 (N_12806,N_12257,N_11684);
or U12807 (N_12807,N_10943,N_12076);
xnor U12808 (N_12808,N_11312,N_11878);
nand U12809 (N_12809,N_10441,N_11050);
nand U12810 (N_12810,N_11144,N_11810);
nor U12811 (N_12811,N_10735,N_11509);
nor U12812 (N_12812,N_10457,N_11595);
xor U12813 (N_12813,N_11666,N_12090);
xor U12814 (N_12814,N_11942,N_10135);
xnor U12815 (N_12815,N_10473,N_11460);
and U12816 (N_12816,N_12472,N_10129);
nor U12817 (N_12817,N_11046,N_11650);
nand U12818 (N_12818,N_11112,N_12338);
nor U12819 (N_12819,N_10089,N_10004);
xor U12820 (N_12820,N_10514,N_12414);
nor U12821 (N_12821,N_10244,N_11222);
xor U12822 (N_12822,N_10303,N_11554);
nor U12823 (N_12823,N_10651,N_12347);
xor U12824 (N_12824,N_11717,N_10347);
or U12825 (N_12825,N_11907,N_12036);
nor U12826 (N_12826,N_10118,N_10988);
or U12827 (N_12827,N_11363,N_11759);
and U12828 (N_12828,N_12258,N_11873);
nor U12829 (N_12829,N_11687,N_10217);
nor U12830 (N_12830,N_11949,N_11228);
and U12831 (N_12831,N_10274,N_11057);
nand U12832 (N_12832,N_10696,N_11082);
nor U12833 (N_12833,N_11123,N_10172);
and U12834 (N_12834,N_10656,N_10498);
and U12835 (N_12835,N_11956,N_10734);
xnor U12836 (N_12836,N_11188,N_10870);
xnor U12837 (N_12837,N_10895,N_10775);
and U12838 (N_12838,N_11410,N_10577);
nand U12839 (N_12839,N_11108,N_12290);
nor U12840 (N_12840,N_10571,N_10492);
nand U12841 (N_12841,N_11950,N_11657);
nand U12842 (N_12842,N_12364,N_11262);
and U12843 (N_12843,N_10472,N_10240);
nand U12844 (N_12844,N_10460,N_11498);
and U12845 (N_12845,N_11600,N_10057);
or U12846 (N_12846,N_10251,N_10071);
and U12847 (N_12847,N_12440,N_11136);
and U12848 (N_12848,N_10758,N_11615);
nor U12849 (N_12849,N_12415,N_11285);
xor U12850 (N_12850,N_11096,N_11027);
nor U12851 (N_12851,N_11771,N_10252);
xnor U12852 (N_12852,N_10123,N_12471);
nand U12853 (N_12853,N_11962,N_11176);
and U12854 (N_12854,N_10648,N_11928);
nor U12855 (N_12855,N_11757,N_10485);
or U12856 (N_12856,N_10746,N_10644);
nor U12857 (N_12857,N_11560,N_11491);
and U12858 (N_12858,N_11246,N_10915);
nor U12859 (N_12859,N_10566,N_10448);
nor U12860 (N_12860,N_11219,N_11494);
nand U12861 (N_12861,N_12054,N_12118);
nor U12862 (N_12862,N_11552,N_11243);
xnor U12863 (N_12863,N_12266,N_11851);
nor U12864 (N_12864,N_11833,N_11310);
nand U12865 (N_12865,N_11021,N_11573);
or U12866 (N_12866,N_10069,N_12113);
or U12867 (N_12867,N_10557,N_11018);
nand U12868 (N_12868,N_12216,N_10736);
and U12869 (N_12869,N_10308,N_10055);
nor U12870 (N_12870,N_11883,N_11066);
nor U12871 (N_12871,N_10495,N_11964);
xnor U12872 (N_12872,N_11521,N_10905);
and U12873 (N_12873,N_10643,N_10728);
xor U12874 (N_12874,N_11352,N_11225);
or U12875 (N_12875,N_10581,N_10322);
nand U12876 (N_12876,N_11288,N_11710);
nand U12877 (N_12877,N_10664,N_10116);
and U12878 (N_12878,N_11268,N_11159);
nor U12879 (N_12879,N_10225,N_10393);
nand U12880 (N_12880,N_11355,N_11948);
nor U12881 (N_12881,N_12131,N_12026);
and U12882 (N_12882,N_11423,N_11143);
nand U12883 (N_12883,N_11371,N_11372);
nor U12884 (N_12884,N_12120,N_10534);
and U12885 (N_12885,N_10836,N_10164);
nor U12886 (N_12886,N_11223,N_11036);
or U12887 (N_12887,N_12469,N_10613);
or U12888 (N_12888,N_11669,N_10128);
or U12889 (N_12889,N_10222,N_11495);
and U12890 (N_12890,N_10952,N_10376);
nor U12891 (N_12891,N_12410,N_12002);
nor U12892 (N_12892,N_11850,N_11929);
xnor U12893 (N_12893,N_10898,N_11737);
nor U12894 (N_12894,N_10352,N_12263);
nand U12895 (N_12895,N_10227,N_10439);
xnor U12896 (N_12896,N_11966,N_10867);
or U12897 (N_12897,N_10107,N_11218);
or U12898 (N_12898,N_12241,N_10253);
nand U12899 (N_12899,N_11628,N_12435);
nor U12900 (N_12900,N_10343,N_10531);
or U12901 (N_12901,N_10803,N_11576);
and U12902 (N_12902,N_11484,N_10976);
or U12903 (N_12903,N_10478,N_10261);
and U12904 (N_12904,N_10226,N_10499);
or U12905 (N_12905,N_11979,N_10094);
and U12906 (N_12906,N_12324,N_10161);
or U12907 (N_12907,N_11213,N_11598);
xor U12908 (N_12908,N_12395,N_10481);
nand U12909 (N_12909,N_11196,N_10101);
nand U12910 (N_12910,N_11445,N_11547);
xnor U12911 (N_12911,N_11995,N_10126);
and U12912 (N_12912,N_11551,N_10515);
or U12913 (N_12913,N_10788,N_11293);
and U12914 (N_12914,N_10184,N_10689);
nand U12915 (N_12915,N_12345,N_11322);
nor U12916 (N_12916,N_10259,N_11420);
nand U12917 (N_12917,N_10155,N_11593);
nor U12918 (N_12918,N_12429,N_11939);
nor U12919 (N_12919,N_11264,N_10137);
nor U12920 (N_12920,N_11404,N_11947);
nand U12921 (N_12921,N_10070,N_10839);
nor U12922 (N_12922,N_10887,N_11591);
and U12923 (N_12923,N_12377,N_11520);
nand U12924 (N_12924,N_10287,N_10649);
and U12925 (N_12925,N_12449,N_10426);
xnor U12926 (N_12926,N_12421,N_12060);
and U12927 (N_12927,N_10519,N_10243);
nand U12928 (N_12928,N_11911,N_10693);
nand U12929 (N_12929,N_11671,N_10899);
or U12930 (N_12930,N_10750,N_12341);
nand U12931 (N_12931,N_10501,N_12203);
nor U12932 (N_12932,N_10401,N_11609);
or U12933 (N_12933,N_10370,N_10309);
xor U12934 (N_12934,N_10296,N_11711);
nor U12935 (N_12935,N_12388,N_11037);
xor U12936 (N_12936,N_12344,N_10562);
nor U12937 (N_12937,N_11006,N_11394);
and U12938 (N_12938,N_10463,N_12053);
nand U12939 (N_12939,N_11764,N_11309);
or U12940 (N_12940,N_10494,N_11639);
nand U12941 (N_12941,N_11183,N_11627);
and U12942 (N_12942,N_12411,N_10191);
or U12943 (N_12943,N_10311,N_12339);
and U12944 (N_12944,N_12190,N_10857);
nand U12945 (N_12945,N_11958,N_11514);
and U12946 (N_12946,N_10512,N_10659);
xor U12947 (N_12947,N_12416,N_12363);
nand U12948 (N_12948,N_10608,N_11570);
xnor U12949 (N_12949,N_11622,N_12066);
or U12950 (N_12950,N_11337,N_10355);
xnor U12951 (N_12951,N_10578,N_11126);
and U12952 (N_12952,N_10030,N_12355);
nand U12953 (N_12953,N_10679,N_10289);
nor U12954 (N_12954,N_10744,N_12029);
and U12955 (N_12955,N_10973,N_11162);
xor U12956 (N_12956,N_11308,N_10314);
nand U12957 (N_12957,N_11704,N_10105);
nor U12958 (N_12958,N_10743,N_11387);
nor U12959 (N_12959,N_11985,N_10326);
nand U12960 (N_12960,N_11849,N_11290);
and U12961 (N_12961,N_12312,N_12451);
nand U12962 (N_12962,N_10794,N_12224);
nand U12963 (N_12963,N_10831,N_11496);
nor U12964 (N_12964,N_10002,N_12035);
nand U12965 (N_12965,N_10453,N_10363);
nand U12966 (N_12966,N_12089,N_10281);
xnor U12967 (N_12967,N_12171,N_12437);
or U12968 (N_12968,N_12088,N_12084);
nor U12969 (N_12969,N_10599,N_10313);
and U12970 (N_12970,N_11284,N_11579);
nor U12971 (N_12971,N_11861,N_10077);
and U12972 (N_12972,N_12269,N_11733);
and U12973 (N_12973,N_11161,N_11304);
xnor U12974 (N_12974,N_10475,N_10365);
and U12975 (N_12975,N_12127,N_12427);
xnor U12976 (N_12976,N_11618,N_10249);
nor U12977 (N_12977,N_11699,N_10489);
xor U12978 (N_12978,N_11207,N_10616);
or U12979 (N_12979,N_11154,N_11081);
and U12980 (N_12980,N_10224,N_10868);
nand U12981 (N_12981,N_10151,N_11296);
xor U12982 (N_12982,N_12398,N_11667);
nor U12983 (N_12983,N_12046,N_11380);
nand U12984 (N_12984,N_10647,N_10122);
nand U12985 (N_12985,N_11043,N_11934);
and U12986 (N_12986,N_10329,N_11384);
and U12987 (N_12987,N_10186,N_11846);
and U12988 (N_12988,N_10998,N_11359);
nand U12989 (N_12989,N_12492,N_12473);
or U12990 (N_12990,N_11085,N_10479);
or U12991 (N_12991,N_12100,N_11209);
nor U12992 (N_12992,N_10563,N_10000);
or U12993 (N_12993,N_11253,N_11534);
and U12994 (N_12994,N_10372,N_10250);
and U12995 (N_12995,N_10835,N_12204);
or U12996 (N_12996,N_12163,N_10888);
nand U12997 (N_12997,N_10843,N_10188);
or U12998 (N_12998,N_10034,N_12372);
and U12999 (N_12999,N_10354,N_12030);
nand U13000 (N_13000,N_12155,N_11575);
nor U13001 (N_13001,N_10671,N_11333);
nand U13002 (N_13002,N_11655,N_11140);
or U13003 (N_13003,N_12438,N_12215);
nand U13004 (N_13004,N_11444,N_10583);
and U13005 (N_13005,N_10909,N_12353);
nand U13006 (N_13006,N_10846,N_10442);
xor U13007 (N_13007,N_11425,N_12378);
and U13008 (N_13008,N_10149,N_12141);
xnor U13009 (N_13009,N_11265,N_10144);
or U13010 (N_13010,N_11983,N_11026);
nand U13011 (N_13011,N_11506,N_12490);
xnor U13012 (N_13012,N_12354,N_10687);
xnor U13013 (N_13013,N_11938,N_11429);
and U13014 (N_13014,N_10533,N_12303);
nor U13015 (N_13015,N_12342,N_11459);
and U13016 (N_13016,N_11470,N_10131);
and U13017 (N_13017,N_10872,N_12122);
xor U13018 (N_13018,N_11480,N_12352);
nor U13019 (N_13019,N_11455,N_11539);
nor U13020 (N_13020,N_12219,N_10003);
or U13021 (N_13021,N_10081,N_10395);
nor U13022 (N_13022,N_11594,N_10143);
xor U13023 (N_13023,N_11005,N_10387);
and U13024 (N_13024,N_11839,N_10051);
or U13025 (N_13025,N_11786,N_11838);
or U13026 (N_13026,N_10342,N_10813);
xnor U13027 (N_13027,N_10653,N_10111);
or U13028 (N_13028,N_11117,N_10046);
and U13029 (N_13029,N_11064,N_12037);
nor U13030 (N_13030,N_11545,N_10054);
nand U13031 (N_13031,N_10397,N_11556);
xor U13032 (N_13032,N_10159,N_11961);
nand U13033 (N_13033,N_10919,N_11386);
nand U13034 (N_13034,N_10766,N_10280);
and U13035 (N_13035,N_11652,N_10820);
nor U13036 (N_13036,N_10650,N_10832);
nor U13037 (N_13037,N_11638,N_10769);
nand U13038 (N_13038,N_10683,N_11847);
nor U13039 (N_13039,N_12297,N_10768);
or U13040 (N_13040,N_11746,N_10854);
and U13041 (N_13041,N_12408,N_12229);
xor U13042 (N_13042,N_11109,N_12013);
xor U13043 (N_13043,N_11887,N_11549);
xnor U13044 (N_13044,N_11255,N_11128);
xnor U13045 (N_13045,N_11252,N_12236);
xnor U13046 (N_13046,N_10646,N_11477);
or U13047 (N_13047,N_10264,N_11760);
xor U13048 (N_13048,N_10042,N_10938);
and U13049 (N_13049,N_10073,N_11300);
and U13050 (N_13050,N_10153,N_10897);
xor U13051 (N_13051,N_11742,N_10294);
xnor U13052 (N_13052,N_10319,N_12177);
xnor U13053 (N_13053,N_11698,N_11167);
nand U13054 (N_13054,N_10482,N_12498);
nor U13055 (N_13055,N_10786,N_10821);
nor U13056 (N_13056,N_10954,N_12150);
xnor U13057 (N_13057,N_11194,N_11168);
and U13058 (N_13058,N_12188,N_11100);
or U13059 (N_13059,N_11518,N_10619);
or U13060 (N_13060,N_11059,N_11133);
xnor U13061 (N_13061,N_11466,N_11499);
and U13062 (N_13062,N_11681,N_10167);
or U13063 (N_13063,N_10638,N_11749);
and U13064 (N_13064,N_11821,N_11785);
nand U13065 (N_13065,N_11328,N_11353);
nor U13066 (N_13066,N_11994,N_12168);
or U13067 (N_13067,N_12380,N_12350);
or U13068 (N_13068,N_10335,N_12205);
xor U13069 (N_13069,N_10043,N_11986);
or U13070 (N_13070,N_11546,N_11663);
xnor U13071 (N_13071,N_11269,N_12382);
xnor U13072 (N_13072,N_12313,N_11317);
and U13073 (N_13073,N_11120,N_12480);
xnor U13074 (N_13074,N_11957,N_11619);
nand U13075 (N_13075,N_11988,N_11906);
and U13076 (N_13076,N_11062,N_11450);
xnor U13077 (N_13077,N_10133,N_11049);
and U13078 (N_13078,N_10248,N_10840);
nor U13079 (N_13079,N_11092,N_11918);
or U13080 (N_13080,N_10219,N_10941);
and U13081 (N_13081,N_10021,N_12027);
xor U13082 (N_13082,N_12389,N_12151);
and U13083 (N_13083,N_10487,N_11633);
nor U13084 (N_13084,N_11045,N_10714);
nand U13085 (N_13085,N_10223,N_10628);
nor U13086 (N_13086,N_10496,N_10110);
nor U13087 (N_13087,N_11973,N_12265);
or U13088 (N_13088,N_10109,N_11553);
or U13089 (N_13089,N_11706,N_10348);
nor U13090 (N_13090,N_11226,N_10944);
nand U13091 (N_13091,N_10306,N_11439);
nor U13092 (N_13092,N_11781,N_10447);
or U13093 (N_13093,N_11976,N_12117);
and U13094 (N_13094,N_12399,N_11843);
or U13095 (N_13095,N_10932,N_11114);
nor U13096 (N_13096,N_11271,N_10708);
nor U13097 (N_13097,N_11678,N_12099);
or U13098 (N_13098,N_12124,N_11408);
xor U13099 (N_13099,N_10266,N_10560);
nand U13100 (N_13100,N_11234,N_11783);
nor U13101 (N_13101,N_11063,N_11084);
nand U13102 (N_13102,N_10535,N_11260);
and U13103 (N_13103,N_12028,N_10039);
xnor U13104 (N_13104,N_11087,N_11876);
nand U13105 (N_13105,N_12323,N_10450);
and U13106 (N_13106,N_10886,N_10333);
nand U13107 (N_13107,N_10513,N_11383);
or U13108 (N_13108,N_11890,N_10849);
xor U13109 (N_13109,N_11904,N_11625);
and U13110 (N_13110,N_11432,N_12014);
xnor U13111 (N_13111,N_12192,N_11370);
nor U13112 (N_13112,N_11349,N_11974);
nor U13113 (N_13113,N_10157,N_10103);
and U13114 (N_13114,N_10980,N_11780);
and U13115 (N_13115,N_10361,N_11604);
nor U13116 (N_13116,N_10049,N_10799);
nand U13117 (N_13117,N_11905,N_10701);
or U13118 (N_13118,N_11239,N_10299);
or U13119 (N_13119,N_10815,N_11148);
nand U13120 (N_13120,N_11131,N_10398);
xnor U13121 (N_13121,N_10293,N_11532);
and U13122 (N_13122,N_11933,N_10552);
nand U13123 (N_13123,N_10510,N_10067);
nor U13124 (N_13124,N_10667,N_11944);
nand U13125 (N_13125,N_12332,N_10674);
nand U13126 (N_13126,N_11587,N_11690);
and U13127 (N_13127,N_10044,N_11010);
nor U13128 (N_13128,N_10195,N_10710);
and U13129 (N_13129,N_12145,N_11311);
nand U13130 (N_13130,N_11040,N_12238);
nand U13131 (N_13131,N_11305,N_11963);
or U13132 (N_13132,N_10436,N_11926);
nand U13133 (N_13133,N_12175,N_12319);
or U13134 (N_13134,N_10271,N_10174);
or U13135 (N_13135,N_10449,N_12447);
and U13136 (N_13136,N_11860,N_10185);
xor U13137 (N_13137,N_10525,N_10916);
nor U13138 (N_13138,N_11584,N_12361);
and U13139 (N_13139,N_10497,N_11315);
nor U13140 (N_13140,N_10469,N_10275);
or U13141 (N_13141,N_12286,N_11430);
xor U13142 (N_13142,N_11418,N_12499);
xnor U13143 (N_13143,N_11180,N_11487);
nand U13144 (N_13144,N_10198,N_12237);
or U13145 (N_13145,N_11842,N_10179);
xnor U13146 (N_13146,N_12135,N_12366);
nand U13147 (N_13147,N_12467,N_11241);
and U13148 (N_13148,N_10214,N_10420);
nor U13149 (N_13149,N_10688,N_12057);
xor U13150 (N_13150,N_10787,N_10627);
xor U13151 (N_13151,N_10145,N_12311);
xnor U13152 (N_13152,N_10862,N_12105);
or U13153 (N_13153,N_11972,N_10351);
and U13154 (N_13154,N_10611,N_11998);
or U13155 (N_13155,N_10705,N_10410);
nand U13156 (N_13156,N_11866,N_11632);
nor U13157 (N_13157,N_10291,N_11683);
and U13158 (N_13158,N_12271,N_10117);
nor U13159 (N_13159,N_10074,N_11826);
xor U13160 (N_13160,N_10414,N_10869);
nor U13161 (N_13161,N_11052,N_12326);
or U13162 (N_13162,N_10088,N_12128);
nor U13163 (N_13163,N_10673,N_11190);
nor U13164 (N_13164,N_10707,N_12454);
nor U13165 (N_13165,N_12033,N_11233);
nor U13166 (N_13166,N_11844,N_12452);
nor U13167 (N_13167,N_10553,N_10975);
nor U13168 (N_13168,N_10747,N_11965);
or U13169 (N_13169,N_10912,N_10585);
nor U13170 (N_13170,N_12172,N_12441);
or U13171 (N_13171,N_12043,N_11574);
nand U13172 (N_13172,N_11069,N_11892);
xor U13173 (N_13173,N_11366,N_11075);
xnor U13174 (N_13174,N_10216,N_10678);
xnor U13175 (N_13175,N_11647,N_10229);
and U13176 (N_13176,N_10896,N_11263);
xnor U13177 (N_13177,N_11303,N_11169);
and U13178 (N_13178,N_11248,N_12358);
xor U13179 (N_13179,N_11467,N_10282);
nor U13180 (N_13180,N_11900,N_10795);
nor U13181 (N_13181,N_12384,N_10677);
nor U13182 (N_13182,N_10102,N_10307);
xnor U13183 (N_13183,N_11338,N_12000);
nand U13184 (N_13184,N_10134,N_10881);
xor U13185 (N_13185,N_11845,N_12244);
nor U13186 (N_13186,N_12301,N_12068);
nand U13187 (N_13187,N_11089,N_11611);
and U13188 (N_13188,N_11129,N_11741);
nor U13189 (N_13189,N_10833,N_11137);
or U13190 (N_13190,N_10330,N_12179);
nor U13191 (N_13191,N_10010,N_11465);
or U13192 (N_13192,N_10375,N_10399);
or U13193 (N_13193,N_10254,N_11483);
nor U13194 (N_13194,N_11452,N_10716);
nand U13195 (N_13195,N_10610,N_12208);
or U13196 (N_13196,N_11896,N_10136);
and U13197 (N_13197,N_10331,N_12455);
nor U13198 (N_13198,N_12330,N_12003);
nor U13199 (N_13199,N_10283,N_11980);
nand U13200 (N_13200,N_10058,N_10524);
or U13201 (N_13201,N_12008,N_10712);
nor U13202 (N_13202,N_11524,N_12249);
xnor U13203 (N_13203,N_10083,N_10663);
or U13204 (N_13204,N_12456,N_11646);
and U13205 (N_13205,N_10292,N_10962);
xnor U13206 (N_13206,N_12260,N_10182);
and U13207 (N_13207,N_12385,N_11559);
xor U13208 (N_13208,N_12308,N_10300);
or U13209 (N_13209,N_11426,N_11865);
xor U13210 (N_13210,N_11336,N_12094);
nor U13211 (N_13211,N_11399,N_10146);
xnor U13212 (N_13212,N_10598,N_11221);
or U13213 (N_13213,N_11134,N_10035);
nor U13214 (N_13214,N_11061,N_10609);
or U13215 (N_13215,N_11000,N_10437);
xor U13216 (N_13216,N_12376,N_10176);
nand U13217 (N_13217,N_12394,N_11581);
nand U13218 (N_13218,N_11003,N_10108);
xor U13219 (N_13219,N_12034,N_10320);
nand U13220 (N_13220,N_11212,N_10383);
nor U13221 (N_13221,N_11316,N_12019);
or U13222 (N_13222,N_10078,N_11198);
nand U13223 (N_13223,N_10409,N_10933);
and U13224 (N_13224,N_12180,N_10324);
or U13225 (N_13225,N_12239,N_12475);
nor U13226 (N_13226,N_12450,N_11071);
nand U13227 (N_13227,N_11734,N_11434);
nor U13228 (N_13228,N_11754,N_11181);
nor U13229 (N_13229,N_11743,N_12111);
xnor U13230 (N_13230,N_11736,N_10703);
and U13231 (N_13231,N_11398,N_10316);
and U13232 (N_13232,N_12140,N_12439);
nor U13233 (N_13233,N_11393,N_12193);
xor U13234 (N_13234,N_10059,N_11784);
or U13235 (N_13235,N_11519,N_11358);
and U13236 (N_13236,N_10416,N_10504);
nand U13237 (N_13237,N_11946,N_11694);
nand U13238 (N_13238,N_11051,N_11662);
xnor U13239 (N_13239,N_10241,N_10800);
or U13240 (N_13240,N_10745,N_11214);
or U13241 (N_13241,N_11184,N_10907);
and U13242 (N_13242,N_12231,N_10221);
nor U13243 (N_13243,N_12334,N_12047);
nor U13244 (N_13244,N_10389,N_11672);
and U13245 (N_13245,N_10446,N_10662);
or U13246 (N_13246,N_10091,N_11321);
and U13247 (N_13247,N_11836,N_11295);
xor U13248 (N_13248,N_12069,N_12011);
or U13249 (N_13249,N_10382,N_10027);
xor U13250 (N_13250,N_12423,N_10380);
nand U13251 (N_13251,N_10033,N_10099);
nand U13252 (N_13252,N_12195,N_10458);
and U13253 (N_13253,N_11621,N_12250);
nand U13254 (N_13254,N_10986,N_11623);
nand U13255 (N_13255,N_10851,N_11206);
xor U13256 (N_13256,N_10165,N_10001);
nor U13257 (N_13257,N_11522,N_11099);
and U13258 (N_13258,N_12091,N_12300);
nor U13259 (N_13259,N_11691,N_10806);
nor U13260 (N_13260,N_11001,N_10925);
or U13261 (N_13261,N_11654,N_12261);
and U13262 (N_13262,N_11607,N_12152);
nor U13263 (N_13263,N_11721,N_12001);
nor U13264 (N_13264,N_11726,N_12270);
xnor U13265 (N_13265,N_10939,N_10015);
or U13266 (N_13266,N_10844,N_11065);
nor U13267 (N_13267,N_10502,N_10593);
and U13268 (N_13268,N_10357,N_12080);
xnor U13269 (N_13269,N_10231,N_11853);
nand U13270 (N_13270,N_10885,N_10477);
nand U13271 (N_13271,N_10547,N_12343);
or U13272 (N_13272,N_10491,N_12491);
and U13273 (N_13273,N_10009,N_12206);
and U13274 (N_13274,N_11745,N_11257);
xor U13275 (N_13275,N_10016,N_12369);
nor U13276 (N_13276,N_11002,N_10160);
and U13277 (N_13277,N_11160,N_11411);
or U13278 (N_13278,N_12295,N_12196);
xnor U13279 (N_13279,N_10722,N_10148);
nand U13280 (N_13280,N_12359,N_10902);
xor U13281 (N_13281,N_11472,N_10908);
nand U13282 (N_13282,N_12194,N_10968);
and U13283 (N_13283,N_11442,N_10127);
xnor U13284 (N_13284,N_11035,N_10452);
and U13285 (N_13285,N_12004,N_11894);
xnor U13286 (N_13286,N_11989,N_11557);
and U13287 (N_13287,N_11340,N_10332);
nor U13288 (N_13288,N_11030,N_11806);
xnor U13289 (N_13289,N_11500,N_10554);
or U13290 (N_13290,N_10443,N_10192);
and U13291 (N_13291,N_11382,N_10162);
or U13292 (N_13292,N_10130,N_11901);
xnor U13293 (N_13293,N_10780,N_10427);
xor U13294 (N_13294,N_10455,N_10205);
and U13295 (N_13295,N_10503,N_11634);
nand U13296 (N_13296,N_11725,N_11086);
or U13297 (N_13297,N_10233,N_11945);
nand U13298 (N_13298,N_11354,N_10367);
and U13299 (N_13299,N_10626,N_10711);
or U13300 (N_13300,N_10097,N_11614);
xor U13301 (N_13301,N_10672,N_11282);
or U13302 (N_13302,N_11888,N_12218);
xor U13303 (N_13303,N_11178,N_10718);
or U13304 (N_13304,N_11244,N_11856);
and U13305 (N_13305,N_11348,N_11195);
or U13306 (N_13306,N_11840,N_11038);
nor U13307 (N_13307,N_10878,N_10947);
nor U13308 (N_13308,N_12259,N_10412);
or U13309 (N_13309,N_11967,N_10462);
nor U13310 (N_13310,N_11164,N_10923);
xnor U13311 (N_13311,N_11564,N_10702);
or U13312 (N_13312,N_10470,N_10603);
nor U13313 (N_13313,N_11543,N_10465);
or U13314 (N_13314,N_11668,N_11897);
nor U13315 (N_13315,N_10323,N_11792);
or U13316 (N_13316,N_10530,N_12169);
xor U13317 (N_13317,N_11583,N_11777);
nor U13318 (N_13318,N_10288,N_11635);
or U13319 (N_13319,N_11577,N_10740);
nor U13320 (N_13320,N_12349,N_10321);
or U13321 (N_13321,N_12478,N_12191);
nand U13322 (N_13322,N_11098,N_10642);
nor U13323 (N_13323,N_12233,N_11490);
or U13324 (N_13324,N_10119,N_10483);
and U13325 (N_13325,N_10891,N_10931);
xor U13326 (N_13326,N_10220,N_10327);
nor U13327 (N_13327,N_10377,N_10751);
or U13328 (N_13328,N_11448,N_11441);
and U13329 (N_13329,N_10173,N_12412);
or U13330 (N_13330,N_12119,N_10699);
or U13331 (N_13331,N_11582,N_11601);
xor U13332 (N_13332,N_10555,N_11696);
and U13333 (N_13333,N_11232,N_10556);
nand U13334 (N_13334,N_12106,N_10549);
nor U13335 (N_13335,N_10428,N_12292);
nand U13336 (N_13336,N_11022,N_11802);
and U13337 (N_13337,N_12071,N_10607);
and U13338 (N_13338,N_11127,N_10177);
xnor U13339 (N_13339,N_12381,N_10911);
and U13340 (N_13340,N_11682,N_12050);
xnor U13341 (N_13341,N_10095,N_12016);
and U13342 (N_13342,N_10087,N_10374);
xnor U13343 (N_13343,N_11403,N_11013);
nand U13344 (N_13344,N_11525,N_10031);
nor U13345 (N_13345,N_12153,N_12222);
xor U13346 (N_13346,N_10573,N_11987);
xor U13347 (N_13347,N_10168,N_12464);
nand U13348 (N_13348,N_11708,N_11565);
nand U13349 (N_13349,N_11438,N_10211);
and U13350 (N_13350,N_12299,N_11476);
and U13351 (N_13351,N_11146,N_10213);
nor U13352 (N_13352,N_11216,N_10785);
xor U13353 (N_13353,N_12281,N_10500);
nand U13354 (N_13354,N_10295,N_10325);
or U13355 (N_13355,N_10772,N_11346);
and U13356 (N_13356,N_11829,N_12161);
xor U13357 (N_13357,N_11877,N_11540);
or U13358 (N_13358,N_11775,N_12197);
and U13359 (N_13359,N_10587,N_11809);
or U13360 (N_13360,N_10804,N_12103);
and U13361 (N_13361,N_12397,N_11984);
nor U13362 (N_13362,N_10537,N_11068);
xor U13363 (N_13363,N_10630,N_10190);
or U13364 (N_13364,N_10789,N_12273);
nor U13365 (N_13365,N_10025,N_11533);
nor U13366 (N_13366,N_11110,N_11854);
nor U13367 (N_13367,N_12256,N_10733);
or U13368 (N_13368,N_11493,N_11811);
xnor U13369 (N_13369,N_10345,N_10419);
nand U13370 (N_13370,N_11715,N_11642);
nor U13371 (N_13371,N_11508,N_11170);
or U13372 (N_13372,N_12444,N_10047);
and U13373 (N_13373,N_11461,N_10617);
or U13374 (N_13374,N_10910,N_11105);
or U13375 (N_13375,N_11924,N_11125);
and U13376 (N_13376,N_10169,N_10305);
nor U13377 (N_13377,N_11463,N_11325);
and U13378 (N_13378,N_10903,N_12129);
nor U13379 (N_13379,N_12024,N_10544);
or U13380 (N_13380,N_11025,N_11732);
or U13381 (N_13381,N_11794,N_12178);
nor U13382 (N_13382,N_12253,N_12433);
xnor U13383 (N_13383,N_12463,N_10764);
xor U13384 (N_13384,N_12007,N_10842);
nand U13385 (N_13385,N_10379,N_11870);
nand U13386 (N_13386,N_10230,N_10356);
nor U13387 (N_13387,N_10855,N_11419);
nand U13388 (N_13388,N_11651,N_11400);
and U13389 (N_13389,N_11094,N_11242);
nand U13390 (N_13390,N_11351,N_10053);
nand U13391 (N_13391,N_11102,N_10641);
nand U13392 (N_13392,N_10421,N_11735);
nor U13393 (N_13393,N_10680,N_10286);
nor U13394 (N_13394,N_12223,N_11535);
nand U13395 (N_13395,N_10848,N_11306);
or U13396 (N_13396,N_11240,N_12287);
or U13397 (N_13397,N_11436,N_10201);
nand U13398 (N_13398,N_11433,N_11779);
and U13399 (N_13399,N_11555,N_11217);
and U13400 (N_13400,N_10425,N_10592);
xor U13401 (N_13401,N_10798,N_12199);
xnor U13402 (N_13402,N_10158,N_11804);
nor U13403 (N_13403,N_12202,N_12402);
and U13404 (N_13404,N_10779,N_11166);
and U13405 (N_13405,N_11709,N_10684);
xnor U13406 (N_13406,N_11177,N_10691);
nor U13407 (N_13407,N_10904,N_12211);
xor U13408 (N_13408,N_10620,N_12351);
xor U13409 (N_13409,N_10955,N_11313);
or U13410 (N_13410,N_11511,N_11714);
xnor U13411 (N_13411,N_11291,N_11613);
and U13412 (N_13412,N_12400,N_11270);
or U13413 (N_13413,N_10797,N_12226);
or U13414 (N_13414,N_10340,N_11200);
nand U13415 (N_13415,N_11392,N_12428);
nor U13416 (N_13416,N_11482,N_11072);
nand U13417 (N_13417,N_10590,N_11319);
xor U13418 (N_13418,N_11782,N_11279);
nor U13419 (N_13419,N_11501,N_11342);
or U13420 (N_13420,N_10632,N_11473);
or U13421 (N_13421,N_10704,N_10508);
or U13422 (N_13422,N_11943,N_11431);
nand U13423 (N_13423,N_11374,N_12182);
nor U13424 (N_13424,N_10948,N_11902);
nand U13425 (N_13425,N_12296,N_11816);
xor U13426 (N_13426,N_12092,N_11859);
or U13427 (N_13427,N_11145,N_11456);
nor U13428 (N_13428,N_11163,N_11249);
nor U13429 (N_13429,N_11538,N_10006);
nand U13430 (N_13430,N_11489,N_11435);
or U13431 (N_13431,N_11231,N_12403);
nor U13432 (N_13432,N_10509,N_11497);
nand U13433 (N_13433,N_11462,N_12307);
and U13434 (N_13434,N_10171,N_12132);
or U13435 (N_13435,N_10737,N_11563);
xor U13436 (N_13436,N_10104,N_10686);
nor U13437 (N_13437,N_11763,N_11024);
xnor U13438 (N_13438,N_10618,N_12018);
and U13439 (N_13439,N_11800,N_11879);
or U13440 (N_13440,N_11201,N_12406);
nor U13441 (N_13441,N_12149,N_12162);
xnor U13442 (N_13442,N_12079,N_11624);
and U13443 (N_13443,N_10404,N_12294);
nor U13444 (N_13444,N_12458,N_11314);
nor U13445 (N_13445,N_11106,N_11510);
nand U13446 (N_13446,N_12055,N_11590);
nand U13447 (N_13447,N_11297,N_10791);
nor U13448 (N_13448,N_11009,N_11999);
nor U13449 (N_13449,N_12387,N_11039);
or U13450 (N_13450,N_11118,N_12240);
xnor U13451 (N_13451,N_11449,N_11774);
xnor U13452 (N_13452,N_11787,N_12282);
and U13453 (N_13453,N_10028,N_10152);
and U13454 (N_13454,N_10802,N_11323);
xor U13455 (N_13455,N_11229,N_10290);
and U13456 (N_13456,N_10518,N_11397);
xor U13457 (N_13457,N_10339,N_10753);
or U13458 (N_13458,N_12371,N_10423);
or U13459 (N_13459,N_10277,N_12434);
or U13460 (N_13460,N_11819,N_10276);
and U13461 (N_13461,N_11215,N_10606);
and U13462 (N_13462,N_11332,N_12365);
nand U13463 (N_13463,N_10966,N_11875);
nand U13464 (N_13464,N_10991,N_11922);
xor U13465 (N_13465,N_11953,N_11960);
or U13466 (N_13466,N_11104,N_12121);
nand U13467 (N_13467,N_10601,N_11513);
or U13468 (N_13468,N_11712,N_11274);
and U13469 (N_13469,N_10586,N_10024);
nand U13470 (N_13470,N_10366,N_11149);
nand U13471 (N_13471,N_11796,N_11097);
xnor U13472 (N_13472,N_12174,N_11936);
nand U13473 (N_13473,N_11855,N_11656);
and U13474 (N_13474,N_11345,N_12031);
nand U13475 (N_13475,N_12225,N_11971);
nor U13476 (N_13476,N_11572,N_11685);
nor U13477 (N_13477,N_12085,N_11758);
xnor U13478 (N_13478,N_10115,N_11055);
xor U13479 (N_13479,N_11631,N_11138);
nand U13480 (N_13480,N_12010,N_12251);
xnor U13481 (N_13481,N_12424,N_10629);
xnor U13482 (N_13482,N_11862,N_12186);
nand U13483 (N_13483,N_10538,N_11457);
and U13484 (N_13484,N_11385,N_12032);
and U13485 (N_13485,N_12370,N_10061);
nor U13486 (N_13486,N_12235,N_11210);
xor U13487 (N_13487,N_10690,N_10527);
xnor U13488 (N_13488,N_11848,N_10037);
or U13489 (N_13489,N_11606,N_10713);
and U13490 (N_13490,N_11909,N_11730);
or U13491 (N_13491,N_11713,N_10841);
nor U13492 (N_13492,N_11331,N_10310);
or U13493 (N_13493,N_10996,N_10124);
nand U13494 (N_13494,N_11531,N_12214);
nor U13495 (N_13495,N_11028,N_11236);
nor U13496 (N_13496,N_11155,N_12207);
nand U13497 (N_13497,N_10698,N_10942);
nor U13498 (N_13498,N_11599,N_11298);
nand U13499 (N_13499,N_11580,N_10694);
and U13500 (N_13500,N_10523,N_10709);
nand U13501 (N_13501,N_10666,N_12025);
nand U13502 (N_13502,N_11391,N_10278);
and U13503 (N_13503,N_12327,N_11421);
nand U13504 (N_13504,N_10655,N_11617);
nand U13505 (N_13505,N_11142,N_10060);
xnor U13506 (N_13506,N_10834,N_10196);
or U13507 (N_13507,N_10369,N_11414);
nand U13508 (N_13508,N_10987,N_12005);
xor U13509 (N_13509,N_11537,N_12078);
nand U13510 (N_13510,N_10900,N_12232);
xor U13511 (N_13511,N_10012,N_10546);
xnor U13512 (N_13512,N_11867,N_10884);
xnor U13513 (N_13513,N_12368,N_10636);
and U13514 (N_13514,N_10700,N_11562);
or U13515 (N_13515,N_10570,N_12493);
nor U13516 (N_13516,N_11858,N_11914);
nor U13517 (N_13517,N_12138,N_11280);
and U13518 (N_13518,N_10392,N_12246);
nand U13519 (N_13519,N_12360,N_12432);
or U13520 (N_13520,N_10532,N_11479);
nand U13521 (N_13521,N_11193,N_11339);
xnor U13522 (N_13522,N_12114,N_11818);
nor U13523 (N_13523,N_12315,N_11413);
xor U13524 (N_13524,N_12346,N_12139);
nand U13525 (N_13525,N_10488,N_12176);
or U13526 (N_13526,N_11751,N_12396);
or U13527 (N_13527,N_10596,N_11417);
nand U13528 (N_13528,N_11722,N_10506);
and U13529 (N_13529,N_11416,N_11750);
nand U13530 (N_13530,N_10759,N_10360);
or U13531 (N_13531,N_12059,N_10237);
nor U13532 (N_13532,N_12157,N_11752);
nor U13533 (N_13533,N_10681,N_11740);
xnor U13534 (N_13534,N_11978,N_10783);
nor U13535 (N_13535,N_10782,N_12293);
nand U13536 (N_13536,N_12098,N_12279);
xor U13537 (N_13537,N_12278,N_12115);
and U13538 (N_13538,N_10852,N_11898);
and U13539 (N_13539,N_10020,N_10568);
xnor U13540 (N_13540,N_10623,N_12375);
and U13541 (N_13541,N_10906,N_11076);
or U13542 (N_13542,N_12148,N_10658);
nand U13543 (N_13543,N_10390,N_10336);
and U13544 (N_13544,N_11882,N_12383);
nand U13545 (N_13545,N_11152,N_12072);
nand U13546 (N_13546,N_11643,N_10005);
nor U13547 (N_13547,N_12474,N_10166);
xor U13548 (N_13548,N_11103,N_10156);
nand U13549 (N_13549,N_11616,N_12125);
and U13550 (N_13550,N_10075,N_10267);
and U13551 (N_13551,N_10040,N_11602);
xnor U13552 (N_13552,N_12116,N_11815);
and U13553 (N_13553,N_10260,N_11665);
or U13554 (N_13554,N_10807,N_10139);
or U13555 (N_13555,N_10970,N_10561);
nor U13556 (N_13556,N_10193,N_10950);
nor U13557 (N_13557,N_10140,N_11405);
nand U13558 (N_13558,N_11661,N_11744);
nand U13559 (N_13559,N_11688,N_10142);
xor U13560 (N_13560,N_10079,N_12061);
or U13561 (N_13561,N_10828,N_11863);
or U13562 (N_13562,N_10371,N_11541);
nor U13563 (N_13563,N_11286,N_10422);
and U13564 (N_13564,N_10315,N_11379);
nand U13565 (N_13565,N_11881,N_10720);
and U13566 (N_13566,N_10468,N_10971);
or U13567 (N_13567,N_12335,N_10861);
nand U13568 (N_13568,N_11923,N_11283);
and U13569 (N_13569,N_10715,N_12426);
and U13570 (N_13570,N_11701,N_10874);
and U13571 (N_13571,N_12110,N_11302);
and U13572 (N_13572,N_11047,N_10528);
nor U13573 (N_13573,N_12247,N_12220);
or U13574 (N_13574,N_10565,N_11341);
xnor U13575 (N_13575,N_11119,N_10183);
nor U13576 (N_13576,N_10270,N_12284);
and U13577 (N_13577,N_10929,N_10635);
or U13578 (N_13578,N_10086,N_11250);
and U13579 (N_13579,N_11825,N_10187);
nor U13580 (N_13580,N_12336,N_12067);
or U13581 (N_13581,N_12331,N_10268);
xor U13582 (N_13582,N_11357,N_12146);
xnor U13583 (N_13583,N_10396,N_11748);
and U13584 (N_13584,N_11023,N_10341);
nand U13585 (N_13585,N_11977,N_10595);
xor U13586 (N_13586,N_10727,N_12102);
or U13587 (N_13587,N_10064,N_11689);
xor U13588 (N_13588,N_11272,N_11959);
xor U13589 (N_13589,N_11182,N_11324);
xnor U13590 (N_13590,N_10985,N_10301);
nor U13591 (N_13591,N_12362,N_11189);
or U13592 (N_13592,N_10215,N_12201);
nor U13593 (N_13593,N_10964,N_10934);
and U13594 (N_13594,N_12038,N_12409);
and U13595 (N_13595,N_12108,N_12276);
and U13596 (N_13596,N_11292,N_11360);
or U13597 (N_13597,N_11659,N_10847);
and U13598 (N_13598,N_10600,N_11208);
nor U13599 (N_13599,N_10466,N_10476);
xor U13600 (N_13600,N_10893,N_10762);
nand U13601 (N_13601,N_11203,N_10018);
nor U13602 (N_13602,N_11113,N_10085);
xor U13603 (N_13603,N_12006,N_11674);
xor U13604 (N_13604,N_10763,N_10373);
nor U13605 (N_13605,N_11832,N_11610);
nor U13606 (N_13606,N_12304,N_10773);
nand U13607 (N_13607,N_11738,N_10242);
nand U13608 (N_13608,N_11165,N_10206);
and U13609 (N_13609,N_11527,N_10318);
nor U13610 (N_13610,N_10661,N_11799);
nor U13611 (N_13611,N_11542,N_11029);
and U13612 (N_13612,N_11294,N_11273);
nand U13613 (N_13613,N_11857,N_11122);
and U13614 (N_13614,N_11034,N_10405);
and U13615 (N_13615,N_12333,N_10937);
and U13616 (N_13616,N_11356,N_11364);
and U13617 (N_13617,N_10228,N_11568);
nand U13618 (N_13618,N_12017,N_11630);
nor U13619 (N_13619,N_11747,N_11503);
xnor U13620 (N_13620,N_11515,N_11475);
nor U13621 (N_13621,N_11041,N_12254);
and U13622 (N_13622,N_12431,N_11569);
and U13623 (N_13623,N_10029,N_10633);
and U13624 (N_13624,N_11347,N_10695);
xnor U13625 (N_13625,N_10809,N_11078);
xor U13626 (N_13626,N_12302,N_12390);
or U13627 (N_13627,N_11191,N_10418);
nor U13628 (N_13628,N_11550,N_10548);
nand U13629 (N_13629,N_11407,N_11729);
nor U13630 (N_13630,N_10913,N_10181);
xnor U13631 (N_13631,N_12142,N_11276);
or U13632 (N_13632,N_12143,N_10550);
nand U13633 (N_13633,N_11629,N_10774);
xnor U13634 (N_13634,N_11277,N_11912);
nand U13635 (N_13635,N_10670,N_10717);
xnor U13636 (N_13636,N_10765,N_12167);
and U13637 (N_13637,N_12147,N_10967);
nor U13638 (N_13638,N_11488,N_11700);
or U13639 (N_13639,N_10045,N_11320);
nand U13640 (N_13640,N_11458,N_10816);
xor U13641 (N_13641,N_11641,N_12039);
and U13642 (N_13642,N_11765,N_11940);
xnor U13643 (N_13643,N_12317,N_11437);
or U13644 (N_13644,N_12466,N_10589);
xor U13645 (N_13645,N_12430,N_10317);
and U13646 (N_13646,N_12446,N_12087);
nand U13647 (N_13647,N_12063,N_10013);
and U13648 (N_13648,N_10918,N_10883);
nor U13649 (N_13649,N_10529,N_10739);
and U13650 (N_13650,N_10435,N_11012);
nand U13651 (N_13651,N_10652,N_12264);
xor U13652 (N_13652,N_12320,N_10871);
nand U13653 (N_13653,N_10245,N_10391);
and U13654 (N_13654,N_10328,N_10540);
xor U13655 (N_13655,N_10265,N_11446);
nand U13656 (N_13656,N_10467,N_10756);
nand U13657 (N_13657,N_10394,N_12367);
nor U13658 (N_13658,N_11016,N_12373);
or U13659 (N_13659,N_12020,N_10011);
and U13660 (N_13660,N_11412,N_11261);
nand U13661 (N_13661,N_12425,N_11528);
nand U13662 (N_13662,N_11603,N_12082);
nand U13663 (N_13663,N_10591,N_12462);
and U13664 (N_13664,N_11791,N_12255);
nand U13665 (N_13665,N_10090,N_10726);
nor U13666 (N_13666,N_11070,N_10979);
or U13667 (N_13667,N_11516,N_10072);
and U13668 (N_13668,N_10992,N_11931);
nor U13669 (N_13669,N_12227,N_11908);
or U13670 (N_13670,N_12065,N_12243);
and U13671 (N_13671,N_12453,N_10752);
nand U13672 (N_13672,N_11790,N_10956);
nor U13673 (N_13673,N_12130,N_10958);
xor U13674 (N_13674,N_10917,N_10050);
xor U13675 (N_13675,N_10386,N_10349);
xor U13676 (N_13676,N_11471,N_10100);
or U13677 (N_13677,N_10873,N_10440);
xor U13678 (N_13678,N_10551,N_10949);
and U13679 (N_13679,N_12283,N_11350);
xnor U13680 (N_13680,N_10614,N_11536);
nor U13681 (N_13681,N_10026,N_11132);
nor U13682 (N_13682,N_11008,N_11703);
xor U13683 (N_13683,N_11077,N_11941);
nor U13684 (N_13684,N_10997,N_11307);
nor U13685 (N_13685,N_11396,N_10113);
or U13686 (N_13686,N_11808,N_10106);
nand U13687 (N_13687,N_11762,N_12056);
xor U13688 (N_13688,N_10853,N_10444);
nand U13689 (N_13689,N_12401,N_10594);
nor U13690 (N_13690,N_11813,N_10430);
nor U13691 (N_13691,N_12407,N_12185);
or U13692 (N_13692,N_11776,N_10114);
nor U13693 (N_13693,N_11653,N_11868);
nor U13694 (N_13694,N_11895,N_10576);
nand U13695 (N_13695,N_11731,N_10273);
and U13696 (N_13696,N_11585,N_12221);
or U13697 (N_13697,N_12133,N_10539);
or U13698 (N_13698,N_10203,N_11588);
and U13699 (N_13699,N_11834,N_11798);
and U13700 (N_13700,N_11199,N_12322);
xor U13701 (N_13701,N_12245,N_10982);
nand U13702 (N_13702,N_10194,N_11969);
or U13703 (N_13703,N_10889,N_10575);
or U13704 (N_13704,N_10993,N_11330);
and U13705 (N_13705,N_10400,N_10637);
nand U13706 (N_13706,N_10163,N_12457);
nor U13707 (N_13707,N_10961,N_10850);
nor U13708 (N_13708,N_10808,N_12166);
xor U13709 (N_13709,N_12074,N_12489);
nand U13710 (N_13710,N_11990,N_10178);
nand U13711 (N_13711,N_10008,N_10065);
and U13712 (N_13712,N_12465,N_12483);
and U13713 (N_13713,N_10719,N_11151);
xnor U13714 (N_13714,N_11899,N_11660);
and U13715 (N_13715,N_11186,N_12405);
and U13716 (N_13716,N_11124,N_10285);
and U13717 (N_13717,N_10384,N_12325);
nand U13718 (N_13718,N_12049,N_12137);
xor U13719 (N_13719,N_10810,N_11204);
or U13720 (N_13720,N_10796,N_11015);
nand U13721 (N_13721,N_10522,N_11586);
nand U13722 (N_13722,N_10431,N_12070);
and U13723 (N_13723,N_10824,N_10147);
nand U13724 (N_13724,N_11761,N_11797);
nor U13725 (N_13725,N_11474,N_12212);
and U13726 (N_13726,N_10777,N_11205);
nor U13727 (N_13727,N_11299,N_11258);
and U13728 (N_13728,N_10963,N_11676);
xor U13729 (N_13729,N_11192,N_12041);
or U13730 (N_13730,N_11478,N_10433);
or U13731 (N_13731,N_11807,N_11916);
xnor U13732 (N_13732,N_10456,N_10771);
or U13733 (N_13733,N_12420,N_10541);
xnor U13734 (N_13734,N_10811,N_12093);
nor U13735 (N_13735,N_11230,N_10279);
or U13736 (N_13736,N_11247,N_10784);
nor U13737 (N_13737,N_10066,N_11991);
and U13738 (N_13738,N_10597,N_11670);
or U13739 (N_13739,N_10507,N_12486);
xor U13740 (N_13740,N_11088,N_10622);
xnor U13741 (N_13741,N_10564,N_11020);
and U13742 (N_13742,N_10200,N_10604);
nand U13743 (N_13743,N_11080,N_11032);
or U13744 (N_13744,N_10892,N_10860);
xnor U13745 (N_13745,N_11395,N_11695);
and U13746 (N_13746,N_12073,N_11982);
and U13747 (N_13747,N_10180,N_10706);
nor U13748 (N_13748,N_12386,N_12280);
and U13749 (N_13749,N_12291,N_10920);
xnor U13750 (N_13750,N_11202,N_10159);
nor U13751 (N_13751,N_11986,N_11230);
nor U13752 (N_13752,N_11851,N_11496);
xnor U13753 (N_13753,N_11084,N_12182);
nand U13754 (N_13754,N_12093,N_11645);
nor U13755 (N_13755,N_11471,N_11378);
and U13756 (N_13756,N_10404,N_10275);
or U13757 (N_13757,N_10806,N_10528);
nand U13758 (N_13758,N_10985,N_10968);
and U13759 (N_13759,N_11439,N_10830);
nor U13760 (N_13760,N_10084,N_10296);
and U13761 (N_13761,N_10388,N_10199);
xor U13762 (N_13762,N_10923,N_12107);
and U13763 (N_13763,N_12156,N_11829);
nor U13764 (N_13764,N_11778,N_12025);
nand U13765 (N_13765,N_11572,N_12282);
nor U13766 (N_13766,N_10852,N_10070);
and U13767 (N_13767,N_11416,N_11014);
nor U13768 (N_13768,N_12344,N_10856);
nor U13769 (N_13769,N_12056,N_11371);
nor U13770 (N_13770,N_11557,N_10203);
nand U13771 (N_13771,N_11856,N_10711);
or U13772 (N_13772,N_11076,N_12180);
and U13773 (N_13773,N_11539,N_12131);
and U13774 (N_13774,N_10059,N_10148);
xnor U13775 (N_13775,N_11769,N_10566);
nand U13776 (N_13776,N_10040,N_11853);
nor U13777 (N_13777,N_10383,N_10283);
nor U13778 (N_13778,N_12488,N_12123);
or U13779 (N_13779,N_12182,N_10694);
or U13780 (N_13780,N_12118,N_11096);
nor U13781 (N_13781,N_12481,N_12085);
and U13782 (N_13782,N_10646,N_11902);
or U13783 (N_13783,N_10446,N_11495);
nand U13784 (N_13784,N_11514,N_11697);
or U13785 (N_13785,N_11339,N_10373);
and U13786 (N_13786,N_11079,N_11520);
and U13787 (N_13787,N_10242,N_11117);
and U13788 (N_13788,N_11801,N_11733);
and U13789 (N_13789,N_10117,N_11708);
nand U13790 (N_13790,N_10467,N_10107);
nand U13791 (N_13791,N_11727,N_12326);
nor U13792 (N_13792,N_10099,N_11422);
or U13793 (N_13793,N_10751,N_11409);
nor U13794 (N_13794,N_10732,N_11082);
xnor U13795 (N_13795,N_10041,N_10928);
xor U13796 (N_13796,N_11703,N_11067);
or U13797 (N_13797,N_10124,N_10308);
and U13798 (N_13798,N_11237,N_11790);
nor U13799 (N_13799,N_12143,N_11414);
and U13800 (N_13800,N_10087,N_10411);
nor U13801 (N_13801,N_11870,N_12366);
xnor U13802 (N_13802,N_10439,N_10884);
nor U13803 (N_13803,N_12321,N_11960);
and U13804 (N_13804,N_11580,N_10519);
xor U13805 (N_13805,N_10217,N_10252);
nand U13806 (N_13806,N_11032,N_10157);
xnor U13807 (N_13807,N_10729,N_12366);
xor U13808 (N_13808,N_11987,N_11877);
nor U13809 (N_13809,N_11420,N_10442);
or U13810 (N_13810,N_11081,N_11314);
nand U13811 (N_13811,N_10071,N_10432);
and U13812 (N_13812,N_10688,N_10216);
xnor U13813 (N_13813,N_12124,N_10230);
nand U13814 (N_13814,N_11816,N_11330);
nor U13815 (N_13815,N_11086,N_10790);
xnor U13816 (N_13816,N_10893,N_11725);
and U13817 (N_13817,N_12277,N_10218);
and U13818 (N_13818,N_11826,N_10070);
nand U13819 (N_13819,N_12220,N_12370);
or U13820 (N_13820,N_10705,N_11689);
or U13821 (N_13821,N_10423,N_10665);
or U13822 (N_13822,N_10375,N_10714);
or U13823 (N_13823,N_10697,N_11278);
and U13824 (N_13824,N_11779,N_11557);
xnor U13825 (N_13825,N_10249,N_11217);
and U13826 (N_13826,N_11382,N_12327);
nand U13827 (N_13827,N_11240,N_10974);
xnor U13828 (N_13828,N_11250,N_11580);
nor U13829 (N_13829,N_11230,N_10985);
nand U13830 (N_13830,N_11765,N_11345);
or U13831 (N_13831,N_10830,N_12438);
xor U13832 (N_13832,N_10794,N_10775);
nor U13833 (N_13833,N_11821,N_10591);
nor U13834 (N_13834,N_11387,N_12488);
nand U13835 (N_13835,N_10928,N_10008);
and U13836 (N_13836,N_11707,N_11050);
or U13837 (N_13837,N_10542,N_12443);
and U13838 (N_13838,N_11404,N_11459);
nor U13839 (N_13839,N_10522,N_11160);
xor U13840 (N_13840,N_11322,N_10629);
and U13841 (N_13841,N_12389,N_11834);
nand U13842 (N_13842,N_11389,N_11627);
and U13843 (N_13843,N_11162,N_11171);
or U13844 (N_13844,N_11966,N_11542);
xor U13845 (N_13845,N_11555,N_10267);
or U13846 (N_13846,N_10025,N_10057);
nand U13847 (N_13847,N_12301,N_12460);
or U13848 (N_13848,N_12283,N_11557);
xor U13849 (N_13849,N_10913,N_11571);
and U13850 (N_13850,N_10826,N_11532);
xor U13851 (N_13851,N_11958,N_11561);
or U13852 (N_13852,N_11365,N_12322);
nor U13853 (N_13853,N_10653,N_10457);
xor U13854 (N_13854,N_11296,N_11519);
or U13855 (N_13855,N_10477,N_10419);
nand U13856 (N_13856,N_11402,N_10862);
or U13857 (N_13857,N_12087,N_10716);
nand U13858 (N_13858,N_10453,N_12080);
and U13859 (N_13859,N_11673,N_12456);
xor U13860 (N_13860,N_11989,N_10660);
nor U13861 (N_13861,N_11666,N_10967);
or U13862 (N_13862,N_11508,N_12304);
xnor U13863 (N_13863,N_12261,N_11555);
nor U13864 (N_13864,N_11082,N_11915);
nand U13865 (N_13865,N_11266,N_11020);
xor U13866 (N_13866,N_11217,N_10104);
and U13867 (N_13867,N_11259,N_11642);
xor U13868 (N_13868,N_10006,N_10558);
nand U13869 (N_13869,N_12045,N_10381);
or U13870 (N_13870,N_10304,N_10560);
xnor U13871 (N_13871,N_11620,N_10793);
and U13872 (N_13872,N_10128,N_11081);
nand U13873 (N_13873,N_12435,N_11567);
or U13874 (N_13874,N_11183,N_11943);
and U13875 (N_13875,N_11109,N_11536);
or U13876 (N_13876,N_11438,N_12090);
nand U13877 (N_13877,N_10987,N_10535);
xor U13878 (N_13878,N_10814,N_11923);
xor U13879 (N_13879,N_12199,N_11295);
nor U13880 (N_13880,N_10636,N_11642);
xnor U13881 (N_13881,N_11009,N_11032);
and U13882 (N_13882,N_10624,N_11260);
nand U13883 (N_13883,N_10051,N_11845);
or U13884 (N_13884,N_11556,N_11199);
xor U13885 (N_13885,N_10773,N_10804);
xor U13886 (N_13886,N_10005,N_11125);
nand U13887 (N_13887,N_12462,N_12198);
nand U13888 (N_13888,N_10002,N_12400);
or U13889 (N_13889,N_12224,N_11734);
nor U13890 (N_13890,N_11125,N_11628);
nand U13891 (N_13891,N_10545,N_11579);
nand U13892 (N_13892,N_12013,N_11049);
xor U13893 (N_13893,N_10385,N_10697);
and U13894 (N_13894,N_10539,N_11697);
or U13895 (N_13895,N_10460,N_11006);
and U13896 (N_13896,N_11114,N_11243);
nor U13897 (N_13897,N_11586,N_12331);
nand U13898 (N_13898,N_10502,N_12232);
and U13899 (N_13899,N_12306,N_10917);
nand U13900 (N_13900,N_12441,N_10396);
xnor U13901 (N_13901,N_11592,N_11440);
and U13902 (N_13902,N_11687,N_11762);
or U13903 (N_13903,N_11147,N_12031);
or U13904 (N_13904,N_12080,N_12382);
xnor U13905 (N_13905,N_10838,N_10368);
nor U13906 (N_13906,N_11465,N_11779);
xor U13907 (N_13907,N_10884,N_10054);
xnor U13908 (N_13908,N_10166,N_12206);
xnor U13909 (N_13909,N_10974,N_11133);
nor U13910 (N_13910,N_10270,N_10470);
and U13911 (N_13911,N_10267,N_10349);
and U13912 (N_13912,N_10654,N_11907);
xnor U13913 (N_13913,N_12162,N_11511);
xnor U13914 (N_13914,N_11986,N_11241);
or U13915 (N_13915,N_10494,N_10228);
nor U13916 (N_13916,N_10244,N_10932);
nor U13917 (N_13917,N_11690,N_12133);
xor U13918 (N_13918,N_11319,N_11977);
nor U13919 (N_13919,N_11931,N_11715);
or U13920 (N_13920,N_10641,N_10626);
nor U13921 (N_13921,N_10534,N_11293);
and U13922 (N_13922,N_10685,N_11066);
and U13923 (N_13923,N_11506,N_10502);
xor U13924 (N_13924,N_11902,N_11778);
nor U13925 (N_13925,N_11679,N_12496);
nand U13926 (N_13926,N_10171,N_12043);
nand U13927 (N_13927,N_11726,N_11535);
xnor U13928 (N_13928,N_11003,N_12340);
xor U13929 (N_13929,N_11435,N_10608);
nand U13930 (N_13930,N_10806,N_11126);
nor U13931 (N_13931,N_11709,N_10189);
nor U13932 (N_13932,N_10145,N_10234);
xnor U13933 (N_13933,N_10788,N_12000);
nor U13934 (N_13934,N_11143,N_11076);
or U13935 (N_13935,N_10400,N_11303);
and U13936 (N_13936,N_10736,N_10686);
and U13937 (N_13937,N_11295,N_11892);
nor U13938 (N_13938,N_11233,N_10771);
xnor U13939 (N_13939,N_10331,N_12177);
xor U13940 (N_13940,N_12130,N_11342);
or U13941 (N_13941,N_11694,N_10163);
or U13942 (N_13942,N_10566,N_10629);
and U13943 (N_13943,N_11026,N_12406);
and U13944 (N_13944,N_10514,N_11839);
xnor U13945 (N_13945,N_10122,N_10727);
and U13946 (N_13946,N_12442,N_11525);
nand U13947 (N_13947,N_10924,N_12429);
or U13948 (N_13948,N_10579,N_11243);
xor U13949 (N_13949,N_11658,N_10153);
xnor U13950 (N_13950,N_12298,N_10408);
nor U13951 (N_13951,N_12263,N_10371);
nor U13952 (N_13952,N_10501,N_10454);
nor U13953 (N_13953,N_11346,N_11367);
and U13954 (N_13954,N_11697,N_12067);
xnor U13955 (N_13955,N_11040,N_10268);
and U13956 (N_13956,N_12399,N_11685);
or U13957 (N_13957,N_11087,N_10684);
nand U13958 (N_13958,N_12390,N_11467);
and U13959 (N_13959,N_11789,N_10438);
nand U13960 (N_13960,N_10840,N_10041);
nand U13961 (N_13961,N_12193,N_11059);
or U13962 (N_13962,N_10811,N_10018);
or U13963 (N_13963,N_10141,N_11374);
or U13964 (N_13964,N_10739,N_12472);
nor U13965 (N_13965,N_10379,N_11896);
nor U13966 (N_13966,N_11707,N_11887);
and U13967 (N_13967,N_11533,N_11468);
nand U13968 (N_13968,N_11127,N_11186);
xor U13969 (N_13969,N_11376,N_10200);
nor U13970 (N_13970,N_10257,N_11691);
xnor U13971 (N_13971,N_10391,N_12393);
xnor U13972 (N_13972,N_10427,N_12476);
nand U13973 (N_13973,N_10162,N_10939);
xor U13974 (N_13974,N_11780,N_10565);
nor U13975 (N_13975,N_10385,N_11047);
nor U13976 (N_13976,N_11930,N_11692);
nand U13977 (N_13977,N_12070,N_10563);
or U13978 (N_13978,N_12208,N_11552);
and U13979 (N_13979,N_11486,N_11793);
xor U13980 (N_13980,N_11842,N_10251);
nor U13981 (N_13981,N_11032,N_11678);
or U13982 (N_13982,N_12479,N_11072);
or U13983 (N_13983,N_10175,N_10504);
nor U13984 (N_13984,N_11965,N_10119);
and U13985 (N_13985,N_10361,N_11718);
and U13986 (N_13986,N_12498,N_10462);
and U13987 (N_13987,N_10370,N_10319);
or U13988 (N_13988,N_10852,N_11837);
xor U13989 (N_13989,N_10068,N_12153);
nor U13990 (N_13990,N_10291,N_12242);
or U13991 (N_13991,N_11923,N_10554);
and U13992 (N_13992,N_11513,N_10996);
or U13993 (N_13993,N_11640,N_11144);
nand U13994 (N_13994,N_10429,N_10056);
xnor U13995 (N_13995,N_12315,N_10809);
nand U13996 (N_13996,N_11099,N_10425);
and U13997 (N_13997,N_11549,N_10736);
or U13998 (N_13998,N_11671,N_10076);
nor U13999 (N_13999,N_11011,N_12189);
and U14000 (N_14000,N_11094,N_11786);
or U14001 (N_14001,N_11867,N_10374);
xnor U14002 (N_14002,N_10140,N_11973);
nand U14003 (N_14003,N_12446,N_10469);
and U14004 (N_14004,N_10652,N_11552);
nand U14005 (N_14005,N_11617,N_11750);
nand U14006 (N_14006,N_11232,N_12333);
or U14007 (N_14007,N_10399,N_11274);
or U14008 (N_14008,N_12427,N_12053);
xnor U14009 (N_14009,N_10443,N_11069);
or U14010 (N_14010,N_12313,N_11089);
and U14011 (N_14011,N_10586,N_12492);
xor U14012 (N_14012,N_10057,N_11811);
nand U14013 (N_14013,N_12014,N_12359);
nor U14014 (N_14014,N_11034,N_10330);
nand U14015 (N_14015,N_10849,N_12050);
nand U14016 (N_14016,N_11786,N_11630);
or U14017 (N_14017,N_10726,N_11155);
xor U14018 (N_14018,N_10857,N_10227);
nor U14019 (N_14019,N_12137,N_12067);
nor U14020 (N_14020,N_10490,N_10963);
nand U14021 (N_14021,N_12390,N_11859);
xor U14022 (N_14022,N_11220,N_10758);
and U14023 (N_14023,N_12351,N_11425);
nor U14024 (N_14024,N_12362,N_10728);
nor U14025 (N_14025,N_11119,N_12399);
or U14026 (N_14026,N_11394,N_10834);
xor U14027 (N_14027,N_10326,N_11215);
xnor U14028 (N_14028,N_10717,N_12268);
nor U14029 (N_14029,N_12496,N_10902);
or U14030 (N_14030,N_10136,N_10396);
or U14031 (N_14031,N_10083,N_11653);
and U14032 (N_14032,N_11490,N_10992);
nand U14033 (N_14033,N_10401,N_10172);
or U14034 (N_14034,N_11284,N_10158);
nor U14035 (N_14035,N_12048,N_10353);
xnor U14036 (N_14036,N_11333,N_12003);
and U14037 (N_14037,N_10763,N_11875);
xor U14038 (N_14038,N_11338,N_11799);
nand U14039 (N_14039,N_11048,N_11465);
or U14040 (N_14040,N_12416,N_10943);
or U14041 (N_14041,N_10668,N_10192);
nand U14042 (N_14042,N_11583,N_11109);
xor U14043 (N_14043,N_11950,N_11681);
and U14044 (N_14044,N_10907,N_10342);
and U14045 (N_14045,N_10786,N_12044);
or U14046 (N_14046,N_10935,N_11348);
xnor U14047 (N_14047,N_11174,N_11068);
xnor U14048 (N_14048,N_11479,N_11334);
nand U14049 (N_14049,N_10928,N_10848);
and U14050 (N_14050,N_11423,N_11861);
and U14051 (N_14051,N_11127,N_10847);
and U14052 (N_14052,N_11724,N_11148);
nor U14053 (N_14053,N_11140,N_10962);
nand U14054 (N_14054,N_12071,N_10075);
nand U14055 (N_14055,N_11514,N_11080);
xor U14056 (N_14056,N_11242,N_11431);
nand U14057 (N_14057,N_11577,N_11352);
and U14058 (N_14058,N_10123,N_11777);
xor U14059 (N_14059,N_10208,N_11439);
nand U14060 (N_14060,N_11111,N_11901);
nor U14061 (N_14061,N_12200,N_12390);
xor U14062 (N_14062,N_11048,N_11112);
xor U14063 (N_14063,N_10390,N_11887);
nor U14064 (N_14064,N_10916,N_12155);
or U14065 (N_14065,N_10035,N_11191);
and U14066 (N_14066,N_12113,N_11607);
nor U14067 (N_14067,N_12132,N_11678);
nor U14068 (N_14068,N_10292,N_10677);
and U14069 (N_14069,N_11511,N_11258);
or U14070 (N_14070,N_12216,N_10571);
nor U14071 (N_14071,N_12397,N_12390);
nor U14072 (N_14072,N_10496,N_11984);
and U14073 (N_14073,N_12368,N_12133);
xor U14074 (N_14074,N_11752,N_11599);
xor U14075 (N_14075,N_10992,N_11902);
and U14076 (N_14076,N_12235,N_10821);
nor U14077 (N_14077,N_11318,N_10738);
xnor U14078 (N_14078,N_10216,N_12217);
nand U14079 (N_14079,N_10969,N_10906);
xnor U14080 (N_14080,N_10676,N_11570);
and U14081 (N_14081,N_12208,N_12261);
or U14082 (N_14082,N_11707,N_10003);
nor U14083 (N_14083,N_11278,N_10130);
xor U14084 (N_14084,N_10614,N_12397);
or U14085 (N_14085,N_10208,N_11173);
nand U14086 (N_14086,N_10908,N_12125);
or U14087 (N_14087,N_11814,N_10588);
nor U14088 (N_14088,N_10853,N_10259);
nor U14089 (N_14089,N_10248,N_10451);
nand U14090 (N_14090,N_11117,N_11744);
xnor U14091 (N_14091,N_10127,N_11987);
and U14092 (N_14092,N_11166,N_10316);
xor U14093 (N_14093,N_11118,N_12337);
nor U14094 (N_14094,N_12191,N_10456);
and U14095 (N_14095,N_10294,N_11046);
nor U14096 (N_14096,N_10635,N_11458);
or U14097 (N_14097,N_11881,N_12310);
nand U14098 (N_14098,N_10003,N_11086);
and U14099 (N_14099,N_11846,N_11498);
or U14100 (N_14100,N_12333,N_12000);
and U14101 (N_14101,N_11096,N_11669);
nor U14102 (N_14102,N_12438,N_11202);
nor U14103 (N_14103,N_10866,N_10026);
nand U14104 (N_14104,N_12396,N_11311);
xnor U14105 (N_14105,N_12463,N_11749);
or U14106 (N_14106,N_11376,N_10184);
or U14107 (N_14107,N_12040,N_10170);
nand U14108 (N_14108,N_11759,N_10533);
or U14109 (N_14109,N_12155,N_10387);
nor U14110 (N_14110,N_10800,N_12130);
xnor U14111 (N_14111,N_10932,N_11769);
or U14112 (N_14112,N_10232,N_11876);
and U14113 (N_14113,N_10688,N_10078);
nand U14114 (N_14114,N_10979,N_10504);
xnor U14115 (N_14115,N_12202,N_10926);
xor U14116 (N_14116,N_11407,N_10576);
xnor U14117 (N_14117,N_11411,N_10945);
and U14118 (N_14118,N_12415,N_11345);
xor U14119 (N_14119,N_10809,N_11396);
nor U14120 (N_14120,N_12300,N_10113);
and U14121 (N_14121,N_12366,N_10926);
nand U14122 (N_14122,N_11651,N_10656);
and U14123 (N_14123,N_12376,N_10923);
nand U14124 (N_14124,N_10111,N_12441);
nand U14125 (N_14125,N_10257,N_11235);
nand U14126 (N_14126,N_11641,N_10388);
nand U14127 (N_14127,N_12465,N_11890);
nand U14128 (N_14128,N_11176,N_11064);
nand U14129 (N_14129,N_12216,N_11009);
and U14130 (N_14130,N_11902,N_10746);
xor U14131 (N_14131,N_11672,N_11831);
nor U14132 (N_14132,N_10204,N_12235);
or U14133 (N_14133,N_11960,N_11129);
xnor U14134 (N_14134,N_11595,N_10248);
nand U14135 (N_14135,N_12462,N_12332);
nand U14136 (N_14136,N_11476,N_12170);
and U14137 (N_14137,N_11937,N_11227);
xor U14138 (N_14138,N_10652,N_10608);
or U14139 (N_14139,N_11572,N_10909);
xnor U14140 (N_14140,N_11651,N_10554);
nor U14141 (N_14141,N_12386,N_11537);
and U14142 (N_14142,N_11703,N_11900);
or U14143 (N_14143,N_10527,N_10076);
and U14144 (N_14144,N_12127,N_12285);
nand U14145 (N_14145,N_12017,N_11593);
xnor U14146 (N_14146,N_10162,N_12265);
or U14147 (N_14147,N_11035,N_10687);
or U14148 (N_14148,N_10939,N_11997);
nand U14149 (N_14149,N_11660,N_11471);
xnor U14150 (N_14150,N_11737,N_10607);
and U14151 (N_14151,N_10210,N_10287);
or U14152 (N_14152,N_10513,N_12127);
and U14153 (N_14153,N_11009,N_10223);
nand U14154 (N_14154,N_12086,N_12255);
nand U14155 (N_14155,N_11022,N_11449);
and U14156 (N_14156,N_11143,N_10729);
xnor U14157 (N_14157,N_11385,N_12454);
xnor U14158 (N_14158,N_11143,N_10128);
xor U14159 (N_14159,N_12049,N_11683);
nand U14160 (N_14160,N_11097,N_11598);
nand U14161 (N_14161,N_10546,N_10630);
xnor U14162 (N_14162,N_11902,N_11112);
and U14163 (N_14163,N_10415,N_11779);
xnor U14164 (N_14164,N_12152,N_11264);
or U14165 (N_14165,N_10939,N_11038);
and U14166 (N_14166,N_11134,N_10487);
xor U14167 (N_14167,N_10992,N_11823);
nand U14168 (N_14168,N_11674,N_10030);
nand U14169 (N_14169,N_10741,N_10501);
nor U14170 (N_14170,N_11500,N_11168);
and U14171 (N_14171,N_11600,N_10472);
nor U14172 (N_14172,N_12458,N_11866);
or U14173 (N_14173,N_11810,N_11608);
and U14174 (N_14174,N_11227,N_10158);
and U14175 (N_14175,N_11194,N_10409);
and U14176 (N_14176,N_11854,N_11306);
nor U14177 (N_14177,N_12339,N_12141);
and U14178 (N_14178,N_12040,N_10241);
or U14179 (N_14179,N_12148,N_10490);
or U14180 (N_14180,N_10619,N_11881);
nor U14181 (N_14181,N_11453,N_10532);
nor U14182 (N_14182,N_11333,N_11727);
or U14183 (N_14183,N_10753,N_10142);
or U14184 (N_14184,N_12268,N_11225);
or U14185 (N_14185,N_11465,N_11469);
and U14186 (N_14186,N_11055,N_10624);
and U14187 (N_14187,N_11974,N_10397);
or U14188 (N_14188,N_12190,N_10944);
nand U14189 (N_14189,N_10134,N_11432);
nand U14190 (N_14190,N_11120,N_10290);
xnor U14191 (N_14191,N_10893,N_10581);
nand U14192 (N_14192,N_10508,N_10763);
or U14193 (N_14193,N_11562,N_11814);
nor U14194 (N_14194,N_10166,N_11842);
or U14195 (N_14195,N_10490,N_10719);
nand U14196 (N_14196,N_11850,N_10101);
nor U14197 (N_14197,N_11180,N_10960);
nor U14198 (N_14198,N_11807,N_10234);
and U14199 (N_14199,N_11556,N_10993);
or U14200 (N_14200,N_12125,N_12441);
nand U14201 (N_14201,N_10442,N_10328);
and U14202 (N_14202,N_11180,N_10784);
or U14203 (N_14203,N_12091,N_11676);
nand U14204 (N_14204,N_11882,N_11280);
nand U14205 (N_14205,N_12013,N_10088);
nand U14206 (N_14206,N_12492,N_11736);
xnor U14207 (N_14207,N_11939,N_11425);
nor U14208 (N_14208,N_10962,N_10348);
and U14209 (N_14209,N_10482,N_11134);
nor U14210 (N_14210,N_11747,N_10311);
nand U14211 (N_14211,N_11508,N_12460);
or U14212 (N_14212,N_11590,N_10068);
or U14213 (N_14213,N_10665,N_11962);
or U14214 (N_14214,N_11983,N_11017);
or U14215 (N_14215,N_10795,N_10996);
and U14216 (N_14216,N_10003,N_10035);
nand U14217 (N_14217,N_10771,N_11909);
nand U14218 (N_14218,N_12413,N_10949);
and U14219 (N_14219,N_11257,N_11911);
and U14220 (N_14220,N_12405,N_10349);
nor U14221 (N_14221,N_11282,N_11782);
and U14222 (N_14222,N_10061,N_10829);
and U14223 (N_14223,N_11421,N_11247);
and U14224 (N_14224,N_11602,N_11338);
and U14225 (N_14225,N_11701,N_11992);
nand U14226 (N_14226,N_11655,N_11585);
and U14227 (N_14227,N_10456,N_10095);
nor U14228 (N_14228,N_11899,N_10232);
nand U14229 (N_14229,N_11939,N_10361);
nand U14230 (N_14230,N_11511,N_12127);
or U14231 (N_14231,N_10871,N_10476);
xnor U14232 (N_14232,N_12499,N_11365);
and U14233 (N_14233,N_12126,N_11602);
xor U14234 (N_14234,N_11779,N_12414);
and U14235 (N_14235,N_10750,N_11239);
xor U14236 (N_14236,N_11841,N_12331);
or U14237 (N_14237,N_11456,N_12497);
and U14238 (N_14238,N_11221,N_11561);
nor U14239 (N_14239,N_11085,N_11190);
nor U14240 (N_14240,N_10720,N_12054);
nand U14241 (N_14241,N_12340,N_11504);
and U14242 (N_14242,N_10298,N_12152);
xor U14243 (N_14243,N_11304,N_10009);
nor U14244 (N_14244,N_10091,N_10006);
and U14245 (N_14245,N_10992,N_11772);
nor U14246 (N_14246,N_11588,N_11244);
xor U14247 (N_14247,N_11596,N_11365);
nor U14248 (N_14248,N_10971,N_12354);
or U14249 (N_14249,N_11975,N_12139);
nor U14250 (N_14250,N_10437,N_10213);
and U14251 (N_14251,N_10956,N_10221);
and U14252 (N_14252,N_10449,N_10442);
nor U14253 (N_14253,N_11505,N_10932);
xor U14254 (N_14254,N_10356,N_12416);
and U14255 (N_14255,N_12333,N_11350);
or U14256 (N_14256,N_12381,N_11177);
nor U14257 (N_14257,N_11494,N_11794);
xnor U14258 (N_14258,N_11212,N_12455);
nor U14259 (N_14259,N_12021,N_11188);
xor U14260 (N_14260,N_11756,N_11095);
and U14261 (N_14261,N_11304,N_12274);
or U14262 (N_14262,N_11924,N_11914);
nand U14263 (N_14263,N_11296,N_10865);
and U14264 (N_14264,N_10448,N_10081);
and U14265 (N_14265,N_12174,N_11364);
nand U14266 (N_14266,N_11362,N_11505);
xnor U14267 (N_14267,N_10728,N_11583);
nor U14268 (N_14268,N_10800,N_11044);
and U14269 (N_14269,N_10111,N_11623);
or U14270 (N_14270,N_11773,N_10994);
nand U14271 (N_14271,N_11388,N_11525);
and U14272 (N_14272,N_11988,N_10803);
nor U14273 (N_14273,N_12075,N_11429);
xnor U14274 (N_14274,N_11956,N_10219);
and U14275 (N_14275,N_11392,N_10628);
or U14276 (N_14276,N_12123,N_10615);
xor U14277 (N_14277,N_11684,N_10236);
nor U14278 (N_14278,N_10380,N_11245);
xor U14279 (N_14279,N_10719,N_10977);
xor U14280 (N_14280,N_10459,N_12232);
or U14281 (N_14281,N_10970,N_10379);
or U14282 (N_14282,N_11153,N_11639);
and U14283 (N_14283,N_11291,N_11362);
xor U14284 (N_14284,N_10652,N_10215);
nor U14285 (N_14285,N_11939,N_11639);
and U14286 (N_14286,N_11180,N_11806);
xnor U14287 (N_14287,N_11536,N_10231);
nand U14288 (N_14288,N_10964,N_10476);
and U14289 (N_14289,N_10005,N_11510);
nand U14290 (N_14290,N_10546,N_11718);
nor U14291 (N_14291,N_10314,N_10142);
nor U14292 (N_14292,N_12051,N_12310);
nand U14293 (N_14293,N_11776,N_10652);
xor U14294 (N_14294,N_11997,N_11760);
xor U14295 (N_14295,N_11390,N_10251);
xor U14296 (N_14296,N_10723,N_10903);
or U14297 (N_14297,N_11336,N_11799);
nor U14298 (N_14298,N_10734,N_10051);
nor U14299 (N_14299,N_10089,N_11075);
and U14300 (N_14300,N_11880,N_11076);
nor U14301 (N_14301,N_12021,N_10615);
or U14302 (N_14302,N_12095,N_11805);
nor U14303 (N_14303,N_11216,N_10977);
nor U14304 (N_14304,N_10644,N_10818);
or U14305 (N_14305,N_11491,N_11290);
or U14306 (N_14306,N_12341,N_11828);
xor U14307 (N_14307,N_11849,N_10873);
xor U14308 (N_14308,N_10820,N_11845);
or U14309 (N_14309,N_10148,N_10265);
and U14310 (N_14310,N_10267,N_11695);
nand U14311 (N_14311,N_10659,N_12178);
and U14312 (N_14312,N_11176,N_11784);
and U14313 (N_14313,N_10606,N_12402);
xor U14314 (N_14314,N_11961,N_11054);
nand U14315 (N_14315,N_12096,N_11767);
or U14316 (N_14316,N_10794,N_12451);
or U14317 (N_14317,N_12419,N_11518);
or U14318 (N_14318,N_11024,N_11332);
nand U14319 (N_14319,N_10805,N_12198);
nor U14320 (N_14320,N_11303,N_10898);
nor U14321 (N_14321,N_11076,N_11522);
xnor U14322 (N_14322,N_11790,N_11365);
nor U14323 (N_14323,N_11302,N_11587);
nor U14324 (N_14324,N_10905,N_10166);
and U14325 (N_14325,N_11124,N_10527);
or U14326 (N_14326,N_12004,N_11108);
nor U14327 (N_14327,N_11522,N_10209);
or U14328 (N_14328,N_10222,N_10499);
nand U14329 (N_14329,N_10092,N_11433);
xnor U14330 (N_14330,N_12408,N_10753);
and U14331 (N_14331,N_10269,N_11746);
nand U14332 (N_14332,N_10187,N_11293);
or U14333 (N_14333,N_10023,N_10096);
and U14334 (N_14334,N_10057,N_12212);
and U14335 (N_14335,N_11766,N_12062);
xnor U14336 (N_14336,N_12089,N_12033);
and U14337 (N_14337,N_10297,N_11445);
nand U14338 (N_14338,N_12100,N_11351);
nand U14339 (N_14339,N_10203,N_11855);
nor U14340 (N_14340,N_12405,N_12047);
nor U14341 (N_14341,N_10705,N_10708);
nand U14342 (N_14342,N_10194,N_11715);
xor U14343 (N_14343,N_10674,N_11482);
nor U14344 (N_14344,N_10589,N_11532);
nand U14345 (N_14345,N_11963,N_10874);
nor U14346 (N_14346,N_11570,N_11189);
xor U14347 (N_14347,N_10470,N_11976);
xnor U14348 (N_14348,N_10119,N_10811);
nand U14349 (N_14349,N_10319,N_12152);
xor U14350 (N_14350,N_10738,N_10200);
or U14351 (N_14351,N_12186,N_12276);
xnor U14352 (N_14352,N_10632,N_11880);
and U14353 (N_14353,N_11653,N_10060);
nand U14354 (N_14354,N_12442,N_11904);
and U14355 (N_14355,N_11146,N_10426);
nand U14356 (N_14356,N_12125,N_11934);
and U14357 (N_14357,N_12491,N_11434);
nand U14358 (N_14358,N_12233,N_12325);
nor U14359 (N_14359,N_10573,N_11690);
nor U14360 (N_14360,N_11634,N_12272);
and U14361 (N_14361,N_10425,N_11114);
nor U14362 (N_14362,N_10118,N_12381);
and U14363 (N_14363,N_12238,N_10313);
or U14364 (N_14364,N_10276,N_11661);
and U14365 (N_14365,N_11759,N_10395);
and U14366 (N_14366,N_11285,N_11317);
nor U14367 (N_14367,N_10579,N_10787);
xnor U14368 (N_14368,N_10745,N_12115);
nor U14369 (N_14369,N_12274,N_11501);
nand U14370 (N_14370,N_10468,N_11281);
nand U14371 (N_14371,N_11323,N_10923);
nand U14372 (N_14372,N_12432,N_10807);
and U14373 (N_14373,N_10031,N_10568);
nand U14374 (N_14374,N_11930,N_11994);
nor U14375 (N_14375,N_10203,N_10225);
nand U14376 (N_14376,N_11818,N_10045);
and U14377 (N_14377,N_10043,N_11531);
nor U14378 (N_14378,N_11246,N_10648);
nor U14379 (N_14379,N_11629,N_12423);
nand U14380 (N_14380,N_12033,N_10802);
nor U14381 (N_14381,N_11218,N_10941);
or U14382 (N_14382,N_11470,N_10702);
or U14383 (N_14383,N_12210,N_11565);
or U14384 (N_14384,N_10754,N_12330);
or U14385 (N_14385,N_11364,N_10731);
nor U14386 (N_14386,N_10236,N_10191);
xor U14387 (N_14387,N_11072,N_12011);
xnor U14388 (N_14388,N_10517,N_10578);
xnor U14389 (N_14389,N_10437,N_12498);
nand U14390 (N_14390,N_10638,N_10963);
nand U14391 (N_14391,N_11920,N_10047);
nand U14392 (N_14392,N_11335,N_10051);
or U14393 (N_14393,N_12293,N_11209);
xnor U14394 (N_14394,N_11122,N_11954);
nor U14395 (N_14395,N_10444,N_11070);
nand U14396 (N_14396,N_12225,N_11667);
and U14397 (N_14397,N_11320,N_11884);
or U14398 (N_14398,N_11390,N_10738);
nor U14399 (N_14399,N_10198,N_12134);
and U14400 (N_14400,N_11891,N_11760);
and U14401 (N_14401,N_10039,N_10145);
or U14402 (N_14402,N_10085,N_10379);
or U14403 (N_14403,N_10714,N_10472);
or U14404 (N_14404,N_10243,N_10194);
xnor U14405 (N_14405,N_12263,N_10049);
or U14406 (N_14406,N_11370,N_10298);
or U14407 (N_14407,N_12444,N_12336);
xnor U14408 (N_14408,N_10533,N_10666);
or U14409 (N_14409,N_11052,N_12202);
nor U14410 (N_14410,N_11798,N_12361);
nor U14411 (N_14411,N_10848,N_12168);
xor U14412 (N_14412,N_11568,N_11040);
or U14413 (N_14413,N_11040,N_11495);
or U14414 (N_14414,N_11871,N_10231);
and U14415 (N_14415,N_12267,N_11781);
and U14416 (N_14416,N_12280,N_12246);
or U14417 (N_14417,N_10406,N_11255);
nor U14418 (N_14418,N_11659,N_11845);
nor U14419 (N_14419,N_12152,N_12238);
and U14420 (N_14420,N_10510,N_11801);
nand U14421 (N_14421,N_10943,N_10403);
or U14422 (N_14422,N_11161,N_10279);
nand U14423 (N_14423,N_10177,N_10232);
nand U14424 (N_14424,N_10000,N_11761);
xor U14425 (N_14425,N_11410,N_11461);
nor U14426 (N_14426,N_11722,N_10434);
nand U14427 (N_14427,N_10827,N_12124);
and U14428 (N_14428,N_10188,N_11933);
xor U14429 (N_14429,N_12485,N_11248);
nand U14430 (N_14430,N_10266,N_12153);
xor U14431 (N_14431,N_12479,N_11842);
nor U14432 (N_14432,N_11410,N_11242);
or U14433 (N_14433,N_10302,N_10245);
nand U14434 (N_14434,N_10581,N_11418);
nand U14435 (N_14435,N_11073,N_10103);
xnor U14436 (N_14436,N_11958,N_10703);
nand U14437 (N_14437,N_12288,N_11747);
and U14438 (N_14438,N_11101,N_12251);
or U14439 (N_14439,N_11144,N_12058);
and U14440 (N_14440,N_11005,N_11028);
and U14441 (N_14441,N_10184,N_12296);
xor U14442 (N_14442,N_10047,N_10733);
or U14443 (N_14443,N_12064,N_10964);
nand U14444 (N_14444,N_10414,N_10303);
nor U14445 (N_14445,N_10241,N_12198);
nor U14446 (N_14446,N_12458,N_12321);
xnor U14447 (N_14447,N_11767,N_12371);
xor U14448 (N_14448,N_12298,N_11192);
xnor U14449 (N_14449,N_10750,N_11049);
and U14450 (N_14450,N_10973,N_11724);
xnor U14451 (N_14451,N_11850,N_12296);
xor U14452 (N_14452,N_10651,N_10300);
xor U14453 (N_14453,N_12451,N_11933);
xnor U14454 (N_14454,N_11788,N_10317);
or U14455 (N_14455,N_10576,N_10032);
nand U14456 (N_14456,N_11185,N_10808);
and U14457 (N_14457,N_10753,N_12092);
or U14458 (N_14458,N_11673,N_10175);
xnor U14459 (N_14459,N_10901,N_10416);
and U14460 (N_14460,N_11308,N_12450);
or U14461 (N_14461,N_12339,N_11046);
nor U14462 (N_14462,N_10630,N_12238);
xnor U14463 (N_14463,N_10977,N_11957);
or U14464 (N_14464,N_11508,N_10846);
or U14465 (N_14465,N_10922,N_12159);
nor U14466 (N_14466,N_11497,N_11804);
nor U14467 (N_14467,N_11795,N_12328);
nand U14468 (N_14468,N_10003,N_11455);
or U14469 (N_14469,N_10297,N_11852);
and U14470 (N_14470,N_11063,N_12420);
xnor U14471 (N_14471,N_11463,N_11053);
nor U14472 (N_14472,N_12420,N_10063);
xnor U14473 (N_14473,N_10611,N_11380);
nand U14474 (N_14474,N_12072,N_10185);
xor U14475 (N_14475,N_12277,N_12025);
nand U14476 (N_14476,N_10031,N_10805);
nor U14477 (N_14477,N_12263,N_10273);
and U14478 (N_14478,N_10945,N_11114);
nand U14479 (N_14479,N_11952,N_11959);
or U14480 (N_14480,N_12311,N_12073);
and U14481 (N_14481,N_11539,N_12449);
nor U14482 (N_14482,N_10209,N_12435);
nand U14483 (N_14483,N_10200,N_11214);
nor U14484 (N_14484,N_10340,N_11333);
or U14485 (N_14485,N_10036,N_11828);
nor U14486 (N_14486,N_11750,N_12298);
and U14487 (N_14487,N_12131,N_12388);
nand U14488 (N_14488,N_12003,N_10861);
xnor U14489 (N_14489,N_12481,N_10098);
or U14490 (N_14490,N_11877,N_12129);
or U14491 (N_14491,N_11280,N_11935);
nand U14492 (N_14492,N_12141,N_11195);
nand U14493 (N_14493,N_12119,N_11530);
xnor U14494 (N_14494,N_11526,N_11765);
xor U14495 (N_14495,N_11678,N_10142);
nor U14496 (N_14496,N_12032,N_10057);
or U14497 (N_14497,N_11569,N_10702);
xor U14498 (N_14498,N_11597,N_12421);
nor U14499 (N_14499,N_12363,N_10995);
and U14500 (N_14500,N_11875,N_12325);
or U14501 (N_14501,N_12321,N_10358);
or U14502 (N_14502,N_10875,N_11744);
nand U14503 (N_14503,N_10432,N_10653);
nor U14504 (N_14504,N_11413,N_10212);
and U14505 (N_14505,N_10797,N_10735);
and U14506 (N_14506,N_12159,N_10822);
nor U14507 (N_14507,N_10883,N_10410);
or U14508 (N_14508,N_12397,N_10378);
xnor U14509 (N_14509,N_11505,N_11353);
xnor U14510 (N_14510,N_12478,N_10680);
and U14511 (N_14511,N_10974,N_11698);
and U14512 (N_14512,N_11559,N_11392);
or U14513 (N_14513,N_11414,N_11710);
and U14514 (N_14514,N_10402,N_10514);
or U14515 (N_14515,N_10977,N_11626);
or U14516 (N_14516,N_11379,N_10925);
xor U14517 (N_14517,N_10621,N_11518);
nand U14518 (N_14518,N_10623,N_10607);
xor U14519 (N_14519,N_10813,N_11969);
xnor U14520 (N_14520,N_11414,N_12490);
or U14521 (N_14521,N_10476,N_12478);
nor U14522 (N_14522,N_10588,N_10674);
xor U14523 (N_14523,N_12254,N_10114);
nand U14524 (N_14524,N_10757,N_10259);
or U14525 (N_14525,N_12199,N_12393);
or U14526 (N_14526,N_11533,N_10805);
nand U14527 (N_14527,N_10579,N_12219);
or U14528 (N_14528,N_11815,N_10373);
nor U14529 (N_14529,N_11658,N_11072);
and U14530 (N_14530,N_10110,N_11809);
and U14531 (N_14531,N_11607,N_10552);
or U14532 (N_14532,N_11849,N_10989);
xnor U14533 (N_14533,N_12229,N_10798);
nor U14534 (N_14534,N_11859,N_10924);
nand U14535 (N_14535,N_12345,N_12347);
nand U14536 (N_14536,N_11831,N_11724);
and U14537 (N_14537,N_12065,N_10685);
nand U14538 (N_14538,N_11307,N_12316);
or U14539 (N_14539,N_10605,N_10760);
and U14540 (N_14540,N_10702,N_11532);
nand U14541 (N_14541,N_10611,N_11751);
and U14542 (N_14542,N_12408,N_12465);
nor U14543 (N_14543,N_12372,N_10822);
or U14544 (N_14544,N_12259,N_11167);
and U14545 (N_14545,N_10266,N_11127);
xor U14546 (N_14546,N_10260,N_11237);
nand U14547 (N_14547,N_11024,N_12063);
or U14548 (N_14548,N_11171,N_11532);
nand U14549 (N_14549,N_10168,N_10515);
or U14550 (N_14550,N_11039,N_10494);
nand U14551 (N_14551,N_10881,N_11069);
and U14552 (N_14552,N_10947,N_11247);
xor U14553 (N_14553,N_10290,N_11208);
and U14554 (N_14554,N_12327,N_11349);
xnor U14555 (N_14555,N_10929,N_11767);
nand U14556 (N_14556,N_10966,N_12447);
nand U14557 (N_14557,N_12057,N_11476);
nand U14558 (N_14558,N_11171,N_10626);
nor U14559 (N_14559,N_11810,N_12404);
and U14560 (N_14560,N_10777,N_10957);
xnor U14561 (N_14561,N_10848,N_11622);
xnor U14562 (N_14562,N_12202,N_11764);
nand U14563 (N_14563,N_10884,N_11645);
nor U14564 (N_14564,N_12082,N_12404);
or U14565 (N_14565,N_12053,N_11297);
nand U14566 (N_14566,N_10901,N_10384);
or U14567 (N_14567,N_11110,N_10582);
nor U14568 (N_14568,N_10584,N_11389);
nor U14569 (N_14569,N_11684,N_10573);
nor U14570 (N_14570,N_10492,N_10669);
or U14571 (N_14571,N_12129,N_11722);
xnor U14572 (N_14572,N_12017,N_10390);
nor U14573 (N_14573,N_11153,N_11517);
xor U14574 (N_14574,N_11471,N_10419);
xnor U14575 (N_14575,N_11719,N_11044);
nor U14576 (N_14576,N_11599,N_10605);
nand U14577 (N_14577,N_11705,N_10597);
or U14578 (N_14578,N_10461,N_11876);
xor U14579 (N_14579,N_10788,N_12137);
or U14580 (N_14580,N_12395,N_11151);
xnor U14581 (N_14581,N_10766,N_10194);
xor U14582 (N_14582,N_11223,N_10919);
or U14583 (N_14583,N_12065,N_11247);
nor U14584 (N_14584,N_11984,N_10979);
nand U14585 (N_14585,N_12427,N_11574);
xnor U14586 (N_14586,N_12260,N_11067);
and U14587 (N_14587,N_10663,N_11019);
nand U14588 (N_14588,N_10296,N_11444);
or U14589 (N_14589,N_11083,N_11938);
and U14590 (N_14590,N_10244,N_11977);
nand U14591 (N_14591,N_10263,N_10220);
nand U14592 (N_14592,N_10503,N_12213);
and U14593 (N_14593,N_11419,N_11322);
or U14594 (N_14594,N_10608,N_12039);
nor U14595 (N_14595,N_10969,N_11390);
nor U14596 (N_14596,N_10726,N_11686);
and U14597 (N_14597,N_10536,N_10228);
nand U14598 (N_14598,N_11739,N_10012);
and U14599 (N_14599,N_10985,N_10658);
nor U14600 (N_14600,N_11249,N_10745);
or U14601 (N_14601,N_12197,N_11854);
or U14602 (N_14602,N_12139,N_12202);
and U14603 (N_14603,N_11133,N_11959);
or U14604 (N_14604,N_10049,N_11492);
or U14605 (N_14605,N_11218,N_10879);
nor U14606 (N_14606,N_10362,N_11216);
xnor U14607 (N_14607,N_11780,N_11394);
xor U14608 (N_14608,N_11381,N_11033);
nor U14609 (N_14609,N_12233,N_10479);
xnor U14610 (N_14610,N_12387,N_12013);
nor U14611 (N_14611,N_10396,N_10846);
xor U14612 (N_14612,N_12456,N_10260);
nand U14613 (N_14613,N_12136,N_11090);
nor U14614 (N_14614,N_12337,N_11173);
or U14615 (N_14615,N_10564,N_11903);
nand U14616 (N_14616,N_10657,N_10977);
xnor U14617 (N_14617,N_11075,N_11658);
nand U14618 (N_14618,N_10319,N_11659);
xnor U14619 (N_14619,N_10545,N_10292);
xor U14620 (N_14620,N_10899,N_12166);
nor U14621 (N_14621,N_12442,N_10249);
nor U14622 (N_14622,N_11087,N_10503);
xnor U14623 (N_14623,N_10034,N_11031);
xnor U14624 (N_14624,N_10295,N_11486);
or U14625 (N_14625,N_12214,N_10692);
xnor U14626 (N_14626,N_12462,N_12438);
nor U14627 (N_14627,N_10589,N_11831);
nand U14628 (N_14628,N_11788,N_12128);
or U14629 (N_14629,N_10625,N_11191);
or U14630 (N_14630,N_10363,N_10214);
xor U14631 (N_14631,N_10450,N_11158);
or U14632 (N_14632,N_11484,N_11449);
xnor U14633 (N_14633,N_10833,N_10203);
or U14634 (N_14634,N_11852,N_10261);
and U14635 (N_14635,N_10310,N_10067);
xor U14636 (N_14636,N_11196,N_11808);
nor U14637 (N_14637,N_11967,N_10057);
or U14638 (N_14638,N_10788,N_10964);
nor U14639 (N_14639,N_11817,N_12438);
xor U14640 (N_14640,N_10987,N_10226);
and U14641 (N_14641,N_12124,N_10128);
nand U14642 (N_14642,N_11690,N_12051);
nand U14643 (N_14643,N_12493,N_10171);
nor U14644 (N_14644,N_10152,N_11931);
and U14645 (N_14645,N_10774,N_10555);
xor U14646 (N_14646,N_10108,N_12232);
nor U14647 (N_14647,N_12035,N_12339);
xor U14648 (N_14648,N_11851,N_10519);
nor U14649 (N_14649,N_11314,N_10564);
nor U14650 (N_14650,N_12163,N_11378);
xor U14651 (N_14651,N_10486,N_10196);
and U14652 (N_14652,N_11230,N_11598);
xnor U14653 (N_14653,N_11185,N_12295);
nand U14654 (N_14654,N_12435,N_12269);
nand U14655 (N_14655,N_11681,N_11692);
nor U14656 (N_14656,N_11549,N_10072);
and U14657 (N_14657,N_11551,N_10101);
or U14658 (N_14658,N_10271,N_10389);
and U14659 (N_14659,N_11585,N_12113);
nand U14660 (N_14660,N_10939,N_10629);
xor U14661 (N_14661,N_11761,N_11052);
nand U14662 (N_14662,N_10507,N_11519);
xor U14663 (N_14663,N_11014,N_12173);
nor U14664 (N_14664,N_10833,N_12416);
nor U14665 (N_14665,N_10233,N_10867);
and U14666 (N_14666,N_12079,N_12385);
or U14667 (N_14667,N_10766,N_10733);
nand U14668 (N_14668,N_11019,N_11926);
and U14669 (N_14669,N_10058,N_10098);
and U14670 (N_14670,N_11653,N_10193);
and U14671 (N_14671,N_11598,N_11690);
nor U14672 (N_14672,N_10888,N_11649);
nor U14673 (N_14673,N_11427,N_10848);
or U14674 (N_14674,N_11611,N_11289);
and U14675 (N_14675,N_10849,N_10308);
or U14676 (N_14676,N_11583,N_10403);
nand U14677 (N_14677,N_11895,N_10344);
nor U14678 (N_14678,N_12162,N_12289);
and U14679 (N_14679,N_11298,N_12470);
nand U14680 (N_14680,N_11633,N_10330);
xnor U14681 (N_14681,N_12312,N_12112);
or U14682 (N_14682,N_10051,N_10804);
or U14683 (N_14683,N_10734,N_11170);
and U14684 (N_14684,N_12121,N_11012);
or U14685 (N_14685,N_11388,N_11585);
nor U14686 (N_14686,N_10389,N_10733);
or U14687 (N_14687,N_11540,N_12467);
or U14688 (N_14688,N_12186,N_10461);
xor U14689 (N_14689,N_10404,N_11178);
xor U14690 (N_14690,N_10790,N_11395);
nor U14691 (N_14691,N_12045,N_10079);
nand U14692 (N_14692,N_10815,N_11141);
nand U14693 (N_14693,N_11472,N_11239);
nor U14694 (N_14694,N_11660,N_11668);
nor U14695 (N_14695,N_11200,N_10109);
nand U14696 (N_14696,N_11253,N_10975);
nand U14697 (N_14697,N_12308,N_11241);
or U14698 (N_14698,N_10982,N_11739);
xnor U14699 (N_14699,N_11743,N_10793);
xor U14700 (N_14700,N_12474,N_11013);
and U14701 (N_14701,N_11882,N_10680);
or U14702 (N_14702,N_11678,N_11872);
or U14703 (N_14703,N_10884,N_11849);
xor U14704 (N_14704,N_11975,N_11934);
and U14705 (N_14705,N_12289,N_10973);
nor U14706 (N_14706,N_10511,N_10537);
and U14707 (N_14707,N_10601,N_12232);
or U14708 (N_14708,N_11650,N_10863);
xnor U14709 (N_14709,N_12134,N_11645);
and U14710 (N_14710,N_11756,N_12220);
nand U14711 (N_14711,N_11015,N_12346);
or U14712 (N_14712,N_10956,N_11369);
xor U14713 (N_14713,N_12021,N_11043);
nand U14714 (N_14714,N_11152,N_10755);
nand U14715 (N_14715,N_10808,N_10390);
nor U14716 (N_14716,N_10173,N_11328);
and U14717 (N_14717,N_10238,N_11172);
or U14718 (N_14718,N_10090,N_11942);
nand U14719 (N_14719,N_11683,N_12288);
nand U14720 (N_14720,N_11348,N_10133);
xor U14721 (N_14721,N_10070,N_10779);
and U14722 (N_14722,N_11161,N_11491);
nor U14723 (N_14723,N_10857,N_11531);
and U14724 (N_14724,N_11989,N_10580);
nor U14725 (N_14725,N_12112,N_12436);
xnor U14726 (N_14726,N_11473,N_11956);
xnor U14727 (N_14727,N_10174,N_10072);
xnor U14728 (N_14728,N_11051,N_11747);
nand U14729 (N_14729,N_11159,N_10227);
nor U14730 (N_14730,N_10878,N_10168);
or U14731 (N_14731,N_10286,N_10942);
xor U14732 (N_14732,N_10435,N_11479);
or U14733 (N_14733,N_11628,N_11395);
xor U14734 (N_14734,N_10477,N_10795);
nand U14735 (N_14735,N_11603,N_12280);
nand U14736 (N_14736,N_12247,N_11924);
xor U14737 (N_14737,N_11501,N_10320);
and U14738 (N_14738,N_12029,N_11869);
xnor U14739 (N_14739,N_11100,N_11612);
xnor U14740 (N_14740,N_12465,N_12128);
nand U14741 (N_14741,N_11738,N_11314);
xnor U14742 (N_14742,N_12402,N_10251);
nand U14743 (N_14743,N_10222,N_10091);
nor U14744 (N_14744,N_10096,N_10779);
and U14745 (N_14745,N_10691,N_10560);
or U14746 (N_14746,N_12190,N_11096);
or U14747 (N_14747,N_11684,N_11727);
xnor U14748 (N_14748,N_10928,N_11354);
nand U14749 (N_14749,N_11707,N_10514);
xnor U14750 (N_14750,N_10639,N_12123);
nand U14751 (N_14751,N_11670,N_10341);
and U14752 (N_14752,N_10044,N_11743);
xor U14753 (N_14753,N_10998,N_10692);
nor U14754 (N_14754,N_12456,N_11244);
or U14755 (N_14755,N_11685,N_10059);
xor U14756 (N_14756,N_10793,N_11378);
nor U14757 (N_14757,N_10275,N_11902);
nand U14758 (N_14758,N_10446,N_10128);
nand U14759 (N_14759,N_11657,N_12240);
nand U14760 (N_14760,N_10588,N_11560);
and U14761 (N_14761,N_11810,N_10074);
and U14762 (N_14762,N_10522,N_11247);
or U14763 (N_14763,N_11047,N_11310);
nand U14764 (N_14764,N_12126,N_11282);
and U14765 (N_14765,N_11016,N_11539);
and U14766 (N_14766,N_10221,N_10330);
nand U14767 (N_14767,N_10327,N_12299);
and U14768 (N_14768,N_11960,N_10655);
and U14769 (N_14769,N_10669,N_11778);
or U14770 (N_14770,N_12125,N_11860);
xnor U14771 (N_14771,N_10104,N_10712);
and U14772 (N_14772,N_12150,N_10074);
nand U14773 (N_14773,N_12276,N_11671);
nand U14774 (N_14774,N_11608,N_10755);
and U14775 (N_14775,N_11861,N_10575);
nand U14776 (N_14776,N_12259,N_12234);
and U14777 (N_14777,N_11042,N_10294);
nand U14778 (N_14778,N_10425,N_10667);
xnor U14779 (N_14779,N_12388,N_11702);
nand U14780 (N_14780,N_12402,N_10654);
xnor U14781 (N_14781,N_10164,N_11834);
or U14782 (N_14782,N_12488,N_10958);
xnor U14783 (N_14783,N_10944,N_10209);
nor U14784 (N_14784,N_12338,N_11219);
nor U14785 (N_14785,N_12090,N_11250);
nor U14786 (N_14786,N_10280,N_10032);
xor U14787 (N_14787,N_11013,N_12169);
nor U14788 (N_14788,N_12225,N_11817);
and U14789 (N_14789,N_11569,N_12356);
nor U14790 (N_14790,N_12105,N_10242);
nor U14791 (N_14791,N_12176,N_12238);
nor U14792 (N_14792,N_11602,N_10062);
nand U14793 (N_14793,N_10561,N_10317);
xnor U14794 (N_14794,N_11896,N_11709);
nor U14795 (N_14795,N_10038,N_11228);
xor U14796 (N_14796,N_10356,N_11667);
nor U14797 (N_14797,N_10115,N_12131);
nor U14798 (N_14798,N_10056,N_11283);
xnor U14799 (N_14799,N_11248,N_12122);
xor U14800 (N_14800,N_10381,N_10332);
and U14801 (N_14801,N_10038,N_10560);
nand U14802 (N_14802,N_10422,N_10465);
xnor U14803 (N_14803,N_10356,N_11520);
xnor U14804 (N_14804,N_11685,N_12226);
nand U14805 (N_14805,N_10071,N_10479);
and U14806 (N_14806,N_10833,N_12105);
nor U14807 (N_14807,N_10437,N_10012);
nor U14808 (N_14808,N_10216,N_11835);
xnor U14809 (N_14809,N_11204,N_12220);
or U14810 (N_14810,N_11286,N_11969);
nor U14811 (N_14811,N_12134,N_11699);
nand U14812 (N_14812,N_11311,N_10244);
xor U14813 (N_14813,N_11591,N_12356);
or U14814 (N_14814,N_12117,N_10035);
xor U14815 (N_14815,N_10638,N_11470);
xor U14816 (N_14816,N_10712,N_11286);
nand U14817 (N_14817,N_10276,N_10280);
nor U14818 (N_14818,N_11588,N_10312);
or U14819 (N_14819,N_10027,N_11118);
nand U14820 (N_14820,N_12106,N_11012);
and U14821 (N_14821,N_11426,N_10134);
or U14822 (N_14822,N_11116,N_12052);
nand U14823 (N_14823,N_11843,N_10703);
nor U14824 (N_14824,N_12460,N_10836);
or U14825 (N_14825,N_12340,N_10798);
xor U14826 (N_14826,N_11770,N_12393);
xor U14827 (N_14827,N_12152,N_11736);
or U14828 (N_14828,N_12141,N_11032);
xnor U14829 (N_14829,N_11168,N_11876);
nand U14830 (N_14830,N_10287,N_11585);
or U14831 (N_14831,N_10626,N_12054);
nand U14832 (N_14832,N_11966,N_12182);
nand U14833 (N_14833,N_12347,N_10687);
xor U14834 (N_14834,N_12076,N_10529);
nand U14835 (N_14835,N_10758,N_11410);
xor U14836 (N_14836,N_11235,N_10401);
nor U14837 (N_14837,N_10822,N_12201);
nor U14838 (N_14838,N_10647,N_11777);
nor U14839 (N_14839,N_10343,N_10415);
and U14840 (N_14840,N_11242,N_10154);
or U14841 (N_14841,N_10542,N_11720);
nand U14842 (N_14842,N_12314,N_12194);
xor U14843 (N_14843,N_10517,N_12413);
nand U14844 (N_14844,N_11971,N_10519);
and U14845 (N_14845,N_10291,N_11981);
or U14846 (N_14846,N_10612,N_11683);
nor U14847 (N_14847,N_12455,N_11522);
or U14848 (N_14848,N_11521,N_10088);
or U14849 (N_14849,N_11010,N_12308);
nand U14850 (N_14850,N_11267,N_11134);
nor U14851 (N_14851,N_12101,N_11870);
and U14852 (N_14852,N_10935,N_12257);
and U14853 (N_14853,N_10220,N_12087);
nand U14854 (N_14854,N_10817,N_10047);
xnor U14855 (N_14855,N_11515,N_12019);
or U14856 (N_14856,N_10784,N_10954);
nor U14857 (N_14857,N_10180,N_11305);
nor U14858 (N_14858,N_11971,N_10335);
nor U14859 (N_14859,N_11326,N_10804);
and U14860 (N_14860,N_10900,N_11606);
nand U14861 (N_14861,N_11862,N_11036);
or U14862 (N_14862,N_12171,N_10471);
nor U14863 (N_14863,N_10612,N_10701);
nor U14864 (N_14864,N_10149,N_10538);
nand U14865 (N_14865,N_10516,N_10717);
nor U14866 (N_14866,N_12091,N_10705);
nor U14867 (N_14867,N_10532,N_12238);
nor U14868 (N_14868,N_12371,N_11542);
and U14869 (N_14869,N_11974,N_11185);
nor U14870 (N_14870,N_11789,N_11767);
or U14871 (N_14871,N_10461,N_11322);
nor U14872 (N_14872,N_10697,N_10999);
nand U14873 (N_14873,N_10946,N_10226);
xor U14874 (N_14874,N_11371,N_10586);
xnor U14875 (N_14875,N_11878,N_10368);
and U14876 (N_14876,N_12301,N_12209);
nand U14877 (N_14877,N_11047,N_10807);
and U14878 (N_14878,N_10382,N_12292);
or U14879 (N_14879,N_11724,N_11154);
nor U14880 (N_14880,N_10675,N_11742);
and U14881 (N_14881,N_10547,N_11051);
or U14882 (N_14882,N_10964,N_12100);
nor U14883 (N_14883,N_10932,N_11064);
or U14884 (N_14884,N_10802,N_11847);
nor U14885 (N_14885,N_11864,N_10164);
nand U14886 (N_14886,N_12159,N_10533);
xnor U14887 (N_14887,N_11007,N_10391);
nand U14888 (N_14888,N_11217,N_12103);
nand U14889 (N_14889,N_10483,N_11504);
or U14890 (N_14890,N_12353,N_11860);
or U14891 (N_14891,N_11584,N_12427);
and U14892 (N_14892,N_12028,N_10642);
and U14893 (N_14893,N_11385,N_11593);
xor U14894 (N_14894,N_10666,N_11565);
xor U14895 (N_14895,N_10354,N_10619);
or U14896 (N_14896,N_10579,N_11234);
and U14897 (N_14897,N_12496,N_11524);
nor U14898 (N_14898,N_12257,N_10908);
nand U14899 (N_14899,N_12000,N_12219);
xnor U14900 (N_14900,N_10503,N_12033);
or U14901 (N_14901,N_12108,N_10023);
and U14902 (N_14902,N_10521,N_10541);
or U14903 (N_14903,N_12441,N_10740);
xnor U14904 (N_14904,N_12092,N_10099);
and U14905 (N_14905,N_10495,N_11541);
and U14906 (N_14906,N_11691,N_10447);
or U14907 (N_14907,N_12143,N_10316);
and U14908 (N_14908,N_10753,N_11010);
nand U14909 (N_14909,N_10975,N_10173);
and U14910 (N_14910,N_10470,N_11061);
or U14911 (N_14911,N_10597,N_11276);
xor U14912 (N_14912,N_12030,N_11762);
nor U14913 (N_14913,N_12413,N_10064);
xor U14914 (N_14914,N_12462,N_10525);
nor U14915 (N_14915,N_10292,N_10653);
nand U14916 (N_14916,N_11948,N_12098);
or U14917 (N_14917,N_11053,N_12117);
and U14918 (N_14918,N_11191,N_12329);
xor U14919 (N_14919,N_12145,N_10247);
nor U14920 (N_14920,N_10126,N_11529);
or U14921 (N_14921,N_10920,N_12369);
and U14922 (N_14922,N_12335,N_11582);
nand U14923 (N_14923,N_10524,N_10424);
or U14924 (N_14924,N_10157,N_10234);
or U14925 (N_14925,N_12155,N_11952);
and U14926 (N_14926,N_11968,N_10087);
and U14927 (N_14927,N_10455,N_11176);
nor U14928 (N_14928,N_10102,N_10701);
xnor U14929 (N_14929,N_11461,N_10284);
nand U14930 (N_14930,N_10239,N_10942);
nor U14931 (N_14931,N_10434,N_10295);
or U14932 (N_14932,N_10666,N_10634);
and U14933 (N_14933,N_11700,N_10141);
nand U14934 (N_14934,N_12386,N_12349);
or U14935 (N_14935,N_10554,N_11868);
xnor U14936 (N_14936,N_12414,N_11753);
nor U14937 (N_14937,N_11810,N_12053);
or U14938 (N_14938,N_10087,N_10199);
or U14939 (N_14939,N_10420,N_10445);
or U14940 (N_14940,N_10867,N_12420);
and U14941 (N_14941,N_11994,N_11269);
xor U14942 (N_14942,N_11978,N_10359);
xnor U14943 (N_14943,N_12027,N_12082);
nor U14944 (N_14944,N_10748,N_10596);
nand U14945 (N_14945,N_12302,N_10174);
nand U14946 (N_14946,N_12323,N_11541);
nor U14947 (N_14947,N_11951,N_10161);
and U14948 (N_14948,N_10792,N_10852);
and U14949 (N_14949,N_10488,N_10158);
xor U14950 (N_14950,N_11926,N_10271);
nand U14951 (N_14951,N_12130,N_12338);
or U14952 (N_14952,N_11028,N_12142);
or U14953 (N_14953,N_10327,N_10699);
xnor U14954 (N_14954,N_10464,N_11785);
or U14955 (N_14955,N_10704,N_10157);
nand U14956 (N_14956,N_12382,N_10663);
and U14957 (N_14957,N_10213,N_10509);
xor U14958 (N_14958,N_10047,N_11746);
or U14959 (N_14959,N_10365,N_11058);
xor U14960 (N_14960,N_11412,N_12181);
and U14961 (N_14961,N_10086,N_11086);
xor U14962 (N_14962,N_10311,N_10983);
nor U14963 (N_14963,N_11385,N_10439);
nor U14964 (N_14964,N_11126,N_10896);
nor U14965 (N_14965,N_11543,N_10585);
xor U14966 (N_14966,N_11849,N_10802);
nor U14967 (N_14967,N_11971,N_11805);
xor U14968 (N_14968,N_11990,N_10160);
xnor U14969 (N_14969,N_11217,N_11112);
or U14970 (N_14970,N_10505,N_10374);
nand U14971 (N_14971,N_11993,N_10296);
xnor U14972 (N_14972,N_11821,N_12308);
nor U14973 (N_14973,N_11423,N_11765);
xnor U14974 (N_14974,N_11997,N_12290);
nand U14975 (N_14975,N_11704,N_10842);
nand U14976 (N_14976,N_12022,N_10509);
xor U14977 (N_14977,N_10359,N_11855);
and U14978 (N_14978,N_12163,N_11911);
nand U14979 (N_14979,N_11799,N_10217);
xnor U14980 (N_14980,N_12440,N_12125);
or U14981 (N_14981,N_11435,N_10398);
xnor U14982 (N_14982,N_10599,N_11429);
xor U14983 (N_14983,N_11759,N_12176);
xnor U14984 (N_14984,N_10883,N_10695);
nand U14985 (N_14985,N_10443,N_11671);
nor U14986 (N_14986,N_12239,N_10070);
xor U14987 (N_14987,N_10957,N_10580);
xor U14988 (N_14988,N_11190,N_10306);
nand U14989 (N_14989,N_12427,N_10701);
nor U14990 (N_14990,N_11417,N_11849);
nor U14991 (N_14991,N_11875,N_10069);
nor U14992 (N_14992,N_11577,N_10660);
nand U14993 (N_14993,N_11889,N_11659);
xnor U14994 (N_14994,N_10759,N_11625);
nor U14995 (N_14995,N_11809,N_10983);
xnor U14996 (N_14996,N_10148,N_11135);
nand U14997 (N_14997,N_12246,N_11190);
or U14998 (N_14998,N_12478,N_10620);
and U14999 (N_14999,N_10477,N_12040);
nor U15000 (N_15000,N_14994,N_12856);
nor U15001 (N_15001,N_14719,N_14833);
xnor U15002 (N_15002,N_12823,N_12527);
nand U15003 (N_15003,N_14393,N_13021);
and U15004 (N_15004,N_13224,N_14985);
nand U15005 (N_15005,N_13691,N_13813);
and U15006 (N_15006,N_12940,N_13930);
or U15007 (N_15007,N_12928,N_13085);
nand U15008 (N_15008,N_12529,N_12615);
nand U15009 (N_15009,N_14845,N_13336);
xor U15010 (N_15010,N_14356,N_12715);
or U15011 (N_15011,N_14226,N_14924);
nor U15012 (N_15012,N_13090,N_12510);
nand U15013 (N_15013,N_14756,N_14515);
or U15014 (N_15014,N_12848,N_13402);
nand U15015 (N_15015,N_13810,N_14647);
nand U15016 (N_15016,N_13095,N_12950);
or U15017 (N_15017,N_14496,N_14714);
nor U15018 (N_15018,N_12839,N_14025);
and U15019 (N_15019,N_12607,N_14904);
xnor U15020 (N_15020,N_13972,N_14355);
nor U15021 (N_15021,N_14630,N_14807);
or U15022 (N_15022,N_13586,N_14029);
and U15023 (N_15023,N_13400,N_14530);
nand U15024 (N_15024,N_12891,N_14000);
nor U15025 (N_15025,N_14829,N_12968);
nor U15026 (N_15026,N_14235,N_13220);
and U15027 (N_15027,N_14342,N_14949);
and U15028 (N_15028,N_13709,N_14230);
nor U15029 (N_15029,N_12994,N_13771);
xnor U15030 (N_15030,N_13523,N_13701);
and U15031 (N_15031,N_13991,N_14576);
nand U15032 (N_15032,N_14173,N_14425);
or U15033 (N_15033,N_12555,N_14652);
nand U15034 (N_15034,N_13529,N_14586);
nor U15035 (N_15035,N_13971,N_13654);
or U15036 (N_15036,N_13260,N_12820);
nor U15037 (N_15037,N_13038,N_14684);
or U15038 (N_15038,N_14916,N_14264);
xnor U15039 (N_15039,N_12772,N_14600);
or U15040 (N_15040,N_14497,N_14942);
or U15041 (N_15041,N_13221,N_13712);
nand U15042 (N_15042,N_13665,N_13408);
and U15043 (N_15043,N_12631,N_14955);
nand U15044 (N_15044,N_13913,N_13265);
and U15045 (N_15045,N_14039,N_12806);
nor U15046 (N_15046,N_13576,N_12796);
nor U15047 (N_15047,N_14122,N_14022);
nand U15048 (N_15048,N_13753,N_12824);
nand U15049 (N_15049,N_14943,N_14086);
or U15050 (N_15050,N_13750,N_14941);
xor U15051 (N_15051,N_14298,N_12870);
nor U15052 (N_15052,N_14844,N_14294);
nand U15053 (N_15053,N_14604,N_12539);
or U15054 (N_15054,N_14927,N_14796);
and U15055 (N_15055,N_13908,N_14026);
and U15056 (N_15056,N_12732,N_13087);
xnor U15057 (N_15057,N_14933,N_12846);
xnor U15058 (N_15058,N_13911,N_14021);
nor U15059 (N_15059,N_14953,N_14826);
or U15060 (N_15060,N_14477,N_13205);
nor U15061 (N_15061,N_12504,N_14655);
nor U15062 (N_15062,N_14893,N_13724);
nor U15063 (N_15063,N_14096,N_12654);
xnor U15064 (N_15064,N_12567,N_14510);
nor U15065 (N_15065,N_12557,N_14853);
and U15066 (N_15066,N_14241,N_13793);
and U15067 (N_15067,N_12652,N_13189);
xnor U15068 (N_15068,N_14367,N_13927);
xnor U15069 (N_15069,N_14403,N_13332);
nand U15070 (N_15070,N_12590,N_13309);
or U15071 (N_15071,N_14897,N_14248);
or U15072 (N_15072,N_14143,N_13326);
or U15073 (N_15073,N_14782,N_13497);
nor U15074 (N_15074,N_13985,N_14761);
or U15075 (N_15075,N_14675,N_14921);
or U15076 (N_15076,N_14704,N_14649);
and U15077 (N_15077,N_13975,N_12955);
xnor U15078 (N_15078,N_12503,N_14887);
nand U15079 (N_15079,N_13471,N_13277);
nand U15080 (N_15080,N_13577,N_13213);
xor U15081 (N_15081,N_14349,N_14598);
or U15082 (N_15082,N_14240,N_14204);
xnor U15083 (N_15083,N_14323,N_14607);
nor U15084 (N_15084,N_12574,N_12711);
or U15085 (N_15085,N_12973,N_14773);
nor U15086 (N_15086,N_14854,N_13510);
nor U15087 (N_15087,N_14163,N_13998);
or U15088 (N_15088,N_14488,N_13001);
and U15089 (N_15089,N_13934,N_12939);
nor U15090 (N_15090,N_14547,N_14485);
or U15091 (N_15091,N_13686,N_13433);
xnor U15092 (N_15092,N_14307,N_12530);
and U15093 (N_15093,N_13719,N_14035);
or U15094 (N_15094,N_14744,N_12683);
or U15095 (N_15095,N_12502,N_13063);
nor U15096 (N_15096,N_12730,N_14005);
or U15097 (N_15097,N_13940,N_13769);
nor U15098 (N_15098,N_13043,N_12680);
nand U15099 (N_15099,N_13049,N_12752);
or U15100 (N_15100,N_14622,N_14841);
and U15101 (N_15101,N_12507,N_12565);
nand U15102 (N_15102,N_14691,N_12674);
nor U15103 (N_15103,N_13776,N_14302);
or U15104 (N_15104,N_13535,N_14753);
nor U15105 (N_15105,N_12884,N_13052);
xor U15106 (N_15106,N_13589,N_14666);
nand U15107 (N_15107,N_14717,N_13821);
nor U15108 (N_15108,N_14708,N_12627);
or U15109 (N_15109,N_13811,N_14973);
nor U15110 (N_15110,N_14919,N_12873);
nand U15111 (N_15111,N_14366,N_14179);
and U15112 (N_15112,N_12681,N_14257);
xor U15113 (N_15113,N_13734,N_14350);
or U15114 (N_15114,N_14615,N_13391);
xor U15115 (N_15115,N_12923,N_13136);
nor U15116 (N_15116,N_13680,N_12748);
nor U15117 (N_15117,N_14238,N_13430);
xnor U15118 (N_15118,N_13415,N_12999);
nand U15119 (N_15119,N_12841,N_14839);
or U15120 (N_15120,N_12943,N_14289);
or U15121 (N_15121,N_13289,N_13527);
or U15122 (N_15122,N_14764,N_13852);
or U15123 (N_15123,N_13375,N_14890);
or U15124 (N_15124,N_14428,N_14514);
xnor U15125 (N_15125,N_14269,N_13357);
nand U15126 (N_15126,N_13915,N_14260);
xor U15127 (N_15127,N_13212,N_14336);
nand U15128 (N_15128,N_14068,N_14244);
or U15129 (N_15129,N_12633,N_12785);
xnor U15130 (N_15130,N_13693,N_14653);
nand U15131 (N_15131,N_14929,N_14676);
nand U15132 (N_15132,N_14690,N_13636);
nand U15133 (N_15133,N_13106,N_13174);
and U15134 (N_15134,N_12684,N_14692);
nand U15135 (N_15135,N_14505,N_14164);
nor U15136 (N_15136,N_12626,N_13086);
xor U15137 (N_15137,N_12718,N_14175);
nand U15138 (N_15138,N_13105,N_13468);
nand U15139 (N_15139,N_13301,N_14781);
nor U15140 (N_15140,N_12546,N_13949);
nand U15141 (N_15141,N_13083,N_12519);
and U15142 (N_15142,N_14406,N_13483);
xor U15143 (N_15143,N_13002,N_12724);
and U15144 (N_15144,N_14037,N_13879);
and U15145 (N_15145,N_13306,N_13302);
xnor U15146 (N_15146,N_12704,N_14689);
and U15147 (N_15147,N_12746,N_14007);
xnor U15148 (N_15148,N_14376,N_12723);
xnor U15149 (N_15149,N_12855,N_13980);
nor U15150 (N_15150,N_12659,N_12564);
nand U15151 (N_15151,N_14458,N_13854);
and U15152 (N_15152,N_13466,N_14042);
xor U15153 (N_15153,N_12766,N_13373);
nor U15154 (N_15154,N_13275,N_14011);
nor U15155 (N_15155,N_14256,N_12887);
nor U15156 (N_15156,N_14389,N_13524);
nand U15157 (N_15157,N_14354,N_12528);
nor U15158 (N_15158,N_12805,N_13041);
nor U15159 (N_15159,N_13084,N_14337);
and U15160 (N_15160,N_13969,N_14283);
or U15161 (N_15161,N_14906,N_12997);
xnor U15162 (N_15162,N_13649,N_14662);
nand U15163 (N_15163,N_14492,N_13469);
nor U15164 (N_15164,N_14987,N_12743);
nand U15165 (N_15165,N_14566,N_12614);
xnor U15166 (N_15166,N_14540,N_12538);
and U15167 (N_15167,N_13185,N_13531);
xnor U15168 (N_15168,N_12547,N_13592);
nor U15169 (N_15169,N_12902,N_13961);
or U15170 (N_15170,N_13801,N_13023);
or U15171 (N_15171,N_13842,N_12798);
or U15172 (N_15172,N_13739,N_14110);
nand U15173 (N_15173,N_13723,N_14718);
xor U15174 (N_15174,N_13008,N_14185);
or U15175 (N_15175,N_13175,N_13595);
nor U15176 (N_15176,N_14080,N_13441);
and U15177 (N_15177,N_13792,N_13662);
nor U15178 (N_15178,N_14333,N_13034);
xor U15179 (N_15179,N_14539,N_12535);
or U15180 (N_15180,N_12998,N_14100);
or U15181 (N_15181,N_14693,N_13903);
nor U15182 (N_15182,N_12906,N_13760);
and U15183 (N_15183,N_14413,N_14819);
and U15184 (N_15184,N_14528,N_14963);
xor U15185 (N_15185,N_12981,N_12882);
nand U15186 (N_15186,N_13905,N_12991);
nand U15187 (N_15187,N_14557,N_13024);
and U15188 (N_15188,N_12886,N_12864);
nand U15189 (N_15189,N_12740,N_12677);
or U15190 (N_15190,N_14707,N_13569);
and U15191 (N_15191,N_13485,N_12531);
xor U15192 (N_15192,N_13138,N_14884);
xor U15193 (N_15193,N_13543,N_12582);
xnor U15194 (N_15194,N_14448,N_13278);
nor U15195 (N_15195,N_14688,N_14951);
nand U15196 (N_15196,N_14135,N_14888);
or U15197 (N_15197,N_14797,N_14755);
xor U15198 (N_15198,N_14316,N_14410);
nor U15199 (N_15199,N_13887,N_13928);
or U15200 (N_15200,N_12753,N_14745);
or U15201 (N_15201,N_12523,N_14751);
or U15202 (N_15202,N_12642,N_14587);
xnor U15203 (N_15203,N_13360,N_13959);
xor U15204 (N_15204,N_14741,N_12733);
nor U15205 (N_15205,N_13721,N_14585);
and U15206 (N_15206,N_14031,N_12990);
xnor U15207 (N_15207,N_13380,N_12629);
xnor U15208 (N_15208,N_14222,N_12602);
nand U15209 (N_15209,N_14049,N_14338);
xor U15210 (N_15210,N_13057,N_13465);
xnor U15211 (N_15211,N_13230,N_12901);
and U15212 (N_15212,N_14267,N_14960);
and U15213 (N_15213,N_12959,N_14468);
nand U15214 (N_15214,N_13005,N_13440);
nor U15215 (N_15215,N_13267,N_13239);
nand U15216 (N_15216,N_13544,N_14093);
or U15217 (N_15217,N_12726,N_13727);
and U15218 (N_15218,N_13645,N_12657);
xor U15219 (N_15219,N_14397,N_13997);
or U15220 (N_15220,N_14142,N_12930);
nand U15221 (N_15221,N_13575,N_12645);
and U15222 (N_15222,N_13520,N_14044);
and U15223 (N_15223,N_13939,N_14885);
xnor U15224 (N_15224,N_12764,N_14003);
nand U15225 (N_15225,N_13486,N_14332);
xnor U15226 (N_15226,N_13037,N_13525);
or U15227 (N_15227,N_12616,N_12637);
nand U15228 (N_15228,N_13366,N_13258);
and U15229 (N_15229,N_13778,N_14721);
nor U15230 (N_15230,N_14494,N_13066);
and U15231 (N_15231,N_14407,N_14117);
or U15232 (N_15232,N_13226,N_14936);
nand U15233 (N_15233,N_13707,N_13682);
nand U15234 (N_15234,N_14119,N_13588);
nand U15235 (N_15235,N_14495,N_14720);
or U15236 (N_15236,N_14664,N_13603);
or U15237 (N_15237,N_13386,N_12697);
and U15238 (N_15238,N_12777,N_14131);
nand U15239 (N_15239,N_13533,N_12807);
nor U15240 (N_15240,N_13312,N_12918);
and U15241 (N_15241,N_14896,N_13015);
xnor U15242 (N_15242,N_14475,N_14006);
xnor U15243 (N_15243,N_14192,N_13947);
and U15244 (N_15244,N_14161,N_14578);
xnor U15245 (N_15245,N_12541,N_13341);
or U15246 (N_15246,N_13599,N_13072);
xor U15247 (N_15247,N_13206,N_14501);
xor U15248 (N_15248,N_14372,N_13722);
or U15249 (N_15249,N_12812,N_14078);
xor U15250 (N_15250,N_13866,N_13029);
and U15251 (N_15251,N_13736,N_14836);
xnor U15252 (N_15252,N_13574,N_14864);
or U15253 (N_15253,N_12983,N_14616);
or U15254 (N_15254,N_14415,N_14591);
or U15255 (N_15255,N_12641,N_14137);
xnor U15256 (N_15256,N_12580,N_14082);
xnor U15257 (N_15257,N_12869,N_14292);
nor U15258 (N_15258,N_14816,N_14127);
and U15259 (N_15259,N_12861,N_13200);
nand U15260 (N_15260,N_13818,N_14926);
nand U15261 (N_15261,N_12854,N_13297);
nor U15262 (N_15262,N_14373,N_12670);
xor U15263 (N_15263,N_14212,N_13229);
or U15264 (N_15264,N_14463,N_14878);
nand U15265 (N_15265,N_14304,N_12653);
nor U15266 (N_15266,N_13847,N_14196);
nand U15267 (N_15267,N_14777,N_13618);
or U15268 (N_15268,N_13311,N_13428);
and U15269 (N_15269,N_12713,N_13246);
nor U15270 (N_15270,N_14038,N_14958);
and U15271 (N_15271,N_12679,N_12905);
or U15272 (N_15272,N_13236,N_13113);
nand U15273 (N_15273,N_13773,N_13878);
nand U15274 (N_15274,N_13704,N_13473);
nor U15275 (N_15275,N_14787,N_13581);
or U15276 (N_15276,N_13674,N_14420);
and U15277 (N_15277,N_14908,N_14780);
or U15278 (N_15278,N_14903,N_14382);
xnor U15279 (N_15279,N_13796,N_13101);
nand U15280 (N_15280,N_13832,N_14710);
nor U15281 (N_15281,N_13917,N_14606);
or U15282 (N_15282,N_13914,N_13779);
or U15283 (N_15283,N_14476,N_14141);
xnor U15284 (N_15284,N_13857,N_13684);
nand U15285 (N_15285,N_14380,N_12736);
nor U15286 (N_15286,N_13899,N_14032);
xnor U15287 (N_15287,N_13337,N_14132);
nand U15288 (N_15288,N_14627,N_13742);
nand U15289 (N_15289,N_12673,N_14769);
and U15290 (N_15290,N_12868,N_13597);
and U15291 (N_15291,N_13952,N_14057);
xnor U15292 (N_15292,N_14983,N_13885);
nand U15293 (N_15293,N_13308,N_14219);
nor U15294 (N_15294,N_13183,N_14459);
xor U15295 (N_15295,N_13192,N_14015);
nand U15296 (N_15296,N_12517,N_12857);
nor U15297 (N_15297,N_13300,N_14984);
and U15298 (N_15298,N_14147,N_14259);
xor U15299 (N_15299,N_13827,N_13040);
nor U15300 (N_15300,N_14808,N_14368);
nand U15301 (N_15301,N_13780,N_12985);
nand U15302 (N_15302,N_14880,N_13694);
or U15303 (N_15303,N_14687,N_13137);
xor U15304 (N_15304,N_14315,N_13889);
and U15305 (N_15305,N_13233,N_13439);
nor U15306 (N_15306,N_12791,N_13142);
or U15307 (N_15307,N_14545,N_13981);
nand U15308 (N_15308,N_14525,N_12871);
nand U15309 (N_15309,N_14213,N_12890);
nand U15310 (N_15310,N_13921,N_12953);
nand U15311 (N_15311,N_13255,N_13006);
nand U15312 (N_15312,N_12776,N_13369);
xor U15313 (N_15313,N_14109,N_13353);
xnor U15314 (N_15314,N_14399,N_13426);
xnor U15315 (N_15315,N_14568,N_13100);
or U15316 (N_15316,N_14471,N_14701);
or U15317 (N_15317,N_13075,N_12872);
nor U15318 (N_15318,N_13330,N_14450);
or U15319 (N_15319,N_13789,N_14931);
and U15320 (N_15320,N_13062,N_14329);
or U15321 (N_15321,N_13990,N_14305);
xor U15322 (N_15322,N_14043,N_13065);
or U15323 (N_15323,N_13240,N_13414);
nor U15324 (N_15324,N_14327,N_14104);
and U15325 (N_15325,N_13349,N_13831);
nand U15326 (N_15326,N_14867,N_14101);
nand U15327 (N_15327,N_14059,N_13663);
nand U15328 (N_15328,N_12979,N_13678);
nand U15329 (N_15329,N_12840,N_14064);
nor U15330 (N_15330,N_14861,N_14763);
nor U15331 (N_15331,N_14205,N_13070);
nor U15332 (N_15332,N_14883,N_13110);
xor U15333 (N_15333,N_14901,N_13896);
xor U15334 (N_15334,N_12501,N_14225);
or U15335 (N_15335,N_14703,N_13966);
and U15336 (N_15336,N_13288,N_13437);
nor U15337 (N_15337,N_13920,N_12795);
nand U15338 (N_15338,N_14200,N_14392);
nor U15339 (N_15339,N_14417,N_14309);
nand U15340 (N_15340,N_13319,N_14479);
or U15341 (N_15341,N_14094,N_13728);
nor U15342 (N_15342,N_14263,N_12600);
nand U15343 (N_15343,N_13248,N_14722);
nor U15344 (N_15344,N_14815,N_12588);
nand U15345 (N_15345,N_14866,N_12705);
nor U15346 (N_15346,N_13602,N_14732);
and U15347 (N_15347,N_14711,N_12698);
nor U15348 (N_15348,N_12608,N_13558);
or U15349 (N_15349,N_14277,N_13279);
xor U15350 (N_15350,N_13111,N_13823);
or U15351 (N_15351,N_12696,N_14818);
xnor U15352 (N_15352,N_13446,N_13315);
nor U15353 (N_15353,N_14930,N_13003);
nor U15354 (N_15354,N_13434,N_13685);
nor U15355 (N_15355,N_14430,N_12784);
nor U15356 (N_15356,N_13436,N_12500);
xnor U15357 (N_15357,N_14679,N_12989);
and U15358 (N_15358,N_14642,N_12957);
or U15359 (N_15359,N_14954,N_13898);
or U15360 (N_15360,N_13039,N_14462);
xor U15361 (N_15361,N_12945,N_12569);
or U15362 (N_15362,N_13303,N_13294);
nand U15363 (N_15363,N_13245,N_13390);
or U15364 (N_15364,N_13715,N_14293);
nor U15365 (N_15365,N_13763,N_14193);
xor U15366 (N_15366,N_12526,N_13667);
nand U15367 (N_15367,N_12621,N_12927);
xnor U15368 (N_15368,N_14651,N_14791);
nand U15369 (N_15369,N_13000,N_14534);
nor U15370 (N_15370,N_13634,N_14178);
xnor U15371 (N_15371,N_14922,N_13243);
xnor U15372 (N_15372,N_14895,N_13339);
nor U15373 (N_15373,N_14639,N_12908);
or U15374 (N_15374,N_13495,N_13676);
nor U15375 (N_15375,N_14577,N_12894);
and U15376 (N_15376,N_14014,N_14899);
xnor U15377 (N_15377,N_13545,N_14151);
or U15378 (N_15378,N_12553,N_14868);
nor U15379 (N_15379,N_13058,N_13091);
and U15380 (N_15380,N_14098,N_14736);
nand U15381 (N_15381,N_14195,N_13210);
xor U15382 (N_15382,N_14377,N_13050);
nand U15383 (N_15383,N_14451,N_12717);
or U15384 (N_15384,N_14234,N_14105);
and U15385 (N_15385,N_13004,N_14997);
and U15386 (N_15386,N_14437,N_14757);
and U15387 (N_15387,N_12536,N_13099);
nor U15388 (N_15388,N_13121,N_14498);
xnor U15389 (N_15389,N_13925,N_12606);
and U15390 (N_15390,N_14385,N_13860);
nor U15391 (N_15391,N_13347,N_13377);
or U15392 (N_15392,N_14776,N_14968);
or U15393 (N_15393,N_14275,N_12875);
nand U15394 (N_15394,N_14159,N_14258);
nand U15395 (N_15395,N_13241,N_13672);
xor U15396 (N_15396,N_13123,N_13026);
or U15397 (N_15397,N_12952,N_14171);
xor U15398 (N_15398,N_14920,N_14353);
xor U15399 (N_15399,N_12895,N_13389);
nand U15400 (N_15400,N_13167,N_13979);
nor U15401 (N_15401,N_14661,N_13276);
and U15402 (N_15402,N_14817,N_12768);
and U15403 (N_15403,N_14254,N_12663);
and U15404 (N_15404,N_14169,N_14176);
xnor U15405 (N_15405,N_13848,N_14249);
and U15406 (N_15406,N_12703,N_13195);
and U15407 (N_15407,N_13042,N_13398);
nor U15408 (N_15408,N_13625,N_13888);
nand U15409 (N_15409,N_13251,N_12549);
nand U15410 (N_15410,N_14313,N_14124);
xnor U15411 (N_15411,N_14500,N_13862);
xnor U15412 (N_15412,N_14830,N_13420);
nor U15413 (N_15413,N_13313,N_13064);
nor U15414 (N_15414,N_13141,N_14646);
nand U15415 (N_15415,N_13331,N_14482);
nor U15416 (N_15416,N_13269,N_13365);
nor U15417 (N_15417,N_12682,N_14474);
nand U15418 (N_15418,N_13350,N_14079);
or U15419 (N_15419,N_13153,N_14970);
or U15420 (N_15420,N_12562,N_12944);
and U15421 (N_15421,N_12623,N_13405);
nor U15422 (N_15422,N_14969,N_12809);
and U15423 (N_15423,N_14914,N_14966);
nand U15424 (N_15424,N_13444,N_13451);
xnor U15425 (N_15425,N_13295,N_13748);
xnor U15426 (N_15426,N_13782,N_12987);
or U15427 (N_15427,N_14971,N_13834);
nor U15428 (N_15428,N_12815,N_13361);
nand U15429 (N_15429,N_12699,N_14357);
nand U15430 (N_15430,N_14621,N_14848);
nand U15431 (N_15431,N_12646,N_14388);
xor U15432 (N_15432,N_14669,N_14593);
xnor U15433 (N_15433,N_13995,N_13968);
and U15434 (N_15434,N_14379,N_13479);
xor U15435 (N_15435,N_12971,N_13250);
xor U15436 (N_15436,N_13614,N_12594);
and U15437 (N_15437,N_12655,N_14558);
nand U15438 (N_15438,N_14282,N_14167);
nor U15439 (N_15439,N_14394,N_13808);
or U15440 (N_15440,N_12783,N_14972);
or U15441 (N_15441,N_14120,N_13035);
or U15442 (N_15442,N_14210,N_13619);
xor U15443 (N_15443,N_12584,N_13127);
nand U15444 (N_15444,N_14599,N_12694);
nand U15445 (N_15445,N_14567,N_14728);
nor U15446 (N_15446,N_14508,N_12767);
or U15447 (N_15447,N_14705,N_14582);
nor U15448 (N_15448,N_12756,N_13561);
nor U15449 (N_15449,N_13355,N_13957);
nor U15450 (N_15450,N_13125,N_13546);
and U15451 (N_15451,N_12545,N_13583);
nand U15452 (N_15452,N_14590,N_14231);
xnor U15453 (N_15453,N_12958,N_13081);
xnor U15454 (N_15454,N_12533,N_12758);
or U15455 (N_15455,N_14145,N_14416);
nand U15456 (N_15456,N_13648,N_13122);
nand U15457 (N_15457,N_14911,N_14838);
nor U15458 (N_15458,N_13978,N_13145);
or U15459 (N_15459,N_12822,N_14401);
and U15460 (N_15460,N_14659,N_14155);
or U15461 (N_15461,N_13600,N_13965);
nor U15462 (N_15462,N_12511,N_12542);
and U15463 (N_15463,N_13982,N_12914);
nand U15464 (N_15464,N_14207,N_13139);
nor U15465 (N_15465,N_14811,N_14150);
xnor U15466 (N_15466,N_14671,N_13011);
nor U15467 (N_15467,N_13162,N_14729);
or U15468 (N_15468,N_14414,N_12828);
nor U15469 (N_15469,N_13538,N_14760);
xor U15470 (N_15470,N_13815,N_12747);
and U15471 (N_15471,N_13673,N_13891);
nand U15472 (N_15472,N_14335,N_13788);
nand U15473 (N_15473,N_13573,N_13130);
and U15474 (N_15474,N_13179,N_12866);
and U15475 (N_15475,N_14735,N_14928);
and U15476 (N_15476,N_13872,N_13247);
or U15477 (N_15477,N_12825,N_13923);
nor U15478 (N_15478,N_13460,N_14330);
nand U15479 (N_15479,N_14674,N_12790);
or U15480 (N_15480,N_12937,N_12599);
or U15481 (N_15481,N_14945,N_13412);
and U15482 (N_15482,N_14873,N_13429);
xnor U15483 (N_15483,N_13653,N_14804);
nor U15484 (N_15484,N_14952,N_12816);
xnor U15485 (N_15485,N_13841,N_12597);
nor U15486 (N_15486,N_13629,N_14077);
nor U15487 (N_15487,N_12725,N_14694);
xnor U15488 (N_15488,N_13897,N_12662);
or U15489 (N_15489,N_14877,N_12716);
xnor U15490 (N_15490,N_13974,N_14976);
nor U15491 (N_15491,N_13633,N_14611);
and U15492 (N_15492,N_14865,N_12585);
nand U15493 (N_15493,N_13781,N_12676);
nor U15494 (N_15494,N_12892,N_13955);
or U15495 (N_15495,N_14803,N_14486);
nor U15496 (N_15496,N_13987,N_13421);
or U15497 (N_15497,N_13910,N_13655);
nand U15498 (N_15498,N_14734,N_13509);
nand U15499 (N_15499,N_14115,N_13967);
nor U15500 (N_15500,N_13354,N_14767);
xnor U15501 (N_15501,N_12829,N_14095);
or U15502 (N_15502,N_12803,N_13218);
nor U15503 (N_15503,N_12687,N_12577);
xor U15504 (N_15504,N_13364,N_12522);
nor U15505 (N_15505,N_13932,N_14834);
nand U15506 (N_15506,N_13334,N_13931);
or U15507 (N_15507,N_12802,N_13924);
nor U15508 (N_15508,N_14395,N_14056);
and U15509 (N_15509,N_12821,N_12850);
or U15510 (N_15510,N_13906,N_13790);
xnor U15511 (N_15511,N_12689,N_13342);
xnor U15512 (N_15512,N_13548,N_13314);
nand U15513 (N_15513,N_14871,N_12789);
and U15514 (N_15514,N_13016,N_13993);
nor U15515 (N_15515,N_13565,N_14114);
xnor U15516 (N_15516,N_12834,N_13596);
nand U15517 (N_15517,N_13092,N_13560);
xnor U15518 (N_15518,N_14431,N_12951);
or U15519 (N_15519,N_13150,N_12591);
nand U15520 (N_15520,N_12671,N_13956);
xnor U15521 (N_15521,N_14784,N_13962);
and U15522 (N_15522,N_14554,N_12786);
or U15523 (N_15523,N_12744,N_13953);
or U15524 (N_15524,N_13082,N_13103);
and U15525 (N_15525,N_14996,N_14010);
or U15526 (N_15526,N_13568,N_13710);
and U15527 (N_15527,N_14506,N_14683);
nand U15528 (N_15528,N_14438,N_12757);
and U15529 (N_15529,N_13746,N_14008);
and U15530 (N_15530,N_14365,N_14177);
or U15531 (N_15531,N_14940,N_12570);
nor U15532 (N_15532,N_14473,N_13608);
xnor U15533 (N_15533,N_13826,N_12978);
nand U15534 (N_15534,N_13147,N_13745);
and U15535 (N_15535,N_12853,N_14529);
and U15536 (N_15536,N_14184,N_13960);
nor U15537 (N_15537,N_13954,N_13472);
xnor U15538 (N_15538,N_14133,N_12508);
or U15539 (N_15539,N_13604,N_13176);
nor U15540 (N_15540,N_13637,N_14944);
and U15541 (N_15541,N_14882,N_13223);
nand U15542 (N_15542,N_14543,N_14346);
nor U15543 (N_15543,N_13411,N_12543);
and U15544 (N_15544,N_14610,N_12912);
nor U15545 (N_15545,N_12817,N_14584);
xnor U15546 (N_15546,N_14339,N_12622);
or U15547 (N_15547,N_13877,N_12701);
xor U15548 (N_15548,N_12589,N_14483);
or U15549 (N_15549,N_12931,N_13025);
nand U15550 (N_15550,N_13134,N_13720);
xor U15551 (N_15551,N_13639,N_12750);
nand U15552 (N_15552,N_14106,N_13563);
and U15553 (N_15553,N_14243,N_14013);
xor U15554 (N_15554,N_14487,N_14418);
nand U15555 (N_15555,N_14320,N_12941);
xnor U15556 (N_15556,N_14938,N_14050);
and U15557 (N_15557,N_12865,N_13941);
and U15558 (N_15558,N_13498,N_14523);
xor U15559 (N_15559,N_13631,N_12578);
or U15560 (N_15560,N_12900,N_13093);
or U15561 (N_15561,N_12773,N_12964);
nor U15562 (N_15562,N_14658,N_14934);
nor U15563 (N_15563,N_13658,N_14575);
xnor U15564 (N_15564,N_14948,N_13868);
and U15565 (N_15565,N_14126,N_13151);
or U15566 (N_15566,N_13871,N_14152);
nand U15567 (N_15567,N_13032,N_12613);
or U15568 (N_15568,N_14111,N_14285);
xor U15569 (N_15569,N_13542,N_13273);
or U15570 (N_15570,N_13256,N_13298);
nor U15571 (N_15571,N_12885,N_13659);
or U15572 (N_15572,N_14876,N_14859);
or U15573 (N_15573,N_14771,N_14605);
or U15574 (N_15574,N_14672,N_13480);
and U15575 (N_15575,N_13856,N_13567);
or U15576 (N_15576,N_14020,N_14191);
xnor U15577 (N_15577,N_13501,N_14381);
nor U15578 (N_15578,N_13989,N_13019);
nor U15579 (N_15579,N_13017,N_14233);
and U15580 (N_15580,N_14635,N_14743);
nand U15581 (N_15581,N_14436,N_13666);
nor U15582 (N_15582,N_14432,N_13253);
xnor U15583 (N_15583,N_14331,N_14456);
xnor U15584 (N_15584,N_14739,N_14686);
nand U15585 (N_15585,N_14738,N_13173);
nand U15586 (N_15586,N_13858,N_13511);
and U15587 (N_15587,N_14967,N_14820);
and U15588 (N_15588,N_13942,N_12942);
xnor U15589 (N_15589,N_14964,N_14995);
xnor U15590 (N_15590,N_14730,N_13464);
nor U15591 (N_15591,N_13876,N_14426);
and U15592 (N_15592,N_13133,N_13804);
nor U15593 (N_15593,N_13117,N_14303);
and U15594 (N_15594,N_12982,N_12844);
nor U15595 (N_15595,N_13143,N_13368);
and U15596 (N_15596,N_13506,N_13711);
or U15597 (N_15597,N_13795,N_12977);
or U15598 (N_15598,N_14467,N_13359);
and U15599 (N_15599,N_13976,N_12573);
and U15600 (N_15600,N_14947,N_12741);
xnor U15601 (N_15601,N_13403,N_14481);
nand U15602 (N_15602,N_13488,N_13837);
xnor U15603 (N_15603,N_14531,N_13481);
and U15604 (N_15604,N_13601,N_12658);
nand U15605 (N_15605,N_13394,N_14291);
nor U15606 (N_15606,N_13009,N_12867);
nand U15607 (N_15607,N_14255,N_14060);
nor U15608 (N_15608,N_14273,N_12540);
xnor U15609 (N_15609,N_13261,N_14832);
or U15610 (N_15610,N_13786,N_12634);
nand U15611 (N_15611,N_13383,N_14140);
and U15612 (N_15612,N_12605,N_13922);
and U15613 (N_15613,N_14237,N_14564);
xor U15614 (N_15614,N_12714,N_13617);
or U15615 (N_15615,N_13168,N_13235);
and U15616 (N_15616,N_13487,N_14165);
and U15617 (N_15617,N_13635,N_14370);
nor U15618 (N_15618,N_12512,N_13644);
xnor U15619 (N_15619,N_14223,N_13517);
xor U15620 (N_15620,N_12624,N_13287);
nand U15621 (N_15621,N_14065,N_14898);
or U15622 (N_15622,N_13124,N_13737);
nor U15623 (N_15623,N_13484,N_14136);
nor U15624 (N_15624,N_13272,N_14770);
nand U15625 (N_15625,N_12810,N_13514);
nor U15626 (N_15626,N_13384,N_13007);
nor U15627 (N_15627,N_14715,N_13973);
or U15628 (N_15628,N_14957,N_12534);
and U15629 (N_15629,N_13371,N_13579);
and U15630 (N_15630,N_13413,N_14364);
nand U15631 (N_15631,N_12640,N_13557);
nor U15632 (N_15632,N_14809,N_13855);
xnor U15633 (N_15633,N_14589,N_14369);
nor U15634 (N_15634,N_14917,N_13363);
nor U15635 (N_15635,N_14580,N_14118);
nor U15636 (N_15636,N_13647,N_14788);
nor U15637 (N_15637,N_12686,N_13222);
nor U15638 (N_15638,N_13886,N_13759);
and U15639 (N_15639,N_13912,N_13859);
nor U15640 (N_15640,N_12851,N_14981);
nand U15641 (N_15641,N_14470,N_13800);
nor U15642 (N_15642,N_13376,N_12788);
and U15643 (N_15643,N_13283,N_13078);
nor U15644 (N_15644,N_12593,N_13054);
and U15645 (N_15645,N_13163,N_13894);
nand U15646 (N_15646,N_13409,N_14640);
nand U15647 (N_15647,N_14352,N_12638);
or U15648 (N_15648,N_14449,N_13304);
and U15649 (N_15649,N_13119,N_12601);
and U15650 (N_15650,N_13216,N_13652);
nand U15651 (N_15651,N_14823,N_13097);
xnor U15652 (N_15652,N_12692,N_12551);
nor U15653 (N_15653,N_14299,N_13274);
nor U15654 (N_15654,N_14061,N_12838);
or U15655 (N_15655,N_14439,N_13169);
or U15656 (N_15656,N_12515,N_14638);
or U15657 (N_15657,N_13193,N_13198);
or U15658 (N_15658,N_14266,N_12513);
or U15659 (N_15659,N_13382,N_12954);
nand U15660 (N_15660,N_13422,N_13281);
and U15661 (N_15661,N_12993,N_12819);
and U15662 (N_15662,N_12975,N_14284);
nand U15663 (N_15663,N_14287,N_12702);
xnor U15664 (N_15664,N_12913,N_14644);
nand U15665 (N_15665,N_12782,N_14047);
nand U15666 (N_15666,N_12727,N_13438);
or U15667 (N_15667,N_14359,N_14656);
and U15668 (N_15668,N_13656,N_13718);
and U15669 (N_15669,N_13044,N_14765);
nor U15670 (N_15670,N_13550,N_12690);
xnor U15671 (N_15671,N_13518,N_12830);
or U15672 (N_15672,N_13901,N_14318);
nor U15673 (N_15673,N_13442,N_13988);
nand U15674 (N_15674,N_14678,N_14837);
or U15675 (N_15675,N_12520,N_14232);
xnor U15676 (N_15676,N_14214,N_14404);
xor U15677 (N_15677,N_14296,N_14270);
or U15678 (N_15678,N_13757,N_14982);
nand U15679 (N_15679,N_12910,N_13585);
or U15680 (N_15680,N_12707,N_14742);
or U15681 (N_15681,N_13146,N_13836);
xnor U15682 (N_15682,N_14560,N_14268);
or U15683 (N_15683,N_12759,N_14434);
or U15684 (N_15684,N_13208,N_13870);
or U15685 (N_15685,N_14400,N_13401);
nand U15686 (N_15686,N_12668,N_14993);
nor U15687 (N_15687,N_14116,N_13045);
or U15688 (N_15688,N_14634,N_13107);
xnor U15689 (N_15689,N_13798,N_13844);
and U15690 (N_15690,N_14053,N_14975);
nor U15691 (N_15691,N_13743,N_13919);
xor U15692 (N_15692,N_14709,N_13244);
nor U15693 (N_15693,N_13918,N_14712);
xor U15694 (N_15694,N_13732,N_13435);
nor U15695 (N_15695,N_12889,N_13387);
xnor U15696 (N_15696,N_14154,N_14454);
xnor U15697 (N_15697,N_14991,N_14261);
xnor U15698 (N_15698,N_12775,N_14391);
nand U15699 (N_15699,N_14680,N_14424);
xor U15700 (N_15700,N_14556,N_14396);
or U15701 (N_15701,N_14023,N_13055);
xor U15702 (N_15702,N_13071,N_13496);
nand U15703 (N_15703,N_12576,N_14572);
and U15704 (N_15704,N_13493,N_14170);
and U15705 (N_15705,N_13482,N_13492);
nand U15706 (N_15706,N_12612,N_14272);
and U15707 (N_15707,N_14092,N_14340);
nor U15708 (N_15708,N_12769,N_14978);
and U15709 (N_15709,N_14378,N_13675);
and U15710 (N_15710,N_14665,N_13950);
nand U15711 (N_15711,N_14113,N_13325);
or U15712 (N_15712,N_14852,N_12966);
and U15713 (N_15713,N_14317,N_14253);
nand U15714 (N_15714,N_14478,N_14160);
nor U15715 (N_15715,N_13768,N_14148);
or U15716 (N_15716,N_14937,N_14216);
nor U15717 (N_15717,N_12751,N_14891);
nand U15718 (N_15718,N_13875,N_14245);
nand U15719 (N_15719,N_14551,N_14677);
and U15720 (N_15720,N_12550,N_13327);
or U15721 (N_15721,N_14752,N_12579);
or U15722 (N_15722,N_13033,N_12595);
nand U15723 (N_15723,N_12664,N_13824);
nand U15724 (N_15724,N_12516,N_13284);
and U15725 (N_15725,N_13606,N_13936);
xor U15726 (N_15726,N_13731,N_14925);
nor U15727 (N_15727,N_14541,N_13470);
nand U15728 (N_15728,N_14172,N_12586);
or U15729 (N_15729,N_14733,N_14297);
nor U15730 (N_15730,N_13129,N_13074);
and U15731 (N_15731,N_14571,N_13512);
and U15732 (N_15732,N_14977,N_14319);
nand U15733 (N_15733,N_13765,N_14247);
or U15734 (N_15734,N_13419,N_13690);
and U15735 (N_15735,N_14103,N_13677);
nor U15736 (N_15736,N_13238,N_13958);
xor U15737 (N_15737,N_13641,N_12827);
or U15738 (N_15738,N_13835,N_13700);
xor U15739 (N_15739,N_14805,N_13348);
nand U15740 (N_15740,N_13622,N_13562);
or U15741 (N_15741,N_13474,N_13263);
nor U15742 (N_15742,N_14546,N_13399);
nor U15743 (N_15743,N_13513,N_13883);
nand U15744 (N_15744,N_13310,N_13340);
xor U15745 (N_15745,N_13764,N_13508);
and U15746 (N_15746,N_12925,N_14218);
and U15747 (N_15747,N_14138,N_14553);
xnor U15748 (N_15748,N_14083,N_14594);
and U15749 (N_15749,N_12560,N_14343);
nand U15750 (N_15750,N_13551,N_13431);
and U15751 (N_15751,N_12661,N_13425);
nor U15752 (N_15752,N_14623,N_13503);
nand U15753 (N_15753,N_13630,N_14563);
and U15754 (N_15754,N_13874,N_13791);
xor U15755 (N_15755,N_14028,N_14070);
and U15756 (N_15756,N_13638,N_12556);
nand U15757 (N_15757,N_14251,N_14618);
nand U15758 (N_15758,N_14835,N_14842);
and U15759 (N_15759,N_13536,N_12537);
nor U15760 (N_15760,N_13504,N_13270);
xnor U15761 (N_15761,N_13929,N_13817);
and U15762 (N_15762,N_12888,N_13098);
xor U15763 (N_15763,N_14295,N_14573);
nand U15764 (N_15764,N_12598,N_14910);
and U15765 (N_15765,N_14288,N_13751);
nand U15766 (N_15766,N_14055,N_14946);
and U15767 (N_15767,N_12787,N_14199);
or U15768 (N_15768,N_12572,N_13570);
or U15769 (N_15769,N_13999,N_14446);
nor U15770 (N_15770,N_13553,N_12722);
or U15771 (N_15771,N_13318,N_14526);
and U15772 (N_15772,N_14465,N_14166);
and U15773 (N_15773,N_14190,N_12709);
and U15774 (N_15774,N_14310,N_12793);
or U15775 (N_15775,N_12610,N_13612);
nand U15776 (N_15776,N_13232,N_12896);
and U15777 (N_15777,N_14139,N_12721);
xnor U15778 (N_15778,N_14822,N_13344);
nand U15779 (N_15779,N_13321,N_12675);
or U15780 (N_15780,N_12797,N_14858);
and U15781 (N_15781,N_13926,N_13028);
xor U15782 (N_15782,N_14509,N_13378);
or U15783 (N_15783,N_13362,N_13102);
or U15784 (N_15784,N_12559,N_13593);
nor U15785 (N_15785,N_12949,N_13393);
or U15786 (N_15786,N_13803,N_13385);
xnor U15787 (N_15787,N_14912,N_14806);
nor U15788 (N_15788,N_14537,N_14052);
nand U15789 (N_15789,N_14660,N_13449);
and U15790 (N_15790,N_12521,N_13455);
or U15791 (N_15791,N_13266,N_14246);
xnor U15792 (N_15792,N_13036,N_12778);
and U15793 (N_15793,N_13708,N_13271);
xnor U15794 (N_15794,N_12708,N_13819);
nor U15795 (N_15795,N_14524,N_13077);
and U15796 (N_15796,N_14555,N_13758);
nand U15797 (N_15797,N_13458,N_14750);
nand U15798 (N_15798,N_12774,N_12917);
xnor U15799 (N_15799,N_13994,N_13159);
nor U15800 (N_15800,N_14112,N_13849);
xnor U15801 (N_15801,N_13296,N_14792);
or U15802 (N_15802,N_14058,N_14198);
nand U15803 (N_15803,N_14048,N_14144);
and U15804 (N_15804,N_13717,N_12632);
xor U15805 (N_15805,N_13772,N_13020);
and U15806 (N_15806,N_14300,N_13329);
and U15807 (N_15807,N_13733,N_12845);
nor U15808 (N_15808,N_13381,N_14033);
and U15809 (N_15809,N_12921,N_13158);
xnor U15810 (N_15810,N_13290,N_13031);
xor U15811 (N_15811,N_13447,N_14932);
nand U15812 (N_15812,N_13598,N_12762);
nand U15813 (N_15813,N_14909,N_12929);
and U15814 (N_15814,N_13706,N_13559);
and U15815 (N_15815,N_13379,N_14511);
or U15816 (N_15816,N_13802,N_13144);
or U15817 (N_15817,N_12881,N_14766);
xnor U15818 (N_15818,N_14324,N_13333);
nand U15819 (N_15819,N_13893,N_12792);
and U15820 (N_15820,N_14134,N_13794);
xnor U15821 (N_15821,N_12581,N_13695);
nand U15822 (N_15822,N_13749,N_14583);
nand U15823 (N_15823,N_12781,N_13351);
nor U15824 (N_15824,N_13767,N_13669);
and U15825 (N_15825,N_13209,N_12926);
xor U15826 (N_15826,N_13191,N_14544);
xor U15827 (N_15827,N_12558,N_14036);
or U15828 (N_15828,N_14875,N_14821);
nor U15829 (N_15829,N_14503,N_12636);
and U15830 (N_15830,N_14961,N_12575);
or U15831 (N_15831,N_13556,N_14682);
nor U15832 (N_15832,N_12712,N_13640);
nand U15833 (N_15833,N_14520,N_12992);
nor U15834 (N_15834,N_14641,N_13320);
nor U15835 (N_15835,N_13014,N_13048);
xnor U15836 (N_15836,N_12749,N_12672);
or U15837 (N_15837,N_14624,N_14128);
nand U15838 (N_15838,N_13689,N_12960);
xor U15839 (N_15839,N_14786,N_14840);
nor U15840 (N_15840,N_12919,N_14443);
or U15841 (N_15841,N_13152,N_13051);
and U15842 (N_15842,N_13683,N_12836);
or U15843 (N_15843,N_13572,N_13907);
or U15844 (N_15844,N_14892,N_14411);
nor U15845 (N_15845,N_13607,N_14802);
or U15846 (N_15846,N_14265,N_14444);
xor U15847 (N_15847,N_13249,N_14918);
nand U15848 (N_15848,N_14188,N_14073);
or U15849 (N_15849,N_14027,N_14851);
and U15850 (N_15850,N_12763,N_12948);
nor U15851 (N_15851,N_14726,N_13214);
or U15852 (N_15852,N_12916,N_14849);
xor U15853 (N_15853,N_12544,N_14522);
nor U15854 (N_15854,N_13424,N_13215);
nand U15855 (N_15855,N_14361,N_13459);
nor U15856 (N_15856,N_13126,N_12620);
xor U15857 (N_15857,N_13984,N_13197);
nand U15858 (N_15858,N_13118,N_13839);
or U15859 (N_15859,N_14490,N_14974);
and U15860 (N_15860,N_12770,N_14162);
or U15861 (N_15861,N_13505,N_14727);
nand U15862 (N_15862,N_14881,N_13404);
and U15863 (N_15863,N_13756,N_14491);
nand U15864 (N_15864,N_12760,N_14447);
or U15865 (N_15865,N_14322,N_14900);
nand U15866 (N_15866,N_13775,N_13867);
and U15867 (N_15867,N_12808,N_14778);
xor U15868 (N_15868,N_13225,N_14696);
nand U15869 (N_15869,N_12678,N_12548);
and U15870 (N_15870,N_12754,N_14228);
nor U15871 (N_15871,N_13610,N_13108);
nor U15872 (N_15872,N_14274,N_14409);
nor U15873 (N_15873,N_13184,N_13547);
nand U15874 (N_15874,N_14980,N_14019);
nand U15875 (N_15875,N_12833,N_12974);
and U15876 (N_15876,N_14016,N_13012);
or U15877 (N_15877,N_14518,N_13013);
xor U15878 (N_15878,N_13478,N_14879);
nand U15879 (N_15879,N_14146,N_13900);
or U15880 (N_15880,N_14202,N_14657);
or U15881 (N_15881,N_14422,N_13164);
or U15882 (N_15882,N_13305,N_13935);
and U15883 (N_15883,N_14314,N_14157);
and U15884 (N_15884,N_13202,N_14030);
and U15885 (N_15885,N_14217,N_14565);
xor U15886 (N_15886,N_12811,N_12524);
or U15887 (N_15887,N_12648,N_14429);
xor U15888 (N_15888,N_14341,N_14846);
nor U15889 (N_15889,N_13986,N_14072);
nor U15890 (N_15890,N_14759,N_13937);
nor U15891 (N_15891,N_12571,N_13820);
or U15892 (N_15892,N_13806,N_13571);
and U15893 (N_15893,N_14206,N_14252);
xor U15894 (N_15894,N_14512,N_14466);
nor U15895 (N_15895,N_13069,N_14180);
nor U15896 (N_15896,N_14886,N_14794);
nor U15897 (N_15897,N_12893,N_14774);
and U15898 (N_15898,N_13738,N_14801);
nor U15899 (N_15899,N_14668,N_13944);
nand U15900 (N_15900,N_13448,N_12988);
nand U15901 (N_15901,N_13902,N_13761);
xnor U15902 (N_15902,N_12719,N_14667);
or U15903 (N_15903,N_14347,N_13713);
xnor U15904 (N_15904,N_12710,N_12835);
nand U15905 (N_15905,N_12996,N_13259);
and U15906 (N_15906,N_14009,N_12837);
nor U15907 (N_15907,N_14813,N_13809);
or U15908 (N_15908,N_13566,N_13996);
nor U15909 (N_15909,N_12984,N_13291);
nor U15910 (N_15910,N_13499,N_12735);
nor U15911 (N_15911,N_13285,N_13234);
nand U15912 (N_15912,N_14187,N_12933);
and U15913 (N_15913,N_14700,N_14074);
nand U15914 (N_15914,N_13699,N_13943);
xnor U15915 (N_15915,N_12630,N_12877);
and U15916 (N_15916,N_14024,N_14869);
or U15917 (N_15917,N_13752,N_13963);
and U15918 (N_15918,N_12899,N_14843);
nand U15919 (N_15919,N_13450,N_13060);
and U15920 (N_15920,N_14905,N_12961);
xnor U15921 (N_15921,N_14828,N_14182);
nor U15922 (N_15922,N_14489,N_13784);
nand U15923 (N_15923,N_14502,N_12794);
and U15924 (N_15924,N_13880,N_14168);
and U15925 (N_15925,N_14872,N_14386);
nor U15926 (N_15926,N_13822,N_13171);
nand U15927 (N_15927,N_14197,N_13282);
xor U15928 (N_15928,N_13845,N_13846);
or U15929 (N_15929,N_13938,N_13651);
and U15930 (N_15930,N_14795,N_14002);
xnor U15931 (N_15931,N_13916,N_13292);
nand U15932 (N_15932,N_12603,N_14989);
or U15933 (N_15933,N_14360,N_12611);
or U15934 (N_15934,N_13135,N_14907);
or U15935 (N_15935,N_14698,N_14408);
or U15936 (N_15936,N_13463,N_14724);
or U15937 (N_15937,N_13177,N_13814);
nand U15938 (N_15938,N_13286,N_12728);
nand U15939 (N_15939,N_13977,N_14321);
xnor U15940 (N_15940,N_14894,N_13754);
and U15941 (N_15941,N_14236,N_13324);
and U15942 (N_15942,N_14189,N_13322);
nor U15943 (N_15943,N_13590,N_13873);
and U15944 (N_15944,N_13515,N_13094);
nor U15945 (N_15945,N_12667,N_14040);
or U15946 (N_15946,N_13725,N_12965);
nor U15947 (N_15947,N_13555,N_12568);
and U15948 (N_15948,N_12947,N_13539);
xor U15949 (N_15949,N_13293,N_14824);
xor U15950 (N_15950,N_12976,N_12862);
and U15951 (N_15951,N_12779,N_12563);
nor U15952 (N_15952,N_13681,N_14800);
or U15953 (N_15953,N_13494,N_12685);
xnor U15954 (N_15954,N_13149,N_14810);
or U15955 (N_15955,N_13194,N_14181);
and U15956 (N_15956,N_12643,N_14099);
nand U15957 (N_15957,N_13864,N_14570);
and U15958 (N_15958,N_13181,N_14421);
or U15959 (N_15959,N_13416,N_13116);
and U15960 (N_15960,N_13115,N_12935);
nand U15961 (N_15961,N_14513,N_12980);
and U15962 (N_15962,N_14208,N_14271);
nand U15963 (N_15963,N_12649,N_14999);
or U15964 (N_15964,N_13642,N_13892);
nand U15965 (N_15965,N_13895,N_14063);
or U15966 (N_15966,N_13714,N_12506);
nand U15967 (N_15967,N_14435,N_13698);
nand U15968 (N_15968,N_14643,N_14783);
nor U15969 (N_15969,N_13552,N_12739);
xor U15970 (N_15970,N_14067,N_12583);
nand U15971 (N_15971,N_14158,N_14183);
xnor U15972 (N_15972,N_13687,N_13816);
nand U15973 (N_15973,N_13061,N_14281);
and U15974 (N_15974,N_13522,N_14279);
and U15975 (N_15975,N_14084,N_12963);
xor U15976 (N_15976,N_14493,N_13352);
nor U15977 (N_15977,N_14088,N_14452);
or U15978 (N_15978,N_14129,N_13869);
xnor U15979 (N_15979,N_13983,N_14860);
nand U15980 (N_15980,N_13237,N_12924);
nand U15981 (N_15981,N_13881,N_14194);
nand U15982 (N_15982,N_13830,N_14250);
nand U15983 (N_15983,N_14469,N_14390);
nor U15984 (N_15984,N_12818,N_12956);
or U15985 (N_15985,N_14348,N_13882);
nor U15986 (N_15986,N_13417,N_14637);
nand U15987 (N_15987,N_14221,N_14939);
nand U15988 (N_15988,N_14071,N_13540);
nor U15989 (N_15989,N_14857,N_13317);
or U15990 (N_15990,N_14405,N_13620);
nand U15991 (N_15991,N_12874,N_14548);
or U15992 (N_15992,N_13370,N_12831);
or U15993 (N_15993,N_14442,N_13946);
xnor U15994 (N_15994,N_14536,N_13521);
and U15995 (N_15995,N_13410,N_13828);
nor U15996 (N_15996,N_13148,N_13165);
and U15997 (N_15997,N_14772,N_13679);
and U15998 (N_15998,N_13621,N_13157);
or U15999 (N_15999,N_14596,N_13367);
nand U16000 (N_16000,N_14533,N_12514);
xor U16001 (N_16001,N_12720,N_13611);
nand U16002 (N_16002,N_14433,N_14220);
nor U16003 (N_16003,N_13696,N_13735);
xor U16004 (N_16004,N_14979,N_12843);
nor U16005 (N_16005,N_13688,N_14532);
nand U16006 (N_16006,N_12936,N_13843);
nand U16007 (N_16007,N_14383,N_13254);
nor U16008 (N_16008,N_14992,N_14785);
nand U16009 (N_16009,N_14562,N_14312);
or U16010 (N_16010,N_13785,N_14602);
nor U16011 (N_16011,N_14581,N_14648);
nor U16012 (N_16012,N_14633,N_13554);
nor U16013 (N_16013,N_12509,N_13627);
nor U16014 (N_16014,N_13580,N_13374);
nand U16015 (N_16015,N_13155,N_14517);
or U16016 (N_16016,N_14085,N_13628);
and U16017 (N_16017,N_14046,N_14457);
nand U16018 (N_16018,N_12700,N_14748);
nor U16019 (N_16019,N_14775,N_12666);
and U16020 (N_16020,N_13392,N_14461);
and U16021 (N_16021,N_14697,N_12826);
and U16022 (N_16022,N_12847,N_14004);
nor U16023 (N_16023,N_12911,N_14280);
xor U16024 (N_16024,N_12969,N_13388);
xor U16025 (N_16025,N_14001,N_13207);
or U16026 (N_16026,N_14419,N_14699);
xnor U16027 (N_16027,N_14504,N_13664);
xnor U16028 (N_16028,N_12552,N_14306);
or U16029 (N_16029,N_13541,N_13172);
and U16030 (N_16030,N_13797,N_13668);
and U16031 (N_16031,N_13395,N_13456);
xnor U16032 (N_16032,N_14737,N_14559);
or U16033 (N_16033,N_14959,N_13467);
and U16034 (N_16034,N_14561,N_14384);
and U16035 (N_16035,N_13053,N_13128);
and U16036 (N_16036,N_13671,N_13396);
xor U16037 (N_16037,N_13461,N_14012);
xor U16038 (N_16038,N_14549,N_13407);
and U16039 (N_16039,N_14334,N_12909);
nand U16040 (N_16040,N_12587,N_14423);
xnor U16041 (N_16041,N_13613,N_13951);
nand U16042 (N_16042,N_12765,N_14499);
xnor U16043 (N_16043,N_13833,N_14629);
nand U16044 (N_16044,N_14519,N_12859);
nand U16045 (N_16045,N_12799,N_12505);
or U16046 (N_16046,N_13783,N_14673);
nand U16047 (N_16047,N_13027,N_12858);
nor U16048 (N_16048,N_12617,N_12554);
or U16049 (N_16049,N_13812,N_13851);
nand U16050 (N_16050,N_14725,N_14108);
nor U16051 (N_16051,N_13477,N_14935);
xnor U16052 (N_16052,N_14625,N_13861);
xnor U16053 (N_16053,N_12849,N_13242);
xor U16054 (N_16054,N_13825,N_13203);
and U16055 (N_16055,N_13068,N_14632);
nor U16056 (N_16056,N_14612,N_12832);
xnor U16057 (N_16057,N_14345,N_13670);
or U16058 (N_16058,N_13530,N_12596);
nand U16059 (N_16059,N_13299,N_12566);
or U16060 (N_16060,N_14286,N_14747);
xor U16061 (N_16061,N_13080,N_13904);
nand U16062 (N_16062,N_13462,N_14923);
xnor U16063 (N_16063,N_12604,N_12986);
nor U16064 (N_16064,N_12938,N_13502);
nand U16065 (N_16065,N_14069,N_12651);
or U16066 (N_16066,N_13182,N_14814);
or U16067 (N_16067,N_12639,N_14527);
and U16068 (N_16068,N_13933,N_13067);
nand U16069 (N_16069,N_12915,N_12619);
nor U16070 (N_16070,N_14402,N_14239);
xnor U16071 (N_16071,N_14018,N_13703);
xor U16072 (N_16072,N_13228,N_12625);
or U16073 (N_16073,N_14740,N_12644);
or U16074 (N_16074,N_13443,N_13089);
nor U16075 (N_16075,N_14716,N_14790);
or U16076 (N_16076,N_13186,N_14915);
xnor U16077 (N_16077,N_13863,N_12814);
xnor U16078 (N_16078,N_13945,N_13605);
nor U16079 (N_16079,N_12813,N_14825);
nor U16080 (N_16080,N_12745,N_13564);
nand U16081 (N_16081,N_14626,N_14153);
nand U16082 (N_16082,N_13526,N_12898);
xnor U16083 (N_16083,N_13204,N_14812);
or U16084 (N_16084,N_14351,N_14308);
nor U16085 (N_16085,N_14017,N_14066);
or U16086 (N_16086,N_13454,N_13584);
xnor U16087 (N_16087,N_12755,N_13406);
xnor U16088 (N_16088,N_14685,N_13418);
nor U16089 (N_16089,N_14507,N_13582);
nor U16090 (N_16090,N_13489,N_13316);
or U16091 (N_16091,N_14681,N_14328);
nor U16092 (N_16092,N_14262,N_14889);
nor U16093 (N_16093,N_13252,N_12995);
xnor U16094 (N_16094,N_12706,N_13838);
or U16095 (N_16095,N_13507,N_14723);
nand U16096 (N_16096,N_14628,N_14174);
nand U16097 (N_16097,N_14998,N_13692);
xor U16098 (N_16098,N_12972,N_13346);
xnor U16099 (N_16099,N_14670,N_14464);
and U16100 (N_16100,N_13970,N_14855);
nand U16101 (N_16101,N_14460,N_13805);
nor U16102 (N_16102,N_12771,N_13338);
and U16103 (N_16103,N_13787,N_13161);
nand U16104 (N_16104,N_14516,N_12897);
or U16105 (N_16105,N_14746,N_13616);
or U16106 (N_16106,N_14290,N_14619);
and U16107 (N_16107,N_13755,N_14484);
nor U16108 (N_16108,N_13096,N_13500);
nand U16109 (N_16109,N_12761,N_13729);
or U16110 (N_16110,N_14440,N_13180);
nand U16111 (N_16111,N_14850,N_13643);
or U16112 (N_16112,N_12800,N_14387);
xnor U16113 (N_16113,N_14412,N_14608);
nand U16114 (N_16114,N_14311,N_14398);
nor U16115 (N_16115,N_12878,N_12880);
or U16116 (N_16116,N_12656,N_14374);
nand U16117 (N_16117,N_13076,N_12525);
and U16118 (N_16118,N_13890,N_12635);
nand U16119 (N_16119,N_14695,N_14278);
or U16120 (N_16120,N_14779,N_13948);
nor U16121 (N_16121,N_13587,N_14123);
or U16122 (N_16122,N_13528,N_14713);
nor U16123 (N_16123,N_14609,N_12738);
nor U16124 (N_16124,N_14075,N_13730);
or U16125 (N_16125,N_13104,N_14827);
xor U16126 (N_16126,N_13323,N_14731);
xor U16127 (N_16127,N_12669,N_12970);
nand U16128 (N_16128,N_12962,N_13532);
or U16129 (N_16129,N_14453,N_13615);
nand U16130 (N_16130,N_14211,N_13170);
or U16131 (N_16131,N_14588,N_13217);
xnor U16132 (N_16132,N_12842,N_13992);
nor U16133 (N_16133,N_12660,N_14427);
nand U16134 (N_16134,N_14702,N_13623);
nand U16135 (N_16135,N_13744,N_12650);
nor U16136 (N_16136,N_14362,N_13046);
nor U16137 (N_16137,N_13646,N_14081);
or U16138 (N_16138,N_14636,N_13231);
and U16139 (N_16139,N_14089,N_14375);
or U16140 (N_16140,N_14186,N_13059);
and U16141 (N_16141,N_14344,N_12883);
xnor U16142 (N_16142,N_14962,N_13519);
or U16143 (N_16143,N_13372,N_13491);
and U16144 (N_16144,N_14229,N_14874);
nor U16145 (N_16145,N_14358,N_12518);
nand U16146 (N_16146,N_13549,N_14542);
or U16147 (N_16147,N_12695,N_14034);
and U16148 (N_16148,N_14990,N_13626);
xor U16149 (N_16149,N_14054,N_12876);
xor U16150 (N_16150,N_13697,N_12729);
nor U16151 (N_16151,N_12801,N_13747);
and U16152 (N_16152,N_14076,N_14768);
xor U16153 (N_16153,N_12879,N_13188);
xor U16154 (N_16154,N_14201,N_13609);
xor U16155 (N_16155,N_13850,N_13660);
nand U16156 (N_16156,N_13594,N_14902);
nand U16157 (N_16157,N_13774,N_14863);
and U16158 (N_16158,N_14574,N_14156);
nor U16159 (N_16159,N_14754,N_14601);
nand U16160 (N_16160,N_12737,N_14956);
or U16161 (N_16161,N_14758,N_14087);
and U16162 (N_16162,N_14326,N_12628);
nor U16163 (N_16163,N_12907,N_13741);
nor U16164 (N_16164,N_14325,N_13762);
and U16165 (N_16165,N_14107,N_12561);
nand U16166 (N_16166,N_13766,N_14091);
and U16167 (N_16167,N_13345,N_14793);
nand U16168 (N_16168,N_14597,N_14950);
nor U16169 (N_16169,N_13650,N_14149);
xnor U16170 (N_16170,N_14569,N_14441);
xnor U16171 (N_16171,N_12780,N_14789);
nor U16172 (N_16172,N_13280,N_14847);
and U16173 (N_16173,N_14579,N_13534);
or U16174 (N_16174,N_12618,N_12904);
xnor U16175 (N_16175,N_14799,N_14209);
xor U16176 (N_16176,N_14862,N_13423);
nand U16177 (N_16177,N_13807,N_12967);
and U16178 (N_16178,N_12920,N_13624);
and U16179 (N_16179,N_14062,N_14538);
nand U16180 (N_16180,N_13201,N_13264);
nor U16181 (N_16181,N_14831,N_13335);
xor U16182 (N_16182,N_14227,N_14749);
nor U16183 (N_16183,N_14125,N_13056);
nor U16184 (N_16184,N_14130,N_13657);
nand U16185 (N_16185,N_14041,N_13356);
xnor U16186 (N_16186,N_13964,N_14965);
nor U16187 (N_16187,N_12647,N_12932);
and U16188 (N_16188,N_12860,N_13047);
nand U16189 (N_16189,N_12922,N_13132);
and U16190 (N_16190,N_13219,N_14617);
nand U16191 (N_16191,N_13109,N_14631);
and U16192 (N_16192,N_13884,N_13632);
or U16193 (N_16193,N_13160,N_14242);
xor U16194 (N_16194,N_13909,N_12734);
and U16195 (N_16195,N_12934,N_12731);
xnor U16196 (N_16196,N_14988,N_14472);
nor U16197 (N_16197,N_13777,N_14550);
and U16198 (N_16198,N_14102,N_14603);
nand U16199 (N_16199,N_14045,N_13079);
nand U16200 (N_16200,N_14121,N_14706);
nand U16201 (N_16201,N_12665,N_14521);
nor U16202 (N_16202,N_14455,N_13154);
nor U16203 (N_16203,N_13853,N_14097);
nor U16204 (N_16204,N_13840,N_13022);
or U16205 (N_16205,N_13358,N_13427);
nor U16206 (N_16206,N_13452,N_14614);
xnor U16207 (N_16207,N_14645,N_14986);
or U16208 (N_16208,N_14798,N_13178);
nand U16209 (N_16209,N_13257,N_13516);
xnor U16210 (N_16210,N_14276,N_13490);
xnor U16211 (N_16211,N_12609,N_13726);
or U16212 (N_16212,N_13187,N_12693);
xor U16213 (N_16213,N_13475,N_13211);
or U16214 (N_16214,N_12742,N_13131);
xor U16215 (N_16215,N_13268,N_14913);
nor U16216 (N_16216,N_12592,N_13166);
xnor U16217 (N_16217,N_14595,N_14203);
and U16218 (N_16218,N_12903,N_14301);
or U16219 (N_16219,N_13018,N_13010);
and U16220 (N_16220,N_14363,N_13476);
or U16221 (N_16221,N_13088,N_13307);
and U16222 (N_16222,N_14215,N_13030);
nand U16223 (N_16223,N_13865,N_14051);
and U16224 (N_16224,N_14535,N_12946);
nand U16225 (N_16225,N_13578,N_13591);
and U16226 (N_16226,N_13227,N_13156);
or U16227 (N_16227,N_13453,N_13661);
or U16228 (N_16228,N_14620,N_13343);
nand U16229 (N_16229,N_14663,N_12532);
nand U16230 (N_16230,N_12691,N_13799);
xor U16231 (N_16231,N_14654,N_13397);
xor U16232 (N_16232,N_13199,N_13073);
nor U16233 (N_16233,N_13740,N_13114);
or U16234 (N_16234,N_14856,N_14762);
xnor U16235 (N_16235,N_14650,N_13112);
xnor U16236 (N_16236,N_13328,N_13457);
nor U16237 (N_16237,N_14592,N_14480);
or U16238 (N_16238,N_12804,N_13702);
or U16239 (N_16239,N_13140,N_13537);
and U16240 (N_16240,N_13196,N_13829);
and U16241 (N_16241,N_14090,N_13262);
or U16242 (N_16242,N_14870,N_13716);
nand U16243 (N_16243,N_14613,N_12863);
and U16244 (N_16244,N_14552,N_12852);
or U16245 (N_16245,N_13190,N_14224);
or U16246 (N_16246,N_12688,N_13705);
or U16247 (N_16247,N_13120,N_13770);
nor U16248 (N_16248,N_13432,N_14445);
nand U16249 (N_16249,N_14371,N_13445);
or U16250 (N_16250,N_12667,N_12702);
or U16251 (N_16251,N_14550,N_13115);
xnor U16252 (N_16252,N_14666,N_12646);
xnor U16253 (N_16253,N_14260,N_14262);
and U16254 (N_16254,N_13768,N_13908);
nor U16255 (N_16255,N_12986,N_13960);
and U16256 (N_16256,N_14823,N_12505);
nor U16257 (N_16257,N_12935,N_13588);
and U16258 (N_16258,N_14856,N_12902);
xor U16259 (N_16259,N_12937,N_13385);
nor U16260 (N_16260,N_12862,N_14537);
nor U16261 (N_16261,N_14082,N_12994);
xor U16262 (N_16262,N_14983,N_14117);
and U16263 (N_16263,N_14734,N_14660);
xnor U16264 (N_16264,N_13848,N_13646);
nand U16265 (N_16265,N_13389,N_12588);
nor U16266 (N_16266,N_13701,N_13655);
nand U16267 (N_16267,N_13777,N_13630);
and U16268 (N_16268,N_13951,N_14296);
and U16269 (N_16269,N_13385,N_14180);
and U16270 (N_16270,N_13514,N_13515);
or U16271 (N_16271,N_14392,N_14651);
xnor U16272 (N_16272,N_12883,N_14564);
xnor U16273 (N_16273,N_14301,N_14925);
or U16274 (N_16274,N_14978,N_13129);
nor U16275 (N_16275,N_12884,N_14747);
xor U16276 (N_16276,N_14340,N_13745);
xor U16277 (N_16277,N_13059,N_14157);
xor U16278 (N_16278,N_12874,N_12588);
nor U16279 (N_16279,N_13569,N_14262);
and U16280 (N_16280,N_13706,N_12906);
and U16281 (N_16281,N_12728,N_14663);
nand U16282 (N_16282,N_14018,N_12769);
or U16283 (N_16283,N_13792,N_12606);
nand U16284 (N_16284,N_13546,N_14637);
or U16285 (N_16285,N_13765,N_13305);
nor U16286 (N_16286,N_14759,N_13407);
nand U16287 (N_16287,N_14745,N_12982);
nor U16288 (N_16288,N_13386,N_14703);
xor U16289 (N_16289,N_12743,N_14475);
and U16290 (N_16290,N_14376,N_13635);
nor U16291 (N_16291,N_14423,N_14352);
and U16292 (N_16292,N_12893,N_13863);
and U16293 (N_16293,N_14255,N_14433);
xnor U16294 (N_16294,N_13434,N_13700);
or U16295 (N_16295,N_12872,N_12617);
nand U16296 (N_16296,N_14304,N_13726);
nor U16297 (N_16297,N_14044,N_13402);
and U16298 (N_16298,N_13911,N_12844);
or U16299 (N_16299,N_12551,N_14613);
nand U16300 (N_16300,N_14090,N_14760);
nor U16301 (N_16301,N_13087,N_14174);
or U16302 (N_16302,N_14328,N_13492);
nor U16303 (N_16303,N_12703,N_14219);
nand U16304 (N_16304,N_14929,N_14467);
or U16305 (N_16305,N_14747,N_13511);
xnor U16306 (N_16306,N_14619,N_14352);
and U16307 (N_16307,N_12984,N_14737);
nor U16308 (N_16308,N_14595,N_14157);
xnor U16309 (N_16309,N_13671,N_14798);
nor U16310 (N_16310,N_12976,N_14043);
nand U16311 (N_16311,N_13105,N_13109);
xor U16312 (N_16312,N_14195,N_12992);
and U16313 (N_16313,N_14061,N_13046);
nand U16314 (N_16314,N_14408,N_14178);
or U16315 (N_16315,N_14946,N_13091);
nand U16316 (N_16316,N_14598,N_13336);
nand U16317 (N_16317,N_14499,N_12672);
xnor U16318 (N_16318,N_14988,N_13329);
nand U16319 (N_16319,N_14565,N_13370);
nor U16320 (N_16320,N_14731,N_12814);
or U16321 (N_16321,N_13633,N_12525);
nand U16322 (N_16322,N_12704,N_12649);
xor U16323 (N_16323,N_13678,N_14833);
or U16324 (N_16324,N_14159,N_13438);
nor U16325 (N_16325,N_14736,N_14195);
xnor U16326 (N_16326,N_14985,N_14735);
or U16327 (N_16327,N_13644,N_12847);
nor U16328 (N_16328,N_12578,N_13821);
or U16329 (N_16329,N_13296,N_14928);
nor U16330 (N_16330,N_13008,N_13378);
xor U16331 (N_16331,N_14580,N_13268);
xnor U16332 (N_16332,N_14376,N_14123);
nor U16333 (N_16333,N_13271,N_14072);
or U16334 (N_16334,N_12705,N_14118);
nor U16335 (N_16335,N_14772,N_12681);
and U16336 (N_16336,N_13157,N_13320);
nand U16337 (N_16337,N_13086,N_12876);
or U16338 (N_16338,N_14916,N_14231);
and U16339 (N_16339,N_13298,N_13230);
nand U16340 (N_16340,N_12796,N_12819);
nand U16341 (N_16341,N_13142,N_14884);
xor U16342 (N_16342,N_12754,N_14767);
nand U16343 (N_16343,N_14653,N_14837);
nand U16344 (N_16344,N_13782,N_13154);
xnor U16345 (N_16345,N_13585,N_12788);
nand U16346 (N_16346,N_13164,N_13606);
nand U16347 (N_16347,N_12996,N_14920);
and U16348 (N_16348,N_12829,N_13093);
nand U16349 (N_16349,N_13508,N_14055);
and U16350 (N_16350,N_12977,N_13103);
and U16351 (N_16351,N_13960,N_14477);
or U16352 (N_16352,N_13966,N_12656);
nor U16353 (N_16353,N_14048,N_14073);
nor U16354 (N_16354,N_13811,N_13814);
nor U16355 (N_16355,N_14687,N_13025);
xor U16356 (N_16356,N_14432,N_14177);
and U16357 (N_16357,N_13765,N_14223);
and U16358 (N_16358,N_12884,N_13784);
or U16359 (N_16359,N_13381,N_14713);
and U16360 (N_16360,N_13003,N_14594);
nor U16361 (N_16361,N_14583,N_13449);
nor U16362 (N_16362,N_13099,N_12512);
or U16363 (N_16363,N_13834,N_13612);
or U16364 (N_16364,N_12973,N_13357);
and U16365 (N_16365,N_12918,N_13452);
nor U16366 (N_16366,N_12607,N_14849);
and U16367 (N_16367,N_13812,N_13696);
or U16368 (N_16368,N_14772,N_12788);
and U16369 (N_16369,N_14429,N_14191);
and U16370 (N_16370,N_12770,N_14297);
and U16371 (N_16371,N_14448,N_14835);
nand U16372 (N_16372,N_13286,N_13757);
and U16373 (N_16373,N_13283,N_12579);
nand U16374 (N_16374,N_13193,N_12759);
or U16375 (N_16375,N_12621,N_12908);
xnor U16376 (N_16376,N_13611,N_14466);
nor U16377 (N_16377,N_12933,N_14030);
nand U16378 (N_16378,N_12782,N_13625);
nor U16379 (N_16379,N_14564,N_14112);
nand U16380 (N_16380,N_14559,N_14794);
xor U16381 (N_16381,N_14755,N_13212);
nand U16382 (N_16382,N_14293,N_14671);
xnor U16383 (N_16383,N_14852,N_13338);
or U16384 (N_16384,N_14608,N_12869);
and U16385 (N_16385,N_12784,N_14612);
xnor U16386 (N_16386,N_13763,N_14475);
xnor U16387 (N_16387,N_14569,N_14507);
or U16388 (N_16388,N_13901,N_14495);
nand U16389 (N_16389,N_14820,N_12571);
or U16390 (N_16390,N_13503,N_14175);
nor U16391 (N_16391,N_14808,N_12797);
or U16392 (N_16392,N_14948,N_13372);
xnor U16393 (N_16393,N_13501,N_14723);
nor U16394 (N_16394,N_14030,N_14705);
or U16395 (N_16395,N_12635,N_14056);
nor U16396 (N_16396,N_14786,N_13103);
or U16397 (N_16397,N_13415,N_13392);
and U16398 (N_16398,N_14082,N_14961);
xor U16399 (N_16399,N_13442,N_14476);
and U16400 (N_16400,N_13246,N_14492);
xor U16401 (N_16401,N_13323,N_14952);
and U16402 (N_16402,N_14806,N_12790);
or U16403 (N_16403,N_13270,N_12865);
nand U16404 (N_16404,N_13816,N_14112);
xnor U16405 (N_16405,N_14679,N_13949);
and U16406 (N_16406,N_12783,N_13407);
and U16407 (N_16407,N_12717,N_13063);
nor U16408 (N_16408,N_14288,N_12862);
nor U16409 (N_16409,N_14657,N_13079);
and U16410 (N_16410,N_14975,N_12503);
nand U16411 (N_16411,N_14574,N_12662);
and U16412 (N_16412,N_14662,N_12517);
or U16413 (N_16413,N_14421,N_12514);
xor U16414 (N_16414,N_14163,N_13317);
and U16415 (N_16415,N_14600,N_13202);
and U16416 (N_16416,N_13954,N_12598);
nor U16417 (N_16417,N_13769,N_14919);
nor U16418 (N_16418,N_14063,N_14518);
xnor U16419 (N_16419,N_13604,N_14906);
xnor U16420 (N_16420,N_13509,N_14177);
and U16421 (N_16421,N_14330,N_13751);
nor U16422 (N_16422,N_12584,N_12815);
and U16423 (N_16423,N_13134,N_12627);
xnor U16424 (N_16424,N_13964,N_14392);
and U16425 (N_16425,N_13127,N_13934);
and U16426 (N_16426,N_14937,N_12650);
and U16427 (N_16427,N_13845,N_13171);
nor U16428 (N_16428,N_14772,N_13103);
nand U16429 (N_16429,N_14712,N_14308);
nor U16430 (N_16430,N_14101,N_13761);
and U16431 (N_16431,N_13795,N_12654);
xor U16432 (N_16432,N_13231,N_13646);
nand U16433 (N_16433,N_12634,N_14388);
nor U16434 (N_16434,N_13495,N_12788);
nand U16435 (N_16435,N_14586,N_13466);
or U16436 (N_16436,N_12822,N_13426);
xor U16437 (N_16437,N_14729,N_13088);
nor U16438 (N_16438,N_13780,N_14891);
and U16439 (N_16439,N_12925,N_13845);
xor U16440 (N_16440,N_13287,N_13981);
and U16441 (N_16441,N_13089,N_14206);
or U16442 (N_16442,N_12532,N_14226);
xnor U16443 (N_16443,N_14625,N_12922);
and U16444 (N_16444,N_13686,N_13331);
nand U16445 (N_16445,N_13401,N_13862);
and U16446 (N_16446,N_13084,N_14214);
or U16447 (N_16447,N_13020,N_12894);
or U16448 (N_16448,N_14296,N_13230);
and U16449 (N_16449,N_13193,N_14227);
or U16450 (N_16450,N_14858,N_14584);
xor U16451 (N_16451,N_13444,N_14581);
nor U16452 (N_16452,N_12665,N_14003);
and U16453 (N_16453,N_13245,N_13944);
nor U16454 (N_16454,N_14024,N_13480);
xnor U16455 (N_16455,N_13301,N_13528);
nor U16456 (N_16456,N_12787,N_13143);
xnor U16457 (N_16457,N_13710,N_13646);
xnor U16458 (N_16458,N_12875,N_13598);
and U16459 (N_16459,N_13649,N_13134);
or U16460 (N_16460,N_13824,N_12874);
nand U16461 (N_16461,N_14057,N_14531);
and U16462 (N_16462,N_13348,N_14701);
or U16463 (N_16463,N_14361,N_14370);
nand U16464 (N_16464,N_13186,N_14898);
xor U16465 (N_16465,N_14664,N_14434);
and U16466 (N_16466,N_13529,N_14745);
xor U16467 (N_16467,N_14508,N_13414);
xnor U16468 (N_16468,N_13291,N_13647);
nor U16469 (N_16469,N_12710,N_14379);
or U16470 (N_16470,N_14126,N_14670);
nand U16471 (N_16471,N_12714,N_14556);
nand U16472 (N_16472,N_14820,N_12882);
nor U16473 (N_16473,N_14122,N_14882);
and U16474 (N_16474,N_13469,N_14585);
and U16475 (N_16475,N_14434,N_14424);
nand U16476 (N_16476,N_14460,N_12621);
xnor U16477 (N_16477,N_13427,N_14510);
nor U16478 (N_16478,N_13965,N_13711);
or U16479 (N_16479,N_13337,N_13734);
nand U16480 (N_16480,N_12810,N_14400);
and U16481 (N_16481,N_14346,N_14851);
and U16482 (N_16482,N_14935,N_13222);
nand U16483 (N_16483,N_14557,N_12915);
nor U16484 (N_16484,N_13980,N_12657);
nand U16485 (N_16485,N_12676,N_14886);
and U16486 (N_16486,N_12958,N_12858);
xnor U16487 (N_16487,N_14244,N_12786);
nand U16488 (N_16488,N_14121,N_13631);
or U16489 (N_16489,N_13286,N_13171);
nor U16490 (N_16490,N_13949,N_12892);
nand U16491 (N_16491,N_13308,N_14751);
nand U16492 (N_16492,N_14676,N_13419);
nand U16493 (N_16493,N_14487,N_12663);
nand U16494 (N_16494,N_14126,N_13036);
xor U16495 (N_16495,N_14109,N_13196);
nand U16496 (N_16496,N_14799,N_14552);
or U16497 (N_16497,N_13498,N_13108);
nand U16498 (N_16498,N_13577,N_13123);
nand U16499 (N_16499,N_13412,N_13527);
or U16500 (N_16500,N_12963,N_14760);
or U16501 (N_16501,N_12556,N_14795);
or U16502 (N_16502,N_13238,N_14246);
or U16503 (N_16503,N_12732,N_13713);
or U16504 (N_16504,N_12932,N_13363);
or U16505 (N_16505,N_14463,N_13195);
nor U16506 (N_16506,N_14410,N_14932);
or U16507 (N_16507,N_14353,N_12697);
nand U16508 (N_16508,N_12866,N_14553);
nor U16509 (N_16509,N_14616,N_12529);
nand U16510 (N_16510,N_12529,N_13941);
and U16511 (N_16511,N_14420,N_13603);
nor U16512 (N_16512,N_13778,N_14312);
nor U16513 (N_16513,N_12676,N_13500);
xor U16514 (N_16514,N_12900,N_12982);
nor U16515 (N_16515,N_14691,N_13856);
nand U16516 (N_16516,N_13500,N_14595);
nor U16517 (N_16517,N_14032,N_13062);
or U16518 (N_16518,N_14963,N_13631);
or U16519 (N_16519,N_14307,N_13728);
nor U16520 (N_16520,N_14555,N_13741);
or U16521 (N_16521,N_13155,N_14605);
xor U16522 (N_16522,N_12514,N_14160);
and U16523 (N_16523,N_12884,N_13101);
xnor U16524 (N_16524,N_14574,N_12705);
xor U16525 (N_16525,N_13583,N_12611);
xor U16526 (N_16526,N_14055,N_13950);
nor U16527 (N_16527,N_13853,N_12815);
xor U16528 (N_16528,N_12826,N_14680);
nor U16529 (N_16529,N_13376,N_14172);
or U16530 (N_16530,N_13215,N_14609);
nor U16531 (N_16531,N_13865,N_13221);
nor U16532 (N_16532,N_14311,N_12505);
nand U16533 (N_16533,N_12564,N_13800);
nor U16534 (N_16534,N_14919,N_12818);
nor U16535 (N_16535,N_12540,N_14332);
xor U16536 (N_16536,N_14062,N_13946);
nor U16537 (N_16537,N_14681,N_13652);
nand U16538 (N_16538,N_14201,N_13102);
xnor U16539 (N_16539,N_13957,N_13871);
xnor U16540 (N_16540,N_14318,N_14577);
or U16541 (N_16541,N_14296,N_13738);
nor U16542 (N_16542,N_14049,N_13104);
or U16543 (N_16543,N_13045,N_14111);
xnor U16544 (N_16544,N_12502,N_12770);
nor U16545 (N_16545,N_12747,N_14176);
xnor U16546 (N_16546,N_13406,N_13626);
and U16547 (N_16547,N_13917,N_14529);
nor U16548 (N_16548,N_13106,N_13926);
or U16549 (N_16549,N_12587,N_14998);
nand U16550 (N_16550,N_14719,N_13741);
nand U16551 (N_16551,N_14939,N_14315);
and U16552 (N_16552,N_13897,N_14697);
and U16553 (N_16553,N_14076,N_13386);
and U16554 (N_16554,N_14739,N_12886);
xor U16555 (N_16555,N_13017,N_13367);
nor U16556 (N_16556,N_12895,N_12628);
xor U16557 (N_16557,N_12603,N_13406);
nand U16558 (N_16558,N_14583,N_13397);
and U16559 (N_16559,N_14458,N_12587);
nor U16560 (N_16560,N_14192,N_13983);
nand U16561 (N_16561,N_12905,N_13453);
or U16562 (N_16562,N_14017,N_13360);
nor U16563 (N_16563,N_14144,N_14357);
nor U16564 (N_16564,N_14025,N_12590);
nor U16565 (N_16565,N_12573,N_14599);
nor U16566 (N_16566,N_12628,N_13801);
and U16567 (N_16567,N_13061,N_14526);
xor U16568 (N_16568,N_13627,N_14390);
nor U16569 (N_16569,N_13547,N_13942);
nand U16570 (N_16570,N_13030,N_13305);
and U16571 (N_16571,N_14458,N_14693);
and U16572 (N_16572,N_13045,N_14173);
or U16573 (N_16573,N_13975,N_13191);
nand U16574 (N_16574,N_12549,N_13919);
and U16575 (N_16575,N_12745,N_12604);
xnor U16576 (N_16576,N_14683,N_12966);
xor U16577 (N_16577,N_14919,N_14305);
nor U16578 (N_16578,N_12582,N_14963);
nor U16579 (N_16579,N_13259,N_13646);
or U16580 (N_16580,N_14736,N_13991);
xnor U16581 (N_16581,N_13387,N_14296);
or U16582 (N_16582,N_12684,N_14700);
and U16583 (N_16583,N_13135,N_14204);
nand U16584 (N_16584,N_13612,N_13844);
or U16585 (N_16585,N_13343,N_13295);
nor U16586 (N_16586,N_14084,N_13886);
xor U16587 (N_16587,N_12859,N_13555);
nor U16588 (N_16588,N_12748,N_14805);
nand U16589 (N_16589,N_14023,N_14383);
or U16590 (N_16590,N_14573,N_14119);
nor U16591 (N_16591,N_14288,N_14318);
nand U16592 (N_16592,N_14162,N_13596);
or U16593 (N_16593,N_13806,N_14318);
nor U16594 (N_16594,N_14256,N_13298);
nand U16595 (N_16595,N_14467,N_14387);
and U16596 (N_16596,N_14389,N_14453);
xnor U16597 (N_16597,N_13265,N_13662);
or U16598 (N_16598,N_13639,N_13877);
or U16599 (N_16599,N_13553,N_12859);
nand U16600 (N_16600,N_12901,N_14672);
nand U16601 (N_16601,N_14596,N_13932);
or U16602 (N_16602,N_12893,N_13725);
and U16603 (N_16603,N_13093,N_14045);
nor U16604 (N_16604,N_14271,N_13725);
nand U16605 (N_16605,N_12905,N_12558);
or U16606 (N_16606,N_12928,N_14988);
or U16607 (N_16607,N_14300,N_12637);
nor U16608 (N_16608,N_13025,N_14241);
or U16609 (N_16609,N_12908,N_14558);
xnor U16610 (N_16610,N_14200,N_13933);
xor U16611 (N_16611,N_13427,N_14431);
nor U16612 (N_16612,N_13612,N_12666);
and U16613 (N_16613,N_14102,N_14008);
or U16614 (N_16614,N_14670,N_14138);
or U16615 (N_16615,N_12550,N_13372);
nand U16616 (N_16616,N_14100,N_12996);
nand U16617 (N_16617,N_13252,N_14360);
or U16618 (N_16618,N_13776,N_13817);
nand U16619 (N_16619,N_13454,N_13644);
or U16620 (N_16620,N_12831,N_12586);
and U16621 (N_16621,N_14967,N_13921);
or U16622 (N_16622,N_14733,N_14809);
nand U16623 (N_16623,N_13855,N_12585);
nor U16624 (N_16624,N_14455,N_13990);
xnor U16625 (N_16625,N_12760,N_13131);
or U16626 (N_16626,N_12803,N_12831);
xor U16627 (N_16627,N_13170,N_13247);
xnor U16628 (N_16628,N_14567,N_13856);
xor U16629 (N_16629,N_13223,N_14851);
nand U16630 (N_16630,N_14792,N_13231);
and U16631 (N_16631,N_14572,N_13917);
and U16632 (N_16632,N_12881,N_13057);
and U16633 (N_16633,N_14063,N_14054);
nor U16634 (N_16634,N_13765,N_13751);
nand U16635 (N_16635,N_12766,N_14906);
or U16636 (N_16636,N_13885,N_12760);
nand U16637 (N_16637,N_13529,N_13187);
nor U16638 (N_16638,N_14669,N_14496);
or U16639 (N_16639,N_13276,N_14361);
or U16640 (N_16640,N_14127,N_14800);
or U16641 (N_16641,N_13801,N_14989);
xnor U16642 (N_16642,N_14429,N_14116);
nand U16643 (N_16643,N_13588,N_14761);
and U16644 (N_16644,N_14261,N_13892);
and U16645 (N_16645,N_13677,N_13247);
or U16646 (N_16646,N_12543,N_13189);
xor U16647 (N_16647,N_13962,N_14675);
or U16648 (N_16648,N_12788,N_13450);
and U16649 (N_16649,N_13478,N_13004);
or U16650 (N_16650,N_13251,N_12909);
or U16651 (N_16651,N_14281,N_14299);
nor U16652 (N_16652,N_14102,N_13670);
nand U16653 (N_16653,N_14408,N_13533);
nand U16654 (N_16654,N_14745,N_12606);
nor U16655 (N_16655,N_14600,N_13200);
nor U16656 (N_16656,N_14236,N_13124);
xor U16657 (N_16657,N_12790,N_12732);
nand U16658 (N_16658,N_12873,N_12654);
nand U16659 (N_16659,N_13695,N_13402);
or U16660 (N_16660,N_13387,N_13260);
or U16661 (N_16661,N_13176,N_14938);
nand U16662 (N_16662,N_12526,N_12966);
xnor U16663 (N_16663,N_13179,N_14891);
nor U16664 (N_16664,N_14417,N_14595);
and U16665 (N_16665,N_13408,N_12564);
nand U16666 (N_16666,N_14935,N_14933);
nand U16667 (N_16667,N_13549,N_13118);
and U16668 (N_16668,N_14682,N_12980);
or U16669 (N_16669,N_13607,N_14369);
nor U16670 (N_16670,N_12990,N_12872);
xnor U16671 (N_16671,N_13718,N_14480);
nand U16672 (N_16672,N_13409,N_13856);
xnor U16673 (N_16673,N_14047,N_13548);
nand U16674 (N_16674,N_14436,N_12744);
and U16675 (N_16675,N_12992,N_13946);
nand U16676 (N_16676,N_13399,N_13236);
or U16677 (N_16677,N_13751,N_14842);
or U16678 (N_16678,N_13090,N_13306);
xor U16679 (N_16679,N_13510,N_14954);
xnor U16680 (N_16680,N_12596,N_14821);
or U16681 (N_16681,N_13500,N_13743);
and U16682 (N_16682,N_14511,N_14377);
nand U16683 (N_16683,N_13075,N_12842);
and U16684 (N_16684,N_13443,N_12933);
or U16685 (N_16685,N_14351,N_13555);
xor U16686 (N_16686,N_14369,N_14402);
nor U16687 (N_16687,N_12945,N_13595);
nor U16688 (N_16688,N_14428,N_13137);
and U16689 (N_16689,N_12693,N_14510);
nor U16690 (N_16690,N_12657,N_12750);
and U16691 (N_16691,N_14185,N_13314);
nor U16692 (N_16692,N_13845,N_12614);
or U16693 (N_16693,N_14566,N_13743);
nand U16694 (N_16694,N_13002,N_14753);
xnor U16695 (N_16695,N_14677,N_12750);
nor U16696 (N_16696,N_14984,N_14140);
nand U16697 (N_16697,N_13910,N_14304);
nor U16698 (N_16698,N_12557,N_14406);
xor U16699 (N_16699,N_14005,N_13122);
nor U16700 (N_16700,N_12572,N_14960);
and U16701 (N_16701,N_13090,N_14351);
and U16702 (N_16702,N_13396,N_14209);
nor U16703 (N_16703,N_14627,N_14549);
nor U16704 (N_16704,N_14972,N_13806);
xnor U16705 (N_16705,N_13601,N_13130);
nor U16706 (N_16706,N_13143,N_14600);
nand U16707 (N_16707,N_13467,N_12739);
and U16708 (N_16708,N_13104,N_14380);
and U16709 (N_16709,N_13335,N_12653);
and U16710 (N_16710,N_14504,N_14322);
nand U16711 (N_16711,N_12719,N_14606);
xnor U16712 (N_16712,N_14160,N_13413);
or U16713 (N_16713,N_12743,N_13723);
or U16714 (N_16714,N_13111,N_13081);
and U16715 (N_16715,N_13225,N_12693);
nor U16716 (N_16716,N_13989,N_12972);
xor U16717 (N_16717,N_14050,N_14889);
nand U16718 (N_16718,N_12840,N_14663);
xor U16719 (N_16719,N_14286,N_14983);
nor U16720 (N_16720,N_12827,N_13717);
and U16721 (N_16721,N_12538,N_14691);
and U16722 (N_16722,N_14091,N_14489);
nor U16723 (N_16723,N_12813,N_12880);
and U16724 (N_16724,N_14275,N_14579);
nand U16725 (N_16725,N_13548,N_13809);
and U16726 (N_16726,N_14268,N_14577);
or U16727 (N_16727,N_13970,N_13373);
and U16728 (N_16728,N_14416,N_13808);
nor U16729 (N_16729,N_12529,N_14898);
nand U16730 (N_16730,N_13427,N_13934);
nor U16731 (N_16731,N_13109,N_14048);
nor U16732 (N_16732,N_14484,N_12947);
and U16733 (N_16733,N_14970,N_12660);
nor U16734 (N_16734,N_12755,N_13253);
xnor U16735 (N_16735,N_12852,N_14668);
xnor U16736 (N_16736,N_13116,N_13976);
nand U16737 (N_16737,N_13920,N_12870);
and U16738 (N_16738,N_13435,N_14596);
nor U16739 (N_16739,N_14474,N_14637);
or U16740 (N_16740,N_14013,N_12674);
nor U16741 (N_16741,N_12632,N_14083);
or U16742 (N_16742,N_14091,N_14428);
xnor U16743 (N_16743,N_13535,N_12964);
and U16744 (N_16744,N_13323,N_13339);
nor U16745 (N_16745,N_14443,N_12578);
nor U16746 (N_16746,N_12567,N_12818);
or U16747 (N_16747,N_13969,N_13321);
or U16748 (N_16748,N_13338,N_14616);
or U16749 (N_16749,N_13322,N_12795);
nor U16750 (N_16750,N_13933,N_13991);
xor U16751 (N_16751,N_13473,N_14890);
xnor U16752 (N_16752,N_14179,N_14354);
or U16753 (N_16753,N_13280,N_14754);
and U16754 (N_16754,N_14223,N_14883);
nor U16755 (N_16755,N_13911,N_13166);
and U16756 (N_16756,N_13618,N_13024);
nor U16757 (N_16757,N_14646,N_12766);
nor U16758 (N_16758,N_14216,N_13896);
and U16759 (N_16759,N_14320,N_14612);
or U16760 (N_16760,N_14156,N_14890);
nand U16761 (N_16761,N_13472,N_13701);
and U16762 (N_16762,N_13268,N_14690);
or U16763 (N_16763,N_13443,N_13078);
nand U16764 (N_16764,N_14632,N_13610);
and U16765 (N_16765,N_14005,N_14348);
xor U16766 (N_16766,N_14898,N_12970);
xor U16767 (N_16767,N_14064,N_13797);
nand U16768 (N_16768,N_12700,N_12554);
nand U16769 (N_16769,N_13000,N_12573);
nor U16770 (N_16770,N_14299,N_12759);
nand U16771 (N_16771,N_14823,N_13691);
nor U16772 (N_16772,N_14649,N_13413);
and U16773 (N_16773,N_12557,N_12861);
xor U16774 (N_16774,N_13765,N_14744);
nand U16775 (N_16775,N_13741,N_12745);
and U16776 (N_16776,N_13289,N_13200);
or U16777 (N_16777,N_13726,N_14153);
or U16778 (N_16778,N_14755,N_14889);
nor U16779 (N_16779,N_13430,N_12817);
or U16780 (N_16780,N_13351,N_14873);
and U16781 (N_16781,N_13604,N_14977);
and U16782 (N_16782,N_13510,N_14765);
and U16783 (N_16783,N_14283,N_14568);
and U16784 (N_16784,N_13903,N_12628);
or U16785 (N_16785,N_13977,N_12734);
or U16786 (N_16786,N_13682,N_14111);
or U16787 (N_16787,N_14991,N_14504);
nand U16788 (N_16788,N_13446,N_14273);
nand U16789 (N_16789,N_12657,N_13623);
and U16790 (N_16790,N_14164,N_14526);
and U16791 (N_16791,N_13804,N_12512);
nor U16792 (N_16792,N_13062,N_12886);
xor U16793 (N_16793,N_14037,N_14699);
and U16794 (N_16794,N_13586,N_14667);
xor U16795 (N_16795,N_13090,N_13897);
or U16796 (N_16796,N_14784,N_12723);
nand U16797 (N_16797,N_13208,N_14176);
nand U16798 (N_16798,N_13458,N_14706);
nand U16799 (N_16799,N_14994,N_13723);
xnor U16800 (N_16800,N_13772,N_14945);
and U16801 (N_16801,N_14837,N_12669);
xnor U16802 (N_16802,N_13425,N_12638);
nand U16803 (N_16803,N_14056,N_14747);
or U16804 (N_16804,N_12876,N_13084);
or U16805 (N_16805,N_13202,N_12685);
nor U16806 (N_16806,N_13718,N_13472);
nor U16807 (N_16807,N_14767,N_13765);
xor U16808 (N_16808,N_12755,N_14626);
xnor U16809 (N_16809,N_12956,N_14648);
nand U16810 (N_16810,N_13710,N_14980);
or U16811 (N_16811,N_14774,N_14258);
or U16812 (N_16812,N_13391,N_13802);
nor U16813 (N_16813,N_13790,N_14333);
nand U16814 (N_16814,N_14347,N_13730);
or U16815 (N_16815,N_14010,N_13786);
nand U16816 (N_16816,N_12617,N_14265);
nand U16817 (N_16817,N_12512,N_12840);
or U16818 (N_16818,N_13579,N_14701);
and U16819 (N_16819,N_14389,N_14951);
nor U16820 (N_16820,N_13014,N_14962);
nand U16821 (N_16821,N_13329,N_13713);
nand U16822 (N_16822,N_14793,N_13591);
xnor U16823 (N_16823,N_14790,N_12804);
nor U16824 (N_16824,N_12701,N_13515);
xnor U16825 (N_16825,N_13381,N_14644);
and U16826 (N_16826,N_14985,N_12523);
or U16827 (N_16827,N_13258,N_12548);
xnor U16828 (N_16828,N_14611,N_12662);
and U16829 (N_16829,N_12562,N_13893);
and U16830 (N_16830,N_13373,N_13932);
nor U16831 (N_16831,N_13235,N_14000);
or U16832 (N_16832,N_12611,N_13156);
xor U16833 (N_16833,N_14032,N_12665);
or U16834 (N_16834,N_13312,N_12535);
nor U16835 (N_16835,N_13855,N_14679);
nand U16836 (N_16836,N_14363,N_14506);
or U16837 (N_16837,N_14421,N_13805);
nor U16838 (N_16838,N_12826,N_14552);
and U16839 (N_16839,N_12957,N_14422);
xnor U16840 (N_16840,N_14392,N_13213);
or U16841 (N_16841,N_13318,N_12927);
nor U16842 (N_16842,N_13808,N_13475);
or U16843 (N_16843,N_14063,N_12882);
nor U16844 (N_16844,N_13337,N_14165);
nand U16845 (N_16845,N_12914,N_13373);
nor U16846 (N_16846,N_13637,N_13036);
or U16847 (N_16847,N_14667,N_14772);
nor U16848 (N_16848,N_12600,N_14809);
or U16849 (N_16849,N_13738,N_12734);
xnor U16850 (N_16850,N_12900,N_14668);
nor U16851 (N_16851,N_13744,N_12972);
nand U16852 (N_16852,N_13575,N_13896);
nand U16853 (N_16853,N_14005,N_14665);
or U16854 (N_16854,N_14778,N_13132);
or U16855 (N_16855,N_12628,N_14458);
and U16856 (N_16856,N_13508,N_14058);
nor U16857 (N_16857,N_13209,N_13336);
and U16858 (N_16858,N_14973,N_13362);
nor U16859 (N_16859,N_12939,N_14271);
or U16860 (N_16860,N_14643,N_13306);
nor U16861 (N_16861,N_13095,N_14315);
nor U16862 (N_16862,N_12852,N_14215);
nor U16863 (N_16863,N_13914,N_12653);
nand U16864 (N_16864,N_13960,N_13846);
and U16865 (N_16865,N_14437,N_13421);
or U16866 (N_16866,N_14908,N_14055);
nor U16867 (N_16867,N_14871,N_13594);
or U16868 (N_16868,N_14773,N_12991);
or U16869 (N_16869,N_14345,N_12551);
nand U16870 (N_16870,N_13903,N_14247);
nand U16871 (N_16871,N_12927,N_12699);
nor U16872 (N_16872,N_12761,N_14782);
nand U16873 (N_16873,N_14002,N_14691);
nor U16874 (N_16874,N_14657,N_12727);
and U16875 (N_16875,N_12759,N_14389);
xnor U16876 (N_16876,N_13519,N_14813);
nor U16877 (N_16877,N_12960,N_13679);
xnor U16878 (N_16878,N_14619,N_13615);
xnor U16879 (N_16879,N_13233,N_14053);
and U16880 (N_16880,N_13166,N_12955);
xnor U16881 (N_16881,N_12520,N_13081);
nand U16882 (N_16882,N_13615,N_12573);
xnor U16883 (N_16883,N_13754,N_13406);
or U16884 (N_16884,N_14568,N_14571);
xor U16885 (N_16885,N_13087,N_13361);
or U16886 (N_16886,N_13159,N_13934);
or U16887 (N_16887,N_14283,N_12787);
xnor U16888 (N_16888,N_13514,N_12748);
or U16889 (N_16889,N_13890,N_12516);
xnor U16890 (N_16890,N_13642,N_14336);
or U16891 (N_16891,N_14086,N_14790);
nor U16892 (N_16892,N_14274,N_13279);
nand U16893 (N_16893,N_13017,N_12844);
or U16894 (N_16894,N_13624,N_13925);
and U16895 (N_16895,N_13886,N_14630);
or U16896 (N_16896,N_14033,N_12872);
nand U16897 (N_16897,N_12849,N_14350);
nor U16898 (N_16898,N_14613,N_13406);
nand U16899 (N_16899,N_14101,N_14306);
or U16900 (N_16900,N_13510,N_13937);
nand U16901 (N_16901,N_12833,N_13096);
xnor U16902 (N_16902,N_12834,N_14419);
and U16903 (N_16903,N_12815,N_12748);
and U16904 (N_16904,N_14641,N_13477);
or U16905 (N_16905,N_13971,N_14680);
xnor U16906 (N_16906,N_14497,N_12927);
or U16907 (N_16907,N_12927,N_13326);
and U16908 (N_16908,N_13568,N_14553);
or U16909 (N_16909,N_13771,N_14336);
xor U16910 (N_16910,N_13480,N_14663);
nor U16911 (N_16911,N_13071,N_13666);
or U16912 (N_16912,N_14781,N_13445);
xnor U16913 (N_16913,N_14876,N_14796);
or U16914 (N_16914,N_13093,N_13686);
nand U16915 (N_16915,N_14926,N_12752);
nor U16916 (N_16916,N_14658,N_14453);
or U16917 (N_16917,N_14960,N_13258);
nor U16918 (N_16918,N_13970,N_13822);
nand U16919 (N_16919,N_12734,N_12743);
xor U16920 (N_16920,N_13529,N_12605);
or U16921 (N_16921,N_12849,N_13203);
nand U16922 (N_16922,N_14454,N_14911);
nor U16923 (N_16923,N_14020,N_14473);
nor U16924 (N_16924,N_14695,N_13652);
or U16925 (N_16925,N_13124,N_13519);
nand U16926 (N_16926,N_12828,N_14089);
or U16927 (N_16927,N_12809,N_13818);
nand U16928 (N_16928,N_14935,N_14748);
nor U16929 (N_16929,N_14074,N_14452);
nor U16930 (N_16930,N_13586,N_14241);
nand U16931 (N_16931,N_14090,N_13314);
nor U16932 (N_16932,N_12886,N_13456);
and U16933 (N_16933,N_13038,N_13651);
or U16934 (N_16934,N_14394,N_14876);
nor U16935 (N_16935,N_14962,N_13304);
and U16936 (N_16936,N_14069,N_14653);
xnor U16937 (N_16937,N_14721,N_13400);
and U16938 (N_16938,N_14757,N_14196);
and U16939 (N_16939,N_14217,N_13129);
or U16940 (N_16940,N_13472,N_14266);
nor U16941 (N_16941,N_14608,N_13515);
or U16942 (N_16942,N_13724,N_13623);
or U16943 (N_16943,N_13591,N_13936);
nand U16944 (N_16944,N_12689,N_13738);
nand U16945 (N_16945,N_12668,N_14773);
xor U16946 (N_16946,N_13925,N_13823);
and U16947 (N_16947,N_13571,N_13706);
xor U16948 (N_16948,N_14551,N_13892);
or U16949 (N_16949,N_12649,N_13571);
and U16950 (N_16950,N_12818,N_13372);
xnor U16951 (N_16951,N_13725,N_14666);
xor U16952 (N_16952,N_14409,N_14688);
or U16953 (N_16953,N_12557,N_13084);
and U16954 (N_16954,N_12815,N_13366);
xnor U16955 (N_16955,N_14382,N_13765);
or U16956 (N_16956,N_13542,N_14192);
nor U16957 (N_16957,N_14641,N_13236);
xnor U16958 (N_16958,N_14396,N_14207);
nor U16959 (N_16959,N_13673,N_14689);
and U16960 (N_16960,N_12724,N_14114);
xnor U16961 (N_16961,N_13181,N_12695);
and U16962 (N_16962,N_14711,N_14358);
xor U16963 (N_16963,N_14755,N_13555);
nor U16964 (N_16964,N_13227,N_13393);
or U16965 (N_16965,N_13520,N_12888);
or U16966 (N_16966,N_13387,N_13029);
nor U16967 (N_16967,N_12981,N_14829);
or U16968 (N_16968,N_12962,N_13449);
and U16969 (N_16969,N_14292,N_14135);
or U16970 (N_16970,N_13310,N_14001);
and U16971 (N_16971,N_14494,N_14750);
and U16972 (N_16972,N_14059,N_14812);
nor U16973 (N_16973,N_14671,N_12940);
nand U16974 (N_16974,N_12996,N_14210);
and U16975 (N_16975,N_13765,N_14240);
nor U16976 (N_16976,N_14356,N_13500);
xor U16977 (N_16977,N_12815,N_12692);
and U16978 (N_16978,N_13218,N_13472);
nor U16979 (N_16979,N_13549,N_14234);
nand U16980 (N_16980,N_14756,N_13732);
nand U16981 (N_16981,N_14161,N_14169);
or U16982 (N_16982,N_12581,N_14099);
and U16983 (N_16983,N_14776,N_13645);
nor U16984 (N_16984,N_12953,N_14187);
xnor U16985 (N_16985,N_12811,N_14818);
and U16986 (N_16986,N_14199,N_14192);
xnor U16987 (N_16987,N_13633,N_14029);
and U16988 (N_16988,N_14491,N_14758);
or U16989 (N_16989,N_14783,N_13840);
xor U16990 (N_16990,N_13538,N_14624);
nor U16991 (N_16991,N_14672,N_14251);
and U16992 (N_16992,N_14090,N_13076);
and U16993 (N_16993,N_13429,N_13301);
nand U16994 (N_16994,N_14228,N_13439);
or U16995 (N_16995,N_12990,N_13014);
and U16996 (N_16996,N_13367,N_12773);
or U16997 (N_16997,N_13303,N_13418);
and U16998 (N_16998,N_13651,N_13093);
and U16999 (N_16999,N_13054,N_14728);
or U17000 (N_17000,N_12722,N_14375);
nor U17001 (N_17001,N_13334,N_12855);
nand U17002 (N_17002,N_13713,N_13218);
or U17003 (N_17003,N_13105,N_12650);
xor U17004 (N_17004,N_13157,N_13092);
nand U17005 (N_17005,N_14456,N_14583);
xor U17006 (N_17006,N_14020,N_12554);
xor U17007 (N_17007,N_14301,N_13783);
and U17008 (N_17008,N_13879,N_13822);
xor U17009 (N_17009,N_14887,N_13776);
nor U17010 (N_17010,N_14845,N_12951);
xnor U17011 (N_17011,N_12782,N_12989);
or U17012 (N_17012,N_13746,N_14493);
nor U17013 (N_17013,N_14355,N_12835);
or U17014 (N_17014,N_12517,N_12930);
or U17015 (N_17015,N_14088,N_12824);
nand U17016 (N_17016,N_14715,N_13132);
xor U17017 (N_17017,N_14722,N_13035);
xnor U17018 (N_17018,N_12879,N_13910);
xor U17019 (N_17019,N_14181,N_14981);
and U17020 (N_17020,N_12994,N_12927);
or U17021 (N_17021,N_14796,N_12683);
xor U17022 (N_17022,N_13165,N_13060);
or U17023 (N_17023,N_14319,N_13957);
or U17024 (N_17024,N_13225,N_13976);
or U17025 (N_17025,N_14766,N_14003);
and U17026 (N_17026,N_13073,N_13621);
nor U17027 (N_17027,N_14989,N_14267);
and U17028 (N_17028,N_13789,N_14677);
xor U17029 (N_17029,N_12508,N_14597);
nor U17030 (N_17030,N_13736,N_14282);
or U17031 (N_17031,N_13752,N_14934);
or U17032 (N_17032,N_13698,N_13132);
nor U17033 (N_17033,N_12542,N_14241);
nand U17034 (N_17034,N_13500,N_13932);
nor U17035 (N_17035,N_13415,N_13390);
nor U17036 (N_17036,N_14466,N_14510);
xor U17037 (N_17037,N_13426,N_13642);
nor U17038 (N_17038,N_14920,N_14155);
nand U17039 (N_17039,N_13866,N_14344);
or U17040 (N_17040,N_14648,N_14708);
nand U17041 (N_17041,N_13285,N_12829);
xnor U17042 (N_17042,N_13209,N_14417);
and U17043 (N_17043,N_14822,N_14858);
xnor U17044 (N_17044,N_12828,N_13578);
or U17045 (N_17045,N_12670,N_14797);
nand U17046 (N_17046,N_14317,N_14011);
xor U17047 (N_17047,N_14595,N_13415);
nor U17048 (N_17048,N_13767,N_14233);
nand U17049 (N_17049,N_14225,N_13609);
nor U17050 (N_17050,N_12758,N_13245);
xor U17051 (N_17051,N_14584,N_12777);
nor U17052 (N_17052,N_14772,N_12989);
xor U17053 (N_17053,N_14704,N_13521);
or U17054 (N_17054,N_13217,N_14505);
and U17055 (N_17055,N_14672,N_13254);
nor U17056 (N_17056,N_14359,N_12573);
nor U17057 (N_17057,N_12506,N_12721);
nand U17058 (N_17058,N_14398,N_14109);
xnor U17059 (N_17059,N_12942,N_14502);
and U17060 (N_17060,N_13531,N_14885);
nand U17061 (N_17061,N_14488,N_14330);
nor U17062 (N_17062,N_13483,N_12893);
nand U17063 (N_17063,N_14401,N_13174);
and U17064 (N_17064,N_14479,N_12957);
nor U17065 (N_17065,N_14887,N_13006);
nand U17066 (N_17066,N_13566,N_12963);
xor U17067 (N_17067,N_13444,N_14008);
and U17068 (N_17068,N_14384,N_14698);
and U17069 (N_17069,N_13898,N_12613);
nor U17070 (N_17070,N_14622,N_14876);
nand U17071 (N_17071,N_14905,N_13861);
or U17072 (N_17072,N_12835,N_14324);
nor U17073 (N_17073,N_12841,N_14921);
and U17074 (N_17074,N_13703,N_12588);
nor U17075 (N_17075,N_13612,N_13262);
nor U17076 (N_17076,N_12809,N_13659);
or U17077 (N_17077,N_14951,N_13614);
and U17078 (N_17078,N_14241,N_14768);
xnor U17079 (N_17079,N_14715,N_13421);
nor U17080 (N_17080,N_12588,N_13890);
or U17081 (N_17081,N_14324,N_13587);
or U17082 (N_17082,N_13133,N_13869);
and U17083 (N_17083,N_12991,N_13482);
nor U17084 (N_17084,N_14979,N_12969);
xor U17085 (N_17085,N_14218,N_14553);
and U17086 (N_17086,N_14501,N_14983);
xor U17087 (N_17087,N_14983,N_13611);
xor U17088 (N_17088,N_13696,N_14514);
nand U17089 (N_17089,N_12972,N_14153);
or U17090 (N_17090,N_13763,N_14880);
and U17091 (N_17091,N_12721,N_13231);
nor U17092 (N_17092,N_12934,N_14294);
or U17093 (N_17093,N_14583,N_14107);
nand U17094 (N_17094,N_14535,N_13790);
nand U17095 (N_17095,N_14544,N_14351);
nand U17096 (N_17096,N_13931,N_13502);
nor U17097 (N_17097,N_14094,N_14431);
nand U17098 (N_17098,N_12928,N_13325);
xor U17099 (N_17099,N_14323,N_12649);
xor U17100 (N_17100,N_14643,N_13453);
or U17101 (N_17101,N_13281,N_14535);
nor U17102 (N_17102,N_13899,N_14494);
xor U17103 (N_17103,N_14857,N_12622);
and U17104 (N_17104,N_14597,N_14529);
nor U17105 (N_17105,N_14573,N_13463);
xor U17106 (N_17106,N_14156,N_14929);
nor U17107 (N_17107,N_13303,N_13018);
xor U17108 (N_17108,N_13179,N_13622);
and U17109 (N_17109,N_14890,N_13621);
nand U17110 (N_17110,N_14643,N_14998);
nor U17111 (N_17111,N_13555,N_12668);
xor U17112 (N_17112,N_14214,N_12833);
and U17113 (N_17113,N_14704,N_12673);
nor U17114 (N_17114,N_12596,N_13992);
nor U17115 (N_17115,N_12643,N_14920);
and U17116 (N_17116,N_13654,N_14555);
nand U17117 (N_17117,N_13679,N_14823);
nor U17118 (N_17118,N_13253,N_13985);
or U17119 (N_17119,N_14136,N_14289);
xnor U17120 (N_17120,N_14241,N_14994);
nor U17121 (N_17121,N_13871,N_13898);
and U17122 (N_17122,N_14325,N_12903);
and U17123 (N_17123,N_14109,N_14399);
nor U17124 (N_17124,N_13062,N_14913);
xnor U17125 (N_17125,N_12968,N_13938);
and U17126 (N_17126,N_12923,N_14962);
and U17127 (N_17127,N_13467,N_14187);
nor U17128 (N_17128,N_13351,N_13846);
or U17129 (N_17129,N_13650,N_14367);
nor U17130 (N_17130,N_12765,N_13990);
nand U17131 (N_17131,N_14146,N_12858);
or U17132 (N_17132,N_13247,N_14968);
and U17133 (N_17133,N_14360,N_13358);
xor U17134 (N_17134,N_14907,N_13374);
and U17135 (N_17135,N_13531,N_14492);
or U17136 (N_17136,N_14325,N_14345);
or U17137 (N_17137,N_12783,N_13540);
xnor U17138 (N_17138,N_14147,N_14769);
or U17139 (N_17139,N_14151,N_13149);
nand U17140 (N_17140,N_12561,N_13754);
and U17141 (N_17141,N_14022,N_14741);
xor U17142 (N_17142,N_12756,N_13585);
nor U17143 (N_17143,N_14236,N_14905);
nor U17144 (N_17144,N_13363,N_14392);
nor U17145 (N_17145,N_14807,N_14058);
xor U17146 (N_17146,N_13883,N_14272);
and U17147 (N_17147,N_12663,N_14012);
or U17148 (N_17148,N_14956,N_14662);
nand U17149 (N_17149,N_12817,N_13306);
and U17150 (N_17150,N_13154,N_14431);
nand U17151 (N_17151,N_14279,N_14506);
xnor U17152 (N_17152,N_14397,N_12601);
nand U17153 (N_17153,N_14912,N_13593);
and U17154 (N_17154,N_13733,N_12968);
nor U17155 (N_17155,N_14538,N_14050);
xor U17156 (N_17156,N_14714,N_12797);
nand U17157 (N_17157,N_14347,N_14944);
or U17158 (N_17158,N_12582,N_12724);
xnor U17159 (N_17159,N_12899,N_13410);
and U17160 (N_17160,N_14889,N_13796);
and U17161 (N_17161,N_14834,N_13793);
or U17162 (N_17162,N_12996,N_14058);
xnor U17163 (N_17163,N_14901,N_13308);
xor U17164 (N_17164,N_14175,N_13465);
nor U17165 (N_17165,N_13383,N_12889);
or U17166 (N_17166,N_12605,N_14310);
and U17167 (N_17167,N_13840,N_13848);
nor U17168 (N_17168,N_14791,N_13235);
nor U17169 (N_17169,N_14706,N_14963);
nor U17170 (N_17170,N_13866,N_14184);
xnor U17171 (N_17171,N_14939,N_13809);
nand U17172 (N_17172,N_13502,N_13499);
xor U17173 (N_17173,N_14722,N_13703);
or U17174 (N_17174,N_13782,N_14859);
nand U17175 (N_17175,N_13887,N_13330);
nand U17176 (N_17176,N_13744,N_14669);
nor U17177 (N_17177,N_13471,N_12984);
nand U17178 (N_17178,N_12690,N_14816);
nor U17179 (N_17179,N_12711,N_14191);
nor U17180 (N_17180,N_13706,N_13117);
or U17181 (N_17181,N_13626,N_13388);
or U17182 (N_17182,N_13925,N_14711);
or U17183 (N_17183,N_14136,N_14887);
nand U17184 (N_17184,N_14980,N_13064);
and U17185 (N_17185,N_13241,N_13051);
or U17186 (N_17186,N_13515,N_14789);
xor U17187 (N_17187,N_13690,N_12994);
and U17188 (N_17188,N_13214,N_13965);
nor U17189 (N_17189,N_13632,N_13945);
or U17190 (N_17190,N_14952,N_13192);
or U17191 (N_17191,N_14916,N_12893);
nand U17192 (N_17192,N_14785,N_14486);
xnor U17193 (N_17193,N_14337,N_13563);
and U17194 (N_17194,N_13007,N_14924);
and U17195 (N_17195,N_14622,N_13424);
xnor U17196 (N_17196,N_12588,N_14767);
or U17197 (N_17197,N_13424,N_12868);
nand U17198 (N_17198,N_14652,N_12500);
and U17199 (N_17199,N_14337,N_13790);
xor U17200 (N_17200,N_13909,N_14488);
nand U17201 (N_17201,N_14410,N_14160);
nor U17202 (N_17202,N_13075,N_12675);
or U17203 (N_17203,N_14248,N_14022);
and U17204 (N_17204,N_13938,N_13930);
or U17205 (N_17205,N_12991,N_12829);
nor U17206 (N_17206,N_13298,N_13675);
and U17207 (N_17207,N_12855,N_14939);
or U17208 (N_17208,N_12504,N_14985);
or U17209 (N_17209,N_14621,N_13404);
nor U17210 (N_17210,N_12517,N_13631);
nand U17211 (N_17211,N_14482,N_12564);
or U17212 (N_17212,N_12901,N_14577);
and U17213 (N_17213,N_14417,N_13609);
nand U17214 (N_17214,N_14506,N_13320);
or U17215 (N_17215,N_12643,N_13330);
or U17216 (N_17216,N_12934,N_13074);
nor U17217 (N_17217,N_13335,N_13448);
and U17218 (N_17218,N_14588,N_14622);
or U17219 (N_17219,N_14797,N_12704);
nand U17220 (N_17220,N_13827,N_14037);
nor U17221 (N_17221,N_13126,N_13651);
or U17222 (N_17222,N_13177,N_13792);
or U17223 (N_17223,N_14635,N_12552);
or U17224 (N_17224,N_12593,N_12941);
or U17225 (N_17225,N_13028,N_13464);
or U17226 (N_17226,N_14165,N_13155);
nor U17227 (N_17227,N_13533,N_14066);
nor U17228 (N_17228,N_14944,N_14611);
or U17229 (N_17229,N_13680,N_13344);
or U17230 (N_17230,N_14101,N_14689);
nand U17231 (N_17231,N_13090,N_12872);
or U17232 (N_17232,N_12893,N_14598);
nor U17233 (N_17233,N_13373,N_13350);
or U17234 (N_17234,N_14302,N_13008);
xnor U17235 (N_17235,N_13797,N_13769);
or U17236 (N_17236,N_14897,N_13735);
or U17237 (N_17237,N_13311,N_14588);
nor U17238 (N_17238,N_14692,N_13004);
nor U17239 (N_17239,N_13403,N_14984);
or U17240 (N_17240,N_12804,N_14834);
nor U17241 (N_17241,N_12963,N_12673);
xor U17242 (N_17242,N_12601,N_12696);
or U17243 (N_17243,N_12611,N_14044);
nand U17244 (N_17244,N_13854,N_13642);
and U17245 (N_17245,N_14551,N_14474);
nand U17246 (N_17246,N_12721,N_13410);
xor U17247 (N_17247,N_13194,N_12517);
and U17248 (N_17248,N_14259,N_14086);
nor U17249 (N_17249,N_13104,N_14063);
nand U17250 (N_17250,N_13482,N_14282);
nor U17251 (N_17251,N_12503,N_13192);
xor U17252 (N_17252,N_13951,N_14023);
nor U17253 (N_17253,N_13970,N_13165);
nor U17254 (N_17254,N_13319,N_13414);
and U17255 (N_17255,N_13464,N_13444);
nor U17256 (N_17256,N_13195,N_13026);
or U17257 (N_17257,N_14515,N_14516);
and U17258 (N_17258,N_14394,N_13208);
nand U17259 (N_17259,N_14632,N_12894);
xor U17260 (N_17260,N_13387,N_13332);
or U17261 (N_17261,N_14364,N_14783);
nor U17262 (N_17262,N_12635,N_13699);
nor U17263 (N_17263,N_12748,N_13004);
or U17264 (N_17264,N_14387,N_14133);
and U17265 (N_17265,N_14404,N_13865);
nand U17266 (N_17266,N_13436,N_13755);
nand U17267 (N_17267,N_14580,N_12692);
xor U17268 (N_17268,N_13338,N_14124);
nand U17269 (N_17269,N_13750,N_12996);
nor U17270 (N_17270,N_14636,N_14779);
nor U17271 (N_17271,N_14806,N_12611);
nor U17272 (N_17272,N_13851,N_13007);
nor U17273 (N_17273,N_14001,N_14306);
xnor U17274 (N_17274,N_12698,N_14801);
or U17275 (N_17275,N_12758,N_13590);
or U17276 (N_17276,N_14231,N_13741);
xor U17277 (N_17277,N_14249,N_13748);
nor U17278 (N_17278,N_13343,N_14844);
or U17279 (N_17279,N_12639,N_14415);
or U17280 (N_17280,N_14398,N_13790);
and U17281 (N_17281,N_14549,N_14676);
nor U17282 (N_17282,N_13170,N_13485);
and U17283 (N_17283,N_14048,N_14288);
nor U17284 (N_17284,N_14982,N_12963);
nor U17285 (N_17285,N_14828,N_14489);
nand U17286 (N_17286,N_14673,N_13403);
xor U17287 (N_17287,N_14680,N_14762);
or U17288 (N_17288,N_13484,N_13151);
xor U17289 (N_17289,N_12795,N_14059);
xor U17290 (N_17290,N_13074,N_14132);
or U17291 (N_17291,N_13482,N_13984);
or U17292 (N_17292,N_14745,N_14785);
or U17293 (N_17293,N_12567,N_14153);
and U17294 (N_17294,N_13760,N_13066);
nand U17295 (N_17295,N_13209,N_13521);
xor U17296 (N_17296,N_12977,N_14695);
nand U17297 (N_17297,N_14751,N_13424);
or U17298 (N_17298,N_13480,N_14179);
nor U17299 (N_17299,N_12560,N_14555);
and U17300 (N_17300,N_14913,N_12925);
xor U17301 (N_17301,N_14912,N_12914);
xor U17302 (N_17302,N_14481,N_14326);
xor U17303 (N_17303,N_13993,N_14451);
nor U17304 (N_17304,N_13529,N_14566);
or U17305 (N_17305,N_14290,N_13046);
xnor U17306 (N_17306,N_12842,N_13066);
or U17307 (N_17307,N_12742,N_14818);
nor U17308 (N_17308,N_13131,N_13159);
or U17309 (N_17309,N_13204,N_12507);
xnor U17310 (N_17310,N_12564,N_14640);
and U17311 (N_17311,N_13614,N_12570);
xnor U17312 (N_17312,N_13028,N_14397);
xnor U17313 (N_17313,N_13633,N_13314);
nand U17314 (N_17314,N_13460,N_14055);
xnor U17315 (N_17315,N_14788,N_13222);
and U17316 (N_17316,N_14134,N_14360);
or U17317 (N_17317,N_12564,N_13476);
xnor U17318 (N_17318,N_14766,N_12595);
nand U17319 (N_17319,N_13500,N_14888);
or U17320 (N_17320,N_14295,N_14198);
nor U17321 (N_17321,N_12875,N_14161);
or U17322 (N_17322,N_13656,N_13197);
nand U17323 (N_17323,N_13237,N_13207);
and U17324 (N_17324,N_14045,N_12710);
and U17325 (N_17325,N_12786,N_12964);
xor U17326 (N_17326,N_14764,N_13650);
nor U17327 (N_17327,N_13506,N_14795);
nand U17328 (N_17328,N_13060,N_14838);
or U17329 (N_17329,N_14827,N_12870);
nand U17330 (N_17330,N_14904,N_14565);
xnor U17331 (N_17331,N_14300,N_12988);
nand U17332 (N_17332,N_13725,N_14691);
or U17333 (N_17333,N_14373,N_12653);
nor U17334 (N_17334,N_14866,N_13297);
nand U17335 (N_17335,N_14566,N_13654);
and U17336 (N_17336,N_12791,N_12570);
nand U17337 (N_17337,N_14302,N_13251);
xnor U17338 (N_17338,N_13416,N_12980);
nand U17339 (N_17339,N_12697,N_14894);
xor U17340 (N_17340,N_13934,N_13333);
nor U17341 (N_17341,N_14749,N_12743);
nand U17342 (N_17342,N_14726,N_14654);
nor U17343 (N_17343,N_13990,N_14064);
or U17344 (N_17344,N_13398,N_13351);
nor U17345 (N_17345,N_13352,N_12763);
and U17346 (N_17346,N_14004,N_12750);
and U17347 (N_17347,N_14136,N_12588);
and U17348 (N_17348,N_14360,N_14551);
and U17349 (N_17349,N_14863,N_12948);
or U17350 (N_17350,N_13911,N_14332);
or U17351 (N_17351,N_13446,N_13562);
xnor U17352 (N_17352,N_13435,N_13906);
and U17353 (N_17353,N_14719,N_13081);
nor U17354 (N_17354,N_14515,N_14612);
and U17355 (N_17355,N_13908,N_14717);
xor U17356 (N_17356,N_14884,N_13504);
nand U17357 (N_17357,N_13475,N_12534);
and U17358 (N_17358,N_14064,N_13615);
nor U17359 (N_17359,N_14000,N_13475);
nor U17360 (N_17360,N_14140,N_14391);
nor U17361 (N_17361,N_12813,N_12916);
nor U17362 (N_17362,N_14989,N_14876);
nor U17363 (N_17363,N_14879,N_12853);
xor U17364 (N_17364,N_13438,N_14585);
nor U17365 (N_17365,N_13733,N_14486);
and U17366 (N_17366,N_13746,N_14670);
and U17367 (N_17367,N_13967,N_14106);
and U17368 (N_17368,N_14648,N_13615);
or U17369 (N_17369,N_12714,N_13769);
nor U17370 (N_17370,N_14877,N_14964);
nor U17371 (N_17371,N_13487,N_12720);
and U17372 (N_17372,N_13588,N_12749);
xor U17373 (N_17373,N_13848,N_12643);
or U17374 (N_17374,N_12580,N_14737);
or U17375 (N_17375,N_13218,N_14157);
xor U17376 (N_17376,N_13225,N_14381);
xnor U17377 (N_17377,N_14009,N_13043);
xor U17378 (N_17378,N_13204,N_13766);
xor U17379 (N_17379,N_14450,N_14192);
nand U17380 (N_17380,N_13577,N_14646);
xor U17381 (N_17381,N_13378,N_14015);
and U17382 (N_17382,N_12786,N_14347);
and U17383 (N_17383,N_14902,N_13662);
xor U17384 (N_17384,N_12795,N_12549);
or U17385 (N_17385,N_12932,N_12810);
or U17386 (N_17386,N_12624,N_14924);
nor U17387 (N_17387,N_13079,N_13477);
xor U17388 (N_17388,N_14458,N_14328);
xnor U17389 (N_17389,N_13830,N_14480);
or U17390 (N_17390,N_13892,N_13406);
xor U17391 (N_17391,N_12715,N_14560);
nor U17392 (N_17392,N_12760,N_14626);
xnor U17393 (N_17393,N_13848,N_14289);
nor U17394 (N_17394,N_13310,N_14052);
and U17395 (N_17395,N_12833,N_14675);
nand U17396 (N_17396,N_12886,N_13095);
nor U17397 (N_17397,N_13380,N_12841);
nor U17398 (N_17398,N_13085,N_14933);
or U17399 (N_17399,N_13743,N_14802);
nand U17400 (N_17400,N_13027,N_12830);
or U17401 (N_17401,N_12977,N_13317);
nand U17402 (N_17402,N_12887,N_13207);
or U17403 (N_17403,N_12820,N_14027);
nor U17404 (N_17404,N_14462,N_13202);
nand U17405 (N_17405,N_14504,N_12579);
and U17406 (N_17406,N_14352,N_14338);
and U17407 (N_17407,N_13148,N_12780);
and U17408 (N_17408,N_12923,N_14519);
xor U17409 (N_17409,N_14218,N_13781);
or U17410 (N_17410,N_13547,N_14163);
xnor U17411 (N_17411,N_13638,N_13517);
and U17412 (N_17412,N_14516,N_13563);
nor U17413 (N_17413,N_13098,N_13439);
nor U17414 (N_17414,N_14100,N_14024);
and U17415 (N_17415,N_14676,N_14202);
and U17416 (N_17416,N_14181,N_14493);
and U17417 (N_17417,N_12947,N_13732);
or U17418 (N_17418,N_14065,N_12921);
xnor U17419 (N_17419,N_13051,N_14645);
nor U17420 (N_17420,N_13591,N_12809);
or U17421 (N_17421,N_12594,N_14634);
or U17422 (N_17422,N_13486,N_12703);
or U17423 (N_17423,N_12916,N_14627);
nand U17424 (N_17424,N_14504,N_12887);
xnor U17425 (N_17425,N_14299,N_13949);
and U17426 (N_17426,N_13061,N_12624);
and U17427 (N_17427,N_13760,N_13796);
xnor U17428 (N_17428,N_12792,N_12794);
xor U17429 (N_17429,N_14108,N_14777);
nand U17430 (N_17430,N_14599,N_12975);
or U17431 (N_17431,N_13685,N_13778);
xor U17432 (N_17432,N_14416,N_14860);
or U17433 (N_17433,N_14593,N_14163);
nor U17434 (N_17434,N_14655,N_12889);
nor U17435 (N_17435,N_14508,N_13906);
xnor U17436 (N_17436,N_13614,N_13987);
nand U17437 (N_17437,N_12835,N_13030);
and U17438 (N_17438,N_14988,N_14365);
xor U17439 (N_17439,N_14636,N_13834);
xor U17440 (N_17440,N_13159,N_13084);
nor U17441 (N_17441,N_12958,N_13424);
nor U17442 (N_17442,N_13404,N_14174);
nand U17443 (N_17443,N_12847,N_14014);
or U17444 (N_17444,N_14748,N_14965);
xnor U17445 (N_17445,N_14695,N_14030);
nor U17446 (N_17446,N_12513,N_14422);
and U17447 (N_17447,N_14033,N_13689);
nor U17448 (N_17448,N_12950,N_12938);
nand U17449 (N_17449,N_14531,N_13693);
xnor U17450 (N_17450,N_14285,N_14259);
and U17451 (N_17451,N_14213,N_13105);
nand U17452 (N_17452,N_12873,N_12693);
nand U17453 (N_17453,N_13795,N_12786);
nor U17454 (N_17454,N_14071,N_13241);
nand U17455 (N_17455,N_14333,N_13005);
or U17456 (N_17456,N_12994,N_13253);
or U17457 (N_17457,N_13886,N_12962);
nor U17458 (N_17458,N_14109,N_13665);
xor U17459 (N_17459,N_13420,N_13926);
or U17460 (N_17460,N_13729,N_14286);
nor U17461 (N_17461,N_14442,N_14983);
xor U17462 (N_17462,N_13991,N_13417);
nor U17463 (N_17463,N_14634,N_14917);
and U17464 (N_17464,N_13753,N_13769);
and U17465 (N_17465,N_14598,N_12907);
or U17466 (N_17466,N_13902,N_14186);
nor U17467 (N_17467,N_14434,N_12841);
or U17468 (N_17468,N_14164,N_14821);
xor U17469 (N_17469,N_14925,N_12815);
xor U17470 (N_17470,N_13296,N_13752);
nor U17471 (N_17471,N_13576,N_12898);
and U17472 (N_17472,N_13259,N_13618);
xor U17473 (N_17473,N_13395,N_13590);
nor U17474 (N_17474,N_14563,N_14387);
and U17475 (N_17475,N_14719,N_13004);
nor U17476 (N_17476,N_12723,N_14733);
nor U17477 (N_17477,N_12657,N_13332);
or U17478 (N_17478,N_14038,N_12791);
or U17479 (N_17479,N_14462,N_12672);
nor U17480 (N_17480,N_14701,N_14695);
or U17481 (N_17481,N_12694,N_13396);
nand U17482 (N_17482,N_14891,N_12529);
nand U17483 (N_17483,N_13874,N_14108);
or U17484 (N_17484,N_14527,N_13691);
nor U17485 (N_17485,N_14438,N_14363);
xnor U17486 (N_17486,N_12680,N_14098);
and U17487 (N_17487,N_12670,N_13088);
nor U17488 (N_17488,N_13987,N_14900);
and U17489 (N_17489,N_12662,N_12919);
and U17490 (N_17490,N_13045,N_14542);
or U17491 (N_17491,N_14075,N_13979);
nor U17492 (N_17492,N_14795,N_13021);
nor U17493 (N_17493,N_14903,N_12629);
or U17494 (N_17494,N_13037,N_12591);
and U17495 (N_17495,N_14860,N_13064);
xnor U17496 (N_17496,N_12588,N_12682);
or U17497 (N_17497,N_13760,N_13197);
nand U17498 (N_17498,N_13070,N_13457);
nand U17499 (N_17499,N_13707,N_13525);
xor U17500 (N_17500,N_15114,N_16857);
nor U17501 (N_17501,N_16456,N_15587);
nand U17502 (N_17502,N_15345,N_16755);
xnor U17503 (N_17503,N_17373,N_17111);
and U17504 (N_17504,N_16869,N_16542);
nand U17505 (N_17505,N_17077,N_15096);
nor U17506 (N_17506,N_15915,N_16984);
nand U17507 (N_17507,N_15285,N_17451);
or U17508 (N_17508,N_17309,N_17032);
nand U17509 (N_17509,N_16180,N_17349);
or U17510 (N_17510,N_16322,N_16788);
nand U17511 (N_17511,N_15333,N_15657);
xnor U17512 (N_17512,N_15985,N_15842);
xnor U17513 (N_17513,N_16021,N_15250);
nand U17514 (N_17514,N_15197,N_15141);
nor U17515 (N_17515,N_16006,N_16162);
xnor U17516 (N_17516,N_16435,N_16175);
xor U17517 (N_17517,N_16752,N_17434);
nand U17518 (N_17518,N_16888,N_15660);
nand U17519 (N_17519,N_15936,N_16278);
and U17520 (N_17520,N_15737,N_15201);
nand U17521 (N_17521,N_17386,N_16813);
nor U17522 (N_17522,N_15779,N_17141);
or U17523 (N_17523,N_17448,N_15738);
and U17524 (N_17524,N_16467,N_15575);
or U17525 (N_17525,N_15110,N_17112);
nor U17526 (N_17526,N_16165,N_16604);
xnor U17527 (N_17527,N_15870,N_17353);
or U17528 (N_17528,N_15594,N_15055);
or U17529 (N_17529,N_15160,N_17043);
xnor U17530 (N_17530,N_15112,N_16818);
and U17531 (N_17531,N_17464,N_15360);
nand U17532 (N_17532,N_16645,N_16969);
nand U17533 (N_17533,N_15579,N_17154);
nor U17534 (N_17534,N_16938,N_16099);
xor U17535 (N_17535,N_15138,N_15644);
nand U17536 (N_17536,N_16035,N_15830);
nand U17537 (N_17537,N_17027,N_15322);
xnor U17538 (N_17538,N_15955,N_15121);
nand U17539 (N_17539,N_16141,N_16594);
nor U17540 (N_17540,N_15558,N_15663);
or U17541 (N_17541,N_15905,N_17136);
nand U17542 (N_17542,N_16854,N_16987);
nor U17543 (N_17543,N_15725,N_15307);
nor U17544 (N_17544,N_16220,N_16721);
and U17545 (N_17545,N_15109,N_16890);
or U17546 (N_17546,N_16269,N_17445);
or U17547 (N_17547,N_17406,N_16886);
nand U17548 (N_17548,N_16423,N_16091);
xor U17549 (N_17549,N_15811,N_16193);
and U17550 (N_17550,N_16921,N_16259);
and U17551 (N_17551,N_16308,N_15760);
xnor U17552 (N_17552,N_15396,N_15505);
or U17553 (N_17553,N_15962,N_15227);
xor U17554 (N_17554,N_16152,N_15045);
and U17555 (N_17555,N_16872,N_15065);
nor U17556 (N_17556,N_16319,N_17232);
xor U17557 (N_17557,N_15049,N_17355);
and U17558 (N_17558,N_15655,N_15762);
and U17559 (N_17559,N_17415,N_17170);
xnor U17560 (N_17560,N_16615,N_17130);
xnor U17561 (N_17561,N_15027,N_16253);
nand U17562 (N_17562,N_17281,N_15642);
nor U17563 (N_17563,N_17437,N_16312);
nand U17564 (N_17564,N_16727,N_15075);
xnor U17565 (N_17565,N_17085,N_15638);
xor U17566 (N_17566,N_16466,N_15826);
or U17567 (N_17567,N_15202,N_16017);
and U17568 (N_17568,N_15132,N_16908);
and U17569 (N_17569,N_16037,N_16298);
xnor U17570 (N_17570,N_16535,N_15422);
nand U17571 (N_17571,N_16765,N_16320);
nor U17572 (N_17572,N_16048,N_17225);
nand U17573 (N_17573,N_15679,N_17219);
and U17574 (N_17574,N_16602,N_15482);
nand U17575 (N_17575,N_16241,N_17041);
nor U17576 (N_17576,N_15091,N_15751);
nand U17577 (N_17577,N_15085,N_16211);
xnor U17578 (N_17578,N_15372,N_15494);
nand U17579 (N_17579,N_15390,N_17311);
nand U17580 (N_17580,N_15446,N_16365);
nand U17581 (N_17581,N_17082,N_16125);
nor U17582 (N_17582,N_16584,N_17006);
and U17583 (N_17583,N_17153,N_16380);
nand U17584 (N_17584,N_15637,N_16049);
xnor U17585 (N_17585,N_16787,N_15604);
and U17586 (N_17586,N_17275,N_16139);
and U17587 (N_17587,N_16889,N_15933);
xor U17588 (N_17588,N_17414,N_15219);
or U17589 (N_17589,N_15136,N_17326);
nor U17590 (N_17590,N_15078,N_17285);
nor U17591 (N_17591,N_16036,N_15692);
nand U17592 (N_17592,N_16541,N_15834);
or U17593 (N_17593,N_17402,N_15528);
or U17594 (N_17594,N_16407,N_15084);
and U17595 (N_17595,N_17139,N_16081);
nor U17596 (N_17596,N_16503,N_15016);
nor U17597 (N_17597,N_16360,N_15506);
xnor U17598 (N_17598,N_17120,N_16285);
xor U17599 (N_17599,N_16197,N_15032);
nand U17600 (N_17600,N_15081,N_17060);
xor U17601 (N_17601,N_17283,N_16323);
nor U17602 (N_17602,N_16714,N_15820);
nor U17603 (N_17603,N_15210,N_16116);
and U17604 (N_17604,N_16379,N_16935);
and U17605 (N_17605,N_15329,N_17103);
xor U17606 (N_17606,N_16279,N_16646);
and U17607 (N_17607,N_15626,N_16679);
nand U17608 (N_17608,N_15028,N_16949);
nor U17609 (N_17609,N_15220,N_16189);
and U17610 (N_17610,N_15546,N_16408);
nor U17611 (N_17611,N_16271,N_17185);
xor U17612 (N_17612,N_16309,N_17473);
nor U17613 (N_17613,N_16415,N_15563);
or U17614 (N_17614,N_16595,N_15847);
nor U17615 (N_17615,N_16354,N_16733);
xnor U17616 (N_17616,N_15861,N_15974);
xnor U17617 (N_17617,N_16839,N_16290);
nand U17618 (N_17618,N_16424,N_16482);
or U17619 (N_17619,N_17391,N_15810);
nand U17620 (N_17620,N_15560,N_17046);
or U17621 (N_17621,N_16807,N_15394);
nand U17622 (N_17622,N_15584,N_16851);
and U17623 (N_17623,N_17378,N_17234);
xnor U17624 (N_17624,N_17132,N_15204);
and U17625 (N_17625,N_15019,N_15559);
xor U17626 (N_17626,N_15901,N_15089);
and U17627 (N_17627,N_15806,N_16922);
xor U17628 (N_17628,N_16593,N_16633);
or U17629 (N_17629,N_15137,N_16459);
nand U17630 (N_17630,N_16896,N_16460);
nand U17631 (N_17631,N_15771,N_16563);
nand U17632 (N_17632,N_17038,N_17255);
nor U17633 (N_17633,N_15258,N_16891);
or U17634 (N_17634,N_17483,N_17004);
xor U17635 (N_17635,N_17229,N_16931);
and U17636 (N_17636,N_15023,N_17056);
or U17637 (N_17637,N_17007,N_15463);
and U17638 (N_17638,N_17020,N_16677);
and U17639 (N_17639,N_16668,N_16263);
nand U17640 (N_17640,N_16700,N_17357);
xnor U17641 (N_17641,N_16304,N_16486);
xnor U17642 (N_17642,N_15095,N_17408);
nor U17643 (N_17643,N_16628,N_16557);
and U17644 (N_17644,N_15489,N_15379);
xnor U17645 (N_17645,N_16723,N_17246);
and U17646 (N_17646,N_17293,N_16427);
nor U17647 (N_17647,N_16123,N_16893);
or U17648 (N_17648,N_15368,N_15367);
or U17649 (N_17649,N_15623,N_16800);
or U17650 (N_17650,N_17364,N_17013);
nand U17651 (N_17651,N_15425,N_15287);
xnor U17652 (N_17652,N_17145,N_16514);
nor U17653 (N_17653,N_17236,N_16485);
xnor U17654 (N_17654,N_16238,N_16926);
or U17655 (N_17655,N_15627,N_15274);
nor U17656 (N_17656,N_17097,N_15350);
xnor U17657 (N_17657,N_17023,N_17462);
and U17658 (N_17658,N_16117,N_16713);
nor U17659 (N_17659,N_16972,N_15851);
and U17660 (N_17660,N_17001,N_16270);
xor U17661 (N_17661,N_16823,N_16816);
nor U17662 (N_17662,N_15813,N_17290);
and U17663 (N_17663,N_17300,N_15491);
and U17664 (N_17664,N_15518,N_16169);
xnor U17665 (N_17665,N_17201,N_15158);
and U17666 (N_17666,N_16802,N_16112);
or U17667 (N_17667,N_16439,N_15526);
nor U17668 (N_17668,N_16578,N_15393);
xor U17669 (N_17669,N_15025,N_15540);
and U17670 (N_17670,N_16867,N_15514);
and U17671 (N_17671,N_17226,N_15195);
nand U17672 (N_17672,N_15495,N_16650);
or U17673 (N_17673,N_15297,N_17159);
or U17674 (N_17674,N_16338,N_15233);
nand U17675 (N_17675,N_15714,N_15880);
nand U17676 (N_17676,N_16256,N_15386);
or U17677 (N_17677,N_15914,N_15791);
nor U17678 (N_17678,N_15080,N_15606);
and U17679 (N_17679,N_16246,N_16096);
and U17680 (N_17680,N_15943,N_16284);
or U17681 (N_17681,N_15572,N_16585);
or U17682 (N_17682,N_16806,N_15739);
nand U17683 (N_17683,N_15823,N_15348);
or U17684 (N_17684,N_15866,N_16441);
xnor U17685 (N_17685,N_15513,N_15708);
xor U17686 (N_17686,N_16072,N_15062);
and U17687 (N_17687,N_16718,N_15459);
nand U17688 (N_17688,N_17323,N_16479);
nor U17689 (N_17689,N_15825,N_16778);
nand U17690 (N_17690,N_15485,N_15770);
nand U17691 (N_17691,N_17140,N_16781);
nor U17692 (N_17692,N_16392,N_16941);
and U17693 (N_17693,N_15289,N_15234);
nand U17694 (N_17694,N_17453,N_16501);
nor U17695 (N_17695,N_16341,N_16178);
nand U17696 (N_17696,N_16609,N_15592);
nand U17697 (N_17697,N_15254,N_15684);
or U17698 (N_17698,N_16487,N_15940);
and U17699 (N_17699,N_17029,N_15247);
nor U17700 (N_17700,N_15891,N_15599);
nand U17701 (N_17701,N_17352,N_15211);
xor U17702 (N_17702,N_17345,N_16237);
nor U17703 (N_17703,N_16145,N_17456);
nand U17704 (N_17704,N_15786,N_16862);
nand U17705 (N_17705,N_16745,N_17447);
and U17706 (N_17706,N_16107,N_17336);
xnor U17707 (N_17707,N_16590,N_15858);
or U17708 (N_17708,N_17274,N_16895);
nand U17709 (N_17709,N_17123,N_16143);
and U17710 (N_17710,N_17237,N_16881);
nor U17711 (N_17711,N_16129,N_16905);
nand U17712 (N_17712,N_16166,N_15403);
xnor U17713 (N_17713,N_16146,N_15843);
xnor U17714 (N_17714,N_16217,N_17129);
nor U17715 (N_17715,N_15266,N_16697);
nand U17716 (N_17716,N_16944,N_16717);
and U17717 (N_17717,N_16024,N_17147);
xnor U17718 (N_17718,N_17403,N_16383);
nand U17719 (N_17719,N_16075,N_15979);
nor U17720 (N_17720,N_16464,N_16042);
and U17721 (N_17721,N_15147,N_16251);
nand U17722 (N_17722,N_15787,N_15547);
or U17723 (N_17723,N_17121,N_17164);
xnor U17724 (N_17724,N_16950,N_16951);
and U17725 (N_17725,N_15719,N_15346);
or U17726 (N_17726,N_16527,N_16450);
xor U17727 (N_17727,N_16915,N_15310);
nor U17728 (N_17728,N_17273,N_15478);
and U17729 (N_17729,N_16254,N_17217);
and U17730 (N_17730,N_16977,N_17411);
nand U17731 (N_17731,N_15423,N_16437);
nor U17732 (N_17732,N_16030,N_16412);
nand U17733 (N_17733,N_16032,N_15500);
and U17734 (N_17734,N_16375,N_15789);
xnor U17735 (N_17735,N_17054,N_15057);
nand U17736 (N_17736,N_16119,N_17190);
nor U17737 (N_17737,N_15166,N_16385);
or U17738 (N_17738,N_17035,N_16328);
or U17739 (N_17739,N_15508,N_15869);
and U17740 (N_17740,N_16429,N_15522);
xor U17741 (N_17741,N_17288,N_16316);
or U17742 (N_17742,N_15864,N_17436);
nand U17743 (N_17743,N_15716,N_16704);
or U17744 (N_17744,N_15315,N_16496);
and U17745 (N_17745,N_16793,N_15300);
or U17746 (N_17746,N_16043,N_15410);
and U17747 (N_17747,N_15126,N_15570);
xnor U17748 (N_17748,N_15596,N_15941);
or U17749 (N_17749,N_15180,N_15653);
xor U17750 (N_17750,N_17016,N_17148);
or U17751 (N_17751,N_17396,N_15853);
nand U17752 (N_17752,N_16586,N_16734);
nor U17753 (N_17753,N_15288,N_16177);
and U17754 (N_17754,N_16127,N_15377);
xor U17755 (N_17755,N_17152,N_15595);
and U17756 (N_17756,N_16000,N_17160);
and U17757 (N_17757,N_17475,N_17157);
nand U17758 (N_17758,N_16780,N_17215);
nor U17759 (N_17759,N_15070,N_16769);
xor U17760 (N_17760,N_16952,N_16834);
and U17761 (N_17761,N_16350,N_17051);
nand U17762 (N_17762,N_15785,N_16689);
nor U17763 (N_17763,N_16861,N_16027);
nand U17764 (N_17764,N_16157,N_16906);
and U17765 (N_17765,N_15142,N_16920);
nand U17766 (N_17766,N_15292,N_15082);
and U17767 (N_17767,N_16858,N_17156);
xor U17768 (N_17768,N_15324,N_16605);
nor U17769 (N_17769,N_15406,N_16786);
nor U17770 (N_17770,N_17360,N_16826);
or U17771 (N_17771,N_15535,N_15688);
nor U17772 (N_17772,N_15854,N_15928);
nor U17773 (N_17773,N_16832,N_15117);
and U17774 (N_17774,N_16314,N_16986);
or U17775 (N_17775,N_15959,N_16004);
nor U17776 (N_17776,N_16104,N_16885);
nor U17777 (N_17777,N_17096,N_17099);
nor U17778 (N_17778,N_16489,N_17481);
or U17779 (N_17779,N_17252,N_16856);
and U17780 (N_17780,N_15800,N_17337);
xor U17781 (N_17781,N_16685,N_17238);
xnor U17782 (N_17782,N_17176,N_16443);
xnor U17783 (N_17783,N_16465,N_15305);
xnor U17784 (N_17784,N_15252,N_16184);
and U17785 (N_17785,N_16364,N_16968);
nand U17786 (N_17786,N_15389,N_16933);
xnor U17787 (N_17787,N_15715,N_15251);
nand U17788 (N_17788,N_15387,N_17346);
nor U17789 (N_17789,N_15674,N_17074);
xor U17790 (N_17790,N_17224,N_16965);
nor U17791 (N_17791,N_17241,N_15337);
nor U17792 (N_17792,N_16821,N_16850);
or U17793 (N_17793,N_16369,N_16919);
nor U17794 (N_17794,N_15051,N_17287);
or U17795 (N_17795,N_16639,N_17119);
nor U17796 (N_17796,N_16398,N_16871);
nand U17797 (N_17797,N_15946,N_15646);
or U17798 (N_17798,N_17491,N_17421);
nor U17799 (N_17799,N_16453,N_16286);
xnor U17800 (N_17800,N_17486,N_16671);
nor U17801 (N_17801,N_16601,N_15256);
xor U17802 (N_17802,N_16789,N_15614);
xnor U17803 (N_17803,N_15897,N_17179);
xnor U17804 (N_17804,N_15354,N_17429);
nand U17805 (N_17805,N_15037,N_15334);
xor U17806 (N_17806,N_17089,N_17459);
nor U17807 (N_17807,N_15629,N_15601);
or U17808 (N_17808,N_16661,N_15246);
and U17809 (N_17809,N_15699,N_16608);
or U17810 (N_17810,N_15910,N_15531);
nor U17811 (N_17811,N_17265,N_15989);
xnor U17812 (N_17812,N_16451,N_16618);
nand U17813 (N_17813,N_16015,N_16221);
nor U17814 (N_17814,N_16702,N_15349);
xnor U17815 (N_17815,N_15371,N_16273);
and U17816 (N_17816,N_15012,N_16698);
xnor U17817 (N_17817,N_16522,N_15155);
xor U17818 (N_17818,N_16653,N_15454);
nor U17819 (N_17819,N_16229,N_15743);
and U17820 (N_17820,N_15146,N_16554);
and U17821 (N_17821,N_17422,N_17369);
nor U17822 (N_17822,N_16736,N_16811);
xnor U17823 (N_17823,N_15544,N_15701);
xor U17824 (N_17824,N_16452,N_16695);
nand U17825 (N_17825,N_17435,N_16321);
nor U17826 (N_17826,N_15471,N_15903);
nand U17827 (N_17827,N_17316,N_15192);
or U17828 (N_17828,N_16331,N_15115);
nand U17829 (N_17829,N_15404,N_15239);
nand U17830 (N_17830,N_16946,N_15432);
or U17831 (N_17831,N_16636,N_17222);
nand U17832 (N_17832,N_16924,N_17375);
and U17833 (N_17833,N_15949,N_15819);
and U17834 (N_17834,N_17042,N_16582);
nand U17835 (N_17835,N_15024,N_17178);
xor U17836 (N_17836,N_15436,N_15460);
or U17837 (N_17837,N_16232,N_16957);
xor U17838 (N_17838,N_16534,N_16829);
nor U17839 (N_17839,N_17173,N_15186);
or U17840 (N_17840,N_17271,N_15932);
or U17841 (N_17841,N_17499,N_16840);
xnor U17842 (N_17842,N_17183,N_15302);
nor U17843 (N_17843,N_17117,N_15600);
xnor U17844 (N_17844,N_15470,N_16327);
and U17845 (N_17845,N_15484,N_17034);
and U17846 (N_17846,N_16822,N_15122);
or U17847 (N_17847,N_15286,N_16100);
and U17848 (N_17848,N_15170,N_15278);
nor U17849 (N_17849,N_16266,N_15273);
nand U17850 (N_17850,N_16703,N_15898);
or U17851 (N_17851,N_15036,N_16070);
nor U17852 (N_17852,N_16190,N_17227);
xnor U17853 (N_17853,N_15061,N_16690);
nor U17854 (N_17854,N_16206,N_17480);
nand U17855 (N_17855,N_15198,N_17008);
nand U17856 (N_17856,N_15174,N_17066);
xnor U17857 (N_17857,N_16518,N_15444);
nand U17858 (N_17858,N_16902,N_17494);
nor U17859 (N_17859,N_15217,N_16025);
or U17860 (N_17860,N_16577,N_15776);
and U17861 (N_17861,N_15295,N_17412);
nor U17862 (N_17862,N_17258,N_16934);
xor U17863 (N_17863,N_16838,N_16962);
and U17864 (N_17864,N_16059,N_17317);
or U17865 (N_17865,N_15822,N_17484);
and U17866 (N_17866,N_16726,N_17325);
nor U17867 (N_17867,N_15413,N_15968);
or U17868 (N_17868,N_17167,N_15257);
and U17869 (N_17869,N_15647,N_16167);
or U17870 (N_17870,N_15009,N_17488);
nor U17871 (N_17871,N_15691,N_15863);
and U17872 (N_17872,N_16124,N_15352);
xor U17873 (N_17873,N_15682,N_17014);
nand U17874 (N_17874,N_17377,N_17211);
nor U17875 (N_17875,N_15995,N_16900);
or U17876 (N_17876,N_15149,N_16046);
or U17877 (N_17877,N_15712,N_16366);
and U17878 (N_17878,N_16979,N_17151);
nand U17879 (N_17879,N_15038,N_17363);
nand U17880 (N_17880,N_17101,N_15721);
and U17881 (N_17881,N_17301,N_16550);
or U17882 (N_17882,N_16108,N_16200);
xnor U17883 (N_17883,N_16672,N_16475);
nor U17884 (N_17884,N_16997,N_15886);
xor U17885 (N_17885,N_16357,N_16057);
xor U17886 (N_17886,N_17230,N_17278);
nor U17887 (N_17887,N_15841,N_15942);
nand U17888 (N_17888,N_15022,N_17127);
nand U17889 (N_17889,N_15060,N_16208);
or U17890 (N_17890,N_16864,N_16681);
nand U17891 (N_17891,N_17022,N_16612);
or U17892 (N_17892,N_15235,N_17228);
and U17893 (N_17893,N_16034,N_15002);
and U17894 (N_17894,N_16186,N_15568);
nor U17895 (N_17895,N_15792,N_16028);
or U17896 (N_17896,N_16343,N_17142);
nand U17897 (N_17897,N_16521,N_16376);
nor U17898 (N_17898,N_17306,N_17387);
nand U17899 (N_17899,N_17181,N_15976);
nor U17900 (N_17900,N_16159,N_16095);
and U17901 (N_17901,N_15705,N_16627);
xnor U17902 (N_17902,N_15336,N_17410);
nor U17903 (N_17903,N_15958,N_16447);
nor U17904 (N_17904,N_17417,N_15885);
xor U17905 (N_17905,N_15734,N_16791);
nor U17906 (N_17906,N_16022,N_16461);
nor U17907 (N_17907,N_15686,N_15151);
xnor U17908 (N_17908,N_15607,N_16611);
nand U17909 (N_17909,N_16973,N_15578);
and U17910 (N_17910,N_16824,N_16288);
or U17911 (N_17911,N_15502,N_16433);
xor U17912 (N_17912,N_17404,N_15669);
or U17913 (N_17913,N_17482,N_16842);
nand U17914 (N_17914,N_16775,N_16102);
xor U17915 (N_17915,N_16892,N_16710);
xnor U17916 (N_17916,N_15145,N_16711);
nor U17917 (N_17917,N_15732,N_15123);
or U17918 (N_17918,N_15380,N_16976);
xnor U17919 (N_17919,N_16654,N_15862);
or U17920 (N_17920,N_15581,N_16005);
nand U17921 (N_17921,N_16648,N_17400);
or U17922 (N_17922,N_16658,N_16236);
or U17923 (N_17923,N_16402,N_17394);
xor U17924 (N_17924,N_16656,N_15753);
xnor U17925 (N_17925,N_15929,N_16137);
nor U17926 (N_17926,N_17084,N_15681);
nand U17927 (N_17927,N_16675,N_15630);
or U17928 (N_17928,N_15722,N_15282);
xor U17929 (N_17929,N_16820,N_16192);
nand U17930 (N_17930,N_15479,N_17188);
nor U17931 (N_17931,N_16085,N_15152);
nand U17932 (N_17932,N_16242,N_15812);
nand U17933 (N_17933,N_16738,N_15097);
xor U17934 (N_17934,N_16060,N_16230);
xor U17935 (N_17935,N_16548,N_16634);
nand U17936 (N_17936,N_16937,N_15215);
or U17937 (N_17937,N_16324,N_16086);
xnor U17938 (N_17938,N_16796,N_17118);
nand U17939 (N_17939,N_17088,N_16448);
and U17940 (N_17940,N_16912,N_15611);
and U17941 (N_17941,N_16699,N_15986);
and U17942 (N_17942,N_16373,N_17460);
or U17943 (N_17943,N_16771,N_17338);
xor U17944 (N_17944,N_15887,N_16568);
and U17945 (N_17945,N_16744,N_15244);
nand U17946 (N_17946,N_15745,N_15496);
or U17947 (N_17947,N_17455,N_15838);
xnor U17948 (N_17948,N_16347,N_16349);
xor U17949 (N_17949,N_17155,N_16458);
nor U17950 (N_17950,N_15969,N_15047);
and U17951 (N_17951,N_16898,N_17045);
nand U17952 (N_17952,N_15649,N_16047);
or U17953 (N_17953,N_17284,N_15018);
or U17954 (N_17954,N_16911,N_16914);
nor U17955 (N_17955,N_16927,N_17427);
or U17956 (N_17956,N_15311,N_16153);
or U17957 (N_17957,N_17202,N_16442);
or U17958 (N_17958,N_15778,N_16272);
nand U17959 (N_17959,N_16436,N_16089);
nand U17960 (N_17960,N_15279,N_15978);
xor U17961 (N_17961,N_17262,N_15951);
or U17962 (N_17962,N_17182,N_16363);
or U17963 (N_17963,N_15397,N_16449);
nand U17964 (N_17964,N_15654,N_15855);
nand U17965 (N_17965,N_16945,N_15856);
nor U17966 (N_17966,N_16434,N_16613);
and U17967 (N_17967,N_16071,N_15179);
or U17968 (N_17968,N_15103,N_15992);
nor U17969 (N_17969,N_15439,N_15005);
nor U17970 (N_17970,N_16795,N_15678);
nand U17971 (N_17971,N_15181,N_15748);
nand U17972 (N_17972,N_16133,N_15620);
nor U17973 (N_17973,N_17005,N_15537);
nor U17974 (N_17974,N_17327,N_17187);
and U17975 (N_17975,N_16989,N_17413);
and U17976 (N_17976,N_15269,N_16670);
nor U17977 (N_17977,N_16731,N_17026);
xnor U17978 (N_17978,N_15996,N_15066);
nor U17979 (N_17979,N_17244,N_15010);
and U17980 (N_17980,N_15556,N_15249);
nor U17981 (N_17981,N_16852,N_16039);
nand U17982 (N_17982,N_17296,N_16170);
nand U17983 (N_17983,N_15799,N_16262);
nand U17984 (N_17984,N_17247,N_16079);
xnor U17985 (N_17985,N_15063,N_15475);
xnor U17986 (N_17986,N_17419,N_16362);
and U17987 (N_17987,N_17389,N_17175);
xor U17988 (N_17988,N_17115,N_16708);
nand U17989 (N_17989,N_15670,N_15782);
or U17990 (N_17990,N_16728,N_15172);
xor U17991 (N_17991,N_17266,N_16985);
nor U17992 (N_17992,N_17367,N_17385);
nand U17993 (N_17993,N_15395,N_17302);
and U17994 (N_17994,N_16746,N_17191);
and U17995 (N_17995,N_16879,N_15481);
and U17996 (N_17996,N_15793,N_16399);
and U17997 (N_17997,N_17002,N_17490);
or U17998 (N_17998,N_15476,N_16110);
or U17999 (N_17999,N_16488,N_16940);
nand U18000 (N_18000,N_17276,N_17206);
nor U18001 (N_18001,N_17242,N_17478);
and U18002 (N_18002,N_15816,N_16883);
and U18003 (N_18003,N_15418,N_15327);
and U18004 (N_18004,N_17442,N_16239);
or U18005 (N_18005,N_15902,N_15453);
nor U18006 (N_18006,N_17295,N_15183);
nor U18007 (N_18007,N_17270,N_16388);
xnor U18008 (N_18008,N_15173,N_16377);
or U18009 (N_18009,N_16478,N_16344);
nand U18010 (N_18010,N_15450,N_16226);
xor U18011 (N_18011,N_15860,N_16396);
or U18012 (N_18012,N_15884,N_15366);
or U18013 (N_18013,N_16828,N_16201);
and U18014 (N_18014,N_15904,N_15298);
and U18015 (N_18015,N_17465,N_15157);
or U18016 (N_18016,N_16983,N_16614);
or U18017 (N_18017,N_15923,N_16836);
and U18018 (N_18018,N_16735,N_15991);
and U18019 (N_18019,N_16353,N_16764);
nor U18020 (N_18020,N_16228,N_15190);
and U18021 (N_18021,N_15056,N_17347);
or U18022 (N_18022,N_16052,N_15736);
nand U18023 (N_18023,N_15467,N_17383);
and U18024 (N_18024,N_16662,N_16497);
xnor U18025 (N_18025,N_16480,N_16549);
and U18026 (N_18026,N_15230,N_17371);
or U18027 (N_18027,N_17365,N_15919);
nand U18028 (N_18028,N_16674,N_17312);
or U18029 (N_18029,N_17090,N_16748);
nand U18030 (N_18030,N_15321,N_16421);
or U18031 (N_18031,N_16995,N_16154);
or U18032 (N_18032,N_16664,N_15375);
xnor U18033 (N_18033,N_16761,N_16430);
or U18034 (N_18034,N_17070,N_16843);
and U18035 (N_18035,N_15385,N_17033);
and U18036 (N_18036,N_15083,N_15775);
xnor U18037 (N_18037,N_16457,N_17072);
xor U18038 (N_18038,N_15156,N_15550);
or U18039 (N_18039,N_16663,N_16757);
xor U18040 (N_18040,N_15261,N_15048);
or U18041 (N_18041,N_17418,N_16741);
nand U18042 (N_18042,N_17291,N_16552);
and U18043 (N_18043,N_16596,N_16195);
xor U18044 (N_18044,N_15845,N_15392);
xnor U18045 (N_18045,N_16569,N_15086);
nand U18046 (N_18046,N_15445,N_15947);
xor U18047 (N_18047,N_17116,N_16964);
or U18048 (N_18048,N_15882,N_17231);
nand U18049 (N_18049,N_16432,N_16469);
and U18050 (N_18050,N_16652,N_15320);
and U18051 (N_18051,N_16260,N_16659);
and U18052 (N_18052,N_15237,N_16367);
and U18053 (N_18053,N_17286,N_16382);
nand U18054 (N_18054,N_17315,N_17304);
and U18055 (N_18055,N_16188,N_17313);
nor U18056 (N_18056,N_16610,N_17405);
or U18057 (N_18057,N_16164,N_16546);
xnor U18058 (N_18058,N_15415,N_16932);
nor U18059 (N_18059,N_16754,N_16676);
xnor U18060 (N_18060,N_17319,N_16198);
xor U18061 (N_18061,N_17095,N_16352);
nand U18062 (N_18062,N_17233,N_15074);
or U18063 (N_18063,N_16887,N_17197);
nand U18064 (N_18064,N_17376,N_15409);
and U18065 (N_18065,N_15740,N_16499);
and U18066 (N_18066,N_15645,N_16406);
and U18067 (N_18067,N_15788,N_15488);
and U18068 (N_18068,N_16848,N_15163);
and U18069 (N_18069,N_16815,N_15814);
nand U18070 (N_18070,N_16841,N_15666);
or U18071 (N_18071,N_17209,N_16084);
or U18072 (N_18072,N_15378,N_16874);
or U18073 (N_18073,N_15232,N_15301);
and U18074 (N_18074,N_16812,N_15007);
nor U18075 (N_18075,N_16058,N_15411);
and U18076 (N_18076,N_15402,N_16389);
and U18077 (N_18077,N_15621,N_16606);
or U18078 (N_18078,N_16556,N_16445);
and U18079 (N_18079,N_17407,N_16307);
or U18080 (N_18080,N_17184,N_15135);
and U18081 (N_18081,N_17441,N_15175);
and U18082 (N_18082,N_16547,N_16318);
nor U18083 (N_18083,N_15583,N_16939);
or U18084 (N_18084,N_15212,N_16740);
nand U18085 (N_18085,N_15591,N_15507);
xor U18086 (N_18086,N_16783,N_17091);
xnor U18087 (N_18087,N_16245,N_15171);
and U18088 (N_18088,N_16073,N_16067);
and U18089 (N_18089,N_16240,N_16054);
and U18090 (N_18090,N_16884,N_16023);
and U18091 (N_18091,N_15930,N_15588);
xor U18092 (N_18092,N_15128,N_16287);
and U18093 (N_18093,N_16991,N_16346);
or U18094 (N_18094,N_17093,N_16008);
nor U18095 (N_18095,N_15801,N_15765);
nor U18096 (N_18096,N_15718,N_15275);
xor U18097 (N_18097,N_17277,N_15006);
or U18098 (N_18098,N_15291,N_16719);
or U18099 (N_18099,N_15076,N_16144);
or U18100 (N_18100,N_16277,N_16468);
nand U18101 (N_18101,N_16515,N_16132);
nor U18102 (N_18102,N_16562,N_17279);
or U18103 (N_18103,N_15104,N_16589);
and U18104 (N_18104,N_16218,N_15248);
or U18105 (N_18105,N_16345,N_17489);
or U18106 (N_18106,N_17370,N_15150);
xnor U18107 (N_18107,N_17053,N_15658);
and U18108 (N_18108,N_15631,N_15031);
xnor U18109 (N_18109,N_16340,N_15807);
and U18110 (N_18110,N_16386,N_15199);
nor U18111 (N_18111,N_15664,N_17398);
nand U18112 (N_18112,N_16974,N_16016);
nor U18113 (N_18113,N_16739,N_17059);
or U18114 (N_18114,N_17021,N_16065);
nor U18115 (N_18115,N_15824,N_16657);
or U18116 (N_18116,N_15213,N_16250);
and U18117 (N_18117,N_17134,N_15222);
nand U18118 (N_18118,N_17372,N_16916);
and U18119 (N_18119,N_15447,N_16525);
or U18120 (N_18120,N_17133,N_17498);
nand U18121 (N_18121,N_16329,N_15340);
nand U18122 (N_18122,N_15519,N_17358);
or U18123 (N_18123,N_15652,N_17298);
and U18124 (N_18124,N_15304,N_16326);
nor U18125 (N_18125,N_15742,N_16474);
and U18126 (N_18126,N_16173,N_16929);
nor U18127 (N_18127,N_15837,N_17049);
nor U18128 (N_18128,N_16798,N_16302);
or U18129 (N_18129,N_15040,N_16640);
or U18130 (N_18130,N_15464,N_17107);
xor U18131 (N_18131,N_16255,N_15878);
nand U18132 (N_18132,N_16624,N_16830);
and U18133 (N_18133,N_15127,N_15408);
xor U18134 (N_18134,N_16289,N_16140);
or U18135 (N_18135,N_17495,N_17163);
and U18136 (N_18136,N_15921,N_15827);
nand U18137 (N_18137,N_17069,N_16538);
or U18138 (N_18138,N_17292,N_16476);
or U18139 (N_18139,N_16234,N_15566);
or U18140 (N_18140,N_15993,N_16910);
nor U18141 (N_18141,N_15729,N_16859);
nand U18142 (N_18142,N_15984,N_15981);
xor U18143 (N_18143,N_15803,N_15900);
nor U18144 (N_18144,N_17479,N_15306);
or U18145 (N_18145,N_17261,N_15303);
and U18146 (N_18146,N_15685,N_15939);
or U18147 (N_18147,N_15609,N_15746);
and U18148 (N_18148,N_16923,N_17094);
nand U18149 (N_18149,N_15209,N_15935);
or U18150 (N_18150,N_16492,N_16975);
xnor U18151 (N_18151,N_15576,N_17012);
or U18152 (N_18152,N_15512,N_15029);
xor U18153 (N_18153,N_15214,N_15690);
nand U18154 (N_18154,N_17039,N_17189);
nor U18155 (N_18155,N_16053,N_16160);
nor U18156 (N_18156,N_16092,N_16371);
nand U18157 (N_18157,N_17324,N_15758);
nand U18158 (N_18158,N_16870,N_15427);
xnor U18159 (N_18159,N_16111,N_15353);
xor U18160 (N_18160,N_15033,N_15613);
xor U18161 (N_18161,N_15755,N_17024);
nor U18162 (N_18162,N_17220,N_15262);
xnor U18163 (N_18163,N_16899,N_15308);
xor U18164 (N_18164,N_15131,N_17472);
or U18165 (N_18165,N_15696,N_17048);
nand U18166 (N_18166,N_15809,N_15892);
and U18167 (N_18167,N_16413,N_15835);
nor U18168 (N_18168,N_15004,N_15477);
and U18169 (N_18169,N_15907,N_16438);
xnor U18170 (N_18170,N_17263,N_16425);
and U18171 (N_18171,N_15756,N_16694);
and U18172 (N_18172,N_16209,N_17332);
xor U18173 (N_18173,N_16730,N_16794);
and U18174 (N_18174,N_15064,N_16384);
or U18175 (N_18175,N_17204,N_15724);
nand U18176 (N_18176,N_16422,N_16519);
and U18177 (N_18177,N_15185,N_15293);
and U18178 (N_18178,N_15922,N_15543);
and U18179 (N_18179,N_16630,N_16325);
or U18180 (N_18180,N_15990,N_15723);
nor U18181 (N_18181,N_17443,N_16512);
nor U18182 (N_18182,N_15087,N_16958);
nor U18183 (N_18183,N_16770,N_15757);
xor U18184 (N_18184,N_16580,N_15693);
nand U18185 (N_18185,N_15373,N_16419);
xnor U18186 (N_18186,N_17424,N_16227);
nor U18187 (N_18187,N_16358,N_16930);
xnor U18188 (N_18188,N_15088,N_15442);
and U18189 (N_18189,N_15918,N_15133);
and U18190 (N_18190,N_16115,N_15603);
and U18191 (N_18191,N_15499,N_15164);
xor U18192 (N_18192,N_17487,N_17073);
nand U18193 (N_18193,N_17063,N_16526);
and U18194 (N_18194,N_16790,N_15804);
nand U18195 (N_18195,N_15967,N_15309);
or U18196 (N_18196,N_15960,N_16007);
nor U18197 (N_18197,N_15384,N_15998);
or U18198 (N_18198,N_15077,N_16833);
or U18199 (N_18199,N_16196,N_16484);
or U18200 (N_18200,N_16504,N_15342);
nor U18201 (N_18201,N_16720,N_15597);
or U18202 (N_18202,N_16295,N_16093);
nand U18203 (N_18203,N_16147,N_16351);
and U18204 (N_18204,N_15511,N_16943);
or U18205 (N_18205,N_15177,N_16051);
nand U18206 (N_18206,N_15982,N_15548);
nand U18207 (N_18207,N_15313,N_15881);
xor U18208 (N_18208,N_15802,N_16971);
xor U18209 (N_18209,N_16077,N_15399);
xor U18210 (N_18210,N_15909,N_17199);
or U18211 (N_18211,N_16641,N_15521);
nand U18212 (N_18212,N_15351,N_17492);
nand U18213 (N_18213,N_15069,N_16638);
and U18214 (N_18214,N_16626,N_15977);
and U18215 (N_18215,N_15053,N_15364);
xor U18216 (N_18216,N_15831,N_17444);
nand U18217 (N_18217,N_16101,N_16715);
xor U18218 (N_18218,N_16768,N_17477);
nand U18219 (N_18219,N_17458,N_16135);
or U18220 (N_18220,N_15972,N_15105);
xor U18221 (N_18221,N_16498,N_17433);
and U18222 (N_18222,N_16961,N_15332);
nand U18223 (N_18223,N_15529,N_15365);
and U18224 (N_18224,N_16774,N_16873);
nand U18225 (N_18225,N_16583,N_16172);
nor U18226 (N_18226,N_16248,N_15245);
or U18227 (N_18227,N_15317,N_15675);
and U18228 (N_18228,N_16216,N_16026);
and U18229 (N_18229,N_16559,N_16076);
xnor U18230 (N_18230,N_15358,N_15781);
nor U18231 (N_18231,N_17052,N_16665);
xnor U18232 (N_18232,N_16809,N_15797);
or U18233 (N_18233,N_16050,N_16330);
nor U18234 (N_18234,N_17259,N_15871);
xnor U18235 (N_18235,N_15593,N_17485);
xnor U18236 (N_18236,N_17137,N_15424);
or U18237 (N_18237,N_17131,N_16574);
nor U18238 (N_18238,N_15253,N_15356);
and U18239 (N_18239,N_15720,N_15330);
or U18240 (N_18240,N_16517,N_16155);
xor U18241 (N_18241,N_15948,N_17339);
and U18242 (N_18242,N_16743,N_16019);
xnor U18243 (N_18243,N_17216,N_16565);
xor U18244 (N_18244,N_16183,N_17098);
or U18245 (N_18245,N_17469,N_16001);
or U18246 (N_18246,N_16481,N_16913);
nand U18247 (N_18247,N_15619,N_15046);
or U18248 (N_18248,N_16683,N_16179);
xor U18249 (N_18249,N_16729,N_15226);
or U18250 (N_18250,N_16428,N_15148);
nand U18251 (N_18251,N_16212,N_15280);
and U18252 (N_18252,N_16773,N_16126);
and U18253 (N_18253,N_17177,N_15341);
xnor U18254 (N_18254,N_15120,N_16342);
xnor U18255 (N_18255,N_15773,N_16235);
or U18256 (N_18256,N_16909,N_15795);
and U18257 (N_18257,N_17210,N_15677);
or U18258 (N_18258,N_17340,N_17196);
and U18259 (N_18259,N_15735,N_16477);
nor U18260 (N_18260,N_16374,N_16540);
nand U18261 (N_18261,N_15938,N_15178);
nand U18262 (N_18262,N_16252,N_16692);
nor U18263 (N_18263,N_15218,N_15107);
and U18264 (N_18264,N_16082,N_16558);
xnor U18265 (N_18265,N_15920,N_15168);
or U18266 (N_18266,N_15963,N_16105);
nor U18267 (N_18267,N_16925,N_15059);
or U18268 (N_18268,N_16960,N_15651);
xor U18269 (N_18269,N_15347,N_15836);
or U18270 (N_18270,N_16516,N_16805);
or U18271 (N_18271,N_16333,N_15916);
nor U18272 (N_18272,N_16524,N_15925);
nand U18273 (N_18273,N_16576,N_17162);
nor U18274 (N_18274,N_17212,N_15533);
xor U18275 (N_18275,N_16121,N_17461);
xnor U18276 (N_18276,N_16956,N_17168);
or U18277 (N_18277,N_15428,N_16470);
and U18278 (N_18278,N_15510,N_17254);
and U18279 (N_18279,N_16564,N_16426);
nand U18280 (N_18280,N_16296,N_16543);
nor U18281 (N_18281,N_17354,N_17331);
nand U18282 (N_18282,N_16303,N_16061);
nor U18283 (N_18283,N_15983,N_17100);
nand U18284 (N_18284,N_17205,N_16215);
nor U18285 (N_18285,N_15462,N_15102);
xnor U18286 (N_18286,N_16660,N_16222);
xor U18287 (N_18287,N_15888,N_15487);
xnor U18288 (N_18288,N_16010,N_16894);
or U18289 (N_18289,N_15430,N_16106);
nand U18290 (N_18290,N_16410,N_16495);
or U18291 (N_18291,N_15931,N_17009);
nor U18292 (N_18292,N_17062,N_16756);
and U18293 (N_18293,N_16598,N_16098);
nand U18294 (N_18294,N_15893,N_15616);
xnor U18295 (N_18295,N_16174,N_15412);
xnor U18296 (N_18296,N_17174,N_15267);
nand U18297 (N_18297,N_15957,N_17018);
or U18298 (N_18298,N_17392,N_17025);
and U18299 (N_18299,N_16018,N_15469);
and U18300 (N_18300,N_16693,N_15182);
xor U18301 (N_18301,N_15839,N_16844);
or U18302 (N_18302,N_15296,N_17390);
and U18303 (N_18303,N_15176,N_16520);
or U18304 (N_18304,N_16507,N_16356);
and U18305 (N_18305,N_16122,N_17067);
nand U18306 (N_18306,N_16163,N_16825);
and U18307 (N_18307,N_15749,N_16249);
nor U18308 (N_18308,N_16033,N_17235);
and U18309 (N_18309,N_16876,N_16142);
or U18310 (N_18310,N_15515,N_17036);
nor U18311 (N_18311,N_15759,N_15265);
or U18312 (N_18312,N_17470,N_15073);
and U18313 (N_18313,N_16336,N_16064);
nand U18314 (N_18314,N_15574,N_16572);
and U18315 (N_18315,N_15090,N_17430);
xnor U18316 (N_18316,N_16758,N_17080);
or U18317 (N_18317,N_17068,N_15255);
nor U18318 (N_18318,N_15727,N_16397);
nand U18319 (N_18319,N_16214,N_15221);
nor U18320 (N_18320,N_15874,N_15896);
nand U18321 (N_18321,N_16903,N_17047);
nand U18322 (N_18322,N_16532,N_16510);
nor U18323 (N_18323,N_16313,N_15554);
xnor U18324 (N_18324,N_17446,N_15608);
nand U18325 (N_18325,N_16138,N_17310);
nor U18326 (N_18326,N_16575,N_16394);
and U18327 (N_18327,N_15790,N_15857);
nor U18328 (N_18328,N_15325,N_15710);
xor U18329 (N_18329,N_15585,N_16651);
xor U18330 (N_18330,N_16090,N_15706);
xor U18331 (N_18331,N_17158,N_15093);
xnor U18332 (N_18332,N_17333,N_15865);
nand U18333 (N_18333,N_15945,N_15501);
and U18334 (N_18334,N_16182,N_16531);
nor U18335 (N_18335,N_15101,N_16666);
nor U18336 (N_18336,N_15035,N_16267);
xnor U18337 (N_18337,N_16801,N_16264);
xor U18338 (N_18338,N_15702,N_17251);
xnor U18339 (N_18339,N_16868,N_17065);
and U18340 (N_18340,N_16629,N_16300);
nor U18341 (N_18341,N_17348,N_15612);
nor U18342 (N_18342,N_15894,N_15707);
or U18343 (N_18343,N_15433,N_17108);
and U18344 (N_18344,N_16947,N_15971);
and U18345 (N_18345,N_17264,N_16310);
xnor U18346 (N_18346,N_16203,N_15465);
nand U18347 (N_18347,N_16505,N_17146);
nor U18348 (N_18348,N_16491,N_15001);
nor U18349 (N_18349,N_15844,N_17128);
xor U18350 (N_18350,N_15414,N_15589);
nand U18351 (N_18351,N_17423,N_15094);
xor U18352 (N_18352,N_16118,N_17268);
xor U18353 (N_18353,N_17463,N_16616);
nor U18354 (N_18354,N_15242,N_17388);
xor U18355 (N_18355,N_15763,N_16390);
nand U18356 (N_18356,N_15331,N_16337);
and U18357 (N_18357,N_16877,N_15420);
or U18358 (N_18358,N_16709,N_15208);
and U18359 (N_18359,N_17454,N_15486);
and U18360 (N_18360,N_17439,N_15161);
nor U18361 (N_18361,N_16387,N_15668);
nor U18362 (N_18362,N_17218,N_17109);
nand U18363 (N_18363,N_15400,N_15270);
or U18364 (N_18364,N_15357,N_16642);
nand U18365 (N_18365,N_16643,N_15241);
xnor U18366 (N_18366,N_16980,N_16202);
or U18367 (N_18367,N_16305,N_17037);
and U18368 (N_18368,N_15294,N_15525);
or U18369 (N_18369,N_16233,N_15238);
nand U18370 (N_18370,N_15119,N_15697);
and U18371 (N_18371,N_15632,N_16620);
or U18372 (N_18372,N_16530,N_15798);
nand U18373 (N_18373,N_17030,N_16391);
nand U18374 (N_18374,N_15975,N_16462);
or U18375 (N_18375,N_16268,N_16409);
xnor U18376 (N_18376,N_16539,N_15189);
xnor U18377 (N_18377,N_17113,N_15867);
and U18378 (N_18378,N_17476,N_17076);
xor U18379 (N_18379,N_16223,N_15276);
nor U18380 (N_18380,N_17169,N_16701);
nand U18381 (N_18381,N_16607,N_15586);
xnor U18382 (N_18382,N_15683,N_15665);
or U18383 (N_18383,N_16959,N_16224);
nor U18384 (N_18384,N_16291,N_16705);
nand U18385 (N_18385,N_16523,N_16803);
nor U18386 (N_18386,N_16282,N_16359);
nand U18387 (N_18387,N_16038,N_15796);
xnor U18388 (N_18388,N_16767,N_15054);
and U18389 (N_18389,N_16083,N_15987);
nand U18390 (N_18390,N_16866,N_16785);
or U18391 (N_18391,N_16749,N_16835);
and U18392 (N_18392,N_16536,N_15689);
xnor U18393 (N_18393,N_15536,N_15391);
nor U18394 (N_18394,N_16213,N_16131);
nand U18395 (N_18395,N_17497,N_17044);
nand U18396 (N_18396,N_16667,N_16444);
xor U18397 (N_18397,N_16545,N_15079);
nor U18398 (N_18398,N_17150,N_15573);
nor U18399 (N_18399,N_15376,N_15316);
or U18400 (N_18400,N_16265,N_16204);
or U18401 (N_18401,N_15106,N_15713);
and U18402 (N_18402,N_17350,N_15567);
nor U18403 (N_18403,N_16103,N_16561);
nor U18404 (N_18404,N_15997,N_15188);
and U18405 (N_18405,N_17249,N_15553);
xnor U18406 (N_18406,N_16827,N_17381);
nor U18407 (N_18407,N_16632,N_16617);
xnor U18408 (N_18408,N_15448,N_15490);
nand U18409 (N_18409,N_17384,N_17399);
or U18410 (N_18410,N_16918,N_15338);
nor U18411 (N_18411,N_17214,N_15184);
nand U18412 (N_18412,N_17194,N_16551);
or U18413 (N_18413,N_15667,N_15369);
and U18414 (N_18414,N_16724,N_15873);
or U18415 (N_18415,N_16281,N_17240);
nor U18416 (N_18416,N_16772,N_16134);
nor U18417 (N_18417,N_16882,N_17195);
nand U18418 (N_18418,N_16990,N_15206);
and U18419 (N_18419,N_16483,N_17071);
and U18420 (N_18420,N_15774,N_15162);
xnor U18421 (N_18421,N_16982,N_15000);
nand U18422 (N_18422,N_15961,N_17314);
nand U18423 (N_18423,N_15140,N_17087);
or U18424 (N_18424,N_15988,N_15440);
nor U18425 (N_18425,N_16055,N_15020);
xnor U18426 (N_18426,N_17409,N_15362);
nand U18427 (N_18427,N_16691,N_16506);
xnor U18428 (N_18428,N_15980,N_15026);
or U18429 (N_18429,N_16080,N_15312);
or U18430 (N_18430,N_16114,N_15846);
nor U18431 (N_18431,N_15200,N_15615);
or U18432 (N_18432,N_16381,N_15203);
nor U18433 (N_18433,N_16431,N_17078);
nor U18434 (N_18434,N_15268,N_15937);
xnor U18435 (N_18435,N_16243,N_16306);
or U18436 (N_18436,N_15924,N_17193);
nand U18437 (N_18437,N_16647,N_16258);
xor U18438 (N_18438,N_15769,N_16579);
nand U18439 (N_18439,N_17341,N_16591);
or U18440 (N_18440,N_16404,N_16760);
or U18441 (N_18441,N_15466,N_15504);
and U18442 (N_18442,N_16276,N_15118);
and U18443 (N_18443,N_15225,N_17061);
xor U18444 (N_18444,N_16777,N_17468);
nand U18445 (N_18445,N_16688,N_15405);
nor U18446 (N_18446,N_15849,N_16014);
or U18447 (N_18447,N_15565,N_15361);
xnor U18448 (N_18448,N_15196,N_16109);
nor U18449 (N_18449,N_17471,N_17368);
and U18450 (N_18450,N_15299,N_15965);
or U18451 (N_18451,N_16455,N_16509);
and U18452 (N_18452,N_16837,N_16649);
and U18453 (N_18453,N_15767,N_15580);
nand U18454 (N_18454,N_16274,N_16753);
xnor U18455 (N_18455,N_16401,N_16751);
and U18456 (N_18456,N_15747,N_15523);
nor U18457 (N_18457,N_17294,N_15875);
nor U18458 (N_18458,N_15872,N_15744);
xnor U18459 (N_18459,N_16571,N_15058);
nor U18460 (N_18460,N_16395,N_15549);
and U18461 (N_18461,N_17297,N_17299);
xnor U18462 (N_18462,N_16472,N_16560);
nand U18463 (N_18463,N_17031,N_16567);
nand U18464 (N_18464,N_15625,N_16766);
nor U18465 (N_18465,N_17125,N_16040);
nor U18466 (N_18466,N_17165,N_17428);
and U18467 (N_18467,N_15562,N_15072);
xnor U18468 (N_18468,N_17393,N_15455);
or U18469 (N_18469,N_15129,N_15134);
nor U18470 (N_18470,N_16420,N_16471);
nand U18471 (N_18471,N_16797,N_17200);
or U18472 (N_18472,N_16370,N_15355);
nor U18473 (N_18473,N_15374,N_15954);
nand U18474 (N_18474,N_16041,N_15633);
xnor U18475 (N_18475,N_17305,N_15534);
nand U18476 (N_18476,N_15449,N_17028);
nand U18477 (N_18477,N_15021,N_15461);
and U18478 (N_18478,N_16181,N_16623);
nand U18479 (N_18479,N_16597,N_17303);
or U18480 (N_18480,N_17431,N_15532);
xor U18481 (N_18481,N_15640,N_15452);
and U18482 (N_18482,N_15551,N_17450);
or U18483 (N_18483,N_16631,N_16191);
and U18484 (N_18484,N_16257,N_15318);
nand U18485 (N_18485,N_16194,N_15236);
and U18486 (N_18486,N_15895,N_16031);
xnor U18487 (N_18487,N_15794,N_15913);
or U18488 (N_18488,N_15343,N_16368);
nor U18489 (N_18489,N_17104,N_16493);
xor U18490 (N_18490,N_16600,N_16074);
and U18491 (N_18491,N_17267,N_15165);
nand U18492 (N_18492,N_16592,N_16292);
or U18493 (N_18493,N_17343,N_16168);
or U18494 (N_18494,N_17452,N_15741);
and U18495 (N_18495,N_16732,N_17203);
and U18496 (N_18496,N_16002,N_17359);
and U18497 (N_18497,N_15557,N_15434);
and U18498 (N_18498,N_16999,N_17086);
xnor U18499 (N_18499,N_17135,N_15610);
nand U18500 (N_18500,N_16348,N_17366);
and U18501 (N_18501,N_15950,N_15877);
nand U18502 (N_18502,N_15071,N_15833);
xnor U18503 (N_18503,N_15228,N_16494);
or U18504 (N_18504,N_16418,N_17379);
and U18505 (N_18505,N_17143,N_15260);
xnor U18506 (N_18506,N_15545,N_16393);
and U18507 (N_18507,N_15144,N_15509);
or U18508 (N_18508,N_17017,N_15205);
nor U18509 (N_18509,N_15429,N_16247);
and U18510 (N_18510,N_16062,N_16417);
and U18511 (N_18511,N_17064,N_15711);
and U18512 (N_18512,N_17208,N_15326);
xor U18513 (N_18513,N_15750,N_15700);
or U18514 (N_18514,N_15098,N_15290);
nand U18515 (N_18515,N_15398,N_15457);
or U18516 (N_18516,N_15473,N_16151);
or U18517 (N_18517,N_16553,N_15973);
xor U18518 (N_18518,N_15890,N_15635);
and U18519 (N_18519,N_16762,N_15416);
nand U18520 (N_18520,N_15264,N_16622);
xor U18521 (N_18521,N_15956,N_17198);
nor U18522 (N_18522,N_15671,N_16625);
or U18523 (N_18523,N_15636,N_16317);
or U18524 (N_18524,N_17050,N_15703);
xor U18525 (N_18525,N_16148,N_17401);
nor U18526 (N_18526,N_17382,N_17260);
nor U18527 (N_18527,N_15966,N_17320);
or U18528 (N_18528,N_15100,N_16996);
nand U18529 (N_18529,N_17496,N_16120);
nand U18530 (N_18530,N_16414,N_15003);
nor U18531 (N_18531,N_15130,N_16936);
or U18532 (N_18532,N_15590,N_17328);
nor U18533 (N_18533,N_17245,N_15879);
xnor U18534 (N_18534,N_17321,N_16161);
and U18535 (N_18535,N_16948,N_15493);
and U18536 (N_18536,N_15694,N_17280);
xnor U18537 (N_18537,N_16853,N_15552);
xor U18538 (N_18538,N_17166,N_17344);
and U18539 (N_18539,N_16339,N_15229);
xnor U18540 (N_18540,N_17186,N_15704);
nand U18541 (N_18541,N_16068,N_15474);
nand U18542 (N_18542,N_15883,N_17282);
nand U18543 (N_18543,N_15008,N_17466);
nor U18544 (N_18544,N_16463,N_15443);
or U18545 (N_18545,N_15994,N_17329);
nor U18546 (N_18546,N_15382,N_15498);
nor U18547 (N_18547,N_16297,N_16513);
nor U18548 (N_18548,N_17192,N_17243);
and U18549 (N_18549,N_16275,N_15673);
xor U18550 (N_18550,N_17272,N_16722);
nor U18551 (N_18551,N_16716,N_16637);
nor U18552 (N_18552,N_17213,N_17356);
nor U18553 (N_18553,N_16207,N_15431);
and U18554 (N_18554,N_17342,N_15030);
or U18555 (N_18555,N_15927,N_16372);
and U18556 (N_18556,N_16810,N_16814);
and U18557 (N_18557,N_15363,N_16817);
nor U18558 (N_18558,N_15876,N_15661);
or U18559 (N_18559,N_15821,N_15271);
nor U18560 (N_18560,N_16669,N_15314);
nor U18561 (N_18561,N_15656,N_16782);
nand U18562 (N_18562,N_17257,N_15730);
xnor U18563 (N_18563,N_17015,N_17426);
or U18564 (N_18564,N_17172,N_15569);
nor U18565 (N_18565,N_15780,N_15628);
and U18566 (N_18566,N_15272,N_15999);
or U18567 (N_18567,N_15648,N_15014);
and U18568 (N_18568,N_16907,N_15015);
nor U18569 (N_18569,N_16500,N_16044);
nand U18570 (N_18570,N_15908,N_15926);
or U18571 (N_18571,N_16011,N_16063);
nor U18572 (N_18572,N_17420,N_15541);
nor U18573 (N_18573,N_15840,N_16742);
and U18574 (N_18574,N_17083,N_16725);
or U18575 (N_18575,N_15154,N_16511);
nand U18576 (N_18576,N_16747,N_15125);
nor U18577 (N_18577,N_15634,N_15911);
or U18578 (N_18578,N_16334,N_15124);
or U18579 (N_18579,N_15828,N_17248);
or U18580 (N_18580,N_16587,N_16846);
nand U18581 (N_18581,N_15817,N_15754);
nor U18582 (N_18582,N_17010,N_15243);
or U18583 (N_18583,N_15944,N_17144);
or U18584 (N_18584,N_15970,N_15344);
nand U18585 (N_18585,N_15456,N_15764);
xor U18586 (N_18586,N_17362,N_16779);
or U18587 (N_18587,N_16130,N_15042);
nor U18588 (N_18588,N_16655,N_16069);
and U18589 (N_18589,N_17361,N_15153);
and U18590 (N_18590,N_15783,N_16544);
nand U18591 (N_18591,N_16988,N_16897);
and U18592 (N_18592,N_17003,N_16875);
nand U18593 (N_18593,N_16860,N_16355);
and U18594 (N_18594,N_15283,N_16799);
and U18595 (N_18595,N_17207,N_16804);
or U18596 (N_18596,N_15050,N_15520);
or U18597 (N_18597,N_16684,N_17149);
xor U18598 (N_18598,N_15417,N_15561);
nand U18599 (N_18599,N_15013,N_17019);
nand U18600 (N_18600,N_15829,N_17124);
or U18601 (N_18601,N_15617,N_15052);
nor U18602 (N_18602,N_16529,N_15768);
xor U18603 (N_18603,N_15043,N_15815);
or U18604 (N_18604,N_16603,N_15516);
nand U18605 (N_18605,N_16750,N_16416);
nand U18606 (N_18606,N_15538,N_15912);
and U18607 (N_18607,N_16205,N_16635);
xor U18608 (N_18608,N_16294,N_15503);
and U18609 (N_18609,N_15934,N_17171);
or U18610 (N_18610,N_16686,N_15564);
or U18611 (N_18611,N_16963,N_16056);
and U18612 (N_18612,N_16012,N_15906);
nor U18613 (N_18613,N_17122,N_16978);
and U18614 (N_18614,N_15598,N_16619);
xnor U18615 (N_18615,N_16555,N_16088);
and U18616 (N_18616,N_15527,N_15709);
or U18617 (N_18617,N_15435,N_16792);
and U18618 (N_18618,N_15034,N_16156);
nand U18619 (N_18619,N_15159,N_16029);
and U18620 (N_18620,N_17330,N_15733);
or U18621 (N_18621,N_16094,N_17114);
and U18622 (N_18622,N_15602,N_16315);
nor U18623 (N_18623,N_17221,N_17269);
nor U18624 (N_18624,N_17161,N_17058);
nand U18625 (N_18625,N_17105,N_15143);
nor U18626 (N_18626,N_15805,N_16621);
xor U18627 (N_18627,N_16003,N_15761);
nor U18628 (N_18628,N_16405,N_16831);
nand U18629 (N_18629,N_16570,N_15041);
and U18630 (N_18630,N_17308,N_16311);
and U18631 (N_18631,N_17449,N_15359);
or U18632 (N_18632,N_15323,N_16954);
or U18633 (N_18633,N_16136,N_15952);
nor U18634 (N_18634,N_17057,N_15044);
nand U18635 (N_18635,N_15850,N_16993);
and U18636 (N_18636,N_17440,N_15848);
and U18637 (N_18637,N_15676,N_16847);
nand U18638 (N_18638,N_16244,N_17457);
nor U18639 (N_18639,N_16678,N_17307);
nor U18640 (N_18640,N_16537,N_16301);
nand U18641 (N_18641,N_16335,N_15555);
and U18642 (N_18642,N_15451,N_15808);
and U18643 (N_18643,N_16581,N_15284);
xor U18644 (N_18644,N_16901,N_15717);
nand U18645 (N_18645,N_15917,N_17223);
nand U18646 (N_18646,N_15421,N_16113);
nor U18647 (N_18647,N_15571,N_17380);
and U18648 (N_18648,N_15092,N_15695);
and U18649 (N_18649,N_16128,N_16845);
or U18650 (N_18650,N_15240,N_15017);
xor U18651 (N_18651,N_16928,N_16808);
nor U18652 (N_18652,N_16097,N_16759);
and U18653 (N_18653,N_15370,N_16737);
xor U18654 (N_18654,N_15953,N_17474);
nor U18655 (N_18655,N_16187,N_16293);
nand U18656 (N_18656,N_15728,N_16776);
nor U18657 (N_18657,N_15167,N_17351);
and U18658 (N_18658,N_15530,N_17322);
nor U18659 (N_18659,N_15108,N_15889);
nand U18660 (N_18660,N_16863,N_15639);
or U18661 (N_18661,N_15039,N_15187);
xor U18662 (N_18662,N_16904,N_17079);
and U18663 (N_18663,N_16176,N_16473);
nand U18664 (N_18664,N_16680,N_16712);
nand U18665 (N_18665,N_15383,N_15169);
nand U18666 (N_18666,N_15259,N_15281);
nand U18667 (N_18667,N_15224,N_17334);
nand U18668 (N_18668,N_15441,N_15680);
xnor U18669 (N_18669,N_16280,N_15067);
xor U18670 (N_18670,N_15662,N_15099);
nor U18671 (N_18671,N_15524,N_16199);
xor U18672 (N_18672,N_15577,N_15191);
nor U18673 (N_18673,N_17467,N_15193);
and U18674 (N_18674,N_15542,N_15437);
and U18675 (N_18675,N_15113,N_16994);
xor U18676 (N_18676,N_17011,N_16158);
and U18677 (N_18677,N_16078,N_16009);
nor U18678 (N_18678,N_15731,N_17416);
or U18679 (N_18679,N_17253,N_17397);
nand U18680 (N_18680,N_16231,N_17374);
nor U18681 (N_18681,N_16687,N_15852);
nand U18682 (N_18682,N_17126,N_17000);
nand U18683 (N_18683,N_16490,N_16981);
and U18684 (N_18684,N_16171,N_17318);
nor U18685 (N_18685,N_16502,N_15111);
nand U18686 (N_18686,N_16819,N_16599);
nor U18687 (N_18687,N_15868,N_16588);
and U18688 (N_18688,N_15458,N_17289);
or U18689 (N_18689,N_15650,N_16454);
and U18690 (N_18690,N_15388,N_16440);
xor U18691 (N_18691,N_15832,N_15068);
xor U18692 (N_18692,N_16261,N_16185);
and U18693 (N_18693,N_15438,N_15818);
or U18694 (N_18694,N_15472,N_15381);
nor U18695 (N_18695,N_16045,N_15659);
xor U18696 (N_18696,N_15011,N_15419);
and U18697 (N_18697,N_16878,N_16855);
nand U18698 (N_18698,N_15277,N_16361);
xor U18699 (N_18699,N_17432,N_15216);
and U18700 (N_18700,N_16917,N_16225);
nand U18701 (N_18701,N_16283,N_17102);
nand U18702 (N_18702,N_15777,N_16966);
xor U18703 (N_18703,N_15207,N_17493);
and U18704 (N_18704,N_16566,N_17250);
xor U18705 (N_18705,N_15772,N_16573);
xor U18706 (N_18706,N_15641,N_16696);
nand U18707 (N_18707,N_16967,N_15726);
nand U18708 (N_18708,N_17425,N_15859);
nand U18709 (N_18709,N_17106,N_15605);
or U18710 (N_18710,N_15339,N_16955);
or U18711 (N_18711,N_15401,N_15194);
or U18712 (N_18712,N_16299,N_17180);
or U18713 (N_18713,N_15582,N_15116);
nand U18714 (N_18714,N_15517,N_16970);
nand U18715 (N_18715,N_16150,N_16149);
xnor U18716 (N_18716,N_15618,N_15483);
and U18717 (N_18717,N_15539,N_16707);
nor U18718 (N_18718,N_16013,N_16378);
nand U18719 (N_18719,N_15139,N_16865);
xor U18720 (N_18720,N_16992,N_15319);
xor U18721 (N_18721,N_17055,N_16784);
nor U18722 (N_18722,N_16411,N_15492);
xnor U18723 (N_18723,N_17335,N_16644);
and U18724 (N_18724,N_17081,N_16528);
xnor U18725 (N_18725,N_16508,N_15784);
nand U18726 (N_18726,N_17138,N_16020);
xor U18727 (N_18727,N_16763,N_15335);
and U18728 (N_18728,N_16219,N_16332);
xnor U18729 (N_18729,N_15426,N_15899);
nor U18730 (N_18730,N_17075,N_15468);
and U18731 (N_18731,N_16849,N_16533);
xor U18732 (N_18732,N_15407,N_15698);
xnor U18733 (N_18733,N_15672,N_16880);
nor U18734 (N_18734,N_16210,N_16706);
and U18735 (N_18735,N_17092,N_16400);
nor U18736 (N_18736,N_17040,N_15497);
nor U18737 (N_18737,N_16403,N_15263);
and U18738 (N_18738,N_16998,N_16953);
xor U18739 (N_18739,N_15328,N_16446);
nand U18740 (N_18740,N_15223,N_16942);
nand U18741 (N_18741,N_15643,N_15622);
and U18742 (N_18742,N_16682,N_15687);
and U18743 (N_18743,N_16673,N_15752);
or U18744 (N_18744,N_16087,N_17239);
nor U18745 (N_18745,N_17438,N_17256);
nor U18746 (N_18746,N_17110,N_15624);
xnor U18747 (N_18747,N_17395,N_15964);
xnor U18748 (N_18748,N_15766,N_15480);
and U18749 (N_18749,N_16066,N_15231);
nand U18750 (N_18750,N_16654,N_15072);
or U18751 (N_18751,N_15638,N_16898);
nand U18752 (N_18752,N_15648,N_17012);
nor U18753 (N_18753,N_16813,N_15308);
xor U18754 (N_18754,N_15810,N_16436);
nand U18755 (N_18755,N_16561,N_15063);
nand U18756 (N_18756,N_16733,N_17166);
and U18757 (N_18757,N_15130,N_15982);
and U18758 (N_18758,N_17361,N_15514);
nand U18759 (N_18759,N_16143,N_16742);
and U18760 (N_18760,N_16665,N_16634);
and U18761 (N_18761,N_17412,N_16818);
nor U18762 (N_18762,N_17455,N_15020);
nand U18763 (N_18763,N_16893,N_17185);
or U18764 (N_18764,N_15668,N_17062);
or U18765 (N_18765,N_16922,N_15545);
or U18766 (N_18766,N_16045,N_16718);
nor U18767 (N_18767,N_15756,N_16703);
nor U18768 (N_18768,N_17093,N_15010);
or U18769 (N_18769,N_16204,N_16768);
or U18770 (N_18770,N_15547,N_15181);
nor U18771 (N_18771,N_15069,N_16002);
nor U18772 (N_18772,N_16924,N_15632);
nand U18773 (N_18773,N_16841,N_16237);
and U18774 (N_18774,N_15635,N_15287);
and U18775 (N_18775,N_15651,N_15749);
nor U18776 (N_18776,N_16368,N_17041);
xor U18777 (N_18777,N_17407,N_15587);
nor U18778 (N_18778,N_15569,N_15856);
nand U18779 (N_18779,N_15829,N_15539);
nand U18780 (N_18780,N_16293,N_16541);
nor U18781 (N_18781,N_15302,N_16463);
and U18782 (N_18782,N_15270,N_17085);
xor U18783 (N_18783,N_16265,N_17365);
xnor U18784 (N_18784,N_16827,N_15836);
and U18785 (N_18785,N_15781,N_15701);
nor U18786 (N_18786,N_17037,N_16524);
xnor U18787 (N_18787,N_15641,N_17304);
xor U18788 (N_18788,N_15395,N_15009);
nor U18789 (N_18789,N_16690,N_16138);
or U18790 (N_18790,N_16288,N_15077);
nand U18791 (N_18791,N_15723,N_17174);
nor U18792 (N_18792,N_17066,N_15153);
or U18793 (N_18793,N_16976,N_16691);
and U18794 (N_18794,N_17158,N_15969);
xnor U18795 (N_18795,N_15111,N_17051);
or U18796 (N_18796,N_15590,N_15446);
or U18797 (N_18797,N_17202,N_15034);
xnor U18798 (N_18798,N_17179,N_16193);
nor U18799 (N_18799,N_15342,N_15284);
and U18800 (N_18800,N_17370,N_15853);
or U18801 (N_18801,N_17075,N_16861);
or U18802 (N_18802,N_15649,N_15856);
nand U18803 (N_18803,N_16188,N_16205);
and U18804 (N_18804,N_17053,N_17284);
nand U18805 (N_18805,N_15189,N_16896);
and U18806 (N_18806,N_15044,N_16088);
nor U18807 (N_18807,N_16019,N_15562);
or U18808 (N_18808,N_15863,N_16677);
nor U18809 (N_18809,N_16572,N_15578);
nor U18810 (N_18810,N_17463,N_15976);
or U18811 (N_18811,N_16501,N_15021);
or U18812 (N_18812,N_16887,N_15199);
nor U18813 (N_18813,N_17367,N_16895);
nor U18814 (N_18814,N_16378,N_15004);
nand U18815 (N_18815,N_15386,N_16995);
or U18816 (N_18816,N_16408,N_16221);
xnor U18817 (N_18817,N_15641,N_16521);
nand U18818 (N_18818,N_15325,N_15813);
nor U18819 (N_18819,N_15479,N_16683);
xor U18820 (N_18820,N_16483,N_15584);
nor U18821 (N_18821,N_15600,N_15693);
xnor U18822 (N_18822,N_17383,N_16179);
nand U18823 (N_18823,N_17003,N_15578);
or U18824 (N_18824,N_16026,N_16041);
nor U18825 (N_18825,N_15279,N_16791);
nor U18826 (N_18826,N_16771,N_15785);
nor U18827 (N_18827,N_16821,N_15364);
nand U18828 (N_18828,N_17487,N_17256);
or U18829 (N_18829,N_16689,N_17104);
nor U18830 (N_18830,N_17156,N_17001);
nor U18831 (N_18831,N_15704,N_15922);
nand U18832 (N_18832,N_17176,N_17490);
xnor U18833 (N_18833,N_17267,N_17262);
or U18834 (N_18834,N_17498,N_16938);
nor U18835 (N_18835,N_15469,N_16711);
nor U18836 (N_18836,N_16357,N_15577);
nor U18837 (N_18837,N_15819,N_16727);
xor U18838 (N_18838,N_16646,N_15106);
xor U18839 (N_18839,N_16583,N_16097);
xnor U18840 (N_18840,N_17218,N_17135);
nand U18841 (N_18841,N_16733,N_15728);
nor U18842 (N_18842,N_16202,N_17012);
and U18843 (N_18843,N_15687,N_15058);
and U18844 (N_18844,N_16936,N_15235);
or U18845 (N_18845,N_16557,N_17127);
or U18846 (N_18846,N_16010,N_16819);
nand U18847 (N_18847,N_15086,N_16605);
nand U18848 (N_18848,N_16506,N_15292);
or U18849 (N_18849,N_15674,N_17327);
nor U18850 (N_18850,N_15084,N_16487);
and U18851 (N_18851,N_16733,N_15652);
and U18852 (N_18852,N_16636,N_15655);
or U18853 (N_18853,N_17412,N_16967);
nor U18854 (N_18854,N_15128,N_16105);
nand U18855 (N_18855,N_17484,N_15841);
nand U18856 (N_18856,N_17190,N_17435);
nand U18857 (N_18857,N_17403,N_16518);
nor U18858 (N_18858,N_17208,N_15722);
xnor U18859 (N_18859,N_16041,N_16331);
or U18860 (N_18860,N_15467,N_17480);
nor U18861 (N_18861,N_15793,N_15704);
nor U18862 (N_18862,N_15421,N_15449);
nand U18863 (N_18863,N_17027,N_15589);
nor U18864 (N_18864,N_15324,N_16369);
xor U18865 (N_18865,N_15016,N_17099);
nand U18866 (N_18866,N_17407,N_16392);
and U18867 (N_18867,N_16154,N_15509);
nand U18868 (N_18868,N_17407,N_15838);
nor U18869 (N_18869,N_16523,N_15903);
or U18870 (N_18870,N_15498,N_15426);
and U18871 (N_18871,N_15126,N_15735);
nand U18872 (N_18872,N_15837,N_15718);
nand U18873 (N_18873,N_16336,N_16672);
xor U18874 (N_18874,N_15127,N_15682);
xnor U18875 (N_18875,N_17083,N_16967);
or U18876 (N_18876,N_15099,N_17003);
or U18877 (N_18877,N_15633,N_17369);
nor U18878 (N_18878,N_15210,N_16113);
or U18879 (N_18879,N_17108,N_15443);
or U18880 (N_18880,N_15031,N_17044);
nor U18881 (N_18881,N_15228,N_16159);
nor U18882 (N_18882,N_15090,N_16394);
xor U18883 (N_18883,N_17228,N_16221);
nor U18884 (N_18884,N_15958,N_16048);
and U18885 (N_18885,N_16553,N_15380);
or U18886 (N_18886,N_15424,N_15347);
xnor U18887 (N_18887,N_15805,N_15427);
nor U18888 (N_18888,N_15682,N_15455);
xnor U18889 (N_18889,N_15884,N_16290);
and U18890 (N_18890,N_16730,N_16721);
xor U18891 (N_18891,N_15611,N_15348);
xnor U18892 (N_18892,N_15499,N_16840);
nand U18893 (N_18893,N_16602,N_16141);
nand U18894 (N_18894,N_16337,N_16391);
nor U18895 (N_18895,N_16873,N_17288);
or U18896 (N_18896,N_16386,N_16549);
nor U18897 (N_18897,N_16188,N_16123);
nand U18898 (N_18898,N_16560,N_15860);
xor U18899 (N_18899,N_15896,N_16795);
and U18900 (N_18900,N_15775,N_16648);
nor U18901 (N_18901,N_15803,N_17444);
nor U18902 (N_18902,N_16267,N_15116);
nand U18903 (N_18903,N_16210,N_16187);
and U18904 (N_18904,N_16932,N_15734);
nor U18905 (N_18905,N_15114,N_15018);
nor U18906 (N_18906,N_16978,N_17054);
nor U18907 (N_18907,N_16376,N_16553);
and U18908 (N_18908,N_15227,N_15252);
or U18909 (N_18909,N_17428,N_16055);
xor U18910 (N_18910,N_17402,N_16453);
or U18911 (N_18911,N_15679,N_15819);
or U18912 (N_18912,N_16733,N_15736);
or U18913 (N_18913,N_15059,N_17386);
and U18914 (N_18914,N_16358,N_17234);
nand U18915 (N_18915,N_15816,N_16347);
xor U18916 (N_18916,N_15684,N_16874);
or U18917 (N_18917,N_15565,N_15442);
nor U18918 (N_18918,N_16314,N_16077);
xnor U18919 (N_18919,N_15764,N_16161);
nand U18920 (N_18920,N_15292,N_17311);
nand U18921 (N_18921,N_16155,N_15163);
nor U18922 (N_18922,N_15647,N_16471);
or U18923 (N_18923,N_17282,N_17034);
or U18924 (N_18924,N_15394,N_15541);
xor U18925 (N_18925,N_16754,N_17401);
xor U18926 (N_18926,N_15402,N_16339);
nand U18927 (N_18927,N_15051,N_17288);
nor U18928 (N_18928,N_15225,N_16529);
nand U18929 (N_18929,N_16972,N_16634);
xor U18930 (N_18930,N_17157,N_15057);
and U18931 (N_18931,N_15967,N_15738);
and U18932 (N_18932,N_17498,N_15529);
nand U18933 (N_18933,N_16054,N_15900);
nor U18934 (N_18934,N_15660,N_16414);
and U18935 (N_18935,N_15387,N_17050);
nor U18936 (N_18936,N_17119,N_17177);
and U18937 (N_18937,N_16977,N_16744);
or U18938 (N_18938,N_15893,N_17083);
nand U18939 (N_18939,N_16493,N_16944);
or U18940 (N_18940,N_17227,N_15246);
nor U18941 (N_18941,N_16693,N_15836);
or U18942 (N_18942,N_16639,N_17044);
and U18943 (N_18943,N_15414,N_17486);
and U18944 (N_18944,N_17336,N_16837);
or U18945 (N_18945,N_16139,N_17452);
xor U18946 (N_18946,N_16839,N_16779);
xor U18947 (N_18947,N_15417,N_15859);
and U18948 (N_18948,N_15810,N_17264);
xor U18949 (N_18949,N_15652,N_15071);
and U18950 (N_18950,N_15131,N_15098);
xnor U18951 (N_18951,N_16110,N_17048);
or U18952 (N_18952,N_16282,N_16477);
nand U18953 (N_18953,N_15156,N_16763);
or U18954 (N_18954,N_16213,N_15175);
xnor U18955 (N_18955,N_16294,N_15954);
and U18956 (N_18956,N_16168,N_17202);
xnor U18957 (N_18957,N_15225,N_16434);
xor U18958 (N_18958,N_15904,N_15728);
xnor U18959 (N_18959,N_16561,N_16513);
or U18960 (N_18960,N_15221,N_15896);
and U18961 (N_18961,N_15841,N_16392);
nor U18962 (N_18962,N_17354,N_15734);
nand U18963 (N_18963,N_15184,N_16133);
xnor U18964 (N_18964,N_15954,N_15012);
xnor U18965 (N_18965,N_15964,N_15060);
nand U18966 (N_18966,N_15066,N_15497);
nor U18967 (N_18967,N_16418,N_15985);
xnor U18968 (N_18968,N_15506,N_16033);
xor U18969 (N_18969,N_15186,N_15871);
nor U18970 (N_18970,N_15453,N_15664);
xnor U18971 (N_18971,N_16184,N_16883);
nor U18972 (N_18972,N_15836,N_17275);
nor U18973 (N_18973,N_15245,N_16719);
nor U18974 (N_18974,N_17067,N_15275);
nand U18975 (N_18975,N_17350,N_17376);
and U18976 (N_18976,N_15295,N_15624);
and U18977 (N_18977,N_15709,N_16753);
nand U18978 (N_18978,N_15318,N_15837);
nand U18979 (N_18979,N_17245,N_16238);
nand U18980 (N_18980,N_16806,N_15222);
or U18981 (N_18981,N_16365,N_16132);
and U18982 (N_18982,N_15515,N_17314);
or U18983 (N_18983,N_15940,N_16219);
and U18984 (N_18984,N_17064,N_16037);
and U18985 (N_18985,N_17467,N_15629);
or U18986 (N_18986,N_15823,N_15063);
and U18987 (N_18987,N_15015,N_16989);
nor U18988 (N_18988,N_16083,N_16204);
or U18989 (N_18989,N_15782,N_16399);
and U18990 (N_18990,N_17467,N_17072);
xnor U18991 (N_18991,N_17166,N_15250);
nor U18992 (N_18992,N_17069,N_16864);
and U18993 (N_18993,N_17216,N_17184);
or U18994 (N_18994,N_15566,N_15016);
and U18995 (N_18995,N_15305,N_16000);
xor U18996 (N_18996,N_15193,N_15814);
nor U18997 (N_18997,N_17055,N_15981);
nor U18998 (N_18998,N_15312,N_17250);
or U18999 (N_18999,N_16409,N_16718);
and U19000 (N_19000,N_16749,N_17236);
nor U19001 (N_19001,N_15041,N_16368);
and U19002 (N_19002,N_16317,N_15741);
or U19003 (N_19003,N_16196,N_17326);
and U19004 (N_19004,N_15875,N_15940);
nor U19005 (N_19005,N_15100,N_15415);
nor U19006 (N_19006,N_15586,N_17155);
and U19007 (N_19007,N_16220,N_17075);
nor U19008 (N_19008,N_16365,N_15289);
and U19009 (N_19009,N_17276,N_16391);
nand U19010 (N_19010,N_15555,N_16940);
and U19011 (N_19011,N_15340,N_17064);
nor U19012 (N_19012,N_15489,N_17067);
nand U19013 (N_19013,N_16604,N_17490);
and U19014 (N_19014,N_17377,N_15302);
xor U19015 (N_19015,N_16640,N_16711);
nand U19016 (N_19016,N_16460,N_17438);
nor U19017 (N_19017,N_15506,N_17004);
nand U19018 (N_19018,N_16636,N_15497);
and U19019 (N_19019,N_16061,N_17139);
xor U19020 (N_19020,N_17234,N_17371);
nand U19021 (N_19021,N_17398,N_17000);
nor U19022 (N_19022,N_16451,N_15547);
nand U19023 (N_19023,N_17160,N_17192);
or U19024 (N_19024,N_16271,N_15873);
nor U19025 (N_19025,N_15673,N_16604);
and U19026 (N_19026,N_16825,N_16217);
and U19027 (N_19027,N_16102,N_17148);
nand U19028 (N_19028,N_15330,N_16298);
xnor U19029 (N_19029,N_15117,N_17054);
nand U19030 (N_19030,N_16919,N_17078);
xnor U19031 (N_19031,N_15354,N_16102);
and U19032 (N_19032,N_16740,N_16423);
xor U19033 (N_19033,N_15892,N_16567);
nor U19034 (N_19034,N_15316,N_15160);
nor U19035 (N_19035,N_16840,N_16126);
nor U19036 (N_19036,N_15654,N_17382);
nor U19037 (N_19037,N_15479,N_15935);
nand U19038 (N_19038,N_16756,N_15344);
xor U19039 (N_19039,N_15380,N_15813);
and U19040 (N_19040,N_16408,N_15114);
nor U19041 (N_19041,N_15950,N_16911);
and U19042 (N_19042,N_16715,N_15874);
xnor U19043 (N_19043,N_16337,N_15400);
xor U19044 (N_19044,N_17016,N_15901);
xor U19045 (N_19045,N_16197,N_17238);
nor U19046 (N_19046,N_15003,N_15401);
nor U19047 (N_19047,N_17000,N_15912);
nor U19048 (N_19048,N_17350,N_15542);
and U19049 (N_19049,N_16128,N_15370);
nand U19050 (N_19050,N_17217,N_17188);
and U19051 (N_19051,N_16681,N_15434);
xnor U19052 (N_19052,N_15461,N_16816);
nor U19053 (N_19053,N_15996,N_15953);
or U19054 (N_19054,N_15417,N_16702);
and U19055 (N_19055,N_17039,N_15717);
and U19056 (N_19056,N_16559,N_15508);
nand U19057 (N_19057,N_15098,N_17363);
and U19058 (N_19058,N_17377,N_16758);
or U19059 (N_19059,N_15338,N_16013);
and U19060 (N_19060,N_17498,N_15116);
or U19061 (N_19061,N_16098,N_15427);
nand U19062 (N_19062,N_15907,N_16214);
nand U19063 (N_19063,N_15256,N_16037);
and U19064 (N_19064,N_15008,N_17307);
and U19065 (N_19065,N_15202,N_16344);
and U19066 (N_19066,N_15623,N_17204);
and U19067 (N_19067,N_17415,N_16919);
nor U19068 (N_19068,N_15996,N_15789);
or U19069 (N_19069,N_15734,N_16376);
nand U19070 (N_19070,N_17098,N_15028);
nor U19071 (N_19071,N_16419,N_16571);
xnor U19072 (N_19072,N_15649,N_15744);
or U19073 (N_19073,N_16118,N_16950);
and U19074 (N_19074,N_15708,N_16168);
and U19075 (N_19075,N_15131,N_16526);
xnor U19076 (N_19076,N_15307,N_15554);
nand U19077 (N_19077,N_17252,N_17260);
nor U19078 (N_19078,N_15483,N_15935);
or U19079 (N_19079,N_16066,N_15531);
nand U19080 (N_19080,N_16850,N_17479);
nand U19081 (N_19081,N_17424,N_17173);
nor U19082 (N_19082,N_16219,N_17221);
nor U19083 (N_19083,N_16628,N_16999);
nand U19084 (N_19084,N_17227,N_16185);
xor U19085 (N_19085,N_15973,N_15735);
xor U19086 (N_19086,N_15227,N_15234);
nor U19087 (N_19087,N_16611,N_15911);
and U19088 (N_19088,N_15512,N_16173);
nand U19089 (N_19089,N_15494,N_17486);
nand U19090 (N_19090,N_15452,N_15930);
xnor U19091 (N_19091,N_16094,N_17298);
or U19092 (N_19092,N_15797,N_16321);
or U19093 (N_19093,N_15730,N_16376);
nor U19094 (N_19094,N_17416,N_17343);
nand U19095 (N_19095,N_16756,N_15991);
or U19096 (N_19096,N_15041,N_15655);
nor U19097 (N_19097,N_15445,N_17405);
and U19098 (N_19098,N_15783,N_16800);
or U19099 (N_19099,N_15911,N_17432);
and U19100 (N_19100,N_15666,N_17206);
nand U19101 (N_19101,N_16194,N_15680);
or U19102 (N_19102,N_15429,N_16141);
nor U19103 (N_19103,N_15868,N_16517);
nor U19104 (N_19104,N_16966,N_16265);
xnor U19105 (N_19105,N_16376,N_16182);
nor U19106 (N_19106,N_15903,N_15258);
and U19107 (N_19107,N_16761,N_16759);
nor U19108 (N_19108,N_16140,N_17122);
nor U19109 (N_19109,N_15238,N_15661);
nand U19110 (N_19110,N_15744,N_16110);
nand U19111 (N_19111,N_15164,N_16613);
and U19112 (N_19112,N_15867,N_16168);
and U19113 (N_19113,N_15754,N_17214);
nor U19114 (N_19114,N_15458,N_16577);
nand U19115 (N_19115,N_15796,N_17043);
xor U19116 (N_19116,N_17152,N_15097);
nor U19117 (N_19117,N_16887,N_15967);
and U19118 (N_19118,N_17188,N_16344);
nor U19119 (N_19119,N_15439,N_17100);
xor U19120 (N_19120,N_15058,N_16074);
or U19121 (N_19121,N_16713,N_16003);
or U19122 (N_19122,N_16299,N_16376);
nor U19123 (N_19123,N_16286,N_15006);
xnor U19124 (N_19124,N_16231,N_17425);
nand U19125 (N_19125,N_17320,N_16261);
and U19126 (N_19126,N_17149,N_15253);
nand U19127 (N_19127,N_15668,N_15640);
xnor U19128 (N_19128,N_15040,N_15728);
and U19129 (N_19129,N_17262,N_16821);
nor U19130 (N_19130,N_16917,N_15528);
nand U19131 (N_19131,N_16111,N_17325);
xor U19132 (N_19132,N_16975,N_16903);
and U19133 (N_19133,N_16553,N_15991);
or U19134 (N_19134,N_16604,N_16349);
and U19135 (N_19135,N_17120,N_15019);
and U19136 (N_19136,N_17167,N_17370);
nand U19137 (N_19137,N_15105,N_16259);
xnor U19138 (N_19138,N_16487,N_15934);
and U19139 (N_19139,N_16622,N_16634);
nand U19140 (N_19140,N_17398,N_16054);
nand U19141 (N_19141,N_15406,N_17084);
xnor U19142 (N_19142,N_15207,N_16393);
or U19143 (N_19143,N_16639,N_16448);
nand U19144 (N_19144,N_16956,N_16526);
or U19145 (N_19145,N_17357,N_17213);
nor U19146 (N_19146,N_16590,N_16827);
xor U19147 (N_19147,N_16195,N_15162);
or U19148 (N_19148,N_17291,N_16358);
xor U19149 (N_19149,N_16784,N_15308);
xor U19150 (N_19150,N_17388,N_17415);
and U19151 (N_19151,N_16518,N_15450);
or U19152 (N_19152,N_17232,N_15521);
or U19153 (N_19153,N_16005,N_16328);
nand U19154 (N_19154,N_17391,N_17114);
xor U19155 (N_19155,N_17260,N_16941);
xnor U19156 (N_19156,N_16607,N_16769);
or U19157 (N_19157,N_17279,N_15211);
nor U19158 (N_19158,N_16944,N_17295);
nand U19159 (N_19159,N_15867,N_16139);
or U19160 (N_19160,N_15183,N_17214);
nand U19161 (N_19161,N_15606,N_15813);
xor U19162 (N_19162,N_16193,N_15665);
and U19163 (N_19163,N_16446,N_16152);
xnor U19164 (N_19164,N_17356,N_15964);
xor U19165 (N_19165,N_15239,N_16921);
or U19166 (N_19166,N_15179,N_17395);
nor U19167 (N_19167,N_16217,N_15022);
nand U19168 (N_19168,N_16481,N_16886);
nor U19169 (N_19169,N_16356,N_15194);
xnor U19170 (N_19170,N_17199,N_17191);
xnor U19171 (N_19171,N_16267,N_16905);
or U19172 (N_19172,N_16281,N_16171);
and U19173 (N_19173,N_16705,N_15179);
or U19174 (N_19174,N_15673,N_17255);
nor U19175 (N_19175,N_15247,N_15380);
and U19176 (N_19176,N_15303,N_16169);
xor U19177 (N_19177,N_17211,N_15993);
nand U19178 (N_19178,N_16351,N_16305);
and U19179 (N_19179,N_15112,N_17478);
nor U19180 (N_19180,N_16684,N_15394);
xnor U19181 (N_19181,N_15330,N_15792);
nor U19182 (N_19182,N_15971,N_15202);
and U19183 (N_19183,N_15389,N_15837);
xor U19184 (N_19184,N_17394,N_15268);
and U19185 (N_19185,N_15442,N_15938);
nand U19186 (N_19186,N_16898,N_15261);
or U19187 (N_19187,N_17435,N_15118);
and U19188 (N_19188,N_15486,N_16870);
and U19189 (N_19189,N_16129,N_15453);
and U19190 (N_19190,N_17260,N_17313);
nand U19191 (N_19191,N_17287,N_16425);
nor U19192 (N_19192,N_16036,N_16346);
xnor U19193 (N_19193,N_16581,N_15520);
nor U19194 (N_19194,N_16133,N_16359);
or U19195 (N_19195,N_17227,N_15170);
nand U19196 (N_19196,N_17187,N_17370);
and U19197 (N_19197,N_17125,N_16657);
xor U19198 (N_19198,N_15907,N_17406);
xor U19199 (N_19199,N_16239,N_16766);
and U19200 (N_19200,N_15851,N_17122);
xor U19201 (N_19201,N_16024,N_15854);
or U19202 (N_19202,N_15017,N_17354);
xnor U19203 (N_19203,N_15610,N_17319);
xnor U19204 (N_19204,N_15122,N_17086);
nor U19205 (N_19205,N_16123,N_17046);
nand U19206 (N_19206,N_17393,N_15265);
and U19207 (N_19207,N_15682,N_15608);
nor U19208 (N_19208,N_15318,N_16363);
and U19209 (N_19209,N_16630,N_17124);
nor U19210 (N_19210,N_15064,N_15014);
xor U19211 (N_19211,N_15908,N_15315);
nand U19212 (N_19212,N_16665,N_16935);
or U19213 (N_19213,N_15906,N_16275);
nand U19214 (N_19214,N_16340,N_15905);
nand U19215 (N_19215,N_15637,N_16381);
xnor U19216 (N_19216,N_17282,N_16067);
and U19217 (N_19217,N_17368,N_16207);
or U19218 (N_19218,N_16403,N_15912);
or U19219 (N_19219,N_17277,N_16783);
nand U19220 (N_19220,N_16345,N_15969);
nor U19221 (N_19221,N_15894,N_15437);
xor U19222 (N_19222,N_15148,N_16728);
nand U19223 (N_19223,N_16477,N_17201);
and U19224 (N_19224,N_15981,N_15176);
or U19225 (N_19225,N_17132,N_16803);
and U19226 (N_19226,N_17479,N_17179);
nand U19227 (N_19227,N_17384,N_16374);
xnor U19228 (N_19228,N_17329,N_16038);
xor U19229 (N_19229,N_16500,N_16759);
xnor U19230 (N_19230,N_15011,N_15483);
or U19231 (N_19231,N_17261,N_16396);
xnor U19232 (N_19232,N_17073,N_16559);
nor U19233 (N_19233,N_15370,N_15495);
xor U19234 (N_19234,N_16359,N_15298);
or U19235 (N_19235,N_16484,N_15228);
xnor U19236 (N_19236,N_16070,N_16206);
xnor U19237 (N_19237,N_16815,N_16971);
xnor U19238 (N_19238,N_17102,N_15650);
and U19239 (N_19239,N_16804,N_16904);
or U19240 (N_19240,N_16820,N_15433);
nor U19241 (N_19241,N_16262,N_15771);
nor U19242 (N_19242,N_15722,N_15964);
and U19243 (N_19243,N_17000,N_15973);
or U19244 (N_19244,N_16720,N_15810);
and U19245 (N_19245,N_16859,N_15803);
nor U19246 (N_19246,N_15904,N_16603);
and U19247 (N_19247,N_15796,N_15414);
nand U19248 (N_19248,N_16195,N_15241);
nand U19249 (N_19249,N_16969,N_16629);
nand U19250 (N_19250,N_17119,N_16452);
xor U19251 (N_19251,N_15778,N_15038);
nor U19252 (N_19252,N_15409,N_15563);
xnor U19253 (N_19253,N_17144,N_15827);
or U19254 (N_19254,N_16031,N_17280);
and U19255 (N_19255,N_16518,N_16973);
nor U19256 (N_19256,N_16737,N_15431);
xor U19257 (N_19257,N_15630,N_15281);
nor U19258 (N_19258,N_16323,N_16111);
or U19259 (N_19259,N_16343,N_16319);
or U19260 (N_19260,N_15579,N_16090);
nor U19261 (N_19261,N_16817,N_15837);
or U19262 (N_19262,N_15120,N_16839);
or U19263 (N_19263,N_16790,N_16839);
nand U19264 (N_19264,N_15424,N_16005);
xor U19265 (N_19265,N_16292,N_17083);
nor U19266 (N_19266,N_15068,N_16763);
nand U19267 (N_19267,N_15974,N_16259);
nand U19268 (N_19268,N_16875,N_16840);
nor U19269 (N_19269,N_15991,N_16293);
or U19270 (N_19270,N_15033,N_16118);
or U19271 (N_19271,N_16054,N_17014);
and U19272 (N_19272,N_15636,N_15386);
xnor U19273 (N_19273,N_15357,N_15165);
nor U19274 (N_19274,N_16012,N_15581);
xnor U19275 (N_19275,N_16818,N_17133);
xnor U19276 (N_19276,N_16103,N_17076);
nor U19277 (N_19277,N_16918,N_16919);
xnor U19278 (N_19278,N_15557,N_16037);
nand U19279 (N_19279,N_15965,N_15629);
xor U19280 (N_19280,N_17152,N_17026);
xnor U19281 (N_19281,N_15164,N_16308);
nand U19282 (N_19282,N_16780,N_15946);
and U19283 (N_19283,N_15668,N_16225);
nor U19284 (N_19284,N_17491,N_15339);
and U19285 (N_19285,N_15939,N_16164);
nand U19286 (N_19286,N_15911,N_15359);
and U19287 (N_19287,N_15349,N_15710);
nor U19288 (N_19288,N_16333,N_15607);
and U19289 (N_19289,N_17459,N_16629);
xnor U19290 (N_19290,N_16131,N_17351);
xor U19291 (N_19291,N_17248,N_16648);
xnor U19292 (N_19292,N_16225,N_16045);
and U19293 (N_19293,N_16197,N_17265);
nor U19294 (N_19294,N_15207,N_17061);
and U19295 (N_19295,N_16594,N_15543);
xnor U19296 (N_19296,N_15387,N_15980);
or U19297 (N_19297,N_15256,N_15575);
or U19298 (N_19298,N_16466,N_15242);
xor U19299 (N_19299,N_16501,N_16184);
nor U19300 (N_19300,N_15870,N_16654);
or U19301 (N_19301,N_15914,N_15770);
xor U19302 (N_19302,N_15482,N_15521);
or U19303 (N_19303,N_15142,N_16757);
nand U19304 (N_19304,N_16590,N_16299);
nand U19305 (N_19305,N_17010,N_15954);
and U19306 (N_19306,N_15923,N_16503);
nor U19307 (N_19307,N_16060,N_16307);
xnor U19308 (N_19308,N_16555,N_16898);
xnor U19309 (N_19309,N_16587,N_17486);
nand U19310 (N_19310,N_16524,N_17376);
and U19311 (N_19311,N_17119,N_15423);
and U19312 (N_19312,N_15710,N_15261);
or U19313 (N_19313,N_16237,N_16353);
or U19314 (N_19314,N_17311,N_17145);
nand U19315 (N_19315,N_16370,N_16420);
xor U19316 (N_19316,N_16374,N_15218);
xnor U19317 (N_19317,N_15147,N_16082);
nor U19318 (N_19318,N_15699,N_15570);
or U19319 (N_19319,N_17313,N_15498);
nor U19320 (N_19320,N_15193,N_17179);
nand U19321 (N_19321,N_16400,N_17008);
nand U19322 (N_19322,N_15131,N_15474);
nand U19323 (N_19323,N_16992,N_15625);
nand U19324 (N_19324,N_16902,N_15772);
xor U19325 (N_19325,N_16165,N_17272);
xnor U19326 (N_19326,N_16044,N_15533);
nor U19327 (N_19327,N_16105,N_15020);
nand U19328 (N_19328,N_15595,N_15931);
nor U19329 (N_19329,N_15490,N_15838);
or U19330 (N_19330,N_15234,N_15034);
nand U19331 (N_19331,N_16936,N_15180);
and U19332 (N_19332,N_15276,N_16871);
nor U19333 (N_19333,N_15411,N_16555);
nor U19334 (N_19334,N_15228,N_16059);
and U19335 (N_19335,N_15746,N_15848);
xor U19336 (N_19336,N_15931,N_15559);
and U19337 (N_19337,N_16228,N_15475);
nor U19338 (N_19338,N_17487,N_16962);
nor U19339 (N_19339,N_16778,N_17408);
and U19340 (N_19340,N_16910,N_15941);
and U19341 (N_19341,N_17417,N_15258);
nand U19342 (N_19342,N_16378,N_15151);
and U19343 (N_19343,N_17171,N_15011);
and U19344 (N_19344,N_17425,N_16884);
or U19345 (N_19345,N_16573,N_16464);
nor U19346 (N_19346,N_16209,N_16024);
nand U19347 (N_19347,N_16828,N_16429);
and U19348 (N_19348,N_15886,N_15204);
nor U19349 (N_19349,N_17113,N_16463);
nand U19350 (N_19350,N_15555,N_15429);
and U19351 (N_19351,N_17470,N_15220);
nor U19352 (N_19352,N_15292,N_17410);
xor U19353 (N_19353,N_16816,N_15923);
nor U19354 (N_19354,N_16947,N_15646);
or U19355 (N_19355,N_16049,N_16769);
nand U19356 (N_19356,N_17047,N_15041);
and U19357 (N_19357,N_17185,N_15857);
and U19358 (N_19358,N_16292,N_16223);
and U19359 (N_19359,N_15335,N_16589);
or U19360 (N_19360,N_17314,N_17412);
xor U19361 (N_19361,N_16317,N_17295);
and U19362 (N_19362,N_16626,N_15898);
xnor U19363 (N_19363,N_15409,N_16418);
and U19364 (N_19364,N_15739,N_17278);
xnor U19365 (N_19365,N_15429,N_15154);
nor U19366 (N_19366,N_15046,N_15888);
xnor U19367 (N_19367,N_15050,N_15698);
xor U19368 (N_19368,N_15824,N_15079);
or U19369 (N_19369,N_16690,N_15432);
or U19370 (N_19370,N_15056,N_15908);
and U19371 (N_19371,N_16367,N_17377);
xnor U19372 (N_19372,N_16187,N_17480);
nand U19373 (N_19373,N_15540,N_16207);
and U19374 (N_19374,N_16013,N_16889);
and U19375 (N_19375,N_16628,N_16814);
xnor U19376 (N_19376,N_17175,N_15154);
xnor U19377 (N_19377,N_15216,N_15903);
nor U19378 (N_19378,N_16900,N_17436);
and U19379 (N_19379,N_16390,N_15079);
or U19380 (N_19380,N_17396,N_15015);
and U19381 (N_19381,N_16765,N_16140);
nand U19382 (N_19382,N_16718,N_15323);
xnor U19383 (N_19383,N_16920,N_17295);
and U19384 (N_19384,N_15216,N_15804);
and U19385 (N_19385,N_17331,N_16812);
nor U19386 (N_19386,N_16661,N_15839);
or U19387 (N_19387,N_16499,N_16808);
xnor U19388 (N_19388,N_15893,N_16258);
nor U19389 (N_19389,N_15762,N_15318);
nor U19390 (N_19390,N_17477,N_16016);
nor U19391 (N_19391,N_15319,N_16024);
nand U19392 (N_19392,N_15298,N_15637);
nand U19393 (N_19393,N_17457,N_15445);
and U19394 (N_19394,N_15036,N_17121);
nand U19395 (N_19395,N_17137,N_16457);
xor U19396 (N_19396,N_16821,N_16702);
nor U19397 (N_19397,N_17118,N_15516);
nor U19398 (N_19398,N_17237,N_16687);
nand U19399 (N_19399,N_16270,N_15188);
nand U19400 (N_19400,N_17060,N_16461);
or U19401 (N_19401,N_16121,N_15774);
or U19402 (N_19402,N_16772,N_16069);
xnor U19403 (N_19403,N_15168,N_16888);
xnor U19404 (N_19404,N_17279,N_15207);
and U19405 (N_19405,N_15902,N_15158);
nand U19406 (N_19406,N_17492,N_17224);
or U19407 (N_19407,N_15570,N_16979);
and U19408 (N_19408,N_15599,N_17164);
nand U19409 (N_19409,N_15070,N_16415);
nor U19410 (N_19410,N_15369,N_15450);
nor U19411 (N_19411,N_15392,N_15290);
nand U19412 (N_19412,N_16533,N_15706);
and U19413 (N_19413,N_17408,N_16300);
and U19414 (N_19414,N_16405,N_17203);
nand U19415 (N_19415,N_16707,N_17304);
and U19416 (N_19416,N_16170,N_16814);
and U19417 (N_19417,N_15194,N_16127);
nor U19418 (N_19418,N_17370,N_17016);
and U19419 (N_19419,N_16681,N_16832);
or U19420 (N_19420,N_16289,N_15902);
xnor U19421 (N_19421,N_15601,N_16755);
nand U19422 (N_19422,N_17097,N_15382);
nor U19423 (N_19423,N_17313,N_17189);
xnor U19424 (N_19424,N_17401,N_16296);
or U19425 (N_19425,N_15855,N_15976);
xor U19426 (N_19426,N_15888,N_15042);
xor U19427 (N_19427,N_15180,N_15003);
nand U19428 (N_19428,N_17118,N_17391);
nor U19429 (N_19429,N_15667,N_15039);
xor U19430 (N_19430,N_17140,N_16699);
nor U19431 (N_19431,N_17414,N_15368);
nor U19432 (N_19432,N_16682,N_15081);
nand U19433 (N_19433,N_16032,N_15240);
nand U19434 (N_19434,N_16185,N_15410);
nor U19435 (N_19435,N_15180,N_16584);
nor U19436 (N_19436,N_15655,N_16678);
nand U19437 (N_19437,N_15648,N_16404);
nand U19438 (N_19438,N_16854,N_16212);
nor U19439 (N_19439,N_17082,N_16626);
nand U19440 (N_19440,N_17017,N_15069);
xnor U19441 (N_19441,N_15531,N_15970);
nor U19442 (N_19442,N_17069,N_16170);
nand U19443 (N_19443,N_15097,N_16743);
xnor U19444 (N_19444,N_17327,N_15824);
nand U19445 (N_19445,N_15807,N_16852);
or U19446 (N_19446,N_15712,N_16684);
or U19447 (N_19447,N_15917,N_15101);
and U19448 (N_19448,N_15263,N_16114);
nor U19449 (N_19449,N_15398,N_16411);
nand U19450 (N_19450,N_15353,N_16150);
and U19451 (N_19451,N_16800,N_16793);
or U19452 (N_19452,N_16735,N_15976);
nor U19453 (N_19453,N_16220,N_15658);
and U19454 (N_19454,N_15271,N_17040);
nand U19455 (N_19455,N_17152,N_16146);
xnor U19456 (N_19456,N_16940,N_15804);
xnor U19457 (N_19457,N_15325,N_15625);
and U19458 (N_19458,N_17440,N_16864);
nand U19459 (N_19459,N_17157,N_15911);
or U19460 (N_19460,N_16696,N_16168);
nand U19461 (N_19461,N_16638,N_16972);
or U19462 (N_19462,N_16969,N_16207);
nor U19463 (N_19463,N_15482,N_16878);
nor U19464 (N_19464,N_16151,N_16364);
and U19465 (N_19465,N_15959,N_17178);
nor U19466 (N_19466,N_17101,N_15845);
and U19467 (N_19467,N_15048,N_16232);
nand U19468 (N_19468,N_15708,N_16635);
nor U19469 (N_19469,N_15104,N_15192);
nor U19470 (N_19470,N_15716,N_16718);
or U19471 (N_19471,N_17198,N_16977);
nand U19472 (N_19472,N_16466,N_16486);
xor U19473 (N_19473,N_16831,N_17244);
xnor U19474 (N_19474,N_16450,N_16251);
xor U19475 (N_19475,N_15401,N_16635);
xor U19476 (N_19476,N_15780,N_15160);
nand U19477 (N_19477,N_15037,N_17112);
or U19478 (N_19478,N_15868,N_16702);
xor U19479 (N_19479,N_16913,N_15388);
nand U19480 (N_19480,N_15103,N_15131);
nand U19481 (N_19481,N_16750,N_16852);
nand U19482 (N_19482,N_16411,N_16706);
and U19483 (N_19483,N_15456,N_16550);
or U19484 (N_19484,N_16192,N_15513);
and U19485 (N_19485,N_15226,N_16565);
nor U19486 (N_19486,N_16032,N_15777);
or U19487 (N_19487,N_16464,N_17153);
or U19488 (N_19488,N_17438,N_15545);
or U19489 (N_19489,N_15514,N_15023);
nand U19490 (N_19490,N_15670,N_15875);
xor U19491 (N_19491,N_15053,N_16657);
or U19492 (N_19492,N_17007,N_15361);
xor U19493 (N_19493,N_16672,N_15410);
nand U19494 (N_19494,N_17020,N_15104);
nor U19495 (N_19495,N_16400,N_17170);
xor U19496 (N_19496,N_15119,N_17173);
or U19497 (N_19497,N_15650,N_15293);
nand U19498 (N_19498,N_15694,N_16232);
nand U19499 (N_19499,N_16938,N_15174);
nand U19500 (N_19500,N_16673,N_15246);
or U19501 (N_19501,N_16608,N_16577);
nor U19502 (N_19502,N_15700,N_17246);
xnor U19503 (N_19503,N_15018,N_16542);
or U19504 (N_19504,N_16981,N_17238);
and U19505 (N_19505,N_17300,N_15014);
nor U19506 (N_19506,N_16173,N_17267);
xor U19507 (N_19507,N_16661,N_16748);
or U19508 (N_19508,N_15835,N_17479);
nor U19509 (N_19509,N_16714,N_17033);
xnor U19510 (N_19510,N_16613,N_15044);
or U19511 (N_19511,N_16614,N_15417);
nor U19512 (N_19512,N_16278,N_15194);
nor U19513 (N_19513,N_16168,N_15195);
xnor U19514 (N_19514,N_15931,N_16986);
or U19515 (N_19515,N_15891,N_16063);
nor U19516 (N_19516,N_16156,N_15823);
or U19517 (N_19517,N_15061,N_15696);
xnor U19518 (N_19518,N_15205,N_16249);
nor U19519 (N_19519,N_16038,N_16968);
nand U19520 (N_19520,N_15183,N_16424);
or U19521 (N_19521,N_15386,N_17049);
and U19522 (N_19522,N_15945,N_15038);
nand U19523 (N_19523,N_15287,N_15311);
nand U19524 (N_19524,N_16949,N_15577);
nand U19525 (N_19525,N_15068,N_17214);
nor U19526 (N_19526,N_16708,N_15738);
xor U19527 (N_19527,N_16154,N_16770);
nor U19528 (N_19528,N_16622,N_16313);
nor U19529 (N_19529,N_16194,N_16168);
nand U19530 (N_19530,N_16151,N_16171);
and U19531 (N_19531,N_17235,N_15306);
and U19532 (N_19532,N_15361,N_16343);
or U19533 (N_19533,N_16906,N_16163);
or U19534 (N_19534,N_17263,N_16679);
nor U19535 (N_19535,N_17389,N_16746);
nand U19536 (N_19536,N_17374,N_16859);
nor U19537 (N_19537,N_17141,N_16390);
nand U19538 (N_19538,N_17328,N_15766);
nor U19539 (N_19539,N_16794,N_16174);
and U19540 (N_19540,N_16854,N_15384);
xor U19541 (N_19541,N_15726,N_15984);
and U19542 (N_19542,N_17148,N_15108);
or U19543 (N_19543,N_16079,N_15829);
or U19544 (N_19544,N_16483,N_15470);
nor U19545 (N_19545,N_15593,N_15535);
xor U19546 (N_19546,N_16975,N_15600);
or U19547 (N_19547,N_17386,N_15030);
and U19548 (N_19548,N_15484,N_17331);
nand U19549 (N_19549,N_15013,N_15514);
nor U19550 (N_19550,N_16083,N_17446);
nand U19551 (N_19551,N_15381,N_15665);
nor U19552 (N_19552,N_17082,N_16379);
and U19553 (N_19553,N_15517,N_16308);
nand U19554 (N_19554,N_17401,N_16199);
and U19555 (N_19555,N_15112,N_16226);
and U19556 (N_19556,N_15432,N_16554);
and U19557 (N_19557,N_15592,N_15473);
or U19558 (N_19558,N_17066,N_17390);
xor U19559 (N_19559,N_16090,N_16187);
nand U19560 (N_19560,N_16005,N_15812);
nor U19561 (N_19561,N_16646,N_15314);
nor U19562 (N_19562,N_15318,N_15693);
nor U19563 (N_19563,N_16382,N_16690);
and U19564 (N_19564,N_16899,N_16614);
xor U19565 (N_19565,N_15134,N_17407);
and U19566 (N_19566,N_15442,N_17271);
nand U19567 (N_19567,N_15519,N_15328);
nand U19568 (N_19568,N_16659,N_16827);
or U19569 (N_19569,N_15370,N_16488);
and U19570 (N_19570,N_17123,N_15365);
and U19571 (N_19571,N_17424,N_16574);
nand U19572 (N_19572,N_17074,N_16330);
nor U19573 (N_19573,N_15522,N_15118);
nand U19574 (N_19574,N_16195,N_15490);
and U19575 (N_19575,N_15239,N_16056);
nor U19576 (N_19576,N_17246,N_16703);
xnor U19577 (N_19577,N_15737,N_15741);
nand U19578 (N_19578,N_15492,N_16751);
nand U19579 (N_19579,N_15538,N_16701);
xnor U19580 (N_19580,N_16201,N_15575);
nand U19581 (N_19581,N_17055,N_17389);
or U19582 (N_19582,N_16548,N_15434);
nor U19583 (N_19583,N_15396,N_17336);
nor U19584 (N_19584,N_15898,N_16753);
and U19585 (N_19585,N_15375,N_15532);
xor U19586 (N_19586,N_16434,N_15139);
and U19587 (N_19587,N_17121,N_15993);
nand U19588 (N_19588,N_16216,N_17319);
and U19589 (N_19589,N_15208,N_15696);
xnor U19590 (N_19590,N_16824,N_17397);
or U19591 (N_19591,N_15728,N_16978);
nor U19592 (N_19592,N_17287,N_15711);
xor U19593 (N_19593,N_16993,N_15659);
or U19594 (N_19594,N_17320,N_17333);
nor U19595 (N_19595,N_16393,N_15102);
xnor U19596 (N_19596,N_15758,N_16004);
nor U19597 (N_19597,N_15329,N_15275);
xnor U19598 (N_19598,N_15059,N_16126);
and U19599 (N_19599,N_15298,N_16464);
or U19600 (N_19600,N_15411,N_16593);
xor U19601 (N_19601,N_16494,N_15457);
nor U19602 (N_19602,N_16572,N_15501);
xor U19603 (N_19603,N_17144,N_16461);
nand U19604 (N_19604,N_15535,N_15862);
nand U19605 (N_19605,N_16641,N_16372);
nand U19606 (N_19606,N_15630,N_16283);
xor U19607 (N_19607,N_17032,N_17036);
nand U19608 (N_19608,N_15892,N_16836);
and U19609 (N_19609,N_16813,N_16285);
xnor U19610 (N_19610,N_16051,N_15535);
or U19611 (N_19611,N_17311,N_16351);
or U19612 (N_19612,N_16832,N_16416);
nor U19613 (N_19613,N_15655,N_16446);
and U19614 (N_19614,N_15824,N_15669);
xor U19615 (N_19615,N_15690,N_17072);
or U19616 (N_19616,N_17081,N_17125);
and U19617 (N_19617,N_15157,N_17212);
or U19618 (N_19618,N_15310,N_17030);
nand U19619 (N_19619,N_15291,N_15990);
nor U19620 (N_19620,N_17011,N_17031);
xor U19621 (N_19621,N_16915,N_16466);
nor U19622 (N_19622,N_16543,N_15824);
nor U19623 (N_19623,N_15060,N_15421);
or U19624 (N_19624,N_16821,N_15475);
or U19625 (N_19625,N_17040,N_15835);
nor U19626 (N_19626,N_15750,N_17127);
xnor U19627 (N_19627,N_15364,N_16093);
xnor U19628 (N_19628,N_16195,N_15165);
or U19629 (N_19629,N_15104,N_16306);
and U19630 (N_19630,N_16626,N_16973);
nand U19631 (N_19631,N_16187,N_15387);
and U19632 (N_19632,N_15626,N_15441);
nor U19633 (N_19633,N_15647,N_15944);
or U19634 (N_19634,N_16781,N_15353);
nand U19635 (N_19635,N_15045,N_16397);
nand U19636 (N_19636,N_16022,N_15575);
nand U19637 (N_19637,N_15463,N_16732);
or U19638 (N_19638,N_16166,N_16647);
or U19639 (N_19639,N_16349,N_17169);
nand U19640 (N_19640,N_17032,N_16861);
nor U19641 (N_19641,N_15305,N_17300);
nand U19642 (N_19642,N_15881,N_15831);
or U19643 (N_19643,N_17060,N_16609);
or U19644 (N_19644,N_15111,N_16460);
nand U19645 (N_19645,N_16443,N_15106);
and U19646 (N_19646,N_15695,N_15778);
and U19647 (N_19647,N_16366,N_16216);
and U19648 (N_19648,N_16235,N_16700);
or U19649 (N_19649,N_16582,N_17172);
xor U19650 (N_19650,N_16993,N_15289);
and U19651 (N_19651,N_17178,N_16882);
nor U19652 (N_19652,N_17340,N_16814);
nor U19653 (N_19653,N_17342,N_15800);
nand U19654 (N_19654,N_17413,N_16753);
nand U19655 (N_19655,N_15874,N_16464);
nor U19656 (N_19656,N_16936,N_16192);
and U19657 (N_19657,N_17131,N_16125);
nor U19658 (N_19658,N_15739,N_16008);
nand U19659 (N_19659,N_17097,N_16653);
and U19660 (N_19660,N_16686,N_16848);
xor U19661 (N_19661,N_16615,N_16589);
and U19662 (N_19662,N_16735,N_16627);
nand U19663 (N_19663,N_15825,N_17289);
nor U19664 (N_19664,N_15090,N_17318);
or U19665 (N_19665,N_16256,N_15700);
xnor U19666 (N_19666,N_16269,N_16970);
or U19667 (N_19667,N_16124,N_16003);
nor U19668 (N_19668,N_16701,N_15023);
xnor U19669 (N_19669,N_16336,N_15159);
or U19670 (N_19670,N_17064,N_16185);
or U19671 (N_19671,N_16124,N_16021);
or U19672 (N_19672,N_17286,N_16739);
nor U19673 (N_19673,N_15343,N_16289);
xnor U19674 (N_19674,N_15690,N_15839);
or U19675 (N_19675,N_15258,N_15674);
nand U19676 (N_19676,N_16848,N_16284);
or U19677 (N_19677,N_15912,N_17304);
nor U19678 (N_19678,N_15719,N_15996);
xnor U19679 (N_19679,N_16932,N_17349);
and U19680 (N_19680,N_16370,N_16778);
nand U19681 (N_19681,N_17215,N_15677);
or U19682 (N_19682,N_16165,N_15749);
and U19683 (N_19683,N_17191,N_17160);
nor U19684 (N_19684,N_15271,N_16644);
or U19685 (N_19685,N_16804,N_15464);
or U19686 (N_19686,N_16329,N_16240);
nand U19687 (N_19687,N_15335,N_15931);
xnor U19688 (N_19688,N_17001,N_15271);
nand U19689 (N_19689,N_15170,N_16822);
nand U19690 (N_19690,N_15490,N_16289);
nor U19691 (N_19691,N_17428,N_16609);
xor U19692 (N_19692,N_15030,N_17136);
or U19693 (N_19693,N_15963,N_15103);
xnor U19694 (N_19694,N_16300,N_16024);
xnor U19695 (N_19695,N_15528,N_15735);
nor U19696 (N_19696,N_17307,N_15290);
xnor U19697 (N_19697,N_16975,N_16235);
and U19698 (N_19698,N_16567,N_15369);
xor U19699 (N_19699,N_15835,N_15946);
or U19700 (N_19700,N_16813,N_15412);
or U19701 (N_19701,N_15435,N_17190);
or U19702 (N_19702,N_15044,N_16921);
xor U19703 (N_19703,N_16279,N_17023);
xor U19704 (N_19704,N_16944,N_16556);
xor U19705 (N_19705,N_16708,N_17286);
xnor U19706 (N_19706,N_15561,N_15199);
nand U19707 (N_19707,N_16453,N_16773);
or U19708 (N_19708,N_16336,N_17487);
and U19709 (N_19709,N_16242,N_17126);
nand U19710 (N_19710,N_17095,N_17333);
or U19711 (N_19711,N_16732,N_17144);
and U19712 (N_19712,N_16631,N_15439);
and U19713 (N_19713,N_16100,N_16366);
xor U19714 (N_19714,N_16754,N_17149);
nor U19715 (N_19715,N_16608,N_16568);
or U19716 (N_19716,N_17245,N_15342);
and U19717 (N_19717,N_17259,N_15673);
nand U19718 (N_19718,N_15626,N_15761);
or U19719 (N_19719,N_16394,N_15818);
nor U19720 (N_19720,N_17176,N_15776);
xor U19721 (N_19721,N_17259,N_16476);
and U19722 (N_19722,N_15105,N_15756);
xor U19723 (N_19723,N_16763,N_15349);
nor U19724 (N_19724,N_16613,N_17249);
and U19725 (N_19725,N_15250,N_16579);
nor U19726 (N_19726,N_16538,N_15094);
and U19727 (N_19727,N_15143,N_16299);
nand U19728 (N_19728,N_16016,N_15023);
nor U19729 (N_19729,N_17153,N_17321);
or U19730 (N_19730,N_17201,N_15496);
or U19731 (N_19731,N_15721,N_16825);
nor U19732 (N_19732,N_16455,N_15879);
and U19733 (N_19733,N_17461,N_15416);
or U19734 (N_19734,N_15794,N_17290);
xnor U19735 (N_19735,N_16278,N_15115);
or U19736 (N_19736,N_15611,N_15752);
or U19737 (N_19737,N_15355,N_17031);
nand U19738 (N_19738,N_15553,N_15600);
and U19739 (N_19739,N_16484,N_16788);
or U19740 (N_19740,N_15297,N_17166);
nor U19741 (N_19741,N_16501,N_15989);
nor U19742 (N_19742,N_16771,N_16273);
and U19743 (N_19743,N_17294,N_15480);
or U19744 (N_19744,N_16577,N_16488);
nor U19745 (N_19745,N_15723,N_15836);
nand U19746 (N_19746,N_15229,N_15044);
nor U19747 (N_19747,N_15067,N_15837);
and U19748 (N_19748,N_16637,N_16390);
or U19749 (N_19749,N_16981,N_17121);
xnor U19750 (N_19750,N_16857,N_16617);
and U19751 (N_19751,N_15391,N_17043);
nor U19752 (N_19752,N_17087,N_17093);
or U19753 (N_19753,N_16972,N_16914);
and U19754 (N_19754,N_15690,N_15075);
nand U19755 (N_19755,N_15561,N_16453);
nor U19756 (N_19756,N_15446,N_17428);
xor U19757 (N_19757,N_16745,N_16201);
or U19758 (N_19758,N_15946,N_16059);
nor U19759 (N_19759,N_15912,N_17493);
nand U19760 (N_19760,N_15752,N_15256);
nand U19761 (N_19761,N_17477,N_16506);
or U19762 (N_19762,N_17339,N_16098);
or U19763 (N_19763,N_16309,N_15985);
nand U19764 (N_19764,N_15202,N_16484);
nor U19765 (N_19765,N_15535,N_17493);
and U19766 (N_19766,N_15368,N_16969);
and U19767 (N_19767,N_16386,N_15501);
or U19768 (N_19768,N_16937,N_16427);
or U19769 (N_19769,N_15027,N_16554);
nor U19770 (N_19770,N_15955,N_16679);
nor U19771 (N_19771,N_15389,N_17406);
and U19772 (N_19772,N_15773,N_15845);
nor U19773 (N_19773,N_16119,N_15022);
and U19774 (N_19774,N_15926,N_15031);
and U19775 (N_19775,N_16562,N_15129);
nand U19776 (N_19776,N_17007,N_15230);
nand U19777 (N_19777,N_15538,N_15854);
xor U19778 (N_19778,N_16603,N_16306);
and U19779 (N_19779,N_15474,N_16122);
nor U19780 (N_19780,N_16124,N_15744);
xor U19781 (N_19781,N_16482,N_16864);
nand U19782 (N_19782,N_16238,N_16827);
nand U19783 (N_19783,N_15471,N_16864);
and U19784 (N_19784,N_16208,N_16222);
and U19785 (N_19785,N_15439,N_15823);
nor U19786 (N_19786,N_16281,N_15975);
nor U19787 (N_19787,N_16624,N_16457);
nor U19788 (N_19788,N_16338,N_17037);
and U19789 (N_19789,N_15961,N_16240);
xnor U19790 (N_19790,N_17334,N_15441);
nand U19791 (N_19791,N_16799,N_16846);
nor U19792 (N_19792,N_17443,N_16428);
or U19793 (N_19793,N_15326,N_15169);
or U19794 (N_19794,N_15198,N_16055);
nand U19795 (N_19795,N_17000,N_16942);
and U19796 (N_19796,N_17362,N_15313);
xor U19797 (N_19797,N_15500,N_16915);
and U19798 (N_19798,N_17465,N_16806);
or U19799 (N_19799,N_15870,N_16219);
nor U19800 (N_19800,N_16597,N_16175);
xor U19801 (N_19801,N_16333,N_16121);
and U19802 (N_19802,N_15990,N_15079);
nor U19803 (N_19803,N_17239,N_16435);
or U19804 (N_19804,N_15696,N_17107);
or U19805 (N_19805,N_16737,N_15295);
xnor U19806 (N_19806,N_16637,N_16618);
xnor U19807 (N_19807,N_16778,N_16960);
or U19808 (N_19808,N_16510,N_16115);
xnor U19809 (N_19809,N_16017,N_17446);
or U19810 (N_19810,N_15981,N_15517);
nand U19811 (N_19811,N_17192,N_15342);
nor U19812 (N_19812,N_15758,N_15558);
nor U19813 (N_19813,N_15721,N_16295);
nand U19814 (N_19814,N_17322,N_16419);
nor U19815 (N_19815,N_15940,N_16393);
and U19816 (N_19816,N_15276,N_15241);
nor U19817 (N_19817,N_16450,N_16806);
nand U19818 (N_19818,N_17366,N_17111);
nor U19819 (N_19819,N_16276,N_15302);
and U19820 (N_19820,N_16647,N_16216);
nand U19821 (N_19821,N_16013,N_16458);
or U19822 (N_19822,N_15560,N_16961);
xor U19823 (N_19823,N_15092,N_17305);
nand U19824 (N_19824,N_15934,N_15795);
nand U19825 (N_19825,N_16314,N_15818);
xor U19826 (N_19826,N_17113,N_16488);
xor U19827 (N_19827,N_16852,N_15685);
and U19828 (N_19828,N_15483,N_16960);
and U19829 (N_19829,N_16019,N_17149);
nand U19830 (N_19830,N_15203,N_15431);
or U19831 (N_19831,N_16756,N_16251);
nand U19832 (N_19832,N_17485,N_15588);
xnor U19833 (N_19833,N_15252,N_17498);
or U19834 (N_19834,N_16470,N_16834);
or U19835 (N_19835,N_16050,N_16953);
nand U19836 (N_19836,N_15157,N_16041);
nor U19837 (N_19837,N_15000,N_15509);
and U19838 (N_19838,N_15770,N_15552);
nand U19839 (N_19839,N_15836,N_16807);
xnor U19840 (N_19840,N_16376,N_16217);
or U19841 (N_19841,N_16217,N_16358);
nand U19842 (N_19842,N_17388,N_17495);
xor U19843 (N_19843,N_17333,N_15498);
xnor U19844 (N_19844,N_17236,N_15486);
nand U19845 (N_19845,N_15669,N_15410);
or U19846 (N_19846,N_16456,N_15347);
xor U19847 (N_19847,N_15850,N_15004);
nor U19848 (N_19848,N_15820,N_16055);
nor U19849 (N_19849,N_15877,N_16594);
or U19850 (N_19850,N_17169,N_16126);
nor U19851 (N_19851,N_16847,N_15338);
xnor U19852 (N_19852,N_16060,N_15244);
and U19853 (N_19853,N_16483,N_16657);
nor U19854 (N_19854,N_15893,N_17052);
xnor U19855 (N_19855,N_16831,N_17052);
nor U19856 (N_19856,N_15668,N_15108);
or U19857 (N_19857,N_17248,N_16783);
nor U19858 (N_19858,N_16676,N_17499);
nand U19859 (N_19859,N_17153,N_15045);
nor U19860 (N_19860,N_17411,N_16112);
nand U19861 (N_19861,N_15740,N_15508);
nand U19862 (N_19862,N_16380,N_16295);
and U19863 (N_19863,N_15227,N_16519);
nand U19864 (N_19864,N_15247,N_17258);
xor U19865 (N_19865,N_17310,N_15776);
and U19866 (N_19866,N_15531,N_15486);
or U19867 (N_19867,N_17411,N_17442);
nor U19868 (N_19868,N_16410,N_16012);
or U19869 (N_19869,N_15150,N_17019);
nor U19870 (N_19870,N_15611,N_15864);
nor U19871 (N_19871,N_15114,N_16738);
nor U19872 (N_19872,N_15481,N_17100);
nand U19873 (N_19873,N_16274,N_16237);
nor U19874 (N_19874,N_15470,N_16154);
nand U19875 (N_19875,N_15560,N_17073);
nor U19876 (N_19876,N_15135,N_16177);
and U19877 (N_19877,N_15769,N_15741);
xnor U19878 (N_19878,N_15646,N_15870);
and U19879 (N_19879,N_17395,N_15891);
xor U19880 (N_19880,N_15168,N_17238);
or U19881 (N_19881,N_15085,N_15203);
or U19882 (N_19882,N_15696,N_15006);
nor U19883 (N_19883,N_16181,N_16058);
nand U19884 (N_19884,N_16288,N_17433);
nand U19885 (N_19885,N_15047,N_16133);
nor U19886 (N_19886,N_16101,N_15134);
or U19887 (N_19887,N_17447,N_15606);
xor U19888 (N_19888,N_15966,N_17306);
or U19889 (N_19889,N_15047,N_15914);
nor U19890 (N_19890,N_15628,N_16931);
nand U19891 (N_19891,N_16372,N_17153);
nor U19892 (N_19892,N_16391,N_17322);
and U19893 (N_19893,N_17186,N_16905);
and U19894 (N_19894,N_15405,N_15721);
nor U19895 (N_19895,N_16118,N_15680);
and U19896 (N_19896,N_15050,N_15906);
and U19897 (N_19897,N_16827,N_17458);
xnor U19898 (N_19898,N_16044,N_15502);
or U19899 (N_19899,N_16405,N_16299);
nor U19900 (N_19900,N_16411,N_16245);
and U19901 (N_19901,N_15674,N_16416);
xnor U19902 (N_19902,N_17267,N_15689);
nor U19903 (N_19903,N_15156,N_15087);
xnor U19904 (N_19904,N_15833,N_17476);
nor U19905 (N_19905,N_16837,N_16965);
or U19906 (N_19906,N_15061,N_17145);
or U19907 (N_19907,N_15258,N_15254);
xor U19908 (N_19908,N_17381,N_15834);
or U19909 (N_19909,N_15494,N_15910);
and U19910 (N_19910,N_16920,N_16672);
and U19911 (N_19911,N_16531,N_16495);
or U19912 (N_19912,N_16005,N_16180);
nor U19913 (N_19913,N_17159,N_16684);
nand U19914 (N_19914,N_15440,N_16032);
and U19915 (N_19915,N_15211,N_15230);
nor U19916 (N_19916,N_15222,N_16378);
nand U19917 (N_19917,N_16490,N_17355);
xnor U19918 (N_19918,N_16179,N_15460);
and U19919 (N_19919,N_15009,N_15218);
nor U19920 (N_19920,N_15899,N_17019);
xor U19921 (N_19921,N_16976,N_16039);
or U19922 (N_19922,N_16403,N_16551);
nor U19923 (N_19923,N_15023,N_16169);
nor U19924 (N_19924,N_16412,N_17138);
nand U19925 (N_19925,N_15018,N_16297);
nand U19926 (N_19926,N_17028,N_16967);
xor U19927 (N_19927,N_17134,N_15481);
nand U19928 (N_19928,N_15913,N_15316);
and U19929 (N_19929,N_15260,N_16489);
nor U19930 (N_19930,N_15258,N_16136);
xor U19931 (N_19931,N_16127,N_16292);
nand U19932 (N_19932,N_15190,N_17366);
nor U19933 (N_19933,N_15961,N_15128);
or U19934 (N_19934,N_16761,N_17326);
nor U19935 (N_19935,N_15498,N_15457);
or U19936 (N_19936,N_15185,N_17412);
xor U19937 (N_19937,N_16877,N_16543);
or U19938 (N_19938,N_16471,N_16139);
nor U19939 (N_19939,N_17307,N_17001);
xnor U19940 (N_19940,N_16270,N_15208);
nand U19941 (N_19941,N_16912,N_15036);
nor U19942 (N_19942,N_16489,N_16393);
nand U19943 (N_19943,N_16913,N_15953);
nor U19944 (N_19944,N_17119,N_15897);
nand U19945 (N_19945,N_17039,N_17267);
or U19946 (N_19946,N_15479,N_16122);
nand U19947 (N_19947,N_16490,N_17386);
and U19948 (N_19948,N_16827,N_16130);
or U19949 (N_19949,N_16083,N_15877);
nand U19950 (N_19950,N_15043,N_17342);
xor U19951 (N_19951,N_15287,N_15146);
or U19952 (N_19952,N_16424,N_15629);
nand U19953 (N_19953,N_16576,N_16374);
nor U19954 (N_19954,N_16415,N_16266);
nor U19955 (N_19955,N_15417,N_16233);
and U19956 (N_19956,N_16768,N_16748);
and U19957 (N_19957,N_16352,N_16087);
xor U19958 (N_19958,N_16607,N_15844);
nor U19959 (N_19959,N_17048,N_16018);
and U19960 (N_19960,N_16714,N_15363);
and U19961 (N_19961,N_16519,N_17285);
or U19962 (N_19962,N_15136,N_16974);
or U19963 (N_19963,N_15793,N_15517);
or U19964 (N_19964,N_15907,N_17059);
nor U19965 (N_19965,N_15263,N_16875);
nand U19966 (N_19966,N_15488,N_15768);
and U19967 (N_19967,N_15780,N_16790);
xnor U19968 (N_19968,N_16704,N_15894);
or U19969 (N_19969,N_17186,N_15802);
and U19970 (N_19970,N_16618,N_15003);
or U19971 (N_19971,N_16186,N_16872);
and U19972 (N_19972,N_16383,N_15651);
or U19973 (N_19973,N_17166,N_16777);
and U19974 (N_19974,N_15731,N_16021);
nor U19975 (N_19975,N_16877,N_16229);
xor U19976 (N_19976,N_15851,N_16217);
nand U19977 (N_19977,N_15434,N_17248);
xor U19978 (N_19978,N_15324,N_16868);
xnor U19979 (N_19979,N_15882,N_16761);
and U19980 (N_19980,N_17047,N_15395);
xnor U19981 (N_19981,N_15729,N_16787);
nor U19982 (N_19982,N_15791,N_16845);
or U19983 (N_19983,N_16024,N_16777);
and U19984 (N_19984,N_16968,N_16916);
nor U19985 (N_19985,N_15029,N_15405);
and U19986 (N_19986,N_15370,N_16255);
xnor U19987 (N_19987,N_17264,N_15807);
nand U19988 (N_19988,N_17301,N_16127);
or U19989 (N_19989,N_15825,N_15332);
or U19990 (N_19990,N_16545,N_15980);
nand U19991 (N_19991,N_16165,N_17072);
xnor U19992 (N_19992,N_16086,N_16442);
and U19993 (N_19993,N_17434,N_16583);
nor U19994 (N_19994,N_16629,N_16055);
and U19995 (N_19995,N_15713,N_15959);
nor U19996 (N_19996,N_16199,N_15224);
and U19997 (N_19997,N_15887,N_15930);
or U19998 (N_19998,N_16990,N_16156);
nor U19999 (N_19999,N_15749,N_15900);
and U20000 (N_20000,N_18143,N_17657);
nand U20001 (N_20001,N_18080,N_18392);
and U20002 (N_20002,N_19761,N_18565);
nor U20003 (N_20003,N_18734,N_18767);
nand U20004 (N_20004,N_18407,N_17866);
nor U20005 (N_20005,N_18519,N_19822);
nor U20006 (N_20006,N_19736,N_19530);
nand U20007 (N_20007,N_19190,N_19378);
or U20008 (N_20008,N_19133,N_19961);
or U20009 (N_20009,N_18712,N_18784);
or U20010 (N_20010,N_19998,N_17585);
nor U20011 (N_20011,N_18893,N_19952);
and U20012 (N_20012,N_18643,N_18016);
nor U20013 (N_20013,N_18679,N_18654);
nand U20014 (N_20014,N_18853,N_18283);
or U20015 (N_20015,N_19446,N_19097);
nor U20016 (N_20016,N_18276,N_19365);
and U20017 (N_20017,N_18810,N_17772);
nand U20018 (N_20018,N_19533,N_17769);
nor U20019 (N_20019,N_18372,N_18668);
nor U20020 (N_20020,N_19629,N_19511);
nand U20021 (N_20021,N_17571,N_19309);
nand U20022 (N_20022,N_18762,N_19211);
nand U20023 (N_20023,N_19785,N_19186);
nand U20024 (N_20024,N_19821,N_19755);
and U20025 (N_20025,N_17629,N_18190);
or U20026 (N_20026,N_19358,N_18239);
and U20027 (N_20027,N_18217,N_18451);
xor U20028 (N_20028,N_19779,N_19687);
or U20029 (N_20029,N_19003,N_18870);
and U20030 (N_20030,N_18349,N_18173);
nor U20031 (N_20031,N_18230,N_17601);
nor U20032 (N_20032,N_17917,N_17622);
or U20033 (N_20033,N_18954,N_19708);
or U20034 (N_20034,N_19644,N_17781);
or U20035 (N_20035,N_18518,N_19974);
nand U20036 (N_20036,N_18901,N_17847);
or U20037 (N_20037,N_19613,N_17596);
and U20038 (N_20038,N_19750,N_17647);
nor U20039 (N_20039,N_19545,N_18562);
nor U20040 (N_20040,N_18161,N_17575);
nor U20041 (N_20041,N_17584,N_19457);
nand U20042 (N_20042,N_18726,N_17790);
or U20043 (N_20043,N_17929,N_19735);
xnor U20044 (N_20044,N_19082,N_19271);
nand U20045 (N_20045,N_17913,N_17993);
and U20046 (N_20046,N_18638,N_17591);
nor U20047 (N_20047,N_19605,N_18076);
xor U20048 (N_20048,N_18699,N_18866);
nor U20049 (N_20049,N_19598,N_17909);
nor U20050 (N_20050,N_18673,N_18412);
and U20051 (N_20051,N_17744,N_18089);
xnor U20052 (N_20052,N_18674,N_18471);
xnor U20053 (N_20053,N_18884,N_19228);
and U20054 (N_20054,N_19017,N_19058);
nor U20055 (N_20055,N_18559,N_19374);
nor U20056 (N_20056,N_19823,N_19321);
or U20057 (N_20057,N_19645,N_17811);
xnor U20058 (N_20058,N_17683,N_17509);
nor U20059 (N_20059,N_17580,N_17655);
xor U20060 (N_20060,N_19329,N_18874);
nor U20061 (N_20061,N_19922,N_17936);
xor U20062 (N_20062,N_19799,N_19224);
and U20063 (N_20063,N_18028,N_18975);
nand U20064 (N_20064,N_19105,N_19999);
xor U20065 (N_20065,N_18871,N_19151);
nand U20066 (N_20066,N_19118,N_18002);
nor U20067 (N_20067,N_18522,N_19559);
nand U20068 (N_20068,N_17882,N_18695);
nand U20069 (N_20069,N_17598,N_19671);
xor U20070 (N_20070,N_18261,N_19023);
nor U20071 (N_20071,N_19618,N_18165);
or U20072 (N_20072,N_19315,N_18065);
xnor U20073 (N_20073,N_17663,N_19754);
or U20074 (N_20074,N_18041,N_18801);
nor U20075 (N_20075,N_19709,N_19425);
and U20076 (N_20076,N_18043,N_17679);
nand U20077 (N_20077,N_19503,N_19656);
nand U20078 (N_20078,N_18444,N_17771);
nor U20079 (N_20079,N_18533,N_18831);
nor U20080 (N_20080,N_18448,N_19883);
nor U20081 (N_20081,N_18434,N_19489);
nor U20082 (N_20082,N_17863,N_18580);
or U20083 (N_20083,N_19440,N_18593);
xor U20084 (N_20084,N_18294,N_19411);
and U20085 (N_20085,N_18129,N_18947);
and U20086 (N_20086,N_19187,N_18828);
xnor U20087 (N_20087,N_17991,N_17524);
xor U20088 (N_20088,N_18716,N_17915);
xor U20089 (N_20089,N_18232,N_17595);
nand U20090 (N_20090,N_18922,N_19371);
nor U20091 (N_20091,N_18855,N_18044);
and U20092 (N_20092,N_18340,N_19609);
nand U20093 (N_20093,N_18697,N_19062);
nand U20094 (N_20094,N_17895,N_18024);
nor U20095 (N_20095,N_19814,N_19432);
nand U20096 (N_20096,N_19292,N_19013);
nand U20097 (N_20097,N_19345,N_18682);
or U20098 (N_20098,N_19188,N_17623);
nand U20099 (N_20099,N_19950,N_19841);
or U20100 (N_20100,N_17904,N_18072);
or U20101 (N_20101,N_17665,N_18493);
or U20102 (N_20102,N_18252,N_19429);
or U20103 (N_20103,N_18182,N_17992);
nand U20104 (N_20104,N_19293,N_19981);
or U20105 (N_20105,N_17688,N_19923);
nand U20106 (N_20106,N_18817,N_19955);
nand U20107 (N_20107,N_18116,N_17540);
xnor U20108 (N_20108,N_19758,N_19124);
and U20109 (N_20109,N_19536,N_19469);
nand U20110 (N_20110,N_19843,N_17971);
nand U20111 (N_20111,N_19653,N_19179);
nor U20112 (N_20112,N_18625,N_18508);
nor U20113 (N_20113,N_19300,N_18030);
xnor U20114 (N_20114,N_18938,N_18620);
nor U20115 (N_20115,N_19091,N_18314);
nand U20116 (N_20116,N_17898,N_18835);
nand U20117 (N_20117,N_18096,N_18888);
xnor U20118 (N_20118,N_19061,N_17833);
nand U20119 (N_20119,N_19453,N_17839);
and U20120 (N_20120,N_17869,N_18147);
and U20121 (N_20121,N_17631,N_17625);
and U20122 (N_20122,N_18704,N_17519);
xnor U20123 (N_20123,N_19126,N_19540);
nand U20124 (N_20124,N_19454,N_18334);
nor U20125 (N_20125,N_19971,N_17633);
nor U20126 (N_20126,N_17919,N_17570);
nor U20127 (N_20127,N_17579,N_18546);
or U20128 (N_20128,N_19339,N_18987);
or U20129 (N_20129,N_17830,N_18589);
nor U20130 (N_20130,N_19128,N_18200);
nand U20131 (N_20131,N_19770,N_19441);
nand U20132 (N_20132,N_18991,N_18951);
nor U20133 (N_20133,N_19220,N_19354);
or U20134 (N_20134,N_17767,N_18369);
nor U20135 (N_20135,N_18007,N_19556);
or U20136 (N_20136,N_17932,N_19278);
xor U20137 (N_20137,N_19256,N_18960);
and U20138 (N_20138,N_19019,N_18093);
or U20139 (N_20139,N_17852,N_18742);
or U20140 (N_20140,N_18282,N_19836);
or U20141 (N_20141,N_19442,N_19793);
and U20142 (N_20142,N_19697,N_19577);
xor U20143 (N_20143,N_19681,N_18541);
and U20144 (N_20144,N_19322,N_18468);
nand U20145 (N_20145,N_19597,N_17953);
and U20146 (N_20146,N_19829,N_19889);
and U20147 (N_20147,N_17567,N_18045);
or U20148 (N_20148,N_19243,N_18743);
nand U20149 (N_20149,N_18733,N_18930);
or U20150 (N_20150,N_18038,N_19016);
nand U20151 (N_20151,N_19415,N_19616);
nor U20152 (N_20152,N_19523,N_17969);
and U20153 (N_20153,N_19934,N_19230);
or U20154 (N_20154,N_17515,N_19980);
and U20155 (N_20155,N_17727,N_17520);
nor U20156 (N_20156,N_19665,N_17930);
and U20157 (N_20157,N_18450,N_18193);
and U20158 (N_20158,N_18957,N_17822);
nor U20159 (N_20159,N_19895,N_19764);
nor U20160 (N_20160,N_19946,N_17713);
and U20161 (N_20161,N_19395,N_18690);
xnor U20162 (N_20162,N_18023,N_18956);
nor U20163 (N_20163,N_19423,N_18356);
nor U20164 (N_20164,N_18184,N_19433);
and U20165 (N_20165,N_19038,N_17548);
nor U20166 (N_20166,N_17711,N_17862);
xor U20167 (N_20167,N_18222,N_19435);
or U20168 (N_20168,N_17805,N_18821);
and U20169 (N_20169,N_17988,N_19943);
or U20170 (N_20170,N_19044,N_18144);
or U20171 (N_20171,N_18621,N_18213);
nor U20172 (N_20172,N_18359,N_19740);
nor U20173 (N_20173,N_18949,N_18219);
and U20174 (N_20174,N_19674,N_19775);
and U20175 (N_20175,N_19888,N_18231);
nand U20176 (N_20176,N_19192,N_18179);
nor U20177 (N_20177,N_18121,N_17561);
and U20178 (N_20178,N_18698,N_19175);
or U20179 (N_20179,N_18770,N_18862);
or U20180 (N_20180,N_19449,N_18148);
nand U20181 (N_20181,N_18812,N_17517);
nor U20182 (N_20182,N_18603,N_19257);
or U20183 (N_20183,N_17998,N_19407);
nor U20184 (N_20184,N_19658,N_19581);
nor U20185 (N_20185,N_19153,N_18727);
nand U20186 (N_20186,N_18268,N_19221);
and U20187 (N_20187,N_19201,N_17942);
nor U20188 (N_20188,N_18145,N_19650);
nand U20189 (N_20189,N_17808,N_17610);
or U20190 (N_20190,N_17944,N_19729);
and U20191 (N_20191,N_19833,N_19619);
nor U20192 (N_20192,N_18858,N_18623);
or U20193 (N_20193,N_18516,N_17947);
nor U20194 (N_20194,N_19076,N_18504);
xnor U20195 (N_20195,N_19504,N_18378);
xnor U20196 (N_20196,N_17533,N_19621);
nor U20197 (N_20197,N_19839,N_18525);
xnor U20198 (N_20198,N_19759,N_18284);
and U20199 (N_20199,N_19984,N_18178);
nor U20200 (N_20200,N_18223,N_17941);
nand U20201 (N_20201,N_18891,N_17576);
nor U20202 (N_20202,N_19342,N_17565);
or U20203 (N_20203,N_18181,N_18249);
or U20204 (N_20204,N_18502,N_18384);
nor U20205 (N_20205,N_18062,N_18234);
xor U20206 (N_20206,N_17568,N_18458);
and U20207 (N_20207,N_18013,N_19002);
or U20208 (N_20208,N_19370,N_18786);
and U20209 (N_20209,N_19343,N_19679);
or U20210 (N_20210,N_17981,N_17554);
nand U20211 (N_20211,N_17880,N_18146);
or U20212 (N_20212,N_19462,N_19314);
and U20213 (N_20213,N_19108,N_19957);
or U20214 (N_20214,N_18296,N_18218);
nor U20215 (N_20215,N_19526,N_18348);
xnor U20216 (N_20216,N_18246,N_19040);
or U20217 (N_20217,N_17597,N_17583);
and U20218 (N_20218,N_19255,N_19788);
and U20219 (N_20219,N_17968,N_19845);
or U20220 (N_20220,N_18629,N_18578);
nor U20221 (N_20221,N_18832,N_19419);
nand U20222 (N_20222,N_19751,N_18887);
or U20223 (N_20223,N_18577,N_17525);
nor U20224 (N_20224,N_19068,N_18609);
nor U20225 (N_20225,N_17518,N_19828);
nor U20226 (N_20226,N_19313,N_19529);
xor U20227 (N_20227,N_18180,N_18467);
nor U20228 (N_20228,N_19887,N_18039);
nand U20229 (N_20229,N_19877,N_19401);
xnor U20230 (N_20230,N_19452,N_19033);
nand U20231 (N_20231,N_18160,N_19916);
and U20232 (N_20232,N_17994,N_19564);
xor U20233 (N_20233,N_18520,N_17938);
or U20234 (N_20234,N_19612,N_17838);
nor U20235 (N_20235,N_17974,N_17723);
xnor U20236 (N_20236,N_17812,N_19000);
nor U20237 (N_20237,N_19047,N_18354);
xnor U20238 (N_20238,N_18605,N_19900);
and U20239 (N_20239,N_19475,N_19647);
xnor U20240 (N_20240,N_18739,N_18355);
xnor U20241 (N_20241,N_17757,N_17680);
or U20242 (N_20242,N_17877,N_18119);
xnor U20243 (N_20243,N_19007,N_19404);
nand U20244 (N_20244,N_19131,N_18996);
and U20245 (N_20245,N_18736,N_17678);
nand U20246 (N_20246,N_18303,N_18807);
or U20247 (N_20247,N_19603,N_18390);
or U20248 (N_20248,N_18191,N_17756);
xor U20249 (N_20249,N_17761,N_17694);
and U20250 (N_20250,N_17910,N_19431);
nor U20251 (N_20251,N_18462,N_19140);
xnor U20252 (N_20252,N_18311,N_17762);
and U20253 (N_20253,N_17807,N_18971);
or U20254 (N_20254,N_19800,N_18436);
nand U20255 (N_20255,N_19566,N_18313);
nand U20256 (N_20256,N_18936,N_19194);
nand U20257 (N_20257,N_17527,N_18758);
nand U20258 (N_20258,N_18694,N_17965);
or U20259 (N_20259,N_17796,N_17724);
or U20260 (N_20260,N_17687,N_17604);
nor U20261 (N_20261,N_19393,N_18657);
and U20262 (N_20262,N_19072,N_18842);
nor U20263 (N_20263,N_19592,N_19661);
xnor U20264 (N_20264,N_18564,N_18970);
and U20265 (N_20265,N_18464,N_18396);
and U20266 (N_20266,N_17948,N_17513);
and U20267 (N_20267,N_19020,N_19218);
nand U20268 (N_20268,N_19333,N_18513);
and U20269 (N_20269,N_19515,N_18479);
nand U20270 (N_20270,N_18337,N_19599);
xnor U20271 (N_20271,N_18243,N_17645);
or U20272 (N_20272,N_19947,N_19326);
or U20273 (N_20273,N_19848,N_18398);
xor U20274 (N_20274,N_18924,N_17977);
nand U20275 (N_20275,N_19477,N_18466);
and U20276 (N_20276,N_19702,N_18262);
or U20277 (N_20277,N_18584,N_18964);
nor U20278 (N_20278,N_18641,N_19274);
xnor U20279 (N_20279,N_17939,N_17721);
and U20280 (N_20280,N_18935,N_17502);
or U20281 (N_20281,N_18574,N_18900);
nand U20282 (N_20282,N_18633,N_18492);
nand U20283 (N_20283,N_18644,N_18585);
nor U20284 (N_20284,N_18630,N_19250);
and U20285 (N_20285,N_18804,N_18523);
or U20286 (N_20286,N_18321,N_17765);
nand U20287 (N_20287,N_18550,N_19884);
or U20288 (N_20288,N_19282,N_17739);
or U20289 (N_20289,N_19390,N_18320);
or U20290 (N_20290,N_18894,N_19853);
xnor U20291 (N_20291,N_18221,N_18664);
or U20292 (N_20292,N_18310,N_19593);
xnor U20293 (N_20293,N_19579,N_17809);
xnor U20294 (N_20294,N_19289,N_19199);
nor U20295 (N_20295,N_17891,N_18588);
nand U20296 (N_20296,N_17656,N_18686);
nor U20297 (N_20297,N_17973,N_19109);
nor U20298 (N_20298,N_17737,N_18558);
or U20299 (N_20299,N_19649,N_19036);
nor U20300 (N_20300,N_18059,N_18174);
nor U20301 (N_20301,N_19630,N_19772);
nor U20302 (N_20302,N_19311,N_17729);
and U20303 (N_20303,N_18087,N_19268);
xor U20304 (N_20304,N_18576,N_17682);
xnor U20305 (N_20305,N_17886,N_19483);
nand U20306 (N_20306,N_18732,N_19026);
or U20307 (N_20307,N_18381,N_19659);
and U20308 (N_20308,N_19569,N_18999);
nand U20309 (N_20309,N_17726,N_19486);
nand U20310 (N_20310,N_17792,N_18435);
and U20311 (N_20311,N_19892,N_18825);
nor U20312 (N_20312,N_19451,N_17900);
nor U20313 (N_20313,N_19997,N_19905);
nor U20314 (N_20314,N_17677,N_18452);
xor U20315 (N_20315,N_18809,N_19870);
and U20316 (N_20316,N_18984,N_19120);
nand U20317 (N_20317,N_18805,N_18319);
and U20318 (N_20318,N_18328,N_19302);
xnor U20319 (N_20319,N_18104,N_19193);
and U20320 (N_20320,N_17572,N_19233);
nand U20321 (N_20321,N_18102,N_19636);
or U20322 (N_20322,N_17701,N_18338);
xor U20323 (N_20323,N_18912,N_18292);
nor U20324 (N_20324,N_19863,N_19854);
nor U20325 (N_20325,N_19111,N_19917);
xnor U20326 (N_20326,N_19262,N_18731);
nand U20327 (N_20327,N_19139,N_17843);
and U20328 (N_20328,N_19757,N_18106);
xor U20329 (N_20329,N_19100,N_19626);
nand U20330 (N_20330,N_19163,N_18815);
xor U20331 (N_20331,N_19488,N_18245);
nand U20332 (N_20332,N_19275,N_19318);
and U20333 (N_20333,N_18800,N_19926);
nand U20334 (N_20334,N_17921,N_18608);
nand U20335 (N_20335,N_18989,N_17528);
nand U20336 (N_20336,N_17635,N_19229);
and U20337 (N_20337,N_19214,N_18031);
or U20338 (N_20338,N_19063,N_19509);
or U20339 (N_20339,N_18109,N_19149);
nor U20340 (N_20340,N_18819,N_18177);
and U20341 (N_20341,N_18130,N_19090);
nand U20342 (N_20342,N_19741,N_18424);
and U20343 (N_20343,N_18696,N_18210);
or U20344 (N_20344,N_18676,N_19198);
xor U20345 (N_20345,N_19572,N_17608);
nand U20346 (N_20346,N_18204,N_17658);
nand U20347 (N_20347,N_18306,N_18791);
nand U20348 (N_20348,N_18683,N_18943);
and U20349 (N_20349,N_17763,N_18868);
or U20350 (N_20350,N_18105,N_17532);
nand U20351 (N_20351,N_18684,N_19573);
xor U20352 (N_20352,N_19876,N_19930);
xor U20353 (N_20353,N_19913,N_17854);
or U20354 (N_20354,N_18881,N_17643);
or U20355 (N_20355,N_19362,N_17885);
nand U20356 (N_20356,N_18138,N_18404);
xor U20357 (N_20357,N_19104,N_19882);
nand U20358 (N_20358,N_18175,N_19516);
nor U20359 (N_20359,N_19001,N_18837);
xor U20360 (N_20360,N_18702,N_18803);
xnor U20361 (N_20361,N_18503,N_17976);
xor U20362 (N_20362,N_19535,N_18430);
nand U20363 (N_20363,N_18665,N_19723);
nand U20364 (N_20364,N_18032,N_19767);
and U20365 (N_20365,N_18267,N_19051);
xnor U20366 (N_20366,N_19168,N_18266);
nor U20367 (N_20367,N_19157,N_19648);
xor U20368 (N_20368,N_18092,N_17881);
or U20369 (N_20369,N_19812,N_19906);
and U20370 (N_20370,N_18042,N_18961);
xnor U20371 (N_20371,N_18409,N_18538);
and U20372 (N_20372,N_18136,N_17523);
nand U20373 (N_20373,N_19651,N_18350);
nor U20374 (N_20374,N_19156,N_19587);
nor U20375 (N_20375,N_18838,N_19398);
nor U20376 (N_20376,N_19541,N_19524);
or U20377 (N_20377,N_17864,N_19748);
nand U20378 (N_20378,N_19677,N_17884);
and U20379 (N_20379,N_19539,N_17578);
and U20380 (N_20380,N_18473,N_18167);
nand U20381 (N_20381,N_17818,N_19964);
xor U20382 (N_20382,N_17791,N_19144);
nand U20383 (N_20383,N_18823,N_19045);
nor U20384 (N_20384,N_19819,N_18126);
xor U20385 (N_20385,N_17960,N_19065);
nand U20386 (N_20386,N_18774,N_18952);
nand U20387 (N_20387,N_18711,N_17990);
nor U20388 (N_20388,N_18046,N_17937);
or U20389 (N_20389,N_17594,N_18188);
xor U20390 (N_20390,N_18555,N_18923);
xnor U20391 (N_20391,N_17972,N_19507);
xnor U20392 (N_20392,N_19127,N_17703);
nor U20393 (N_20393,N_17605,N_19437);
or U20394 (N_20394,N_17779,N_19041);
xnor U20395 (N_20395,N_19739,N_19915);
xor U20396 (N_20396,N_17616,N_19513);
nand U20397 (N_20397,N_19304,N_18457);
or U20398 (N_20398,N_19253,N_19388);
xnor U20399 (N_20399,N_19207,N_18848);
nand U20400 (N_20400,N_17624,N_19238);
and U20401 (N_20401,N_18826,N_17755);
nand U20402 (N_20402,N_18759,N_18818);
nand U20403 (N_20403,N_17603,N_18291);
xnor U20404 (N_20404,N_19944,N_18199);
nor U20405 (N_20405,N_19975,N_18652);
or U20406 (N_20406,N_19624,N_19319);
nand U20407 (N_20407,N_19548,N_17943);
and U20408 (N_20408,N_19176,N_17975);
nand U20409 (N_20409,N_18864,N_18708);
nand U20410 (N_20410,N_19791,N_19032);
nor U20411 (N_20411,N_17883,N_19424);
nor U20412 (N_20412,N_19578,N_19574);
and U20413 (N_20413,N_17835,N_18709);
or U20414 (N_20414,N_19147,N_19991);
or U20415 (N_20415,N_19412,N_19938);
or U20416 (N_20416,N_17670,N_18680);
xnor U20417 (N_20417,N_18005,N_17933);
xnor U20418 (N_20418,N_19846,N_18055);
and U20419 (N_20419,N_18972,N_19286);
nand U20420 (N_20420,N_17710,N_18744);
xnor U20421 (N_20421,N_18751,N_19078);
nand U20422 (N_20422,N_17950,N_18738);
nand U20423 (N_20423,N_18012,N_19356);
or U20424 (N_20424,N_17815,N_19323);
nand U20425 (N_20425,N_18714,N_18557);
and U20426 (N_20426,N_18678,N_18681);
xor U20427 (N_20427,N_18248,N_19869);
nor U20428 (N_20428,N_19405,N_19896);
and U20429 (N_20429,N_18391,N_17699);
xor U20430 (N_20430,N_17510,N_17979);
or U20431 (N_20431,N_18808,N_17743);
and U20432 (N_20432,N_19949,N_19347);
nor U20433 (N_20433,N_18981,N_18427);
and U20434 (N_20434,N_18250,N_18419);
nor U20435 (N_20435,N_18710,N_17555);
nand U20436 (N_20436,N_17742,N_17868);
or U20437 (N_20437,N_17961,N_18082);
and U20438 (N_20438,N_18554,N_19350);
xnor U20439 (N_20439,N_18365,N_19602);
nor U20440 (N_20440,N_17607,N_19396);
nor U20441 (N_20441,N_19792,N_18986);
nor U20442 (N_20442,N_17639,N_18216);
nand U20443 (N_20443,N_19831,N_18685);
nand U20444 (N_20444,N_18207,N_18021);
nand U20445 (N_20445,N_19400,N_18241);
xor U20446 (N_20446,N_19382,N_18084);
or U20447 (N_20447,N_19506,N_19549);
and U20448 (N_20448,N_19461,N_19561);
nor U20449 (N_20449,N_19240,N_19379);
and U20450 (N_20450,N_19355,N_18247);
or U20451 (N_20451,N_18280,N_19258);
and U20452 (N_20452,N_17716,N_19988);
xor U20453 (N_20453,N_18344,N_17501);
nand U20454 (N_20454,N_18095,N_18439);
xor U20455 (N_20455,N_19482,N_18902);
nand U20456 (N_20456,N_19673,N_18364);
and U20457 (N_20457,N_18877,N_18067);
and U20458 (N_20458,N_19746,N_17897);
xor U20459 (N_20459,N_18187,N_19633);
or U20460 (N_20460,N_19264,N_18861);
xnor U20461 (N_20461,N_18061,N_18691);
nand U20462 (N_20462,N_18257,N_17887);
or U20463 (N_20463,N_18865,N_18950);
nand U20464 (N_20464,N_19583,N_19886);
and U20465 (N_20465,N_18273,N_17507);
and U20466 (N_20466,N_19209,N_19614);
or U20467 (N_20467,N_17700,N_18839);
or U20468 (N_20468,N_18152,N_18103);
and U20469 (N_20469,N_19987,N_19325);
and U20470 (N_20470,N_17764,N_18166);
nor U20471 (N_20471,N_19685,N_18033);
or U20472 (N_20472,N_19570,N_19641);
and U20473 (N_20473,N_18526,N_18967);
or U20474 (N_20474,N_18373,N_19890);
nor U20475 (N_20475,N_19150,N_18052);
or U20476 (N_20476,N_19805,N_18570);
nor U20477 (N_20477,N_18383,N_17987);
nand U20478 (N_20478,N_18368,N_18153);
xor U20479 (N_20479,N_19861,N_19180);
nand U20480 (N_20480,N_19024,N_19083);
nand U20481 (N_20481,N_17731,N_19171);
xnor U20482 (N_20482,N_19181,N_18753);
xnor U20483 (N_20483,N_18869,N_17931);
xnor U20484 (N_20484,N_18057,N_18761);
and U20485 (N_20485,N_19196,N_19901);
nand U20486 (N_20486,N_17628,N_19450);
xnor U20487 (N_20487,N_18966,N_18913);
nor U20488 (N_20488,N_19920,N_18772);
nor U20489 (N_20489,N_17732,N_17752);
nand U20490 (N_20490,N_19776,N_17542);
nand U20491 (N_20491,N_19459,N_18854);
nor U20492 (N_20492,N_19306,N_18561);
nor U20493 (N_20493,N_18393,N_17735);
or U20494 (N_20494,N_18551,N_19727);
nor U20495 (N_20495,N_18485,N_19928);
nor U20496 (N_20496,N_18534,N_19472);
xnor U20497 (N_20497,N_18488,N_17952);
nand U20498 (N_20498,N_19141,N_18982);
and U20499 (N_20499,N_18658,N_19012);
xor U20500 (N_20500,N_18196,N_18075);
nand U20501 (N_20501,N_17892,N_18494);
nor U20502 (N_20502,N_17696,N_17559);
or U20503 (N_20503,N_18445,N_18414);
nor U20504 (N_20504,N_17827,N_18380);
or U20505 (N_20505,N_19361,N_18164);
xnor U20506 (N_20506,N_18163,N_19115);
and U20507 (N_20507,N_19352,N_18244);
nand U20508 (N_20508,N_18937,N_19931);
nand U20509 (N_20509,N_18070,N_17521);
nor U20510 (N_20510,N_18358,N_17956);
or U20511 (N_20511,N_18054,N_19639);
or U20512 (N_20512,N_18026,N_19704);
nor U20513 (N_20513,N_19035,N_17935);
xor U20514 (N_20514,N_18777,N_19699);
xor U20515 (N_20515,N_19978,N_17853);
and U20516 (N_20516,N_18940,N_18640);
or U20517 (N_20517,N_19011,N_19114);
or U20518 (N_20518,N_17780,N_19288);
or U20519 (N_20519,N_19308,N_19490);
xnor U20520 (N_20520,N_18018,N_19344);
nor U20521 (N_20521,N_17775,N_18719);
and U20522 (N_20522,N_19635,N_17845);
xor U20523 (N_20523,N_19208,N_19413);
nor U20524 (N_20524,N_19226,N_18512);
or U20525 (N_20525,N_17544,N_18139);
or U20526 (N_20526,N_17758,N_17661);
or U20527 (N_20527,N_19303,N_19856);
nand U20528 (N_20528,N_19427,N_18617);
and U20529 (N_20529,N_19738,N_17745);
or U20530 (N_20530,N_19341,N_19670);
nand U20531 (N_20531,N_19086,N_19103);
or U20532 (N_20532,N_19711,N_19722);
nor U20533 (N_20533,N_19668,N_19242);
nor U20534 (N_20534,N_18019,N_18860);
or U20535 (N_20535,N_18659,N_17673);
or U20536 (N_20536,N_19919,N_18737);
nand U20537 (N_20537,N_19688,N_17650);
or U20538 (N_20538,N_17824,N_17782);
nand U20539 (N_20539,N_17773,N_17671);
nor U20540 (N_20540,N_18740,N_18125);
nor U20541 (N_20541,N_18360,N_18499);
nand U20542 (N_20542,N_18226,N_19716);
and U20543 (N_20543,N_19239,N_19173);
or U20544 (N_20544,N_19125,N_19122);
and U20545 (N_20545,N_17800,N_17834);
xnor U20546 (N_20546,N_17707,N_17849);
and U20547 (N_20547,N_17719,N_17664);
and U20548 (N_20548,N_19119,N_19055);
nand U20549 (N_20549,N_19801,N_18915);
nand U20550 (N_20550,N_19745,N_17653);
or U20551 (N_20551,N_17672,N_17747);
or U20552 (N_20552,N_19728,N_19628);
xnor U20553 (N_20553,N_17995,N_19070);
nor U20554 (N_20554,N_18426,N_17865);
nand U20555 (N_20555,N_18845,N_19678);
or U20556 (N_20556,N_17529,N_18829);
and U20557 (N_20557,N_18361,N_19021);
and U20558 (N_20558,N_18903,N_19682);
and U20559 (N_20559,N_18718,N_19734);
nor U20560 (N_20560,N_18980,N_19492);
nor U20561 (N_20561,N_19560,N_19977);
xnor U20562 (N_20562,N_18571,N_18212);
xor U20563 (N_20563,N_18497,N_17530);
xnor U20564 (N_20564,N_18081,N_19376);
xor U20565 (N_20565,N_19835,N_19137);
nand U20566 (N_20566,N_18600,N_18788);
nand U20567 (N_20567,N_19460,N_19696);
or U20568 (N_20568,N_17872,N_19172);
nor U20569 (N_20569,N_18521,N_17927);
xnor U20570 (N_20570,N_18496,N_18581);
or U20571 (N_20571,N_17632,N_17798);
and U20572 (N_20572,N_18487,N_18863);
or U20573 (N_20573,N_18265,N_19695);
nand U20574 (N_20574,N_19582,N_18242);
nand U20575 (N_20575,N_18706,N_19527);
xnor U20576 (N_20576,N_18532,N_19005);
and U20577 (N_20577,N_19710,N_19471);
nand U20578 (N_20578,N_18529,N_18655);
nand U20579 (N_20579,N_19970,N_19837);
nor U20580 (N_20580,N_18651,N_18675);
xor U20581 (N_20581,N_19331,N_18723);
nand U20582 (N_20582,N_19006,N_18269);
nor U20583 (N_20583,N_18477,N_18615);
or U20584 (N_20584,N_19528,N_19443);
and U20585 (N_20585,N_19204,N_19079);
nor U20586 (N_20586,N_17674,N_18189);
nor U20587 (N_20587,N_19053,N_19134);
nand U20588 (N_20588,N_19046,N_19054);
or U20589 (N_20589,N_17582,N_18820);
and U20590 (N_20590,N_18274,N_18509);
and U20591 (N_20591,N_17718,N_17557);
xnor U20592 (N_20592,N_19766,N_19543);
or U20593 (N_20593,N_17543,N_18009);
nand U20594 (N_20594,N_18293,N_17846);
or U20595 (N_20595,N_17651,N_19074);
nand U20596 (N_20596,N_19731,N_17534);
nor U20597 (N_20597,N_17712,N_19244);
nor U20598 (N_20598,N_17870,N_18645);
or U20599 (N_20599,N_19334,N_18846);
nand U20600 (N_20600,N_19908,N_18185);
or U20601 (N_20601,N_18836,N_19241);
and U20602 (N_20602,N_18128,N_19121);
or U20603 (N_20603,N_17828,N_18305);
or U20604 (N_20604,N_19925,N_17954);
nand U20605 (N_20605,N_18456,N_18498);
or U20606 (N_20606,N_19620,N_17871);
and U20607 (N_20607,N_17506,N_19279);
nor U20608 (N_20608,N_18785,N_19899);
nand U20609 (N_20609,N_19634,N_17722);
or U20610 (N_20610,N_18834,N_18780);
and U20611 (N_20611,N_19254,N_18064);
nor U20612 (N_20612,N_19167,N_19010);
or U20613 (N_20613,N_17778,N_18208);
and U20614 (N_20614,N_19669,N_17541);
and U20615 (N_20615,N_19584,N_19525);
nand U20616 (N_20616,N_19718,N_19717);
xnor U20617 (N_20617,N_18386,N_18850);
and U20618 (N_20618,N_18299,N_19760);
nor U20619 (N_20619,N_17702,N_19232);
or U20620 (N_20620,N_18636,N_19375);
xor U20621 (N_20621,N_19468,N_19742);
nand U20622 (N_20622,N_18990,N_19898);
nand U20623 (N_20623,N_18978,N_18123);
and U20624 (N_20624,N_18206,N_17894);
nand U20625 (N_20625,N_18979,N_17685);
nand U20626 (N_20626,N_17906,N_19715);
nand U20627 (N_20627,N_19165,N_19298);
nor U20628 (N_20628,N_18432,N_19087);
nor U20629 (N_20629,N_19030,N_18689);
xnor U20630 (N_20630,N_19249,N_19519);
nor U20631 (N_20631,N_19265,N_19684);
nor U20632 (N_20632,N_18056,N_18725);
or U20633 (N_20633,N_19458,N_19774);
nor U20634 (N_20634,N_19807,N_19713);
nand U20635 (N_20635,N_19394,N_19847);
nand U20636 (N_20636,N_17648,N_18921);
xnor U20637 (N_20637,N_19166,N_19495);
or U20638 (N_20638,N_19769,N_19842);
nor U20639 (N_20639,N_18151,N_18069);
nor U20640 (N_20640,N_17748,N_17989);
nand U20641 (N_20641,N_19518,N_17888);
xnor U20642 (N_20642,N_19806,N_17801);
and U20643 (N_20643,N_19098,N_17831);
and U20644 (N_20644,N_18263,N_18671);
and U20645 (N_20645,N_19392,N_17705);
and U20646 (N_20646,N_18346,N_19595);
nor U20647 (N_20647,N_18931,N_19505);
xnor U20648 (N_20648,N_18566,N_19048);
and U20649 (N_20649,N_19034,N_19744);
or U20650 (N_20650,N_18677,N_19826);
nor U20651 (N_20651,N_18766,N_18648);
or U20652 (N_20652,N_18073,N_19478);
nor U20653 (N_20653,N_17613,N_17599);
or U20654 (N_20654,N_17982,N_19247);
or U20655 (N_20655,N_19691,N_17770);
nand U20656 (N_20656,N_19816,N_18911);
or U20657 (N_20657,N_18347,N_19600);
nor U20658 (N_20658,N_18667,N_18653);
nand U20659 (N_20659,N_19191,N_17826);
nor U20660 (N_20660,N_17776,N_17511);
or U20661 (N_20661,N_19485,N_19042);
nand U20662 (N_20662,N_19797,N_18460);
or U20663 (N_20663,N_17612,N_17660);
and U20664 (N_20664,N_17814,N_18079);
nor U20665 (N_20665,N_17636,N_19290);
nand U20666 (N_20666,N_18569,N_18131);
or U20667 (N_20667,N_17785,N_19773);
and U20668 (N_20668,N_18783,N_18822);
xor U20669 (N_20669,N_17615,N_17905);
nor U20670 (N_20670,N_19712,N_17500);
xnor U20671 (N_20671,N_19855,N_19297);
xnor U20672 (N_20672,N_18169,N_17573);
and U20673 (N_20673,N_18757,N_19552);
or U20674 (N_20674,N_19640,N_17574);
or U20675 (N_20675,N_18335,N_18524);
xor U20676 (N_20676,N_19312,N_19986);
xnor U20677 (N_20677,N_19263,N_18475);
nand U20678 (N_20678,N_19107,N_18339);
nand U20679 (N_20679,N_18939,N_18323);
nand U20680 (N_20680,N_18048,N_18352);
or U20681 (N_20681,N_19164,N_18309);
or U20682 (N_20682,N_18549,N_19520);
xor U20683 (N_20683,N_19940,N_19692);
nand U20684 (N_20684,N_18379,N_18469);
and U20685 (N_20685,N_19840,N_19962);
nand U20686 (N_20686,N_19830,N_18539);
xnor U20687 (N_20687,N_18672,N_19409);
and U20688 (N_20688,N_18341,N_18530);
nand U20689 (N_20689,N_17819,N_19236);
xnor U20690 (N_20690,N_18480,N_19060);
xnor U20691 (N_20691,N_19660,N_18531);
or U20692 (N_20692,N_18195,N_18150);
nand U20693 (N_20693,N_19367,N_19148);
or U20694 (N_20694,N_17816,N_19844);
or U20695 (N_20695,N_17691,N_17963);
nand U20696 (N_20696,N_18317,N_17955);
xnor U20697 (N_20697,N_18371,N_18211);
nor U20698 (N_20698,N_18097,N_18505);
nand U20699 (N_20699,N_19532,N_18316);
and U20700 (N_20700,N_18490,N_18332);
or U20701 (N_20701,N_18878,N_18162);
nor U20702 (N_20702,N_18500,N_19075);
or U20703 (N_20703,N_19652,N_18110);
nand U20704 (N_20704,N_19422,N_18308);
or U20705 (N_20705,N_17926,N_19299);
xnor U20706 (N_20706,N_19749,N_17549);
and U20707 (N_20707,N_19123,N_17978);
nor U20708 (N_20708,N_17788,N_19498);
and U20709 (N_20709,N_19170,N_18168);
nand U20710 (N_20710,N_18394,N_18318);
or U20711 (N_20711,N_18120,N_19102);
nand U20712 (N_20712,N_18433,N_18304);
and U20713 (N_20713,N_18049,N_18916);
or U20714 (N_20714,N_18259,N_17786);
nand U20715 (N_20715,N_19571,N_19248);
xor U20716 (N_20716,N_19225,N_19818);
nand U20717 (N_20717,N_18973,N_17536);
or U20718 (N_20718,N_19765,N_18399);
xnor U20719 (N_20719,N_18437,N_19195);
nor U20720 (N_20720,N_18553,N_19714);
or U20721 (N_20721,N_18068,N_17802);
nor U20722 (N_20722,N_19958,N_17638);
nor U20723 (N_20723,N_18688,N_19756);
or U20724 (N_20724,N_19996,N_17508);
or U20725 (N_20725,N_19627,N_19227);
nor U20726 (N_20726,N_19939,N_18214);
and U20727 (N_20727,N_19317,N_19733);
nor U20728 (N_20728,N_18745,N_19064);
and U20729 (N_20729,N_18662,N_19663);
xnor U20730 (N_20730,N_19878,N_19284);
nor U20731 (N_20731,N_18944,N_19436);
xnor U20732 (N_20732,N_18254,N_19834);
nor U20733 (N_20733,N_18856,N_18256);
and U20734 (N_20734,N_19130,N_18833);
or U20735 (N_20735,N_18429,N_19081);
nand U20736 (N_20736,N_18724,N_18000);
xnor U20737 (N_20737,N_18085,N_17999);
nor U20738 (N_20738,N_18882,N_18778);
nand U20739 (N_20739,N_19049,N_18802);
nor U20740 (N_20740,N_19662,N_18573);
and U20741 (N_20741,N_19782,N_18568);
xnor U20742 (N_20742,N_19666,N_19270);
or U20743 (N_20743,N_19360,N_18506);
nand U20744 (N_20744,N_18896,N_17654);
or U20745 (N_20745,N_17569,N_19169);
and U20746 (N_20746,N_18906,N_18277);
nand U20747 (N_20747,N_18425,N_19676);
nand U20748 (N_20748,N_18071,N_18983);
nor U20749 (N_20749,N_19448,N_19637);
or U20750 (N_20750,N_19643,N_19631);
and U20751 (N_20751,N_19106,N_19402);
nand U20752 (N_20752,N_17889,N_18816);
nor U20753 (N_20753,N_19719,N_18976);
xor U20754 (N_20754,N_18851,N_18118);
and U20755 (N_20755,N_18591,N_18094);
nand U20756 (N_20756,N_19056,N_19683);
nor U20757 (N_20757,N_18765,N_18773);
nor U20758 (N_20758,N_18406,N_17626);
xor U20759 (N_20759,N_18388,N_18074);
nand U20760 (N_20760,N_18730,N_19617);
and U20761 (N_20761,N_17551,N_19787);
nor U20762 (N_20762,N_19512,N_19992);
or U20763 (N_20763,N_17630,N_18198);
and U20764 (N_20764,N_18370,N_19491);
and U20765 (N_20765,N_18376,N_17617);
nor U20766 (N_20766,N_19080,N_19494);
or U20767 (N_20767,N_19976,N_18985);
or U20768 (N_20768,N_19348,N_18992);
xnor U20769 (N_20769,N_17602,N_17704);
and U20770 (N_20770,N_19784,N_18728);
nand U20771 (N_20771,N_18363,N_18717);
nand U20772 (N_20772,N_18579,N_19794);
nor U20773 (N_20773,N_19726,N_18463);
and U20774 (N_20774,N_18582,N_19990);
nor U20775 (N_20775,N_19953,N_18227);
nand U20776 (N_20776,N_18544,N_19789);
xor U20777 (N_20777,N_18928,N_17740);
nor U20778 (N_20778,N_17531,N_18618);
and U20779 (N_20779,N_17690,N_19096);
xor U20780 (N_20780,N_18417,N_19825);
nand U20781 (N_20781,N_18117,N_18050);
nand U20782 (N_20782,N_18597,N_17985);
xor U20783 (N_20783,N_18287,N_19389);
and U20784 (N_20784,N_18183,N_19933);
nor U20785 (N_20785,N_19657,N_19827);
or U20786 (N_20786,N_17851,N_19576);
or U20787 (N_20787,N_17940,N_18760);
and U20788 (N_20788,N_18020,N_17908);
and U20789 (N_20789,N_19349,N_18843);
xnor U20790 (N_20790,N_18501,N_18051);
nand U20791 (N_20791,N_18635,N_19363);
or U20792 (N_20792,N_19655,N_18631);
and U20793 (N_20793,N_19132,N_19979);
nand U20794 (N_20794,N_18953,N_18289);
nand U20795 (N_20795,N_19879,N_18022);
xnor U20796 (N_20796,N_19385,N_19880);
and U20797 (N_20797,N_19099,N_17560);
xnor U20798 (N_20798,N_18910,N_19408);
xnor U20799 (N_20799,N_18890,N_19296);
or U20800 (N_20800,N_19780,N_18171);
nand U20801 (N_20801,N_19089,N_18789);
or U20802 (N_20802,N_18873,N_17934);
nand U20803 (N_20803,N_18443,N_19008);
or U20804 (N_20804,N_19786,N_19594);
nor U20805 (N_20805,N_18403,N_18613);
nor U20806 (N_20806,N_18124,N_18484);
or U20807 (N_20807,N_17966,N_19790);
nor U20808 (N_20808,N_17983,N_19924);
and U20809 (N_20809,N_18077,N_19514);
and U20810 (N_20810,N_19273,N_19328);
and U20811 (N_20811,N_18602,N_19009);
nand U20812 (N_20812,N_19307,N_18209);
nand U20813 (N_20813,N_19973,N_18053);
nand U20814 (N_20814,N_18595,N_19808);
xor U20815 (N_20815,N_17820,N_19138);
nand U20816 (N_20816,N_19499,N_18112);
xnor U20817 (N_20817,N_17760,N_18752);
and U20818 (N_20818,N_19897,N_19027);
or U20819 (N_20819,N_19604,N_18895);
and U20820 (N_20820,N_18594,N_17911);
nor U20821 (N_20821,N_18741,N_19989);
and U20822 (N_20822,N_17844,N_18133);
xor U20823 (N_20823,N_17855,N_19881);
nor U20824 (N_20824,N_19417,N_18270);
nand U20825 (N_20825,N_18720,N_19177);
xor U20826 (N_20826,N_17514,N_18763);
nor U20827 (N_20827,N_17618,N_18563);
xor U20828 (N_20828,N_17642,N_18511);
or U20829 (N_20829,N_17750,N_18592);
and U20830 (N_20830,N_18813,N_19357);
nor U20831 (N_20831,N_19022,N_19873);
nor U20832 (N_20832,N_18197,N_19555);
nand U20833 (N_20833,N_18769,N_18830);
nand U20834 (N_20834,N_18586,N_17875);
nand U20835 (N_20835,N_17577,N_18781);
xnor U20836 (N_20836,N_19956,N_18357);
or U20837 (N_20837,N_19910,N_19416);
xnor U20838 (N_20838,N_18478,N_19234);
or U20839 (N_20839,N_19993,N_19479);
nand U20840 (N_20840,N_19463,N_19285);
nor U20841 (N_20841,N_18955,N_17693);
and U20842 (N_20842,N_19562,N_19963);
or U20843 (N_20843,N_19622,N_19547);
and U20844 (N_20844,N_19675,N_19553);
nand U20845 (N_20845,N_17564,N_18793);
or U20846 (N_20846,N_18034,N_18637);
xor U20847 (N_20847,N_18914,N_17962);
nand U20848 (N_20848,N_19907,N_18962);
nor U20849 (N_20849,N_18933,N_18279);
or U20850 (N_20850,N_19476,N_19205);
or U20851 (N_20851,N_18994,N_18298);
and U20852 (N_20852,N_19092,N_18192);
or U20853 (N_20853,N_19406,N_18806);
nor U20854 (N_20854,N_18977,N_18707);
nand U20855 (N_20855,N_18852,N_19259);
or U20856 (N_20856,N_18796,N_19216);
or U20857 (N_20857,N_17754,N_18271);
xor U20858 (N_20858,N_19470,N_17749);
nand U20859 (N_20859,N_19110,N_19399);
nor U20860 (N_20860,N_19778,N_18926);
nand U20861 (N_20861,N_18134,N_18330);
or U20862 (N_20862,N_19567,N_17503);
nand U20863 (N_20863,N_18400,N_19865);
nor U20864 (N_20864,N_19517,N_19004);
xnor U20865 (N_20865,N_19261,N_19936);
xnor U20866 (N_20866,N_19703,N_18236);
nor U20867 (N_20867,N_18560,N_18543);
and U20868 (N_20868,N_19798,N_19589);
nand U20869 (N_20869,N_18342,N_17997);
and U20870 (N_20870,N_17715,N_17914);
nor U20871 (N_20871,N_17588,N_19159);
nand U20872 (N_20872,N_19135,N_17803);
xor U20873 (N_20873,N_18418,N_18748);
nor U20874 (N_20874,N_19500,N_17717);
nand U20875 (N_20875,N_17545,N_19335);
nor U20876 (N_20876,N_19305,N_19568);
nor U20877 (N_20877,N_19174,N_19705);
nand U20878 (N_20878,N_18157,N_18088);
xor U20879 (N_20879,N_18315,N_18713);
or U20880 (N_20880,N_19725,N_18840);
and U20881 (N_20881,N_19625,N_18385);
nand U20882 (N_20882,N_18746,N_19724);
nor U20883 (N_20883,N_19142,N_18201);
and U20884 (N_20884,N_17925,N_17873);
or U20885 (N_20885,N_17806,N_18295);
nand U20886 (N_20886,N_18327,N_19212);
nand U20887 (N_20887,N_19085,N_17512);
or U20888 (N_20888,N_17552,N_19610);
nand U20889 (N_20889,N_18929,N_17832);
and U20890 (N_20890,N_17874,N_19935);
nand U20891 (N_20891,N_18889,N_18768);
or U20892 (N_20892,N_19563,N_18510);
nor U20893 (N_20893,N_17640,N_19580);
and U20894 (N_20894,N_19185,N_18703);
and U20895 (N_20895,N_18411,N_18782);
xor U20896 (N_20896,N_19995,N_19050);
or U20897 (N_20897,N_19015,N_18326);
and U20898 (N_20898,N_17970,N_18194);
and U20899 (N_20899,N_19364,N_19857);
xor U20900 (N_20900,N_18669,N_19368);
xnor U20901 (N_20901,N_17945,N_19084);
xnor U20902 (N_20902,N_18415,N_17825);
xor U20903 (N_20903,N_19069,N_19590);
or U20904 (N_20904,N_18362,N_19706);
nand U20905 (N_20905,N_19824,N_19465);
nand U20906 (N_20906,N_18642,N_18449);
and U20907 (N_20907,N_19380,N_18438);
nand U20908 (N_20908,N_19815,N_19267);
xor U20909 (N_20909,N_17797,N_17641);
and U20910 (N_20910,N_18476,N_19183);
and U20911 (N_20911,N_19391,N_18345);
or U20912 (N_20912,N_19372,N_18322);
or U20913 (N_20913,N_18035,N_18754);
nand U20914 (N_20914,N_17787,N_17689);
and U20915 (N_20915,N_18735,N_19359);
nor U20916 (N_20916,N_18898,N_18228);
xnor U20917 (N_20917,N_18423,N_18047);
and U20918 (N_20918,N_17860,N_19743);
xnor U20919 (N_20919,N_19885,N_17996);
nand U20920 (N_20920,N_18156,N_18646);
and U20921 (N_20921,N_19686,N_19295);
or U20922 (N_20922,N_19222,N_17558);
nor U20923 (N_20923,N_19531,N_17856);
or U20924 (N_20924,N_18948,N_19129);
nor U20925 (N_20925,N_19340,N_18507);
nand U20926 (N_20926,N_19795,N_17918);
nor U20927 (N_20927,N_18663,N_18060);
nand U20928 (N_20928,N_18892,N_17619);
nand U20929 (N_20929,N_18945,N_18612);
xnor U20930 (N_20930,N_18749,N_17730);
or U20931 (N_20931,N_19945,N_18974);
and U20932 (N_20932,N_17766,N_19983);
and U20933 (N_20933,N_17504,N_18382);
nor U20934 (N_20934,N_19039,N_18107);
nor U20935 (N_20935,N_18285,N_19025);
nor U20936 (N_20936,N_18421,N_18883);
or U20937 (N_20937,N_19330,N_19667);
and U20938 (N_20938,N_18278,N_19377);
and U20939 (N_20939,N_17903,N_18442);
and U20940 (N_20940,N_18108,N_18333);
or U20941 (N_20941,N_18764,N_17902);
or U20942 (N_20942,N_18715,N_19680);
xnor U20943 (N_20943,N_19753,N_18100);
and U20944 (N_20944,N_18875,N_18606);
nor U20945 (N_20945,N_18599,N_19960);
nand U20946 (N_20946,N_18408,N_18907);
nand U20947 (N_20947,N_18729,N_17964);
nand U20948 (N_20948,N_19982,N_17627);
nand U20949 (N_20949,N_18010,N_19921);
and U20950 (N_20950,N_19213,N_19608);
nand U20951 (N_20951,N_19337,N_18919);
nor U20952 (N_20952,N_17980,N_18988);
nor U20953 (N_20953,N_17698,N_18932);
or U20954 (N_20954,N_18351,N_17957);
nand U20955 (N_20955,N_19796,N_19994);
xor U20956 (N_20956,N_19215,N_19904);
or U20957 (N_20957,N_19903,N_17813);
or U20958 (N_20958,N_19324,N_19591);
and U20959 (N_20959,N_18857,N_19366);
or U20960 (N_20960,N_17959,N_18037);
nand U20961 (N_20961,N_17516,N_19466);
and U20962 (N_20962,N_17810,N_19152);
or U20963 (N_20963,N_17600,N_19246);
nand U20964 (N_20964,N_18927,N_19281);
xor U20965 (N_20965,N_18240,N_19642);
nand U20966 (N_20966,N_18824,N_19783);
or U20967 (N_20967,N_19615,N_19937);
or U20968 (N_20968,N_19551,N_18747);
or U20969 (N_20969,N_18995,N_18481);
xor U20970 (N_20970,N_19747,N_18011);
xnor U20971 (N_20971,N_18428,N_19320);
xor U20972 (N_20972,N_18537,N_19860);
or U20973 (N_20973,N_19294,N_19430);
and U20974 (N_20974,N_19852,N_19866);
nand U20975 (N_20975,N_19810,N_19480);
and U20976 (N_20976,N_18416,N_19445);
nor U20977 (N_20977,N_18255,N_18004);
nand U20978 (N_20978,N_18660,N_19353);
nand U20979 (N_20979,N_18474,N_17609);
or U20980 (N_20980,N_17620,N_19632);
nor U20981 (N_20981,N_18587,N_19721);
or U20982 (N_20982,N_19932,N_19737);
xor U20983 (N_20983,N_19859,N_18827);
xor U20984 (N_20984,N_19203,N_17706);
nor U20985 (N_20985,N_17986,N_19397);
xnor U20986 (N_20986,N_18375,N_19864);
xnor U20987 (N_20987,N_18779,N_19066);
nor U20988 (N_20988,N_18628,N_19014);
nand U20989 (N_20989,N_19588,N_19689);
or U20990 (N_20990,N_18963,N_17738);
and U20991 (N_20991,N_19558,N_19646);
nand U20992 (N_20992,N_18489,N_17861);
and U20993 (N_20993,N_19768,N_17823);
xnor U20994 (N_20994,N_18811,N_17563);
nand U20995 (N_20995,N_18798,N_18312);
and U20996 (N_20996,N_17837,N_19269);
nand U20997 (N_20997,N_17668,N_17793);
xnor U20998 (N_20998,N_18482,N_19948);
xor U20999 (N_20999,N_18908,N_19850);
or U21000 (N_21000,N_17799,N_18141);
or U21001 (N_21001,N_18260,N_18091);
nor U21002 (N_21002,N_19467,N_19316);
nand U21003 (N_21003,N_18969,N_18453);
and U21004 (N_21004,N_19781,N_18025);
nor U21005 (N_21005,N_17652,N_18616);
xnor U21006 (N_21006,N_18331,N_19200);
xnor U21007 (N_21007,N_19607,N_18993);
and U21008 (N_21008,N_19057,N_18575);
xnor U21009 (N_21009,N_18622,N_18885);
or U21010 (N_21010,N_18301,N_19557);
nor U21011 (N_21011,N_19762,N_18905);
nor U21012 (N_21012,N_19918,N_18377);
nor U21013 (N_21013,N_18495,N_18771);
nand U21014 (N_21014,N_18958,N_17614);
and U21015 (N_21015,N_19664,N_18583);
xnor U21016 (N_21016,N_19052,N_17587);
or U21017 (N_21017,N_18607,N_17667);
or U21018 (N_21018,N_19875,N_18547);
xor U21019 (N_21019,N_19439,N_18286);
nor U21020 (N_21020,N_17538,N_18401);
xor U21021 (N_21021,N_18203,N_18098);
nor U21022 (N_21022,N_18431,N_18925);
xnor U21023 (N_21023,N_18814,N_19707);
and U21024 (N_21024,N_18155,N_18205);
xnor U21025 (N_21025,N_19447,N_19820);
or U21026 (N_21026,N_19972,N_19277);
xnor U21027 (N_21027,N_19690,N_19542);
nor U21028 (N_21028,N_19260,N_18611);
nand U21029 (N_21029,N_18705,N_19804);
or U21030 (N_21030,N_19077,N_17784);
nand U21031 (N_21031,N_17646,N_18776);
nand U21032 (N_21032,N_18447,N_18632);
or U21033 (N_21033,N_18015,N_19464);
or U21034 (N_21034,N_19178,N_18101);
and U21035 (N_21035,N_18918,N_19496);
xor U21036 (N_21036,N_19031,N_19310);
nand U21037 (N_21037,N_18297,N_19487);
xnor U21038 (N_21038,N_19336,N_17669);
xnor U21039 (N_21039,N_19752,N_19929);
or U21040 (N_21040,N_19280,N_19985);
nand U21041 (N_21041,N_19474,N_17859);
nand U21042 (N_21042,N_18238,N_18036);
xor U21043 (N_21043,N_18787,N_18693);
or U21044 (N_21044,N_19426,N_18535);
nor U21045 (N_21045,N_19155,N_18459);
and U21046 (N_21046,N_18775,N_19777);
nand U21047 (N_21047,N_18387,N_18090);
or U21048 (N_21048,N_18841,N_18470);
nor U21049 (N_21049,N_18465,N_18880);
xnor U21050 (N_21050,N_19813,N_19586);
or U21051 (N_21051,N_18413,N_17644);
nand U21052 (N_21052,N_18258,N_17734);
xor U21053 (N_21053,N_18307,N_18142);
and U21054 (N_21054,N_17841,N_19136);
and U21055 (N_21055,N_19969,N_19565);
or U21056 (N_21056,N_17922,N_18656);
xor U21057 (N_21057,N_19763,N_17590);
xor U21058 (N_21058,N_19037,N_17539);
nor U21059 (N_21059,N_18797,N_19832);
or U21060 (N_21060,N_18799,N_17753);
xnor U21061 (N_21061,N_18542,N_19601);
and U21062 (N_21062,N_18336,N_17923);
nor U21063 (N_21063,N_19606,N_18614);
and U21064 (N_21064,N_19954,N_18790);
nor U21065 (N_21065,N_17621,N_18290);
nor U21066 (N_21066,N_19867,N_19481);
xor U21067 (N_21067,N_19585,N_18300);
and U21068 (N_21068,N_18215,N_18886);
nand U21069 (N_21069,N_18941,N_18078);
nor U21070 (N_21070,N_18486,N_18619);
or U21071 (N_21071,N_19510,N_18795);
and U21072 (N_21072,N_18540,N_18634);
or U21073 (N_21073,N_18624,N_18132);
xnor U21074 (N_21074,N_19386,N_17817);
nor U21075 (N_21075,N_17714,N_17901);
and U21076 (N_21076,N_17920,N_19966);
xnor U21077 (N_21077,N_19508,N_18343);
xnor U21078 (N_21078,N_19874,N_18692);
and U21079 (N_21079,N_18750,N_19438);
xnor U21080 (N_21080,N_18472,N_18127);
xor U21081 (N_21081,N_18849,N_17535);
nor U21082 (N_21082,N_19521,N_17842);
xor U21083 (N_21083,N_18111,N_17850);
xor U21084 (N_21084,N_17720,N_19403);
or U21085 (N_21085,N_18934,N_17505);
nor U21086 (N_21086,N_17878,N_19116);
or U21087 (N_21087,N_18687,N_18063);
nand U21088 (N_21088,N_19951,N_17907);
nor U21089 (N_21089,N_18722,N_18946);
nand U21090 (N_21090,N_19672,N_18959);
or U21091 (N_21091,N_18170,N_17637);
and U21092 (N_21092,N_17537,N_19272);
xor U21093 (N_21093,N_17649,N_19410);
nor U21094 (N_21094,N_19018,N_18601);
or U21095 (N_21095,N_19029,N_18366);
nand U21096 (N_21096,N_18968,N_17768);
nand U21097 (N_21097,N_17550,N_18700);
nor U21098 (N_21098,N_19700,N_18590);
nand U21099 (N_21099,N_19502,N_18027);
or U21100 (N_21100,N_17546,N_17795);
nand U21101 (N_21101,N_18454,N_17951);
nor U21102 (N_21102,N_17666,N_17967);
nand U21103 (N_21103,N_19959,N_18572);
or U21104 (N_21104,N_19694,N_18225);
xnor U21105 (N_21105,N_19911,N_19862);
and U21106 (N_21106,N_18661,N_18008);
xor U21107 (N_21107,N_19383,N_18876);
or U21108 (N_21108,N_18627,N_19418);
or U21109 (N_21109,N_18253,N_17840);
or U21110 (N_21110,N_17857,N_19113);
or U21111 (N_21111,N_19554,N_18159);
nand U21112 (N_21112,N_19146,N_17709);
nand U21113 (N_21113,N_18528,N_18066);
or U21114 (N_21114,N_17867,N_18545);
and U21115 (N_21115,N_18137,N_19251);
nor U21116 (N_21116,N_19550,N_19338);
or U21117 (N_21117,N_18140,N_18596);
and U21118 (N_21118,N_19575,N_18844);
nor U21119 (N_21119,N_18329,N_17876);
nor U21120 (N_21120,N_19891,N_17697);
and U21121 (N_21121,N_19158,N_18233);
nand U21122 (N_21122,N_18422,N_19384);
and U21123 (N_21123,N_18441,N_18229);
xor U21124 (N_21124,N_18324,N_17774);
nand U21125 (N_21125,N_17662,N_17804);
nand U21126 (N_21126,N_18897,N_18794);
and U21127 (N_21127,N_19927,N_18461);
nor U21128 (N_21128,N_17634,N_18014);
nor U21129 (N_21129,N_17759,N_17848);
xor U21130 (N_21130,N_18536,N_17958);
and U21131 (N_21131,N_18867,N_17821);
or U21132 (N_21132,N_19596,N_18556);
xnor U21133 (N_21133,N_17984,N_19202);
nor U21134 (N_21134,N_17858,N_19217);
or U21135 (N_21135,N_19638,N_19544);
or U21136 (N_21136,N_19162,N_18998);
xor U21137 (N_21137,N_18920,N_18402);
nor U21138 (N_21138,N_17522,N_18006);
or U21139 (N_21139,N_19473,N_17912);
xnor U21140 (N_21140,N_19809,N_19043);
xor U21141 (N_21141,N_17695,N_17725);
nand U21142 (N_21142,N_18029,N_17789);
xor U21143 (N_21143,N_19088,N_19028);
xnor U21144 (N_21144,N_18666,N_19223);
nor U21145 (N_21145,N_19332,N_19160);
or U21146 (N_21146,N_18420,N_17684);
and U21147 (N_21147,N_18701,N_19231);
xnor U21148 (N_21148,N_19872,N_19858);
xor U21149 (N_21149,N_18264,N_18483);
xor U21150 (N_21150,N_19245,N_18917);
and U21151 (N_21151,N_19197,N_19967);
nor U21152 (N_21152,N_18670,N_18086);
and U21153 (N_21153,N_18154,N_18847);
nor U21154 (N_21154,N_17593,N_19210);
and U21155 (N_21155,N_17783,N_18272);
xor U21156 (N_21156,N_18567,N_18001);
and U21157 (N_21157,N_17611,N_19093);
or U21158 (N_21158,N_19546,N_19387);
and U21159 (N_21159,N_18281,N_18237);
or U21160 (N_21160,N_19534,N_18756);
xor U21161 (N_21161,N_18650,N_17741);
xor U21162 (N_21162,N_19902,N_17946);
and U21163 (N_21163,N_19771,N_19803);
nand U21164 (N_21164,N_18397,N_17526);
xor U21165 (N_21165,N_17547,N_19811);
nor U21166 (N_21166,N_19802,N_19071);
or U21167 (N_21167,N_18389,N_17592);
xor U21168 (N_21168,N_19351,N_19346);
xor U21169 (N_21169,N_19206,N_18405);
or U21170 (N_21170,N_18158,N_18235);
nor U21171 (N_21171,N_17581,N_17928);
nand U21172 (N_21172,N_18374,N_19838);
nor U21173 (N_21173,N_19283,N_19732);
or U21174 (N_21174,N_19912,N_17751);
and U21175 (N_21175,N_19184,N_18598);
xnor U21176 (N_21176,N_19522,N_17692);
or U21177 (N_21177,N_17675,N_19693);
xor U21178 (N_21178,N_18186,N_18610);
xnor U21179 (N_21179,N_19327,N_17681);
and U21180 (N_21180,N_18514,N_19941);
or U21181 (N_21181,N_19456,N_17606);
and U21182 (N_21182,N_18003,N_19266);
nor U21183 (N_21183,N_18491,N_18639);
or U21184 (N_21184,N_19073,N_19094);
or U21185 (N_21185,N_17836,N_17676);
nand U21186 (N_21186,N_17794,N_19252);
nor U21187 (N_21187,N_19654,N_17589);
and U21188 (N_21188,N_19117,N_18114);
xor U21189 (N_21189,N_18515,N_19914);
and U21190 (N_21190,N_19095,N_19537);
nand U21191 (N_21191,N_19219,N_18275);
and U21192 (N_21192,N_19434,N_18899);
nand U21193 (N_21193,N_18942,N_18149);
or U21194 (N_21194,N_18395,N_19059);
nand U21195 (N_21195,N_19161,N_18122);
or U21196 (N_21196,N_19444,N_18604);
or U21197 (N_21197,N_18251,N_18527);
nor U21198 (N_21198,N_19720,N_19237);
xnor U21199 (N_21199,N_18410,N_19849);
xnor U21200 (N_21200,N_17736,N_19182);
xor U21201 (N_21201,N_19871,N_18552);
and U21202 (N_21202,N_17586,N_19484);
nand U21203 (N_21203,N_18517,N_19968);
nor U21204 (N_21204,N_19373,N_18859);
or U21205 (N_21205,N_19154,N_19909);
xnor U21206 (N_21206,N_18220,N_19698);
nor U21207 (N_21207,N_19942,N_17879);
nand U21208 (N_21208,N_18353,N_18176);
and U21209 (N_21209,N_19965,N_17924);
nand U21210 (N_21210,N_19894,N_17562);
nand U21211 (N_21211,N_17746,N_18224);
nor U21212 (N_21212,N_17708,N_18099);
xnor U21213 (N_21213,N_18202,N_18288);
and U21214 (N_21214,N_19538,N_19455);
nand U21215 (N_21215,N_17896,N_19287);
xor U21216 (N_21216,N_17733,N_19701);
xor U21217 (N_21217,N_17949,N_19817);
and U21218 (N_21218,N_19101,N_19851);
and U21219 (N_21219,N_19730,N_18965);
and U21220 (N_21220,N_19067,N_19291);
nand U21221 (N_21221,N_19493,N_19381);
or U21222 (N_21222,N_18721,N_18649);
or U21223 (N_21223,N_17829,N_19501);
nor U21224 (N_21224,N_17899,N_18367);
nor U21225 (N_21225,N_19235,N_18755);
and U21226 (N_21226,N_19276,N_17553);
xnor U21227 (N_21227,N_17916,N_18040);
xor U21228 (N_21228,N_18172,N_18879);
or U21229 (N_21229,N_19868,N_18997);
or U21230 (N_21230,N_18440,N_19112);
or U21231 (N_21231,N_18792,N_18113);
nor U21232 (N_21232,N_19428,N_18325);
xnor U21233 (N_21233,N_18083,N_17566);
xnor U21234 (N_21234,N_19497,N_17893);
nor U21235 (N_21235,N_19189,N_18058);
xor U21236 (N_21236,N_18455,N_19414);
nand U21237 (N_21237,N_18909,N_18302);
nor U21238 (N_21238,N_17659,N_19301);
xor U21239 (N_21239,N_18904,N_19420);
or U21240 (N_21240,N_18647,N_17777);
and U21241 (N_21241,N_18115,N_18135);
nand U21242 (N_21242,N_19369,N_17728);
and U21243 (N_21243,N_19143,N_17890);
or U21244 (N_21244,N_18446,N_18626);
nand U21245 (N_21245,N_18872,N_18548);
xnor U21246 (N_21246,N_17556,N_19145);
xor U21247 (N_21247,N_19623,N_19611);
and U21248 (N_21248,N_17686,N_18017);
nor U21249 (N_21249,N_19893,N_19421);
and U21250 (N_21250,N_18217,N_19135);
xnor U21251 (N_21251,N_19822,N_18419);
xnor U21252 (N_21252,N_19023,N_19944);
and U21253 (N_21253,N_17555,N_17771);
nand U21254 (N_21254,N_19517,N_17945);
or U21255 (N_21255,N_19288,N_18481);
or U21256 (N_21256,N_17777,N_18541);
or U21257 (N_21257,N_19338,N_19961);
nand U21258 (N_21258,N_18384,N_18832);
nand U21259 (N_21259,N_17923,N_18698);
or U21260 (N_21260,N_18606,N_18518);
and U21261 (N_21261,N_17990,N_19925);
nor U21262 (N_21262,N_17517,N_19156);
or U21263 (N_21263,N_19824,N_18300);
xor U21264 (N_21264,N_19193,N_17737);
nand U21265 (N_21265,N_19203,N_17570);
nand U21266 (N_21266,N_19411,N_17578);
nand U21267 (N_21267,N_18156,N_18349);
xor U21268 (N_21268,N_17859,N_17628);
nor U21269 (N_21269,N_18088,N_17851);
or U21270 (N_21270,N_19765,N_19184);
xnor U21271 (N_21271,N_19390,N_17767);
and U21272 (N_21272,N_19497,N_18273);
or U21273 (N_21273,N_19247,N_18768);
nand U21274 (N_21274,N_19358,N_19580);
and U21275 (N_21275,N_17894,N_19747);
nand U21276 (N_21276,N_18782,N_19942);
and U21277 (N_21277,N_18670,N_19923);
or U21278 (N_21278,N_19709,N_19435);
nor U21279 (N_21279,N_19767,N_19616);
xnor U21280 (N_21280,N_17735,N_17678);
or U21281 (N_21281,N_19766,N_18516);
nand U21282 (N_21282,N_18146,N_18449);
and U21283 (N_21283,N_19489,N_19681);
xor U21284 (N_21284,N_17679,N_17729);
and U21285 (N_21285,N_18926,N_19273);
or U21286 (N_21286,N_17813,N_19498);
xor U21287 (N_21287,N_17793,N_18517);
nand U21288 (N_21288,N_18963,N_19224);
nand U21289 (N_21289,N_19848,N_17612);
nand U21290 (N_21290,N_18169,N_17729);
nor U21291 (N_21291,N_19218,N_17567);
nor U21292 (N_21292,N_17625,N_17710);
nand U21293 (N_21293,N_17635,N_19361);
nor U21294 (N_21294,N_18556,N_18879);
nor U21295 (N_21295,N_19235,N_18868);
nor U21296 (N_21296,N_19881,N_19190);
or U21297 (N_21297,N_19592,N_19699);
nand U21298 (N_21298,N_19733,N_17716);
and U21299 (N_21299,N_17538,N_18926);
xor U21300 (N_21300,N_19932,N_17687);
nor U21301 (N_21301,N_19944,N_17684);
or U21302 (N_21302,N_18310,N_19081);
or U21303 (N_21303,N_18518,N_19052);
nor U21304 (N_21304,N_19424,N_19405);
nand U21305 (N_21305,N_18236,N_17565);
xor U21306 (N_21306,N_19076,N_18417);
nor U21307 (N_21307,N_17877,N_19298);
nor U21308 (N_21308,N_19688,N_18682);
and U21309 (N_21309,N_19276,N_19244);
nor U21310 (N_21310,N_18459,N_19372);
nand U21311 (N_21311,N_19569,N_17714);
or U21312 (N_21312,N_19748,N_17589);
nor U21313 (N_21313,N_18283,N_18879);
and U21314 (N_21314,N_18417,N_18027);
nor U21315 (N_21315,N_18997,N_18592);
nand U21316 (N_21316,N_18013,N_18847);
or U21317 (N_21317,N_18266,N_19337);
xor U21318 (N_21318,N_19392,N_19728);
xnor U21319 (N_21319,N_19799,N_19566);
nand U21320 (N_21320,N_19163,N_18023);
nor U21321 (N_21321,N_18770,N_19947);
nand U21322 (N_21322,N_19333,N_17638);
and U21323 (N_21323,N_18503,N_17961);
nor U21324 (N_21324,N_19442,N_19714);
nand U21325 (N_21325,N_18710,N_19740);
and U21326 (N_21326,N_19209,N_19638);
or U21327 (N_21327,N_19349,N_18591);
nor U21328 (N_21328,N_18666,N_17795);
or U21329 (N_21329,N_18524,N_19433);
or U21330 (N_21330,N_19660,N_18240);
xor U21331 (N_21331,N_18197,N_19692);
xor U21332 (N_21332,N_18077,N_18200);
nor U21333 (N_21333,N_18167,N_18169);
xnor U21334 (N_21334,N_18408,N_18836);
nand U21335 (N_21335,N_19827,N_18749);
nor U21336 (N_21336,N_18135,N_19006);
nand U21337 (N_21337,N_19827,N_17501);
and U21338 (N_21338,N_19221,N_18201);
and U21339 (N_21339,N_18441,N_19543);
and U21340 (N_21340,N_19836,N_18822);
or U21341 (N_21341,N_19331,N_18928);
nor U21342 (N_21342,N_17861,N_19627);
nand U21343 (N_21343,N_19904,N_18420);
xor U21344 (N_21344,N_18398,N_18760);
or U21345 (N_21345,N_18242,N_18677);
nor U21346 (N_21346,N_19216,N_19070);
nor U21347 (N_21347,N_19697,N_19107);
xor U21348 (N_21348,N_18588,N_19912);
or U21349 (N_21349,N_18023,N_19584);
xnor U21350 (N_21350,N_18865,N_17947);
and U21351 (N_21351,N_19460,N_17525);
xor U21352 (N_21352,N_19433,N_19673);
and U21353 (N_21353,N_18649,N_17995);
and U21354 (N_21354,N_17661,N_18257);
xor U21355 (N_21355,N_18815,N_18641);
nand U21356 (N_21356,N_19833,N_19411);
nor U21357 (N_21357,N_17650,N_18218);
nand U21358 (N_21358,N_18539,N_18795);
or U21359 (N_21359,N_19339,N_19954);
xnor U21360 (N_21360,N_19711,N_19742);
or U21361 (N_21361,N_17834,N_19074);
or U21362 (N_21362,N_19042,N_19253);
or U21363 (N_21363,N_18732,N_17801);
and U21364 (N_21364,N_19579,N_19350);
xor U21365 (N_21365,N_17668,N_18533);
or U21366 (N_21366,N_19189,N_18042);
and U21367 (N_21367,N_18301,N_19165);
xnor U21368 (N_21368,N_18314,N_19783);
xnor U21369 (N_21369,N_18573,N_18487);
nor U21370 (N_21370,N_17747,N_18680);
nor U21371 (N_21371,N_19735,N_18361);
xor U21372 (N_21372,N_18009,N_19172);
xor U21373 (N_21373,N_19573,N_19219);
or U21374 (N_21374,N_19819,N_19346);
nand U21375 (N_21375,N_18854,N_17873);
xor U21376 (N_21376,N_19772,N_18115);
and U21377 (N_21377,N_19991,N_17524);
xor U21378 (N_21378,N_17940,N_18730);
nor U21379 (N_21379,N_18840,N_19298);
nand U21380 (N_21380,N_17899,N_19938);
or U21381 (N_21381,N_19627,N_18234);
and U21382 (N_21382,N_19966,N_18417);
nor U21383 (N_21383,N_17524,N_19235);
or U21384 (N_21384,N_17859,N_19247);
and U21385 (N_21385,N_18940,N_17737);
nand U21386 (N_21386,N_17704,N_18184);
or U21387 (N_21387,N_18100,N_19610);
xnor U21388 (N_21388,N_19291,N_17899);
and U21389 (N_21389,N_19454,N_19500);
nor U21390 (N_21390,N_18774,N_17763);
nand U21391 (N_21391,N_17891,N_19602);
xnor U21392 (N_21392,N_19984,N_19894);
nor U21393 (N_21393,N_19658,N_19834);
xnor U21394 (N_21394,N_19809,N_18578);
nand U21395 (N_21395,N_19039,N_18731);
or U21396 (N_21396,N_19323,N_19512);
nor U21397 (N_21397,N_19517,N_19845);
nand U21398 (N_21398,N_19326,N_18056);
xnor U21399 (N_21399,N_19285,N_18700);
nor U21400 (N_21400,N_17824,N_18041);
or U21401 (N_21401,N_19065,N_19498);
and U21402 (N_21402,N_19331,N_19020);
and U21403 (N_21403,N_19009,N_18400);
or U21404 (N_21404,N_19700,N_19004);
nand U21405 (N_21405,N_18380,N_18171);
and U21406 (N_21406,N_19613,N_19694);
or U21407 (N_21407,N_19676,N_18396);
xor U21408 (N_21408,N_19226,N_18257);
and U21409 (N_21409,N_19827,N_18318);
nand U21410 (N_21410,N_18451,N_19166);
nand U21411 (N_21411,N_17965,N_19807);
and U21412 (N_21412,N_19091,N_17968);
and U21413 (N_21413,N_18124,N_17902);
and U21414 (N_21414,N_18582,N_18899);
xor U21415 (N_21415,N_18281,N_17894);
nand U21416 (N_21416,N_17616,N_17837);
nand U21417 (N_21417,N_17891,N_18840);
xnor U21418 (N_21418,N_19852,N_18508);
and U21419 (N_21419,N_18296,N_18830);
and U21420 (N_21420,N_17515,N_18504);
and U21421 (N_21421,N_19396,N_17628);
nor U21422 (N_21422,N_17895,N_17780);
and U21423 (N_21423,N_18914,N_18230);
xnor U21424 (N_21424,N_17500,N_18298);
or U21425 (N_21425,N_19015,N_19504);
xor U21426 (N_21426,N_19169,N_17718);
xor U21427 (N_21427,N_18353,N_18117);
xnor U21428 (N_21428,N_17500,N_17565);
xnor U21429 (N_21429,N_18473,N_17848);
or U21430 (N_21430,N_18496,N_19700);
nand U21431 (N_21431,N_18082,N_18381);
xnor U21432 (N_21432,N_17910,N_17582);
nor U21433 (N_21433,N_19196,N_19229);
xnor U21434 (N_21434,N_19880,N_18670);
and U21435 (N_21435,N_18651,N_18635);
nor U21436 (N_21436,N_18507,N_18593);
and U21437 (N_21437,N_18552,N_19287);
xnor U21438 (N_21438,N_17853,N_17672);
nand U21439 (N_21439,N_19343,N_18405);
and U21440 (N_21440,N_18406,N_17700);
and U21441 (N_21441,N_19668,N_19226);
nand U21442 (N_21442,N_17968,N_18921);
or U21443 (N_21443,N_17502,N_17849);
or U21444 (N_21444,N_19575,N_18788);
nand U21445 (N_21445,N_19721,N_18925);
xnor U21446 (N_21446,N_19170,N_17641);
nor U21447 (N_21447,N_18116,N_18332);
xnor U21448 (N_21448,N_17671,N_19583);
nor U21449 (N_21449,N_18719,N_19295);
xnor U21450 (N_21450,N_19774,N_19193);
nor U21451 (N_21451,N_19506,N_19364);
or U21452 (N_21452,N_18820,N_18029);
nand U21453 (N_21453,N_19675,N_18492);
nand U21454 (N_21454,N_19460,N_19774);
xor U21455 (N_21455,N_17972,N_18806);
xnor U21456 (N_21456,N_18300,N_17891);
and U21457 (N_21457,N_19956,N_19807);
nor U21458 (N_21458,N_18983,N_18970);
nand U21459 (N_21459,N_19094,N_18516);
and U21460 (N_21460,N_17774,N_19257);
nor U21461 (N_21461,N_19740,N_19689);
nor U21462 (N_21462,N_19889,N_19962);
xor U21463 (N_21463,N_17815,N_18883);
and U21464 (N_21464,N_18402,N_17734);
or U21465 (N_21465,N_19991,N_18498);
or U21466 (N_21466,N_18941,N_19151);
and U21467 (N_21467,N_19624,N_19018);
xnor U21468 (N_21468,N_17609,N_19946);
nor U21469 (N_21469,N_19127,N_19470);
xnor U21470 (N_21470,N_19129,N_18001);
nand U21471 (N_21471,N_19727,N_18596);
xor U21472 (N_21472,N_19070,N_19202);
and U21473 (N_21473,N_19900,N_18851);
nor U21474 (N_21474,N_18350,N_19115);
nand U21475 (N_21475,N_18552,N_18362);
or U21476 (N_21476,N_18613,N_19205);
xnor U21477 (N_21477,N_19455,N_17678);
nand U21478 (N_21478,N_19761,N_19821);
and U21479 (N_21479,N_19306,N_17721);
and U21480 (N_21480,N_19952,N_17678);
xor U21481 (N_21481,N_19407,N_19683);
nor U21482 (N_21482,N_19132,N_18616);
nor U21483 (N_21483,N_19084,N_19475);
xor U21484 (N_21484,N_17762,N_17899);
xor U21485 (N_21485,N_17793,N_18937);
or U21486 (N_21486,N_18827,N_19538);
nor U21487 (N_21487,N_18174,N_19174);
and U21488 (N_21488,N_18450,N_18614);
nor U21489 (N_21489,N_18463,N_18434);
or U21490 (N_21490,N_18142,N_18451);
or U21491 (N_21491,N_17665,N_18104);
nor U21492 (N_21492,N_18990,N_19506);
and U21493 (N_21493,N_18035,N_18250);
and U21494 (N_21494,N_19607,N_19139);
and U21495 (N_21495,N_19548,N_19353);
nor U21496 (N_21496,N_19441,N_19018);
nor U21497 (N_21497,N_19771,N_19541);
nor U21498 (N_21498,N_19262,N_17690);
or U21499 (N_21499,N_19401,N_18282);
and U21500 (N_21500,N_19851,N_18363);
or U21501 (N_21501,N_17533,N_17682);
xor U21502 (N_21502,N_19963,N_17609);
xor U21503 (N_21503,N_19375,N_19736);
nor U21504 (N_21504,N_17858,N_19546);
or U21505 (N_21505,N_19105,N_18265);
or U21506 (N_21506,N_19322,N_18632);
or U21507 (N_21507,N_17932,N_18719);
or U21508 (N_21508,N_18784,N_17818);
or U21509 (N_21509,N_18530,N_18868);
or U21510 (N_21510,N_18052,N_17888);
nor U21511 (N_21511,N_19050,N_18433);
and U21512 (N_21512,N_19685,N_18435);
or U21513 (N_21513,N_19589,N_18448);
and U21514 (N_21514,N_18398,N_18353);
or U21515 (N_21515,N_19895,N_18740);
nand U21516 (N_21516,N_19855,N_19419);
and U21517 (N_21517,N_17792,N_19910);
or U21518 (N_21518,N_19743,N_19664);
and U21519 (N_21519,N_19016,N_18679);
nor U21520 (N_21520,N_18996,N_19221);
or U21521 (N_21521,N_19147,N_19194);
nand U21522 (N_21522,N_18963,N_19208);
or U21523 (N_21523,N_17737,N_19184);
nor U21524 (N_21524,N_18151,N_18080);
xnor U21525 (N_21525,N_19050,N_18010);
nor U21526 (N_21526,N_18930,N_18544);
or U21527 (N_21527,N_19595,N_19054);
nor U21528 (N_21528,N_19766,N_17542);
xnor U21529 (N_21529,N_18223,N_19568);
or U21530 (N_21530,N_19072,N_18389);
and U21531 (N_21531,N_18997,N_18764);
or U21532 (N_21532,N_18276,N_18172);
and U21533 (N_21533,N_19272,N_19707);
and U21534 (N_21534,N_19775,N_18184);
nand U21535 (N_21535,N_18359,N_18238);
xnor U21536 (N_21536,N_17501,N_18243);
nor U21537 (N_21537,N_18069,N_18408);
nor U21538 (N_21538,N_18593,N_18077);
xor U21539 (N_21539,N_18582,N_19982);
nor U21540 (N_21540,N_18414,N_19063);
nand U21541 (N_21541,N_18957,N_18677);
or U21542 (N_21542,N_18155,N_17923);
nand U21543 (N_21543,N_18254,N_17595);
nor U21544 (N_21544,N_17593,N_17888);
xnor U21545 (N_21545,N_19814,N_19403);
or U21546 (N_21546,N_18211,N_18137);
xnor U21547 (N_21547,N_18198,N_19904);
and U21548 (N_21548,N_18759,N_19297);
or U21549 (N_21549,N_19015,N_19556);
nand U21550 (N_21550,N_18871,N_18903);
nand U21551 (N_21551,N_19710,N_19087);
xor U21552 (N_21552,N_17845,N_18543);
and U21553 (N_21553,N_19786,N_19752);
nor U21554 (N_21554,N_18542,N_18359);
and U21555 (N_21555,N_19599,N_18353);
xor U21556 (N_21556,N_19979,N_18508);
nand U21557 (N_21557,N_18803,N_19916);
and U21558 (N_21558,N_18920,N_18616);
xor U21559 (N_21559,N_18271,N_19485);
or U21560 (N_21560,N_18624,N_19174);
xor U21561 (N_21561,N_18908,N_18630);
or U21562 (N_21562,N_17830,N_17676);
nand U21563 (N_21563,N_18730,N_19097);
nand U21564 (N_21564,N_19396,N_18636);
and U21565 (N_21565,N_18633,N_18160);
nand U21566 (N_21566,N_18214,N_18864);
xor U21567 (N_21567,N_17633,N_19015);
nand U21568 (N_21568,N_18358,N_19357);
nor U21569 (N_21569,N_19278,N_19394);
or U21570 (N_21570,N_18836,N_18381);
nor U21571 (N_21571,N_19536,N_19467);
and U21572 (N_21572,N_18972,N_18409);
xnor U21573 (N_21573,N_19878,N_18212);
nor U21574 (N_21574,N_19777,N_17650);
or U21575 (N_21575,N_19956,N_19689);
nor U21576 (N_21576,N_18478,N_19365);
nand U21577 (N_21577,N_18002,N_18833);
nand U21578 (N_21578,N_17993,N_18407);
or U21579 (N_21579,N_19765,N_18064);
nor U21580 (N_21580,N_17558,N_18061);
and U21581 (N_21581,N_19771,N_18637);
and U21582 (N_21582,N_18250,N_17630);
or U21583 (N_21583,N_19249,N_18088);
and U21584 (N_21584,N_19791,N_19085);
and U21585 (N_21585,N_17830,N_18100);
nand U21586 (N_21586,N_19088,N_18219);
xnor U21587 (N_21587,N_19923,N_18090);
or U21588 (N_21588,N_17699,N_18409);
xor U21589 (N_21589,N_19403,N_19130);
nand U21590 (N_21590,N_17505,N_19873);
and U21591 (N_21591,N_19553,N_18847);
nand U21592 (N_21592,N_18697,N_17765);
nor U21593 (N_21593,N_18271,N_18009);
nor U21594 (N_21594,N_17726,N_19990);
nand U21595 (N_21595,N_19902,N_19945);
and U21596 (N_21596,N_19350,N_19224);
and U21597 (N_21597,N_19902,N_17853);
and U21598 (N_21598,N_19004,N_19492);
or U21599 (N_21599,N_19489,N_17518);
nand U21600 (N_21600,N_17766,N_18188);
nor U21601 (N_21601,N_18276,N_18082);
nor U21602 (N_21602,N_19812,N_19882);
or U21603 (N_21603,N_19510,N_17789);
nor U21604 (N_21604,N_18287,N_18154);
xnor U21605 (N_21605,N_19715,N_18191);
or U21606 (N_21606,N_17852,N_19524);
nor U21607 (N_21607,N_18853,N_18892);
and U21608 (N_21608,N_17603,N_19767);
nor U21609 (N_21609,N_18892,N_19404);
or U21610 (N_21610,N_18686,N_18335);
nor U21611 (N_21611,N_19628,N_19909);
xor U21612 (N_21612,N_18653,N_19663);
or U21613 (N_21613,N_19970,N_18258);
nor U21614 (N_21614,N_19702,N_17539);
or U21615 (N_21615,N_19694,N_17715);
and U21616 (N_21616,N_19446,N_18706);
and U21617 (N_21617,N_19743,N_19921);
nor U21618 (N_21618,N_17577,N_19398);
xor U21619 (N_21619,N_18345,N_17850);
nand U21620 (N_21620,N_19663,N_19782);
nor U21621 (N_21621,N_17971,N_19579);
nand U21622 (N_21622,N_17559,N_18471);
nor U21623 (N_21623,N_18463,N_18220);
or U21624 (N_21624,N_19817,N_19938);
nor U21625 (N_21625,N_17592,N_19204);
and U21626 (N_21626,N_19898,N_19765);
xnor U21627 (N_21627,N_19760,N_17716);
nor U21628 (N_21628,N_18237,N_19763);
and U21629 (N_21629,N_17768,N_18019);
xnor U21630 (N_21630,N_18030,N_19447);
nor U21631 (N_21631,N_18353,N_17659);
nand U21632 (N_21632,N_19239,N_17644);
and U21633 (N_21633,N_18850,N_18997);
nor U21634 (N_21634,N_19286,N_18505);
or U21635 (N_21635,N_19293,N_19613);
nand U21636 (N_21636,N_18578,N_18872);
nor U21637 (N_21637,N_19076,N_18243);
or U21638 (N_21638,N_18647,N_18551);
xnor U21639 (N_21639,N_18969,N_18361);
or U21640 (N_21640,N_18873,N_17504);
or U21641 (N_21641,N_18500,N_19449);
or U21642 (N_21642,N_19975,N_17878);
and U21643 (N_21643,N_19593,N_19204);
or U21644 (N_21644,N_17932,N_19835);
and U21645 (N_21645,N_18359,N_18342);
xnor U21646 (N_21646,N_19631,N_18810);
and U21647 (N_21647,N_19972,N_19279);
xnor U21648 (N_21648,N_17720,N_17815);
xnor U21649 (N_21649,N_17946,N_17572);
nor U21650 (N_21650,N_17931,N_19500);
nor U21651 (N_21651,N_17517,N_18795);
nand U21652 (N_21652,N_17756,N_18562);
xnor U21653 (N_21653,N_18322,N_18137);
nor U21654 (N_21654,N_18107,N_18846);
nand U21655 (N_21655,N_19312,N_19113);
xor U21656 (N_21656,N_17775,N_19343);
xor U21657 (N_21657,N_19401,N_18356);
xnor U21658 (N_21658,N_18794,N_18672);
or U21659 (N_21659,N_18033,N_18358);
and U21660 (N_21660,N_19727,N_18070);
xor U21661 (N_21661,N_18707,N_19691);
xnor U21662 (N_21662,N_18487,N_18101);
and U21663 (N_21663,N_18656,N_18993);
nor U21664 (N_21664,N_17753,N_19899);
nand U21665 (N_21665,N_18255,N_18247);
or U21666 (N_21666,N_18985,N_19196);
and U21667 (N_21667,N_18493,N_17964);
xor U21668 (N_21668,N_17989,N_18619);
nor U21669 (N_21669,N_19897,N_17944);
or U21670 (N_21670,N_18755,N_19107);
xnor U21671 (N_21671,N_18243,N_19616);
nor U21672 (N_21672,N_19813,N_17882);
and U21673 (N_21673,N_18495,N_19677);
xnor U21674 (N_21674,N_19023,N_19853);
nand U21675 (N_21675,N_18345,N_19619);
xor U21676 (N_21676,N_18349,N_18992);
xor U21677 (N_21677,N_18748,N_17830);
xor U21678 (N_21678,N_18321,N_18300);
and U21679 (N_21679,N_18850,N_18273);
xnor U21680 (N_21680,N_19958,N_17848);
or U21681 (N_21681,N_18834,N_18317);
nor U21682 (N_21682,N_19668,N_18209);
nand U21683 (N_21683,N_19209,N_17759);
nor U21684 (N_21684,N_18751,N_18400);
nand U21685 (N_21685,N_19283,N_19230);
and U21686 (N_21686,N_19768,N_19933);
nand U21687 (N_21687,N_18283,N_17620);
or U21688 (N_21688,N_19241,N_19308);
nor U21689 (N_21689,N_18856,N_19878);
or U21690 (N_21690,N_17606,N_18769);
nand U21691 (N_21691,N_19037,N_19091);
or U21692 (N_21692,N_19005,N_17789);
nand U21693 (N_21693,N_19326,N_18281);
xnor U21694 (N_21694,N_19443,N_18938);
nand U21695 (N_21695,N_18167,N_19550);
nor U21696 (N_21696,N_18421,N_19845);
or U21697 (N_21697,N_18137,N_18476);
nor U21698 (N_21698,N_19305,N_17644);
nand U21699 (N_21699,N_17861,N_19435);
xor U21700 (N_21700,N_17566,N_18739);
nor U21701 (N_21701,N_18668,N_19377);
nand U21702 (N_21702,N_19903,N_19263);
or U21703 (N_21703,N_19329,N_18610);
or U21704 (N_21704,N_19452,N_18444);
or U21705 (N_21705,N_18185,N_17756);
or U21706 (N_21706,N_18570,N_17627);
or U21707 (N_21707,N_17990,N_17587);
nand U21708 (N_21708,N_17788,N_19763);
nor U21709 (N_21709,N_19976,N_18235);
or U21710 (N_21710,N_19386,N_18164);
xor U21711 (N_21711,N_17780,N_19732);
xnor U21712 (N_21712,N_18798,N_17516);
nand U21713 (N_21713,N_17632,N_18543);
or U21714 (N_21714,N_18189,N_17998);
and U21715 (N_21715,N_17851,N_17512);
nand U21716 (N_21716,N_18765,N_18326);
or U21717 (N_21717,N_18214,N_18806);
nor U21718 (N_21718,N_17505,N_17736);
nand U21719 (N_21719,N_17771,N_18349);
nand U21720 (N_21720,N_18008,N_18870);
and U21721 (N_21721,N_18614,N_19272);
and U21722 (N_21722,N_19958,N_19073);
and U21723 (N_21723,N_19407,N_17534);
nand U21724 (N_21724,N_19234,N_18293);
nor U21725 (N_21725,N_19776,N_18345);
nand U21726 (N_21726,N_19820,N_17872);
and U21727 (N_21727,N_18789,N_17998);
or U21728 (N_21728,N_19833,N_19326);
or U21729 (N_21729,N_18078,N_18996);
nor U21730 (N_21730,N_18923,N_18496);
and U21731 (N_21731,N_18565,N_18310);
xnor U21732 (N_21732,N_18019,N_18075);
and U21733 (N_21733,N_18464,N_19692);
nand U21734 (N_21734,N_17627,N_17660);
xor U21735 (N_21735,N_18084,N_18758);
nor U21736 (N_21736,N_17951,N_17613);
or U21737 (N_21737,N_18309,N_19232);
xnor U21738 (N_21738,N_18151,N_17784);
or U21739 (N_21739,N_18123,N_18823);
or U21740 (N_21740,N_17532,N_17581);
xnor U21741 (N_21741,N_18268,N_19082);
and U21742 (N_21742,N_19258,N_17743);
nand U21743 (N_21743,N_17565,N_18098);
nor U21744 (N_21744,N_19343,N_18905);
or U21745 (N_21745,N_18366,N_17650);
and U21746 (N_21746,N_19825,N_17667);
nor U21747 (N_21747,N_17570,N_18926);
and U21748 (N_21748,N_19432,N_18606);
or U21749 (N_21749,N_19453,N_18892);
or U21750 (N_21750,N_19664,N_18993);
nor U21751 (N_21751,N_18008,N_18749);
and U21752 (N_21752,N_19270,N_19536);
or U21753 (N_21753,N_19918,N_18058);
and U21754 (N_21754,N_18040,N_18193);
nor U21755 (N_21755,N_18416,N_18948);
and U21756 (N_21756,N_18150,N_18322);
or U21757 (N_21757,N_19720,N_18118);
nor U21758 (N_21758,N_18805,N_18432);
nand U21759 (N_21759,N_19977,N_17831);
xnor U21760 (N_21760,N_18554,N_17680);
nor U21761 (N_21761,N_18311,N_19736);
nand U21762 (N_21762,N_18407,N_17986);
nand U21763 (N_21763,N_18220,N_18405);
and U21764 (N_21764,N_19519,N_19830);
nand U21765 (N_21765,N_18172,N_19494);
and U21766 (N_21766,N_19478,N_17827);
or U21767 (N_21767,N_17602,N_18347);
nor U21768 (N_21768,N_18549,N_18889);
nor U21769 (N_21769,N_19898,N_18826);
nor U21770 (N_21770,N_18103,N_19645);
and U21771 (N_21771,N_19769,N_19167);
and U21772 (N_21772,N_19054,N_17973);
nor U21773 (N_21773,N_19462,N_19026);
nand U21774 (N_21774,N_18448,N_19045);
nand U21775 (N_21775,N_19776,N_18595);
and U21776 (N_21776,N_18802,N_19535);
xor U21777 (N_21777,N_19269,N_18817);
xor U21778 (N_21778,N_19547,N_19854);
or U21779 (N_21779,N_17545,N_17526);
and U21780 (N_21780,N_19352,N_18158);
nand U21781 (N_21781,N_18435,N_19857);
and U21782 (N_21782,N_18563,N_17707);
xnor U21783 (N_21783,N_17614,N_19765);
and U21784 (N_21784,N_18152,N_18391);
nand U21785 (N_21785,N_17850,N_18564);
and U21786 (N_21786,N_18664,N_17724);
or U21787 (N_21787,N_19600,N_18738);
nand U21788 (N_21788,N_18352,N_19567);
nor U21789 (N_21789,N_17921,N_18534);
nor U21790 (N_21790,N_18726,N_18567);
or U21791 (N_21791,N_17771,N_18514);
nand U21792 (N_21792,N_18782,N_18553);
nor U21793 (N_21793,N_18305,N_18805);
nand U21794 (N_21794,N_17684,N_17905);
nor U21795 (N_21795,N_18115,N_18452);
nor U21796 (N_21796,N_19154,N_19563);
nor U21797 (N_21797,N_19442,N_17730);
or U21798 (N_21798,N_18010,N_18100);
nor U21799 (N_21799,N_19266,N_17614);
nand U21800 (N_21800,N_18752,N_18228);
or U21801 (N_21801,N_18886,N_18326);
xnor U21802 (N_21802,N_18230,N_18246);
or U21803 (N_21803,N_17598,N_18101);
nor U21804 (N_21804,N_19381,N_18308);
and U21805 (N_21805,N_18335,N_19139);
nand U21806 (N_21806,N_19965,N_19067);
or U21807 (N_21807,N_19281,N_17731);
or U21808 (N_21808,N_19508,N_17781);
xor U21809 (N_21809,N_18264,N_19897);
and U21810 (N_21810,N_19688,N_19425);
nor U21811 (N_21811,N_17787,N_19940);
xnor U21812 (N_21812,N_18316,N_19026);
nor U21813 (N_21813,N_17678,N_18663);
nand U21814 (N_21814,N_18838,N_18345);
nand U21815 (N_21815,N_17669,N_19214);
nor U21816 (N_21816,N_18409,N_18158);
or U21817 (N_21817,N_17874,N_17564);
nor U21818 (N_21818,N_19725,N_18019);
nor U21819 (N_21819,N_19343,N_18573);
nor U21820 (N_21820,N_18491,N_19707);
nand U21821 (N_21821,N_19788,N_17799);
and U21822 (N_21822,N_18675,N_19046);
nor U21823 (N_21823,N_18833,N_19477);
or U21824 (N_21824,N_19653,N_18300);
and U21825 (N_21825,N_18366,N_19555);
or U21826 (N_21826,N_19382,N_19741);
xnor U21827 (N_21827,N_18640,N_17833);
nor U21828 (N_21828,N_19278,N_17900);
and U21829 (N_21829,N_18712,N_18338);
or U21830 (N_21830,N_17779,N_19901);
and U21831 (N_21831,N_18493,N_18978);
nor U21832 (N_21832,N_19596,N_17946);
nor U21833 (N_21833,N_18717,N_18660);
nor U21834 (N_21834,N_17931,N_19535);
xor U21835 (N_21835,N_18751,N_18036);
and U21836 (N_21836,N_18144,N_19273);
and U21837 (N_21837,N_18490,N_18668);
nor U21838 (N_21838,N_19721,N_18991);
or U21839 (N_21839,N_18210,N_18826);
xor U21840 (N_21840,N_19543,N_18265);
nand U21841 (N_21841,N_18144,N_18183);
or U21842 (N_21842,N_19174,N_18952);
nor U21843 (N_21843,N_18929,N_17669);
nor U21844 (N_21844,N_18886,N_19272);
xnor U21845 (N_21845,N_17907,N_19653);
or U21846 (N_21846,N_18489,N_19583);
nor U21847 (N_21847,N_18863,N_19683);
and U21848 (N_21848,N_19803,N_18762);
nand U21849 (N_21849,N_19068,N_18750);
and U21850 (N_21850,N_18104,N_19928);
nor U21851 (N_21851,N_19730,N_19238);
and U21852 (N_21852,N_19672,N_18399);
or U21853 (N_21853,N_19413,N_18779);
nand U21854 (N_21854,N_18996,N_18812);
or U21855 (N_21855,N_18551,N_19313);
nor U21856 (N_21856,N_19594,N_17661);
nor U21857 (N_21857,N_19190,N_18123);
xnor U21858 (N_21858,N_19665,N_17536);
nor U21859 (N_21859,N_18471,N_18264);
or U21860 (N_21860,N_19486,N_17867);
xnor U21861 (N_21861,N_18859,N_18705);
nor U21862 (N_21862,N_19785,N_19657);
xor U21863 (N_21863,N_19585,N_19117);
xor U21864 (N_21864,N_18267,N_19012);
xnor U21865 (N_21865,N_18073,N_18793);
nand U21866 (N_21866,N_18425,N_17682);
nor U21867 (N_21867,N_19881,N_18848);
and U21868 (N_21868,N_17703,N_17981);
xnor U21869 (N_21869,N_19313,N_19377);
or U21870 (N_21870,N_19208,N_19407);
nand U21871 (N_21871,N_19990,N_19403);
nand U21872 (N_21872,N_19605,N_19777);
nand U21873 (N_21873,N_17941,N_17728);
nand U21874 (N_21874,N_19733,N_19927);
nand U21875 (N_21875,N_18426,N_18536);
xnor U21876 (N_21876,N_18940,N_18744);
and U21877 (N_21877,N_19129,N_18125);
xnor U21878 (N_21878,N_19604,N_18421);
nor U21879 (N_21879,N_18852,N_17599);
or U21880 (N_21880,N_19465,N_18582);
nand U21881 (N_21881,N_17664,N_19858);
nor U21882 (N_21882,N_19484,N_17929);
or U21883 (N_21883,N_18492,N_18420);
xnor U21884 (N_21884,N_19628,N_17698);
nand U21885 (N_21885,N_17511,N_19020);
nand U21886 (N_21886,N_18584,N_19960);
nand U21887 (N_21887,N_18065,N_19219);
and U21888 (N_21888,N_18048,N_18188);
xnor U21889 (N_21889,N_17933,N_19975);
nor U21890 (N_21890,N_19584,N_19082);
and U21891 (N_21891,N_18840,N_19543);
nor U21892 (N_21892,N_18540,N_17963);
xnor U21893 (N_21893,N_19685,N_19666);
nor U21894 (N_21894,N_17630,N_18099);
and U21895 (N_21895,N_17647,N_19313);
nor U21896 (N_21896,N_17978,N_19587);
nand U21897 (N_21897,N_17858,N_18520);
xor U21898 (N_21898,N_19723,N_19613);
nor U21899 (N_21899,N_17782,N_19995);
and U21900 (N_21900,N_19312,N_18329);
xnor U21901 (N_21901,N_18369,N_18398);
and U21902 (N_21902,N_18973,N_19199);
and U21903 (N_21903,N_18166,N_17678);
and U21904 (N_21904,N_18969,N_19974);
nor U21905 (N_21905,N_18040,N_19008);
nor U21906 (N_21906,N_17689,N_19447);
nor U21907 (N_21907,N_19365,N_17564);
or U21908 (N_21908,N_19386,N_17979);
nor U21909 (N_21909,N_17904,N_19371);
and U21910 (N_21910,N_18297,N_18288);
or U21911 (N_21911,N_18139,N_19745);
or U21912 (N_21912,N_19042,N_18041);
and U21913 (N_21913,N_18384,N_18224);
nand U21914 (N_21914,N_18630,N_19670);
or U21915 (N_21915,N_19438,N_18340);
xor U21916 (N_21916,N_17914,N_19898);
nand U21917 (N_21917,N_19632,N_17876);
nor U21918 (N_21918,N_17569,N_17539);
and U21919 (N_21919,N_19991,N_18920);
nand U21920 (N_21920,N_19827,N_19148);
xnor U21921 (N_21921,N_18356,N_19649);
nand U21922 (N_21922,N_18982,N_18090);
nand U21923 (N_21923,N_18405,N_19811);
nand U21924 (N_21924,N_19742,N_19452);
xor U21925 (N_21925,N_18357,N_18514);
xor U21926 (N_21926,N_17728,N_19258);
and U21927 (N_21927,N_18944,N_19718);
or U21928 (N_21928,N_17664,N_17622);
xor U21929 (N_21929,N_18827,N_18975);
nand U21930 (N_21930,N_19017,N_18754);
nor U21931 (N_21931,N_18489,N_17977);
or U21932 (N_21932,N_19896,N_18112);
nor U21933 (N_21933,N_18118,N_19722);
xor U21934 (N_21934,N_18476,N_19797);
xnor U21935 (N_21935,N_19946,N_18628);
and U21936 (N_21936,N_18655,N_18764);
nand U21937 (N_21937,N_19093,N_19089);
nand U21938 (N_21938,N_18627,N_18706);
xnor U21939 (N_21939,N_19323,N_18578);
or U21940 (N_21940,N_17794,N_18643);
or U21941 (N_21941,N_19508,N_17762);
nand U21942 (N_21942,N_17708,N_17518);
xor U21943 (N_21943,N_18058,N_18459);
and U21944 (N_21944,N_19485,N_19129);
nor U21945 (N_21945,N_19466,N_17617);
xnor U21946 (N_21946,N_19830,N_17771);
and U21947 (N_21947,N_19261,N_18931);
and U21948 (N_21948,N_17520,N_18095);
xnor U21949 (N_21949,N_17792,N_19170);
nor U21950 (N_21950,N_18410,N_19491);
or U21951 (N_21951,N_17948,N_17803);
xnor U21952 (N_21952,N_19284,N_18615);
nand U21953 (N_21953,N_18557,N_18240);
and U21954 (N_21954,N_19606,N_19412);
xnor U21955 (N_21955,N_17794,N_19241);
nor U21956 (N_21956,N_19614,N_18719);
nand U21957 (N_21957,N_18963,N_18671);
and U21958 (N_21958,N_17821,N_18477);
and U21959 (N_21959,N_17670,N_17756);
nand U21960 (N_21960,N_19663,N_18964);
and U21961 (N_21961,N_17586,N_19975);
nor U21962 (N_21962,N_19454,N_17552);
xor U21963 (N_21963,N_18907,N_17971);
nand U21964 (N_21964,N_17618,N_17705);
xor U21965 (N_21965,N_19980,N_19399);
xor U21966 (N_21966,N_18281,N_18769);
nand U21967 (N_21967,N_19409,N_18590);
xnor U21968 (N_21968,N_18664,N_19510);
xor U21969 (N_21969,N_19099,N_19479);
or U21970 (N_21970,N_17521,N_19623);
nand U21971 (N_21971,N_18280,N_18168);
nor U21972 (N_21972,N_19703,N_18591);
and U21973 (N_21973,N_18709,N_19242);
xnor U21974 (N_21974,N_18522,N_19223);
nand U21975 (N_21975,N_19586,N_18782);
nor U21976 (N_21976,N_17695,N_17598);
xnor U21977 (N_21977,N_19642,N_18881);
and U21978 (N_21978,N_17776,N_17705);
nand U21979 (N_21979,N_18152,N_17796);
xor U21980 (N_21980,N_19945,N_18367);
or U21981 (N_21981,N_18258,N_19112);
or U21982 (N_21982,N_18918,N_18540);
nor U21983 (N_21983,N_18548,N_18066);
and U21984 (N_21984,N_17899,N_19425);
and U21985 (N_21985,N_17963,N_19559);
or U21986 (N_21986,N_19643,N_19337);
nor U21987 (N_21987,N_18941,N_19869);
nor U21988 (N_21988,N_18348,N_19908);
nand U21989 (N_21989,N_19636,N_17952);
nor U21990 (N_21990,N_19898,N_19011);
nor U21991 (N_21991,N_17536,N_19471);
and U21992 (N_21992,N_18174,N_18547);
nor U21993 (N_21993,N_18078,N_18111);
nor U21994 (N_21994,N_19230,N_19714);
xnor U21995 (N_21995,N_18233,N_17761);
nand U21996 (N_21996,N_19420,N_18958);
and U21997 (N_21997,N_18013,N_17665);
nand U21998 (N_21998,N_17739,N_18769);
or U21999 (N_21999,N_19871,N_17939);
and U22000 (N_22000,N_17554,N_17636);
and U22001 (N_22001,N_19375,N_18577);
xor U22002 (N_22002,N_17862,N_18501);
or U22003 (N_22003,N_19587,N_17549);
and U22004 (N_22004,N_17742,N_19105);
or U22005 (N_22005,N_18609,N_18505);
nor U22006 (N_22006,N_19615,N_17666);
and U22007 (N_22007,N_18075,N_18321);
or U22008 (N_22008,N_17977,N_17779);
or U22009 (N_22009,N_19069,N_17527);
nor U22010 (N_22010,N_18907,N_19794);
and U22011 (N_22011,N_18125,N_17687);
or U22012 (N_22012,N_19471,N_18785);
or U22013 (N_22013,N_18573,N_18627);
nand U22014 (N_22014,N_19204,N_18293);
or U22015 (N_22015,N_18817,N_18670);
or U22016 (N_22016,N_19561,N_19122);
or U22017 (N_22017,N_19784,N_17651);
or U22018 (N_22018,N_19058,N_17654);
and U22019 (N_22019,N_18840,N_18676);
and U22020 (N_22020,N_18026,N_19090);
and U22021 (N_22021,N_18570,N_18314);
and U22022 (N_22022,N_18200,N_19174);
or U22023 (N_22023,N_18966,N_18206);
nor U22024 (N_22024,N_18182,N_18013);
or U22025 (N_22025,N_18234,N_17558);
xnor U22026 (N_22026,N_18210,N_17905);
or U22027 (N_22027,N_17974,N_19461);
nand U22028 (N_22028,N_17668,N_18137);
nor U22029 (N_22029,N_18202,N_19435);
xor U22030 (N_22030,N_19831,N_17903);
xnor U22031 (N_22031,N_19873,N_18674);
or U22032 (N_22032,N_18251,N_18037);
or U22033 (N_22033,N_17535,N_19532);
xor U22034 (N_22034,N_18766,N_19451);
and U22035 (N_22035,N_19660,N_17764);
or U22036 (N_22036,N_19939,N_19765);
nand U22037 (N_22037,N_17709,N_18216);
or U22038 (N_22038,N_19505,N_19032);
xnor U22039 (N_22039,N_18358,N_18055);
or U22040 (N_22040,N_17888,N_18931);
xnor U22041 (N_22041,N_19990,N_18036);
xnor U22042 (N_22042,N_19433,N_18905);
nand U22043 (N_22043,N_19620,N_18414);
and U22044 (N_22044,N_18196,N_17953);
or U22045 (N_22045,N_18651,N_18766);
xor U22046 (N_22046,N_18084,N_18011);
nor U22047 (N_22047,N_19643,N_19659);
or U22048 (N_22048,N_19961,N_19385);
nor U22049 (N_22049,N_19753,N_17840);
xnor U22050 (N_22050,N_18234,N_19995);
and U22051 (N_22051,N_18061,N_18362);
xor U22052 (N_22052,N_17968,N_18370);
nand U22053 (N_22053,N_19995,N_19748);
nor U22054 (N_22054,N_19539,N_19505);
xnor U22055 (N_22055,N_18916,N_17541);
nand U22056 (N_22056,N_19997,N_19222);
and U22057 (N_22057,N_19534,N_17897);
nand U22058 (N_22058,N_19147,N_17596);
nand U22059 (N_22059,N_18704,N_18906);
xnor U22060 (N_22060,N_19110,N_19393);
nand U22061 (N_22061,N_19186,N_18518);
or U22062 (N_22062,N_17682,N_18194);
nor U22063 (N_22063,N_18905,N_19810);
or U22064 (N_22064,N_19554,N_17822);
or U22065 (N_22065,N_19001,N_18391);
or U22066 (N_22066,N_18549,N_19647);
xor U22067 (N_22067,N_18973,N_17709);
nand U22068 (N_22068,N_18139,N_17516);
xor U22069 (N_22069,N_19180,N_17855);
nor U22070 (N_22070,N_17575,N_18519);
nor U22071 (N_22071,N_17825,N_18331);
nand U22072 (N_22072,N_19213,N_19579);
xor U22073 (N_22073,N_18956,N_18046);
or U22074 (N_22074,N_18216,N_19303);
and U22075 (N_22075,N_18514,N_19920);
or U22076 (N_22076,N_19590,N_19847);
xnor U22077 (N_22077,N_17813,N_18895);
nand U22078 (N_22078,N_19037,N_18879);
and U22079 (N_22079,N_19148,N_19690);
xor U22080 (N_22080,N_19827,N_18087);
or U22081 (N_22081,N_17655,N_18346);
nor U22082 (N_22082,N_18380,N_19286);
xor U22083 (N_22083,N_19021,N_19860);
nor U22084 (N_22084,N_18332,N_19498);
nand U22085 (N_22085,N_19305,N_17777);
or U22086 (N_22086,N_19386,N_18939);
nand U22087 (N_22087,N_17783,N_18030);
nor U22088 (N_22088,N_19247,N_18012);
nand U22089 (N_22089,N_18019,N_18144);
nand U22090 (N_22090,N_19586,N_19687);
or U22091 (N_22091,N_17977,N_19854);
and U22092 (N_22092,N_18073,N_18554);
xnor U22093 (N_22093,N_19282,N_18198);
xor U22094 (N_22094,N_19196,N_19879);
nand U22095 (N_22095,N_19587,N_18522);
nor U22096 (N_22096,N_19192,N_18835);
or U22097 (N_22097,N_19244,N_19231);
and U22098 (N_22098,N_18283,N_19810);
and U22099 (N_22099,N_17774,N_19597);
or U22100 (N_22100,N_18658,N_19335);
nor U22101 (N_22101,N_19146,N_18184);
or U22102 (N_22102,N_19277,N_19502);
nor U22103 (N_22103,N_19979,N_19419);
nand U22104 (N_22104,N_19610,N_19146);
nor U22105 (N_22105,N_18214,N_17907);
or U22106 (N_22106,N_18527,N_19887);
and U22107 (N_22107,N_18525,N_17927);
nor U22108 (N_22108,N_18525,N_17683);
nand U22109 (N_22109,N_17991,N_18855);
and U22110 (N_22110,N_19459,N_17598);
nor U22111 (N_22111,N_17979,N_18510);
nor U22112 (N_22112,N_17896,N_19452);
xnor U22113 (N_22113,N_19067,N_17608);
and U22114 (N_22114,N_18549,N_18189);
or U22115 (N_22115,N_19654,N_17647);
or U22116 (N_22116,N_19540,N_18753);
and U22117 (N_22117,N_18027,N_19798);
nand U22118 (N_22118,N_19824,N_18556);
and U22119 (N_22119,N_18025,N_19541);
nor U22120 (N_22120,N_18528,N_17906);
xor U22121 (N_22121,N_18274,N_18960);
or U22122 (N_22122,N_18616,N_18552);
xor U22123 (N_22123,N_18220,N_18795);
xnor U22124 (N_22124,N_19870,N_18551);
nand U22125 (N_22125,N_19827,N_19446);
xor U22126 (N_22126,N_18587,N_18006);
nand U22127 (N_22127,N_19941,N_17735);
nor U22128 (N_22128,N_18476,N_19382);
nor U22129 (N_22129,N_19759,N_18004);
nand U22130 (N_22130,N_18681,N_18990);
nor U22131 (N_22131,N_19923,N_18593);
or U22132 (N_22132,N_17887,N_18636);
nor U22133 (N_22133,N_18106,N_19152);
or U22134 (N_22134,N_18685,N_18976);
nor U22135 (N_22135,N_17737,N_19575);
and U22136 (N_22136,N_19241,N_18758);
nor U22137 (N_22137,N_18470,N_18974);
nor U22138 (N_22138,N_19282,N_18170);
nand U22139 (N_22139,N_19378,N_18145);
or U22140 (N_22140,N_17621,N_18155);
nand U22141 (N_22141,N_17515,N_19015);
nor U22142 (N_22142,N_17999,N_18452);
and U22143 (N_22143,N_18538,N_18268);
nand U22144 (N_22144,N_19218,N_17654);
nor U22145 (N_22145,N_18008,N_17710);
or U22146 (N_22146,N_19346,N_17743);
and U22147 (N_22147,N_17596,N_19321);
xor U22148 (N_22148,N_19519,N_19404);
nor U22149 (N_22149,N_18301,N_19228);
nand U22150 (N_22150,N_18672,N_19443);
and U22151 (N_22151,N_18063,N_19929);
nand U22152 (N_22152,N_17785,N_19620);
or U22153 (N_22153,N_17810,N_18090);
or U22154 (N_22154,N_17681,N_18506);
and U22155 (N_22155,N_17509,N_18649);
or U22156 (N_22156,N_17632,N_19836);
nand U22157 (N_22157,N_18761,N_19668);
xnor U22158 (N_22158,N_18610,N_19969);
or U22159 (N_22159,N_18870,N_19445);
and U22160 (N_22160,N_17962,N_18445);
and U22161 (N_22161,N_18949,N_17925);
and U22162 (N_22162,N_18920,N_18195);
xor U22163 (N_22163,N_18119,N_18142);
xnor U22164 (N_22164,N_18532,N_19748);
nor U22165 (N_22165,N_19335,N_19665);
nor U22166 (N_22166,N_18260,N_18905);
xor U22167 (N_22167,N_18517,N_18928);
nand U22168 (N_22168,N_19132,N_19448);
nand U22169 (N_22169,N_19273,N_18733);
and U22170 (N_22170,N_18262,N_17937);
or U22171 (N_22171,N_19587,N_18663);
and U22172 (N_22172,N_19074,N_18189);
nand U22173 (N_22173,N_19738,N_17962);
xnor U22174 (N_22174,N_17680,N_18803);
and U22175 (N_22175,N_18383,N_18227);
nor U22176 (N_22176,N_19429,N_17576);
nor U22177 (N_22177,N_17854,N_17696);
or U22178 (N_22178,N_19565,N_19526);
nor U22179 (N_22179,N_19202,N_18987);
nor U22180 (N_22180,N_18526,N_19597);
nor U22181 (N_22181,N_19201,N_19228);
and U22182 (N_22182,N_17951,N_18799);
and U22183 (N_22183,N_17897,N_18218);
and U22184 (N_22184,N_19362,N_17699);
nand U22185 (N_22185,N_18198,N_19213);
nor U22186 (N_22186,N_19864,N_19243);
nand U22187 (N_22187,N_19573,N_18038);
nor U22188 (N_22188,N_18385,N_17831);
and U22189 (N_22189,N_18116,N_17671);
nand U22190 (N_22190,N_19729,N_19938);
and U22191 (N_22191,N_18856,N_19024);
xnor U22192 (N_22192,N_19746,N_17898);
and U22193 (N_22193,N_18944,N_18562);
nand U22194 (N_22194,N_18292,N_18917);
and U22195 (N_22195,N_17592,N_19698);
nor U22196 (N_22196,N_18592,N_18986);
nor U22197 (N_22197,N_17847,N_19563);
nor U22198 (N_22198,N_18635,N_19771);
nand U22199 (N_22199,N_19682,N_18736);
nand U22200 (N_22200,N_17648,N_19127);
and U22201 (N_22201,N_18789,N_19280);
nor U22202 (N_22202,N_19878,N_18867);
nand U22203 (N_22203,N_19847,N_19624);
nand U22204 (N_22204,N_18299,N_18593);
or U22205 (N_22205,N_18131,N_18099);
nor U22206 (N_22206,N_18311,N_19989);
nand U22207 (N_22207,N_18495,N_19525);
nor U22208 (N_22208,N_19760,N_19377);
nor U22209 (N_22209,N_17758,N_19964);
nand U22210 (N_22210,N_18550,N_17803);
and U22211 (N_22211,N_18115,N_18131);
nand U22212 (N_22212,N_19035,N_19121);
nand U22213 (N_22213,N_19588,N_18913);
xor U22214 (N_22214,N_18125,N_17760);
or U22215 (N_22215,N_19564,N_18839);
and U22216 (N_22216,N_19670,N_17554);
nor U22217 (N_22217,N_18096,N_19220);
and U22218 (N_22218,N_17600,N_18497);
nor U22219 (N_22219,N_18629,N_18470);
and U22220 (N_22220,N_17734,N_18292);
xor U22221 (N_22221,N_19271,N_17554);
nor U22222 (N_22222,N_19535,N_17602);
nand U22223 (N_22223,N_18827,N_18764);
nand U22224 (N_22224,N_19689,N_19957);
and U22225 (N_22225,N_18694,N_19758);
and U22226 (N_22226,N_19481,N_17616);
and U22227 (N_22227,N_18455,N_18958);
nand U22228 (N_22228,N_18047,N_19623);
and U22229 (N_22229,N_18835,N_18002);
nor U22230 (N_22230,N_18673,N_19398);
xor U22231 (N_22231,N_19082,N_17915);
and U22232 (N_22232,N_18939,N_18433);
and U22233 (N_22233,N_18585,N_19631);
or U22234 (N_22234,N_19374,N_18140);
or U22235 (N_22235,N_17981,N_19867);
nand U22236 (N_22236,N_19819,N_19381);
xor U22237 (N_22237,N_18087,N_17720);
or U22238 (N_22238,N_18910,N_19673);
nor U22239 (N_22239,N_17872,N_17563);
nor U22240 (N_22240,N_18203,N_19435);
or U22241 (N_22241,N_19943,N_18594);
xor U22242 (N_22242,N_19684,N_19482);
nand U22243 (N_22243,N_18208,N_19521);
or U22244 (N_22244,N_18037,N_19331);
or U22245 (N_22245,N_19614,N_18090);
nand U22246 (N_22246,N_17537,N_17831);
xnor U22247 (N_22247,N_18115,N_19824);
nand U22248 (N_22248,N_17519,N_18419);
and U22249 (N_22249,N_18544,N_19805);
and U22250 (N_22250,N_18166,N_18325);
or U22251 (N_22251,N_18290,N_19437);
xnor U22252 (N_22252,N_19418,N_18769);
and U22253 (N_22253,N_17643,N_18061);
and U22254 (N_22254,N_19356,N_19046);
xor U22255 (N_22255,N_19188,N_18008);
nor U22256 (N_22256,N_18559,N_19011);
and U22257 (N_22257,N_18190,N_18104);
nor U22258 (N_22258,N_18182,N_18752);
or U22259 (N_22259,N_19946,N_18773);
nor U22260 (N_22260,N_18000,N_18407);
nand U22261 (N_22261,N_18285,N_19707);
nand U22262 (N_22262,N_19903,N_17502);
nand U22263 (N_22263,N_18788,N_17842);
or U22264 (N_22264,N_19538,N_17673);
xnor U22265 (N_22265,N_18898,N_18400);
nor U22266 (N_22266,N_19036,N_19283);
nand U22267 (N_22267,N_18350,N_19330);
nand U22268 (N_22268,N_17927,N_19913);
xor U22269 (N_22269,N_18329,N_19635);
and U22270 (N_22270,N_17997,N_17620);
and U22271 (N_22271,N_19435,N_18890);
or U22272 (N_22272,N_18223,N_18627);
nor U22273 (N_22273,N_18237,N_18677);
xor U22274 (N_22274,N_19684,N_17732);
or U22275 (N_22275,N_18013,N_19644);
and U22276 (N_22276,N_18375,N_18506);
or U22277 (N_22277,N_18633,N_17920);
nand U22278 (N_22278,N_19653,N_19039);
nor U22279 (N_22279,N_19473,N_18367);
nor U22280 (N_22280,N_17645,N_18057);
nor U22281 (N_22281,N_19771,N_18286);
or U22282 (N_22282,N_19707,N_18308);
or U22283 (N_22283,N_19491,N_19326);
and U22284 (N_22284,N_19727,N_17647);
nor U22285 (N_22285,N_19810,N_17700);
nand U22286 (N_22286,N_19594,N_17719);
nor U22287 (N_22287,N_19491,N_17826);
nand U22288 (N_22288,N_18674,N_19452);
nor U22289 (N_22289,N_19155,N_17702);
and U22290 (N_22290,N_18107,N_18970);
and U22291 (N_22291,N_18270,N_19955);
or U22292 (N_22292,N_19832,N_18781);
xor U22293 (N_22293,N_18279,N_18438);
xor U22294 (N_22294,N_17936,N_18986);
and U22295 (N_22295,N_19480,N_18429);
or U22296 (N_22296,N_17767,N_17993);
or U22297 (N_22297,N_18219,N_17604);
or U22298 (N_22298,N_19282,N_19026);
and U22299 (N_22299,N_17917,N_18088);
xnor U22300 (N_22300,N_18925,N_17853);
and U22301 (N_22301,N_19107,N_18892);
nand U22302 (N_22302,N_19108,N_18307);
nand U22303 (N_22303,N_18612,N_19748);
nand U22304 (N_22304,N_19828,N_19038);
or U22305 (N_22305,N_18230,N_17674);
nand U22306 (N_22306,N_17684,N_19643);
xnor U22307 (N_22307,N_17610,N_17889);
nor U22308 (N_22308,N_18020,N_19104);
xnor U22309 (N_22309,N_19684,N_19333);
and U22310 (N_22310,N_19044,N_18733);
and U22311 (N_22311,N_18220,N_18523);
nor U22312 (N_22312,N_19708,N_18646);
nor U22313 (N_22313,N_17837,N_18910);
or U22314 (N_22314,N_18474,N_17584);
and U22315 (N_22315,N_19058,N_18881);
nand U22316 (N_22316,N_19971,N_18828);
nand U22317 (N_22317,N_17989,N_18087);
nand U22318 (N_22318,N_18085,N_19368);
nor U22319 (N_22319,N_19556,N_17860);
or U22320 (N_22320,N_18582,N_18171);
or U22321 (N_22321,N_18730,N_19194);
or U22322 (N_22322,N_19885,N_18796);
xor U22323 (N_22323,N_17507,N_17815);
xnor U22324 (N_22324,N_19420,N_18889);
or U22325 (N_22325,N_19471,N_18286);
nor U22326 (N_22326,N_17766,N_19075);
or U22327 (N_22327,N_18167,N_17697);
nand U22328 (N_22328,N_18927,N_18656);
nand U22329 (N_22329,N_17594,N_19949);
nand U22330 (N_22330,N_18609,N_17514);
or U22331 (N_22331,N_19417,N_19977);
nand U22332 (N_22332,N_17786,N_18850);
and U22333 (N_22333,N_19288,N_17818);
nor U22334 (N_22334,N_18175,N_18563);
nand U22335 (N_22335,N_17783,N_19837);
and U22336 (N_22336,N_19364,N_19965);
and U22337 (N_22337,N_19002,N_17554);
nand U22338 (N_22338,N_19023,N_17803);
or U22339 (N_22339,N_17556,N_19815);
nor U22340 (N_22340,N_17749,N_18376);
nand U22341 (N_22341,N_19634,N_19274);
nor U22342 (N_22342,N_17758,N_18373);
xnor U22343 (N_22343,N_18309,N_18264);
nand U22344 (N_22344,N_19605,N_18670);
nor U22345 (N_22345,N_18190,N_18012);
nor U22346 (N_22346,N_19765,N_19716);
and U22347 (N_22347,N_18821,N_18286);
nand U22348 (N_22348,N_17708,N_19398);
or U22349 (N_22349,N_18553,N_19355);
or U22350 (N_22350,N_19940,N_19893);
or U22351 (N_22351,N_19883,N_17991);
nor U22352 (N_22352,N_18286,N_18773);
nand U22353 (N_22353,N_17505,N_18617);
nand U22354 (N_22354,N_18585,N_18537);
xor U22355 (N_22355,N_18813,N_18108);
nand U22356 (N_22356,N_18131,N_19855);
xor U22357 (N_22357,N_19795,N_18155);
nand U22358 (N_22358,N_17942,N_18169);
and U22359 (N_22359,N_18204,N_17891);
xnor U22360 (N_22360,N_18940,N_18355);
nand U22361 (N_22361,N_18161,N_19575);
nand U22362 (N_22362,N_17948,N_18228);
nand U22363 (N_22363,N_18319,N_17509);
or U22364 (N_22364,N_18309,N_19305);
nor U22365 (N_22365,N_18283,N_17931);
or U22366 (N_22366,N_19134,N_19125);
nand U22367 (N_22367,N_18668,N_18408);
xor U22368 (N_22368,N_19381,N_19273);
nand U22369 (N_22369,N_17882,N_19847);
nor U22370 (N_22370,N_18732,N_19220);
nor U22371 (N_22371,N_19107,N_17812);
xor U22372 (N_22372,N_19232,N_19658);
and U22373 (N_22373,N_19412,N_18060);
xor U22374 (N_22374,N_18885,N_18853);
nor U22375 (N_22375,N_19013,N_19469);
and U22376 (N_22376,N_19763,N_18527);
or U22377 (N_22377,N_19665,N_17882);
or U22378 (N_22378,N_19506,N_17897);
nor U22379 (N_22379,N_18482,N_18036);
nor U22380 (N_22380,N_19762,N_19098);
nand U22381 (N_22381,N_17888,N_19127);
xnor U22382 (N_22382,N_17839,N_17544);
xnor U22383 (N_22383,N_17583,N_19312);
nand U22384 (N_22384,N_18229,N_18004);
nor U22385 (N_22385,N_18710,N_17922);
xor U22386 (N_22386,N_18361,N_18853);
xor U22387 (N_22387,N_18141,N_17574);
and U22388 (N_22388,N_18109,N_19019);
nand U22389 (N_22389,N_19964,N_18577);
nor U22390 (N_22390,N_19913,N_17876);
nor U22391 (N_22391,N_17819,N_17871);
xor U22392 (N_22392,N_19175,N_17563);
nor U22393 (N_22393,N_19896,N_18966);
and U22394 (N_22394,N_17543,N_18487);
nor U22395 (N_22395,N_17682,N_18869);
nor U22396 (N_22396,N_19134,N_17541);
and U22397 (N_22397,N_18069,N_18978);
or U22398 (N_22398,N_17663,N_18374);
or U22399 (N_22399,N_19241,N_17682);
xnor U22400 (N_22400,N_18614,N_18615);
or U22401 (N_22401,N_19977,N_19772);
and U22402 (N_22402,N_18847,N_19867);
or U22403 (N_22403,N_17721,N_18172);
nor U22404 (N_22404,N_19431,N_17796);
nor U22405 (N_22405,N_18349,N_18575);
and U22406 (N_22406,N_19955,N_17635);
nor U22407 (N_22407,N_18588,N_18064);
nand U22408 (N_22408,N_19851,N_19321);
and U22409 (N_22409,N_17890,N_19672);
nand U22410 (N_22410,N_18100,N_18266);
nand U22411 (N_22411,N_18560,N_19228);
nand U22412 (N_22412,N_18491,N_18662);
and U22413 (N_22413,N_19029,N_18802);
nand U22414 (N_22414,N_19224,N_19701);
or U22415 (N_22415,N_17901,N_18721);
or U22416 (N_22416,N_19544,N_19692);
nor U22417 (N_22417,N_17997,N_17576);
xor U22418 (N_22418,N_19195,N_19714);
and U22419 (N_22419,N_19891,N_17811);
and U22420 (N_22420,N_17650,N_19792);
and U22421 (N_22421,N_17854,N_19013);
xor U22422 (N_22422,N_17893,N_18582);
nand U22423 (N_22423,N_18163,N_18440);
or U22424 (N_22424,N_18469,N_19187);
xor U22425 (N_22425,N_19197,N_19340);
xnor U22426 (N_22426,N_19369,N_19722);
nor U22427 (N_22427,N_17990,N_18473);
nand U22428 (N_22428,N_19173,N_17804);
xnor U22429 (N_22429,N_18921,N_18151);
or U22430 (N_22430,N_18447,N_17783);
or U22431 (N_22431,N_18894,N_19909);
nand U22432 (N_22432,N_19872,N_17902);
xnor U22433 (N_22433,N_19579,N_18450);
nand U22434 (N_22434,N_19590,N_18188);
nor U22435 (N_22435,N_18354,N_19314);
nor U22436 (N_22436,N_19653,N_17504);
or U22437 (N_22437,N_18635,N_18388);
or U22438 (N_22438,N_18710,N_19072);
and U22439 (N_22439,N_17889,N_19711);
xnor U22440 (N_22440,N_19544,N_17623);
nor U22441 (N_22441,N_18002,N_19332);
or U22442 (N_22442,N_17858,N_19218);
xnor U22443 (N_22443,N_17971,N_19136);
nor U22444 (N_22444,N_17869,N_18594);
or U22445 (N_22445,N_17509,N_19394);
xnor U22446 (N_22446,N_19587,N_18584);
xor U22447 (N_22447,N_18865,N_19314);
nor U22448 (N_22448,N_17574,N_17756);
and U22449 (N_22449,N_18864,N_19507);
xor U22450 (N_22450,N_19195,N_17911);
nand U22451 (N_22451,N_18956,N_19451);
and U22452 (N_22452,N_18753,N_19693);
and U22453 (N_22453,N_18547,N_19874);
nand U22454 (N_22454,N_17870,N_19075);
and U22455 (N_22455,N_19724,N_17877);
and U22456 (N_22456,N_19434,N_18387);
xnor U22457 (N_22457,N_18265,N_18242);
and U22458 (N_22458,N_17883,N_18745);
xnor U22459 (N_22459,N_19833,N_18784);
nor U22460 (N_22460,N_18064,N_18094);
and U22461 (N_22461,N_18433,N_17537);
and U22462 (N_22462,N_19547,N_19276);
nor U22463 (N_22463,N_17901,N_19292);
and U22464 (N_22464,N_19131,N_18516);
or U22465 (N_22465,N_19409,N_18064);
xnor U22466 (N_22466,N_19587,N_19835);
and U22467 (N_22467,N_19257,N_17942);
nor U22468 (N_22468,N_18391,N_19108);
xnor U22469 (N_22469,N_18165,N_19960);
nand U22470 (N_22470,N_18898,N_19883);
nand U22471 (N_22471,N_18366,N_19969);
nor U22472 (N_22472,N_18625,N_19703);
and U22473 (N_22473,N_18897,N_18131);
nand U22474 (N_22474,N_18382,N_18778);
and U22475 (N_22475,N_19933,N_19057);
nor U22476 (N_22476,N_18241,N_19429);
nor U22477 (N_22477,N_19908,N_19267);
nor U22478 (N_22478,N_18654,N_18789);
and U22479 (N_22479,N_17884,N_17930);
nor U22480 (N_22480,N_19896,N_17532);
nand U22481 (N_22481,N_19701,N_18295);
and U22482 (N_22482,N_18205,N_19195);
xnor U22483 (N_22483,N_18464,N_18843);
and U22484 (N_22484,N_19211,N_18610);
and U22485 (N_22485,N_19458,N_18713);
nand U22486 (N_22486,N_18037,N_19956);
nand U22487 (N_22487,N_18178,N_18081);
or U22488 (N_22488,N_19342,N_18028);
or U22489 (N_22489,N_19376,N_19314);
or U22490 (N_22490,N_17849,N_18639);
nand U22491 (N_22491,N_18913,N_18730);
xor U22492 (N_22492,N_19354,N_18682);
nor U22493 (N_22493,N_18031,N_18540);
nand U22494 (N_22494,N_17636,N_18804);
xnor U22495 (N_22495,N_17597,N_19488);
nor U22496 (N_22496,N_18255,N_19928);
nor U22497 (N_22497,N_18272,N_18413);
and U22498 (N_22498,N_19164,N_19950);
and U22499 (N_22499,N_19689,N_19385);
nor U22500 (N_22500,N_21215,N_20719);
nand U22501 (N_22501,N_22437,N_20106);
nor U22502 (N_22502,N_22242,N_20123);
nor U22503 (N_22503,N_21499,N_21203);
nor U22504 (N_22504,N_21111,N_20386);
xor U22505 (N_22505,N_22189,N_21565);
or U22506 (N_22506,N_22366,N_20000);
nand U22507 (N_22507,N_20656,N_21289);
nand U22508 (N_22508,N_22054,N_20335);
nor U22509 (N_22509,N_22383,N_21938);
nand U22510 (N_22510,N_20264,N_21720);
nand U22511 (N_22511,N_20032,N_20233);
xor U22512 (N_22512,N_22435,N_22055);
and U22513 (N_22513,N_22467,N_22352);
xor U22514 (N_22514,N_20870,N_20808);
and U22515 (N_22515,N_21612,N_21534);
or U22516 (N_22516,N_21162,N_20073);
or U22517 (N_22517,N_20469,N_20336);
xor U22518 (N_22518,N_21878,N_21476);
nand U22519 (N_22519,N_21653,N_21036);
xor U22520 (N_22520,N_21320,N_20216);
and U22521 (N_22521,N_22147,N_20684);
or U22522 (N_22522,N_21072,N_20943);
nor U22523 (N_22523,N_22248,N_22334);
and U22524 (N_22524,N_20732,N_21809);
and U22525 (N_22525,N_20434,N_20798);
nand U22526 (N_22526,N_21924,N_22221);
nand U22527 (N_22527,N_21290,N_21970);
nor U22528 (N_22528,N_20292,N_21796);
nor U22529 (N_22529,N_21827,N_20270);
nor U22530 (N_22530,N_21168,N_20312);
nand U22531 (N_22531,N_21728,N_22476);
nor U22532 (N_22532,N_21460,N_20999);
xnor U22533 (N_22533,N_21706,N_21884);
xnor U22534 (N_22534,N_22003,N_21444);
and U22535 (N_22535,N_20874,N_21234);
xor U22536 (N_22536,N_21637,N_22203);
or U22537 (N_22537,N_20321,N_20851);
or U22538 (N_22538,N_20401,N_20407);
or U22539 (N_22539,N_21449,N_20086);
or U22540 (N_22540,N_20496,N_22041);
or U22541 (N_22541,N_20856,N_20437);
and U22542 (N_22542,N_20093,N_20906);
nor U22543 (N_22543,N_20937,N_21647);
nor U22544 (N_22544,N_21031,N_21395);
xnor U22545 (N_22545,N_20258,N_21708);
or U22546 (N_22546,N_22239,N_22330);
or U22547 (N_22547,N_20368,N_20826);
or U22548 (N_22548,N_21436,N_20111);
nor U22549 (N_22549,N_20955,N_20338);
and U22550 (N_22550,N_21972,N_20900);
xnor U22551 (N_22551,N_22421,N_20374);
or U22552 (N_22552,N_20962,N_21258);
or U22553 (N_22553,N_22089,N_21097);
and U22554 (N_22554,N_22496,N_21863);
nand U22555 (N_22555,N_22103,N_21439);
nor U22556 (N_22556,N_21580,N_21002);
or U22557 (N_22557,N_22118,N_21159);
nand U22558 (N_22558,N_22349,N_21944);
or U22559 (N_22559,N_20712,N_20546);
and U22560 (N_22560,N_20717,N_20588);
xnor U22561 (N_22561,N_21759,N_22200);
xor U22562 (N_22562,N_22324,N_22303);
and U22563 (N_22563,N_21251,N_22184);
and U22564 (N_22564,N_21994,N_21898);
xnor U22565 (N_22565,N_20057,N_22283);
and U22566 (N_22566,N_20433,N_21688);
nor U22567 (N_22567,N_20326,N_20281);
nand U22568 (N_22568,N_22379,N_21362);
or U22569 (N_22569,N_20606,N_21054);
nand U22570 (N_22570,N_20161,N_20080);
nand U22571 (N_22571,N_20709,N_20979);
and U22572 (N_22572,N_21426,N_20317);
nand U22573 (N_22573,N_21236,N_22127);
or U22574 (N_22574,N_21849,N_20942);
nor U22575 (N_22575,N_20240,N_21158);
or U22576 (N_22576,N_20625,N_21797);
nand U22577 (N_22577,N_21075,N_22025);
nor U22578 (N_22578,N_20740,N_22305);
or U22579 (N_22579,N_20307,N_21262);
nand U22580 (N_22580,N_21324,N_20099);
nand U22581 (N_22581,N_20484,N_21358);
nor U22582 (N_22582,N_21364,N_21604);
or U22583 (N_22583,N_20518,N_20695);
nor U22584 (N_22584,N_22377,N_21520);
and U22585 (N_22585,N_20363,N_20403);
and U22586 (N_22586,N_21462,N_20616);
xor U22587 (N_22587,N_21427,N_21034);
nand U22588 (N_22588,N_21600,N_20542);
nor U22589 (N_22589,N_22053,N_21223);
nand U22590 (N_22590,N_22424,N_20998);
xnor U22591 (N_22591,N_21558,N_21933);
or U22592 (N_22592,N_21519,N_20824);
xor U22593 (N_22593,N_20485,N_22380);
xor U22594 (N_22594,N_21895,N_21343);
xnor U22595 (N_22595,N_20738,N_20662);
nor U22596 (N_22596,N_21213,N_21006);
and U22597 (N_22597,N_20245,N_21789);
xnor U22598 (N_22598,N_22155,N_20482);
nor U22599 (N_22599,N_20842,N_21387);
or U22600 (N_22600,N_20822,N_20373);
xnor U22601 (N_22601,N_20750,N_20811);
and U22602 (N_22602,N_21452,N_21421);
or U22603 (N_22603,N_21183,N_21498);
nand U22604 (N_22604,N_21308,N_21722);
and U22605 (N_22605,N_21160,N_21035);
nor U22606 (N_22606,N_20090,N_21335);
and U22607 (N_22607,N_22241,N_20521);
nand U22608 (N_22608,N_20038,N_20021);
xnor U22609 (N_22609,N_21388,N_20427);
and U22610 (N_22610,N_22206,N_20072);
or U22611 (N_22611,N_20014,N_22316);
and U22612 (N_22612,N_21910,N_21350);
and U22613 (N_22613,N_20002,N_20071);
nand U22614 (N_22614,N_20443,N_20609);
nand U22615 (N_22615,N_21384,N_20409);
and U22616 (N_22616,N_21840,N_22104);
xor U22617 (N_22617,N_20487,N_20253);
nor U22618 (N_22618,N_21955,N_21968);
xor U22619 (N_22619,N_21352,N_20827);
and U22620 (N_22620,N_21877,N_22255);
nand U22621 (N_22621,N_20215,N_20890);
nor U22622 (N_22622,N_21030,N_20917);
nand U22623 (N_22623,N_20379,N_20968);
nor U22624 (N_22624,N_20658,N_20790);
and U22625 (N_22625,N_21546,N_21367);
or U22626 (N_22626,N_20211,N_21517);
and U22627 (N_22627,N_20758,N_20408);
nor U22628 (N_22628,N_21004,N_21224);
or U22629 (N_22629,N_21567,N_20939);
and U22630 (N_22630,N_20938,N_21516);
xor U22631 (N_22631,N_20949,N_20774);
or U22632 (N_22632,N_22293,N_21331);
xnor U22633 (N_22633,N_22042,N_21046);
nor U22634 (N_22634,N_21577,N_21828);
nor U22635 (N_22635,N_21529,N_21678);
nor U22636 (N_22636,N_20866,N_20107);
and U22637 (N_22637,N_21091,N_22331);
or U22638 (N_22638,N_20686,N_20532);
nand U22639 (N_22639,N_20399,N_20491);
nand U22640 (N_22640,N_21470,N_20529);
xor U22641 (N_22641,N_20604,N_21463);
or U22642 (N_22642,N_21068,N_21853);
nor U22643 (N_22643,N_20982,N_21411);
and U22644 (N_22644,N_20088,N_20242);
or U22645 (N_22645,N_21680,N_22181);
xor U22646 (N_22646,N_20599,N_20903);
xnor U22647 (N_22647,N_21661,N_22073);
nand U22648 (N_22648,N_21208,N_20537);
xnor U22649 (N_22649,N_22064,N_21889);
nor U22650 (N_22650,N_20557,N_21099);
and U22651 (N_22651,N_21151,N_22492);
or U22652 (N_22652,N_20558,N_20507);
and U22653 (N_22653,N_21887,N_21926);
nor U22654 (N_22654,N_21113,N_22268);
or U22655 (N_22655,N_22230,N_22205);
nand U22656 (N_22656,N_20023,N_20204);
and U22657 (N_22657,N_21284,N_21406);
and U22658 (N_22658,N_21305,N_21978);
nor U22659 (N_22659,N_20715,N_21711);
or U22660 (N_22660,N_21486,N_20018);
nand U22661 (N_22661,N_22277,N_20193);
nand U22662 (N_22662,N_21953,N_21128);
and U22663 (N_22663,N_21296,N_21820);
nor U22664 (N_22664,N_22005,N_22083);
nor U22665 (N_22665,N_20116,N_22016);
and U22666 (N_22666,N_20648,N_20430);
xor U22667 (N_22667,N_21599,N_21611);
xnor U22668 (N_22668,N_20305,N_21836);
xor U22669 (N_22669,N_20118,N_21310);
and U22670 (N_22670,N_20197,N_20573);
or U22671 (N_22671,N_20461,N_20297);
or U22672 (N_22672,N_20497,N_22397);
and U22673 (N_22673,N_22347,N_20355);
or U22674 (N_22674,N_21266,N_22436);
or U22675 (N_22675,N_20871,N_20875);
xor U22676 (N_22676,N_21222,N_21958);
nor U22677 (N_22677,N_20711,N_21105);
and U22678 (N_22678,N_21843,N_20283);
or U22679 (N_22679,N_21148,N_20825);
nor U22680 (N_22680,N_21245,N_21174);
xnor U22681 (N_22681,N_20170,N_21240);
and U22682 (N_22682,N_20592,N_22111);
nand U22683 (N_22683,N_21503,N_20272);
nor U22684 (N_22684,N_20751,N_20419);
nand U22685 (N_22685,N_22082,N_21202);
and U22686 (N_22686,N_20294,N_22006);
nor U22687 (N_22687,N_21477,N_21620);
nor U22688 (N_22688,N_20760,N_20725);
and U22689 (N_22689,N_21846,N_20296);
xor U22690 (N_22690,N_22001,N_21133);
or U22691 (N_22691,N_20769,N_20762);
or U22692 (N_22692,N_20003,N_21301);
nor U22693 (N_22693,N_20803,N_20405);
or U22694 (N_22694,N_20202,N_20855);
nand U22695 (N_22695,N_20535,N_21020);
nand U22696 (N_22696,N_20571,N_20044);
and U22697 (N_22697,N_22350,N_20423);
or U22698 (N_22698,N_22098,N_21504);
or U22699 (N_22699,N_22307,N_22237);
and U22700 (N_22700,N_20172,N_22318);
xnor U22701 (N_22701,N_22427,N_20972);
and U22702 (N_22702,N_20356,N_21010);
nor U22703 (N_22703,N_20454,N_22049);
nand U22704 (N_22704,N_20584,N_21608);
or U22705 (N_22705,N_20350,N_21531);
or U22706 (N_22706,N_22369,N_21725);
xnor U22707 (N_22707,N_21014,N_22299);
and U22708 (N_22708,N_22168,N_20314);
nor U22709 (N_22709,N_21242,N_22039);
nand U22710 (N_22710,N_20575,N_20665);
nor U22711 (N_22711,N_21300,N_20873);
xor U22712 (N_22712,N_21227,N_22321);
nor U22713 (N_22713,N_21701,N_20340);
and U22714 (N_22714,N_21141,N_22218);
or U22715 (N_22715,N_20862,N_22478);
or U22716 (N_22716,N_20153,N_20361);
and U22717 (N_22717,N_21501,N_21261);
and U22718 (N_22718,N_20545,N_20891);
and U22719 (N_22719,N_20612,N_20964);
nand U22720 (N_22720,N_22363,N_20449);
nor U22721 (N_22721,N_20817,N_20160);
or U22722 (N_22722,N_20781,N_21859);
nor U22723 (N_22723,N_22153,N_20672);
xor U22724 (N_22724,N_21749,N_21757);
and U22725 (N_22725,N_21140,N_21287);
xor U22726 (N_22726,N_20953,N_22361);
nor U22727 (N_22727,N_20691,N_22004);
or U22728 (N_22728,N_21229,N_20411);
nand U22729 (N_22729,N_21587,N_22240);
and U22730 (N_22730,N_21682,N_21751);
nor U22731 (N_22731,N_20907,N_21966);
nand U22732 (N_22732,N_22138,N_20650);
and U22733 (N_22733,N_21093,N_21042);
nand U22734 (N_22734,N_21856,N_21790);
xor U22735 (N_22735,N_21942,N_21475);
and U22736 (N_22736,N_22123,N_21574);
xnor U22737 (N_22737,N_22133,N_21466);
xor U22738 (N_22738,N_20494,N_20499);
nor U22739 (N_22739,N_20619,N_21731);
nand U22740 (N_22740,N_20112,N_20693);
or U22741 (N_22741,N_21794,N_21694);
nor U22742 (N_22742,N_21595,N_20570);
or U22743 (N_22743,N_20467,N_22183);
nor U22744 (N_22744,N_20572,N_21636);
xnor U22745 (N_22745,N_21319,N_21511);
nor U22746 (N_22746,N_21448,N_22010);
xnor U22747 (N_22747,N_21218,N_20113);
xor U22748 (N_22748,N_21339,N_20789);
xnor U22749 (N_22749,N_20520,N_21078);
xnor U22750 (N_22750,N_20591,N_22164);
xor U22751 (N_22751,N_20782,N_20101);
or U22752 (N_22752,N_20661,N_21313);
nor U22753 (N_22753,N_22099,N_22449);
and U22754 (N_22754,N_21084,N_22308);
and U22755 (N_22755,N_21250,N_20940);
nand U22756 (N_22756,N_22429,N_20426);
nor U22757 (N_22757,N_21351,N_22490);
nand U22758 (N_22758,N_20383,N_20671);
or U22759 (N_22759,N_21408,N_21814);
nand U22760 (N_22760,N_21169,N_20841);
nor U22761 (N_22761,N_20508,N_20514);
nor U22762 (N_22762,N_21737,N_20327);
xnor U22763 (N_22763,N_22253,N_21521);
or U22764 (N_22764,N_20192,N_20230);
or U22765 (N_22765,N_21788,N_20325);
nor U22766 (N_22766,N_21542,N_21293);
or U22767 (N_22767,N_20158,N_21564);
nor U22768 (N_22768,N_21667,N_20928);
xnor U22769 (N_22769,N_21629,N_21642);
nand U22770 (N_22770,N_21440,N_21800);
xor U22771 (N_22771,N_22415,N_21530);
nor U22772 (N_22772,N_20448,N_22149);
xnor U22773 (N_22773,N_21954,N_21355);
and U22774 (N_22774,N_21095,N_21917);
xnor U22775 (N_22775,N_20420,N_22079);
nor U22776 (N_22776,N_21657,N_20334);
xor U22777 (N_22777,N_20990,N_21817);
and U22778 (N_22778,N_21412,N_22442);
and U22779 (N_22779,N_22210,N_20320);
xnor U22780 (N_22780,N_21309,N_21370);
or U22781 (N_22781,N_20269,N_21645);
or U22782 (N_22782,N_21923,N_20649);
nor U22783 (N_22783,N_20353,N_20477);
xor U22784 (N_22784,N_20306,N_22312);
and U22785 (N_22785,N_21810,N_22368);
and U22786 (N_22786,N_21246,N_22217);
nand U22787 (N_22787,N_20277,N_20867);
or U22788 (N_22788,N_22052,N_20451);
xnor U22789 (N_22789,N_21192,N_22245);
or U22790 (N_22790,N_20688,N_20188);
and U22791 (N_22791,N_22482,N_22438);
and U22792 (N_22792,N_20965,N_21114);
nand U22793 (N_22793,N_20352,N_20043);
xnor U22794 (N_22794,N_22145,N_21443);
xor U22795 (N_22795,N_21874,N_20371);
and U22796 (N_22796,N_20190,N_20095);
nand U22797 (N_22797,N_21743,N_22443);
or U22798 (N_22798,N_20198,N_22086);
nor U22799 (N_22799,N_21323,N_22493);
and U22800 (N_22800,N_20179,N_21256);
or U22801 (N_22801,N_21485,N_20007);
xnor U22802 (N_22802,N_20837,N_21812);
nor U22803 (N_22803,N_21392,N_21755);
and U22804 (N_22804,N_20015,N_22199);
xnor U22805 (N_22805,N_21959,N_21570);
nor U22806 (N_22806,N_22178,N_21649);
xor U22807 (N_22807,N_20039,N_22469);
or U22808 (N_22808,N_21249,N_20651);
or U22809 (N_22809,N_20033,N_20341);
xor U22810 (N_22810,N_20624,N_20562);
nor U22811 (N_22811,N_20354,N_20655);
xor U22812 (N_22812,N_20696,N_20452);
and U22813 (N_22813,N_20110,N_22117);
nand U22814 (N_22814,N_20142,N_21956);
xnor U22815 (N_22815,N_20675,N_21527);
and U22816 (N_22816,N_20797,N_20077);
or U22817 (N_22817,N_21920,N_21062);
or U22818 (N_22818,N_21484,N_20315);
or U22819 (N_22819,N_20780,N_22002);
nand U22820 (N_22820,N_22284,N_21007);
nand U22821 (N_22821,N_22074,N_21163);
and U22822 (N_22822,N_20159,N_21915);
nand U22823 (N_22823,N_20309,N_20605);
or U22824 (N_22824,N_20530,N_20201);
nor U22825 (N_22825,N_21146,N_20303);
nand U22826 (N_22826,N_20929,N_21416);
nand U22827 (N_22827,N_22141,N_20767);
or U22828 (N_22828,N_22087,N_20257);
nor U22829 (N_22829,N_20611,N_20898);
xor U22830 (N_22830,N_20385,N_20276);
and U22831 (N_22831,N_20578,N_22109);
xnor U22832 (N_22832,N_20091,N_20249);
nand U22833 (N_22833,N_22475,N_20722);
and U22834 (N_22834,N_21523,N_22256);
and U22835 (N_22835,N_20474,N_21196);
and U22836 (N_22836,N_20028,N_21945);
nor U22837 (N_22837,N_21115,N_21278);
or U22838 (N_22838,N_20902,N_20041);
xor U22839 (N_22839,N_20777,N_21764);
nand U22840 (N_22840,N_20214,N_21627);
or U22841 (N_22841,N_21779,N_20271);
and U22842 (N_22842,N_21110,N_20236);
or U22843 (N_22843,N_20417,N_20935);
or U22844 (N_22844,N_20422,N_20613);
nand U22845 (N_22845,N_21615,N_22214);
and U22846 (N_22846,N_21098,N_20127);
nand U22847 (N_22847,N_22365,N_22468);
and U22848 (N_22848,N_20210,N_22357);
nand U22849 (N_22849,N_20641,N_20831);
xnor U22850 (N_22850,N_20846,N_20540);
or U22851 (N_22851,N_20328,N_20582);
nand U22852 (N_22852,N_20676,N_21023);
and U22853 (N_22853,N_21535,N_21109);
or U22854 (N_22854,N_21712,N_22121);
nand U22855 (N_22855,N_21494,N_22048);
or U22856 (N_22856,N_22372,N_21777);
and U22857 (N_22857,N_20428,N_20848);
xnor U22858 (N_22858,N_20820,N_21458);
xnor U22859 (N_22859,N_22198,N_20680);
xor U22860 (N_22860,N_20527,N_20199);
or U22861 (N_22861,N_21606,N_22119);
or U22862 (N_22862,N_21383,N_20748);
xor U22863 (N_22863,N_20012,N_21487);
xnor U22864 (N_22864,N_22332,N_20629);
nand U22865 (N_22865,N_22174,N_22453);
nor U22866 (N_22866,N_21260,N_20079);
xor U22867 (N_22867,N_21132,N_22414);
xnor U22868 (N_22868,N_20255,N_21964);
nor U22869 (N_22869,N_20724,N_21893);
nor U22870 (N_22870,N_21778,N_21671);
nor U22871 (N_22871,N_20109,N_22207);
or U22872 (N_22872,N_21943,N_21316);
and U22873 (N_22873,N_20047,N_20429);
or U22874 (N_22874,N_20714,N_21340);
nor U22875 (N_22875,N_22296,N_21268);
or U22876 (N_22876,N_21610,N_20122);
and U22877 (N_22877,N_20146,N_20960);
or U22878 (N_22878,N_21700,N_20246);
and U22879 (N_22879,N_21134,N_20476);
xnor U22880 (N_22880,N_21125,N_20016);
xnor U22881 (N_22881,N_20138,N_22474);
or U22882 (N_22882,N_20905,N_20961);
xor U22883 (N_22883,N_20515,N_22439);
and U22884 (N_22884,N_20225,N_20776);
nand U22885 (N_22885,N_21597,N_22246);
nor U22886 (N_22886,N_21407,N_22445);
or U22887 (N_22887,N_22481,N_20351);
or U22888 (N_22888,N_20683,N_21995);
or U22889 (N_22889,N_22250,N_20463);
and U22890 (N_22890,N_20627,N_21337);
nand U22891 (N_22891,N_22432,N_20205);
xnor U22892 (N_22892,N_22498,N_21526);
and U22893 (N_22893,N_20128,N_21304);
nand U22894 (N_22894,N_22354,N_22345);
nand U22895 (N_22895,N_20522,N_21438);
or U22896 (N_22896,N_22459,N_20918);
nand U22897 (N_22897,N_20988,N_22219);
xor U22898 (N_22898,N_22208,N_20533);
or U22899 (N_22899,N_21419,N_21903);
nor U22900 (N_22900,N_20730,N_22322);
and U22901 (N_22901,N_21235,N_22272);
nor U22902 (N_22902,N_20559,N_20729);
or U22903 (N_22903,N_21121,N_21973);
xnor U22904 (N_22904,N_22077,N_21157);
and U22905 (N_22905,N_22384,N_20194);
nand U22906 (N_22906,N_20300,N_21461);
and U22907 (N_22907,N_22461,N_20728);
nor U22908 (N_22908,N_20547,N_20085);
or U22909 (N_22909,N_21135,N_20096);
nor U22910 (N_22910,N_20025,N_20506);
and U22911 (N_22911,N_21210,N_20059);
and U22912 (N_22912,N_22197,N_21857);
nand U22913 (N_22913,N_22146,N_21518);
nand U22914 (N_22914,N_22460,N_20785);
xnor U22915 (N_22915,N_22234,N_20697);
nand U22916 (N_22916,N_21333,N_21758);
or U22917 (N_22917,N_21080,N_20332);
or U22918 (N_22918,N_21022,N_21451);
xnor U22919 (N_22919,N_21211,N_21239);
and U22920 (N_22920,N_21417,N_20897);
and U22921 (N_22921,N_20839,N_21404);
xnor U22922 (N_22922,N_22340,N_20156);
and U22923 (N_22923,N_21602,N_20997);
and U22924 (N_22924,N_22222,N_21118);
and U22925 (N_22925,N_21858,N_21635);
and U22926 (N_22926,N_20069,N_22097);
nand U22927 (N_22927,N_20944,N_21361);
and U22928 (N_22928,N_22051,N_20238);
nand U22929 (N_22929,N_20791,N_22209);
and U22930 (N_22930,N_21745,N_21559);
and U22931 (N_22931,N_22311,N_22182);
or U22932 (N_22932,N_21540,N_22408);
nor U22933 (N_22933,N_21232,N_22489);
nand U22934 (N_22934,N_21150,N_21182);
nand U22935 (N_22935,N_20930,N_20395);
nor U22936 (N_22936,N_20698,N_20501);
and U22937 (N_22937,N_21543,N_20920);
xnor U22938 (N_22938,N_21058,N_21490);
or U22939 (N_22939,N_22423,N_21515);
and U22940 (N_22940,N_20082,N_22069);
nand U22941 (N_22941,N_22446,N_22126);
nor U22942 (N_22942,N_21549,N_22407);
xnor U22943 (N_22943,N_21489,N_21738);
nor U22944 (N_22944,N_20816,N_21292);
xnor U22945 (N_22945,N_21969,N_21129);
or U22946 (N_22946,N_22374,N_20478);
and U22947 (N_22947,N_21867,N_20889);
and U22948 (N_22948,N_22094,N_21430);
nor U22949 (N_22949,N_21935,N_22401);
or U22950 (N_22950,N_22251,N_21879);
xnor U22951 (N_22951,N_20794,N_21069);
xnor U22952 (N_22952,N_20313,N_20319);
or U22953 (N_22953,N_21456,N_21767);
or U22954 (N_22954,N_21663,N_21435);
nor U22955 (N_22955,N_21727,N_20726);
xor U22956 (N_22956,N_20548,N_21666);
nand U22957 (N_22957,N_21643,N_21550);
or U22958 (N_22958,N_20094,N_20853);
xor U22959 (N_22959,N_20983,N_21868);
nor U22960 (N_22960,N_21414,N_21117);
xor U22961 (N_22961,N_21116,N_21345);
xnor U22962 (N_22962,N_20195,N_21689);
xor U22963 (N_22963,N_22297,N_22247);
nand U22964 (N_22964,N_21353,N_22270);
nor U22965 (N_22965,N_22488,N_21659);
and U22966 (N_22966,N_21692,N_20177);
nor U22967 (N_22967,N_21673,N_21782);
and U22968 (N_22968,N_21616,N_22269);
nand U22969 (N_22969,N_22433,N_21492);
nor U22970 (N_22970,N_21660,N_20349);
and U22971 (N_22971,N_21376,N_20931);
and U22972 (N_22972,N_21382,N_22391);
nor U22973 (N_22973,N_20690,N_22046);
nand U22974 (N_22974,N_20217,N_21664);
nand U22975 (N_22975,N_20348,N_21593);
and U22976 (N_22976,N_22327,N_21713);
xnor U22977 (N_22977,N_20049,N_21894);
nand U22978 (N_22978,N_21613,N_22281);
nor U22979 (N_22979,N_20125,N_20904);
or U22980 (N_22980,N_21209,N_21601);
or U22981 (N_22981,N_22080,N_21997);
nor U22982 (N_22982,N_21735,N_21582);
xnor U22983 (N_22983,N_21379,N_22151);
or U22984 (N_22984,N_22409,N_21070);
xor U22985 (N_22985,N_22011,N_20343);
or U22986 (N_22986,N_21124,N_22233);
and U22987 (N_22987,N_21061,N_21269);
nor U22988 (N_22988,N_20001,N_21907);
xnor U22989 (N_22989,N_22226,N_21391);
and U22990 (N_22990,N_21328,N_20908);
nand U22991 (N_22991,N_22314,N_22425);
or U22992 (N_22992,N_20286,N_21420);
nand U22993 (N_22993,N_20062,N_20489);
nand U22994 (N_22994,N_21152,N_21094);
and U22995 (N_22995,N_21573,N_20861);
xor U22996 (N_22996,N_21509,N_22390);
and U22997 (N_22997,N_20436,N_21424);
and U22998 (N_22998,N_21488,N_20947);
xor U22999 (N_22999,N_22291,N_21177);
nand U23000 (N_23000,N_22114,N_20432);
nor U23001 (N_23001,N_20759,N_21244);
nor U23002 (N_23002,N_20102,N_22419);
nor U23003 (N_23003,N_21880,N_20565);
and U23004 (N_23004,N_20219,N_20011);
nand U23005 (N_23005,N_22466,N_21690);
nand U23006 (N_23006,N_22454,N_21831);
or U23007 (N_23007,N_22388,N_20035);
and U23008 (N_23008,N_20322,N_22170);
xnor U23009 (N_23009,N_20134,N_22201);
nand U23010 (N_23010,N_21403,N_21916);
and U23011 (N_23011,N_21555,N_22342);
nor U23012 (N_23012,N_21841,N_20845);
nand U23013 (N_23013,N_22047,N_20027);
nand U23014 (N_23014,N_22406,N_20615);
nand U23015 (N_23015,N_21622,N_22457);
or U23016 (N_23016,N_20912,N_22285);
nor U23017 (N_23017,N_20115,N_21123);
nor U23018 (N_23018,N_20589,N_20132);
nor U23019 (N_23019,N_21992,N_21307);
nand U23020 (N_23020,N_21609,N_20168);
nor U23021 (N_23021,N_22115,N_22140);
or U23022 (N_23022,N_20455,N_21628);
xnor U23023 (N_23023,N_21001,N_22040);
or U23024 (N_23024,N_21698,N_21869);
nand U23025 (N_23025,N_20865,N_21056);
or U23026 (N_23026,N_21130,N_20135);
and U23027 (N_23027,N_22030,N_20282);
xnor U23028 (N_23028,N_22456,N_22485);
nand U23029 (N_23029,N_21178,N_20768);
or U23030 (N_23030,N_22403,N_22173);
nor U23031 (N_23031,N_20736,N_20129);
or U23032 (N_23032,N_21327,N_20223);
xnor U23033 (N_23033,N_21630,N_21928);
or U23034 (N_23034,N_20886,N_21537);
xnor U23035 (N_23035,N_21285,N_22271);
or U23036 (N_23036,N_20669,N_21716);
nand U23037 (N_23037,N_21100,N_21592);
or U23038 (N_23038,N_20973,N_20681);
and U23039 (N_23039,N_20203,N_21065);
xor U23040 (N_23040,N_22187,N_20752);
nand U23041 (N_23041,N_20707,N_21422);
and U23042 (N_23042,N_21963,N_20439);
or U23043 (N_23043,N_22020,N_21255);
nor U23044 (N_23044,N_20076,N_21156);
xnor U23045 (N_23045,N_21977,N_20869);
nand U23046 (N_23046,N_21119,N_21142);
xor U23047 (N_23047,N_22033,N_21808);
xor U23048 (N_23048,N_21805,N_22068);
and U23049 (N_23049,N_21584,N_20390);
nand U23050 (N_23050,N_21066,N_21044);
nand U23051 (N_23051,N_20745,N_21747);
and U23052 (N_23052,N_22280,N_20381);
xor U23053 (N_23053,N_22066,N_21979);
nor U23054 (N_23054,N_21219,N_20008);
nand U23055 (N_23055,N_22487,N_22009);
and U23056 (N_23056,N_22032,N_22093);
nand U23057 (N_23057,N_21672,N_21514);
and U23058 (N_23058,N_21848,N_20783);
or U23059 (N_23059,N_21165,N_20359);
nor U23060 (N_23060,N_22394,N_20863);
nand U23061 (N_23061,N_21974,N_20534);
nor U23062 (N_23062,N_21579,N_22274);
or U23063 (N_23063,N_22252,N_21144);
and U23064 (N_23064,N_22348,N_21940);
and U23065 (N_23065,N_20318,N_21480);
xnor U23066 (N_23066,N_20224,N_21639);
nor U23067 (N_23067,N_21341,N_21164);
nor U23068 (N_23068,N_21468,N_22220);
or U23069 (N_23069,N_21539,N_20206);
xor U23070 (N_23070,N_20273,N_20976);
xnor U23071 (N_23071,N_20460,N_21413);
nor U23072 (N_23072,N_22278,N_20844);
nor U23073 (N_23073,N_21786,N_20879);
or U23074 (N_23074,N_20054,N_20812);
nand U23075 (N_23075,N_20458,N_20652);
nand U23076 (N_23076,N_21281,N_21077);
or U23077 (N_23077,N_21998,N_21453);
and U23078 (N_23078,N_20843,N_20576);
nor U23079 (N_23079,N_22084,N_22152);
and U23080 (N_23080,N_20823,N_21000);
nor U23081 (N_23081,N_21332,N_21060);
and U23082 (N_23082,N_21623,N_21282);
xor U23083 (N_23083,N_21389,N_20992);
nand U23084 (N_23084,N_20175,N_22328);
nand U23085 (N_23085,N_22440,N_20017);
nor U23086 (N_23086,N_21108,N_21154);
and U23087 (N_23087,N_21882,N_21029);
and U23088 (N_23088,N_21906,N_22216);
xor U23089 (N_23089,N_21041,N_20596);
and U23090 (N_23090,N_22260,N_20525);
nor U23091 (N_23091,N_21045,N_21482);
nor U23092 (N_23092,N_21598,N_20259);
nor U23093 (N_23093,N_22238,N_20813);
or U23094 (N_23094,N_22422,N_20208);
or U23095 (N_23095,N_21247,N_21750);
nor U23096 (N_23096,N_21771,N_21982);
and U23097 (N_23097,N_22185,N_21371);
or U23098 (N_23098,N_22276,N_20144);
nand U23099 (N_23099,N_22279,N_21603);
nor U23100 (N_23100,N_20289,N_20786);
nand U23101 (N_23101,N_21005,N_20637);
and U23102 (N_23102,N_22008,N_21948);
nor U23103 (N_23103,N_22150,N_22204);
nor U23104 (N_23104,N_20066,N_20554);
xnor U23105 (N_23105,N_20950,N_20254);
or U23106 (N_23106,N_21225,N_22371);
and U23107 (N_23107,N_22050,N_22463);
xor U23108 (N_23108,N_21173,N_20754);
and U23109 (N_23109,N_22302,N_21633);
nor U23110 (N_23110,N_22249,N_21562);
and U23111 (N_23111,N_21908,N_20104);
and U23112 (N_23112,N_20150,N_22258);
nand U23113 (N_23113,N_20967,N_20105);
or U23114 (N_23114,N_21762,N_20868);
nand U23115 (N_23115,N_21829,N_22395);
or U23116 (N_23116,N_20013,N_22315);
xnor U23117 (N_23117,N_20922,N_21699);
xor U23118 (N_23118,N_21557,N_20796);
xnor U23119 (N_23119,N_20311,N_21568);
or U23120 (N_23120,N_21905,N_21264);
xnor U23121 (N_23121,N_21703,N_22313);
xor U23122 (N_23122,N_21143,N_21206);
nand U23123 (N_23123,N_20004,N_20787);
xnor U23124 (N_23124,N_21506,N_20169);
and U23125 (N_23125,N_21838,N_20706);
or U23126 (N_23126,N_22072,N_21781);
and U23127 (N_23127,N_21252,N_21053);
xnor U23128 (N_23128,N_21662,N_22451);
and U23129 (N_23129,N_21259,N_20958);
nor U23130 (N_23130,N_20218,N_21932);
nor U23131 (N_23131,N_21936,N_22416);
and U23132 (N_23132,N_21106,N_20678);
nand U23133 (N_23133,N_21648,N_21990);
nor U23134 (N_23134,N_21265,N_20376);
or U23135 (N_23135,N_21563,N_20833);
nand U23136 (N_23136,N_20747,N_22262);
or U23137 (N_23137,N_21742,N_22091);
and U23138 (N_23138,N_21194,N_21696);
nand U23139 (N_23139,N_21798,N_20486);
or U23140 (N_23140,N_20183,N_20945);
xor U23141 (N_23141,N_20561,N_20810);
and U23142 (N_23142,N_21638,N_20524);
and U23143 (N_23143,N_21483,N_22356);
xor U23144 (N_23144,N_20366,N_21822);
nor U23145 (N_23145,N_20544,N_21746);
and U23146 (N_23146,N_21866,N_20620);
xnor U23147 (N_23147,N_20574,N_22085);
xor U23148 (N_23148,N_22063,N_22113);
xnor U23149 (N_23149,N_21803,N_20378);
nor U23150 (N_23150,N_21090,N_20773);
or U23151 (N_23151,N_20959,N_20700);
and U23152 (N_23152,N_20749,N_20626);
and U23153 (N_23153,N_21588,N_22061);
nand U23154 (N_23154,N_22358,N_20415);
xnor U23155 (N_23155,N_21583,N_20659);
or U23156 (N_23156,N_20806,N_21533);
xnor U23157 (N_23157,N_21832,N_21280);
and U23158 (N_23158,N_20182,N_21038);
nand U23159 (N_23159,N_20167,N_20957);
or U23160 (N_23160,N_21631,N_20878);
xnor U23161 (N_23161,N_21188,N_21548);
and U23162 (N_23162,N_21719,N_21983);
nand U23163 (N_23163,N_21214,N_20597);
or U23164 (N_23164,N_20744,N_20053);
and U23165 (N_23165,N_20721,N_22287);
or U23166 (N_23166,N_21377,N_21496);
xnor U23167 (N_23167,N_20598,N_20595);
or U23168 (N_23168,N_20640,N_22112);
nor U23169 (N_23169,N_20603,N_22023);
xnor U23170 (N_23170,N_20391,N_22136);
and U23171 (N_23171,N_22171,N_21122);
xnor U23172 (N_23172,N_22130,N_20555);
xnor U23173 (N_23173,N_20809,N_22062);
nor U23174 (N_23174,N_20145,N_20131);
nor U23175 (N_23175,N_22470,N_21683);
or U23176 (N_23176,N_21765,N_20425);
nand U23177 (N_23177,N_22329,N_20392);
and U23178 (N_23178,N_20453,N_20268);
or U23179 (N_23179,N_20850,N_20985);
nor U23180 (N_23180,N_22060,N_22161);
or U23181 (N_23181,N_20256,N_22355);
xnor U23182 (N_23182,N_21048,N_22343);
nand U23183 (N_23183,N_20472,N_21221);
nor U23184 (N_23184,N_21952,N_21043);
or U23185 (N_23185,N_20916,N_22065);
nand U23186 (N_23186,N_21500,N_21120);
and U23187 (N_23187,N_21575,N_21009);
nand U23188 (N_23188,N_21721,N_21295);
and U23189 (N_23189,N_20860,N_20178);
and U23190 (N_23190,N_20157,N_22142);
or U23191 (N_23191,N_22095,N_20050);
or U23192 (N_23192,N_21198,N_21248);
or U23193 (N_23193,N_22034,N_20893);
nor U23194 (N_23194,N_20852,N_21525);
nor U23195 (N_23195,N_20926,N_21896);
nand U23196 (N_23196,N_21199,N_21189);
or U23197 (N_23197,N_21640,N_21946);
and U23198 (N_23198,N_21441,N_22037);
or U23199 (N_23199,N_21815,N_20070);
xnor U23200 (N_23200,N_21085,N_20673);
xnor U23201 (N_23201,N_21147,N_21459);
nor U23202 (N_23202,N_21270,N_21748);
nor U23203 (N_23203,N_20723,N_22447);
xor U23204 (N_23204,N_21754,N_21913);
or U23205 (N_23205,N_20733,N_21318);
nor U23206 (N_23206,N_20293,N_22228);
and U23207 (N_23207,N_20566,N_21204);
and U23208 (N_23208,N_21847,N_21545);
nor U23209 (N_23209,N_21704,N_20872);
nand U23210 (N_23210,N_22480,N_20670);
xnor U23211 (N_23211,N_21715,N_21071);
xnor U23212 (N_23212,N_21784,N_21912);
nor U23213 (N_23213,N_20165,N_22159);
xor U23214 (N_23214,N_21176,N_20372);
nand U23215 (N_23215,N_21450,N_22154);
nand U23216 (N_23216,N_21658,N_21378);
or U23217 (N_23217,N_21734,N_21844);
and U23218 (N_23218,N_20795,N_20468);
or U23219 (N_23219,N_22106,N_21027);
nand U23220 (N_23220,N_22071,N_20884);
xor U23221 (N_23221,N_21685,N_22180);
or U23222 (N_23222,N_21513,N_21442);
nor U23223 (N_23223,N_22323,N_20480);
nand U23224 (N_23224,N_21886,N_22132);
xnor U23225 (N_23225,N_20876,N_20471);
nor U23226 (N_23226,N_22310,N_20667);
nor U23227 (N_23227,N_21830,N_21074);
xor U23228 (N_23228,N_21544,N_20541);
nand U23229 (N_23229,N_20196,N_21510);
nor U23230 (N_23230,N_20213,N_21399);
nand U23231 (N_23231,N_20152,N_21679);
or U23232 (N_23232,N_21471,N_20229);
nand U23233 (N_23233,N_20222,N_20414);
nor U23234 (N_23234,N_20187,N_20761);
and U23235 (N_23235,N_21052,N_20438);
xor U23236 (N_23236,N_20668,N_20583);
and U23237 (N_23237,N_20466,N_21230);
nor U23238 (N_23238,N_20642,N_22124);
nand U23239 (N_23239,N_22202,N_20089);
and U23240 (N_23240,N_21775,N_21541);
and U23241 (N_23241,N_21446,N_22497);
or U23242 (N_23242,N_20830,N_22231);
xor U23243 (N_23243,N_20377,N_22289);
and U23244 (N_23244,N_20228,N_22398);
or U23245 (N_23245,N_20247,N_21818);
nor U23246 (N_23246,N_21137,N_22232);
nand U23247 (N_23247,N_21410,N_20657);
nor U23248 (N_23248,N_20818,N_20045);
or U23249 (N_23249,N_21656,N_20237);
and U23250 (N_23250,N_21740,N_20097);
and U23251 (N_23251,N_21409,N_21233);
nor U23252 (N_23252,N_21479,N_20560);
and U23253 (N_23253,N_20299,N_21816);
nand U23254 (N_23254,N_21092,N_20720);
and U23255 (N_23255,N_20511,N_22426);
nor U23256 (N_23256,N_20954,N_20763);
nand U23257 (N_23257,N_20261,N_22188);
nand U23258 (N_23258,N_21175,N_22341);
nand U23259 (N_23259,N_20705,N_20819);
nand U23260 (N_23260,N_21674,N_21373);
nor U23261 (N_23261,N_20406,N_21842);
nor U23262 (N_23262,N_21497,N_20633);
or U23263 (N_23263,N_21049,N_20357);
or U23264 (N_23264,N_21984,N_21714);
xnor U23265 (N_23265,N_20367,N_21845);
nor U23266 (N_23266,N_21346,N_20737);
xnor U23267 (N_23267,N_21271,N_22192);
xnor U23268 (N_23268,N_21507,N_20263);
and U23269 (N_23269,N_20221,N_20009);
nor U23270 (N_23270,N_20171,N_20046);
xnor U23271 (N_23271,N_21238,N_21187);
xnor U23272 (N_23272,N_21670,N_22417);
nor U23273 (N_23273,N_21756,N_21733);
xor U23274 (N_23274,N_20260,N_20645);
nand U23275 (N_23275,N_20838,N_20800);
xnor U23276 (N_23276,N_20513,N_22351);
xor U23277 (N_23277,N_20384,N_21149);
nor U23278 (N_23278,N_20617,N_20279);
or U23279 (N_23279,N_21941,N_21621);
nor U23280 (N_23280,N_22288,N_22101);
or U23281 (N_23281,N_20569,N_20504);
nor U23282 (N_23282,N_22035,N_22370);
or U23283 (N_23283,N_21228,N_21929);
nand U23284 (N_23284,N_20250,N_21651);
and U23285 (N_23285,N_20840,N_21181);
and U23286 (N_23286,N_22484,N_21329);
or U23287 (N_23287,N_22265,N_20989);
or U23288 (N_23288,N_21019,N_20019);
xor U23289 (N_23289,N_20450,N_21291);
nand U23290 (N_23290,N_21418,N_21821);
xor U23291 (N_23291,N_21297,N_22418);
xor U23292 (N_23292,N_20784,N_21999);
nand U23293 (N_23293,N_22028,N_20601);
and U23294 (N_23294,N_22193,N_20755);
xor U23295 (N_23295,N_21474,N_21312);
xnor U23296 (N_23296,N_21707,N_21852);
or U23297 (N_23297,N_21338,N_20987);
nand U23298 (N_23298,N_20022,N_22134);
and U23299 (N_23299,N_22190,N_22367);
nand U23300 (N_23300,N_21314,N_20026);
and U23301 (N_23301,N_21922,N_20490);
or U23302 (N_23302,N_20996,N_21274);
xnor U23303 (N_23303,N_22166,N_20509);
nand U23304 (N_23304,N_21652,N_20910);
and U23305 (N_23305,N_21051,N_21625);
nor U23306 (N_23306,N_21325,N_21996);
xnor U23307 (N_23307,N_21677,N_20971);
or U23308 (N_23308,N_21883,N_20682);
xnor U23309 (N_23309,N_21962,N_21806);
or U23310 (N_23310,N_20731,N_21554);
and U23311 (N_23311,N_21695,N_20117);
and U23312 (N_23312,N_21032,N_20631);
xor U23313 (N_23313,N_20174,N_21890);
or U23314 (N_23314,N_20644,N_20885);
nor U23315 (N_23315,N_20442,N_21478);
xnor U23316 (N_23316,N_22045,N_20934);
and U23317 (N_23317,N_21632,N_20936);
nand U23318 (N_23318,N_21381,N_20495);
nand U23319 (N_23319,N_21493,N_21021);
nand U23320 (N_23320,N_21988,N_22129);
nor U23321 (N_23321,N_21947,N_22385);
nand U23322 (N_23322,N_20854,N_20739);
xor U23323 (N_23323,N_21170,N_20465);
nand U23324 (N_23324,N_20539,N_20139);
or U23325 (N_23325,N_20741,N_20778);
and U23326 (N_23326,N_22021,N_20946);
xnor U23327 (N_23327,N_21760,N_21987);
nand U23328 (N_23328,N_22412,N_21804);
nand U23329 (N_23329,N_22301,N_22088);
xor U23330 (N_23330,N_21835,N_20986);
nand U23331 (N_23331,N_21457,N_22491);
or U23332 (N_23332,N_22186,N_20503);
xor U23333 (N_23333,N_22452,N_21207);
nand U23334 (N_23334,N_21572,N_22472);
or U23335 (N_23335,N_21865,N_20991);
xor U23336 (N_23336,N_20804,N_20074);
nand U23337 (N_23337,N_22100,N_21089);
xor U23338 (N_23338,N_20440,N_21283);
or U23339 (N_23339,N_22344,N_21949);
nand U23340 (N_23340,N_20473,N_20124);
nor U23341 (N_23341,N_21617,N_22326);
nand U23342 (N_23342,N_21911,N_20184);
nor U23343 (N_23343,N_20756,N_21991);
nor U23344 (N_23344,N_20679,N_21684);
nand U23345 (N_23345,N_21675,N_22325);
and U23346 (N_23346,N_21254,N_21981);
and U23347 (N_23347,N_21040,N_21243);
and U23348 (N_23348,N_21434,N_21311);
and U23349 (N_23349,N_21791,N_21200);
and U23350 (N_23350,N_21139,N_20024);
or U23351 (N_23351,N_21342,N_20410);
nor U23352 (N_23352,N_20151,N_22364);
nor U23353 (N_23353,N_22162,N_20674);
and U23354 (N_23354,N_20226,N_21083);
nand U23355 (N_23355,N_22157,N_21927);
nor U23356 (N_23356,N_20829,N_21465);
and U23357 (N_23357,N_21566,N_22179);
nand U23358 (N_23358,N_20621,N_20251);
nor U23359 (N_23359,N_21374,N_21975);
xor U23360 (N_23360,N_21980,N_20280);
nor U23361 (N_23361,N_21298,N_21015);
or U23362 (N_23362,N_20666,N_21145);
xor U23363 (N_23363,N_21096,N_20799);
and U23364 (N_23364,N_22462,N_22254);
xor U23365 (N_23365,N_21763,N_21082);
or U23366 (N_23366,N_20006,N_21013);
nor U23367 (N_23367,N_22375,N_22125);
xnor U23368 (N_23368,N_20290,N_20994);
nor U23369 (N_23369,N_20037,N_21288);
xor U23370 (N_23370,N_20052,N_21131);
xnor U23371 (N_23371,N_20010,N_20913);
and U23372 (N_23372,N_20743,N_21286);
or U23373 (N_23373,N_22434,N_20030);
or U23374 (N_23374,N_20970,N_20821);
and U23375 (N_23375,N_20239,N_22413);
and U23376 (N_23376,N_20488,N_21366);
nor U23377 (N_23377,N_21039,N_21957);
xnor U23378 (N_23378,N_21851,N_22483);
nand U23379 (N_23379,N_20636,N_20646);
xnor U23380 (N_23380,N_20618,N_20516);
and U23381 (N_23381,N_20653,N_21241);
and U23382 (N_23382,N_21195,N_21536);
xnor U23383 (N_23383,N_20241,N_21578);
xor U23384 (N_23384,N_21590,N_20398);
or U23385 (N_23385,N_20864,N_22057);
nor U23386 (N_23386,N_21365,N_20828);
nand U23387 (N_23387,N_21161,N_21872);
nor U23388 (N_23388,N_20858,N_22373);
xor U23389 (N_23389,N_22116,N_20551);
and U23390 (N_23390,N_21547,N_20227);
and U23391 (N_23391,N_22018,N_22448);
nand U23392 (N_23392,N_21423,N_20543);
or U23393 (N_23393,N_22076,N_22386);
and U23394 (N_23394,N_20523,N_22267);
and U23395 (N_23395,N_21753,N_22455);
nor U23396 (N_23396,N_20492,N_22381);
and U23397 (N_23397,N_22044,N_22135);
nand U23398 (N_23398,N_21862,N_21467);
nand U23399 (N_23399,N_21303,N_20029);
xnor U23400 (N_23400,N_22306,N_20552);
nand U23401 (N_23401,N_22211,N_21726);
xnor U23402 (N_23402,N_20051,N_21086);
or U23403 (N_23403,N_20288,N_21472);
nand U23404 (N_23404,N_21669,N_20120);
or U23405 (N_23405,N_21774,N_22378);
and U23406 (N_23406,N_21201,N_21855);
nor U23407 (N_23407,N_22458,N_21985);
or U23408 (N_23408,N_21101,N_22261);
and U23409 (N_23409,N_20608,N_21349);
xor U23410 (N_23410,N_22137,N_20346);
nor U23411 (N_23411,N_21326,N_20149);
nand U23412 (N_23412,N_21697,N_20563);
nor U23413 (N_23413,N_22031,N_20189);
nor U23414 (N_23414,N_21191,N_20103);
nor U23415 (N_23415,N_21397,N_22194);
or U23416 (N_23416,N_21033,N_21909);
nor U23417 (N_23417,N_20232,N_20362);
or U23418 (N_23418,N_20538,N_22360);
and U23419 (N_23419,N_20301,N_20382);
xor U23420 (N_23420,N_20528,N_20278);
and U23421 (N_23421,N_21398,N_22471);
xor U23422 (N_23422,N_21402,N_21184);
or U23423 (N_23423,N_22019,N_20975);
xor U23424 (N_23424,N_21986,N_20063);
and U23425 (N_23425,N_21429,N_21646);
nor U23426 (N_23426,N_20248,N_22295);
nor U23427 (N_23427,N_20896,N_21112);
nor U23428 (N_23428,N_21012,N_20483);
nor U23429 (N_23429,N_22128,N_22362);
or U23430 (N_23430,N_21823,N_20753);
nand U23431 (N_23431,N_20330,N_20607);
nor U23432 (N_23432,N_22017,N_20100);
and U23433 (N_23433,N_21914,N_20447);
or U23434 (N_23434,N_20126,N_22172);
xor U23435 (N_23435,N_21897,N_22212);
or U23436 (N_23436,N_21581,N_21088);
xor U23437 (N_23437,N_20344,N_21138);
and U23438 (N_23438,N_21028,N_20164);
xnor U23439 (N_23439,N_22393,N_20287);
nand U23440 (N_23440,N_20284,N_21103);
nand U23441 (N_23441,N_21390,N_22078);
nand U23442 (N_23442,N_21495,N_21594);
nor U23443 (N_23443,N_20186,N_21237);
and U23444 (N_23444,N_20628,N_21741);
nor U23445 (N_23445,N_20083,N_21605);
xor U23446 (N_23446,N_21079,N_20963);
xnor U23447 (N_23447,N_21919,N_21315);
nor U23448 (N_23448,N_22430,N_22473);
xnor U23449 (N_23449,N_21216,N_22450);
nor U23450 (N_23450,N_22346,N_20067);
or U23451 (N_23451,N_21860,N_20772);
xor U23452 (N_23452,N_20358,N_20663);
nand U23453 (N_23453,N_21155,N_21837);
or U23454 (N_23454,N_20771,N_22404);
or U23455 (N_23455,N_20087,N_20857);
nand U23456 (N_23456,N_22320,N_20519);
nand U23457 (N_23457,N_21357,N_21172);
xor U23458 (N_23458,N_20654,N_21447);
or U23459 (N_23459,N_22464,N_20899);
and U23460 (N_23460,N_20412,N_21925);
xnor U23461 (N_23461,N_20924,N_20166);
nor U23462 (N_23462,N_20342,N_21665);
xnor U23463 (N_23463,N_22102,N_20369);
nand U23464 (N_23464,N_20517,N_21873);
nor U23465 (N_23465,N_22499,N_21787);
xnor U23466 (N_23466,N_22014,N_20677);
nand U23467 (N_23467,N_20234,N_22405);
nand U23468 (N_23468,N_20331,N_20580);
xor U23469 (N_23469,N_22389,N_21037);
nor U23470 (N_23470,N_20081,N_22191);
nand U23471 (N_23471,N_22012,N_22335);
nand U23472 (N_23472,N_22013,N_21081);
nand U23473 (N_23473,N_20285,N_20710);
or U23474 (N_23474,N_20788,N_20005);
nand U23475 (N_23475,N_20579,N_20735);
xor U23476 (N_23476,N_21976,N_22105);
nand U23477 (N_23477,N_21650,N_22015);
nand U23478 (N_23478,N_20207,N_21073);
nand U23479 (N_23479,N_20911,N_20396);
nand U23480 (N_23480,N_21076,N_20130);
nand U23481 (N_23481,N_22176,N_20921);
nand U23482 (N_23482,N_20444,N_22070);
nor U23483 (N_23483,N_21591,N_20500);
or U23484 (N_23484,N_20742,N_20431);
nand U23485 (N_23485,N_21931,N_20140);
and U23486 (N_23486,N_22235,N_21624);
nor U23487 (N_23487,N_20388,N_22195);
or U23488 (N_23488,N_21267,N_20304);
xnor U23489 (N_23489,N_20075,N_20553);
or U23490 (N_23490,N_21888,N_22336);
or U23491 (N_23491,N_21811,N_21299);
xor U23492 (N_23492,N_21354,N_22257);
or U23493 (N_23493,N_21768,N_20098);
nand U23494 (N_23494,N_21585,N_20347);
nand U23495 (N_23495,N_20393,N_20639);
nand U23496 (N_23496,N_22038,N_21127);
xnor U23497 (N_23497,N_21825,N_22317);
nand U23498 (N_23498,N_21380,N_21359);
xor U23499 (N_23499,N_22495,N_20602);
nand U23500 (N_23500,N_20713,N_20779);
and U23501 (N_23501,N_20901,N_21394);
xnor U23502 (N_23502,N_21802,N_20770);
nor U23503 (N_23503,N_20859,N_20147);
nand U23504 (N_23504,N_20892,N_21561);
nand U23505 (N_23505,N_22110,N_22175);
xnor U23506 (N_23506,N_20252,N_20092);
xnor U23507 (N_23507,N_21770,N_21971);
and U23508 (N_23508,N_20727,N_21766);
and U23509 (N_23509,N_20687,N_20231);
nand U23510 (N_23510,N_20068,N_21532);
xor U23511 (N_23511,N_21813,N_21834);
and U23512 (N_23512,N_20512,N_21321);
and U23513 (N_23513,N_21654,N_21016);
or U23514 (N_23514,N_20757,N_21003);
xor U23515 (N_23515,N_22144,N_21273);
nand U23516 (N_23516,N_21614,N_22304);
xnor U23517 (N_23517,N_20966,N_20995);
nand U23518 (N_23518,N_21302,N_20446);
or U23519 (N_23519,N_20660,N_21686);
nand U23520 (N_23520,N_20464,N_22223);
and U23521 (N_23521,N_20308,N_21275);
and U23522 (N_23522,N_20941,N_21344);
nor U23523 (N_23523,N_21505,N_21902);
or U23524 (N_23524,N_21571,N_21870);
xnor U23525 (N_23525,N_20040,N_21607);
nand U23526 (N_23526,N_20181,N_20927);
nand U23527 (N_23527,N_22275,N_21375);
xor U23528 (N_23528,N_22411,N_20031);
and U23529 (N_23529,N_21892,N_21063);
xnor U23530 (N_23530,N_21064,N_21538);
nand U23531 (N_23531,N_21801,N_21415);
nor U23532 (N_23532,N_20416,N_22043);
nor U23533 (N_23533,N_22273,N_21231);
and U23534 (N_23534,N_21217,N_21552);
nand U23535 (N_23535,N_20418,N_21718);
or U23536 (N_23536,N_21589,N_20061);
or U23537 (N_23537,N_21641,N_21739);
or U23538 (N_23538,N_22376,N_21676);
and U23539 (N_23539,N_21876,N_20042);
nand U23540 (N_23540,N_21433,N_20630);
xor U23541 (N_23541,N_22213,N_21437);
nand U23542 (N_23542,N_22264,N_21769);
and U23543 (N_23543,N_20703,N_21067);
xnor U23544 (N_23544,N_21226,N_20814);
nand U23545 (N_23545,N_21705,N_20162);
xnor U23546 (N_23546,N_20914,N_20925);
or U23547 (N_23547,N_20634,N_21330);
and U23548 (N_23548,N_20441,N_20173);
xor U23549 (N_23549,N_22353,N_21356);
or U23550 (N_23550,N_21050,N_21634);
or U23551 (N_23551,N_21348,N_21560);
nor U23552 (N_23552,N_20262,N_20577);
or U23553 (N_23553,N_21136,N_21193);
nor U23554 (N_23554,N_20200,N_22092);
nor U23555 (N_23555,N_20549,N_21428);
nor U23556 (N_23556,N_20324,N_20664);
nand U23557 (N_23557,N_20708,N_20881);
or U23558 (N_23558,N_21960,N_22400);
xor U23559 (N_23559,N_21386,N_20380);
or U23560 (N_23560,N_22243,N_21294);
nand U23561 (N_23561,N_21522,N_21405);
or U23562 (N_23562,N_21709,N_20163);
and U23563 (N_23563,N_20581,N_21785);
xnor U23564 (N_23564,N_21761,N_21950);
xor U23565 (N_23565,N_21839,N_20815);
or U23566 (N_23566,N_21693,N_20413);
xnor U23567 (N_23567,N_20969,N_21875);
or U23568 (N_23568,N_20556,N_20295);
nand U23569 (N_23569,N_21961,N_21263);
nand U23570 (N_23570,N_20316,N_21186);
and U23571 (N_23571,N_21393,N_22229);
or U23572 (N_23572,N_20479,N_21939);
nand U23573 (N_23573,N_20734,N_20180);
nand U23574 (N_23574,N_22339,N_21360);
and U23575 (N_23575,N_21455,N_21744);
nand U23576 (N_23576,N_20586,N_22337);
nor U23577 (N_23577,N_21185,N_22022);
nor U23578 (N_23578,N_22420,N_21179);
xnor U23579 (N_23579,N_20265,N_21008);
and U23580 (N_23580,N_21277,N_21508);
nand U23581 (N_23581,N_21317,N_22227);
or U23582 (N_23582,N_22059,N_22333);
or U23583 (N_23583,N_22024,N_20424);
nand U23584 (N_23584,N_20462,N_22158);
nor U23585 (N_23585,N_21276,N_20632);
or U23586 (N_23586,N_21681,N_20685);
and U23587 (N_23587,N_21752,N_21854);
or U23588 (N_23588,N_20243,N_22056);
xor U23589 (N_23589,N_21736,N_20136);
and U23590 (N_23590,N_22026,N_20060);
and U23591 (N_23591,N_21899,N_22298);
and U23592 (N_23592,N_20333,N_21469);
nor U23593 (N_23593,N_21723,N_21464);
nand U23594 (N_23594,N_22036,N_21553);
xor U23595 (N_23595,N_20034,N_22165);
and U23596 (N_23596,N_20610,N_20274);
nor U23597 (N_23597,N_22236,N_21445);
nor U23598 (N_23598,N_21793,N_22122);
and U23599 (N_23599,N_20764,N_21807);
xor U23600 (N_23600,N_20877,N_20805);
xnor U23601 (N_23601,N_22486,N_21011);
and U23602 (N_23602,N_20801,N_20564);
or U23603 (N_23603,N_21819,N_21024);
nand U23604 (N_23604,N_21904,N_21795);
nor U23605 (N_23605,N_20337,N_22402);
xor U23606 (N_23606,N_20065,N_20526);
nand U23607 (N_23607,N_20716,N_21596);
nand U23608 (N_23608,N_20365,N_21569);
nor U23609 (N_23609,N_21773,N_22410);
and U23610 (N_23610,N_20114,N_21334);
nand U23611 (N_23611,N_21717,N_21153);
or U23612 (N_23612,N_21772,N_21824);
or U23613 (N_23613,N_21626,N_22309);
xnor U23614 (N_23614,N_22196,N_20339);
nand U23615 (N_23615,N_20323,N_20143);
nor U23616 (N_23616,N_20933,N_20699);
and U23617 (N_23617,N_20694,N_20647);
and U23618 (N_23618,N_21018,N_21431);
nor U23619 (N_23619,N_20882,N_21502);
and U23620 (N_23620,N_22000,N_22215);
nand U23621 (N_23621,N_22382,N_20133);
or U23622 (N_23622,N_20402,N_20880);
xor U23623 (N_23623,N_21026,N_22282);
xor U23624 (N_23624,N_21729,N_21396);
xnor U23625 (N_23625,N_20718,N_21881);
or U23626 (N_23626,N_20394,N_20121);
or U23627 (N_23627,N_22131,N_20585);
xor U23628 (N_23628,N_20956,N_21833);
nand U23629 (N_23629,N_22096,N_22399);
xnor U23630 (N_23630,N_22290,N_20244);
and U23631 (N_23631,N_21644,N_20568);
xnor U23632 (N_23632,N_21336,N_22244);
nor U23633 (N_23633,N_21257,N_20148);
nand U23634 (N_23634,N_20505,N_21732);
nor U23635 (N_23635,N_22075,N_21322);
and U23636 (N_23636,N_22027,N_20587);
or U23637 (N_23637,N_20643,N_21057);
nand U23638 (N_23638,N_20974,N_21372);
nand U23639 (N_23639,N_20493,N_21850);
nor U23640 (N_23640,N_21691,N_20235);
nand U23641 (N_23641,N_22143,N_21473);
or U23642 (N_23642,N_20622,N_21104);
xor U23643 (N_23643,N_22338,N_20475);
and U23644 (N_23644,N_21528,N_21347);
or U23645 (N_23645,N_22259,N_22160);
nand U23646 (N_23646,N_21272,N_20909);
xnor U23647 (N_23647,N_20212,N_21668);
nand U23648 (N_23648,N_20291,N_22286);
xor U23649 (N_23649,N_20036,N_21454);
or U23650 (N_23650,N_22108,N_20456);
or U23651 (N_23651,N_22387,N_20457);
or U23652 (N_23652,N_20510,N_22263);
nand U23653 (N_23653,N_20952,N_20064);
and U23654 (N_23654,N_22465,N_22479);
or U23655 (N_23655,N_20345,N_20894);
xnor U23656 (N_23656,N_22081,N_21107);
nand U23657 (N_23657,N_20364,N_20154);
and U23658 (N_23658,N_21368,N_22007);
xnor U23659 (N_23659,N_22292,N_20689);
xnor U23660 (N_23660,N_20835,N_22444);
nand U23661 (N_23661,N_20567,N_21126);
nand U23662 (N_23662,N_21780,N_21967);
xnor U23663 (N_23663,N_20176,N_20360);
xnor U23664 (N_23664,N_21197,N_22167);
nor U23665 (N_23665,N_20191,N_21934);
or U23666 (N_23666,N_20498,N_21047);
or U23667 (N_23667,N_20302,N_21619);
nor U23668 (N_23668,N_21055,N_21826);
xnor U23669 (N_23669,N_21918,N_20266);
xnor U23670 (N_23670,N_20919,N_20981);
xor U23671 (N_23671,N_20887,N_20400);
or U23672 (N_23672,N_22428,N_21087);
xor U23673 (N_23673,N_20923,N_20704);
xor U23674 (N_23674,N_21655,N_20310);
or U23675 (N_23675,N_22294,N_22300);
nor U23676 (N_23676,N_20387,N_21190);
and U23677 (N_23677,N_20951,N_21400);
nand U23678 (N_23678,N_20635,N_20701);
nor U23679 (N_23679,N_20421,N_20792);
xor U23680 (N_23680,N_20766,N_20267);
and U23681 (N_23681,N_20802,N_21432);
xor U23682 (N_23682,N_22319,N_20984);
xnor U23683 (N_23683,N_21212,N_20590);
and U23684 (N_23684,N_20220,N_22177);
nand U23685 (N_23685,N_20832,N_20459);
nor U23686 (N_23686,N_21059,N_20594);
or U23687 (N_23687,N_20593,N_20397);
nor U23688 (N_23688,N_21369,N_22359);
nand U23689 (N_23689,N_20932,N_20980);
nand U23690 (N_23690,N_22494,N_20775);
nand U23691 (N_23691,N_20119,N_20108);
and U23692 (N_23692,N_22396,N_20084);
or U23693 (N_23693,N_20638,N_20370);
nand U23694 (N_23694,N_20536,N_20470);
or U23695 (N_23695,N_22090,N_21965);
and U23696 (N_23696,N_20978,N_20948);
xor U23697 (N_23697,N_20883,N_21025);
nand U23698 (N_23698,N_21792,N_21205);
or U23699 (N_23699,N_22431,N_22225);
and U23700 (N_23700,N_21171,N_20141);
and U23701 (N_23701,N_20275,N_20298);
nand U23702 (N_23702,N_20048,N_20807);
nand U23703 (N_23703,N_20445,N_20375);
xnor U23704 (N_23704,N_20793,N_21776);
or U23705 (N_23705,N_20502,N_22392);
nor U23706 (N_23706,N_22163,N_21167);
xor U23707 (N_23707,N_20746,N_21618);
or U23708 (N_23708,N_20765,N_20550);
xor U23709 (N_23709,N_20849,N_20056);
or U23710 (N_23710,N_20185,N_21861);
xnor U23711 (N_23711,N_20834,N_20055);
and U23712 (N_23712,N_22029,N_20888);
or U23713 (N_23713,N_21512,N_20600);
nor U23714 (N_23714,N_21425,N_20481);
xnor U23715 (N_23715,N_22169,N_22120);
xnor U23716 (N_23716,N_21401,N_21306);
and U23717 (N_23717,N_20209,N_21993);
and U23718 (N_23718,N_21017,N_20847);
or U23719 (N_23719,N_21901,N_20329);
xor U23720 (N_23720,N_21102,N_21363);
or U23721 (N_23721,N_21864,N_21724);
xnor U23722 (N_23722,N_21576,N_21710);
xnor U23723 (N_23723,N_20977,N_21279);
xnor U23724 (N_23724,N_20020,N_21180);
nand U23725 (N_23725,N_20389,N_21687);
nand U23726 (N_23726,N_20078,N_20915);
or U23727 (N_23727,N_22156,N_21385);
xor U23728 (N_23728,N_20692,N_22067);
xnor U23729 (N_23729,N_21783,N_21220);
and U23730 (N_23730,N_21989,N_22058);
and U23731 (N_23731,N_20895,N_21556);
and U23732 (N_23732,N_21524,N_21253);
xor U23733 (N_23733,N_21921,N_21900);
nand U23734 (N_23734,N_21930,N_20531);
nor U23735 (N_23735,N_21586,N_20623);
or U23736 (N_23736,N_21481,N_21730);
nor U23737 (N_23737,N_21166,N_20058);
or U23738 (N_23738,N_21551,N_21799);
and U23739 (N_23739,N_20155,N_20702);
nor U23740 (N_23740,N_20435,N_22224);
nand U23741 (N_23741,N_20836,N_20137);
nand U23742 (N_23742,N_20404,N_22441);
xnor U23743 (N_23743,N_21937,N_22477);
xor U23744 (N_23744,N_21491,N_21885);
xor U23745 (N_23745,N_21891,N_20993);
xnor U23746 (N_23746,N_21702,N_21871);
xnor U23747 (N_23747,N_22107,N_20614);
and U23748 (N_23748,N_22266,N_21951);
nand U23749 (N_23749,N_22148,N_22139);
and U23750 (N_23750,N_21069,N_22319);
or U23751 (N_23751,N_21794,N_20797);
xnor U23752 (N_23752,N_21528,N_21165);
nand U23753 (N_23753,N_20090,N_20540);
nand U23754 (N_23754,N_21047,N_20804);
xor U23755 (N_23755,N_20651,N_21190);
or U23756 (N_23756,N_20336,N_22468);
xnor U23757 (N_23757,N_21045,N_20005);
nand U23758 (N_23758,N_20491,N_21063);
nor U23759 (N_23759,N_21974,N_21302);
and U23760 (N_23760,N_21086,N_22217);
and U23761 (N_23761,N_22068,N_20456);
or U23762 (N_23762,N_20130,N_21662);
nor U23763 (N_23763,N_22146,N_22335);
and U23764 (N_23764,N_20753,N_22309);
nor U23765 (N_23765,N_21140,N_22456);
nor U23766 (N_23766,N_21945,N_20764);
nand U23767 (N_23767,N_22175,N_20200);
nand U23768 (N_23768,N_20085,N_21753);
nor U23769 (N_23769,N_20352,N_21832);
xor U23770 (N_23770,N_22369,N_22317);
nand U23771 (N_23771,N_20447,N_21540);
and U23772 (N_23772,N_20610,N_21388);
or U23773 (N_23773,N_20172,N_20915);
or U23774 (N_23774,N_21840,N_21094);
and U23775 (N_23775,N_20430,N_22495);
nand U23776 (N_23776,N_22426,N_20011);
nor U23777 (N_23777,N_20550,N_21900);
and U23778 (N_23778,N_20832,N_21319);
nand U23779 (N_23779,N_20088,N_20140);
xor U23780 (N_23780,N_20495,N_21165);
xnor U23781 (N_23781,N_21997,N_20699);
nor U23782 (N_23782,N_22387,N_20273);
or U23783 (N_23783,N_20127,N_22398);
nor U23784 (N_23784,N_22423,N_20652);
or U23785 (N_23785,N_21114,N_22466);
nand U23786 (N_23786,N_20899,N_22147);
or U23787 (N_23787,N_20715,N_22106);
nand U23788 (N_23788,N_21862,N_20693);
or U23789 (N_23789,N_22206,N_20300);
and U23790 (N_23790,N_20340,N_21314);
nor U23791 (N_23791,N_22040,N_20702);
nand U23792 (N_23792,N_20187,N_22499);
nand U23793 (N_23793,N_21906,N_20403);
nor U23794 (N_23794,N_20829,N_22445);
and U23795 (N_23795,N_21041,N_20436);
and U23796 (N_23796,N_21737,N_22442);
and U23797 (N_23797,N_20377,N_21137);
xor U23798 (N_23798,N_22055,N_22314);
xor U23799 (N_23799,N_22226,N_20346);
nor U23800 (N_23800,N_21028,N_20927);
and U23801 (N_23801,N_20415,N_22329);
nand U23802 (N_23802,N_20615,N_21181);
xnor U23803 (N_23803,N_22391,N_21653);
and U23804 (N_23804,N_21088,N_21105);
or U23805 (N_23805,N_20308,N_21863);
nand U23806 (N_23806,N_20226,N_20476);
nor U23807 (N_23807,N_20835,N_22086);
xnor U23808 (N_23808,N_20137,N_20501);
and U23809 (N_23809,N_21604,N_20549);
nor U23810 (N_23810,N_22081,N_21451);
nand U23811 (N_23811,N_21729,N_20315);
nor U23812 (N_23812,N_20605,N_22493);
nor U23813 (N_23813,N_20893,N_20414);
nand U23814 (N_23814,N_21419,N_21696);
nor U23815 (N_23815,N_21865,N_21004);
nand U23816 (N_23816,N_21487,N_20984);
nor U23817 (N_23817,N_20722,N_20078);
nor U23818 (N_23818,N_21470,N_20334);
nand U23819 (N_23819,N_21872,N_20861);
and U23820 (N_23820,N_21916,N_21257);
and U23821 (N_23821,N_20868,N_21274);
xor U23822 (N_23822,N_21192,N_22211);
xor U23823 (N_23823,N_21916,N_20225);
nand U23824 (N_23824,N_22276,N_20947);
or U23825 (N_23825,N_20706,N_20624);
nand U23826 (N_23826,N_22206,N_21603);
or U23827 (N_23827,N_20778,N_21682);
nor U23828 (N_23828,N_20246,N_22041);
nor U23829 (N_23829,N_21606,N_21760);
nor U23830 (N_23830,N_20132,N_20834);
or U23831 (N_23831,N_20975,N_21408);
or U23832 (N_23832,N_22383,N_21972);
xnor U23833 (N_23833,N_20686,N_21580);
or U23834 (N_23834,N_21019,N_21924);
or U23835 (N_23835,N_21420,N_21121);
xnor U23836 (N_23836,N_20745,N_22217);
and U23837 (N_23837,N_20277,N_21111);
or U23838 (N_23838,N_20077,N_21498);
or U23839 (N_23839,N_21887,N_20608);
nor U23840 (N_23840,N_20240,N_20024);
nor U23841 (N_23841,N_21948,N_22176);
or U23842 (N_23842,N_20971,N_21412);
and U23843 (N_23843,N_21923,N_20864);
xor U23844 (N_23844,N_20057,N_20424);
xnor U23845 (N_23845,N_21851,N_21289);
xnor U23846 (N_23846,N_22161,N_22353);
or U23847 (N_23847,N_21089,N_20922);
and U23848 (N_23848,N_20236,N_22321);
nand U23849 (N_23849,N_22276,N_22284);
xor U23850 (N_23850,N_20683,N_21301);
and U23851 (N_23851,N_20227,N_20984);
nor U23852 (N_23852,N_22287,N_20498);
nor U23853 (N_23853,N_21628,N_20963);
nand U23854 (N_23854,N_21807,N_22090);
nand U23855 (N_23855,N_20562,N_20563);
nor U23856 (N_23856,N_21937,N_22465);
nand U23857 (N_23857,N_22218,N_22479);
or U23858 (N_23858,N_22142,N_21239);
and U23859 (N_23859,N_20564,N_21043);
nand U23860 (N_23860,N_21012,N_21977);
nor U23861 (N_23861,N_21450,N_22473);
xor U23862 (N_23862,N_20366,N_21585);
xor U23863 (N_23863,N_21982,N_20533);
nand U23864 (N_23864,N_21637,N_21861);
or U23865 (N_23865,N_21446,N_20245);
nand U23866 (N_23866,N_22332,N_20128);
xnor U23867 (N_23867,N_20819,N_20132);
nor U23868 (N_23868,N_20501,N_21168);
nand U23869 (N_23869,N_20113,N_20539);
nand U23870 (N_23870,N_22268,N_22499);
and U23871 (N_23871,N_20411,N_20750);
nor U23872 (N_23872,N_21452,N_20285);
or U23873 (N_23873,N_22282,N_22098);
or U23874 (N_23874,N_20371,N_21069);
and U23875 (N_23875,N_20278,N_22076);
nor U23876 (N_23876,N_21759,N_20354);
nand U23877 (N_23877,N_21669,N_21865);
xor U23878 (N_23878,N_21266,N_22414);
nand U23879 (N_23879,N_22113,N_20337);
or U23880 (N_23880,N_20136,N_20880);
xor U23881 (N_23881,N_20933,N_20428);
or U23882 (N_23882,N_21880,N_21610);
xnor U23883 (N_23883,N_20300,N_20614);
or U23884 (N_23884,N_20159,N_21380);
and U23885 (N_23885,N_22095,N_21708);
and U23886 (N_23886,N_21776,N_21273);
nand U23887 (N_23887,N_20465,N_21085);
or U23888 (N_23888,N_21750,N_20731);
or U23889 (N_23889,N_20874,N_20011);
and U23890 (N_23890,N_20730,N_20091);
and U23891 (N_23891,N_22064,N_22222);
xnor U23892 (N_23892,N_21781,N_20964);
nor U23893 (N_23893,N_20955,N_22253);
nor U23894 (N_23894,N_22443,N_21257);
or U23895 (N_23895,N_21139,N_21572);
xnor U23896 (N_23896,N_21710,N_21893);
and U23897 (N_23897,N_21625,N_21432);
nor U23898 (N_23898,N_21468,N_21001);
and U23899 (N_23899,N_20836,N_21885);
xnor U23900 (N_23900,N_20349,N_22347);
nand U23901 (N_23901,N_21066,N_21697);
or U23902 (N_23902,N_21884,N_22327);
nor U23903 (N_23903,N_21594,N_21219);
or U23904 (N_23904,N_20372,N_21576);
or U23905 (N_23905,N_20484,N_21680);
nor U23906 (N_23906,N_20992,N_20453);
and U23907 (N_23907,N_21682,N_20505);
or U23908 (N_23908,N_21867,N_22221);
and U23909 (N_23909,N_21185,N_20192);
xnor U23910 (N_23910,N_20058,N_20275);
nand U23911 (N_23911,N_20051,N_20216);
nand U23912 (N_23912,N_21287,N_21337);
nor U23913 (N_23913,N_20560,N_22236);
nand U23914 (N_23914,N_20129,N_22157);
and U23915 (N_23915,N_21297,N_22095);
xnor U23916 (N_23916,N_20754,N_21492);
and U23917 (N_23917,N_20645,N_20232);
xnor U23918 (N_23918,N_22055,N_20655);
xor U23919 (N_23919,N_21693,N_20548);
xor U23920 (N_23920,N_21547,N_22120);
or U23921 (N_23921,N_22008,N_22488);
nor U23922 (N_23922,N_21668,N_20549);
and U23923 (N_23923,N_21975,N_21990);
nor U23924 (N_23924,N_21141,N_22142);
nor U23925 (N_23925,N_22021,N_20035);
xnor U23926 (N_23926,N_21263,N_22036);
or U23927 (N_23927,N_21488,N_22117);
nor U23928 (N_23928,N_21161,N_22479);
and U23929 (N_23929,N_21858,N_21387);
and U23930 (N_23930,N_21232,N_21892);
or U23931 (N_23931,N_20623,N_20246);
nor U23932 (N_23932,N_20841,N_21358);
xor U23933 (N_23933,N_20241,N_21837);
nor U23934 (N_23934,N_21729,N_20747);
nand U23935 (N_23935,N_21053,N_20510);
or U23936 (N_23936,N_22118,N_22443);
xor U23937 (N_23937,N_20784,N_22285);
xnor U23938 (N_23938,N_20162,N_21905);
nor U23939 (N_23939,N_20142,N_22315);
xor U23940 (N_23940,N_21493,N_21009);
xor U23941 (N_23941,N_21532,N_21474);
nand U23942 (N_23942,N_20271,N_22198);
or U23943 (N_23943,N_21615,N_20915);
nand U23944 (N_23944,N_20582,N_21468);
and U23945 (N_23945,N_21325,N_20494);
and U23946 (N_23946,N_20261,N_20646);
nor U23947 (N_23947,N_20523,N_21080);
nand U23948 (N_23948,N_22377,N_21919);
or U23949 (N_23949,N_21314,N_21958);
xor U23950 (N_23950,N_21527,N_21341);
and U23951 (N_23951,N_22271,N_21249);
nand U23952 (N_23952,N_20765,N_20304);
and U23953 (N_23953,N_20733,N_20023);
and U23954 (N_23954,N_22411,N_22173);
or U23955 (N_23955,N_21049,N_20597);
xor U23956 (N_23956,N_20642,N_20501);
or U23957 (N_23957,N_20427,N_20013);
nand U23958 (N_23958,N_20559,N_20364);
nor U23959 (N_23959,N_20324,N_21757);
and U23960 (N_23960,N_20286,N_21180);
nand U23961 (N_23961,N_20825,N_21764);
and U23962 (N_23962,N_21179,N_20112);
nor U23963 (N_23963,N_20682,N_22428);
nand U23964 (N_23964,N_21126,N_20840);
or U23965 (N_23965,N_21053,N_22259);
nand U23966 (N_23966,N_20156,N_20836);
xor U23967 (N_23967,N_21776,N_21769);
xor U23968 (N_23968,N_20866,N_20650);
xor U23969 (N_23969,N_22275,N_22406);
nand U23970 (N_23970,N_21575,N_22161);
xnor U23971 (N_23971,N_20383,N_21248);
xor U23972 (N_23972,N_22207,N_21629);
xnor U23973 (N_23973,N_20978,N_22320);
xor U23974 (N_23974,N_21641,N_22306);
nor U23975 (N_23975,N_20659,N_20460);
and U23976 (N_23976,N_20706,N_20547);
or U23977 (N_23977,N_20051,N_22232);
and U23978 (N_23978,N_21462,N_21100);
or U23979 (N_23979,N_21506,N_20110);
or U23980 (N_23980,N_22249,N_20411);
or U23981 (N_23981,N_21279,N_21331);
and U23982 (N_23982,N_20491,N_20627);
xnor U23983 (N_23983,N_21792,N_21870);
xor U23984 (N_23984,N_21147,N_21745);
and U23985 (N_23985,N_20447,N_20615);
xor U23986 (N_23986,N_21483,N_20455);
nand U23987 (N_23987,N_22063,N_22052);
or U23988 (N_23988,N_20946,N_21381);
xor U23989 (N_23989,N_20791,N_20515);
and U23990 (N_23990,N_20812,N_20397);
or U23991 (N_23991,N_20371,N_22315);
nor U23992 (N_23992,N_20710,N_21745);
and U23993 (N_23993,N_20537,N_21387);
nor U23994 (N_23994,N_21192,N_22217);
and U23995 (N_23995,N_21355,N_21434);
and U23996 (N_23996,N_20898,N_21058);
nor U23997 (N_23997,N_22286,N_20139);
and U23998 (N_23998,N_21317,N_20365);
or U23999 (N_23999,N_22235,N_20979);
or U24000 (N_24000,N_20817,N_20708);
xnor U24001 (N_24001,N_21898,N_21471);
and U24002 (N_24002,N_20722,N_21974);
and U24003 (N_24003,N_21220,N_20082);
and U24004 (N_24004,N_22161,N_21678);
nor U24005 (N_24005,N_21892,N_20346);
xor U24006 (N_24006,N_20544,N_20755);
or U24007 (N_24007,N_21354,N_21419);
and U24008 (N_24008,N_22140,N_21045);
nand U24009 (N_24009,N_21753,N_20277);
or U24010 (N_24010,N_22374,N_21349);
nor U24011 (N_24011,N_21205,N_20593);
nand U24012 (N_24012,N_21901,N_21204);
xnor U24013 (N_24013,N_20302,N_21336);
xnor U24014 (N_24014,N_20084,N_20604);
nand U24015 (N_24015,N_22465,N_20583);
nand U24016 (N_24016,N_21495,N_20992);
and U24017 (N_24017,N_21015,N_21420);
and U24018 (N_24018,N_21362,N_22191);
xnor U24019 (N_24019,N_21693,N_22246);
or U24020 (N_24020,N_20316,N_20294);
and U24021 (N_24021,N_21343,N_20054);
or U24022 (N_24022,N_21540,N_21410);
nand U24023 (N_24023,N_22287,N_20162);
and U24024 (N_24024,N_20308,N_22063);
nor U24025 (N_24025,N_21581,N_20467);
and U24026 (N_24026,N_20809,N_21075);
and U24027 (N_24027,N_20718,N_21414);
or U24028 (N_24028,N_20832,N_22173);
and U24029 (N_24029,N_20846,N_22288);
xnor U24030 (N_24030,N_21202,N_21192);
or U24031 (N_24031,N_20831,N_20896);
nor U24032 (N_24032,N_21302,N_20589);
nor U24033 (N_24033,N_22310,N_20845);
and U24034 (N_24034,N_20317,N_20403);
and U24035 (N_24035,N_21962,N_22488);
nor U24036 (N_24036,N_21502,N_20488);
nand U24037 (N_24037,N_22467,N_21721);
xnor U24038 (N_24038,N_20835,N_22036);
or U24039 (N_24039,N_21493,N_20876);
xor U24040 (N_24040,N_20513,N_20085);
xor U24041 (N_24041,N_20826,N_20595);
nor U24042 (N_24042,N_22183,N_21649);
nor U24043 (N_24043,N_22116,N_21219);
nor U24044 (N_24044,N_20882,N_22005);
nand U24045 (N_24045,N_21324,N_20389);
xnor U24046 (N_24046,N_20827,N_21104);
nand U24047 (N_24047,N_20386,N_22473);
nand U24048 (N_24048,N_21952,N_22400);
xnor U24049 (N_24049,N_20962,N_20683);
nor U24050 (N_24050,N_22390,N_20969);
nor U24051 (N_24051,N_21032,N_20445);
or U24052 (N_24052,N_22017,N_20066);
xnor U24053 (N_24053,N_20278,N_21440);
xor U24054 (N_24054,N_21230,N_20012);
nor U24055 (N_24055,N_21817,N_21152);
and U24056 (N_24056,N_20952,N_20052);
or U24057 (N_24057,N_21253,N_21079);
xor U24058 (N_24058,N_21177,N_20499);
nor U24059 (N_24059,N_21433,N_20664);
or U24060 (N_24060,N_20737,N_21066);
or U24061 (N_24061,N_20440,N_20799);
nand U24062 (N_24062,N_20254,N_20405);
or U24063 (N_24063,N_21016,N_22055);
or U24064 (N_24064,N_20153,N_22006);
nor U24065 (N_24065,N_20831,N_20030);
or U24066 (N_24066,N_21394,N_21658);
xnor U24067 (N_24067,N_21632,N_21600);
nand U24068 (N_24068,N_21465,N_20879);
or U24069 (N_24069,N_20041,N_21445);
and U24070 (N_24070,N_20184,N_22169);
and U24071 (N_24071,N_21875,N_20981);
nor U24072 (N_24072,N_21380,N_20481);
xor U24073 (N_24073,N_21548,N_21907);
nor U24074 (N_24074,N_20485,N_22475);
xor U24075 (N_24075,N_21971,N_21293);
xnor U24076 (N_24076,N_20892,N_21107);
or U24077 (N_24077,N_21215,N_21312);
nand U24078 (N_24078,N_20444,N_20941);
nand U24079 (N_24079,N_20293,N_21813);
xor U24080 (N_24080,N_21563,N_21013);
and U24081 (N_24081,N_22354,N_20810);
or U24082 (N_24082,N_20907,N_20673);
nor U24083 (N_24083,N_21218,N_21597);
or U24084 (N_24084,N_20677,N_21119);
nor U24085 (N_24085,N_22203,N_20050);
or U24086 (N_24086,N_21681,N_20039);
xnor U24087 (N_24087,N_21872,N_21210);
or U24088 (N_24088,N_22218,N_20291);
nand U24089 (N_24089,N_20033,N_22282);
nand U24090 (N_24090,N_22152,N_21571);
xnor U24091 (N_24091,N_20017,N_22027);
or U24092 (N_24092,N_20343,N_20768);
and U24093 (N_24093,N_20734,N_20882);
or U24094 (N_24094,N_20752,N_20921);
or U24095 (N_24095,N_20631,N_21399);
nor U24096 (N_24096,N_20334,N_21686);
and U24097 (N_24097,N_20538,N_21815);
and U24098 (N_24098,N_22166,N_21052);
nor U24099 (N_24099,N_20119,N_21232);
nand U24100 (N_24100,N_20544,N_20232);
nand U24101 (N_24101,N_21266,N_20439);
nand U24102 (N_24102,N_20614,N_20266);
nor U24103 (N_24103,N_22270,N_20965);
xor U24104 (N_24104,N_20303,N_22436);
and U24105 (N_24105,N_21086,N_21688);
nor U24106 (N_24106,N_21563,N_20369);
nor U24107 (N_24107,N_21777,N_20139);
nand U24108 (N_24108,N_22006,N_20483);
nor U24109 (N_24109,N_20418,N_21676);
xor U24110 (N_24110,N_20542,N_20628);
and U24111 (N_24111,N_22383,N_21287);
or U24112 (N_24112,N_21535,N_22281);
or U24113 (N_24113,N_22060,N_20248);
nor U24114 (N_24114,N_21885,N_22292);
nor U24115 (N_24115,N_21032,N_21015);
or U24116 (N_24116,N_22428,N_20777);
nand U24117 (N_24117,N_20076,N_21315);
xnor U24118 (N_24118,N_20411,N_20403);
nand U24119 (N_24119,N_20481,N_22104);
xnor U24120 (N_24120,N_20607,N_20452);
nor U24121 (N_24121,N_22344,N_21592);
nor U24122 (N_24122,N_21452,N_20691);
nand U24123 (N_24123,N_22265,N_21665);
nand U24124 (N_24124,N_21963,N_21049);
nand U24125 (N_24125,N_21382,N_21833);
nand U24126 (N_24126,N_21502,N_20732);
or U24127 (N_24127,N_20111,N_21953);
and U24128 (N_24128,N_21029,N_22258);
or U24129 (N_24129,N_22021,N_21733);
nand U24130 (N_24130,N_21823,N_21980);
and U24131 (N_24131,N_20342,N_21352);
and U24132 (N_24132,N_20161,N_21919);
xor U24133 (N_24133,N_20348,N_20403);
xnor U24134 (N_24134,N_20812,N_20882);
nand U24135 (N_24135,N_21388,N_20799);
and U24136 (N_24136,N_21191,N_21830);
or U24137 (N_24137,N_20075,N_20259);
or U24138 (N_24138,N_21055,N_20103);
nand U24139 (N_24139,N_20519,N_22050);
nor U24140 (N_24140,N_20797,N_20784);
nand U24141 (N_24141,N_22035,N_22093);
nand U24142 (N_24142,N_22249,N_20342);
xnor U24143 (N_24143,N_21608,N_20028);
xnor U24144 (N_24144,N_20234,N_21033);
nor U24145 (N_24145,N_20675,N_20035);
nand U24146 (N_24146,N_20911,N_22447);
nand U24147 (N_24147,N_20925,N_21562);
xor U24148 (N_24148,N_20325,N_21989);
xor U24149 (N_24149,N_20823,N_21227);
xor U24150 (N_24150,N_22007,N_21591);
xnor U24151 (N_24151,N_20091,N_20813);
nor U24152 (N_24152,N_21331,N_21814);
or U24153 (N_24153,N_21106,N_20580);
and U24154 (N_24154,N_22290,N_21186);
or U24155 (N_24155,N_21434,N_20110);
nor U24156 (N_24156,N_21045,N_20356);
and U24157 (N_24157,N_21527,N_20503);
or U24158 (N_24158,N_22423,N_21322);
nand U24159 (N_24159,N_20158,N_21325);
nand U24160 (N_24160,N_21618,N_22252);
and U24161 (N_24161,N_22045,N_21410);
nor U24162 (N_24162,N_20934,N_20666);
or U24163 (N_24163,N_21717,N_21942);
nor U24164 (N_24164,N_20712,N_21353);
xor U24165 (N_24165,N_21693,N_21841);
xnor U24166 (N_24166,N_20470,N_22034);
xor U24167 (N_24167,N_21835,N_20398);
nand U24168 (N_24168,N_20118,N_21582);
and U24169 (N_24169,N_22159,N_20413);
nand U24170 (N_24170,N_22436,N_20504);
xnor U24171 (N_24171,N_21550,N_20949);
and U24172 (N_24172,N_21374,N_20356);
xor U24173 (N_24173,N_22162,N_22290);
nor U24174 (N_24174,N_20460,N_20550);
or U24175 (N_24175,N_21994,N_21740);
xnor U24176 (N_24176,N_21660,N_20475);
and U24177 (N_24177,N_20265,N_20315);
and U24178 (N_24178,N_21366,N_21062);
nand U24179 (N_24179,N_20558,N_20178);
xnor U24180 (N_24180,N_21560,N_21671);
and U24181 (N_24181,N_21386,N_21309);
nand U24182 (N_24182,N_21271,N_22287);
nor U24183 (N_24183,N_22306,N_22488);
or U24184 (N_24184,N_22018,N_21770);
and U24185 (N_24185,N_21687,N_21166);
nand U24186 (N_24186,N_21160,N_22272);
and U24187 (N_24187,N_22401,N_22364);
and U24188 (N_24188,N_21189,N_21814);
and U24189 (N_24189,N_21388,N_20997);
xor U24190 (N_24190,N_21428,N_20809);
nand U24191 (N_24191,N_20599,N_21367);
or U24192 (N_24192,N_20744,N_22433);
and U24193 (N_24193,N_21792,N_21453);
xor U24194 (N_24194,N_20818,N_21573);
or U24195 (N_24195,N_22155,N_20832);
and U24196 (N_24196,N_22246,N_21008);
nor U24197 (N_24197,N_21063,N_20210);
and U24198 (N_24198,N_20755,N_22059);
or U24199 (N_24199,N_21480,N_21093);
or U24200 (N_24200,N_22442,N_21879);
xnor U24201 (N_24201,N_20505,N_20029);
and U24202 (N_24202,N_21584,N_20502);
xnor U24203 (N_24203,N_21878,N_21460);
nor U24204 (N_24204,N_22127,N_21987);
or U24205 (N_24205,N_21188,N_21218);
or U24206 (N_24206,N_21034,N_21952);
or U24207 (N_24207,N_20902,N_21914);
or U24208 (N_24208,N_20691,N_20267);
xnor U24209 (N_24209,N_20965,N_21688);
or U24210 (N_24210,N_22099,N_20608);
nor U24211 (N_24211,N_20487,N_20717);
nor U24212 (N_24212,N_22006,N_20085);
and U24213 (N_24213,N_20447,N_22469);
nor U24214 (N_24214,N_22371,N_21000);
nor U24215 (N_24215,N_22156,N_21374);
and U24216 (N_24216,N_22136,N_20521);
or U24217 (N_24217,N_20771,N_20318);
or U24218 (N_24218,N_20758,N_21928);
nor U24219 (N_24219,N_20883,N_21220);
and U24220 (N_24220,N_22098,N_20107);
or U24221 (N_24221,N_21879,N_21011);
or U24222 (N_24222,N_20512,N_21223);
nand U24223 (N_24223,N_21188,N_21306);
xnor U24224 (N_24224,N_22204,N_20879);
and U24225 (N_24225,N_22031,N_21773);
xor U24226 (N_24226,N_21837,N_21127);
or U24227 (N_24227,N_21604,N_21241);
nor U24228 (N_24228,N_22315,N_22050);
and U24229 (N_24229,N_20654,N_21854);
or U24230 (N_24230,N_22269,N_21261);
and U24231 (N_24231,N_20087,N_20321);
and U24232 (N_24232,N_20268,N_22076);
nand U24233 (N_24233,N_22450,N_21558);
xnor U24234 (N_24234,N_21786,N_20807);
xnor U24235 (N_24235,N_21464,N_21215);
and U24236 (N_24236,N_21122,N_22337);
or U24237 (N_24237,N_20771,N_22398);
xor U24238 (N_24238,N_20092,N_20559);
nand U24239 (N_24239,N_21281,N_21704);
nor U24240 (N_24240,N_21565,N_21856);
xor U24241 (N_24241,N_22280,N_21868);
xor U24242 (N_24242,N_22042,N_22277);
nor U24243 (N_24243,N_22478,N_21252);
xor U24244 (N_24244,N_20792,N_20994);
and U24245 (N_24245,N_21929,N_22318);
and U24246 (N_24246,N_20644,N_20193);
xor U24247 (N_24247,N_20819,N_21692);
nand U24248 (N_24248,N_21745,N_22477);
nand U24249 (N_24249,N_21107,N_20227);
and U24250 (N_24250,N_22358,N_20922);
and U24251 (N_24251,N_20120,N_20746);
nand U24252 (N_24252,N_21878,N_20070);
xor U24253 (N_24253,N_22279,N_20277);
or U24254 (N_24254,N_22153,N_20250);
or U24255 (N_24255,N_20267,N_21795);
xor U24256 (N_24256,N_21153,N_22156);
nand U24257 (N_24257,N_21316,N_20992);
xor U24258 (N_24258,N_20504,N_21129);
or U24259 (N_24259,N_22399,N_20503);
or U24260 (N_24260,N_20499,N_21642);
nand U24261 (N_24261,N_21583,N_20630);
or U24262 (N_24262,N_20648,N_21571);
xor U24263 (N_24263,N_20586,N_22219);
xor U24264 (N_24264,N_20566,N_21511);
xor U24265 (N_24265,N_20793,N_20664);
nor U24266 (N_24266,N_22065,N_21299);
or U24267 (N_24267,N_20932,N_20626);
nor U24268 (N_24268,N_20096,N_20668);
xor U24269 (N_24269,N_22330,N_21590);
and U24270 (N_24270,N_20325,N_21779);
nor U24271 (N_24271,N_21714,N_20498);
or U24272 (N_24272,N_20360,N_20001);
and U24273 (N_24273,N_20194,N_20565);
nand U24274 (N_24274,N_21441,N_22240);
nand U24275 (N_24275,N_20521,N_20427);
xor U24276 (N_24276,N_20928,N_21448);
and U24277 (N_24277,N_21608,N_20850);
and U24278 (N_24278,N_21311,N_20455);
or U24279 (N_24279,N_20145,N_22118);
nand U24280 (N_24280,N_20058,N_20277);
and U24281 (N_24281,N_22090,N_21272);
or U24282 (N_24282,N_21930,N_20459);
nand U24283 (N_24283,N_21010,N_21764);
nor U24284 (N_24284,N_20945,N_20080);
and U24285 (N_24285,N_20736,N_22445);
nand U24286 (N_24286,N_21064,N_20425);
and U24287 (N_24287,N_20509,N_21533);
nor U24288 (N_24288,N_21077,N_22056);
nand U24289 (N_24289,N_20527,N_22469);
xnor U24290 (N_24290,N_22027,N_20379);
and U24291 (N_24291,N_21479,N_20382);
xnor U24292 (N_24292,N_20957,N_20320);
or U24293 (N_24293,N_20914,N_21546);
nor U24294 (N_24294,N_22192,N_21153);
nor U24295 (N_24295,N_21143,N_21215);
and U24296 (N_24296,N_22456,N_21669);
or U24297 (N_24297,N_21767,N_22065);
and U24298 (N_24298,N_20284,N_20490);
nand U24299 (N_24299,N_20827,N_20481);
nor U24300 (N_24300,N_22239,N_22076);
nand U24301 (N_24301,N_21329,N_20401);
and U24302 (N_24302,N_20937,N_20825);
nor U24303 (N_24303,N_20429,N_20419);
nor U24304 (N_24304,N_20017,N_20899);
and U24305 (N_24305,N_20882,N_22098);
nor U24306 (N_24306,N_22221,N_20920);
and U24307 (N_24307,N_20129,N_21161);
nor U24308 (N_24308,N_21061,N_21396);
nand U24309 (N_24309,N_21969,N_20255);
nor U24310 (N_24310,N_20347,N_20133);
xnor U24311 (N_24311,N_22256,N_20730);
nor U24312 (N_24312,N_21450,N_22418);
nand U24313 (N_24313,N_20023,N_22247);
and U24314 (N_24314,N_21751,N_22047);
nand U24315 (N_24315,N_21438,N_21556);
nand U24316 (N_24316,N_21424,N_20093);
nor U24317 (N_24317,N_21659,N_20291);
nor U24318 (N_24318,N_20230,N_20217);
or U24319 (N_24319,N_20704,N_22084);
xnor U24320 (N_24320,N_21646,N_22006);
or U24321 (N_24321,N_22211,N_20516);
nor U24322 (N_24322,N_20369,N_21164);
nand U24323 (N_24323,N_21953,N_21160);
nor U24324 (N_24324,N_22073,N_20093);
nor U24325 (N_24325,N_20106,N_22444);
nor U24326 (N_24326,N_20468,N_21845);
nor U24327 (N_24327,N_21715,N_20066);
xor U24328 (N_24328,N_20577,N_21029);
nor U24329 (N_24329,N_21934,N_22188);
and U24330 (N_24330,N_21492,N_21104);
nand U24331 (N_24331,N_22197,N_21126);
xnor U24332 (N_24332,N_20028,N_20258);
nand U24333 (N_24333,N_20819,N_20776);
xor U24334 (N_24334,N_21294,N_22382);
xnor U24335 (N_24335,N_20952,N_22300);
xor U24336 (N_24336,N_21474,N_21407);
xnor U24337 (N_24337,N_21347,N_21318);
nor U24338 (N_24338,N_21170,N_20570);
nand U24339 (N_24339,N_22436,N_20485);
xor U24340 (N_24340,N_22148,N_22271);
or U24341 (N_24341,N_20371,N_20303);
and U24342 (N_24342,N_22068,N_20985);
or U24343 (N_24343,N_22315,N_20467);
nor U24344 (N_24344,N_22325,N_22235);
or U24345 (N_24345,N_21670,N_20990);
nand U24346 (N_24346,N_21306,N_20125);
xnor U24347 (N_24347,N_22215,N_21130);
or U24348 (N_24348,N_20394,N_22276);
xnor U24349 (N_24349,N_21481,N_22021);
or U24350 (N_24350,N_21004,N_20186);
or U24351 (N_24351,N_20124,N_21877);
or U24352 (N_24352,N_22127,N_20391);
nor U24353 (N_24353,N_20725,N_20692);
or U24354 (N_24354,N_20503,N_20085);
or U24355 (N_24355,N_20852,N_22014);
xnor U24356 (N_24356,N_21155,N_21643);
nor U24357 (N_24357,N_21733,N_20034);
nor U24358 (N_24358,N_21599,N_21002);
nand U24359 (N_24359,N_21615,N_20944);
xnor U24360 (N_24360,N_21827,N_21616);
or U24361 (N_24361,N_21243,N_20787);
nor U24362 (N_24362,N_20646,N_20218);
nor U24363 (N_24363,N_21176,N_20834);
or U24364 (N_24364,N_20461,N_20276);
and U24365 (N_24365,N_21390,N_20413);
nor U24366 (N_24366,N_22049,N_21621);
or U24367 (N_24367,N_21542,N_21402);
or U24368 (N_24368,N_20739,N_20633);
or U24369 (N_24369,N_21064,N_22399);
and U24370 (N_24370,N_21262,N_20094);
and U24371 (N_24371,N_20660,N_20239);
and U24372 (N_24372,N_20160,N_20433);
xnor U24373 (N_24373,N_21623,N_21646);
nand U24374 (N_24374,N_21473,N_20274);
xnor U24375 (N_24375,N_21742,N_20394);
and U24376 (N_24376,N_22225,N_21218);
or U24377 (N_24377,N_21518,N_22473);
xnor U24378 (N_24378,N_20014,N_20802);
nand U24379 (N_24379,N_20840,N_21393);
and U24380 (N_24380,N_20437,N_21837);
xor U24381 (N_24381,N_21400,N_22382);
nor U24382 (N_24382,N_21450,N_20754);
or U24383 (N_24383,N_22185,N_21879);
nor U24384 (N_24384,N_20103,N_21790);
xor U24385 (N_24385,N_20418,N_21415);
nand U24386 (N_24386,N_22325,N_21860);
nor U24387 (N_24387,N_22432,N_21548);
nand U24388 (N_24388,N_21746,N_20408);
nand U24389 (N_24389,N_20692,N_21658);
or U24390 (N_24390,N_21963,N_20157);
nor U24391 (N_24391,N_22164,N_21620);
xor U24392 (N_24392,N_21382,N_22464);
xnor U24393 (N_24393,N_22127,N_21157);
and U24394 (N_24394,N_20143,N_21200);
nand U24395 (N_24395,N_20699,N_21422);
nor U24396 (N_24396,N_21389,N_22042);
or U24397 (N_24397,N_21021,N_20222);
nor U24398 (N_24398,N_22159,N_21553);
nor U24399 (N_24399,N_21839,N_21057);
and U24400 (N_24400,N_21848,N_21979);
or U24401 (N_24401,N_21329,N_20768);
nand U24402 (N_24402,N_20705,N_20812);
or U24403 (N_24403,N_21826,N_21460);
or U24404 (N_24404,N_21053,N_20840);
xnor U24405 (N_24405,N_21516,N_21263);
or U24406 (N_24406,N_21590,N_20630);
nor U24407 (N_24407,N_22287,N_21456);
xnor U24408 (N_24408,N_20968,N_20139);
or U24409 (N_24409,N_20334,N_21292);
xnor U24410 (N_24410,N_22220,N_22178);
and U24411 (N_24411,N_21960,N_21127);
or U24412 (N_24412,N_22236,N_21017);
and U24413 (N_24413,N_20315,N_21184);
and U24414 (N_24414,N_21252,N_21698);
xnor U24415 (N_24415,N_20676,N_21717);
and U24416 (N_24416,N_21652,N_21473);
nor U24417 (N_24417,N_21837,N_22031);
xor U24418 (N_24418,N_21751,N_20566);
nor U24419 (N_24419,N_20261,N_21979);
xor U24420 (N_24420,N_21079,N_22326);
or U24421 (N_24421,N_22286,N_22211);
nor U24422 (N_24422,N_22493,N_20637);
and U24423 (N_24423,N_20366,N_21531);
or U24424 (N_24424,N_22434,N_21511);
xor U24425 (N_24425,N_20729,N_20517);
nor U24426 (N_24426,N_21052,N_21083);
nand U24427 (N_24427,N_20358,N_20235);
and U24428 (N_24428,N_21297,N_21954);
or U24429 (N_24429,N_20648,N_21566);
xor U24430 (N_24430,N_20242,N_20477);
nor U24431 (N_24431,N_22218,N_20409);
xnor U24432 (N_24432,N_20627,N_20255);
xor U24433 (N_24433,N_20765,N_20115);
nand U24434 (N_24434,N_21590,N_21591);
nand U24435 (N_24435,N_20174,N_21195);
nor U24436 (N_24436,N_20023,N_22319);
nor U24437 (N_24437,N_21162,N_20700);
and U24438 (N_24438,N_21988,N_20923);
nor U24439 (N_24439,N_21777,N_20379);
nor U24440 (N_24440,N_21797,N_20754);
or U24441 (N_24441,N_20037,N_20981);
nand U24442 (N_24442,N_20774,N_20911);
and U24443 (N_24443,N_22076,N_20288);
and U24444 (N_24444,N_22429,N_20968);
xor U24445 (N_24445,N_20347,N_21383);
nor U24446 (N_24446,N_22117,N_21961);
and U24447 (N_24447,N_20411,N_21423);
nand U24448 (N_24448,N_21359,N_22216);
nand U24449 (N_24449,N_20392,N_21076);
or U24450 (N_24450,N_20298,N_22256);
nand U24451 (N_24451,N_21855,N_20511);
xor U24452 (N_24452,N_20337,N_21393);
xnor U24453 (N_24453,N_20942,N_21039);
nand U24454 (N_24454,N_20645,N_21878);
xor U24455 (N_24455,N_20911,N_22138);
nor U24456 (N_24456,N_20190,N_21934);
nand U24457 (N_24457,N_20585,N_21662);
nand U24458 (N_24458,N_20718,N_21600);
nand U24459 (N_24459,N_20211,N_20289);
nand U24460 (N_24460,N_21607,N_21969);
nand U24461 (N_24461,N_21476,N_21238);
nand U24462 (N_24462,N_21614,N_20187);
nor U24463 (N_24463,N_20348,N_20499);
xor U24464 (N_24464,N_21958,N_20211);
or U24465 (N_24465,N_21103,N_20886);
and U24466 (N_24466,N_20899,N_21087);
or U24467 (N_24467,N_20966,N_21854);
xnor U24468 (N_24468,N_21367,N_22274);
xor U24469 (N_24469,N_21696,N_20061);
xnor U24470 (N_24470,N_22039,N_21138);
and U24471 (N_24471,N_20783,N_21366);
nand U24472 (N_24472,N_22181,N_22068);
nand U24473 (N_24473,N_21927,N_22368);
xor U24474 (N_24474,N_21000,N_22194);
and U24475 (N_24475,N_21056,N_21263);
nor U24476 (N_24476,N_21570,N_20970);
nor U24477 (N_24477,N_22092,N_21547);
xor U24478 (N_24478,N_20714,N_21332);
and U24479 (N_24479,N_21426,N_20839);
or U24480 (N_24480,N_20372,N_20560);
nor U24481 (N_24481,N_21344,N_20030);
or U24482 (N_24482,N_21000,N_21934);
and U24483 (N_24483,N_20070,N_21236);
nor U24484 (N_24484,N_20827,N_22307);
or U24485 (N_24485,N_20358,N_20054);
nor U24486 (N_24486,N_21231,N_20320);
and U24487 (N_24487,N_20541,N_20821);
nand U24488 (N_24488,N_22011,N_21858);
nor U24489 (N_24489,N_21903,N_20811);
and U24490 (N_24490,N_21431,N_20464);
nor U24491 (N_24491,N_20528,N_20385);
nor U24492 (N_24492,N_21078,N_21966);
nor U24493 (N_24493,N_20475,N_20860);
nand U24494 (N_24494,N_21567,N_20879);
nor U24495 (N_24495,N_21021,N_20592);
nor U24496 (N_24496,N_20532,N_21072);
and U24497 (N_24497,N_22232,N_22211);
nor U24498 (N_24498,N_21647,N_20833);
or U24499 (N_24499,N_22287,N_20722);
and U24500 (N_24500,N_21706,N_20762);
nand U24501 (N_24501,N_21576,N_21480);
xor U24502 (N_24502,N_22350,N_22313);
or U24503 (N_24503,N_21871,N_22331);
xor U24504 (N_24504,N_22448,N_21865);
nand U24505 (N_24505,N_20519,N_20106);
xor U24506 (N_24506,N_21353,N_20009);
nand U24507 (N_24507,N_21606,N_21187);
xnor U24508 (N_24508,N_20381,N_21823);
nand U24509 (N_24509,N_20037,N_21512);
or U24510 (N_24510,N_20001,N_21058);
xor U24511 (N_24511,N_22210,N_21693);
and U24512 (N_24512,N_20989,N_21058);
xnor U24513 (N_24513,N_21457,N_21298);
xor U24514 (N_24514,N_21927,N_21201);
and U24515 (N_24515,N_22499,N_21889);
xor U24516 (N_24516,N_20480,N_21629);
nor U24517 (N_24517,N_20758,N_20199);
nor U24518 (N_24518,N_22221,N_21685);
nor U24519 (N_24519,N_21873,N_21764);
xor U24520 (N_24520,N_20522,N_20314);
nand U24521 (N_24521,N_22240,N_20379);
xnor U24522 (N_24522,N_20047,N_21722);
xor U24523 (N_24523,N_20326,N_21543);
xnor U24524 (N_24524,N_20448,N_21615);
xor U24525 (N_24525,N_22421,N_22196);
xor U24526 (N_24526,N_22351,N_21802);
xor U24527 (N_24527,N_22243,N_20959);
or U24528 (N_24528,N_20141,N_21945);
xnor U24529 (N_24529,N_22375,N_20717);
nor U24530 (N_24530,N_21853,N_20743);
xor U24531 (N_24531,N_20924,N_20493);
and U24532 (N_24532,N_20954,N_21052);
and U24533 (N_24533,N_21788,N_20102);
or U24534 (N_24534,N_20110,N_21313);
xnor U24535 (N_24535,N_21713,N_21799);
nand U24536 (N_24536,N_20861,N_21845);
xor U24537 (N_24537,N_20704,N_20675);
xor U24538 (N_24538,N_21218,N_20386);
xor U24539 (N_24539,N_21897,N_20177);
xnor U24540 (N_24540,N_22487,N_21990);
nor U24541 (N_24541,N_21391,N_20013);
nor U24542 (N_24542,N_21107,N_21866);
nor U24543 (N_24543,N_20035,N_20351);
nor U24544 (N_24544,N_22158,N_20648);
nand U24545 (N_24545,N_20402,N_20819);
nor U24546 (N_24546,N_20932,N_20294);
or U24547 (N_24547,N_21016,N_21504);
nand U24548 (N_24548,N_20478,N_21330);
nor U24549 (N_24549,N_21686,N_20100);
nor U24550 (N_24550,N_22350,N_22081);
or U24551 (N_24551,N_22402,N_20284);
and U24552 (N_24552,N_20624,N_20774);
or U24553 (N_24553,N_21021,N_20212);
and U24554 (N_24554,N_22458,N_22024);
and U24555 (N_24555,N_20977,N_22463);
and U24556 (N_24556,N_22221,N_21904);
nor U24557 (N_24557,N_21834,N_21013);
or U24558 (N_24558,N_21920,N_21585);
and U24559 (N_24559,N_21249,N_22346);
xor U24560 (N_24560,N_20127,N_20403);
nor U24561 (N_24561,N_20140,N_22313);
nor U24562 (N_24562,N_22439,N_22250);
or U24563 (N_24563,N_20488,N_21612);
nand U24564 (N_24564,N_21010,N_21466);
xnor U24565 (N_24565,N_21580,N_21112);
or U24566 (N_24566,N_22433,N_22303);
nand U24567 (N_24567,N_21181,N_21417);
nand U24568 (N_24568,N_20001,N_20588);
nor U24569 (N_24569,N_20877,N_22082);
nor U24570 (N_24570,N_20627,N_20536);
xnor U24571 (N_24571,N_20884,N_20635);
nand U24572 (N_24572,N_22334,N_21464);
or U24573 (N_24573,N_22428,N_20488);
nand U24574 (N_24574,N_20290,N_20906);
nor U24575 (N_24575,N_20068,N_21065);
and U24576 (N_24576,N_20896,N_21453);
nand U24577 (N_24577,N_21117,N_20329);
nor U24578 (N_24578,N_21829,N_22100);
nor U24579 (N_24579,N_22114,N_21308);
or U24580 (N_24580,N_20652,N_21226);
nor U24581 (N_24581,N_21072,N_20359);
or U24582 (N_24582,N_20678,N_21102);
and U24583 (N_24583,N_20616,N_21664);
nor U24584 (N_24584,N_20091,N_21606);
xor U24585 (N_24585,N_21145,N_22382);
nand U24586 (N_24586,N_22194,N_21423);
nor U24587 (N_24587,N_20636,N_20925);
nand U24588 (N_24588,N_20065,N_21635);
and U24589 (N_24589,N_20870,N_22081);
or U24590 (N_24590,N_20091,N_21632);
nor U24591 (N_24591,N_20522,N_22420);
nor U24592 (N_24592,N_21103,N_21156);
nor U24593 (N_24593,N_21330,N_20730);
xor U24594 (N_24594,N_22014,N_20069);
nand U24595 (N_24595,N_22265,N_21590);
xnor U24596 (N_24596,N_20313,N_21599);
or U24597 (N_24597,N_22030,N_22091);
nand U24598 (N_24598,N_20119,N_21184);
nand U24599 (N_24599,N_21017,N_20917);
xor U24600 (N_24600,N_21967,N_21689);
or U24601 (N_24601,N_22344,N_20983);
xnor U24602 (N_24602,N_21059,N_22236);
nor U24603 (N_24603,N_21002,N_22063);
or U24604 (N_24604,N_21862,N_21073);
nand U24605 (N_24605,N_22200,N_22007);
or U24606 (N_24606,N_22190,N_20871);
and U24607 (N_24607,N_20150,N_22002);
and U24608 (N_24608,N_22156,N_22329);
xor U24609 (N_24609,N_20652,N_20367);
xor U24610 (N_24610,N_20354,N_21214);
or U24611 (N_24611,N_22276,N_21964);
nor U24612 (N_24612,N_21216,N_21833);
or U24613 (N_24613,N_21305,N_21600);
and U24614 (N_24614,N_20341,N_21757);
nor U24615 (N_24615,N_21594,N_21271);
xnor U24616 (N_24616,N_20092,N_22060);
nor U24617 (N_24617,N_21542,N_21226);
nand U24618 (N_24618,N_22387,N_20357);
nand U24619 (N_24619,N_21918,N_21359);
and U24620 (N_24620,N_20025,N_21725);
xnor U24621 (N_24621,N_21493,N_21701);
or U24622 (N_24622,N_22109,N_20723);
nand U24623 (N_24623,N_22064,N_20396);
xor U24624 (N_24624,N_22267,N_20406);
or U24625 (N_24625,N_20528,N_21101);
xnor U24626 (N_24626,N_21240,N_20392);
nor U24627 (N_24627,N_21433,N_20625);
and U24628 (N_24628,N_22013,N_20514);
and U24629 (N_24629,N_20503,N_20704);
nand U24630 (N_24630,N_21930,N_22219);
and U24631 (N_24631,N_22088,N_21108);
xnor U24632 (N_24632,N_20862,N_22130);
or U24633 (N_24633,N_21111,N_21340);
nor U24634 (N_24634,N_21990,N_22076);
nand U24635 (N_24635,N_21684,N_20968);
nor U24636 (N_24636,N_20093,N_22258);
xnor U24637 (N_24637,N_20363,N_21123);
and U24638 (N_24638,N_21419,N_20640);
nand U24639 (N_24639,N_22392,N_21902);
and U24640 (N_24640,N_20453,N_21288);
or U24641 (N_24641,N_21539,N_22254);
xnor U24642 (N_24642,N_22198,N_21148);
xnor U24643 (N_24643,N_20193,N_22496);
nand U24644 (N_24644,N_20620,N_21769);
and U24645 (N_24645,N_21728,N_21265);
nand U24646 (N_24646,N_20539,N_21532);
or U24647 (N_24647,N_20291,N_20382);
nor U24648 (N_24648,N_21825,N_20680);
or U24649 (N_24649,N_21916,N_22188);
nor U24650 (N_24650,N_21842,N_21017);
nor U24651 (N_24651,N_21554,N_21755);
or U24652 (N_24652,N_20022,N_20096);
xnor U24653 (N_24653,N_20391,N_20264);
nand U24654 (N_24654,N_20274,N_20907);
nor U24655 (N_24655,N_20957,N_20041);
and U24656 (N_24656,N_21605,N_20985);
nor U24657 (N_24657,N_22479,N_20840);
and U24658 (N_24658,N_21909,N_20704);
xnor U24659 (N_24659,N_21412,N_21990);
xnor U24660 (N_24660,N_20843,N_22011);
and U24661 (N_24661,N_21271,N_20452);
nand U24662 (N_24662,N_21953,N_21264);
xor U24663 (N_24663,N_21539,N_21131);
xor U24664 (N_24664,N_21522,N_20360);
or U24665 (N_24665,N_20025,N_20189);
nand U24666 (N_24666,N_20110,N_21287);
nand U24667 (N_24667,N_20685,N_21480);
nand U24668 (N_24668,N_22038,N_20693);
xnor U24669 (N_24669,N_21817,N_21841);
nand U24670 (N_24670,N_21563,N_20015);
or U24671 (N_24671,N_22081,N_20943);
or U24672 (N_24672,N_21850,N_20496);
nor U24673 (N_24673,N_21943,N_22441);
nand U24674 (N_24674,N_20677,N_22243);
xnor U24675 (N_24675,N_20884,N_20488);
nand U24676 (N_24676,N_21010,N_20633);
or U24677 (N_24677,N_21418,N_21288);
nand U24678 (N_24678,N_21483,N_20660);
or U24679 (N_24679,N_20445,N_20267);
and U24680 (N_24680,N_21579,N_20562);
nor U24681 (N_24681,N_21056,N_21505);
and U24682 (N_24682,N_21155,N_22137);
nor U24683 (N_24683,N_20904,N_22238);
or U24684 (N_24684,N_22097,N_21832);
xnor U24685 (N_24685,N_21316,N_22126);
nor U24686 (N_24686,N_21590,N_21573);
and U24687 (N_24687,N_20987,N_20495);
and U24688 (N_24688,N_22018,N_20739);
nor U24689 (N_24689,N_20348,N_20855);
xor U24690 (N_24690,N_20168,N_20181);
nand U24691 (N_24691,N_20113,N_21758);
or U24692 (N_24692,N_21327,N_21484);
or U24693 (N_24693,N_21306,N_20005);
nand U24694 (N_24694,N_22299,N_20470);
or U24695 (N_24695,N_21503,N_20794);
xor U24696 (N_24696,N_20091,N_21390);
nand U24697 (N_24697,N_21339,N_20290);
nand U24698 (N_24698,N_21993,N_21576);
or U24699 (N_24699,N_21951,N_21572);
nor U24700 (N_24700,N_20338,N_22460);
or U24701 (N_24701,N_20018,N_22260);
and U24702 (N_24702,N_22397,N_20536);
or U24703 (N_24703,N_21647,N_21888);
nor U24704 (N_24704,N_22365,N_22183);
nor U24705 (N_24705,N_21950,N_21690);
or U24706 (N_24706,N_20086,N_21086);
nand U24707 (N_24707,N_21328,N_21363);
and U24708 (N_24708,N_22360,N_20472);
nor U24709 (N_24709,N_20843,N_20432);
nand U24710 (N_24710,N_20469,N_22258);
nor U24711 (N_24711,N_21031,N_22452);
nand U24712 (N_24712,N_20933,N_21200);
and U24713 (N_24713,N_20807,N_21854);
nor U24714 (N_24714,N_20164,N_21792);
nor U24715 (N_24715,N_20600,N_21951);
nor U24716 (N_24716,N_22323,N_21534);
and U24717 (N_24717,N_22484,N_21244);
nand U24718 (N_24718,N_22265,N_20402);
and U24719 (N_24719,N_20868,N_22000);
or U24720 (N_24720,N_21579,N_22408);
or U24721 (N_24721,N_21439,N_21694);
and U24722 (N_24722,N_20111,N_21677);
nand U24723 (N_24723,N_22287,N_20891);
xnor U24724 (N_24724,N_20678,N_22371);
and U24725 (N_24725,N_21921,N_20532);
or U24726 (N_24726,N_21319,N_21596);
xor U24727 (N_24727,N_20648,N_20397);
nor U24728 (N_24728,N_20480,N_21631);
xor U24729 (N_24729,N_21987,N_22419);
nor U24730 (N_24730,N_20790,N_21689);
and U24731 (N_24731,N_21361,N_22331);
and U24732 (N_24732,N_20472,N_21395);
and U24733 (N_24733,N_21712,N_20999);
nand U24734 (N_24734,N_20126,N_22473);
or U24735 (N_24735,N_20117,N_20542);
nand U24736 (N_24736,N_20772,N_22305);
and U24737 (N_24737,N_22365,N_20018);
and U24738 (N_24738,N_22268,N_22303);
or U24739 (N_24739,N_21382,N_21499);
xnor U24740 (N_24740,N_22417,N_22297);
and U24741 (N_24741,N_21311,N_20525);
nand U24742 (N_24742,N_22311,N_20399);
nor U24743 (N_24743,N_20640,N_20426);
xnor U24744 (N_24744,N_21869,N_21649);
xor U24745 (N_24745,N_20105,N_20504);
nand U24746 (N_24746,N_21801,N_20765);
or U24747 (N_24747,N_22438,N_20994);
and U24748 (N_24748,N_21910,N_20267);
xnor U24749 (N_24749,N_21661,N_20561);
nor U24750 (N_24750,N_21880,N_20309);
or U24751 (N_24751,N_22102,N_20358);
or U24752 (N_24752,N_22263,N_21183);
xnor U24753 (N_24753,N_20749,N_21391);
xor U24754 (N_24754,N_21652,N_21754);
or U24755 (N_24755,N_22393,N_20026);
nand U24756 (N_24756,N_21248,N_22464);
and U24757 (N_24757,N_21325,N_20344);
or U24758 (N_24758,N_20402,N_20319);
nor U24759 (N_24759,N_20995,N_21325);
or U24760 (N_24760,N_21488,N_21880);
xor U24761 (N_24761,N_20483,N_20611);
nand U24762 (N_24762,N_21000,N_20897);
xor U24763 (N_24763,N_21808,N_21768);
nand U24764 (N_24764,N_22248,N_21496);
and U24765 (N_24765,N_21253,N_22379);
nand U24766 (N_24766,N_20213,N_22368);
and U24767 (N_24767,N_21448,N_21266);
nor U24768 (N_24768,N_20756,N_21529);
and U24769 (N_24769,N_21568,N_20682);
nand U24770 (N_24770,N_20015,N_21731);
nor U24771 (N_24771,N_20002,N_21767);
nor U24772 (N_24772,N_21288,N_22323);
nand U24773 (N_24773,N_20407,N_20751);
nor U24774 (N_24774,N_20504,N_21336);
nand U24775 (N_24775,N_20265,N_20489);
xnor U24776 (N_24776,N_20702,N_20706);
xnor U24777 (N_24777,N_20400,N_21047);
and U24778 (N_24778,N_22164,N_21642);
or U24779 (N_24779,N_21030,N_21660);
nor U24780 (N_24780,N_21396,N_20087);
xor U24781 (N_24781,N_22326,N_20139);
and U24782 (N_24782,N_20253,N_20521);
xnor U24783 (N_24783,N_20655,N_20755);
or U24784 (N_24784,N_20809,N_22068);
nand U24785 (N_24785,N_20831,N_21058);
nand U24786 (N_24786,N_21451,N_20350);
and U24787 (N_24787,N_21544,N_21932);
nor U24788 (N_24788,N_20344,N_21363);
nand U24789 (N_24789,N_20702,N_21267);
xnor U24790 (N_24790,N_21459,N_20161);
or U24791 (N_24791,N_20621,N_22301);
or U24792 (N_24792,N_21839,N_22410);
nand U24793 (N_24793,N_21624,N_21467);
xor U24794 (N_24794,N_20106,N_21719);
nand U24795 (N_24795,N_20757,N_20054);
nand U24796 (N_24796,N_20888,N_21600);
or U24797 (N_24797,N_20696,N_22419);
and U24798 (N_24798,N_22106,N_22351);
nor U24799 (N_24799,N_20371,N_20896);
nand U24800 (N_24800,N_21340,N_21670);
nor U24801 (N_24801,N_20205,N_20274);
or U24802 (N_24802,N_20450,N_20227);
and U24803 (N_24803,N_21081,N_21909);
and U24804 (N_24804,N_21007,N_20274);
or U24805 (N_24805,N_21870,N_21375);
xor U24806 (N_24806,N_22411,N_21065);
nor U24807 (N_24807,N_21963,N_20882);
or U24808 (N_24808,N_21717,N_21888);
nand U24809 (N_24809,N_21445,N_21783);
or U24810 (N_24810,N_20298,N_20794);
nor U24811 (N_24811,N_22253,N_22064);
xnor U24812 (N_24812,N_20069,N_20920);
nand U24813 (N_24813,N_21736,N_21827);
nor U24814 (N_24814,N_21304,N_20831);
xnor U24815 (N_24815,N_22116,N_21315);
nor U24816 (N_24816,N_22291,N_22235);
xor U24817 (N_24817,N_21854,N_21056);
xnor U24818 (N_24818,N_21167,N_20501);
or U24819 (N_24819,N_20250,N_20831);
and U24820 (N_24820,N_22184,N_22462);
or U24821 (N_24821,N_21590,N_20267);
and U24822 (N_24822,N_22313,N_22198);
nor U24823 (N_24823,N_21411,N_20558);
and U24824 (N_24824,N_20254,N_22295);
or U24825 (N_24825,N_22481,N_22320);
nor U24826 (N_24826,N_21523,N_21801);
nand U24827 (N_24827,N_20158,N_20457);
and U24828 (N_24828,N_20683,N_21547);
xnor U24829 (N_24829,N_20732,N_21155);
xor U24830 (N_24830,N_20558,N_21112);
and U24831 (N_24831,N_20237,N_21172);
nand U24832 (N_24832,N_20931,N_21611);
xor U24833 (N_24833,N_22387,N_22201);
and U24834 (N_24834,N_21595,N_22119);
nand U24835 (N_24835,N_22473,N_21420);
and U24836 (N_24836,N_20303,N_20532);
or U24837 (N_24837,N_20370,N_20725);
nand U24838 (N_24838,N_22050,N_20560);
or U24839 (N_24839,N_20580,N_20901);
nand U24840 (N_24840,N_21413,N_20630);
xor U24841 (N_24841,N_21782,N_20623);
nand U24842 (N_24842,N_22444,N_21551);
or U24843 (N_24843,N_21945,N_20090);
and U24844 (N_24844,N_20180,N_22292);
xor U24845 (N_24845,N_21897,N_21313);
or U24846 (N_24846,N_22341,N_21945);
and U24847 (N_24847,N_20979,N_20171);
and U24848 (N_24848,N_20557,N_20514);
or U24849 (N_24849,N_21120,N_20549);
xnor U24850 (N_24850,N_21994,N_20542);
nand U24851 (N_24851,N_21805,N_21432);
xor U24852 (N_24852,N_21555,N_20247);
and U24853 (N_24853,N_20838,N_20297);
and U24854 (N_24854,N_21673,N_21268);
and U24855 (N_24855,N_20529,N_22315);
nand U24856 (N_24856,N_21839,N_20181);
xnor U24857 (N_24857,N_20028,N_21177);
and U24858 (N_24858,N_20161,N_21506);
or U24859 (N_24859,N_20640,N_22309);
or U24860 (N_24860,N_21078,N_20603);
and U24861 (N_24861,N_21991,N_22344);
nor U24862 (N_24862,N_22479,N_21340);
nand U24863 (N_24863,N_20268,N_20562);
xor U24864 (N_24864,N_22281,N_20463);
nor U24865 (N_24865,N_21530,N_21383);
or U24866 (N_24866,N_21678,N_21932);
or U24867 (N_24867,N_22045,N_22332);
or U24868 (N_24868,N_22303,N_21118);
and U24869 (N_24869,N_22032,N_22356);
nand U24870 (N_24870,N_21525,N_21368);
or U24871 (N_24871,N_20550,N_21000);
nor U24872 (N_24872,N_21110,N_21676);
and U24873 (N_24873,N_20139,N_21938);
nand U24874 (N_24874,N_20574,N_20234);
and U24875 (N_24875,N_20886,N_20537);
and U24876 (N_24876,N_20549,N_20850);
or U24877 (N_24877,N_20298,N_22445);
and U24878 (N_24878,N_22110,N_20247);
xor U24879 (N_24879,N_20399,N_20213);
and U24880 (N_24880,N_21754,N_22493);
or U24881 (N_24881,N_21236,N_22118);
xor U24882 (N_24882,N_21638,N_20220);
and U24883 (N_24883,N_21486,N_20259);
and U24884 (N_24884,N_21234,N_22164);
nor U24885 (N_24885,N_20014,N_21879);
and U24886 (N_24886,N_21522,N_20285);
nor U24887 (N_24887,N_21427,N_20249);
nand U24888 (N_24888,N_20285,N_20584);
and U24889 (N_24889,N_21959,N_22193);
nor U24890 (N_24890,N_22485,N_21603);
and U24891 (N_24891,N_21788,N_22424);
nand U24892 (N_24892,N_21873,N_20036);
nand U24893 (N_24893,N_21004,N_21031);
xor U24894 (N_24894,N_21072,N_20573);
xnor U24895 (N_24895,N_22483,N_20008);
and U24896 (N_24896,N_21044,N_21484);
or U24897 (N_24897,N_21750,N_22224);
nor U24898 (N_24898,N_22241,N_20264);
nor U24899 (N_24899,N_20250,N_21708);
and U24900 (N_24900,N_22253,N_21563);
and U24901 (N_24901,N_21024,N_22035);
or U24902 (N_24902,N_20673,N_21486);
or U24903 (N_24903,N_20615,N_21827);
or U24904 (N_24904,N_21202,N_22374);
nor U24905 (N_24905,N_21744,N_20043);
or U24906 (N_24906,N_21917,N_21691);
nor U24907 (N_24907,N_21063,N_20950);
nor U24908 (N_24908,N_21612,N_20786);
and U24909 (N_24909,N_20091,N_22228);
xor U24910 (N_24910,N_22247,N_20239);
nor U24911 (N_24911,N_20237,N_20617);
xnor U24912 (N_24912,N_21019,N_20849);
nand U24913 (N_24913,N_21217,N_22140);
or U24914 (N_24914,N_21314,N_22097);
xor U24915 (N_24915,N_21266,N_20743);
or U24916 (N_24916,N_21386,N_20437);
nand U24917 (N_24917,N_21606,N_21863);
nand U24918 (N_24918,N_21111,N_21214);
nor U24919 (N_24919,N_20730,N_21122);
nand U24920 (N_24920,N_21792,N_22376);
nor U24921 (N_24921,N_22213,N_20201);
and U24922 (N_24922,N_21898,N_21991);
nand U24923 (N_24923,N_20074,N_20630);
and U24924 (N_24924,N_21957,N_21324);
xnor U24925 (N_24925,N_21785,N_20349);
nand U24926 (N_24926,N_20284,N_20001);
nor U24927 (N_24927,N_22333,N_20667);
nor U24928 (N_24928,N_21861,N_20383);
or U24929 (N_24929,N_22278,N_21937);
xnor U24930 (N_24930,N_20561,N_21323);
nor U24931 (N_24931,N_21514,N_22103);
nor U24932 (N_24932,N_20499,N_21506);
xor U24933 (N_24933,N_22065,N_21132);
nor U24934 (N_24934,N_21937,N_20326);
or U24935 (N_24935,N_20782,N_20093);
nor U24936 (N_24936,N_21984,N_21111);
xnor U24937 (N_24937,N_22223,N_20356);
xnor U24938 (N_24938,N_20198,N_21769);
nand U24939 (N_24939,N_22384,N_22327);
nand U24940 (N_24940,N_21061,N_21105);
or U24941 (N_24941,N_21959,N_20154);
or U24942 (N_24942,N_20192,N_21582);
and U24943 (N_24943,N_22175,N_20324);
and U24944 (N_24944,N_21774,N_20490);
nand U24945 (N_24945,N_22474,N_20075);
and U24946 (N_24946,N_20341,N_21576);
nor U24947 (N_24947,N_20328,N_21522);
and U24948 (N_24948,N_22466,N_21393);
or U24949 (N_24949,N_20555,N_21272);
and U24950 (N_24950,N_22110,N_22425);
xnor U24951 (N_24951,N_21755,N_21502);
or U24952 (N_24952,N_21066,N_21591);
or U24953 (N_24953,N_20546,N_20158);
nand U24954 (N_24954,N_22441,N_20514);
or U24955 (N_24955,N_22448,N_21559);
nand U24956 (N_24956,N_20098,N_21540);
xnor U24957 (N_24957,N_21185,N_20208);
xnor U24958 (N_24958,N_20445,N_21630);
and U24959 (N_24959,N_21099,N_20065);
xnor U24960 (N_24960,N_20042,N_20561);
xor U24961 (N_24961,N_20087,N_20191);
nor U24962 (N_24962,N_22133,N_21496);
xor U24963 (N_24963,N_21458,N_21955);
xor U24964 (N_24964,N_20807,N_22162);
nor U24965 (N_24965,N_20085,N_20670);
or U24966 (N_24966,N_22121,N_21872);
and U24967 (N_24967,N_20860,N_21059);
xnor U24968 (N_24968,N_20071,N_21578);
xnor U24969 (N_24969,N_20376,N_20972);
or U24970 (N_24970,N_21201,N_20353);
nor U24971 (N_24971,N_21143,N_22350);
and U24972 (N_24972,N_22355,N_21843);
and U24973 (N_24973,N_21128,N_21894);
xor U24974 (N_24974,N_20660,N_22239);
and U24975 (N_24975,N_21911,N_21822);
or U24976 (N_24976,N_21317,N_20235);
nand U24977 (N_24977,N_20618,N_21070);
or U24978 (N_24978,N_21301,N_21861);
xnor U24979 (N_24979,N_21608,N_20935);
xnor U24980 (N_24980,N_20592,N_20029);
nand U24981 (N_24981,N_21752,N_22334);
nor U24982 (N_24982,N_21835,N_22034);
and U24983 (N_24983,N_20978,N_21909);
nand U24984 (N_24984,N_21865,N_22361);
xor U24985 (N_24985,N_21513,N_21379);
xor U24986 (N_24986,N_20246,N_21536);
xnor U24987 (N_24987,N_21701,N_20988);
xor U24988 (N_24988,N_22433,N_20211);
or U24989 (N_24989,N_21713,N_21518);
nor U24990 (N_24990,N_20483,N_20554);
xnor U24991 (N_24991,N_21477,N_21781);
or U24992 (N_24992,N_21237,N_21556);
nand U24993 (N_24993,N_20046,N_21344);
or U24994 (N_24994,N_22022,N_21973);
nor U24995 (N_24995,N_20384,N_21534);
or U24996 (N_24996,N_22269,N_21183);
and U24997 (N_24997,N_20876,N_21562);
xor U24998 (N_24998,N_20064,N_20787);
nor U24999 (N_24999,N_21465,N_21069);
or U25000 (N_25000,N_23484,N_24199);
or U25001 (N_25001,N_22816,N_23314);
nand U25002 (N_25002,N_24764,N_23480);
nor U25003 (N_25003,N_22958,N_22806);
or U25004 (N_25004,N_24293,N_23332);
xnor U25005 (N_25005,N_23953,N_24019);
nor U25006 (N_25006,N_23989,N_23329);
nor U25007 (N_25007,N_24458,N_24406);
nand U25008 (N_25008,N_23138,N_22839);
or U25009 (N_25009,N_24770,N_24776);
or U25010 (N_25010,N_23583,N_23994);
or U25011 (N_25011,N_23101,N_22683);
or U25012 (N_25012,N_23882,N_23053);
and U25013 (N_25013,N_22543,N_23768);
xor U25014 (N_25014,N_23561,N_24800);
or U25015 (N_25015,N_23373,N_22717);
nand U25016 (N_25016,N_22504,N_24677);
or U25017 (N_25017,N_23607,N_23950);
and U25018 (N_25018,N_22945,N_23401);
nor U25019 (N_25019,N_24837,N_24174);
or U25020 (N_25020,N_24734,N_22517);
xor U25021 (N_25021,N_22557,N_23837);
or U25022 (N_25022,N_23115,N_23374);
or U25023 (N_25023,N_22848,N_23127);
nor U25024 (N_25024,N_22722,N_22752);
or U25025 (N_25025,N_22876,N_23615);
xor U25026 (N_25026,N_23553,N_24222);
nand U25027 (N_25027,N_24866,N_23995);
nand U25028 (N_25028,N_24785,N_23354);
xnor U25029 (N_25029,N_22679,N_24420);
nor U25030 (N_25030,N_22596,N_23214);
nor U25031 (N_25031,N_24249,N_24438);
and U25032 (N_25032,N_23830,N_24742);
nor U25033 (N_25033,N_24204,N_24018);
nand U25034 (N_25034,N_24404,N_23161);
or U25035 (N_25035,N_23941,N_24951);
nor U25036 (N_25036,N_23513,N_24806);
nand U25037 (N_25037,N_24993,N_23205);
nor U25038 (N_25038,N_23176,N_24361);
nand U25039 (N_25039,N_24384,N_24339);
or U25040 (N_25040,N_24394,N_24049);
xor U25041 (N_25041,N_22874,N_23915);
or U25042 (N_25042,N_23103,N_22592);
xor U25043 (N_25043,N_22818,N_22743);
and U25044 (N_25044,N_24484,N_23009);
xor U25045 (N_25045,N_24954,N_22828);
nor U25046 (N_25046,N_23520,N_23250);
and U25047 (N_25047,N_24156,N_24383);
xor U25048 (N_25048,N_24098,N_23661);
or U25049 (N_25049,N_24213,N_24869);
or U25050 (N_25050,N_23604,N_23828);
xnor U25051 (N_25051,N_23310,N_24263);
or U25052 (N_25052,N_23134,N_22558);
or U25053 (N_25053,N_23588,N_22900);
or U25054 (N_25054,N_24259,N_24364);
and U25055 (N_25055,N_24336,N_22613);
or U25056 (N_25056,N_22979,N_24190);
or U25057 (N_25057,N_24914,N_24166);
nor U25058 (N_25058,N_23086,N_24781);
or U25059 (N_25059,N_24714,N_23946);
nor U25060 (N_25060,N_23307,N_23706);
and U25061 (N_25061,N_22823,N_24240);
nor U25062 (N_25062,N_24159,N_23933);
xor U25063 (N_25063,N_22616,N_24242);
nor U25064 (N_25064,N_24091,N_23562);
nand U25065 (N_25065,N_23699,N_23461);
or U25066 (N_25066,N_24856,N_22849);
or U25067 (N_25067,N_24120,N_24984);
nor U25068 (N_25068,N_24437,N_22924);
or U25069 (N_25069,N_22676,N_23185);
xnor U25070 (N_25070,N_23534,N_24141);
xnor U25071 (N_25071,N_23133,N_23640);
and U25072 (N_25072,N_22782,N_24121);
and U25073 (N_25073,N_24606,N_24890);
nand U25074 (N_25074,N_24173,N_23456);
or U25075 (N_25075,N_23523,N_23398);
and U25076 (N_25076,N_22603,N_22608);
and U25077 (N_25077,N_24235,N_22977);
xor U25078 (N_25078,N_24532,N_23068);
or U25079 (N_25079,N_23780,N_22912);
nand U25080 (N_25080,N_24381,N_24231);
or U25081 (N_25081,N_23939,N_22980);
or U25082 (N_25082,N_24185,N_23501);
and U25083 (N_25083,N_23741,N_22946);
or U25084 (N_25084,N_23696,N_22508);
nor U25085 (N_25085,N_24371,N_22646);
and U25086 (N_25086,N_22858,N_24071);
nor U25087 (N_25087,N_23611,N_24322);
and U25088 (N_25088,N_24841,N_24503);
or U25089 (N_25089,N_24473,N_24378);
nand U25090 (N_25090,N_24843,N_22801);
xor U25091 (N_25091,N_23648,N_23364);
or U25092 (N_25092,N_23548,N_23436);
nand U25093 (N_25093,N_23568,N_24833);
nand U25094 (N_25094,N_23217,N_24981);
and U25095 (N_25095,N_22634,N_24539);
and U25096 (N_25096,N_24630,N_24319);
or U25097 (N_25097,N_24502,N_22527);
nand U25098 (N_25098,N_23171,N_23111);
nand U25099 (N_25099,N_24106,N_23430);
xnor U25100 (N_25100,N_24139,N_22591);
and U25101 (N_25101,N_24063,N_24766);
xor U25102 (N_25102,N_23884,N_23312);
or U25103 (N_25103,N_22626,N_23427);
and U25104 (N_25104,N_24906,N_22664);
nor U25105 (N_25105,N_23844,N_22642);
or U25106 (N_25106,N_23049,N_23324);
or U25107 (N_25107,N_24513,N_24635);
nor U25108 (N_25108,N_24119,N_23452);
xor U25109 (N_25109,N_23984,N_23424);
xnor U25110 (N_25110,N_24909,N_24672);
nand U25111 (N_25111,N_24789,N_24899);
nor U25112 (N_25112,N_24868,N_23034);
nand U25113 (N_25113,N_23449,N_22878);
nand U25114 (N_25114,N_22619,N_23985);
nor U25115 (N_25115,N_22810,N_24146);
or U25116 (N_25116,N_22851,N_24418);
xnor U25117 (N_25117,N_24634,N_24817);
nor U25118 (N_25118,N_23505,N_22789);
nand U25119 (N_25119,N_23090,N_23108);
nand U25120 (N_25120,N_23089,N_23740);
nand U25121 (N_25121,N_23067,N_24356);
or U25122 (N_25122,N_22716,N_23435);
xor U25123 (N_25123,N_23123,N_23499);
xnor U25124 (N_25124,N_23971,N_22767);
xnor U25125 (N_25125,N_23193,N_22565);
or U25126 (N_25126,N_24597,N_24186);
nor U25127 (N_25127,N_23457,N_22750);
xor U25128 (N_25128,N_22880,N_23496);
nor U25129 (N_25129,N_24352,N_23580);
xor U25130 (N_25130,N_23126,N_24609);
nor U25131 (N_25131,N_23316,N_22844);
and U25132 (N_25132,N_22667,N_24250);
nand U25133 (N_25133,N_24123,N_23151);
or U25134 (N_25134,N_23766,N_23709);
nand U25135 (N_25135,N_22726,N_23077);
and U25136 (N_25136,N_24508,N_24517);
nand U25137 (N_25137,N_23596,N_23061);
nand U25138 (N_25138,N_23085,N_24402);
nor U25139 (N_25139,N_23519,N_22872);
nand U25140 (N_25140,N_22533,N_23441);
xor U25141 (N_25141,N_22788,N_24689);
xor U25142 (N_25142,N_23448,N_23491);
nand U25143 (N_25143,N_23947,N_24160);
xor U25144 (N_25144,N_24820,N_23730);
and U25145 (N_25145,N_23243,N_23259);
nand U25146 (N_25146,N_23614,N_24592);
nand U25147 (N_25147,N_24345,N_23397);
or U25148 (N_25148,N_23206,N_24940);
nand U25149 (N_25149,N_23573,N_22837);
and U25150 (N_25150,N_24929,N_23464);
nand U25151 (N_25151,N_24246,N_23210);
nand U25152 (N_25152,N_23380,N_24772);
or U25153 (N_25153,N_22868,N_23535);
nand U25154 (N_25154,N_23536,N_23302);
nand U25155 (N_25155,N_23582,N_24663);
nand U25156 (N_25156,N_24978,N_23707);
and U25157 (N_25157,N_24970,N_22864);
and U25158 (N_25158,N_24538,N_23292);
or U25159 (N_25159,N_23843,N_24003);
nand U25160 (N_25160,N_24457,N_24005);
nand U25161 (N_25161,N_23684,N_23381);
or U25162 (N_25162,N_23518,N_24399);
and U25163 (N_25163,N_24587,N_24276);
or U25164 (N_25164,N_23031,N_22775);
and U25165 (N_25165,N_22700,N_23997);
or U25166 (N_25166,N_24939,N_23925);
nor U25167 (N_25167,N_22915,N_22635);
nand U25168 (N_25168,N_22822,N_23445);
or U25169 (N_25169,N_23306,N_24310);
or U25170 (N_25170,N_22771,N_23690);
nor U25171 (N_25171,N_24533,N_24673);
xor U25172 (N_25172,N_23966,N_23695);
nand U25173 (N_25173,N_23466,N_23271);
and U25174 (N_25174,N_24857,N_24715);
nand U25175 (N_25175,N_22781,N_24549);
nor U25176 (N_25176,N_23320,N_23043);
and U25177 (N_25177,N_24441,N_23195);
nand U25178 (N_25178,N_22925,N_24266);
and U25179 (N_25179,N_22833,N_23409);
or U25180 (N_25180,N_24616,N_24150);
nor U25181 (N_25181,N_24892,N_24813);
or U25182 (N_25182,N_23136,N_24669);
and U25183 (N_25183,N_24144,N_23679);
or U25184 (N_25184,N_24481,N_22836);
nor U25185 (N_25185,N_23112,N_23325);
nor U25186 (N_25186,N_23952,N_24783);
nand U25187 (N_25187,N_22831,N_24493);
or U25188 (N_25188,N_23825,N_22871);
nor U25189 (N_25189,N_22959,N_23152);
nand U25190 (N_25190,N_23581,N_24226);
or U25191 (N_25191,N_23092,N_24787);
xor U25192 (N_25192,N_22516,N_22827);
and U25193 (N_25193,N_24957,N_23621);
or U25194 (N_25194,N_23014,N_22933);
nand U25195 (N_25195,N_23039,N_24370);
nor U25196 (N_25196,N_24086,N_23608);
and U25197 (N_25197,N_23265,N_23635);
and U25198 (N_25198,N_23290,N_24456);
and U25199 (N_25199,N_24175,N_24492);
nor U25200 (N_25200,N_22681,N_23500);
and U25201 (N_25201,N_23274,N_22786);
or U25202 (N_25202,N_22918,N_24959);
and U25203 (N_25203,N_22675,N_24919);
nand U25204 (N_25204,N_22672,N_24720);
nand U25205 (N_25205,N_23718,N_22522);
xor U25206 (N_25206,N_24382,N_23973);
nand U25207 (N_25207,N_24923,N_23564);
and U25208 (N_25208,N_23649,N_23175);
xnor U25209 (N_25209,N_23450,N_23379);
nand U25210 (N_25210,N_22510,N_24969);
nand U25211 (N_25211,N_23164,N_23071);
nand U25212 (N_25212,N_23143,N_23342);
nand U25213 (N_25213,N_23428,N_24004);
and U25214 (N_25214,N_24330,N_24055);
or U25215 (N_25215,N_23743,N_24559);
nand U25216 (N_25216,N_24047,N_23815);
xor U25217 (N_25217,N_24862,N_24670);
and U25218 (N_25218,N_24229,N_23928);
nand U25219 (N_25219,N_24884,N_24271);
and U25220 (N_25220,N_24350,N_23128);
xnor U25221 (N_25221,N_24192,N_22597);
nor U25222 (N_25222,N_24140,N_22923);
and U25223 (N_25223,N_22873,N_24888);
nand U25224 (N_25224,N_23688,N_24595);
nor U25225 (N_25225,N_22559,N_22708);
and U25226 (N_25226,N_22554,N_23686);
nand U25227 (N_25227,N_24234,N_24851);
or U25228 (N_25228,N_24903,N_23764);
nand U25229 (N_25229,N_23600,N_24988);
or U25230 (N_25230,N_22567,N_24927);
nand U25231 (N_25231,N_23352,N_23572);
and U25232 (N_25232,N_22825,N_24994);
or U25233 (N_25233,N_24972,N_23189);
xnor U25234 (N_25234,N_23822,N_23145);
xnor U25235 (N_25235,N_24209,N_24829);
or U25236 (N_25236,N_23967,N_23685);
xor U25237 (N_25237,N_24839,N_23856);
xor U25238 (N_25238,N_24176,N_23159);
nand U25239 (N_25239,N_24499,N_24882);
nand U25240 (N_25240,N_23514,N_23318);
or U25241 (N_25241,N_24759,N_22986);
nand U25242 (N_25242,N_23204,N_24380);
nor U25243 (N_25243,N_22651,N_23808);
xor U25244 (N_25244,N_23305,N_22706);
nor U25245 (N_25245,N_22588,N_23129);
or U25246 (N_25246,N_23879,N_23862);
and U25247 (N_25247,N_23299,N_23948);
and U25248 (N_25248,N_24719,N_22714);
nand U25249 (N_25249,N_23030,N_23716);
xor U25250 (N_25250,N_24088,N_24550);
and U25251 (N_25251,N_23041,N_22698);
and U25252 (N_25252,N_24069,N_23473);
xor U25253 (N_25253,N_23551,N_22612);
nor U25254 (N_25254,N_22561,N_24389);
nor U25255 (N_25255,N_24385,N_22749);
nor U25256 (N_25256,N_24840,N_24621);
nand U25257 (N_25257,N_24908,N_23378);
nor U25258 (N_25258,N_23416,N_24497);
xnor U25259 (N_25259,N_23691,N_22660);
xnor U25260 (N_25260,N_24111,N_23917);
xor U25261 (N_25261,N_23747,N_22515);
and U25262 (N_25262,N_23539,N_22703);
nand U25263 (N_25263,N_23173,N_23836);
and U25264 (N_25264,N_24602,N_24642);
nand U25265 (N_25265,N_24082,N_23062);
xnor U25266 (N_25266,N_22916,N_24327);
or U25267 (N_25267,N_24318,N_23601);
or U25268 (N_25268,N_23227,N_23857);
nor U25269 (N_25269,N_22528,N_24943);
or U25270 (N_25270,N_23183,N_23664);
or U25271 (N_25271,N_24865,N_24053);
nand U25272 (N_25272,N_23717,N_22845);
and U25273 (N_25273,N_23390,N_24590);
nor U25274 (N_25274,N_24221,N_24022);
xnor U25275 (N_25275,N_23120,N_24396);
nand U25276 (N_25276,N_24237,N_23330);
and U25277 (N_25277,N_22766,N_23182);
or U25278 (N_25278,N_23872,N_23811);
and U25279 (N_25279,N_24596,N_23326);
or U25280 (N_25280,N_23238,N_23420);
nand U25281 (N_25281,N_22855,N_22539);
or U25282 (N_25282,N_23668,N_22610);
or U25283 (N_25283,N_24712,N_24081);
xnor U25284 (N_25284,N_24223,N_22802);
or U25285 (N_25285,N_22756,N_23272);
xor U25286 (N_25286,N_22884,N_22658);
xor U25287 (N_25287,N_23069,N_24520);
nand U25288 (N_25288,N_24207,N_23415);
and U25289 (N_25289,N_22746,N_22576);
nand U25290 (N_25290,N_24414,N_23345);
xor U25291 (N_25291,N_24200,N_24507);
nor U25292 (N_25292,N_24955,N_23074);
xnor U25293 (N_25293,N_24072,N_22637);
and U25294 (N_25294,N_24416,N_23486);
or U25295 (N_25295,N_24135,N_24067);
nor U25296 (N_25296,N_24126,N_24733);
nand U25297 (N_25297,N_24002,N_24485);
nand U25298 (N_25298,N_23525,N_24065);
xnor U25299 (N_25299,N_23976,N_23006);
nand U25300 (N_25300,N_24031,N_22704);
nor U25301 (N_25301,N_23926,N_24946);
and U25302 (N_25302,N_24683,N_24247);
xor U25303 (N_25303,N_24129,N_23076);
or U25304 (N_25304,N_23807,N_23019);
and U25305 (N_25305,N_23891,N_23021);
and U25306 (N_25306,N_24182,N_24703);
xnor U25307 (N_25307,N_23460,N_22908);
nor U25308 (N_25308,N_23512,N_23447);
or U25309 (N_25309,N_23052,N_24171);
or U25310 (N_25310,N_23774,N_22870);
xor U25311 (N_25311,N_24656,N_23005);
nor U25312 (N_25312,N_23760,N_24828);
nor U25313 (N_25313,N_23547,N_23488);
xor U25314 (N_25314,N_22906,N_23286);
or U25315 (N_25315,N_23493,N_22575);
and U25316 (N_25316,N_23529,N_24664);
and U25317 (N_25317,N_23404,N_24593);
nor U25318 (N_25318,N_22817,N_24832);
nor U25319 (N_25319,N_23890,N_23241);
or U25320 (N_25320,N_23870,N_22699);
xor U25321 (N_25321,N_22652,N_24046);
nand U25322 (N_25322,N_24024,N_22500);
nand U25323 (N_25323,N_24353,N_22982);
or U25324 (N_25324,N_24184,N_24536);
and U25325 (N_25325,N_24328,N_24277);
or U25326 (N_25326,N_24960,N_22725);
and U25327 (N_25327,N_24010,N_23483);
nor U25328 (N_25328,N_23284,N_23754);
nand U25329 (N_25329,N_23748,N_24372);
nor U25330 (N_25330,N_24580,N_23413);
nand U25331 (N_25331,N_24653,N_24627);
nor U25332 (N_25332,N_24285,N_22692);
or U25333 (N_25333,N_24208,N_24230);
nor U25334 (N_25334,N_23213,N_22795);
and U25335 (N_25335,N_23623,N_24478);
nand U25336 (N_25336,N_23226,N_23467);
xnor U25337 (N_25337,N_24858,N_22991);
xor U25338 (N_25338,N_24393,N_24962);
or U25339 (N_25339,N_23722,N_23405);
or U25340 (N_25340,N_24804,N_23749);
xnor U25341 (N_25341,N_22984,N_24085);
xnor U25342 (N_25342,N_24700,N_22955);
or U25343 (N_25343,N_24995,N_23918);
xnor U25344 (N_25344,N_24131,N_23975);
nor U25345 (N_25345,N_22742,N_24425);
nand U25346 (N_25346,N_24486,N_23659);
or U25347 (N_25347,N_22897,N_23794);
nor U25348 (N_25348,N_23365,N_23239);
nor U25349 (N_25349,N_24895,N_22800);
nand U25350 (N_25350,N_22883,N_24985);
and U25351 (N_25351,N_22663,N_23375);
nor U25352 (N_25352,N_24579,N_23526);
and U25353 (N_25353,N_22898,N_22744);
nand U25354 (N_25354,N_24203,N_24831);
nor U25355 (N_25355,N_24125,N_23293);
and U25356 (N_25356,N_24245,N_24138);
and U25357 (N_25357,N_23104,N_23280);
xor U25358 (N_25358,N_24116,N_23395);
or U25359 (N_25359,N_23058,N_22584);
and U25360 (N_25360,N_23554,N_22730);
xor U25361 (N_25361,N_24705,N_22776);
or U25362 (N_25362,N_23671,N_24886);
nand U25363 (N_25363,N_22785,N_24822);
or U25364 (N_25364,N_22830,N_23609);
nand U25365 (N_25365,N_24871,N_22525);
nor U25366 (N_25366,N_22702,N_24629);
or U25367 (N_25367,N_23056,N_22541);
xor U25368 (N_25368,N_23212,N_22920);
nor U25369 (N_25369,N_22620,N_24729);
nor U25370 (N_25370,N_22931,N_22896);
or U25371 (N_25371,N_22548,N_24922);
nand U25372 (N_25372,N_22987,N_24527);
xor U25373 (N_25373,N_23156,N_24183);
and U25374 (N_25374,N_22529,N_23494);
nor U25375 (N_25375,N_22573,N_23929);
xnor U25376 (N_25376,N_22507,N_24562);
and U25377 (N_25377,N_23383,N_22812);
xor U25378 (N_25378,N_23542,N_24608);
or U25379 (N_25379,N_23781,N_23093);
nand U25380 (N_25380,N_23869,N_23442);
or U25381 (N_25381,N_22772,N_23055);
nand U25382 (N_25382,N_23795,N_23957);
and U25383 (N_25383,N_24522,N_24738);
xnor U25384 (N_25384,N_23620,N_23935);
or U25385 (N_25385,N_24574,N_23046);
and U25386 (N_25386,N_24543,N_23225);
xor U25387 (N_25387,N_23786,N_23260);
xnor U25388 (N_25388,N_24750,N_24180);
xor U25389 (N_25389,N_23462,N_22994);
nor U25390 (N_25390,N_23969,N_24751);
xor U25391 (N_25391,N_24045,N_24289);
xor U25392 (N_25392,N_24278,N_22531);
xor U25393 (N_25393,N_24686,N_23389);
nor U25394 (N_25394,N_23240,N_24791);
nand U25395 (N_25395,N_24659,N_24913);
xor U25396 (N_25396,N_24101,N_24170);
and U25397 (N_25397,N_23465,N_24329);
nand U25398 (N_25398,N_24465,N_24523);
and U25399 (N_25399,N_23847,N_22627);
nor U25400 (N_25400,N_24386,N_22950);
xnor U25401 (N_25401,N_22583,N_22922);
or U25402 (N_25402,N_24287,N_23663);
or U25403 (N_25403,N_22857,N_23469);
xor U25404 (N_25404,N_23908,N_24638);
or U25405 (N_25405,N_23751,N_24479);
nand U25406 (N_25406,N_23453,N_24260);
nand U25407 (N_25407,N_23849,N_23516);
nor U25408 (N_25408,N_23258,N_23248);
and U25409 (N_25409,N_24525,N_22917);
and U25410 (N_25410,N_24976,N_24584);
or U25411 (N_25411,N_22606,N_24571);
and U25412 (N_25412,N_23081,N_24462);
nand U25413 (N_25413,N_24267,N_23013);
nor U25414 (N_25414,N_23017,N_24702);
and U25415 (N_25415,N_24104,N_22894);
nand U25416 (N_25416,N_22947,N_23082);
nand U25417 (N_25417,N_24557,N_23083);
nand U25418 (N_25418,N_24935,N_23059);
nor U25419 (N_25419,N_23924,N_23323);
and U25420 (N_25420,N_23921,N_24472);
and U25421 (N_25421,N_24324,N_22580);
nand U25422 (N_25422,N_24745,N_23545);
nand U25423 (N_25423,N_24652,N_23681);
nand U25424 (N_25424,N_23066,N_23683);
or U25425 (N_25425,N_23027,N_24586);
or U25426 (N_25426,N_24253,N_22589);
nand U25427 (N_25427,N_22919,N_23277);
or U25428 (N_25428,N_23692,N_23842);
nor U25429 (N_25429,N_24990,N_23713);
or U25430 (N_25430,N_24323,N_23698);
xnor U25431 (N_25431,N_24375,N_24818);
and U25432 (N_25432,N_24965,N_22526);
xnor U25433 (N_25433,N_23731,N_24007);
nand U25434 (N_25434,N_23287,N_23218);
nor U25435 (N_25435,N_24398,N_23744);
and U25436 (N_25436,N_22807,N_24035);
nor U25437 (N_25437,N_24690,N_24961);
nor U25438 (N_25438,N_24179,N_23657);
nor U25439 (N_25439,N_23602,N_22594);
nand U25440 (N_25440,N_23328,N_22733);
nor U25441 (N_25441,N_22555,N_24169);
or U25442 (N_25442,N_24915,N_24313);
and U25443 (N_25443,N_22768,N_23191);
and U25444 (N_25444,N_23281,N_24735);
xnor U25445 (N_25445,N_24448,N_23167);
nand U25446 (N_25446,N_23940,N_23508);
nor U25447 (N_25447,N_24570,N_24282);
nor U25448 (N_25448,N_23255,N_23215);
xor U25449 (N_25449,N_24708,N_23880);
or U25450 (N_25450,N_24092,N_22774);
and U25451 (N_25451,N_24573,N_24360);
xor U25452 (N_25452,N_24341,N_23920);
and U25453 (N_25453,N_22905,N_24337);
and U25454 (N_25454,N_23868,N_24124);
nor U25455 (N_25455,N_24717,N_24761);
nor U25456 (N_25456,N_23153,N_23362);
nand U25457 (N_25457,N_24647,N_24219);
xnor U25458 (N_25458,N_24605,N_23658);
and U25459 (N_25459,N_24303,N_22881);
nand U25460 (N_25460,N_24826,N_23451);
xnor U25461 (N_25461,N_24167,N_22893);
nand U25462 (N_25462,N_24793,N_24417);
nor U25463 (N_25463,N_24151,N_22755);
and U25464 (N_25464,N_24801,N_24796);
nor U25465 (N_25465,N_22617,N_23219);
xnor U25466 (N_25466,N_24216,N_23653);
and U25467 (N_25467,N_24636,N_23130);
nand U25468 (N_25468,N_22713,N_23567);
nand U25469 (N_25469,N_22909,N_22741);
or U25470 (N_25470,N_23454,N_23854);
xor U25471 (N_25471,N_23885,N_23767);
and U25472 (N_25472,N_24949,N_24655);
and U25473 (N_25473,N_23961,N_24925);
and U25474 (N_25474,N_23998,N_23650);
xnor U25475 (N_25475,N_24461,N_23407);
xnor U25476 (N_25476,N_23595,N_24515);
and U25477 (N_25477,N_23301,N_22934);
nor U25478 (N_25478,N_24881,N_23775);
nor U25479 (N_25479,N_22989,N_23367);
and U25480 (N_25480,N_23871,N_24015);
and U25481 (N_25481,N_23898,N_23630);
or U25482 (N_25482,N_23000,N_22645);
nand U25483 (N_25483,N_22939,N_23188);
and U25484 (N_25484,N_24924,N_24727);
nor U25485 (N_25485,N_22949,N_23142);
nor U25486 (N_25486,N_24463,N_23154);
or U25487 (N_25487,N_23119,N_23824);
and U25488 (N_25488,N_23433,N_24732);
xnor U25489 (N_25489,N_23303,N_23311);
or U25490 (N_25490,N_24901,N_22932);
nor U25491 (N_25491,N_23801,N_23359);
or U25492 (N_25492,N_24821,N_23654);
nor U25493 (N_25493,N_24512,N_23439);
xor U25494 (N_25494,N_23753,N_23011);
or U25495 (N_25495,N_23728,N_24083);
nor U25496 (N_25496,N_24701,N_23769);
and U25497 (N_25497,N_22805,N_22997);
nor U25498 (N_25498,N_24261,N_23968);
and U25499 (N_25499,N_24134,N_24528);
nor U25500 (N_25500,N_23875,N_23181);
nand U25501 (N_25501,N_22808,N_23791);
xor U25502 (N_25502,N_24471,N_22595);
nor U25503 (N_25503,N_23727,N_24191);
nand U25504 (N_25504,N_23773,N_24780);
and U25505 (N_25505,N_24556,N_22556);
or U25506 (N_25506,N_23308,N_24028);
or U25507 (N_25507,N_23641,N_23201);
and U25508 (N_25508,N_24401,N_23987);
and U25509 (N_25509,N_23423,N_23266);
xnor U25510 (N_25510,N_23252,N_22953);
nand U25511 (N_25511,N_24423,N_24311);
xnor U25512 (N_25512,N_24201,N_23251);
nor U25513 (N_25513,N_23804,N_24823);
xnor U25514 (N_25514,N_24215,N_23712);
nand U25515 (N_25515,N_23393,N_24650);
and U25516 (N_25516,N_22501,N_22737);
and U25517 (N_25517,N_23033,N_23835);
or U25518 (N_25518,N_23122,N_24933);
xor U25519 (N_25519,N_23900,N_23892);
and U25520 (N_25520,N_23833,N_22835);
and U25521 (N_25521,N_24968,N_22748);
nand U25522 (N_25522,N_23937,N_23687);
nand U25523 (N_25523,N_23100,N_23028);
nand U25524 (N_25524,N_22655,N_22863);
xor U25525 (N_25525,N_23858,N_23517);
xnor U25526 (N_25526,N_22866,N_22758);
nand U25527 (N_25527,N_22965,N_23376);
xor U25528 (N_25528,N_24657,N_23593);
xor U25529 (N_25529,N_24628,N_23549);
nor U25530 (N_25530,N_24181,N_24427);
nand U25531 (N_25531,N_22764,N_22803);
xor U25532 (N_25532,N_22899,N_22678);
nand U25533 (N_25533,N_24711,N_22738);
nand U25534 (N_25534,N_23363,N_23355);
nand U25535 (N_25535,N_22773,N_24387);
and U25536 (N_25536,N_24059,N_23812);
nand U25537 (N_25537,N_22724,N_23261);
nand U25538 (N_25538,N_22889,N_24376);
or U25539 (N_25539,N_23852,N_23809);
and U25540 (N_25540,N_24958,N_23208);
xnor U25541 (N_25541,N_24849,N_23282);
xnor U25542 (N_25542,N_24754,N_24681);
nand U25543 (N_25543,N_23656,N_24145);
and U25544 (N_25544,N_22579,N_24062);
nor U25545 (N_25545,N_24626,N_24644);
and U25546 (N_25546,N_23992,N_23121);
and U25547 (N_25547,N_23887,N_23710);
nor U25548 (N_25548,N_23669,N_24090);
or U25549 (N_25549,N_24920,N_22892);
and U25550 (N_25550,N_23911,N_24846);
or U25551 (N_25551,N_23356,N_22719);
or U25552 (N_25552,N_24774,N_23247);
and U25553 (N_25553,N_24432,N_24495);
xor U25554 (N_25554,N_23432,N_23366);
and U25555 (N_25555,N_23160,N_24446);
nand U25556 (N_25556,N_24565,N_22821);
xor U25557 (N_25557,N_24093,N_22992);
or U25558 (N_25558,N_23300,N_22914);
xnor U25559 (N_25559,N_22978,N_22936);
or U25560 (N_25560,N_24105,N_23230);
or U25561 (N_25561,N_23861,N_24975);
and U25562 (N_25562,N_24688,N_22628);
nand U25563 (N_25563,N_23422,N_23165);
or U25564 (N_25564,N_23297,N_23636);
and U25565 (N_25565,N_23024,N_24519);
and U25566 (N_25566,N_23411,N_23617);
or U25567 (N_25567,N_23012,N_23256);
nor U25568 (N_25568,N_22666,N_23958);
and U25569 (N_25569,N_23106,N_23232);
or U25570 (N_25570,N_24454,N_23789);
or U25571 (N_25571,N_23632,N_24997);
and U25572 (N_25572,N_24443,N_23682);
xor U25573 (N_25573,N_22879,N_23772);
nand U25574 (N_25574,N_22586,N_24094);
xor U25575 (N_25575,N_22969,N_23702);
xnor U25576 (N_25576,N_23531,N_23347);
nor U25577 (N_25577,N_23304,N_23521);
nor U25578 (N_25578,N_23003,N_23045);
xnor U25579 (N_25579,N_24421,N_24769);
xnor U25580 (N_25580,N_24305,N_24252);
or U25581 (N_25581,N_22552,N_23954);
xor U25582 (N_25582,N_22673,N_23637);
xor U25583 (N_25583,N_23203,N_24567);
nand U25584 (N_25584,N_24749,N_24115);
nor U25585 (N_25585,N_22792,N_22762);
and U25586 (N_25586,N_24424,N_24679);
nand U25587 (N_25587,N_24675,N_24986);
nor U25588 (N_25588,N_22563,N_24668);
or U25589 (N_25589,N_24177,N_23674);
and U25590 (N_25590,N_24706,N_22654);
nand U25591 (N_25591,N_24206,N_23371);
nand U25592 (N_25592,N_24077,N_24704);
nor U25593 (N_25593,N_24898,N_23231);
nand U25594 (N_25594,N_23233,N_22624);
or U25595 (N_25595,N_23587,N_24848);
nand U25596 (N_25596,N_22587,N_24911);
and U25597 (N_25597,N_24651,N_23402);
nand U25598 (N_25598,N_24468,N_24623);
xnor U25599 (N_25599,N_23313,N_24051);
nand U25600 (N_25600,N_23916,N_24023);
or U25601 (N_25601,N_24773,N_24080);
nor U25602 (N_25602,N_22740,N_24331);
nor U25603 (N_25603,N_23336,N_24143);
or U25604 (N_25604,N_23180,N_24102);
or U25605 (N_25605,N_23978,N_22705);
nor U25606 (N_25606,N_22550,N_24127);
and U25607 (N_25607,N_22720,N_23889);
or U25608 (N_25608,N_24054,N_22865);
xor U25609 (N_25609,N_23988,N_24283);
nand U25610 (N_25610,N_23116,N_24718);
or U25611 (N_25611,N_24265,N_23118);
and U25612 (N_25612,N_23612,N_22553);
nor U25613 (N_25613,N_24057,N_23007);
nor U25614 (N_25614,N_23403,N_22813);
xor U25615 (N_25615,N_24113,N_23788);
nor U25616 (N_25616,N_24475,N_22618);
nor U25617 (N_25617,N_24588,N_24168);
or U25618 (N_25618,N_24814,N_24390);
and U25619 (N_25619,N_24349,N_23834);
and U25620 (N_25620,N_23981,N_24482);
or U25621 (N_25621,N_23859,N_23131);
and U25622 (N_25622,N_22999,N_24763);
or U25623 (N_25623,N_22694,N_23755);
nand U25624 (N_25624,N_23221,N_23346);
nand U25625 (N_25625,N_24753,N_22581);
and U25626 (N_25626,N_22777,N_24142);
or U25627 (N_25627,N_24405,N_24694);
nor U25628 (N_25628,N_22629,N_23827);
xor U25629 (N_25629,N_23294,N_23438);
nor U25630 (N_25630,N_23477,N_24099);
or U25631 (N_25631,N_23558,N_24740);
and U25632 (N_25632,N_24660,N_24295);
nand U25633 (N_25633,N_24428,N_24540);
xor U25634 (N_25634,N_22650,N_24163);
nand U25635 (N_25635,N_24779,N_24444);
and U25636 (N_25636,N_24309,N_23114);
nor U25637 (N_25637,N_24953,N_24239);
and U25638 (N_25638,N_23590,N_24347);
and U25639 (N_25639,N_24193,N_24838);
nand U25640 (N_25640,N_24541,N_24744);
nor U25641 (N_25641,N_24334,N_23002);
or U25642 (N_25642,N_23510,N_24490);
or U25643 (N_25643,N_24578,N_22966);
nand U25644 (N_25644,N_24152,N_23964);
and U25645 (N_25645,N_24130,N_22570);
nor U25646 (N_25646,N_24558,N_23348);
or U25647 (N_25647,N_23140,N_24816);
or U25648 (N_25648,N_23502,N_24274);
and U25649 (N_25649,N_23816,N_22747);
nand U25650 (N_25650,N_24904,N_24068);
nor U25651 (N_25651,N_24032,N_24332);
or U25652 (N_25652,N_24162,N_23341);
xnor U25653 (N_25653,N_22971,N_22599);
nor U25654 (N_25654,N_22721,N_22630);
xor U25655 (N_25655,N_22895,N_24030);
nand U25656 (N_25656,N_24076,N_22847);
and U25657 (N_25657,N_23170,N_24600);
nand U25658 (N_25658,N_24368,N_24992);
and U25659 (N_25659,N_22537,N_23972);
nand U25660 (N_25660,N_23613,N_23418);
or U25661 (N_25661,N_22600,N_24687);
nand U25662 (N_25662,N_24211,N_23038);
or U25663 (N_25663,N_23643,N_23873);
or U25664 (N_25664,N_23877,N_22913);
or U25665 (N_25665,N_23563,N_24999);
and U25666 (N_25666,N_24244,N_23864);
or U25667 (N_25667,N_24496,N_23557);
xnor U25668 (N_25668,N_23207,N_24710);
and U25669 (N_25669,N_23700,N_23174);
or U25670 (N_25670,N_24286,N_22988);
nand U25671 (N_25671,N_23708,N_23394);
nor U25672 (N_25672,N_24613,N_22601);
or U25673 (N_25673,N_24132,N_23736);
or U25674 (N_25674,N_22952,N_23392);
nor U25675 (N_25675,N_23584,N_24980);
and U25676 (N_25676,N_22718,N_23723);
nor U25677 (N_25677,N_22656,N_23472);
or U25678 (N_25678,N_23334,N_23524);
or U25679 (N_25679,N_23579,N_24164);
nor U25680 (N_25680,N_24505,N_23026);
and U25681 (N_25681,N_23639,N_22975);
xor U25682 (N_25682,N_23357,N_23015);
nor U25683 (N_25683,N_24601,N_24944);
or U25684 (N_25684,N_24542,N_23737);
nand U25685 (N_25685,N_24374,N_23410);
or U25686 (N_25686,N_23559,N_23618);
and U25687 (N_25687,N_24728,N_24534);
or U25688 (N_25688,N_24784,N_22572);
and U25689 (N_25689,N_23360,N_23945);
nand U25690 (N_25690,N_24971,N_23257);
nor U25691 (N_25691,N_22842,N_23485);
nand U25692 (N_25692,N_23719,N_24695);
nor U25693 (N_25693,N_23550,N_23527);
nor U25694 (N_25694,N_23912,N_24631);
or U25695 (N_25695,N_24149,N_22546);
nor U25696 (N_25696,N_24009,N_24566);
xor U25697 (N_25697,N_22944,N_24692);
nor U25698 (N_25698,N_22697,N_23064);
nor U25699 (N_25699,N_23270,N_23490);
nor U25700 (N_25700,N_24291,N_24696);
nand U25701 (N_25701,N_24036,N_24870);
nand U25702 (N_25702,N_24815,N_24885);
or U25703 (N_25703,N_24316,N_24844);
nor U25704 (N_25704,N_23785,N_24874);
nor U25705 (N_25705,N_24469,N_22513);
or U25706 (N_25706,N_24907,N_22731);
or U25707 (N_25707,N_22974,N_24639);
or U25708 (N_25708,N_24952,N_22793);
xnor U25709 (N_25709,N_23178,N_23361);
and U25710 (N_25710,N_22903,N_24662);
xor U25711 (N_25711,N_24897,N_22545);
nor U25712 (N_25712,N_23846,N_23018);
or U25713 (N_25713,N_23829,N_24736);
and U25714 (N_25714,N_24128,N_23678);
xnor U25715 (N_25715,N_23965,N_22985);
or U25716 (N_25716,N_23776,N_24615);
and U25717 (N_25717,N_24464,N_23511);
and U25718 (N_25718,N_22745,N_24395);
and U25719 (N_25719,N_23057,N_23813);
and U25720 (N_25720,N_24510,N_24433);
xor U25721 (N_25721,N_24373,N_24852);
xnor U25722 (N_25722,N_22942,N_23818);
nor U25723 (N_25723,N_23384,N_23970);
xnor U25724 (N_25724,N_24637,N_24157);
or U25725 (N_25725,N_24109,N_23515);
nand U25726 (N_25726,N_23495,N_24270);
nor U25727 (N_25727,N_23959,N_24297);
nor U25728 (N_25728,N_23735,N_24262);
or U25729 (N_25729,N_24877,N_22711);
nor U25730 (N_25730,N_24320,N_23425);
nor U25731 (N_25731,N_24863,N_23589);
nand U25732 (N_25732,N_24743,N_24762);
nor U25733 (N_25733,N_24802,N_23288);
and U25734 (N_25734,N_23762,N_24854);
or U25735 (N_25735,N_22723,N_23276);
xor U25736 (N_25736,N_24155,N_23025);
xnor U25737 (N_25737,N_23619,N_24220);
nor U25738 (N_25738,N_22503,N_24034);
nand U25739 (N_25739,N_24805,N_24233);
nor U25740 (N_25740,N_23711,N_23315);
or U25741 (N_25741,N_24618,N_24296);
nor U25742 (N_25742,N_23406,N_24537);
nor U25743 (N_25743,N_24758,N_23666);
nor U25744 (N_25744,N_23821,N_23761);
xor U25745 (N_25745,N_23638,N_23874);
nand U25746 (N_25746,N_23309,N_23387);
or U25747 (N_25747,N_23273,N_24066);
and U25748 (N_25748,N_23672,N_24290);
and U25749 (N_25749,N_22787,N_24467);
and U25750 (N_25750,N_22566,N_24620);
xnor U25751 (N_25751,N_23246,N_23196);
and U25752 (N_25752,N_23327,N_22970);
nor U25753 (N_25753,N_24114,N_22910);
nand U25754 (N_25754,N_24358,N_23820);
or U25755 (N_25755,N_22648,N_22882);
or U25756 (N_25756,N_24936,N_22682);
and U25757 (N_25757,N_23382,N_23335);
nand U25758 (N_25758,N_22680,N_24012);
or U25759 (N_25759,N_23268,N_22861);
nand U25760 (N_25760,N_24000,N_22964);
and U25761 (N_25761,N_24661,N_23876);
or U25762 (N_25762,N_24355,N_23338);
and U25763 (N_25763,N_23202,N_22796);
and U25764 (N_25764,N_24470,N_23029);
nor U25765 (N_25765,N_23800,N_22904);
and U25766 (N_25766,N_24707,N_23901);
nand U25767 (N_25767,N_23552,N_24926);
and U25768 (N_25768,N_22674,N_23832);
xor U25769 (N_25769,N_22506,N_24682);
and U25770 (N_25770,N_23662,N_24867);
xnor U25771 (N_25771,N_22636,N_22891);
xnor U25772 (N_25772,N_24103,N_24308);
nand U25773 (N_25773,N_24447,N_24950);
xor U25774 (N_25774,N_24912,N_24314);
nand U25775 (N_25775,N_23278,N_23344);
or U25776 (N_25776,N_24027,N_24379);
or U25777 (N_25777,N_23487,N_23839);
nor U25778 (N_25778,N_24366,N_23155);
xor U25779 (N_25779,N_23168,N_24346);
or U25780 (N_25780,N_23974,N_24321);
xnor U25781 (N_25781,N_24521,N_22643);
nor U25782 (N_25782,N_24243,N_22571);
or U25783 (N_25783,N_23035,N_24697);
and U25784 (N_25784,N_22615,N_23904);
and U25785 (N_25785,N_24782,N_24307);
xnor U25786 (N_25786,N_22921,N_24790);
xnor U25787 (N_25787,N_24449,N_24477);
nand U25788 (N_25788,N_24365,N_24269);
and U25789 (N_25789,N_23113,N_24604);
nand U25790 (N_25790,N_22778,N_24610);
and U25791 (N_25791,N_24498,N_24850);
xnor U25792 (N_25792,N_23893,N_22995);
and U25793 (N_25793,N_23881,N_24722);
xor U25794 (N_25794,N_24487,N_23732);
nor U25795 (N_25795,N_24810,N_24607);
or U25796 (N_25796,N_23431,N_24476);
or U25797 (N_25797,N_24232,N_23888);
or U25798 (N_25798,N_24304,N_24598);
nor U25799 (N_25799,N_22509,N_22689);
and U25800 (N_25800,N_24633,N_23986);
nor U25801 (N_25801,N_24989,N_22691);
xor U25802 (N_25802,N_23867,N_23492);
nand U25803 (N_25803,N_23137,N_23044);
xnor U25804 (N_25804,N_22614,N_24987);
xor U25805 (N_25805,N_24359,N_24794);
xnor U25806 (N_25806,N_24006,N_24225);
xor U25807 (N_25807,N_24812,N_23733);
xnor U25808 (N_25808,N_24894,N_23863);
and U25809 (N_25809,N_24354,N_24016);
or U25810 (N_25810,N_24755,N_24859);
or U25811 (N_25811,N_22649,N_23162);
xnor U25812 (N_25812,N_24529,N_23470);
nand U25813 (N_25813,N_23096,N_23042);
and U25814 (N_25814,N_23481,N_23234);
nor U25815 (N_25815,N_22799,N_24569);
nand U25816 (N_25816,N_24442,N_22549);
and U25817 (N_25817,N_22536,N_24439);
nor U25818 (N_25818,N_24964,N_22757);
nand U25819 (N_25819,N_24967,N_24516);
or U25820 (N_25820,N_23802,N_24878);
and U25821 (N_25821,N_23377,N_24415);
nor U25822 (N_25822,N_24453,N_23169);
xor U25823 (N_25823,N_23646,N_23388);
nor U25824 (N_25824,N_22856,N_23919);
nor U25825 (N_25825,N_23236,N_23091);
nand U25826 (N_25826,N_22852,N_22514);
xnor U25827 (N_25827,N_23040,N_22686);
nand U25828 (N_25828,N_23396,N_24474);
nand U25829 (N_25829,N_23629,N_23980);
nand U25830 (N_25830,N_22804,N_23726);
nand U25831 (N_25831,N_23860,N_23538);
or U25832 (N_25832,N_23097,N_24665);
and U25833 (N_25833,N_23269,N_23110);
nand U25834 (N_25834,N_23242,N_24996);
or U25835 (N_25835,N_22790,N_24187);
xnor U25836 (N_25836,N_23673,N_24136);
nand U25837 (N_25837,N_24910,N_24431);
xor U25838 (N_25838,N_22843,N_24148);
and U25839 (N_25839,N_24778,N_24459);
and U25840 (N_25840,N_24827,N_22765);
or U25841 (N_25841,N_24357,N_23224);
or U25842 (N_25842,N_24768,N_22569);
and U25843 (N_25843,N_23211,N_24873);
nand U25844 (N_25844,N_22840,N_24466);
and U25845 (N_25845,N_23738,N_23459);
nand U25846 (N_25846,N_24572,N_22622);
nand U25847 (N_25847,N_24966,N_23883);
nand U25848 (N_25848,N_24367,N_23507);
xor U25849 (N_25849,N_23546,N_24842);
nor U25850 (N_25850,N_24218,N_23616);
nor U25851 (N_25851,N_23001,N_22770);
or U25852 (N_25852,N_24872,N_22954);
nor U25853 (N_25853,N_24741,N_24654);
or U25854 (N_25854,N_24617,N_22973);
or U25855 (N_25855,N_23977,N_24575);
nor U25856 (N_25856,N_24563,N_24847);
xor U25857 (N_25857,N_24594,N_24491);
nand U25858 (N_25858,N_22739,N_24891);
nor U25859 (N_25859,N_24811,N_24430);
nand U25860 (N_25860,N_24195,N_24238);
nand U25861 (N_25861,N_22972,N_23094);
and U25862 (N_25862,N_23627,N_23158);
xor U25863 (N_25863,N_24643,N_24451);
nor U25864 (N_25864,N_23936,N_23198);
nor U25865 (N_25865,N_24730,N_24001);
xnor U25866 (N_25866,N_22677,N_22877);
xor U25867 (N_25867,N_23023,N_23372);
and U25868 (N_25868,N_24480,N_24640);
xor U25869 (N_25869,N_24280,N_23792);
xor U25870 (N_25870,N_22668,N_22732);
nand U25871 (N_25871,N_24340,N_22885);
or U25872 (N_25872,N_24172,N_24641);
xnor U25873 (N_25873,N_24158,N_22598);
nor U25874 (N_25874,N_23179,N_22661);
or U25875 (N_25875,N_24440,N_23353);
nor U25876 (N_25876,N_24258,N_24264);
xnor U25877 (N_25877,N_24112,N_24413);
and U25878 (N_25878,N_22523,N_22814);
nor U25879 (N_25879,N_23676,N_24052);
or U25880 (N_25880,N_22948,N_23771);
xnor U25881 (N_25881,N_24344,N_22511);
or U25882 (N_25882,N_24025,N_24189);
nor U25883 (N_25883,N_23783,N_22859);
nand U25884 (N_25884,N_24552,N_23528);
nor U25885 (N_25885,N_24546,N_22760);
nor U25886 (N_25886,N_23903,N_24227);
or U25887 (N_25887,N_23417,N_24095);
or U25888 (N_25888,N_22929,N_24100);
or U25889 (N_25889,N_22577,N_22784);
nand U25890 (N_25890,N_23625,N_24147);
and U25891 (N_25891,N_22590,N_24455);
nor U25892 (N_25892,N_23610,N_24335);
nand U25893 (N_25893,N_24918,N_23894);
nand U25894 (N_25894,N_23951,N_23541);
xnor U25895 (N_25895,N_23400,N_22623);
and U25896 (N_25896,N_24896,N_23784);
nand U25897 (N_25897,N_24721,N_23752);
and U25898 (N_25898,N_24834,N_24887);
nand U25899 (N_25899,N_24803,N_22638);
nor U25900 (N_25900,N_24693,N_24301);
and U25901 (N_25901,N_23927,N_24268);
xor U25902 (N_25902,N_23229,N_23626);
nand U25903 (N_25903,N_24514,N_22990);
nand U25904 (N_25904,N_23228,N_23223);
nand U25905 (N_25905,N_24979,N_23184);
or U25906 (N_25906,N_23117,N_23782);
and U25907 (N_25907,N_24257,N_23149);
or U25908 (N_25908,N_24788,N_23831);
nand U25909 (N_25909,N_22809,N_23471);
or U25910 (N_25910,N_24524,N_23177);
and U25911 (N_25911,N_24577,N_23279);
nor U25912 (N_25912,N_22544,N_24900);
nand U25913 (N_25913,N_22798,N_22834);
nor U25914 (N_25914,N_23216,N_23931);
nand U25915 (N_25915,N_22937,N_24050);
nor U25916 (N_25916,N_24079,N_22826);
nor U25917 (N_25917,N_24746,N_23996);
and U25918 (N_25918,N_23983,N_23645);
and U25919 (N_25919,N_23739,N_24317);
xor U25920 (N_25920,N_24589,N_23597);
xor U25921 (N_25921,N_24306,N_22727);
nor U25922 (N_25922,N_22633,N_22957);
nand U25923 (N_25923,N_23530,N_24723);
and U25924 (N_25924,N_23982,N_24509);
nor U25925 (N_25925,N_24713,N_23677);
nor U25926 (N_25926,N_23955,N_23575);
or U25927 (N_25927,N_23729,N_22888);
and U25928 (N_25928,N_22927,N_22653);
nor U25929 (N_25929,N_24760,N_22911);
nand U25930 (N_25930,N_24591,N_24333);
xor U25931 (N_25931,N_23840,N_22853);
nor U25932 (N_25932,N_24893,N_22941);
nor U25933 (N_25933,N_23497,N_24561);
xnor U25934 (N_25934,N_23050,N_23569);
and U25935 (N_25935,N_24786,N_22520);
or U25936 (N_25936,N_23426,N_22644);
or U25937 (N_25937,N_24033,N_22562);
nand U25938 (N_25938,N_22578,N_24154);
or U25939 (N_25939,N_24044,N_22512);
xor U25940 (N_25940,N_22521,N_24678);
xnor U25941 (N_25941,N_23956,N_24666);
or U25942 (N_25942,N_23421,N_24725);
nor U25943 (N_25943,N_23923,N_23999);
or U25944 (N_25944,N_22815,N_24041);
and U25945 (N_25945,N_23902,N_22631);
and U25946 (N_25946,N_24934,N_23369);
nor U25947 (N_25947,N_24084,N_24400);
nand U25948 (N_25948,N_23806,N_23197);
or U25949 (N_25949,N_23004,N_24450);
xnor U25950 (N_25950,N_24748,N_24599);
and U25951 (N_25951,N_23599,N_23187);
nand U25952 (N_25952,N_22593,N_24921);
xor U25953 (N_25953,N_23680,N_24326);
nor U25954 (N_25954,N_24408,N_22551);
nor U25955 (N_25955,N_23295,N_24941);
and U25956 (N_25956,N_24013,N_23148);
nand U25957 (N_25957,N_24798,N_22535);
nand U25958 (N_25958,N_23823,N_24646);
or U25959 (N_25959,N_23109,N_22582);
and U25960 (N_25960,N_24363,N_22735);
nor U25961 (N_25961,N_23060,N_22647);
xnor U25962 (N_25962,N_24315,N_22659);
and U25963 (N_25963,N_23135,N_23333);
or U25964 (N_25964,N_23078,N_23721);
nor U25965 (N_25965,N_24489,N_24568);
xor U25966 (N_25966,N_23032,N_23899);
xnor U25967 (N_25967,N_23343,N_22669);
or U25968 (N_25968,N_24956,N_23628);
nor U25969 (N_25969,N_23803,N_22779);
xnor U25970 (N_25970,N_23555,N_23319);
nand U25971 (N_25971,N_22665,N_23644);
or U25972 (N_25972,N_23855,N_23262);
nand U25973 (N_25973,N_23476,N_23909);
nor U25974 (N_25974,N_24272,N_23544);
nor U25975 (N_25975,N_24855,N_22671);
xnor U25976 (N_25976,N_23048,N_24757);
and U25977 (N_25977,N_23095,N_24535);
nand U25978 (N_25978,N_24576,N_22542);
or U25979 (N_25979,N_23482,N_23560);
xor U25980 (N_25980,N_24325,N_22983);
xnor U25981 (N_25981,N_23866,N_24224);
or U25982 (N_25982,N_23633,N_22860);
and U25983 (N_25983,N_23693,N_22938);
or U25984 (N_25984,N_24671,N_23598);
nor U25985 (N_25985,N_23897,N_24835);
and U25986 (N_25986,N_24864,N_24792);
nor U25987 (N_25987,N_23385,N_22657);
nor U25988 (N_25988,N_24097,N_23022);
or U25989 (N_25989,N_23758,N_23339);
xor U25990 (N_25990,N_23578,N_24254);
or U25991 (N_25991,N_23139,N_23934);
nor U25992 (N_25992,N_24973,N_23283);
xor U25993 (N_25993,N_24392,N_24501);
nor U25994 (N_25994,N_24188,N_23853);
and U25995 (N_25995,N_23150,N_22928);
nor U25996 (N_25996,N_24096,N_23990);
xnor U25997 (N_25997,N_22604,N_24752);
and U25998 (N_25998,N_24214,N_23102);
nand U25999 (N_25999,N_23429,N_22687);
nand U26000 (N_26000,N_23099,N_24554);
xnor U26001 (N_26001,N_23504,N_22887);
nor U26002 (N_26002,N_23455,N_22797);
and U26003 (N_26003,N_23585,N_23370);
nor U26004 (N_26004,N_23793,N_24928);
and U26005 (N_26005,N_23163,N_23647);
nand U26006 (N_26006,N_23566,N_23697);
or U26007 (N_26007,N_22998,N_24795);
nor U26008 (N_26008,N_24407,N_24060);
xnor U26009 (N_26009,N_24945,N_23264);
and U26010 (N_26010,N_24716,N_24983);
nand U26011 (N_26011,N_23080,N_23010);
nor U26012 (N_26012,N_24991,N_23419);
xnor U26013 (N_26013,N_22951,N_23979);
or U26014 (N_26014,N_22524,N_24419);
nand U26015 (N_26015,N_22729,N_23073);
xnor U26016 (N_26016,N_24603,N_24338);
nand U26017 (N_26017,N_23634,N_23543);
nand U26018 (N_26018,N_23631,N_24302);
and U26019 (N_26019,N_24948,N_22568);
nand U26020 (N_26020,N_24073,N_24667);
nor U26021 (N_26021,N_22574,N_23592);
nand U26022 (N_26022,N_23778,N_24452);
nor U26023 (N_26023,N_24042,N_24391);
xor U26024 (N_26024,N_24075,N_23070);
nor U26025 (N_26025,N_24110,N_24583);
or U26026 (N_26026,N_24020,N_22968);
or U26027 (N_26027,N_22611,N_24236);
or U26028 (N_26028,N_24058,N_23603);
xor U26029 (N_26029,N_23478,N_23576);
xor U26030 (N_26030,N_24860,N_23750);
xor U26031 (N_26031,N_24504,N_24411);
and U26032 (N_26032,N_24724,N_23340);
and U26033 (N_26033,N_22869,N_24942);
xnor U26034 (N_26034,N_24397,N_24165);
and U26035 (N_26035,N_22956,N_24021);
xor U26036 (N_26036,N_22560,N_23291);
and U26037 (N_26037,N_23665,N_23079);
xnor U26038 (N_26038,N_22960,N_23845);
nor U26039 (N_26039,N_23440,N_22625);
nand U26040 (N_26040,N_23141,N_24809);
and U26041 (N_26041,N_23065,N_24403);
nor U26042 (N_26042,N_24488,N_24875);
and U26043 (N_26043,N_23914,N_23905);
nand U26044 (N_26044,N_23704,N_23317);
or U26045 (N_26045,N_23913,N_23878);
xor U26046 (N_26046,N_23759,N_23235);
xor U26047 (N_26047,N_24255,N_24853);
or U26048 (N_26048,N_23838,N_22693);
or U26049 (N_26049,N_24362,N_22819);
nor U26050 (N_26050,N_22850,N_24228);
xor U26051 (N_26051,N_23249,N_23756);
nor U26052 (N_26052,N_24292,N_23244);
xor U26053 (N_26053,N_24251,N_23689);
nor U26054 (N_26054,N_23991,N_24674);
nor U26055 (N_26055,N_24412,N_22632);
and U26056 (N_26056,N_24830,N_24008);
and U26057 (N_26057,N_23660,N_24108);
nor U26058 (N_26058,N_23556,N_24836);
nand U26059 (N_26059,N_23798,N_22538);
nor U26060 (N_26060,N_23850,N_24348);
nor U26061 (N_26061,N_23624,N_23540);
and U26062 (N_26062,N_24938,N_23570);
xnor U26063 (N_26063,N_23605,N_24241);
xor U26064 (N_26064,N_24548,N_24698);
xor U26065 (N_26065,N_22641,N_23886);
and U26066 (N_26066,N_23817,N_23960);
and U26067 (N_26067,N_24248,N_24930);
xnor U26068 (N_26068,N_24434,N_22502);
xnor U26069 (N_26069,N_24545,N_24676);
xnor U26070 (N_26070,N_23446,N_22963);
xor U26071 (N_26071,N_23943,N_24551);
nand U26072 (N_26072,N_23498,N_23826);
nor U26073 (N_26073,N_22564,N_23088);
nand U26074 (N_26074,N_22976,N_23399);
nand U26075 (N_26075,N_22967,N_23506);
nand U26076 (N_26076,N_24281,N_22532);
nor U26077 (N_26077,N_22846,N_24494);
and U26078 (N_26078,N_23132,N_23993);
nor U26079 (N_26079,N_22783,N_23745);
nand U26080 (N_26080,N_22875,N_23848);
xor U26081 (N_26081,N_22841,N_23746);
or U26082 (N_26082,N_24845,N_23186);
and U26083 (N_26083,N_24685,N_22701);
nor U26084 (N_26084,N_22690,N_23285);
nand U26085 (N_26085,N_23594,N_22761);
xnor U26086 (N_26086,N_23368,N_23437);
or U26087 (N_26087,N_22996,N_23574);
xnor U26088 (N_26088,N_22811,N_24932);
or U26089 (N_26089,N_23200,N_24284);
xor U26090 (N_26090,N_22763,N_23063);
and U26091 (N_26091,N_23144,N_23932);
xnor U26092 (N_26092,N_24797,N_24624);
xor U26093 (N_26093,N_24963,N_22935);
nor U26094 (N_26094,N_24917,N_23703);
nand U26095 (N_26095,N_22609,N_24581);
nor U26096 (N_26096,N_24544,N_24429);
nor U26097 (N_26097,N_22547,N_24861);
nand U26098 (N_26098,N_22907,N_24074);
or U26099 (N_26099,N_24256,N_24982);
or U26100 (N_26100,N_24889,N_24048);
xor U26101 (N_26101,N_23263,N_23245);
or U26102 (N_26102,N_23715,N_24087);
nor U26103 (N_26103,N_22505,N_24435);
nor U26104 (N_26104,N_24153,N_23675);
and U26105 (N_26105,N_24064,N_24824);
nand U26106 (N_26106,N_23322,N_23087);
nor U26107 (N_26107,N_24070,N_24756);
xnor U26108 (N_26108,N_23124,N_22715);
nor U26109 (N_26109,N_23350,N_23577);
and U26110 (N_26110,N_23051,N_22530);
nor U26111 (N_26111,N_24460,N_23765);
and U26112 (N_26112,N_23237,N_22754);
xor U26113 (N_26113,N_24611,N_24118);
or U26114 (N_26114,N_22930,N_23787);
xor U26115 (N_26115,N_24526,N_23075);
nand U26116 (N_26116,N_24931,N_22886);
or U26117 (N_26117,N_24029,N_23358);
nor U26118 (N_26118,N_24137,N_23810);
nor U26119 (N_26119,N_23797,N_23125);
nor U26120 (N_26120,N_24312,N_22518);
or U26121 (N_26121,N_22695,N_23190);
and U26122 (N_26122,N_24555,N_24731);
xnor U26123 (N_26123,N_24808,N_23655);
xnor U26124 (N_26124,N_22540,N_22940);
and U26125 (N_26125,N_22688,N_23105);
xor U26126 (N_26126,N_22890,N_24388);
or U26127 (N_26127,N_22751,N_23533);
or U26128 (N_26128,N_23963,N_22832);
and U26129 (N_26129,N_23642,N_23331);
and U26130 (N_26130,N_22867,N_23907);
nor U26131 (N_26131,N_24056,N_23349);
xnor U26132 (N_26132,N_23796,N_24977);
and U26133 (N_26133,N_24279,N_23757);
xnor U26134 (N_26134,N_23321,N_22838);
xor U26135 (N_26135,N_23020,N_24658);
xnor U26136 (N_26136,N_23172,N_23192);
nand U26137 (N_26137,N_24649,N_23895);
or U26138 (N_26138,N_23906,N_23036);
nand U26139 (N_26139,N_22707,N_23275);
or U26140 (N_26140,N_24680,N_24619);
or U26141 (N_26141,N_23944,N_24506);
xor U26142 (N_26142,N_24625,N_23606);
nand U26143 (N_26143,N_24876,N_24178);
xor U26144 (N_26144,N_24039,N_23408);
and U26145 (N_26145,N_24122,N_24117);
nand U26146 (N_26146,N_24275,N_23667);
xnor U26147 (N_26147,N_24409,N_23586);
nand U26148 (N_26148,N_24648,N_23434);
nor U26149 (N_26149,N_23479,N_23930);
xnor U26150 (N_26150,N_22962,N_24531);
or U26151 (N_26151,N_23047,N_24298);
nor U26152 (N_26152,N_24369,N_24299);
xnor U26153 (N_26153,N_23841,N_22684);
nor U26154 (N_26154,N_23267,N_24014);
nand U26155 (N_26155,N_24061,N_23008);
xor U26156 (N_26156,N_24426,N_24511);
nand U26157 (N_26157,N_23720,N_22670);
or U26158 (N_26158,N_23571,N_23509);
nor U26159 (N_26159,N_24089,N_24445);
or U26160 (N_26160,N_23622,N_22854);
nand U26161 (N_26161,N_22829,N_23146);
nor U26162 (N_26162,N_22791,N_22709);
and U26163 (N_26163,N_24273,N_23701);
and U26164 (N_26164,N_23962,N_23694);
xnor U26165 (N_26165,N_23463,N_24217);
nor U26166 (N_26166,N_23805,N_24560);
nor U26167 (N_26167,N_23799,N_23734);
and U26168 (N_26168,N_23705,N_23670);
xnor U26169 (N_26169,N_24198,N_23199);
or U26170 (N_26170,N_22824,N_22585);
nor U26171 (N_26171,N_23351,N_23444);
or U26172 (N_26172,N_24294,N_23298);
nor U26173 (N_26173,N_22685,N_22862);
xor U26174 (N_26174,N_23289,N_24879);
or U26175 (N_26175,N_23652,N_22753);
or U26176 (N_26176,N_23725,N_23220);
xor U26177 (N_26177,N_24202,N_24799);
nand U26178 (N_26178,N_23054,N_22902);
xor U26179 (N_26179,N_22728,N_22780);
and U26180 (N_26180,N_23391,N_22662);
xnor U26181 (N_26181,N_22961,N_23443);
nand U26182 (N_26182,N_23565,N_23651);
nor U26183 (N_26183,N_22607,N_23865);
nor U26184 (N_26184,N_22769,N_24530);
nor U26185 (N_26185,N_22639,N_22712);
xor U26186 (N_26186,N_23147,N_24133);
or U26187 (N_26187,N_24422,N_24747);
nand U26188 (N_26188,N_24026,N_23742);
xor U26189 (N_26189,N_24518,N_24043);
xor U26190 (N_26190,N_24974,N_23942);
xnor U26191 (N_26191,N_22794,N_23475);
or U26192 (N_26192,N_23790,N_23770);
and U26193 (N_26193,N_23037,N_23537);
nand U26194 (N_26194,N_24078,N_22696);
nand U26195 (N_26195,N_23777,N_24342);
nor U26196 (N_26196,N_24775,N_22640);
xnor U26197 (N_26197,N_24777,N_23386);
or U26198 (N_26198,N_24197,N_22981);
or U26199 (N_26199,N_24351,N_24040);
and U26200 (N_26200,N_24582,N_22820);
and U26201 (N_26201,N_23474,N_23222);
xor U26202 (N_26202,N_22993,N_24632);
xnor U26203 (N_26203,N_24699,N_23938);
or U26204 (N_26204,N_23107,N_24883);
nand U26205 (N_26205,N_24771,N_24564);
and U26206 (N_26206,N_24038,N_23724);
nor U26207 (N_26207,N_24300,N_22943);
nand U26208 (N_26208,N_24194,N_23922);
xnor U26209 (N_26209,N_23412,N_24880);
and U26210 (N_26210,N_24739,N_23819);
or U26211 (N_26211,N_23468,N_24547);
nor U26212 (N_26212,N_24709,N_22926);
nor U26213 (N_26213,N_22710,N_24947);
or U26214 (N_26214,N_24410,N_24205);
xnor U26215 (N_26215,N_24767,N_23072);
nand U26216 (N_26216,N_24819,N_23157);
and U26217 (N_26217,N_23910,N_23522);
or U26218 (N_26218,N_24553,N_24161);
and U26219 (N_26219,N_23814,N_24377);
nor U26220 (N_26220,N_23209,N_23503);
nor U26221 (N_26221,N_23084,N_24436);
or U26222 (N_26222,N_24500,N_23414);
or U26223 (N_26223,N_23016,N_24614);
nor U26224 (N_26224,N_24905,N_24902);
nand U26225 (N_26225,N_24998,N_23458);
nor U26226 (N_26226,N_24011,N_23763);
xnor U26227 (N_26227,N_23337,N_24210);
nor U26228 (N_26228,N_22901,N_24765);
nand U26229 (N_26229,N_24017,N_23591);
and U26230 (N_26230,N_24585,N_24807);
xnor U26231 (N_26231,N_23098,N_22759);
or U26232 (N_26232,N_24737,N_22734);
xor U26233 (N_26233,N_23489,N_24622);
nor U26234 (N_26234,N_24645,N_24037);
or U26235 (N_26235,N_24684,N_23166);
or U26236 (N_26236,N_23532,N_23296);
xnor U26237 (N_26237,N_24107,N_22621);
or U26238 (N_26238,N_23851,N_23896);
or U26239 (N_26239,N_24343,N_24483);
or U26240 (N_26240,N_23194,N_24691);
or U26241 (N_26241,N_24196,N_23254);
or U26242 (N_26242,N_24937,N_23949);
xnor U26243 (N_26243,N_23779,N_24212);
xnor U26244 (N_26244,N_22602,N_23714);
and U26245 (N_26245,N_22519,N_22534);
nand U26246 (N_26246,N_24726,N_24288);
nor U26247 (N_26247,N_22605,N_24916);
nand U26248 (N_26248,N_24825,N_22736);
or U26249 (N_26249,N_23253,N_24612);
xnor U26250 (N_26250,N_23650,N_24254);
or U26251 (N_26251,N_24017,N_22958);
and U26252 (N_26252,N_24814,N_22926);
or U26253 (N_26253,N_24285,N_24623);
xnor U26254 (N_26254,N_23909,N_24934);
nand U26255 (N_26255,N_23680,N_22894);
nand U26256 (N_26256,N_24367,N_23438);
or U26257 (N_26257,N_22935,N_23774);
nor U26258 (N_26258,N_24315,N_23327);
nand U26259 (N_26259,N_24560,N_24743);
and U26260 (N_26260,N_23033,N_23393);
xor U26261 (N_26261,N_24303,N_24570);
and U26262 (N_26262,N_24731,N_23944);
xor U26263 (N_26263,N_22805,N_24089);
nor U26264 (N_26264,N_23111,N_23627);
xnor U26265 (N_26265,N_23649,N_22965);
and U26266 (N_26266,N_23458,N_23004);
nand U26267 (N_26267,N_23111,N_24009);
xnor U26268 (N_26268,N_23961,N_22976);
and U26269 (N_26269,N_23485,N_22500);
xor U26270 (N_26270,N_23786,N_22761);
and U26271 (N_26271,N_24973,N_22894);
xnor U26272 (N_26272,N_23939,N_23591);
and U26273 (N_26273,N_24938,N_24516);
and U26274 (N_26274,N_24552,N_23092);
nand U26275 (N_26275,N_24416,N_24724);
xnor U26276 (N_26276,N_24619,N_24954);
xor U26277 (N_26277,N_22827,N_23244);
or U26278 (N_26278,N_23518,N_24262);
xnor U26279 (N_26279,N_23062,N_24473);
or U26280 (N_26280,N_24708,N_23614);
nor U26281 (N_26281,N_24958,N_24288);
or U26282 (N_26282,N_22884,N_24494);
nor U26283 (N_26283,N_23864,N_24225);
or U26284 (N_26284,N_24706,N_24473);
nand U26285 (N_26285,N_23560,N_22555);
and U26286 (N_26286,N_24460,N_22982);
nor U26287 (N_26287,N_24233,N_23008);
nand U26288 (N_26288,N_22584,N_24659);
nor U26289 (N_26289,N_22980,N_24144);
and U26290 (N_26290,N_22980,N_24184);
xnor U26291 (N_26291,N_22710,N_24570);
nand U26292 (N_26292,N_22632,N_23951);
nand U26293 (N_26293,N_24811,N_23931);
and U26294 (N_26294,N_23393,N_24825);
nor U26295 (N_26295,N_23087,N_23826);
nand U26296 (N_26296,N_23443,N_23624);
nand U26297 (N_26297,N_22866,N_23364);
and U26298 (N_26298,N_24869,N_23203);
nand U26299 (N_26299,N_23556,N_24113);
nand U26300 (N_26300,N_24054,N_22987);
and U26301 (N_26301,N_23983,N_23359);
or U26302 (N_26302,N_23159,N_22558);
nor U26303 (N_26303,N_23397,N_24321);
nor U26304 (N_26304,N_23395,N_24357);
xor U26305 (N_26305,N_24846,N_24001);
and U26306 (N_26306,N_23672,N_24938);
nor U26307 (N_26307,N_22814,N_23036);
nor U26308 (N_26308,N_22764,N_24868);
nor U26309 (N_26309,N_23300,N_22998);
nand U26310 (N_26310,N_23505,N_24919);
xor U26311 (N_26311,N_24134,N_22971);
nand U26312 (N_26312,N_22848,N_23397);
and U26313 (N_26313,N_23818,N_23551);
or U26314 (N_26314,N_23808,N_22579);
and U26315 (N_26315,N_23941,N_22541);
or U26316 (N_26316,N_24387,N_23507);
nor U26317 (N_26317,N_24627,N_24666);
nand U26318 (N_26318,N_23473,N_24151);
nand U26319 (N_26319,N_24594,N_24202);
nand U26320 (N_26320,N_24884,N_22714);
or U26321 (N_26321,N_22736,N_22764);
nor U26322 (N_26322,N_23147,N_24364);
nor U26323 (N_26323,N_23651,N_23357);
or U26324 (N_26324,N_23241,N_24584);
xnor U26325 (N_26325,N_24749,N_23717);
xnor U26326 (N_26326,N_23000,N_23918);
nor U26327 (N_26327,N_24339,N_23827);
xor U26328 (N_26328,N_23965,N_24630);
or U26329 (N_26329,N_24558,N_23744);
nor U26330 (N_26330,N_24255,N_23384);
and U26331 (N_26331,N_24991,N_24639);
or U26332 (N_26332,N_24981,N_24178);
nor U26333 (N_26333,N_23211,N_24123);
nor U26334 (N_26334,N_23719,N_23074);
and U26335 (N_26335,N_24101,N_24082);
nor U26336 (N_26336,N_23275,N_23757);
or U26337 (N_26337,N_24699,N_23237);
xnor U26338 (N_26338,N_22821,N_24932);
or U26339 (N_26339,N_22835,N_24159);
xor U26340 (N_26340,N_24086,N_22690);
and U26341 (N_26341,N_23762,N_23076);
nor U26342 (N_26342,N_23661,N_24348);
nand U26343 (N_26343,N_24367,N_24006);
xor U26344 (N_26344,N_24066,N_23043);
and U26345 (N_26345,N_23427,N_23457);
nand U26346 (N_26346,N_24054,N_23327);
nor U26347 (N_26347,N_24670,N_23695);
and U26348 (N_26348,N_24149,N_22710);
or U26349 (N_26349,N_24837,N_24316);
nor U26350 (N_26350,N_23164,N_23069);
nand U26351 (N_26351,N_24221,N_23344);
xor U26352 (N_26352,N_23916,N_24679);
or U26353 (N_26353,N_22909,N_23753);
and U26354 (N_26354,N_24383,N_23549);
and U26355 (N_26355,N_23301,N_24606);
or U26356 (N_26356,N_23252,N_24179);
xnor U26357 (N_26357,N_24489,N_23673);
or U26358 (N_26358,N_24001,N_23060);
nor U26359 (N_26359,N_23530,N_23390);
nor U26360 (N_26360,N_23307,N_23027);
nand U26361 (N_26361,N_24506,N_24752);
xor U26362 (N_26362,N_23226,N_22904);
nor U26363 (N_26363,N_24627,N_22672);
and U26364 (N_26364,N_22509,N_23398);
nor U26365 (N_26365,N_22692,N_23486);
xor U26366 (N_26366,N_23438,N_23031);
nand U26367 (N_26367,N_23595,N_24022);
and U26368 (N_26368,N_22963,N_23699);
nand U26369 (N_26369,N_24317,N_23309);
and U26370 (N_26370,N_24003,N_24154);
nand U26371 (N_26371,N_22592,N_22887);
xnor U26372 (N_26372,N_24875,N_24948);
nor U26373 (N_26373,N_23177,N_23113);
and U26374 (N_26374,N_24012,N_24194);
nand U26375 (N_26375,N_23569,N_23529);
nand U26376 (N_26376,N_22811,N_24227);
and U26377 (N_26377,N_24124,N_24451);
xor U26378 (N_26378,N_22786,N_23308);
and U26379 (N_26379,N_24001,N_24314);
nor U26380 (N_26380,N_23313,N_24224);
nor U26381 (N_26381,N_23429,N_24933);
and U26382 (N_26382,N_22967,N_24259);
xor U26383 (N_26383,N_22998,N_24059);
nor U26384 (N_26384,N_23059,N_24150);
nand U26385 (N_26385,N_23108,N_23953);
xor U26386 (N_26386,N_23013,N_23448);
and U26387 (N_26387,N_23504,N_22972);
nor U26388 (N_26388,N_23427,N_23100);
or U26389 (N_26389,N_24374,N_23963);
xnor U26390 (N_26390,N_23317,N_24666);
nor U26391 (N_26391,N_22804,N_22911);
and U26392 (N_26392,N_24058,N_23948);
or U26393 (N_26393,N_22518,N_22987);
or U26394 (N_26394,N_23718,N_22999);
or U26395 (N_26395,N_24684,N_24734);
xor U26396 (N_26396,N_23015,N_22612);
and U26397 (N_26397,N_22852,N_24850);
nand U26398 (N_26398,N_23711,N_24735);
or U26399 (N_26399,N_22949,N_24084);
nor U26400 (N_26400,N_22851,N_23489);
nor U26401 (N_26401,N_23650,N_23443);
nand U26402 (N_26402,N_22633,N_23556);
nand U26403 (N_26403,N_24946,N_24432);
nor U26404 (N_26404,N_22685,N_23899);
nand U26405 (N_26405,N_24734,N_24533);
or U26406 (N_26406,N_24873,N_23768);
nand U26407 (N_26407,N_24126,N_22735);
nor U26408 (N_26408,N_24079,N_23626);
xnor U26409 (N_26409,N_24111,N_23039);
nand U26410 (N_26410,N_24059,N_23916);
nand U26411 (N_26411,N_24128,N_22835);
or U26412 (N_26412,N_24373,N_24684);
xor U26413 (N_26413,N_23415,N_24887);
nor U26414 (N_26414,N_23484,N_23899);
or U26415 (N_26415,N_24887,N_23679);
or U26416 (N_26416,N_23431,N_23078);
nor U26417 (N_26417,N_24321,N_22995);
xnor U26418 (N_26418,N_24210,N_24139);
nor U26419 (N_26419,N_24308,N_24021);
or U26420 (N_26420,N_22730,N_24082);
nand U26421 (N_26421,N_22707,N_23330);
xnor U26422 (N_26422,N_23039,N_24163);
and U26423 (N_26423,N_24636,N_23924);
and U26424 (N_26424,N_22637,N_22517);
nor U26425 (N_26425,N_24639,N_24350);
nand U26426 (N_26426,N_22969,N_23740);
nor U26427 (N_26427,N_24039,N_23156);
nand U26428 (N_26428,N_23249,N_23155);
nand U26429 (N_26429,N_23319,N_22647);
nand U26430 (N_26430,N_22617,N_22532);
nand U26431 (N_26431,N_22974,N_23285);
or U26432 (N_26432,N_23303,N_24218);
or U26433 (N_26433,N_23480,N_24404);
nor U26434 (N_26434,N_23717,N_24420);
or U26435 (N_26435,N_24240,N_23236);
xor U26436 (N_26436,N_24036,N_22769);
and U26437 (N_26437,N_23101,N_24681);
nor U26438 (N_26438,N_22858,N_23578);
and U26439 (N_26439,N_22772,N_23097);
and U26440 (N_26440,N_23324,N_24270);
and U26441 (N_26441,N_23096,N_24432);
nand U26442 (N_26442,N_23724,N_22835);
or U26443 (N_26443,N_23302,N_23549);
or U26444 (N_26444,N_23621,N_22935);
nand U26445 (N_26445,N_23333,N_22958);
and U26446 (N_26446,N_24738,N_23162);
nor U26447 (N_26447,N_24740,N_24936);
xnor U26448 (N_26448,N_23675,N_24599);
xnor U26449 (N_26449,N_24740,N_24945);
or U26450 (N_26450,N_22966,N_24138);
nor U26451 (N_26451,N_22768,N_24016);
nor U26452 (N_26452,N_24899,N_24518);
nor U26453 (N_26453,N_23498,N_22801);
and U26454 (N_26454,N_22956,N_23059);
nand U26455 (N_26455,N_24554,N_24760);
and U26456 (N_26456,N_22921,N_23528);
xor U26457 (N_26457,N_23717,N_22854);
nor U26458 (N_26458,N_24907,N_23380);
or U26459 (N_26459,N_24061,N_24352);
nand U26460 (N_26460,N_24406,N_23902);
or U26461 (N_26461,N_24078,N_23423);
xor U26462 (N_26462,N_23537,N_24068);
and U26463 (N_26463,N_24567,N_22787);
and U26464 (N_26464,N_23608,N_23474);
and U26465 (N_26465,N_23752,N_24391);
xnor U26466 (N_26466,N_22850,N_23376);
or U26467 (N_26467,N_22696,N_23848);
and U26468 (N_26468,N_23329,N_23334);
xor U26469 (N_26469,N_23350,N_24815);
or U26470 (N_26470,N_22661,N_23976);
nor U26471 (N_26471,N_23484,N_24797);
nor U26472 (N_26472,N_22825,N_24942);
and U26473 (N_26473,N_24379,N_23073);
or U26474 (N_26474,N_22774,N_23994);
nand U26475 (N_26475,N_24128,N_22899);
and U26476 (N_26476,N_24567,N_23876);
nor U26477 (N_26477,N_24521,N_24327);
and U26478 (N_26478,N_24365,N_23918);
and U26479 (N_26479,N_22526,N_23952);
xor U26480 (N_26480,N_22884,N_22822);
xnor U26481 (N_26481,N_24748,N_22760);
xor U26482 (N_26482,N_23478,N_22639);
xor U26483 (N_26483,N_24503,N_23802);
nor U26484 (N_26484,N_22823,N_23330);
nand U26485 (N_26485,N_23758,N_23849);
and U26486 (N_26486,N_23298,N_22804);
xor U26487 (N_26487,N_24904,N_24979);
nand U26488 (N_26488,N_23086,N_22902);
or U26489 (N_26489,N_23453,N_24901);
nand U26490 (N_26490,N_24613,N_24170);
and U26491 (N_26491,N_23884,N_23718);
or U26492 (N_26492,N_23959,N_24867);
nand U26493 (N_26493,N_22619,N_22757);
xnor U26494 (N_26494,N_23540,N_24887);
and U26495 (N_26495,N_22765,N_23307);
xor U26496 (N_26496,N_22694,N_23139);
nand U26497 (N_26497,N_24279,N_24421);
and U26498 (N_26498,N_24569,N_23003);
or U26499 (N_26499,N_24935,N_24689);
and U26500 (N_26500,N_23548,N_24498);
nand U26501 (N_26501,N_24341,N_23747);
and U26502 (N_26502,N_22652,N_24023);
nand U26503 (N_26503,N_23704,N_22966);
or U26504 (N_26504,N_23727,N_24537);
nor U26505 (N_26505,N_24930,N_24330);
or U26506 (N_26506,N_22775,N_24455);
nand U26507 (N_26507,N_24077,N_22676);
nor U26508 (N_26508,N_22947,N_23120);
nand U26509 (N_26509,N_23835,N_24689);
nand U26510 (N_26510,N_23962,N_24136);
and U26511 (N_26511,N_23268,N_22784);
nor U26512 (N_26512,N_22828,N_23638);
or U26513 (N_26513,N_23970,N_24082);
and U26514 (N_26514,N_22915,N_23223);
and U26515 (N_26515,N_23107,N_22632);
xnor U26516 (N_26516,N_24895,N_22934);
and U26517 (N_26517,N_22999,N_23950);
and U26518 (N_26518,N_23045,N_24508);
and U26519 (N_26519,N_24098,N_23234);
nor U26520 (N_26520,N_23292,N_22685);
or U26521 (N_26521,N_24813,N_23977);
and U26522 (N_26522,N_23691,N_23419);
or U26523 (N_26523,N_23191,N_23320);
xor U26524 (N_26524,N_24696,N_23771);
and U26525 (N_26525,N_23081,N_22553);
nor U26526 (N_26526,N_23332,N_23430);
xnor U26527 (N_26527,N_23226,N_24120);
xor U26528 (N_26528,N_23465,N_22531);
xor U26529 (N_26529,N_23788,N_24611);
nor U26530 (N_26530,N_23424,N_24737);
nor U26531 (N_26531,N_24733,N_24179);
nor U26532 (N_26532,N_24896,N_22768);
nor U26533 (N_26533,N_22616,N_24510);
nor U26534 (N_26534,N_23684,N_22575);
xnor U26535 (N_26535,N_24931,N_24421);
nand U26536 (N_26536,N_23285,N_24109);
xnor U26537 (N_26537,N_23901,N_23078);
nand U26538 (N_26538,N_23989,N_23187);
or U26539 (N_26539,N_23905,N_24322);
or U26540 (N_26540,N_23190,N_24180);
nor U26541 (N_26541,N_24849,N_22515);
and U26542 (N_26542,N_23045,N_23238);
nor U26543 (N_26543,N_23550,N_22819);
and U26544 (N_26544,N_23481,N_24545);
or U26545 (N_26545,N_23644,N_22673);
xnor U26546 (N_26546,N_24236,N_24590);
or U26547 (N_26547,N_22722,N_24987);
or U26548 (N_26548,N_22699,N_22785);
and U26549 (N_26549,N_23580,N_23727);
nand U26550 (N_26550,N_23278,N_24559);
or U26551 (N_26551,N_23904,N_23978);
nand U26552 (N_26552,N_22762,N_24853);
xor U26553 (N_26553,N_23779,N_23462);
or U26554 (N_26554,N_23718,N_22854);
xor U26555 (N_26555,N_23281,N_22863);
xnor U26556 (N_26556,N_24867,N_23124);
xor U26557 (N_26557,N_22596,N_24398);
xnor U26558 (N_26558,N_23303,N_23491);
and U26559 (N_26559,N_24096,N_23774);
nand U26560 (N_26560,N_22519,N_22961);
and U26561 (N_26561,N_24827,N_23962);
nand U26562 (N_26562,N_22975,N_24404);
nand U26563 (N_26563,N_24082,N_23035);
xnor U26564 (N_26564,N_23047,N_23876);
nand U26565 (N_26565,N_24526,N_23084);
nand U26566 (N_26566,N_24973,N_22715);
and U26567 (N_26567,N_23487,N_22803);
and U26568 (N_26568,N_24061,N_23860);
nor U26569 (N_26569,N_23808,N_24400);
and U26570 (N_26570,N_23072,N_23406);
nand U26571 (N_26571,N_23536,N_24626);
and U26572 (N_26572,N_24918,N_23308);
xor U26573 (N_26573,N_23097,N_23239);
or U26574 (N_26574,N_24261,N_23886);
nor U26575 (N_26575,N_24630,N_23121);
nand U26576 (N_26576,N_24568,N_24977);
nand U26577 (N_26577,N_24336,N_22701);
or U26578 (N_26578,N_23255,N_22773);
xnor U26579 (N_26579,N_24022,N_24788);
xnor U26580 (N_26580,N_22796,N_24336);
nor U26581 (N_26581,N_24470,N_23138);
nand U26582 (N_26582,N_23167,N_22641);
nor U26583 (N_26583,N_22755,N_23966);
xnor U26584 (N_26584,N_24236,N_23347);
or U26585 (N_26585,N_24077,N_22979);
xor U26586 (N_26586,N_23124,N_24732);
nor U26587 (N_26587,N_22671,N_24029);
or U26588 (N_26588,N_24312,N_24021);
xnor U26589 (N_26589,N_24699,N_23107);
nor U26590 (N_26590,N_24589,N_24677);
and U26591 (N_26591,N_24140,N_22981);
and U26592 (N_26592,N_23115,N_24286);
nor U26593 (N_26593,N_24293,N_22651);
and U26594 (N_26594,N_23183,N_23304);
nor U26595 (N_26595,N_24923,N_24124);
nand U26596 (N_26596,N_24510,N_24475);
xor U26597 (N_26597,N_23188,N_23133);
xor U26598 (N_26598,N_23839,N_24981);
nand U26599 (N_26599,N_24528,N_24873);
or U26600 (N_26600,N_23949,N_24976);
nand U26601 (N_26601,N_24535,N_23043);
or U26602 (N_26602,N_22770,N_22842);
nand U26603 (N_26603,N_24784,N_23216);
nor U26604 (N_26604,N_22815,N_23796);
and U26605 (N_26605,N_24923,N_23921);
or U26606 (N_26606,N_23432,N_24640);
and U26607 (N_26607,N_24431,N_24252);
or U26608 (N_26608,N_23916,N_23875);
or U26609 (N_26609,N_24487,N_22997);
nor U26610 (N_26610,N_23644,N_23920);
nand U26611 (N_26611,N_24375,N_23444);
nand U26612 (N_26612,N_24005,N_23562);
nand U26613 (N_26613,N_23417,N_23173);
or U26614 (N_26614,N_24947,N_23210);
nor U26615 (N_26615,N_24153,N_24462);
and U26616 (N_26616,N_24223,N_23856);
or U26617 (N_26617,N_24602,N_24801);
nand U26618 (N_26618,N_24468,N_23796);
and U26619 (N_26619,N_24135,N_22611);
and U26620 (N_26620,N_23908,N_22616);
nand U26621 (N_26621,N_23856,N_22557);
nor U26622 (N_26622,N_24493,N_24668);
nor U26623 (N_26623,N_24223,N_22511);
nand U26624 (N_26624,N_23724,N_22525);
or U26625 (N_26625,N_24454,N_23810);
xor U26626 (N_26626,N_22817,N_23964);
or U26627 (N_26627,N_23124,N_23085);
nand U26628 (N_26628,N_23117,N_23020);
nand U26629 (N_26629,N_24278,N_24930);
or U26630 (N_26630,N_24128,N_23105);
or U26631 (N_26631,N_23722,N_23436);
nand U26632 (N_26632,N_22575,N_24365);
nor U26633 (N_26633,N_24503,N_23289);
xor U26634 (N_26634,N_24324,N_23496);
xor U26635 (N_26635,N_24787,N_24061);
and U26636 (N_26636,N_22584,N_24441);
nor U26637 (N_26637,N_24499,N_23509);
xnor U26638 (N_26638,N_24530,N_24712);
nor U26639 (N_26639,N_24730,N_24799);
xnor U26640 (N_26640,N_23207,N_22729);
nand U26641 (N_26641,N_23957,N_24486);
xor U26642 (N_26642,N_23194,N_23251);
xnor U26643 (N_26643,N_22653,N_23835);
nand U26644 (N_26644,N_24698,N_23889);
nand U26645 (N_26645,N_22930,N_22833);
nor U26646 (N_26646,N_24056,N_23516);
nand U26647 (N_26647,N_23440,N_24297);
xnor U26648 (N_26648,N_24419,N_24714);
xor U26649 (N_26649,N_24144,N_23578);
nand U26650 (N_26650,N_24267,N_22555);
nor U26651 (N_26651,N_24906,N_22829);
nand U26652 (N_26652,N_24570,N_23274);
or U26653 (N_26653,N_22874,N_23869);
and U26654 (N_26654,N_23249,N_23737);
and U26655 (N_26655,N_23226,N_23186);
and U26656 (N_26656,N_22794,N_22748);
nor U26657 (N_26657,N_24268,N_24054);
nand U26658 (N_26658,N_23631,N_22777);
nand U26659 (N_26659,N_24635,N_24860);
xor U26660 (N_26660,N_24016,N_22549);
xnor U26661 (N_26661,N_23301,N_23711);
or U26662 (N_26662,N_23817,N_24907);
or U26663 (N_26663,N_23929,N_23789);
xnor U26664 (N_26664,N_24472,N_22593);
xor U26665 (N_26665,N_22771,N_23906);
nor U26666 (N_26666,N_24922,N_22966);
nand U26667 (N_26667,N_23085,N_24683);
or U26668 (N_26668,N_23794,N_24398);
nor U26669 (N_26669,N_24745,N_23498);
nor U26670 (N_26670,N_23569,N_22683);
and U26671 (N_26671,N_24373,N_23154);
xnor U26672 (N_26672,N_24753,N_23565);
nor U26673 (N_26673,N_24163,N_24249);
or U26674 (N_26674,N_22777,N_23419);
or U26675 (N_26675,N_23467,N_24917);
nor U26676 (N_26676,N_23377,N_24307);
and U26677 (N_26677,N_23273,N_24015);
nand U26678 (N_26678,N_24007,N_24935);
nand U26679 (N_26679,N_24298,N_22593);
nand U26680 (N_26680,N_24945,N_23092);
xnor U26681 (N_26681,N_22976,N_23586);
nor U26682 (N_26682,N_24104,N_23200);
and U26683 (N_26683,N_22508,N_24157);
xnor U26684 (N_26684,N_24070,N_24408);
nand U26685 (N_26685,N_24354,N_23469);
nor U26686 (N_26686,N_23320,N_23238);
or U26687 (N_26687,N_24432,N_24283);
and U26688 (N_26688,N_24203,N_24680);
or U26689 (N_26689,N_23719,N_23312);
and U26690 (N_26690,N_24953,N_23308);
nand U26691 (N_26691,N_23468,N_22761);
nand U26692 (N_26692,N_23560,N_23459);
nand U26693 (N_26693,N_23173,N_24436);
xnor U26694 (N_26694,N_23698,N_23004);
nand U26695 (N_26695,N_23614,N_24570);
xor U26696 (N_26696,N_22616,N_22917);
xnor U26697 (N_26697,N_24531,N_24368);
and U26698 (N_26698,N_23348,N_22769);
or U26699 (N_26699,N_22514,N_23317);
and U26700 (N_26700,N_22965,N_23084);
nand U26701 (N_26701,N_24438,N_24290);
or U26702 (N_26702,N_22570,N_23195);
xor U26703 (N_26703,N_24225,N_23525);
and U26704 (N_26704,N_24091,N_24480);
or U26705 (N_26705,N_23887,N_24032);
xor U26706 (N_26706,N_24143,N_22612);
or U26707 (N_26707,N_23654,N_22970);
or U26708 (N_26708,N_23405,N_22522);
or U26709 (N_26709,N_23326,N_24745);
and U26710 (N_26710,N_23754,N_24994);
nand U26711 (N_26711,N_22664,N_22643);
and U26712 (N_26712,N_23889,N_24155);
nor U26713 (N_26713,N_23070,N_24912);
or U26714 (N_26714,N_23343,N_24278);
and U26715 (N_26715,N_22799,N_23506);
xnor U26716 (N_26716,N_23148,N_23806);
and U26717 (N_26717,N_23529,N_22775);
and U26718 (N_26718,N_23256,N_22727);
and U26719 (N_26719,N_24990,N_24529);
and U26720 (N_26720,N_24424,N_22672);
nor U26721 (N_26721,N_23783,N_22641);
nand U26722 (N_26722,N_24087,N_22592);
xnor U26723 (N_26723,N_24393,N_24746);
xor U26724 (N_26724,N_24963,N_24206);
xnor U26725 (N_26725,N_23995,N_23199);
xor U26726 (N_26726,N_24969,N_22638);
nor U26727 (N_26727,N_24158,N_24586);
or U26728 (N_26728,N_23219,N_24838);
and U26729 (N_26729,N_23870,N_24059);
or U26730 (N_26730,N_24522,N_22754);
nand U26731 (N_26731,N_22892,N_23275);
nor U26732 (N_26732,N_24330,N_23657);
nand U26733 (N_26733,N_24940,N_23094);
or U26734 (N_26734,N_22971,N_23582);
nand U26735 (N_26735,N_24853,N_24628);
nand U26736 (N_26736,N_23080,N_22820);
xnor U26737 (N_26737,N_22888,N_23078);
and U26738 (N_26738,N_24818,N_23161);
nand U26739 (N_26739,N_23869,N_24221);
and U26740 (N_26740,N_24064,N_23463);
and U26741 (N_26741,N_22527,N_23448);
or U26742 (N_26742,N_24390,N_23138);
nor U26743 (N_26743,N_24295,N_22885);
xnor U26744 (N_26744,N_24625,N_23819);
and U26745 (N_26745,N_23104,N_23429);
and U26746 (N_26746,N_24467,N_23867);
xor U26747 (N_26747,N_23819,N_24448);
nor U26748 (N_26748,N_24376,N_23382);
nand U26749 (N_26749,N_23690,N_23423);
nand U26750 (N_26750,N_23859,N_24595);
and U26751 (N_26751,N_23368,N_23471);
nor U26752 (N_26752,N_22824,N_23023);
nand U26753 (N_26753,N_24640,N_23229);
nor U26754 (N_26754,N_24892,N_22902);
and U26755 (N_26755,N_22865,N_23655);
and U26756 (N_26756,N_24731,N_23135);
nor U26757 (N_26757,N_23944,N_23662);
or U26758 (N_26758,N_24240,N_23547);
nand U26759 (N_26759,N_24448,N_22856);
nand U26760 (N_26760,N_23790,N_22599);
nand U26761 (N_26761,N_23807,N_23010);
xnor U26762 (N_26762,N_24758,N_23817);
xnor U26763 (N_26763,N_23356,N_23331);
xnor U26764 (N_26764,N_24418,N_24539);
xnor U26765 (N_26765,N_22664,N_24972);
xnor U26766 (N_26766,N_22556,N_22566);
or U26767 (N_26767,N_22583,N_23955);
nor U26768 (N_26768,N_22559,N_23334);
nor U26769 (N_26769,N_23533,N_24766);
xor U26770 (N_26770,N_23707,N_23332);
and U26771 (N_26771,N_24480,N_23360);
and U26772 (N_26772,N_23670,N_24011);
or U26773 (N_26773,N_23724,N_22522);
and U26774 (N_26774,N_24524,N_23846);
and U26775 (N_26775,N_24253,N_23790);
nor U26776 (N_26776,N_23089,N_24309);
and U26777 (N_26777,N_24839,N_24450);
nand U26778 (N_26778,N_24443,N_23385);
and U26779 (N_26779,N_24469,N_22503);
nand U26780 (N_26780,N_23276,N_24532);
and U26781 (N_26781,N_24158,N_23084);
nor U26782 (N_26782,N_22751,N_22930);
and U26783 (N_26783,N_23279,N_24814);
and U26784 (N_26784,N_23999,N_24428);
nor U26785 (N_26785,N_24875,N_24859);
nor U26786 (N_26786,N_24874,N_23246);
nand U26787 (N_26787,N_23263,N_23942);
nor U26788 (N_26788,N_23735,N_24550);
or U26789 (N_26789,N_24197,N_23316);
or U26790 (N_26790,N_22865,N_22758);
xor U26791 (N_26791,N_24024,N_22603);
and U26792 (N_26792,N_23918,N_23838);
xnor U26793 (N_26793,N_23167,N_23086);
and U26794 (N_26794,N_23404,N_22797);
nor U26795 (N_26795,N_23896,N_24188);
nor U26796 (N_26796,N_24896,N_24535);
nor U26797 (N_26797,N_24898,N_23336);
and U26798 (N_26798,N_22828,N_24395);
nor U26799 (N_26799,N_23638,N_23443);
nor U26800 (N_26800,N_24234,N_24662);
and U26801 (N_26801,N_23954,N_23256);
or U26802 (N_26802,N_23357,N_23029);
nand U26803 (N_26803,N_22538,N_23957);
nor U26804 (N_26804,N_24053,N_22802);
and U26805 (N_26805,N_24110,N_22598);
nand U26806 (N_26806,N_24101,N_23780);
nand U26807 (N_26807,N_23862,N_22758);
nand U26808 (N_26808,N_24227,N_22872);
or U26809 (N_26809,N_22531,N_22537);
or U26810 (N_26810,N_24550,N_24560);
or U26811 (N_26811,N_22871,N_23422);
and U26812 (N_26812,N_23971,N_22698);
xor U26813 (N_26813,N_23173,N_24661);
or U26814 (N_26814,N_23467,N_24138);
and U26815 (N_26815,N_22802,N_24448);
and U26816 (N_26816,N_22635,N_23631);
and U26817 (N_26817,N_24394,N_23885);
nor U26818 (N_26818,N_23307,N_24165);
xor U26819 (N_26819,N_23369,N_22624);
nor U26820 (N_26820,N_24130,N_22779);
and U26821 (N_26821,N_24006,N_22920);
nor U26822 (N_26822,N_23831,N_24696);
and U26823 (N_26823,N_24610,N_24933);
and U26824 (N_26824,N_24460,N_24247);
nand U26825 (N_26825,N_24941,N_24106);
xnor U26826 (N_26826,N_24168,N_24241);
nand U26827 (N_26827,N_23601,N_23359);
nor U26828 (N_26828,N_24335,N_22732);
and U26829 (N_26829,N_22622,N_24465);
nand U26830 (N_26830,N_23840,N_22793);
and U26831 (N_26831,N_23235,N_24109);
and U26832 (N_26832,N_23521,N_23244);
nand U26833 (N_26833,N_23324,N_22671);
and U26834 (N_26834,N_23530,N_24093);
or U26835 (N_26835,N_23847,N_23024);
xnor U26836 (N_26836,N_23500,N_24304);
nand U26837 (N_26837,N_24575,N_24759);
or U26838 (N_26838,N_24333,N_23968);
nand U26839 (N_26839,N_22572,N_22669);
and U26840 (N_26840,N_22844,N_23452);
nor U26841 (N_26841,N_23565,N_24015);
and U26842 (N_26842,N_24173,N_23588);
xnor U26843 (N_26843,N_24284,N_23068);
or U26844 (N_26844,N_24447,N_22571);
nor U26845 (N_26845,N_24047,N_24887);
xor U26846 (N_26846,N_23005,N_23871);
or U26847 (N_26847,N_23709,N_24859);
nor U26848 (N_26848,N_22502,N_24638);
xnor U26849 (N_26849,N_22521,N_24366);
nand U26850 (N_26850,N_23930,N_24553);
and U26851 (N_26851,N_23245,N_23428);
nor U26852 (N_26852,N_24597,N_23537);
xnor U26853 (N_26853,N_24553,N_23415);
nand U26854 (N_26854,N_24193,N_22570);
or U26855 (N_26855,N_22622,N_24229);
xor U26856 (N_26856,N_24682,N_23914);
nand U26857 (N_26857,N_22650,N_22619);
or U26858 (N_26858,N_23980,N_23399);
xnor U26859 (N_26859,N_23884,N_24810);
nand U26860 (N_26860,N_23919,N_24818);
xnor U26861 (N_26861,N_23363,N_24946);
nor U26862 (N_26862,N_23233,N_23771);
or U26863 (N_26863,N_24069,N_24421);
nand U26864 (N_26864,N_23151,N_23328);
and U26865 (N_26865,N_22731,N_24212);
and U26866 (N_26866,N_24305,N_23683);
and U26867 (N_26867,N_22780,N_23570);
nor U26868 (N_26868,N_22733,N_23819);
nand U26869 (N_26869,N_22977,N_24141);
nand U26870 (N_26870,N_24362,N_23554);
nor U26871 (N_26871,N_23060,N_24178);
or U26872 (N_26872,N_24739,N_22981);
xnor U26873 (N_26873,N_22563,N_22684);
xor U26874 (N_26874,N_24578,N_23655);
or U26875 (N_26875,N_23602,N_23689);
and U26876 (N_26876,N_24163,N_24713);
xor U26877 (N_26877,N_22558,N_23843);
nand U26878 (N_26878,N_24490,N_24009);
nor U26879 (N_26879,N_24705,N_24691);
xnor U26880 (N_26880,N_22895,N_22950);
xor U26881 (N_26881,N_24505,N_24953);
or U26882 (N_26882,N_23834,N_24581);
xor U26883 (N_26883,N_22726,N_23042);
and U26884 (N_26884,N_22940,N_24830);
nand U26885 (N_26885,N_23369,N_23267);
xor U26886 (N_26886,N_24641,N_22764);
and U26887 (N_26887,N_22821,N_22528);
nand U26888 (N_26888,N_22792,N_23982);
and U26889 (N_26889,N_23884,N_24267);
nor U26890 (N_26890,N_22501,N_24934);
and U26891 (N_26891,N_23663,N_24735);
nand U26892 (N_26892,N_23721,N_22793);
and U26893 (N_26893,N_22645,N_23681);
nand U26894 (N_26894,N_24905,N_22903);
xnor U26895 (N_26895,N_24887,N_23135);
and U26896 (N_26896,N_22644,N_23794);
nand U26897 (N_26897,N_24642,N_23814);
or U26898 (N_26898,N_24042,N_24370);
nor U26899 (N_26899,N_24649,N_23679);
xnor U26900 (N_26900,N_24437,N_23787);
and U26901 (N_26901,N_24596,N_22792);
or U26902 (N_26902,N_22882,N_23599);
or U26903 (N_26903,N_23027,N_22629);
nor U26904 (N_26904,N_23304,N_24860);
nand U26905 (N_26905,N_22921,N_23190);
and U26906 (N_26906,N_24474,N_24744);
and U26907 (N_26907,N_22631,N_23029);
nand U26908 (N_26908,N_24962,N_24130);
or U26909 (N_26909,N_24229,N_24635);
and U26910 (N_26910,N_24022,N_22593);
or U26911 (N_26911,N_23139,N_23638);
nand U26912 (N_26912,N_22930,N_24329);
or U26913 (N_26913,N_23996,N_22915);
nor U26914 (N_26914,N_23521,N_22641);
nand U26915 (N_26915,N_22969,N_24134);
or U26916 (N_26916,N_23658,N_24112);
and U26917 (N_26917,N_24551,N_23599);
nor U26918 (N_26918,N_22542,N_22943);
nand U26919 (N_26919,N_24807,N_22927);
nor U26920 (N_26920,N_24453,N_24104);
xnor U26921 (N_26921,N_23849,N_23874);
nor U26922 (N_26922,N_24952,N_22754);
xor U26923 (N_26923,N_22697,N_23595);
or U26924 (N_26924,N_24966,N_23053);
nand U26925 (N_26925,N_24400,N_24449);
nand U26926 (N_26926,N_22627,N_24942);
nand U26927 (N_26927,N_22931,N_24633);
or U26928 (N_26928,N_23119,N_23273);
or U26929 (N_26929,N_24748,N_23160);
xor U26930 (N_26930,N_23822,N_23394);
or U26931 (N_26931,N_24790,N_24996);
and U26932 (N_26932,N_22625,N_23028);
nor U26933 (N_26933,N_23245,N_23722);
and U26934 (N_26934,N_23606,N_22910);
nand U26935 (N_26935,N_22603,N_23859);
nor U26936 (N_26936,N_22592,N_24648);
and U26937 (N_26937,N_24817,N_23228);
and U26938 (N_26938,N_22785,N_23819);
and U26939 (N_26939,N_22622,N_23219);
nor U26940 (N_26940,N_24219,N_23731);
or U26941 (N_26941,N_22637,N_22974);
nor U26942 (N_26942,N_24525,N_23517);
or U26943 (N_26943,N_24765,N_23627);
nand U26944 (N_26944,N_23775,N_23909);
or U26945 (N_26945,N_24709,N_22858);
and U26946 (N_26946,N_22863,N_24045);
or U26947 (N_26947,N_22717,N_24896);
and U26948 (N_26948,N_22565,N_23865);
and U26949 (N_26949,N_22634,N_22527);
and U26950 (N_26950,N_22814,N_24965);
and U26951 (N_26951,N_24994,N_24120);
nor U26952 (N_26952,N_22550,N_24536);
and U26953 (N_26953,N_24960,N_23181);
or U26954 (N_26954,N_24847,N_24154);
xnor U26955 (N_26955,N_24175,N_24537);
nand U26956 (N_26956,N_22797,N_22668);
or U26957 (N_26957,N_23200,N_24840);
nor U26958 (N_26958,N_22995,N_24592);
and U26959 (N_26959,N_24214,N_23228);
nand U26960 (N_26960,N_23979,N_22930);
nand U26961 (N_26961,N_23083,N_23980);
or U26962 (N_26962,N_23691,N_23823);
xnor U26963 (N_26963,N_22910,N_24648);
xnor U26964 (N_26964,N_22721,N_23790);
or U26965 (N_26965,N_22531,N_22813);
and U26966 (N_26966,N_24436,N_23244);
and U26967 (N_26967,N_24728,N_24283);
and U26968 (N_26968,N_23498,N_24375);
and U26969 (N_26969,N_24649,N_23279);
nor U26970 (N_26970,N_24618,N_24006);
or U26971 (N_26971,N_24366,N_24024);
or U26972 (N_26972,N_24336,N_24511);
nor U26973 (N_26973,N_23449,N_24199);
and U26974 (N_26974,N_24195,N_23218);
xnor U26975 (N_26975,N_22666,N_23921);
or U26976 (N_26976,N_23297,N_23076);
and U26977 (N_26977,N_24320,N_23025);
or U26978 (N_26978,N_23968,N_24723);
or U26979 (N_26979,N_23148,N_22906);
nand U26980 (N_26980,N_22924,N_24307);
or U26981 (N_26981,N_23164,N_22533);
xor U26982 (N_26982,N_22815,N_24408);
and U26983 (N_26983,N_24553,N_23191);
xor U26984 (N_26984,N_24348,N_24770);
nor U26985 (N_26985,N_23490,N_24443);
nand U26986 (N_26986,N_23727,N_23238);
xnor U26987 (N_26987,N_22597,N_24467);
nand U26988 (N_26988,N_24781,N_22766);
nand U26989 (N_26989,N_23772,N_23993);
xnor U26990 (N_26990,N_22622,N_24793);
and U26991 (N_26991,N_23879,N_24319);
nor U26992 (N_26992,N_24502,N_23894);
nor U26993 (N_26993,N_22785,N_23279);
xnor U26994 (N_26994,N_24887,N_22841);
xor U26995 (N_26995,N_23824,N_24474);
xnor U26996 (N_26996,N_24376,N_24016);
nand U26997 (N_26997,N_23193,N_24140);
and U26998 (N_26998,N_23605,N_24523);
or U26999 (N_26999,N_24162,N_23156);
and U27000 (N_27000,N_24298,N_22993);
nor U27001 (N_27001,N_23373,N_24095);
and U27002 (N_27002,N_24453,N_24847);
and U27003 (N_27003,N_24042,N_22533);
and U27004 (N_27004,N_23569,N_24562);
nand U27005 (N_27005,N_24029,N_24278);
or U27006 (N_27006,N_23059,N_22856);
nor U27007 (N_27007,N_22560,N_23162);
or U27008 (N_27008,N_24820,N_23137);
nand U27009 (N_27009,N_24717,N_23417);
xor U27010 (N_27010,N_22754,N_23269);
nor U27011 (N_27011,N_24602,N_24297);
nor U27012 (N_27012,N_23114,N_23913);
or U27013 (N_27013,N_24567,N_24702);
or U27014 (N_27014,N_23693,N_22565);
nor U27015 (N_27015,N_22694,N_24616);
and U27016 (N_27016,N_24291,N_24930);
nand U27017 (N_27017,N_24012,N_24267);
and U27018 (N_27018,N_24862,N_22764);
nor U27019 (N_27019,N_23407,N_23950);
and U27020 (N_27020,N_24088,N_22749);
and U27021 (N_27021,N_22866,N_24013);
and U27022 (N_27022,N_24785,N_24513);
or U27023 (N_27023,N_24681,N_23509);
nand U27024 (N_27024,N_23880,N_23533);
nand U27025 (N_27025,N_22829,N_23800);
nand U27026 (N_27026,N_23827,N_23900);
nand U27027 (N_27027,N_23625,N_23778);
nand U27028 (N_27028,N_24556,N_23077);
or U27029 (N_27029,N_22574,N_24294);
and U27030 (N_27030,N_22557,N_24706);
and U27031 (N_27031,N_24877,N_24339);
nor U27032 (N_27032,N_22689,N_22931);
xnor U27033 (N_27033,N_22725,N_24379);
nor U27034 (N_27034,N_24578,N_22583);
or U27035 (N_27035,N_23676,N_23792);
or U27036 (N_27036,N_23445,N_23707);
and U27037 (N_27037,N_23079,N_24477);
xor U27038 (N_27038,N_22510,N_23356);
xor U27039 (N_27039,N_23423,N_23966);
xnor U27040 (N_27040,N_23105,N_23150);
nor U27041 (N_27041,N_24771,N_22606);
nor U27042 (N_27042,N_24601,N_23331);
nor U27043 (N_27043,N_24680,N_24460);
or U27044 (N_27044,N_24557,N_24797);
and U27045 (N_27045,N_22798,N_24145);
nor U27046 (N_27046,N_23630,N_23559);
xor U27047 (N_27047,N_23727,N_24688);
nand U27048 (N_27048,N_22989,N_24576);
nor U27049 (N_27049,N_24423,N_24596);
xor U27050 (N_27050,N_24897,N_24493);
nor U27051 (N_27051,N_23575,N_22752);
nand U27052 (N_27052,N_24611,N_23276);
or U27053 (N_27053,N_23664,N_22838);
xnor U27054 (N_27054,N_24354,N_24768);
or U27055 (N_27055,N_23115,N_23466);
nand U27056 (N_27056,N_23882,N_23613);
nand U27057 (N_27057,N_23109,N_23529);
or U27058 (N_27058,N_24224,N_24725);
and U27059 (N_27059,N_23257,N_24870);
nor U27060 (N_27060,N_23106,N_23653);
or U27061 (N_27061,N_23631,N_22541);
xor U27062 (N_27062,N_23669,N_24821);
or U27063 (N_27063,N_24206,N_23737);
nor U27064 (N_27064,N_22838,N_24728);
nor U27065 (N_27065,N_22658,N_23715);
nand U27066 (N_27066,N_22566,N_23685);
or U27067 (N_27067,N_23609,N_23332);
nand U27068 (N_27068,N_24739,N_23660);
and U27069 (N_27069,N_23166,N_22711);
xor U27070 (N_27070,N_23535,N_23429);
nor U27071 (N_27071,N_23397,N_22620);
nand U27072 (N_27072,N_24748,N_22924);
nor U27073 (N_27073,N_22771,N_24226);
xor U27074 (N_27074,N_23301,N_24777);
nor U27075 (N_27075,N_23866,N_23913);
xor U27076 (N_27076,N_23537,N_24457);
and U27077 (N_27077,N_24701,N_24155);
xor U27078 (N_27078,N_24469,N_23289);
and U27079 (N_27079,N_23964,N_24094);
nand U27080 (N_27080,N_23212,N_22529);
nor U27081 (N_27081,N_24225,N_23203);
nor U27082 (N_27082,N_23824,N_24469);
xor U27083 (N_27083,N_24265,N_24764);
and U27084 (N_27084,N_24258,N_22662);
xor U27085 (N_27085,N_24670,N_23113);
and U27086 (N_27086,N_22726,N_24432);
or U27087 (N_27087,N_24037,N_22991);
and U27088 (N_27088,N_23001,N_23770);
and U27089 (N_27089,N_24061,N_23917);
nand U27090 (N_27090,N_24747,N_24823);
and U27091 (N_27091,N_23624,N_23069);
xnor U27092 (N_27092,N_22731,N_23436);
nor U27093 (N_27093,N_23320,N_24023);
and U27094 (N_27094,N_23863,N_24001);
and U27095 (N_27095,N_24564,N_22754);
xnor U27096 (N_27096,N_24435,N_24554);
or U27097 (N_27097,N_23321,N_23594);
or U27098 (N_27098,N_22894,N_23046);
nor U27099 (N_27099,N_24834,N_23414);
nor U27100 (N_27100,N_23132,N_23561);
or U27101 (N_27101,N_23601,N_24168);
nand U27102 (N_27102,N_23374,N_24288);
or U27103 (N_27103,N_22880,N_24581);
nor U27104 (N_27104,N_24380,N_24734);
nand U27105 (N_27105,N_23006,N_23503);
nor U27106 (N_27106,N_23188,N_24031);
and U27107 (N_27107,N_23962,N_24975);
nand U27108 (N_27108,N_22651,N_24609);
xor U27109 (N_27109,N_24520,N_23537);
xnor U27110 (N_27110,N_22576,N_24781);
nor U27111 (N_27111,N_24565,N_24824);
xnor U27112 (N_27112,N_24628,N_24732);
nand U27113 (N_27113,N_24659,N_22635);
nand U27114 (N_27114,N_24672,N_22776);
nand U27115 (N_27115,N_22603,N_22896);
and U27116 (N_27116,N_24030,N_24083);
nand U27117 (N_27117,N_22547,N_23696);
and U27118 (N_27118,N_22613,N_24557);
nand U27119 (N_27119,N_23320,N_24070);
and U27120 (N_27120,N_22997,N_22561);
xnor U27121 (N_27121,N_22793,N_24622);
or U27122 (N_27122,N_23341,N_24454);
nor U27123 (N_27123,N_24787,N_23790);
or U27124 (N_27124,N_22945,N_24211);
nor U27125 (N_27125,N_24319,N_22831);
nor U27126 (N_27126,N_23656,N_23209);
nor U27127 (N_27127,N_24615,N_22777);
or U27128 (N_27128,N_22841,N_22697);
nand U27129 (N_27129,N_23438,N_23117);
or U27130 (N_27130,N_24025,N_24137);
or U27131 (N_27131,N_22928,N_23821);
nor U27132 (N_27132,N_24993,N_24921);
and U27133 (N_27133,N_24354,N_24486);
xnor U27134 (N_27134,N_23456,N_22884);
nor U27135 (N_27135,N_22844,N_24821);
xnor U27136 (N_27136,N_24545,N_23485);
and U27137 (N_27137,N_22997,N_23383);
and U27138 (N_27138,N_24245,N_23503);
nor U27139 (N_27139,N_23007,N_24811);
xor U27140 (N_27140,N_24253,N_23742);
and U27141 (N_27141,N_23097,N_24642);
nor U27142 (N_27142,N_22597,N_24569);
nor U27143 (N_27143,N_24804,N_23758);
xor U27144 (N_27144,N_22802,N_24978);
and U27145 (N_27145,N_24181,N_24841);
xnor U27146 (N_27146,N_23204,N_22586);
nand U27147 (N_27147,N_24955,N_23861);
or U27148 (N_27148,N_24344,N_23143);
or U27149 (N_27149,N_23808,N_24078);
or U27150 (N_27150,N_23162,N_24802);
xnor U27151 (N_27151,N_24310,N_24084);
or U27152 (N_27152,N_22937,N_22562);
nand U27153 (N_27153,N_23861,N_24281);
or U27154 (N_27154,N_22929,N_24252);
xor U27155 (N_27155,N_23212,N_23127);
xor U27156 (N_27156,N_23908,N_24621);
xor U27157 (N_27157,N_24860,N_23435);
and U27158 (N_27158,N_23434,N_24091);
and U27159 (N_27159,N_23665,N_23245);
and U27160 (N_27160,N_23420,N_22818);
or U27161 (N_27161,N_23518,N_24327);
nor U27162 (N_27162,N_23659,N_24581);
xor U27163 (N_27163,N_22613,N_24554);
or U27164 (N_27164,N_22681,N_22507);
and U27165 (N_27165,N_22786,N_24251);
nor U27166 (N_27166,N_23305,N_23788);
nor U27167 (N_27167,N_23655,N_23594);
xnor U27168 (N_27168,N_22574,N_24450);
xor U27169 (N_27169,N_24525,N_24635);
or U27170 (N_27170,N_23737,N_22558);
nor U27171 (N_27171,N_23841,N_24350);
nor U27172 (N_27172,N_24328,N_23546);
xor U27173 (N_27173,N_22984,N_24066);
or U27174 (N_27174,N_24910,N_23600);
and U27175 (N_27175,N_24084,N_24180);
nor U27176 (N_27176,N_23918,N_24221);
xnor U27177 (N_27177,N_24831,N_23629);
and U27178 (N_27178,N_22622,N_24168);
nor U27179 (N_27179,N_23713,N_23051);
nand U27180 (N_27180,N_22913,N_24362);
xnor U27181 (N_27181,N_24574,N_24046);
nand U27182 (N_27182,N_23437,N_24499);
or U27183 (N_27183,N_24241,N_22742);
xnor U27184 (N_27184,N_24858,N_23886);
or U27185 (N_27185,N_24664,N_24147);
and U27186 (N_27186,N_22677,N_24604);
nand U27187 (N_27187,N_24235,N_22800);
nor U27188 (N_27188,N_23121,N_22859);
nor U27189 (N_27189,N_24803,N_24547);
or U27190 (N_27190,N_23648,N_23119);
nand U27191 (N_27191,N_23861,N_24673);
xnor U27192 (N_27192,N_24023,N_24912);
nand U27193 (N_27193,N_24268,N_23476);
nor U27194 (N_27194,N_24464,N_22924);
xnor U27195 (N_27195,N_22721,N_22735);
nor U27196 (N_27196,N_23621,N_23262);
nor U27197 (N_27197,N_24482,N_22667);
or U27198 (N_27198,N_22526,N_23219);
nand U27199 (N_27199,N_24810,N_24042);
xor U27200 (N_27200,N_22943,N_22868);
or U27201 (N_27201,N_23940,N_22964);
nor U27202 (N_27202,N_24424,N_22522);
nand U27203 (N_27203,N_23262,N_24313);
nand U27204 (N_27204,N_24667,N_24041);
nor U27205 (N_27205,N_23555,N_22633);
nor U27206 (N_27206,N_22974,N_23316);
xor U27207 (N_27207,N_23678,N_22704);
or U27208 (N_27208,N_24064,N_23798);
nand U27209 (N_27209,N_23459,N_22554);
nand U27210 (N_27210,N_23450,N_22830);
or U27211 (N_27211,N_23170,N_24803);
nand U27212 (N_27212,N_24576,N_23508);
nor U27213 (N_27213,N_24828,N_24210);
nor U27214 (N_27214,N_22897,N_22740);
and U27215 (N_27215,N_23674,N_23601);
and U27216 (N_27216,N_24991,N_24949);
or U27217 (N_27217,N_24058,N_24743);
nor U27218 (N_27218,N_22832,N_24124);
nor U27219 (N_27219,N_24989,N_22539);
xnor U27220 (N_27220,N_24629,N_22561);
and U27221 (N_27221,N_24261,N_23407);
nor U27222 (N_27222,N_24931,N_22866);
xor U27223 (N_27223,N_23717,N_24130);
nor U27224 (N_27224,N_22858,N_23402);
or U27225 (N_27225,N_24322,N_24760);
or U27226 (N_27226,N_22743,N_23214);
and U27227 (N_27227,N_24989,N_23847);
or U27228 (N_27228,N_24079,N_24476);
nor U27229 (N_27229,N_24561,N_24352);
nand U27230 (N_27230,N_24671,N_24778);
nand U27231 (N_27231,N_22933,N_23827);
or U27232 (N_27232,N_23437,N_24276);
and U27233 (N_27233,N_24518,N_24984);
nand U27234 (N_27234,N_22874,N_24562);
nand U27235 (N_27235,N_23252,N_22581);
or U27236 (N_27236,N_23599,N_23413);
xnor U27237 (N_27237,N_24974,N_22697);
nor U27238 (N_27238,N_22811,N_23830);
xnor U27239 (N_27239,N_22969,N_24976);
and U27240 (N_27240,N_22812,N_24996);
xnor U27241 (N_27241,N_24903,N_24553);
nor U27242 (N_27242,N_23030,N_23887);
and U27243 (N_27243,N_22542,N_22525);
nor U27244 (N_27244,N_22957,N_24200);
or U27245 (N_27245,N_23226,N_23430);
or U27246 (N_27246,N_23590,N_24866);
nand U27247 (N_27247,N_22573,N_24595);
xor U27248 (N_27248,N_22956,N_24112);
xor U27249 (N_27249,N_23891,N_24394);
nor U27250 (N_27250,N_24553,N_24309);
nand U27251 (N_27251,N_23418,N_24980);
or U27252 (N_27252,N_22972,N_24013);
or U27253 (N_27253,N_23631,N_24791);
nor U27254 (N_27254,N_23766,N_22964);
nand U27255 (N_27255,N_22587,N_24730);
nand U27256 (N_27256,N_23157,N_22734);
nor U27257 (N_27257,N_23330,N_24819);
and U27258 (N_27258,N_22928,N_23699);
nor U27259 (N_27259,N_23124,N_23925);
xor U27260 (N_27260,N_22621,N_24895);
xor U27261 (N_27261,N_22797,N_24692);
nand U27262 (N_27262,N_23742,N_23133);
or U27263 (N_27263,N_23350,N_23797);
nand U27264 (N_27264,N_24136,N_24471);
nand U27265 (N_27265,N_23811,N_23005);
nor U27266 (N_27266,N_24889,N_23883);
nand U27267 (N_27267,N_23330,N_24298);
nor U27268 (N_27268,N_22996,N_23247);
xor U27269 (N_27269,N_22571,N_24715);
and U27270 (N_27270,N_23754,N_23910);
xor U27271 (N_27271,N_24668,N_24971);
and U27272 (N_27272,N_23156,N_23350);
or U27273 (N_27273,N_23692,N_23073);
xor U27274 (N_27274,N_24355,N_23063);
xnor U27275 (N_27275,N_24362,N_24972);
nand U27276 (N_27276,N_23255,N_24104);
and U27277 (N_27277,N_24957,N_22663);
xnor U27278 (N_27278,N_23677,N_23994);
and U27279 (N_27279,N_24252,N_22950);
or U27280 (N_27280,N_22753,N_22500);
and U27281 (N_27281,N_23650,N_24830);
xor U27282 (N_27282,N_22544,N_24592);
xor U27283 (N_27283,N_23564,N_23556);
xor U27284 (N_27284,N_23141,N_24208);
nand U27285 (N_27285,N_23574,N_24804);
xor U27286 (N_27286,N_23269,N_22588);
nor U27287 (N_27287,N_23130,N_24768);
nor U27288 (N_27288,N_23923,N_22593);
nand U27289 (N_27289,N_24319,N_24121);
nor U27290 (N_27290,N_23075,N_22777);
and U27291 (N_27291,N_23446,N_23624);
or U27292 (N_27292,N_24464,N_22581);
or U27293 (N_27293,N_23748,N_24653);
nand U27294 (N_27294,N_23354,N_23636);
nand U27295 (N_27295,N_23833,N_24721);
nor U27296 (N_27296,N_24271,N_24673);
or U27297 (N_27297,N_22698,N_24314);
xor U27298 (N_27298,N_23493,N_23021);
xor U27299 (N_27299,N_23146,N_23653);
xor U27300 (N_27300,N_23416,N_22748);
nor U27301 (N_27301,N_23141,N_23341);
nand U27302 (N_27302,N_22841,N_23091);
and U27303 (N_27303,N_22849,N_23608);
or U27304 (N_27304,N_23913,N_24757);
and U27305 (N_27305,N_22868,N_23864);
and U27306 (N_27306,N_23968,N_22933);
and U27307 (N_27307,N_23403,N_22642);
xor U27308 (N_27308,N_22752,N_23683);
nor U27309 (N_27309,N_24727,N_22812);
nand U27310 (N_27310,N_24741,N_22621);
and U27311 (N_27311,N_22652,N_23855);
or U27312 (N_27312,N_23435,N_23130);
or U27313 (N_27313,N_23992,N_24370);
or U27314 (N_27314,N_22545,N_24692);
nand U27315 (N_27315,N_22598,N_24410);
nor U27316 (N_27316,N_24974,N_23319);
nand U27317 (N_27317,N_23476,N_24906);
xor U27318 (N_27318,N_24865,N_22952);
nor U27319 (N_27319,N_23602,N_23439);
nor U27320 (N_27320,N_24430,N_23511);
nand U27321 (N_27321,N_22806,N_23552);
or U27322 (N_27322,N_23932,N_23718);
and U27323 (N_27323,N_23621,N_23129);
or U27324 (N_27324,N_23889,N_24748);
and U27325 (N_27325,N_24594,N_23494);
nand U27326 (N_27326,N_23466,N_23121);
or U27327 (N_27327,N_23797,N_24899);
nand U27328 (N_27328,N_22839,N_22806);
and U27329 (N_27329,N_23876,N_24379);
xor U27330 (N_27330,N_23254,N_24232);
xnor U27331 (N_27331,N_23826,N_23597);
or U27332 (N_27332,N_24241,N_23962);
nor U27333 (N_27333,N_24499,N_24061);
and U27334 (N_27334,N_23211,N_23015);
nand U27335 (N_27335,N_22562,N_24517);
or U27336 (N_27336,N_24900,N_23404);
or U27337 (N_27337,N_24416,N_24464);
nor U27338 (N_27338,N_22616,N_24535);
nor U27339 (N_27339,N_24188,N_23190);
nor U27340 (N_27340,N_23398,N_23998);
xor U27341 (N_27341,N_24798,N_24133);
and U27342 (N_27342,N_23569,N_23736);
or U27343 (N_27343,N_24593,N_22764);
nor U27344 (N_27344,N_24469,N_23567);
xor U27345 (N_27345,N_23705,N_22669);
nand U27346 (N_27346,N_22861,N_22637);
nand U27347 (N_27347,N_24655,N_24049);
nor U27348 (N_27348,N_23012,N_22782);
and U27349 (N_27349,N_24518,N_23898);
xor U27350 (N_27350,N_24733,N_23317);
nand U27351 (N_27351,N_23189,N_23048);
xnor U27352 (N_27352,N_22911,N_22584);
nor U27353 (N_27353,N_24029,N_22976);
xnor U27354 (N_27354,N_23599,N_24187);
and U27355 (N_27355,N_22566,N_22657);
nand U27356 (N_27356,N_24576,N_23535);
xor U27357 (N_27357,N_24264,N_22930);
xnor U27358 (N_27358,N_24549,N_22788);
nor U27359 (N_27359,N_22883,N_24574);
nor U27360 (N_27360,N_24736,N_24407);
or U27361 (N_27361,N_23390,N_23214);
and U27362 (N_27362,N_23213,N_24055);
nor U27363 (N_27363,N_24299,N_24073);
nand U27364 (N_27364,N_24726,N_23709);
and U27365 (N_27365,N_24425,N_24680);
nor U27366 (N_27366,N_23684,N_23873);
nand U27367 (N_27367,N_23284,N_24951);
xor U27368 (N_27368,N_23444,N_24340);
nor U27369 (N_27369,N_22910,N_24027);
or U27370 (N_27370,N_24196,N_24965);
nor U27371 (N_27371,N_22716,N_23240);
xnor U27372 (N_27372,N_24804,N_23495);
nand U27373 (N_27373,N_23399,N_24541);
nand U27374 (N_27374,N_24891,N_24006);
nand U27375 (N_27375,N_23875,N_22987);
nor U27376 (N_27376,N_24306,N_23922);
nor U27377 (N_27377,N_24248,N_22917);
or U27378 (N_27378,N_23601,N_24331);
nand U27379 (N_27379,N_22570,N_23284);
or U27380 (N_27380,N_24519,N_24035);
nor U27381 (N_27381,N_24311,N_23209);
nand U27382 (N_27382,N_24815,N_22627);
and U27383 (N_27383,N_24938,N_24357);
and U27384 (N_27384,N_23714,N_24951);
and U27385 (N_27385,N_24934,N_23899);
nand U27386 (N_27386,N_24601,N_23301);
and U27387 (N_27387,N_23006,N_24080);
nand U27388 (N_27388,N_24358,N_22758);
nand U27389 (N_27389,N_24039,N_23094);
nand U27390 (N_27390,N_24845,N_22520);
nor U27391 (N_27391,N_23812,N_24157);
and U27392 (N_27392,N_23367,N_24252);
nand U27393 (N_27393,N_24800,N_22710);
nand U27394 (N_27394,N_22775,N_23782);
nor U27395 (N_27395,N_24334,N_23889);
nor U27396 (N_27396,N_23707,N_22529);
and U27397 (N_27397,N_24198,N_23677);
xor U27398 (N_27398,N_24410,N_24815);
or U27399 (N_27399,N_23892,N_24388);
xnor U27400 (N_27400,N_24900,N_23119);
xor U27401 (N_27401,N_23966,N_23517);
nand U27402 (N_27402,N_23790,N_23431);
or U27403 (N_27403,N_22583,N_23289);
or U27404 (N_27404,N_24403,N_24962);
nand U27405 (N_27405,N_23154,N_23872);
xor U27406 (N_27406,N_24562,N_24187);
and U27407 (N_27407,N_24940,N_22639);
and U27408 (N_27408,N_23229,N_22843);
or U27409 (N_27409,N_24734,N_23166);
and U27410 (N_27410,N_22784,N_24916);
nor U27411 (N_27411,N_24552,N_24248);
and U27412 (N_27412,N_22861,N_24942);
and U27413 (N_27413,N_24557,N_22685);
and U27414 (N_27414,N_23004,N_24760);
or U27415 (N_27415,N_24684,N_23671);
and U27416 (N_27416,N_24148,N_24398);
nand U27417 (N_27417,N_24056,N_22789);
nand U27418 (N_27418,N_23690,N_24172);
xor U27419 (N_27419,N_24506,N_23207);
nor U27420 (N_27420,N_22573,N_23925);
xor U27421 (N_27421,N_24428,N_24403);
and U27422 (N_27422,N_23718,N_23581);
nand U27423 (N_27423,N_23574,N_24894);
xor U27424 (N_27424,N_23664,N_24160);
xor U27425 (N_27425,N_24564,N_24506);
nand U27426 (N_27426,N_24641,N_23915);
xor U27427 (N_27427,N_24054,N_24848);
and U27428 (N_27428,N_23180,N_22757);
or U27429 (N_27429,N_22824,N_24034);
nor U27430 (N_27430,N_24032,N_24901);
and U27431 (N_27431,N_23065,N_24063);
and U27432 (N_27432,N_24436,N_24000);
xor U27433 (N_27433,N_23091,N_22834);
nand U27434 (N_27434,N_23345,N_23941);
or U27435 (N_27435,N_23229,N_22822);
or U27436 (N_27436,N_23749,N_22721);
and U27437 (N_27437,N_23257,N_24721);
xor U27438 (N_27438,N_24404,N_22546);
and U27439 (N_27439,N_22989,N_22773);
or U27440 (N_27440,N_24484,N_23624);
xor U27441 (N_27441,N_24555,N_23063);
and U27442 (N_27442,N_22535,N_24418);
xor U27443 (N_27443,N_23607,N_23391);
nor U27444 (N_27444,N_23493,N_24036);
nand U27445 (N_27445,N_22756,N_23207);
xor U27446 (N_27446,N_24218,N_23831);
nor U27447 (N_27447,N_24216,N_22735);
nor U27448 (N_27448,N_24840,N_23712);
or U27449 (N_27449,N_23386,N_24282);
and U27450 (N_27450,N_24447,N_22501);
nand U27451 (N_27451,N_23417,N_24474);
nand U27452 (N_27452,N_22695,N_23572);
xor U27453 (N_27453,N_22825,N_23573);
nor U27454 (N_27454,N_22942,N_24410);
nand U27455 (N_27455,N_24570,N_24673);
and U27456 (N_27456,N_23570,N_23213);
nand U27457 (N_27457,N_24889,N_22703);
and U27458 (N_27458,N_24092,N_22896);
nor U27459 (N_27459,N_23196,N_24924);
nor U27460 (N_27460,N_22726,N_23525);
nor U27461 (N_27461,N_24331,N_24590);
or U27462 (N_27462,N_22638,N_24701);
nand U27463 (N_27463,N_24216,N_23996);
xor U27464 (N_27464,N_24370,N_23326);
and U27465 (N_27465,N_24646,N_24704);
and U27466 (N_27466,N_23540,N_24220);
xor U27467 (N_27467,N_22695,N_24428);
nand U27468 (N_27468,N_23681,N_22855);
xnor U27469 (N_27469,N_24492,N_24489);
or U27470 (N_27470,N_24825,N_23687);
xnor U27471 (N_27471,N_23764,N_24523);
xnor U27472 (N_27472,N_24045,N_23147);
or U27473 (N_27473,N_24282,N_24252);
and U27474 (N_27474,N_24467,N_23828);
xor U27475 (N_27475,N_23722,N_23184);
nor U27476 (N_27476,N_22620,N_22775);
or U27477 (N_27477,N_23529,N_24797);
xnor U27478 (N_27478,N_23104,N_24957);
nand U27479 (N_27479,N_24770,N_23519);
xor U27480 (N_27480,N_24123,N_24069);
nor U27481 (N_27481,N_23700,N_22565);
or U27482 (N_27482,N_23450,N_23861);
and U27483 (N_27483,N_23329,N_23599);
and U27484 (N_27484,N_23594,N_23806);
xor U27485 (N_27485,N_22512,N_23179);
and U27486 (N_27486,N_23774,N_22872);
nor U27487 (N_27487,N_22556,N_23899);
nand U27488 (N_27488,N_22913,N_22595);
nand U27489 (N_27489,N_24356,N_23136);
nor U27490 (N_27490,N_24105,N_22927);
and U27491 (N_27491,N_23353,N_23197);
or U27492 (N_27492,N_22636,N_22609);
and U27493 (N_27493,N_24844,N_23235);
xor U27494 (N_27494,N_22809,N_24787);
xor U27495 (N_27495,N_24086,N_24348);
xnor U27496 (N_27496,N_23558,N_23212);
nor U27497 (N_27497,N_24752,N_23234);
or U27498 (N_27498,N_22948,N_23634);
or U27499 (N_27499,N_24076,N_22823);
or U27500 (N_27500,N_26929,N_25667);
nor U27501 (N_27501,N_26319,N_26143);
and U27502 (N_27502,N_27353,N_27017);
xnor U27503 (N_27503,N_25360,N_25485);
nand U27504 (N_27504,N_26775,N_25015);
xnor U27505 (N_27505,N_25666,N_27496);
nor U27506 (N_27506,N_27143,N_26126);
nor U27507 (N_27507,N_25287,N_27080);
nor U27508 (N_27508,N_26555,N_26470);
xor U27509 (N_27509,N_26202,N_25433);
xor U27510 (N_27510,N_26419,N_26615);
or U27511 (N_27511,N_25642,N_26974);
xor U27512 (N_27512,N_26950,N_26004);
xnor U27513 (N_27513,N_25641,N_25332);
nor U27514 (N_27514,N_27213,N_27413);
nor U27515 (N_27515,N_26531,N_25868);
and U27516 (N_27516,N_26030,N_25558);
and U27517 (N_27517,N_26608,N_26289);
nor U27518 (N_27518,N_26204,N_27276);
nor U27519 (N_27519,N_25810,N_25971);
nand U27520 (N_27520,N_26494,N_25095);
xor U27521 (N_27521,N_27472,N_26768);
and U27522 (N_27522,N_25804,N_27437);
and U27523 (N_27523,N_25704,N_26607);
nand U27524 (N_27524,N_25163,N_25061);
nand U27525 (N_27525,N_27156,N_25482);
nor U27526 (N_27526,N_26542,N_26315);
xor U27527 (N_27527,N_26762,N_26725);
or U27528 (N_27528,N_26627,N_26798);
nand U27529 (N_27529,N_27023,N_27222);
xor U27530 (N_27530,N_25238,N_26569);
nor U27531 (N_27531,N_26948,N_26696);
and U27532 (N_27532,N_25937,N_26525);
or U27533 (N_27533,N_25324,N_25016);
xnor U27534 (N_27534,N_27089,N_26394);
or U27535 (N_27535,N_25984,N_25613);
and U27536 (N_27536,N_27033,N_25721);
nor U27537 (N_27537,N_26671,N_26300);
or U27538 (N_27538,N_26943,N_25784);
or U27539 (N_27539,N_26084,N_26576);
nand U27540 (N_27540,N_27122,N_26796);
or U27541 (N_27541,N_26399,N_27274);
xor U27542 (N_27542,N_27331,N_27417);
and U27543 (N_27543,N_27452,N_27208);
nor U27544 (N_27544,N_27497,N_27139);
nand U27545 (N_27545,N_26593,N_26583);
xnor U27546 (N_27546,N_26164,N_26041);
or U27547 (N_27547,N_26913,N_25671);
and U27548 (N_27548,N_25409,N_25137);
or U27549 (N_27549,N_25614,N_26409);
and U27550 (N_27550,N_27463,N_25024);
or U27551 (N_27551,N_26447,N_25323);
nand U27552 (N_27552,N_25110,N_25996);
nor U27553 (N_27553,N_25056,N_27412);
or U27554 (N_27554,N_25689,N_25473);
or U27555 (N_27555,N_26735,N_26769);
nor U27556 (N_27556,N_25959,N_25242);
xnor U27557 (N_27557,N_26076,N_27319);
or U27558 (N_27558,N_25940,N_26311);
nand U27559 (N_27559,N_25303,N_26752);
nand U27560 (N_27560,N_27293,N_26770);
or U27561 (N_27561,N_26960,N_26630);
and U27562 (N_27562,N_25275,N_27249);
nand U27563 (N_27563,N_25833,N_26586);
or U27564 (N_27564,N_25091,N_25021);
nor U27565 (N_27565,N_25060,N_26666);
nor U27566 (N_27566,N_25847,N_25801);
or U27567 (N_27567,N_26867,N_25157);
or U27568 (N_27568,N_26171,N_27197);
xnor U27569 (N_27569,N_27205,N_27086);
xnor U27570 (N_27570,N_26170,N_26424);
or U27571 (N_27571,N_25223,N_27339);
xnor U27572 (N_27572,N_25445,N_26129);
nand U27573 (N_27573,N_25310,N_25298);
and U27574 (N_27574,N_25697,N_27016);
xor U27575 (N_27575,N_25053,N_26290);
nand U27576 (N_27576,N_25322,N_25987);
and U27577 (N_27577,N_26242,N_26585);
and U27578 (N_27578,N_26642,N_26907);
xnor U27579 (N_27579,N_27409,N_26556);
nand U27580 (N_27580,N_26108,N_27231);
and U27581 (N_27581,N_25909,N_25679);
nor U27582 (N_27582,N_26089,N_25559);
nand U27583 (N_27583,N_25738,N_25006);
and U27584 (N_27584,N_25557,N_26596);
nand U27585 (N_27585,N_25610,N_26883);
nand U27586 (N_27586,N_26254,N_25737);
nand U27587 (N_27587,N_27400,N_26916);
xor U27588 (N_27588,N_27165,N_25032);
xnor U27589 (N_27589,N_26207,N_26905);
xnor U27590 (N_27590,N_25716,N_26141);
nand U27591 (N_27591,N_26110,N_25342);
nand U27592 (N_27592,N_26001,N_25663);
xor U27593 (N_27593,N_25866,N_25403);
nand U27594 (N_27594,N_27467,N_25706);
or U27595 (N_27595,N_25200,N_27011);
xor U27596 (N_27596,N_25428,N_26610);
nor U27597 (N_27597,N_26540,N_25715);
xor U27598 (N_27598,N_25526,N_27354);
xnor U27599 (N_27599,N_26908,N_26454);
xor U27600 (N_27600,N_26625,N_25218);
nor U27601 (N_27601,N_26155,N_27352);
nor U27602 (N_27602,N_26348,N_25354);
xor U27603 (N_27603,N_26329,N_27022);
nand U27604 (N_27604,N_27286,N_25941);
xor U27605 (N_27605,N_25796,N_25086);
and U27606 (N_27606,N_25780,N_27041);
or U27607 (N_27607,N_26065,N_25012);
xor U27608 (N_27608,N_26807,N_25608);
xnor U27609 (N_27609,N_25915,N_25731);
nor U27610 (N_27610,N_25636,N_25257);
xor U27611 (N_27611,N_25654,N_26467);
xor U27612 (N_27612,N_25890,N_25264);
xnor U27613 (N_27613,N_26417,N_26362);
and U27614 (N_27614,N_25945,N_26732);
and U27615 (N_27615,N_26079,N_26487);
xnor U27616 (N_27616,N_25455,N_25373);
nand U27617 (N_27617,N_27120,N_25683);
nand U27618 (N_27618,N_26680,N_25074);
xnor U27619 (N_27619,N_25818,N_25949);
and U27620 (N_27620,N_25284,N_25420);
nand U27621 (N_27621,N_27104,N_26841);
nand U27622 (N_27622,N_26102,N_26476);
nand U27623 (N_27623,N_26081,N_25822);
nor U27624 (N_27624,N_25270,N_25861);
xor U27625 (N_27625,N_25897,N_25094);
or U27626 (N_27626,N_27367,N_26457);
xnor U27627 (N_27627,N_25970,N_25411);
xnor U27628 (N_27628,N_26521,N_25117);
nor U27629 (N_27629,N_27432,N_26982);
xor U27630 (N_27630,N_25229,N_27494);
and U27631 (N_27631,N_26431,N_25050);
and U27632 (N_27632,N_25406,N_27220);
xnor U27633 (N_27633,N_25700,N_27349);
xor U27634 (N_27634,N_26972,N_26008);
nor U27635 (N_27635,N_26167,N_25874);
nand U27636 (N_27636,N_25438,N_26993);
nor U27637 (N_27637,N_26379,N_25000);
and U27638 (N_27638,N_25691,N_26364);
xor U27639 (N_27639,N_26223,N_26378);
nand U27640 (N_27640,N_25025,N_25856);
and U27641 (N_27641,N_25175,N_26448);
nand U27642 (N_27642,N_26293,N_26322);
and U27643 (N_27643,N_25985,N_25151);
nor U27644 (N_27644,N_25809,N_26876);
xor U27645 (N_27645,N_25076,N_27038);
and U27646 (N_27646,N_25577,N_26658);
nor U27647 (N_27647,N_26480,N_26381);
nor U27648 (N_27648,N_25924,N_26574);
xor U27649 (N_27649,N_26387,N_26548);
and U27650 (N_27650,N_26321,N_26034);
nand U27651 (N_27651,N_26063,N_25521);
or U27652 (N_27652,N_27479,N_27262);
nor U27653 (N_27653,N_26243,N_27121);
nor U27654 (N_27654,N_26301,N_25158);
and U27655 (N_27655,N_26549,N_26229);
and U27656 (N_27656,N_26154,N_26923);
xor U27657 (N_27657,N_27183,N_26022);
or U27658 (N_27658,N_27492,N_26208);
nor U27659 (N_27659,N_26451,N_27272);
and U27660 (N_27660,N_25197,N_25246);
and U27661 (N_27661,N_26991,N_25400);
or U27662 (N_27662,N_26554,N_26622);
nand U27663 (N_27663,N_25168,N_25994);
and U27664 (N_27664,N_26591,N_25720);
xor U27665 (N_27665,N_27337,N_26595);
and U27666 (N_27666,N_25954,N_25556);
and U27667 (N_27667,N_25415,N_25840);
or U27668 (N_27668,N_26640,N_25293);
nand U27669 (N_27669,N_25509,N_27090);
or U27670 (N_27670,N_27054,N_25172);
xor U27671 (N_27671,N_25686,N_25670);
nand U27672 (N_27672,N_26432,N_25724);
or U27673 (N_27673,N_26949,N_26811);
and U27674 (N_27674,N_25525,N_27252);
nor U27675 (N_27675,N_25385,N_25593);
nand U27676 (N_27676,N_25358,N_27067);
xor U27677 (N_27677,N_25041,N_25146);
or U27678 (N_27678,N_25534,N_25602);
and U27679 (N_27679,N_26897,N_25936);
nand U27680 (N_27680,N_27307,N_26600);
nand U27681 (N_27681,N_26862,N_25267);
and U27682 (N_27682,N_25318,N_25101);
nand U27683 (N_27683,N_26205,N_27049);
xnor U27684 (N_27684,N_26994,N_25368);
nor U27685 (N_27685,N_25426,N_26511);
xor U27686 (N_27686,N_26450,N_25208);
xnor U27687 (N_27687,N_25450,N_26423);
xnor U27688 (N_27688,N_25719,N_26848);
xor U27689 (N_27689,N_25471,N_27106);
nand U27690 (N_27690,N_26503,N_26460);
xnor U27691 (N_27691,N_25756,N_25746);
and U27692 (N_27692,N_25040,N_25637);
nor U27693 (N_27693,N_26571,N_25790);
or U27694 (N_27694,N_26425,N_26504);
or U27695 (N_27695,N_26541,N_25429);
and U27696 (N_27696,N_25315,N_26453);
xnor U27697 (N_27697,N_25118,N_26355);
or U27698 (N_27698,N_27364,N_26727);
xnor U27699 (N_27699,N_25881,N_25533);
nand U27700 (N_27700,N_26096,N_26634);
or U27701 (N_27701,N_25961,N_27001);
xor U27702 (N_27702,N_25550,N_25205);
and U27703 (N_27703,N_26174,N_25826);
nor U27704 (N_27704,N_26602,N_25545);
nand U27705 (N_27705,N_25188,N_26612);
or U27706 (N_27706,N_26830,N_27167);
nand U27707 (N_27707,N_26466,N_25687);
nor U27708 (N_27708,N_25106,N_27326);
nand U27709 (N_27709,N_26478,N_26125);
xor U27710 (N_27710,N_25435,N_25206);
or U27711 (N_27711,N_26446,N_25806);
nand U27712 (N_27712,N_25444,N_27046);
nand U27713 (N_27713,N_26550,N_27282);
and U27714 (N_27714,N_25480,N_26097);
xor U27715 (N_27715,N_27332,N_25594);
and U27716 (N_27716,N_27253,N_25313);
nand U27717 (N_27717,N_26175,N_25918);
and U27718 (N_27718,N_25647,N_25842);
and U27719 (N_27719,N_26698,N_26890);
or U27720 (N_27720,N_26979,N_25690);
and U27721 (N_27721,N_26920,N_25034);
and U27722 (N_27722,N_25404,N_26393);
nand U27723 (N_27723,N_26048,N_25121);
nor U27724 (N_27724,N_26543,N_27107);
or U27725 (N_27725,N_25199,N_26064);
nand U27726 (N_27726,N_26353,N_27314);
or U27727 (N_27727,N_26462,N_25317);
or U27728 (N_27728,N_27447,N_26358);
xnor U27729 (N_27729,N_25841,N_25729);
and U27730 (N_27730,N_27099,N_25266);
nand U27731 (N_27731,N_25906,N_25725);
nor U27732 (N_27732,N_27110,N_25919);
or U27733 (N_27733,N_26077,N_25467);
nor U27734 (N_27734,N_27373,N_25692);
nor U27735 (N_27735,N_26985,N_25033);
nand U27736 (N_27736,N_26323,N_26059);
nor U27737 (N_27737,N_25005,N_26191);
or U27738 (N_27738,N_25308,N_26606);
and U27739 (N_27739,N_26418,N_27395);
and U27740 (N_27740,N_27004,N_25183);
nand U27741 (N_27741,N_27053,N_26169);
xnor U27742 (N_27742,N_25828,N_27397);
or U27743 (N_27743,N_26429,N_26116);
nor U27744 (N_27744,N_25999,N_25454);
nand U27745 (N_27745,N_25527,N_26562);
nand U27746 (N_27746,N_26224,N_26415);
xor U27747 (N_27747,N_27064,N_27018);
and U27748 (N_27748,N_25997,N_25736);
and U27749 (N_27749,N_26376,N_25343);
and U27750 (N_27750,N_26405,N_25529);
nand U27751 (N_27751,N_27009,N_25102);
nor U27752 (N_27752,N_26751,N_26513);
xnor U27753 (N_27753,N_25653,N_25138);
xnor U27754 (N_27754,N_26973,N_27118);
and U27755 (N_27755,N_26927,N_26705);
and U27756 (N_27756,N_26018,N_26468);
or U27757 (N_27757,N_27423,N_26702);
xnor U27758 (N_27758,N_27248,N_26672);
and U27759 (N_27759,N_26816,N_26032);
and U27760 (N_27760,N_25084,N_26857);
nor U27761 (N_27761,N_27116,N_26684);
nand U27762 (N_27762,N_26391,N_26995);
nor U27763 (N_27763,N_27435,N_27238);
nand U27764 (N_27764,N_26214,N_27379);
and U27765 (N_27765,N_25126,N_26469);
xnor U27766 (N_27766,N_27474,N_27133);
and U27767 (N_27767,N_27174,N_25245);
nand U27768 (N_27768,N_26828,N_25506);
and U27769 (N_27769,N_26225,N_26784);
or U27770 (N_27770,N_26964,N_26967);
nor U27771 (N_27771,N_27465,N_25466);
xor U27772 (N_27772,N_25609,N_26286);
or U27773 (N_27773,N_26072,N_25112);
nor U27774 (N_27774,N_25808,N_26020);
nand U27775 (N_27775,N_27198,N_26695);
and U27776 (N_27776,N_25789,N_27266);
nor U27777 (N_27777,N_25359,N_26568);
nand U27778 (N_27778,N_25156,N_27137);
and U27779 (N_27779,N_26365,N_27215);
nand U27780 (N_27780,N_26433,N_25489);
and U27781 (N_27781,N_26430,N_25283);
xnor U27782 (N_27782,N_25619,N_26369);
or U27783 (N_27783,N_25143,N_27020);
xnor U27784 (N_27784,N_25803,N_26863);
nor U27785 (N_27785,N_25171,N_26152);
nor U27786 (N_27786,N_26320,N_26551);
nor U27787 (N_27787,N_25244,N_26936);
and U27788 (N_27788,N_25669,N_27301);
and U27789 (N_27789,N_26189,N_25779);
or U27790 (N_27790,N_27281,N_26098);
nand U27791 (N_27791,N_26019,N_27230);
nand U27792 (N_27792,N_26975,N_25226);
or U27793 (N_27793,N_26790,N_26287);
xor U27794 (N_27794,N_25591,N_26713);
and U27795 (N_27795,N_27278,N_25078);
or U27796 (N_27796,N_27195,N_25470);
nor U27797 (N_27797,N_26304,N_27141);
nor U27798 (N_27798,N_26215,N_26157);
nor U27799 (N_27799,N_25329,N_26226);
and U27800 (N_27800,N_26199,N_25778);
or U27801 (N_27801,N_25772,N_25944);
and U27802 (N_27802,N_26998,N_26946);
nand U27803 (N_27803,N_27157,N_25402);
and U27804 (N_27804,N_26618,N_26147);
nand U27805 (N_27805,N_26136,N_25612);
xnor U27806 (N_27806,N_25998,N_25440);
or U27807 (N_27807,N_25885,N_26987);
xor U27808 (N_27808,N_26316,N_26813);
nor U27809 (N_27809,N_25794,N_25496);
xnor U27810 (N_27810,N_25295,N_25090);
nor U27811 (N_27811,N_26795,N_25864);
or U27812 (N_27812,N_26273,N_25544);
or U27813 (N_27813,N_25113,N_25272);
or U27814 (N_27814,N_25708,N_27045);
and U27815 (N_27815,N_25104,N_26485);
nand U27816 (N_27816,N_27036,N_25823);
xor U27817 (N_27817,N_26755,N_26027);
nor U27818 (N_27818,N_25222,N_25447);
nand U27819 (N_27819,N_26919,N_25198);
xor U27820 (N_27820,N_25049,N_25611);
or U27821 (N_27821,N_27458,N_25982);
nand U27822 (N_27822,N_25029,N_26587);
and U27823 (N_27823,N_27221,N_26603);
and U27824 (N_27824,N_26659,N_26194);
nand U27825 (N_27825,N_27269,N_25517);
nor U27826 (N_27826,N_25805,N_25328);
nor U27827 (N_27827,N_26655,N_26690);
xor U27828 (N_27828,N_25912,N_27264);
nor U27829 (N_27829,N_25010,N_26427);
xor U27830 (N_27830,N_25170,N_26743);
nand U27831 (N_27831,N_25107,N_25478);
xor U27832 (N_27832,N_26673,N_26342);
nand U27833 (N_27833,N_25981,N_27283);
or U27834 (N_27834,N_27480,N_26221);
xor U27835 (N_27835,N_25728,N_27444);
nor U27836 (N_27836,N_25978,N_27271);
nand U27837 (N_27837,N_25727,N_26283);
or U27838 (N_27838,N_27384,N_25371);
nor U27839 (N_27839,N_26888,N_25933);
and U27840 (N_27840,N_26477,N_25564);
and U27841 (N_27841,N_26664,N_26999);
or U27842 (N_27842,N_26829,N_27217);
nor U27843 (N_27843,N_26760,N_26660);
nor U27844 (N_27844,N_25853,N_25030);
nand U27845 (N_27845,N_25757,N_26663);
nand U27846 (N_27846,N_25388,N_26406);
or U27847 (N_27847,N_26281,N_27015);
or U27848 (N_27848,N_26781,N_25018);
or U27849 (N_27849,N_26874,N_25307);
or U27850 (N_27850,N_26216,N_25802);
nand U27851 (N_27851,N_26121,N_25396);
and U27852 (N_27852,N_25857,N_25325);
or U27853 (N_27853,N_25484,N_27154);
nand U27854 (N_27854,N_25665,N_26968);
nand U27855 (N_27855,N_25688,N_25320);
xnor U27856 (N_27856,N_27370,N_26421);
nand U27857 (N_27857,N_25290,N_25265);
xnor U27858 (N_27858,N_25066,N_26722);
or U27859 (N_27859,N_25661,N_27433);
and U27860 (N_27860,N_26101,N_25286);
nand U27861 (N_27861,N_25817,N_25520);
or U27862 (N_27862,N_26187,N_26780);
or U27863 (N_27863,N_25748,N_25570);
nand U27864 (N_27864,N_25753,N_27387);
and U27865 (N_27865,N_27124,N_27219);
nor U27866 (N_27866,N_26963,N_26183);
nand U27867 (N_27867,N_25500,N_25169);
nor U27868 (N_27868,N_25943,N_25414);
or U27869 (N_27869,N_25660,N_26611);
nor U27870 (N_27870,N_26017,N_25291);
or U27871 (N_27871,N_25993,N_25600);
or U27872 (N_27872,N_26088,N_25668);
and U27873 (N_27873,N_26288,N_25657);
xor U27874 (N_27874,N_26234,N_25696);
nor U27875 (N_27875,N_26881,N_27242);
xnor U27876 (N_27876,N_26507,N_26073);
or U27877 (N_27877,N_25749,N_26895);
nor U27878 (N_27878,N_27410,N_26815);
and U27879 (N_27879,N_26986,N_25972);
nand U27880 (N_27880,N_25991,N_25136);
nand U27881 (N_27881,N_26127,N_26605);
nand U27882 (N_27882,N_26213,N_25951);
xnor U27883 (N_27883,N_25344,N_26822);
or U27884 (N_27884,N_26056,N_27383);
or U27885 (N_27885,N_25253,N_27241);
or U27886 (N_27886,N_26653,N_26616);
xor U27887 (N_27887,N_26730,N_26681);
nand U27888 (N_27888,N_26710,N_26133);
or U27889 (N_27889,N_26024,N_25569);
nand U27890 (N_27890,N_27040,N_25758);
or U27891 (N_27891,N_25263,N_26918);
or U27892 (N_27892,N_25492,N_25073);
nor U27893 (N_27893,N_25896,N_25174);
nand U27894 (N_27894,N_26344,N_27443);
or U27895 (N_27895,N_27176,N_25097);
or U27896 (N_27896,N_27322,N_27002);
nand U27897 (N_27897,N_25571,N_26445);
or U27898 (N_27898,N_26516,N_26012);
nor U27899 (N_27899,N_25221,N_26720);
or U27900 (N_27900,N_26662,N_26724);
nor U27901 (N_27901,N_25588,N_27098);
nand U27902 (N_27902,N_26613,N_27330);
and U27903 (N_27903,N_26514,N_25767);
and U27904 (N_27904,N_25189,N_25336);
and U27905 (N_27905,N_26679,N_26801);
or U27906 (N_27906,N_27029,N_25921);
and U27907 (N_27907,N_26797,N_27087);
and U27908 (N_27908,N_26859,N_25887);
nand U27909 (N_27909,N_27464,N_25228);
xor U27910 (N_27910,N_25381,N_26495);
xnor U27911 (N_27911,N_27109,N_27280);
or U27912 (N_27912,N_25001,N_25192);
nand U27913 (N_27913,N_25045,N_25518);
nor U27914 (N_27914,N_25583,N_25132);
or U27915 (N_27915,N_25079,N_26230);
nor U27916 (N_27916,N_27345,N_26414);
or U27917 (N_27917,N_25081,N_26708);
nor U27918 (N_27918,N_27055,N_27371);
nand U27919 (N_27919,N_26437,N_26165);
nor U27920 (N_27920,N_27477,N_26176);
nor U27921 (N_27921,N_26715,N_27068);
or U27922 (N_27922,N_26493,N_25184);
or U27923 (N_27923,N_25093,N_26834);
or U27924 (N_27924,N_25065,N_27390);
nor U27925 (N_27925,N_25734,N_25764);
nor U27926 (N_27926,N_26519,N_27305);
nand U27927 (N_27927,N_25140,N_26915);
and U27928 (N_27928,N_26107,N_25515);
xor U27929 (N_27929,N_27228,N_25563);
or U27930 (N_27930,N_25990,N_26729);
nor U27931 (N_27931,N_27489,N_25644);
nor U27932 (N_27932,N_26172,N_25100);
xnor U27933 (N_27933,N_26026,N_26850);
nand U27934 (N_27934,N_25412,N_25379);
or U27935 (N_27935,N_26648,N_25195);
nand U27936 (N_27936,N_26509,N_26464);
and U27937 (N_27937,N_27000,N_27450);
xor U27938 (N_27938,N_26337,N_26604);
and U27939 (N_27939,N_25139,N_25063);
xnor U27940 (N_27940,N_27406,N_26989);
nor U27941 (N_27941,N_27359,N_25333);
or U27942 (N_27942,N_25760,N_26832);
and U27943 (N_27943,N_26961,N_26851);
and U27944 (N_27944,N_26232,N_27028);
xnor U27945 (N_27945,N_26518,N_26646);
or U27946 (N_27946,N_27250,N_26294);
nand U27947 (N_27947,N_27386,N_25128);
and U27948 (N_27948,N_27042,N_25481);
or U27949 (N_27949,N_27196,N_26845);
nand U27950 (N_27950,N_25491,N_27014);
and U27951 (N_27951,N_27333,N_27405);
xor U27952 (N_27952,N_27062,N_26545);
nor U27953 (N_27953,N_25540,N_26384);
nor U27954 (N_27954,N_26435,N_25992);
and U27955 (N_27955,N_25395,N_25819);
and U27956 (N_27956,N_27096,N_26794);
nor U27957 (N_27957,N_26884,N_26422);
nor U27958 (N_27958,N_26893,N_25087);
nor U27959 (N_27959,N_27057,N_26856);
xor U27960 (N_27960,N_25294,N_25262);
and U27961 (N_27961,N_26131,N_26035);
and U27962 (N_27962,N_27190,N_25119);
nand U27963 (N_27963,N_27051,N_26956);
and U27964 (N_27964,N_27255,N_26522);
or U27965 (N_27965,N_27439,N_26906);
and U27966 (N_27966,N_26547,N_25269);
xnor U27967 (N_27967,N_27358,N_26629);
and U27968 (N_27968,N_25144,N_26250);
nor U27969 (N_27969,N_25979,N_25516);
or U27970 (N_27970,N_25215,N_26268);
nand U27971 (N_27971,N_25676,N_25398);
or U27972 (N_27972,N_26909,N_25243);
nor U27973 (N_27973,N_25829,N_25838);
nand U27974 (N_27974,N_25085,N_26295);
nand U27975 (N_27975,N_26528,N_25069);
or U27976 (N_27976,N_26340,N_25193);
nand U27977 (N_27977,N_25432,N_27294);
nor U27978 (N_27978,N_27499,N_27491);
nand U27979 (N_27979,N_25791,N_26506);
and U27980 (N_27980,N_27034,N_25249);
nand U27981 (N_27981,N_27428,N_26951);
nand U27982 (N_27982,N_26397,N_26314);
xor U27983 (N_27983,N_26758,N_27211);
and U27984 (N_27984,N_25370,N_25186);
and U27985 (N_27985,N_26669,N_25781);
and U27986 (N_27986,N_27418,N_27394);
nand U27987 (N_27987,N_25009,N_26552);
xnor U27988 (N_27988,N_26817,N_27475);
nor U27989 (N_27989,N_27338,N_25098);
nor U27990 (N_27990,N_27091,N_26969);
or U27991 (N_27991,N_27347,N_25129);
nand U27992 (N_27992,N_26517,N_26879);
or U27993 (N_27993,N_27187,N_26307);
or U27994 (N_27994,N_25133,N_26390);
or U27995 (N_27995,N_27100,N_26650);
or U27996 (N_27996,N_25623,N_25177);
or U27997 (N_27997,N_25761,N_26266);
and U27998 (N_27998,N_25234,N_27177);
nor U27999 (N_27999,N_26510,N_26324);
or U28000 (N_28000,N_27210,N_26990);
xnor U28001 (N_28001,N_26410,N_26045);
nand U28002 (N_28002,N_26357,N_26092);
xnor U28003 (N_28003,N_25347,N_25542);
nor U28004 (N_28004,N_25877,N_25413);
or U28005 (N_28005,N_26105,N_26196);
and U28006 (N_28006,N_25858,N_25714);
and U28007 (N_28007,N_27012,N_27341);
xor U28008 (N_28008,N_25083,N_26326);
nor U28009 (N_28009,N_25769,N_25920);
nand U28010 (N_28010,N_25710,N_26382);
or U28011 (N_28011,N_27247,N_26118);
nor U28012 (N_28012,N_25421,N_26263);
or U28013 (N_28013,N_25519,N_27071);
nand U28014 (N_28014,N_25309,N_26043);
xnor U28015 (N_28015,N_26068,N_26188);
or U28016 (N_28016,N_27377,N_26484);
or U28017 (N_28017,N_26463,N_27035);
nor U28018 (N_28018,N_26443,N_26370);
or U28019 (N_28019,N_25182,N_26746);
xnor U28020 (N_28020,N_26624,N_27229);
and U28021 (N_28021,N_25123,N_27461);
or U28022 (N_28022,N_25827,N_27298);
or U28023 (N_28023,N_25051,N_26911);
and U28024 (N_28024,N_27289,N_27076);
nor U28025 (N_28025,N_25865,N_26748);
nor U28026 (N_28026,N_26039,N_25196);
xnor U28027 (N_28027,N_27212,N_25530);
or U28028 (N_28028,N_25930,N_27237);
nand U28029 (N_28029,N_25486,N_25080);
nand U28030 (N_28030,N_27408,N_27292);
or U28031 (N_28031,N_27369,N_26942);
nor U28032 (N_28032,N_27194,N_25792);
nor U28033 (N_28033,N_26886,N_26827);
or U28034 (N_28034,N_26738,N_25952);
or U28035 (N_28035,N_27327,N_25942);
nand U28036 (N_28036,N_27146,N_25037);
nand U28037 (N_28037,N_26292,N_26346);
or U28038 (N_28038,N_26529,N_26661);
and U28039 (N_28039,N_25645,N_25130);
nor U28040 (N_28040,N_25312,N_26299);
nor U28041 (N_28041,N_26589,N_25111);
nor U28042 (N_28042,N_26959,N_25386);
and U28043 (N_28043,N_25020,N_25574);
nand U28044 (N_28044,N_25348,N_25305);
and U28045 (N_28045,N_27003,N_25726);
or U28046 (N_28046,N_25296,N_25524);
nor U28047 (N_28047,N_25705,N_25439);
and U28048 (N_28048,N_25573,N_26413);
nand U28049 (N_28049,N_25552,N_25946);
and U28050 (N_28050,N_27285,N_27125);
xor U28051 (N_28051,N_25255,N_26246);
xor U28052 (N_28052,N_25026,N_26347);
nand U28053 (N_28053,N_25423,N_27169);
or U28054 (N_28054,N_25147,N_25595);
and U28055 (N_28055,N_25089,N_25462);
or U28056 (N_28056,N_25239,N_25597);
nand U28057 (N_28057,N_25566,N_26941);
or U28058 (N_28058,N_25476,N_26178);
or U28059 (N_28059,N_25211,N_25161);
and U28060 (N_28060,N_27324,N_26306);
nand U28061 (N_28061,N_26312,N_27457);
or U28062 (N_28062,N_26310,N_26334);
or U28063 (N_28063,N_25816,N_25397);
nor U28064 (N_28064,N_26082,N_26338);
xnor U28065 (N_28065,N_27380,N_25225);
xor U28066 (N_28066,N_26436,N_26336);
or U28067 (N_28067,N_25456,N_25273);
nor U28068 (N_28068,N_25375,N_26614);
nand U28069 (N_28069,N_26692,N_26536);
and U28070 (N_28070,N_27260,N_26497);
or U28071 (N_28071,N_26471,N_25958);
nand U28072 (N_28072,N_26523,N_25768);
or U28073 (N_28073,N_25883,N_25490);
and U28074 (N_28074,N_26734,N_27427);
or U28075 (N_28075,N_27470,N_25254);
nand U28076 (N_28076,N_25219,N_25625);
nand U28077 (N_28077,N_25314,N_26109);
or U28078 (N_28078,N_27246,N_26527);
and U28079 (N_28079,N_25418,N_27275);
nor U28080 (N_28080,N_26219,N_27265);
xor U28081 (N_28081,N_26579,N_26965);
xor U28082 (N_28082,N_25795,N_26426);
xnor U28083 (N_28083,N_26654,N_26594);
and U28084 (N_28084,N_27344,N_26386);
nor U28085 (N_28085,N_26952,N_25003);
or U28086 (N_28086,N_26235,N_26298);
xor U28087 (N_28087,N_26047,N_27161);
and U28088 (N_28088,N_26804,N_26163);
and U28089 (N_28089,N_27163,N_27297);
xor U28090 (N_28090,N_25664,N_26499);
and U28091 (N_28091,N_26474,N_25054);
or U28092 (N_28092,N_25194,N_26553);
xnor U28093 (N_28093,N_27058,N_25292);
nor U28094 (N_28094,N_26778,N_27069);
nor U28095 (N_28095,N_27420,N_25586);
and U28096 (N_28096,N_25884,N_26577);
or U28097 (N_28097,N_27153,N_26860);
and U28098 (N_28098,N_25852,N_25067);
nand U28099 (N_28099,N_26244,N_25900);
nand U28100 (N_28100,N_27478,N_26526);
nor U28101 (N_28101,N_26754,N_27473);
or U28102 (N_28102,N_26209,N_27239);
or U28103 (N_28103,N_25622,N_26524);
nor U28104 (N_28104,N_25274,N_27218);
nor U28105 (N_28105,N_26623,N_27469);
xnor U28106 (N_28106,N_26864,N_26277);
nor U28107 (N_28107,N_26566,N_26771);
nand U28108 (N_28108,N_26256,N_26937);
nand U28109 (N_28109,N_25717,N_25043);
and U28110 (N_28110,N_25974,N_27206);
or U28111 (N_28111,N_26707,N_27173);
nor U28112 (N_28112,N_26880,N_27436);
or U28113 (N_28113,N_27245,N_27052);
and U28114 (N_28114,N_26670,N_26069);
nand U28115 (N_28115,N_26318,N_26675);
or U28116 (N_28116,N_26558,N_25537);
nor U28117 (N_28117,N_25701,N_26597);
nor U28118 (N_28118,N_27466,N_27140);
and U28119 (N_28119,N_26668,N_25382);
and U28120 (N_28120,N_27019,N_25154);
xnor U28121 (N_28121,N_27366,N_26538);
nand U28122 (N_28122,N_26570,N_27268);
xor U28123 (N_28123,N_27152,N_25207);
or U28124 (N_28124,N_25504,N_26275);
nand U28125 (N_28125,N_25836,N_25300);
nand U28126 (N_28126,N_26134,N_25536);
or U28127 (N_28127,N_26062,N_27398);
or U28128 (N_28128,N_26737,N_25543);
or U28129 (N_28129,N_25848,N_26345);
nor U28130 (N_28130,N_25926,N_25913);
or U28131 (N_28131,N_25535,N_27008);
and U28132 (N_28132,N_25546,N_26428);
or U28133 (N_28133,N_25917,N_27193);
xnor U28134 (N_28134,N_26104,N_25616);
or U28135 (N_28135,N_26392,N_26687);
nor U28136 (N_28136,N_26251,N_26628);
nor U28137 (N_28137,N_27425,N_25458);
nor U28138 (N_28138,N_26388,N_26789);
and U28139 (N_28139,N_26434,N_26953);
nand U28140 (N_28140,N_27006,N_25916);
nor U28141 (N_28141,N_25331,N_25902);
and U28142 (N_28142,N_27340,N_26486);
nor U28143 (N_28143,N_26716,N_27414);
xnor U28144 (N_28144,N_25567,N_26142);
xor U28145 (N_28145,N_26278,N_26015);
nand U28146 (N_28146,N_25072,N_25289);
nand U28147 (N_28147,N_25811,N_26882);
or U28148 (N_28148,N_27468,N_25461);
nand U28149 (N_28149,N_25633,N_26945);
and U28150 (N_28150,N_25815,N_26006);
nor U28151 (N_28151,N_27063,N_27027);
or U28152 (N_28152,N_25782,N_26401);
or U28153 (N_28153,N_25606,N_25762);
nor U28154 (N_28154,N_26617,N_26253);
nor U28155 (N_28155,N_25431,N_27316);
nor U28156 (N_28156,N_26501,N_25765);
nor U28157 (N_28157,N_25202,N_27117);
xor U28158 (N_28158,N_26981,N_26626);
nor U28159 (N_28159,N_27399,N_25356);
or U28160 (N_28160,N_27348,N_26091);
and U28161 (N_28161,N_25477,N_26563);
nor U28162 (N_28162,N_27227,N_27456);
or U28163 (N_28163,N_26800,N_25256);
nand U28164 (N_28164,N_25297,N_26598);
nor U28165 (N_28165,N_26100,N_26887);
nor U28166 (N_28166,N_25777,N_25754);
nand U28167 (N_28167,N_25341,N_26682);
and U28168 (N_28168,N_26820,N_27066);
and U28169 (N_28169,N_25363,N_25425);
or U28170 (N_28170,N_25585,N_25443);
or U28171 (N_28171,N_26117,N_27424);
or U28172 (N_28172,N_25862,N_25389);
nand U28173 (N_28173,N_25038,N_25210);
nand U28174 (N_28174,N_25793,N_25640);
xnor U28175 (N_28175,N_25741,N_26700);
or U28176 (N_28176,N_25966,N_25590);
or U28177 (N_28177,N_26185,N_26877);
or U28178 (N_28178,N_25070,N_27256);
xor U28179 (N_28179,N_26739,N_26944);
nand U28180 (N_28180,N_25582,N_26054);
nand U28181 (N_28181,N_25148,N_25759);
xnor U28182 (N_28182,N_25630,N_25434);
or U28183 (N_28183,N_25217,N_25967);
or U28184 (N_28184,N_26233,N_26071);
nor U28185 (N_28185,N_25892,N_27132);
xor U28186 (N_28186,N_27490,N_25891);
nand U28187 (N_28187,N_27378,N_26377);
and U28188 (N_28188,N_25430,N_25587);
and U28189 (N_28189,N_25326,N_26619);
nor U28190 (N_28190,N_26135,N_26631);
and U28191 (N_28191,N_26011,N_25751);
xnor U28192 (N_28192,N_27372,N_25742);
xor U28193 (N_28193,N_26498,N_25446);
xor U28194 (N_28194,N_26677,N_25821);
and U28195 (N_28195,N_26704,N_25786);
nand U28196 (N_28196,N_27415,N_26124);
and U28197 (N_28197,N_25820,N_25763);
xor U28198 (N_28198,N_26033,N_25956);
nor U28199 (N_28199,N_26258,N_25299);
nand U28200 (N_28200,N_25361,N_26067);
nand U28201 (N_28201,N_27070,N_25702);
or U28202 (N_28202,N_26137,N_25372);
xor U28203 (N_28203,N_26939,N_25565);
nor U28204 (N_28204,N_27375,N_25023);
or U28205 (N_28205,N_25145,N_26544);
nand U28206 (N_28206,N_26441,N_26930);
xnor U28207 (N_28207,N_27065,N_27113);
or U28208 (N_28208,N_26398,N_25392);
nand U28209 (N_28209,N_25699,N_27317);
or U28210 (N_28210,N_27485,N_26195);
nand U28211 (N_28211,N_25187,N_25351);
nor U28212 (N_28212,N_26297,N_26792);
or U28213 (N_28213,N_27312,N_26128);
or U28214 (N_28214,N_27024,N_25596);
and U28215 (N_28215,N_25349,N_26590);
or U28216 (N_28216,N_26279,N_25216);
xor U28217 (N_28217,N_25427,N_25127);
xnor U28218 (N_28218,N_25288,N_25988);
xnor U28219 (N_28219,N_25575,N_26249);
nor U28220 (N_28220,N_26756,N_26638);
xor U28221 (N_28221,N_27179,N_26761);
xor U28222 (N_28222,N_25316,N_25532);
nand U28223 (N_28223,N_27083,N_27130);
or U28224 (N_28224,N_25643,N_25713);
xnor U28225 (N_28225,N_25977,N_26824);
xor U28226 (N_28226,N_25134,N_26160);
xnor U28227 (N_28227,N_26855,N_25453);
xor U28228 (N_28228,N_27182,N_26481);
and U28229 (N_28229,N_25488,N_26036);
or U28230 (N_28230,N_27095,N_25082);
and U28231 (N_28231,N_26933,N_26898);
xor U28232 (N_28232,N_25876,N_26237);
or U28233 (N_28233,N_26291,N_25551);
and U28234 (N_28234,N_27482,N_27445);
and U28235 (N_28235,N_25160,N_26052);
nand U28236 (N_28236,N_26359,N_26639);
and U28237 (N_28237,N_26854,N_25366);
nand U28238 (N_28238,N_27234,N_25562);
and U28239 (N_28239,N_25834,N_26005);
and U28240 (N_28240,N_26805,N_27093);
or U28241 (N_28241,N_26458,N_25417);
and U28242 (N_28242,N_25058,N_27323);
nand U28243 (N_28243,N_25159,N_25605);
and U28244 (N_28244,N_26731,N_25362);
nand U28245 (N_28245,N_25464,N_26330);
nor U28246 (N_28246,N_26599,N_27175);
xnor U28247 (N_28247,N_25497,N_26575);
nor U28248 (N_28248,N_26728,N_26095);
nor U28249 (N_28249,N_25553,N_25939);
or U28250 (N_28250,N_26122,N_26144);
nor U28251 (N_28251,N_25135,N_26455);
xnor U28252 (N_28252,N_26080,N_25592);
xor U28253 (N_28253,N_25235,N_26111);
nand U28254 (N_28254,N_26372,N_26350);
and U28255 (N_28255,N_27321,N_26274);
xnor U28256 (N_28256,N_26184,N_25014);
xnor U28257 (N_28257,N_25346,N_26385);
nor U28258 (N_28258,N_26149,N_26957);
and U28259 (N_28259,N_26803,N_26055);
and U28260 (N_28260,N_27431,N_26853);
nor U28261 (N_28261,N_25549,N_26861);
nand U28262 (N_28262,N_25495,N_27336);
nand U28263 (N_28263,N_26935,N_26354);
xnor U28264 (N_28264,N_27440,N_26439);
and U28265 (N_28265,N_25812,N_25579);
or U28266 (N_28266,N_26057,N_26231);
and U28267 (N_28267,N_27303,N_26849);
nor U28268 (N_28268,N_26028,N_26181);
nor U28269 (N_28269,N_27074,N_26061);
or U28270 (N_28270,N_26085,N_25510);
and U28271 (N_28271,N_25953,N_26361);
nor U28272 (N_28272,N_27493,N_26885);
and U28273 (N_28273,N_26644,N_26988);
nand U28274 (N_28274,N_25905,N_26984);
nor U28275 (N_28275,N_27365,N_26228);
or U28276 (N_28276,N_25561,N_27200);
nor U28277 (N_28277,N_25783,N_25584);
and U28278 (N_28278,N_27350,N_25498);
nor U28279 (N_28279,N_27360,N_27362);
nor U28280 (N_28280,N_27476,N_25062);
xnor U28281 (N_28281,N_27115,N_27302);
nand U28282 (N_28282,N_27081,N_26534);
and U28283 (N_28283,N_25843,N_26240);
xnor U28284 (N_28284,N_25149,N_26356);
and U28285 (N_28285,N_26787,N_25825);
xnor U28286 (N_28286,N_25122,N_27315);
and U28287 (N_28287,N_25950,N_25166);
and U28288 (N_28288,N_25888,N_27328);
or U28289 (N_28289,N_25203,N_25908);
and U28290 (N_28290,N_27313,N_25311);
nor U28291 (N_28291,N_25365,N_27047);
or U28292 (N_28292,N_25460,N_25276);
and U28293 (N_28293,N_27170,N_25452);
and U28294 (N_28294,N_26349,N_25830);
nand U28295 (N_28295,N_26186,N_25752);
nand U28296 (N_28296,N_26866,N_25968);
xnor U28297 (N_28297,N_26106,N_27421);
or U28298 (N_28298,N_25261,N_25424);
nor U28299 (N_28299,N_26153,N_27481);
and U28300 (N_28300,N_26978,N_25190);
xnor U28301 (N_28301,N_26685,N_26201);
xor U28302 (N_28302,N_25773,N_26697);
or U28303 (N_28303,N_27136,N_25511);
nor U28304 (N_28304,N_27363,N_25755);
nand U28305 (N_28305,N_25733,N_27498);
nor U28306 (N_28306,N_26633,N_26699);
xor U28307 (N_28307,N_26539,N_25882);
or U28308 (N_28308,N_25850,N_26473);
xnor U28309 (N_28309,N_27446,N_26572);
xor U28310 (N_28310,N_25576,N_26496);
nor U28311 (N_28311,N_26383,N_27235);
or U28312 (N_28312,N_26560,N_25539);
and U28313 (N_28313,N_25180,N_25258);
or U28314 (N_28314,N_26053,N_27257);
nor U28315 (N_28315,N_26162,N_26678);
or U28316 (N_28316,N_25044,N_26396);
and U28317 (N_28317,N_27309,N_25384);
xnor U28318 (N_28318,N_26582,N_25330);
and U28319 (N_28319,N_27126,N_27416);
and U28320 (N_28320,N_25280,N_25278);
xnor U28321 (N_28321,N_26875,N_26757);
nand U28322 (N_28322,N_27407,N_25872);
nor U28323 (N_28323,N_25904,N_25634);
or U28324 (N_28324,N_26179,N_26745);
xor U28325 (N_28325,N_25547,N_27135);
nand U28326 (N_28326,N_27078,N_25938);
xnor U28327 (N_28327,N_25285,N_25948);
xnor U28328 (N_28328,N_26733,N_27112);
nand U28329 (N_28329,N_25648,N_25680);
or U28330 (N_28330,N_26023,N_26505);
and U28331 (N_28331,N_26502,N_26046);
nor U28332 (N_28332,N_25247,N_25889);
and U28333 (N_28333,N_26609,N_26198);
nand U28334 (N_28334,N_27335,N_26029);
nor U28335 (N_28335,N_25873,N_25451);
nand U28336 (N_28336,N_26371,N_25813);
nor U28337 (N_28337,N_26726,N_25011);
or U28338 (N_28338,N_27180,N_25377);
nor U28339 (N_28339,N_25835,N_27155);
nor U28340 (N_28340,N_26955,N_26366);
xnor U28341 (N_28341,N_26564,N_25740);
and U28342 (N_28342,N_25201,N_26565);
nand U28343 (N_28343,N_27092,N_26686);
nand U28344 (N_28344,N_25621,N_26472);
xnor U28345 (N_28345,N_25947,N_26826);
xor U28346 (N_28346,N_27376,N_25744);
xor U28347 (N_28347,N_25335,N_26578);
nor U28348 (N_28348,N_25807,N_26621);
and U28349 (N_28349,N_25851,N_26139);
and U28350 (N_28350,N_25173,N_25814);
and U28351 (N_28351,N_25338,N_26688);
nor U28352 (N_28352,N_26368,N_25869);
xor U28353 (N_28353,N_25155,N_27320);
nand U28354 (N_28354,N_26058,N_25408);
nand U28355 (N_28355,N_27199,N_26050);
or U28356 (N_28356,N_26835,N_25059);
nand U28357 (N_28357,N_26922,N_25650);
nand U28358 (N_28358,N_26269,N_26764);
and U28359 (N_28359,N_25380,N_26532);
xor U28360 (N_28360,N_27148,N_26271);
nor U28361 (N_28361,N_25934,N_26093);
nand U28362 (N_28362,N_25419,N_26900);
nor U28363 (N_28363,N_26763,N_27159);
and U28364 (N_28364,N_27060,N_25879);
nand U28365 (N_28365,N_26712,N_26025);
xnor U28366 (N_28366,N_25035,N_27374);
and U28367 (N_28367,N_25164,N_27318);
and U28368 (N_28368,N_27441,N_25004);
or U28369 (N_28369,N_25684,N_25376);
xor U28370 (N_28370,N_26335,N_27178);
and U28371 (N_28371,N_25008,N_26168);
xor U28372 (N_28372,N_25124,N_27402);
xnor U28373 (N_28373,N_27189,N_25800);
nor U28374 (N_28374,N_27072,N_25581);
xor U28375 (N_28375,N_25013,N_25964);
or U28376 (N_28376,N_26925,N_26774);
nor U28377 (N_28377,N_26588,N_26940);
nor U28378 (N_28378,N_25505,N_25711);
and U28379 (N_28379,N_25743,N_25077);
or U28380 (N_28380,N_25282,N_25775);
or U28381 (N_28381,N_26924,N_26412);
nand U28382 (N_28382,N_26878,N_26561);
and U28383 (N_28383,N_25989,N_26869);
nor U28384 (N_28384,N_25831,N_25867);
nor U28385 (N_28385,N_26220,N_26099);
and U28386 (N_28386,N_25321,N_25319);
nand U28387 (N_28387,N_25391,N_25845);
xor U28388 (N_28388,N_25167,N_25209);
or U28389 (N_28389,N_27128,N_26280);
nor U28390 (N_28390,N_27460,N_26645);
xnor U28391 (N_28391,N_25832,N_27075);
and U28392 (N_28392,N_26926,N_25620);
nor U28393 (N_28393,N_26416,N_26075);
nor U28394 (N_28394,N_27346,N_27419);
nand U28395 (N_28395,N_25522,N_25538);
xor U28396 (N_28396,N_27236,N_26021);
nand U28397 (N_28397,N_26010,N_27226);
nand U28398 (N_28398,N_26452,N_25142);
nor U28399 (N_28399,N_25682,N_25677);
nand U28400 (N_28400,N_26765,N_26592);
nand U28401 (N_28401,N_27031,N_27396);
nor U28402 (N_28402,N_26210,N_26711);
and U28403 (N_28403,N_27119,N_26709);
nor U28404 (N_28404,N_27097,N_27342);
or U28405 (N_28405,N_26013,N_25512);
and U28406 (N_28406,N_25191,N_27288);
nand U28407 (N_28407,N_25632,N_26222);
and U28408 (N_28408,N_27488,N_26146);
and U28409 (N_28409,N_26389,N_25703);
nand U28410 (N_28410,N_26742,N_27351);
nor U28411 (N_28411,N_26947,N_25957);
nand U28412 (N_28412,N_25248,N_27279);
and U28413 (N_28413,N_25103,N_26831);
nand U28414 (N_28414,N_25162,N_26156);
nor U28415 (N_28415,N_26112,N_25383);
nor U28416 (N_28416,N_26367,N_27188);
nand U28417 (N_28417,N_27483,N_26837);
or U28418 (N_28418,N_26331,N_26203);
or U28419 (N_28419,N_26962,N_25604);
or U28420 (N_28420,N_25448,N_26044);
nor U28421 (N_28421,N_25875,N_26693);
xor U28422 (N_28422,N_26103,N_26317);
or U28423 (N_28423,N_26060,N_25659);
xor U28424 (N_28424,N_26002,N_25931);
nor U28425 (N_28425,N_26308,N_25493);
and U28426 (N_28426,N_27007,N_26456);
xnor U28427 (N_28427,N_26512,N_27296);
nand U28428 (N_28428,N_26252,N_26928);
or U28429 (N_28429,N_26719,N_26475);
or U28430 (N_28430,N_25722,N_26843);
nand U28431 (N_28431,N_26921,N_26783);
nor U28432 (N_28432,N_25886,N_26159);
and U28433 (N_28433,N_27304,N_27273);
nand U28434 (N_28434,N_26343,N_27295);
xor U28435 (N_28435,N_26302,N_27484);
nor U28436 (N_28436,N_25739,N_26491);
xnor U28437 (N_28437,N_26776,N_26773);
nor U28438 (N_28438,N_25465,N_25658);
nand U28439 (N_28439,N_25681,N_27214);
nand U28440 (N_28440,N_25863,N_25236);
xor U28441 (N_28441,N_26809,N_25787);
or U28442 (N_28442,N_27451,N_26740);
nand U28443 (N_28443,N_26665,N_25709);
nor U28444 (N_28444,N_26325,N_25878);
and U28445 (N_28445,N_26479,N_26508);
or U28446 (N_28446,N_25075,N_27391);
or U28447 (N_28447,N_27449,N_25036);
xor U28448 (N_28448,N_26255,N_27061);
nand U28449 (N_28449,N_25350,N_26996);
nand U28450 (N_28450,N_27361,N_25799);
xnor U28451 (N_28451,N_25560,N_25922);
nor U28452 (N_28452,N_26407,N_27357);
nor U28453 (N_28453,N_25459,N_25893);
and U28454 (N_28454,N_26852,N_26276);
xnor U28455 (N_28455,N_26042,N_26899);
xnor U28456 (N_28456,N_25855,N_25694);
xor U28457 (N_28457,N_25635,N_26248);
nand U28458 (N_28458,N_26636,N_26753);
or U28459 (N_28459,N_26810,N_27158);
nand U28460 (N_28460,N_26197,N_27032);
xnor U28461 (N_28461,N_25437,N_25973);
xor U28462 (N_28462,N_26844,N_27310);
and U28463 (N_28463,N_26649,N_25027);
nand U28464 (N_28464,N_25501,N_27085);
xnor U28465 (N_28465,N_26657,N_26090);
or U28466 (N_28466,N_26483,N_26736);
nor U28467 (N_28467,N_27392,N_26808);
nand U28468 (N_28468,N_27240,N_26408);
xnor U28469 (N_28469,N_27261,N_26932);
and U28470 (N_28470,N_25306,N_25387);
nand U28471 (N_28471,N_25108,N_25357);
xor U28472 (N_28472,N_25105,N_25120);
or U28473 (N_28473,N_25629,N_26000);
xnor U28474 (N_28474,N_25252,N_27181);
and U28475 (N_28475,N_25955,N_25693);
nor U28476 (N_28476,N_25983,N_26917);
or U28477 (N_28477,N_25903,N_25064);
nor U28478 (N_28478,N_27389,N_26714);
xor U28479 (N_28479,N_25364,N_25479);
nor U28480 (N_28480,N_26150,N_25302);
nor U28481 (N_28481,N_26193,N_26360);
xor U28482 (N_28482,N_26741,N_26520);
and U28483 (N_28483,N_27164,N_25281);
and U28484 (N_28484,N_26218,N_27233);
or U28485 (N_28485,N_27145,N_27277);
nand U28486 (N_28486,N_26931,N_26689);
nor U28487 (N_28487,N_25047,N_27108);
nand U28488 (N_28488,N_25116,N_25141);
and U28489 (N_28489,N_25152,N_27171);
xor U28490 (N_28490,N_25176,N_26759);
and U28491 (N_28491,N_26791,N_25631);
nand U28492 (N_28492,N_25627,N_27426);
nand U28493 (N_28493,N_25007,N_25055);
nor U28494 (N_28494,N_27186,N_27105);
nor U28495 (N_28495,N_26902,N_27150);
nand U28496 (N_28496,N_26192,N_25624);
or U28497 (N_28497,N_25031,N_25935);
nand U28498 (N_28498,N_27142,N_26490);
and U28499 (N_28499,N_27203,N_25554);
nand U28500 (N_28500,N_26257,N_26839);
or U28501 (N_28501,N_26819,N_25185);
and U28502 (N_28502,N_25407,N_26151);
or U28503 (N_28503,N_27102,N_26375);
nor U28504 (N_28504,N_25541,N_27073);
xor U28505 (N_28505,N_25723,N_25548);
xnor U28506 (N_28506,N_25735,N_25601);
xor U28507 (N_28507,N_26489,N_26903);
and U28508 (N_28508,N_26449,N_26305);
or U28509 (N_28509,N_25181,N_26910);
nand U28510 (N_28510,N_25178,N_27263);
and U28511 (N_28511,N_25367,N_25339);
and U28512 (N_28512,N_26037,N_26123);
and U28513 (N_28513,N_27311,N_27044);
xor U28514 (N_28514,N_25962,N_26442);
nand U28515 (N_28515,N_25963,N_25969);
xnor U28516 (N_28516,N_25771,N_26701);
and U28517 (N_28517,N_26236,N_26267);
nor U28518 (N_28518,N_26825,N_25340);
xor U28519 (N_28519,N_25436,N_25502);
and U28520 (N_28520,N_27134,N_25649);
nand U28521 (N_28521,N_27192,N_25844);
nor U28522 (N_28522,N_25057,N_27138);
nand U28523 (N_28523,N_27459,N_25224);
nand U28524 (N_28524,N_26272,N_26007);
or U28525 (N_28525,N_25150,N_25923);
nor U28526 (N_28526,N_27388,N_25337);
or U28527 (N_28527,N_26440,N_26958);
nand U28528 (N_28528,N_27026,N_26647);
nand U28529 (N_28529,N_26557,N_25233);
nand U28530 (N_28530,N_27287,N_26601);
or U28531 (N_28531,N_26718,N_25475);
nor U28532 (N_28532,N_26515,N_27306);
nor U28533 (N_28533,N_25698,N_26694);
and U28534 (N_28534,N_27103,N_25854);
nand U28535 (N_28535,N_27232,N_26833);
nor U28536 (N_28536,N_26767,N_25531);
nand U28537 (N_28537,N_26115,N_27021);
or U28538 (N_28538,N_26581,N_26889);
nand U28539 (N_28539,N_25022,N_27254);
or U28540 (N_28540,N_26031,N_26559);
xnor U28541 (N_28541,N_25503,N_25237);
or U28542 (N_28542,N_26114,N_26846);
nand U28543 (N_28543,N_26546,N_26786);
nand U28544 (N_28544,N_27486,N_27487);
nand U28545 (N_28545,N_27251,N_25369);
nand U28546 (N_28546,N_27191,N_26537);
or U28547 (N_28547,N_25712,N_25469);
or U28548 (N_28548,N_27244,N_26040);
and U28549 (N_28549,N_26744,N_25096);
xnor U28550 (N_28550,N_27123,N_25378);
nand U28551 (N_28551,N_27223,N_25092);
nor U28552 (N_28552,N_25678,N_26980);
nor U28553 (N_28553,N_26403,N_26465);
and U28554 (N_28554,N_25925,N_25639);
nor U28555 (N_28555,N_27005,N_26078);
and U28556 (N_28556,N_27084,N_26285);
or U28557 (N_28557,N_26461,N_25932);
xor U28558 (N_28558,N_25914,N_27129);
or U28559 (N_28559,N_25508,N_25259);
nor U28560 (N_28560,N_25399,N_26912);
or U28561 (N_28561,N_26094,N_26766);
or U28562 (N_28562,N_27290,N_25730);
or U28563 (N_28563,N_26870,N_26873);
nand U28564 (N_28564,N_26821,N_26132);
nand U28565 (N_28565,N_25662,N_25250);
nand U28566 (N_28566,N_27037,N_27184);
xnor U28567 (N_28567,N_26086,N_27454);
nand U28568 (N_28568,N_27082,N_27114);
xnor U28569 (N_28569,N_25251,N_27267);
nand U28570 (N_28570,N_27025,N_26087);
and U28571 (N_28571,N_26901,N_25975);
and U28572 (N_28572,N_25472,N_25114);
nand U28573 (N_28573,N_25019,N_27151);
nor U28574 (N_28574,N_27160,N_27299);
and U28575 (N_28575,N_26872,N_27356);
and U28576 (N_28576,N_25355,N_27204);
and U28577 (N_28577,N_26074,N_26066);
nor U28578 (N_28578,N_25901,N_26313);
and U28579 (N_28579,N_26488,N_26793);
xor U28580 (N_28580,N_26865,N_26145);
nand U28581 (N_28581,N_25131,N_26904);
nand U28582 (N_28582,N_25046,N_26217);
nand U28583 (N_28583,N_26812,N_27448);
xnor U28584 (N_28584,N_25277,N_26777);
nand U28585 (N_28585,N_27147,N_25580);
xnor U28586 (N_28586,N_25028,N_26782);
nand U28587 (N_28587,N_27382,N_26747);
nor U28588 (N_28588,N_26954,N_26683);
and U28589 (N_28589,N_26977,N_27404);
xnor U28590 (N_28590,N_26785,N_25220);
nand U28591 (N_28591,N_26182,N_26530);
nand U28592 (N_28592,N_25240,N_27168);
and U28593 (N_28593,N_26641,N_26282);
xnor U28594 (N_28594,N_26138,N_25718);
and U28595 (N_28595,N_25785,N_26836);
and U28596 (N_28596,N_27162,N_25214);
nand U28597 (N_28597,N_25766,N_27308);
nand U28598 (N_28598,N_25068,N_26158);
nand U28599 (N_28599,N_25405,N_25071);
and U28600 (N_28600,N_25824,N_25212);
xnor U28601 (N_28601,N_27430,N_26190);
xnor U28602 (N_28602,N_27216,N_26635);
nor U28603 (N_28603,N_26380,N_25894);
and U28604 (N_28604,N_27127,N_25017);
or U28605 (N_28605,N_25732,N_25499);
or U28606 (N_28606,N_25673,N_25555);
and U28607 (N_28607,N_25837,N_25279);
xor U28608 (N_28608,N_25599,N_27050);
and U28609 (N_28609,N_26620,N_25774);
or U28610 (N_28610,N_27243,N_26656);
xnor U28611 (N_28611,N_26038,N_25750);
nor U28612 (N_28612,N_26166,N_26651);
nor U28613 (N_28613,N_25410,N_25895);
nor U28614 (N_28614,N_27225,N_26049);
xnor U28615 (N_28615,N_26976,N_26938);
and U28616 (N_28616,N_26750,N_25390);
nor U28617 (N_28617,N_25422,N_26420);
xor U28618 (N_28618,N_25685,N_26332);
or U28619 (N_28619,N_27343,N_26806);
or U28620 (N_28620,N_25088,N_27088);
xor U28621 (N_28621,N_26120,N_26003);
and U28622 (N_28622,N_25880,N_26260);
and U28623 (N_28623,N_26721,N_26896);
or U28624 (N_28624,N_25656,N_27462);
and U28625 (N_28625,N_26206,N_26161);
nand U28626 (N_28626,N_27270,N_27224);
or U28627 (N_28627,N_26891,N_25907);
xor U28628 (N_28628,N_26934,N_26130);
nor U28629 (N_28629,N_25568,N_25002);
or U28630 (N_28630,N_25231,N_26140);
nor U28631 (N_28631,N_25651,N_26363);
nor U28632 (N_28632,N_26411,N_26717);
xnor U28633 (N_28633,N_27258,N_26341);
nand U28634 (N_28634,N_26373,N_26212);
xor U28635 (N_28635,N_26573,N_27201);
nor U28636 (N_28636,N_25638,N_25899);
and U28637 (N_28637,N_25115,N_25965);
or U28638 (N_28638,N_25846,N_25672);
and U28639 (N_28639,N_25507,N_25468);
nor U28640 (N_28640,N_25747,N_27291);
nand U28641 (N_28641,N_26799,N_25483);
nand U28642 (N_28642,N_26070,N_25927);
or U28643 (N_28643,N_26265,N_26404);
nor U28644 (N_28644,N_25652,N_27202);
nor U28645 (N_28645,N_26051,N_27094);
nor U28646 (N_28646,N_27056,N_25301);
nor U28647 (N_28647,N_26667,N_27209);
and U28648 (N_28648,N_26992,N_26303);
xor U28649 (N_28649,N_27401,N_27393);
nor U28650 (N_28650,N_25695,N_27434);
nor U28651 (N_28651,N_25788,N_25268);
nor U28652 (N_28652,N_25513,N_25995);
nand U28653 (N_28653,N_26241,N_25745);
or U28654 (N_28654,N_25227,N_25334);
xnor U28655 (N_28655,N_25165,N_27442);
nor U28656 (N_28656,N_26632,N_25213);
and U28657 (N_28657,N_25675,N_25457);
nor U28658 (N_28658,N_26580,N_27039);
and U28659 (N_28659,N_25617,N_25514);
and U28660 (N_28660,N_26858,N_25598);
xor U28661 (N_28661,N_26180,N_26402);
nand U28662 (N_28662,N_27300,N_25394);
and U28663 (N_28663,N_26239,N_26238);
or U28664 (N_28664,N_25960,N_27149);
or U28665 (N_28665,N_26723,N_25401);
nand U28666 (N_28666,N_25929,N_26148);
xnor U28667 (N_28667,N_26842,N_25474);
nand U28668 (N_28668,N_25345,N_25646);
and U28669 (N_28669,N_25230,N_26374);
or U28670 (N_28670,N_26818,N_25976);
or U28671 (N_28671,N_25798,N_26970);
nand U28672 (N_28672,N_25849,N_26296);
nor U28673 (N_28673,N_26567,N_26270);
xnor U28674 (N_28674,N_25204,N_26652);
nor U28675 (N_28675,N_27166,N_26177);
or U28676 (N_28676,N_26706,N_27284);
xor U28677 (N_28677,N_27077,N_25179);
and U28678 (N_28678,N_26444,N_25797);
nor U28679 (N_28679,N_25327,N_25839);
nand U28680 (N_28680,N_27010,N_27455);
and U28681 (N_28681,N_25776,N_25528);
and U28682 (N_28682,N_25494,N_26691);
nand U28683 (N_28683,N_25039,N_27403);
and U28684 (N_28684,N_25871,N_25870);
nand U28685 (N_28685,N_26840,N_26894);
nor U28686 (N_28686,N_26823,N_26113);
nor U28687 (N_28687,N_26327,N_26200);
nor U28688 (N_28688,N_26259,N_27111);
or U28689 (N_28689,N_25260,N_27422);
xnor U28690 (N_28690,N_25910,N_27334);
nor U28691 (N_28691,N_25980,N_26400);
xor U28692 (N_28692,N_26779,N_26814);
nand U28693 (N_28693,N_27329,N_26892);
or U28694 (N_28694,N_25615,N_25618);
xor U28695 (N_28695,N_27453,N_25770);
nor U28696 (N_28696,N_26227,N_25416);
and U28697 (N_28697,N_26772,N_25052);
and U28698 (N_28698,N_26328,N_25674);
xnor U28699 (N_28699,N_27429,N_25589);
nand U28700 (N_28700,N_25271,N_26438);
nor U28701 (N_28701,N_27101,N_26871);
xnor U28702 (N_28702,N_25898,N_26983);
xnor U28703 (N_28703,N_27438,N_26284);
and U28704 (N_28704,N_25304,N_27030);
and U28705 (N_28705,N_25441,N_27385);
nor U28706 (N_28706,N_27048,N_25241);
nor U28707 (N_28707,N_26339,N_26309);
and U28708 (N_28708,N_26584,N_25607);
or U28709 (N_28709,N_26261,N_27144);
nor U28710 (N_28710,N_25707,N_26262);
nor U28711 (N_28711,N_26802,N_25353);
nand U28712 (N_28712,N_26119,N_25572);
xnor U28713 (N_28713,N_26247,N_26637);
nor U28714 (N_28714,N_26643,N_25463);
nor U28715 (N_28715,N_25628,N_25626);
xnor U28716 (N_28716,N_26703,N_27013);
nor U28717 (N_28717,N_25928,N_26868);
xnor U28718 (N_28718,N_26788,N_27471);
xor U28719 (N_28719,N_27411,N_26492);
and U28720 (N_28720,N_27172,N_26838);
nor U28721 (N_28721,N_25986,N_25860);
and U28722 (N_28722,N_26083,N_25655);
nand U28723 (N_28723,N_26395,N_26914);
and U28724 (N_28724,N_26500,N_27355);
xnor U28725 (N_28725,N_26014,N_26459);
nand U28726 (N_28726,N_26245,N_26674);
nor U28727 (N_28727,N_26211,N_25911);
nand U28728 (N_28728,N_25578,N_27207);
or U28729 (N_28729,N_25042,N_25603);
nand U28730 (N_28730,N_26264,N_27131);
xnor U28731 (N_28731,N_26009,N_27043);
xnor U28732 (N_28732,N_25442,N_27495);
and U28733 (N_28733,N_27079,N_25109);
nor U28734 (N_28734,N_27325,N_27259);
nand U28735 (N_28735,N_25048,N_26533);
nand U28736 (N_28736,N_26749,N_25352);
nor U28737 (N_28737,N_26997,N_25859);
or U28738 (N_28738,N_26535,N_25099);
xor U28739 (N_28739,N_26482,N_25393);
nor U28740 (N_28740,N_26016,N_26971);
nor U28741 (N_28741,N_26966,N_25523);
nor U28742 (N_28742,N_25449,N_26333);
or U28743 (N_28743,N_25153,N_27185);
nor U28744 (N_28744,N_26847,N_27368);
nand U28745 (N_28745,N_27059,N_26352);
xor U28746 (N_28746,N_26351,N_25487);
and U28747 (N_28747,N_25125,N_27381);
or U28748 (N_28748,N_25232,N_26676);
and U28749 (N_28749,N_26173,N_25374);
xnor U28750 (N_28750,N_26142,N_25589);
or U28751 (N_28751,N_26413,N_25318);
nand U28752 (N_28752,N_26267,N_25091);
nor U28753 (N_28753,N_25609,N_25558);
and U28754 (N_28754,N_27020,N_25010);
and U28755 (N_28755,N_27343,N_27007);
nor U28756 (N_28756,N_25057,N_26624);
nor U28757 (N_28757,N_25345,N_25711);
xnor U28758 (N_28758,N_26440,N_26655);
or U28759 (N_28759,N_25543,N_25301);
or U28760 (N_28760,N_25817,N_25831);
or U28761 (N_28761,N_25638,N_25841);
or U28762 (N_28762,N_26955,N_26127);
and U28763 (N_28763,N_27082,N_25421);
nor U28764 (N_28764,N_25612,N_26198);
xnor U28765 (N_28765,N_27039,N_27137);
nor U28766 (N_28766,N_27201,N_25854);
nand U28767 (N_28767,N_25045,N_26217);
xnor U28768 (N_28768,N_26049,N_25348);
xor U28769 (N_28769,N_26773,N_26174);
and U28770 (N_28770,N_25061,N_26760);
xor U28771 (N_28771,N_25293,N_25531);
and U28772 (N_28772,N_26240,N_26845);
and U28773 (N_28773,N_26109,N_26899);
or U28774 (N_28774,N_25289,N_25432);
xor U28775 (N_28775,N_27039,N_27325);
nand U28776 (N_28776,N_25165,N_26342);
nor U28777 (N_28777,N_27487,N_26159);
xnor U28778 (N_28778,N_26699,N_27063);
nor U28779 (N_28779,N_25775,N_26340);
or U28780 (N_28780,N_26909,N_26305);
and U28781 (N_28781,N_27451,N_27127);
nand U28782 (N_28782,N_26821,N_27131);
and U28783 (N_28783,N_25828,N_25949);
or U28784 (N_28784,N_27413,N_27371);
xor U28785 (N_28785,N_25014,N_26453);
xor U28786 (N_28786,N_27397,N_25565);
xor U28787 (N_28787,N_25289,N_27264);
or U28788 (N_28788,N_25897,N_27201);
or U28789 (N_28789,N_25311,N_25438);
and U28790 (N_28790,N_26993,N_25008);
xor U28791 (N_28791,N_26536,N_25545);
nor U28792 (N_28792,N_26973,N_26461);
and U28793 (N_28793,N_26929,N_25009);
or U28794 (N_28794,N_25123,N_26868);
xor U28795 (N_28795,N_26275,N_26760);
nand U28796 (N_28796,N_25704,N_25730);
and U28797 (N_28797,N_25818,N_27137);
or U28798 (N_28798,N_26482,N_25785);
and U28799 (N_28799,N_27186,N_25216);
xor U28800 (N_28800,N_25281,N_26769);
and U28801 (N_28801,N_25291,N_25686);
or U28802 (N_28802,N_25576,N_26209);
xnor U28803 (N_28803,N_27039,N_26254);
and U28804 (N_28804,N_26546,N_25071);
or U28805 (N_28805,N_25645,N_27478);
xor U28806 (N_28806,N_26383,N_27198);
nor U28807 (N_28807,N_25055,N_25978);
nor U28808 (N_28808,N_27147,N_25909);
xor U28809 (N_28809,N_27279,N_26601);
nor U28810 (N_28810,N_26486,N_26170);
nor U28811 (N_28811,N_25076,N_25872);
nand U28812 (N_28812,N_26256,N_26459);
xnor U28813 (N_28813,N_26501,N_27084);
xor U28814 (N_28814,N_26729,N_25705);
and U28815 (N_28815,N_26123,N_27092);
and U28816 (N_28816,N_26900,N_26587);
nand U28817 (N_28817,N_25998,N_26680);
nand U28818 (N_28818,N_26833,N_27112);
nand U28819 (N_28819,N_26805,N_26369);
nor U28820 (N_28820,N_25441,N_27117);
nor U28821 (N_28821,N_27258,N_27364);
nor U28822 (N_28822,N_25191,N_25890);
or U28823 (N_28823,N_25608,N_26225);
xnor U28824 (N_28824,N_27205,N_26318);
nor U28825 (N_28825,N_25926,N_26631);
or U28826 (N_28826,N_26942,N_25180);
and U28827 (N_28827,N_26092,N_25413);
or U28828 (N_28828,N_25662,N_26009);
or U28829 (N_28829,N_25635,N_27459);
and U28830 (N_28830,N_26229,N_25205);
nand U28831 (N_28831,N_25281,N_25098);
or U28832 (N_28832,N_25812,N_26344);
and U28833 (N_28833,N_27383,N_26976);
or U28834 (N_28834,N_25076,N_25293);
xor U28835 (N_28835,N_27455,N_26054);
nand U28836 (N_28836,N_26617,N_25050);
xnor U28837 (N_28837,N_26038,N_26703);
or U28838 (N_28838,N_25823,N_25579);
nor U28839 (N_28839,N_26007,N_26310);
xor U28840 (N_28840,N_27224,N_26358);
xor U28841 (N_28841,N_27034,N_25895);
nor U28842 (N_28842,N_25395,N_26976);
or U28843 (N_28843,N_26700,N_27415);
nor U28844 (N_28844,N_26203,N_25912);
nor U28845 (N_28845,N_25073,N_26044);
xnor U28846 (N_28846,N_26815,N_25585);
nor U28847 (N_28847,N_25986,N_27203);
xor U28848 (N_28848,N_25876,N_27173);
nand U28849 (N_28849,N_25771,N_26162);
xor U28850 (N_28850,N_26238,N_26583);
nor U28851 (N_28851,N_25595,N_26554);
nor U28852 (N_28852,N_27219,N_25279);
and U28853 (N_28853,N_27174,N_26945);
and U28854 (N_28854,N_25434,N_27112);
and U28855 (N_28855,N_27039,N_25024);
xnor U28856 (N_28856,N_26260,N_25289);
xnor U28857 (N_28857,N_26928,N_25502);
xnor U28858 (N_28858,N_25192,N_27011);
nand U28859 (N_28859,N_26871,N_26859);
nand U28860 (N_28860,N_25462,N_26073);
or U28861 (N_28861,N_25100,N_26899);
or U28862 (N_28862,N_27069,N_25729);
or U28863 (N_28863,N_26251,N_26690);
or U28864 (N_28864,N_25628,N_26632);
nor U28865 (N_28865,N_25811,N_27138);
or U28866 (N_28866,N_25562,N_25988);
nor U28867 (N_28867,N_25791,N_25547);
nand U28868 (N_28868,N_26141,N_25710);
nor U28869 (N_28869,N_26469,N_27057);
nor U28870 (N_28870,N_27142,N_26940);
nor U28871 (N_28871,N_26135,N_27291);
and U28872 (N_28872,N_26765,N_26076);
xnor U28873 (N_28873,N_26336,N_27018);
xor U28874 (N_28874,N_25712,N_25953);
nor U28875 (N_28875,N_26972,N_25866);
nand U28876 (N_28876,N_27233,N_26939);
nand U28877 (N_28877,N_26987,N_27323);
nand U28878 (N_28878,N_26757,N_25968);
nor U28879 (N_28879,N_25559,N_26504);
and U28880 (N_28880,N_25074,N_26257);
nand U28881 (N_28881,N_26206,N_27112);
xor U28882 (N_28882,N_27422,N_26909);
xor U28883 (N_28883,N_25893,N_25105);
xor U28884 (N_28884,N_25273,N_27112);
nor U28885 (N_28885,N_26048,N_26890);
or U28886 (N_28886,N_25541,N_27102);
nand U28887 (N_28887,N_25187,N_26774);
xor U28888 (N_28888,N_26747,N_26499);
xor U28889 (N_28889,N_26911,N_25783);
or U28890 (N_28890,N_26994,N_25977);
xnor U28891 (N_28891,N_26837,N_26465);
or U28892 (N_28892,N_25582,N_26314);
and U28893 (N_28893,N_25385,N_26952);
or U28894 (N_28894,N_26776,N_26821);
or U28895 (N_28895,N_25222,N_26420);
and U28896 (N_28896,N_25290,N_25796);
and U28897 (N_28897,N_25485,N_26246);
or U28898 (N_28898,N_25162,N_27398);
xnor U28899 (N_28899,N_25582,N_25615);
xor U28900 (N_28900,N_25234,N_25440);
nor U28901 (N_28901,N_25490,N_26056);
or U28902 (N_28902,N_25558,N_27461);
or U28903 (N_28903,N_26083,N_25113);
and U28904 (N_28904,N_25651,N_26472);
or U28905 (N_28905,N_27040,N_26951);
nand U28906 (N_28906,N_25039,N_25728);
and U28907 (N_28907,N_25127,N_25355);
xnor U28908 (N_28908,N_25324,N_25226);
nand U28909 (N_28909,N_25820,N_27069);
xnor U28910 (N_28910,N_26887,N_26377);
nand U28911 (N_28911,N_26037,N_25849);
and U28912 (N_28912,N_25724,N_26612);
nand U28913 (N_28913,N_25392,N_25905);
xnor U28914 (N_28914,N_25493,N_25192);
and U28915 (N_28915,N_27037,N_25841);
and U28916 (N_28916,N_25262,N_26640);
nand U28917 (N_28917,N_26244,N_25650);
or U28918 (N_28918,N_27337,N_27482);
xor U28919 (N_28919,N_27296,N_27198);
nand U28920 (N_28920,N_27354,N_25686);
or U28921 (N_28921,N_26448,N_25875);
nand U28922 (N_28922,N_26912,N_25543);
and U28923 (N_28923,N_26052,N_25382);
or U28924 (N_28924,N_25928,N_25196);
or U28925 (N_28925,N_26382,N_26325);
xnor U28926 (N_28926,N_25230,N_25998);
nor U28927 (N_28927,N_25924,N_26322);
xnor U28928 (N_28928,N_25647,N_25262);
and U28929 (N_28929,N_25261,N_25269);
xnor U28930 (N_28930,N_25326,N_25052);
nand U28931 (N_28931,N_26030,N_27367);
or U28932 (N_28932,N_25764,N_25762);
xnor U28933 (N_28933,N_25847,N_26642);
nor U28934 (N_28934,N_25594,N_26837);
or U28935 (N_28935,N_25473,N_25072);
nor U28936 (N_28936,N_25636,N_25174);
or U28937 (N_28937,N_26716,N_26901);
nor U28938 (N_28938,N_25337,N_26177);
nor U28939 (N_28939,N_27387,N_27216);
nand U28940 (N_28940,N_25843,N_25482);
or U28941 (N_28941,N_26141,N_25251);
or U28942 (N_28942,N_25875,N_25081);
xor U28943 (N_28943,N_26706,N_26153);
or U28944 (N_28944,N_26082,N_26796);
nand U28945 (N_28945,N_25845,N_25029);
nor U28946 (N_28946,N_26830,N_26681);
nand U28947 (N_28947,N_26763,N_26006);
nand U28948 (N_28948,N_26184,N_26451);
or U28949 (N_28949,N_26347,N_25281);
or U28950 (N_28950,N_26588,N_26203);
or U28951 (N_28951,N_25077,N_27004);
and U28952 (N_28952,N_25512,N_27099);
xor U28953 (N_28953,N_26620,N_25682);
or U28954 (N_28954,N_25809,N_27408);
xor U28955 (N_28955,N_26645,N_26738);
xnor U28956 (N_28956,N_26866,N_25429);
nand U28957 (N_28957,N_27400,N_26095);
xor U28958 (N_28958,N_27037,N_26701);
nand U28959 (N_28959,N_26175,N_26166);
or U28960 (N_28960,N_26417,N_26070);
nand U28961 (N_28961,N_27133,N_26028);
and U28962 (N_28962,N_25306,N_26990);
or U28963 (N_28963,N_26676,N_27409);
nor U28964 (N_28964,N_25682,N_26384);
nor U28965 (N_28965,N_27306,N_26864);
xor U28966 (N_28966,N_25820,N_27150);
and U28967 (N_28967,N_25188,N_27490);
nor U28968 (N_28968,N_25566,N_25414);
nor U28969 (N_28969,N_25767,N_26254);
and U28970 (N_28970,N_26981,N_26887);
xnor U28971 (N_28971,N_26607,N_26288);
nand U28972 (N_28972,N_26417,N_26439);
or U28973 (N_28973,N_25130,N_27151);
and U28974 (N_28974,N_25155,N_26695);
nor U28975 (N_28975,N_26474,N_25048);
xnor U28976 (N_28976,N_26853,N_26725);
xor U28977 (N_28977,N_26394,N_26752);
xor U28978 (N_28978,N_25923,N_25592);
nand U28979 (N_28979,N_25270,N_26994);
nand U28980 (N_28980,N_25900,N_25512);
or U28981 (N_28981,N_25634,N_25564);
nand U28982 (N_28982,N_26587,N_26015);
nor U28983 (N_28983,N_25986,N_26403);
xor U28984 (N_28984,N_27440,N_25503);
nand U28985 (N_28985,N_26835,N_25636);
or U28986 (N_28986,N_26677,N_25520);
and U28987 (N_28987,N_27166,N_26703);
or U28988 (N_28988,N_25323,N_27297);
nor U28989 (N_28989,N_27126,N_25468);
nand U28990 (N_28990,N_26083,N_26384);
nand U28991 (N_28991,N_27460,N_26733);
nor U28992 (N_28992,N_27064,N_26632);
and U28993 (N_28993,N_27007,N_25865);
nor U28994 (N_28994,N_26342,N_25161);
and U28995 (N_28995,N_25787,N_25647);
xor U28996 (N_28996,N_25375,N_26305);
nor U28997 (N_28997,N_26932,N_26204);
xor U28998 (N_28998,N_26202,N_26473);
and U28999 (N_28999,N_25935,N_25952);
or U29000 (N_29000,N_27431,N_26167);
and U29001 (N_29001,N_26246,N_27456);
nand U29002 (N_29002,N_26826,N_26339);
and U29003 (N_29003,N_25414,N_25477);
nand U29004 (N_29004,N_25865,N_25003);
nor U29005 (N_29005,N_25440,N_25241);
xor U29006 (N_29006,N_26223,N_25098);
xnor U29007 (N_29007,N_25690,N_25556);
or U29008 (N_29008,N_26064,N_26107);
or U29009 (N_29009,N_27196,N_25796);
nand U29010 (N_29010,N_26233,N_26610);
nor U29011 (N_29011,N_26975,N_25660);
nor U29012 (N_29012,N_26012,N_26550);
or U29013 (N_29013,N_27240,N_25363);
nor U29014 (N_29014,N_27030,N_25484);
nor U29015 (N_29015,N_25158,N_26334);
or U29016 (N_29016,N_27091,N_27318);
nor U29017 (N_29017,N_25750,N_26582);
nor U29018 (N_29018,N_25588,N_25901);
and U29019 (N_29019,N_25197,N_25136);
nand U29020 (N_29020,N_25966,N_25108);
nand U29021 (N_29021,N_25286,N_25644);
or U29022 (N_29022,N_25205,N_27320);
nand U29023 (N_29023,N_26091,N_26948);
or U29024 (N_29024,N_26332,N_25793);
and U29025 (N_29025,N_27085,N_26099);
or U29026 (N_29026,N_27445,N_26316);
or U29027 (N_29027,N_25589,N_26988);
nand U29028 (N_29028,N_25667,N_25156);
and U29029 (N_29029,N_25877,N_26686);
and U29030 (N_29030,N_26941,N_26741);
nand U29031 (N_29031,N_25039,N_25356);
xor U29032 (N_29032,N_27495,N_27429);
or U29033 (N_29033,N_26820,N_25354);
nor U29034 (N_29034,N_25534,N_27161);
xor U29035 (N_29035,N_25388,N_26314);
nor U29036 (N_29036,N_26987,N_26378);
or U29037 (N_29037,N_25869,N_27248);
xor U29038 (N_29038,N_26863,N_25683);
xor U29039 (N_29039,N_25114,N_25895);
nor U29040 (N_29040,N_25211,N_26467);
and U29041 (N_29041,N_27260,N_25592);
xor U29042 (N_29042,N_26509,N_26300);
nand U29043 (N_29043,N_25620,N_26618);
or U29044 (N_29044,N_25439,N_26897);
xor U29045 (N_29045,N_25298,N_25300);
nand U29046 (N_29046,N_26408,N_25082);
nor U29047 (N_29047,N_26314,N_25593);
or U29048 (N_29048,N_27084,N_25231);
nor U29049 (N_29049,N_25848,N_25584);
xor U29050 (N_29050,N_25207,N_26917);
nor U29051 (N_29051,N_26650,N_26495);
and U29052 (N_29052,N_26076,N_26339);
nand U29053 (N_29053,N_27329,N_26433);
or U29054 (N_29054,N_25272,N_27153);
nor U29055 (N_29055,N_25054,N_27076);
and U29056 (N_29056,N_26189,N_25659);
nand U29057 (N_29057,N_26497,N_26684);
or U29058 (N_29058,N_25242,N_27402);
xnor U29059 (N_29059,N_26715,N_25527);
nor U29060 (N_29060,N_27004,N_26687);
nor U29061 (N_29061,N_25906,N_26586);
nor U29062 (N_29062,N_25977,N_25887);
nand U29063 (N_29063,N_26228,N_27080);
nor U29064 (N_29064,N_26883,N_26454);
xor U29065 (N_29065,N_25704,N_26035);
nand U29066 (N_29066,N_27460,N_27070);
xnor U29067 (N_29067,N_25371,N_25514);
and U29068 (N_29068,N_26230,N_25448);
nand U29069 (N_29069,N_26395,N_25129);
nand U29070 (N_29070,N_26705,N_25033);
nor U29071 (N_29071,N_25974,N_25895);
and U29072 (N_29072,N_26333,N_25140);
nand U29073 (N_29073,N_25133,N_25766);
nor U29074 (N_29074,N_27057,N_26834);
and U29075 (N_29075,N_25889,N_26666);
xnor U29076 (N_29076,N_26468,N_25391);
and U29077 (N_29077,N_25404,N_25192);
or U29078 (N_29078,N_25521,N_26772);
nor U29079 (N_29079,N_25576,N_26126);
nand U29080 (N_29080,N_26166,N_27385);
and U29081 (N_29081,N_26509,N_25034);
and U29082 (N_29082,N_26213,N_25991);
nor U29083 (N_29083,N_25513,N_25556);
xor U29084 (N_29084,N_26078,N_25118);
nor U29085 (N_29085,N_25789,N_25301);
and U29086 (N_29086,N_26840,N_25958);
or U29087 (N_29087,N_25749,N_25643);
nor U29088 (N_29088,N_26142,N_27213);
xor U29089 (N_29089,N_25553,N_25556);
nand U29090 (N_29090,N_25317,N_27278);
and U29091 (N_29091,N_25238,N_27285);
or U29092 (N_29092,N_26450,N_26396);
and U29093 (N_29093,N_25020,N_26703);
or U29094 (N_29094,N_26020,N_25254);
xnor U29095 (N_29095,N_25347,N_26928);
nor U29096 (N_29096,N_26672,N_25649);
nand U29097 (N_29097,N_26023,N_25275);
and U29098 (N_29098,N_25864,N_25928);
nand U29099 (N_29099,N_27020,N_26425);
and U29100 (N_29100,N_25905,N_25601);
or U29101 (N_29101,N_27048,N_27399);
nor U29102 (N_29102,N_26728,N_25185);
xor U29103 (N_29103,N_25779,N_26519);
nand U29104 (N_29104,N_25185,N_25879);
or U29105 (N_29105,N_25998,N_26324);
nor U29106 (N_29106,N_26760,N_27359);
and U29107 (N_29107,N_25431,N_26374);
nor U29108 (N_29108,N_26547,N_26020);
nand U29109 (N_29109,N_25841,N_26625);
or U29110 (N_29110,N_26787,N_25489);
xor U29111 (N_29111,N_25492,N_25111);
and U29112 (N_29112,N_25812,N_25192);
xnor U29113 (N_29113,N_25733,N_27318);
and U29114 (N_29114,N_25895,N_27431);
or U29115 (N_29115,N_27403,N_25323);
nand U29116 (N_29116,N_26387,N_27124);
nand U29117 (N_29117,N_25678,N_27192);
or U29118 (N_29118,N_27064,N_25813);
or U29119 (N_29119,N_26301,N_25600);
xnor U29120 (N_29120,N_25626,N_27487);
nor U29121 (N_29121,N_26922,N_26683);
nand U29122 (N_29122,N_26766,N_25741);
nor U29123 (N_29123,N_26185,N_27233);
nand U29124 (N_29124,N_25692,N_27133);
and U29125 (N_29125,N_26504,N_25390);
or U29126 (N_29126,N_26773,N_27409);
and U29127 (N_29127,N_27411,N_25113);
nor U29128 (N_29128,N_25968,N_27063);
nor U29129 (N_29129,N_27024,N_26735);
xnor U29130 (N_29130,N_25253,N_27305);
nand U29131 (N_29131,N_26086,N_26863);
nand U29132 (N_29132,N_25277,N_27357);
nand U29133 (N_29133,N_26054,N_25799);
xor U29134 (N_29134,N_27063,N_25378);
xor U29135 (N_29135,N_27363,N_25944);
nand U29136 (N_29136,N_26959,N_26935);
nand U29137 (N_29137,N_26890,N_25180);
and U29138 (N_29138,N_25735,N_26437);
nor U29139 (N_29139,N_25978,N_25561);
or U29140 (N_29140,N_25347,N_26650);
and U29141 (N_29141,N_25108,N_27144);
and U29142 (N_29142,N_27068,N_26102);
xnor U29143 (N_29143,N_26914,N_27364);
xor U29144 (N_29144,N_25142,N_25527);
xnor U29145 (N_29145,N_25307,N_25604);
and U29146 (N_29146,N_27253,N_26938);
xnor U29147 (N_29147,N_25084,N_26319);
and U29148 (N_29148,N_25063,N_26874);
nor U29149 (N_29149,N_27318,N_25960);
nand U29150 (N_29150,N_25462,N_25648);
and U29151 (N_29151,N_25287,N_26037);
and U29152 (N_29152,N_25477,N_26479);
or U29153 (N_29153,N_26453,N_26664);
or U29154 (N_29154,N_27349,N_25607);
xnor U29155 (N_29155,N_27444,N_26500);
nor U29156 (N_29156,N_26197,N_25525);
or U29157 (N_29157,N_26907,N_26865);
nor U29158 (N_29158,N_27344,N_26680);
xor U29159 (N_29159,N_27057,N_26499);
nor U29160 (N_29160,N_26977,N_26124);
and U29161 (N_29161,N_25972,N_25389);
nor U29162 (N_29162,N_27348,N_25782);
nor U29163 (N_29163,N_25372,N_26832);
or U29164 (N_29164,N_25909,N_26134);
nand U29165 (N_29165,N_25923,N_27497);
nand U29166 (N_29166,N_26170,N_26306);
nor U29167 (N_29167,N_26324,N_25329);
nor U29168 (N_29168,N_25419,N_25929);
and U29169 (N_29169,N_27385,N_27086);
nand U29170 (N_29170,N_26688,N_26799);
nand U29171 (N_29171,N_26779,N_25292);
nand U29172 (N_29172,N_25735,N_26794);
and U29173 (N_29173,N_26585,N_26714);
or U29174 (N_29174,N_26320,N_25289);
nand U29175 (N_29175,N_27160,N_27361);
nand U29176 (N_29176,N_26333,N_27007);
nand U29177 (N_29177,N_26252,N_25165);
nand U29178 (N_29178,N_26415,N_26447);
xor U29179 (N_29179,N_26574,N_26337);
xnor U29180 (N_29180,N_25675,N_26545);
xor U29181 (N_29181,N_26603,N_27290);
or U29182 (N_29182,N_25205,N_27066);
nand U29183 (N_29183,N_25247,N_27306);
or U29184 (N_29184,N_26858,N_25026);
nor U29185 (N_29185,N_25579,N_25401);
nor U29186 (N_29186,N_26127,N_26136);
and U29187 (N_29187,N_27121,N_27306);
nor U29188 (N_29188,N_26623,N_26706);
nand U29189 (N_29189,N_25199,N_25979);
or U29190 (N_29190,N_25633,N_26876);
and U29191 (N_29191,N_26249,N_25232);
and U29192 (N_29192,N_25029,N_27208);
nand U29193 (N_29193,N_26069,N_27408);
or U29194 (N_29194,N_26390,N_26226);
nand U29195 (N_29195,N_27334,N_26887);
nor U29196 (N_29196,N_26714,N_27203);
or U29197 (N_29197,N_26414,N_26226);
nor U29198 (N_29198,N_25800,N_25365);
or U29199 (N_29199,N_26564,N_25162);
and U29200 (N_29200,N_25033,N_27136);
nand U29201 (N_29201,N_25846,N_27235);
nand U29202 (N_29202,N_27417,N_26299);
and U29203 (N_29203,N_26400,N_26860);
xor U29204 (N_29204,N_25806,N_27357);
or U29205 (N_29205,N_27254,N_25705);
or U29206 (N_29206,N_27346,N_25351);
nor U29207 (N_29207,N_27049,N_25877);
nor U29208 (N_29208,N_27403,N_26190);
or U29209 (N_29209,N_27036,N_25335);
nor U29210 (N_29210,N_26462,N_25781);
nor U29211 (N_29211,N_25853,N_26415);
nand U29212 (N_29212,N_26978,N_25172);
or U29213 (N_29213,N_25321,N_25295);
xor U29214 (N_29214,N_25720,N_25850);
or U29215 (N_29215,N_26484,N_25221);
or U29216 (N_29216,N_25088,N_26465);
and U29217 (N_29217,N_27226,N_25263);
or U29218 (N_29218,N_27017,N_25727);
nor U29219 (N_29219,N_25358,N_27427);
xnor U29220 (N_29220,N_26455,N_25811);
or U29221 (N_29221,N_25963,N_26781);
nand U29222 (N_29222,N_27297,N_25842);
or U29223 (N_29223,N_26817,N_27235);
nor U29224 (N_29224,N_25872,N_27137);
xor U29225 (N_29225,N_26357,N_25505);
and U29226 (N_29226,N_27163,N_26457);
xnor U29227 (N_29227,N_26321,N_27378);
xor U29228 (N_29228,N_25644,N_25745);
and U29229 (N_29229,N_26465,N_26200);
nor U29230 (N_29230,N_25228,N_26609);
xnor U29231 (N_29231,N_25302,N_25131);
or U29232 (N_29232,N_26566,N_25146);
xnor U29233 (N_29233,N_25088,N_26410);
xor U29234 (N_29234,N_26499,N_25000);
nand U29235 (N_29235,N_25317,N_26647);
nand U29236 (N_29236,N_26197,N_25401);
xor U29237 (N_29237,N_26499,N_26346);
or U29238 (N_29238,N_25132,N_26543);
nor U29239 (N_29239,N_26851,N_26916);
or U29240 (N_29240,N_25254,N_25374);
nor U29241 (N_29241,N_27109,N_25177);
xor U29242 (N_29242,N_25897,N_26637);
xnor U29243 (N_29243,N_25890,N_26859);
nand U29244 (N_29244,N_27039,N_25686);
or U29245 (N_29245,N_25793,N_26595);
and U29246 (N_29246,N_26171,N_26848);
nor U29247 (N_29247,N_26701,N_26174);
or U29248 (N_29248,N_25876,N_26031);
and U29249 (N_29249,N_25788,N_26795);
xnor U29250 (N_29250,N_25691,N_27427);
and U29251 (N_29251,N_26913,N_27047);
nor U29252 (N_29252,N_27166,N_26111);
nor U29253 (N_29253,N_26334,N_26659);
or U29254 (N_29254,N_27266,N_25400);
nor U29255 (N_29255,N_27458,N_25119);
nor U29256 (N_29256,N_26300,N_27366);
or U29257 (N_29257,N_25785,N_26526);
or U29258 (N_29258,N_25371,N_26275);
or U29259 (N_29259,N_26805,N_25318);
xor U29260 (N_29260,N_25703,N_27422);
or U29261 (N_29261,N_25296,N_26779);
and U29262 (N_29262,N_25958,N_25746);
nor U29263 (N_29263,N_25896,N_25877);
nor U29264 (N_29264,N_27496,N_26264);
or U29265 (N_29265,N_26099,N_26796);
or U29266 (N_29266,N_25997,N_25820);
nor U29267 (N_29267,N_25057,N_26435);
nand U29268 (N_29268,N_27289,N_26074);
or U29269 (N_29269,N_25161,N_26508);
nor U29270 (N_29270,N_25003,N_25529);
xnor U29271 (N_29271,N_27378,N_25947);
and U29272 (N_29272,N_27273,N_25679);
nor U29273 (N_29273,N_25050,N_25929);
nor U29274 (N_29274,N_26679,N_25617);
xor U29275 (N_29275,N_27206,N_27233);
or U29276 (N_29276,N_26859,N_25491);
nand U29277 (N_29277,N_26935,N_25688);
nor U29278 (N_29278,N_27002,N_27239);
nor U29279 (N_29279,N_26217,N_26437);
and U29280 (N_29280,N_27301,N_26602);
nand U29281 (N_29281,N_27324,N_25963);
xor U29282 (N_29282,N_25828,N_25048);
or U29283 (N_29283,N_26673,N_26036);
nand U29284 (N_29284,N_27144,N_25770);
nor U29285 (N_29285,N_25810,N_25449);
nand U29286 (N_29286,N_26512,N_27339);
xor U29287 (N_29287,N_25929,N_26042);
or U29288 (N_29288,N_27336,N_25239);
and U29289 (N_29289,N_26703,N_25091);
nor U29290 (N_29290,N_26718,N_27157);
xnor U29291 (N_29291,N_25088,N_26453);
nor U29292 (N_29292,N_27006,N_25709);
or U29293 (N_29293,N_27374,N_26541);
or U29294 (N_29294,N_26015,N_27272);
and U29295 (N_29295,N_25878,N_26342);
nand U29296 (N_29296,N_26165,N_25806);
nor U29297 (N_29297,N_25079,N_27398);
or U29298 (N_29298,N_26019,N_26347);
and U29299 (N_29299,N_25388,N_25609);
and U29300 (N_29300,N_27152,N_25050);
xnor U29301 (N_29301,N_26099,N_26121);
xor U29302 (N_29302,N_25029,N_26127);
and U29303 (N_29303,N_25414,N_26400);
or U29304 (N_29304,N_26195,N_26818);
nor U29305 (N_29305,N_27477,N_26802);
nor U29306 (N_29306,N_25330,N_27325);
nand U29307 (N_29307,N_27110,N_27212);
nor U29308 (N_29308,N_26504,N_26712);
nor U29309 (N_29309,N_27027,N_26652);
xor U29310 (N_29310,N_25700,N_26267);
nand U29311 (N_29311,N_27003,N_26953);
and U29312 (N_29312,N_27304,N_26177);
xor U29313 (N_29313,N_26607,N_26192);
and U29314 (N_29314,N_25679,N_27186);
xor U29315 (N_29315,N_26967,N_25449);
xor U29316 (N_29316,N_25226,N_27436);
or U29317 (N_29317,N_26126,N_27127);
nor U29318 (N_29318,N_25823,N_26920);
xnor U29319 (N_29319,N_26798,N_25003);
or U29320 (N_29320,N_25105,N_25156);
nor U29321 (N_29321,N_26911,N_26155);
or U29322 (N_29322,N_25450,N_27180);
and U29323 (N_29323,N_26049,N_25188);
xnor U29324 (N_29324,N_25774,N_25883);
and U29325 (N_29325,N_26355,N_25164);
xnor U29326 (N_29326,N_25188,N_25383);
and U29327 (N_29327,N_26236,N_26356);
nor U29328 (N_29328,N_25488,N_26332);
nor U29329 (N_29329,N_26413,N_25374);
nand U29330 (N_29330,N_27075,N_27164);
or U29331 (N_29331,N_26337,N_25908);
nor U29332 (N_29332,N_26298,N_26872);
or U29333 (N_29333,N_25144,N_26266);
or U29334 (N_29334,N_25247,N_26313);
and U29335 (N_29335,N_27365,N_26350);
and U29336 (N_29336,N_26851,N_27499);
nor U29337 (N_29337,N_25913,N_25900);
nand U29338 (N_29338,N_25099,N_27382);
nor U29339 (N_29339,N_27412,N_27137);
or U29340 (N_29340,N_26034,N_25619);
nor U29341 (N_29341,N_25013,N_27065);
and U29342 (N_29342,N_25663,N_27429);
or U29343 (N_29343,N_27113,N_25161);
and U29344 (N_29344,N_26805,N_26054);
nand U29345 (N_29345,N_27390,N_25018);
and U29346 (N_29346,N_26869,N_26692);
xor U29347 (N_29347,N_27148,N_26330);
and U29348 (N_29348,N_25883,N_27055);
and U29349 (N_29349,N_25786,N_26723);
nand U29350 (N_29350,N_25635,N_25512);
xor U29351 (N_29351,N_26056,N_26543);
xnor U29352 (N_29352,N_27403,N_26220);
nand U29353 (N_29353,N_25598,N_27423);
nand U29354 (N_29354,N_26715,N_26915);
or U29355 (N_29355,N_26204,N_25114);
nand U29356 (N_29356,N_25969,N_26010);
or U29357 (N_29357,N_25998,N_26371);
xnor U29358 (N_29358,N_26644,N_25395);
xnor U29359 (N_29359,N_27198,N_27106);
or U29360 (N_29360,N_27481,N_25890);
xor U29361 (N_29361,N_25953,N_25899);
and U29362 (N_29362,N_26645,N_26599);
or U29363 (N_29363,N_27499,N_25503);
nor U29364 (N_29364,N_26887,N_25501);
nor U29365 (N_29365,N_26470,N_25615);
xnor U29366 (N_29366,N_25085,N_25534);
nor U29367 (N_29367,N_25632,N_25097);
or U29368 (N_29368,N_25143,N_26825);
and U29369 (N_29369,N_25096,N_25905);
nand U29370 (N_29370,N_25227,N_25762);
or U29371 (N_29371,N_26214,N_26970);
or U29372 (N_29372,N_27059,N_25061);
and U29373 (N_29373,N_26825,N_27292);
nor U29374 (N_29374,N_25341,N_25754);
nand U29375 (N_29375,N_25952,N_26843);
xor U29376 (N_29376,N_26322,N_27225);
xor U29377 (N_29377,N_27253,N_27348);
xor U29378 (N_29378,N_25147,N_25139);
nand U29379 (N_29379,N_25401,N_26170);
or U29380 (N_29380,N_26376,N_26539);
nor U29381 (N_29381,N_26574,N_26094);
xnor U29382 (N_29382,N_27320,N_26621);
xor U29383 (N_29383,N_27070,N_25736);
and U29384 (N_29384,N_25015,N_25102);
or U29385 (N_29385,N_26055,N_26046);
nand U29386 (N_29386,N_25227,N_25397);
or U29387 (N_29387,N_26453,N_27439);
nor U29388 (N_29388,N_27492,N_26765);
nand U29389 (N_29389,N_26552,N_26322);
and U29390 (N_29390,N_25023,N_26973);
xor U29391 (N_29391,N_26052,N_26307);
xnor U29392 (N_29392,N_26999,N_26039);
nand U29393 (N_29393,N_27374,N_25189);
and U29394 (N_29394,N_27295,N_27154);
nor U29395 (N_29395,N_25801,N_25072);
nor U29396 (N_29396,N_27176,N_27394);
or U29397 (N_29397,N_26992,N_26579);
nor U29398 (N_29398,N_25154,N_25368);
xor U29399 (N_29399,N_26925,N_25502);
or U29400 (N_29400,N_26173,N_25335);
nand U29401 (N_29401,N_26434,N_26286);
xor U29402 (N_29402,N_25287,N_27257);
and U29403 (N_29403,N_26645,N_26708);
nand U29404 (N_29404,N_27489,N_27212);
and U29405 (N_29405,N_27276,N_27207);
xor U29406 (N_29406,N_26523,N_25597);
xor U29407 (N_29407,N_26625,N_26719);
nor U29408 (N_29408,N_26203,N_27168);
and U29409 (N_29409,N_25187,N_26647);
nand U29410 (N_29410,N_27193,N_25358);
and U29411 (N_29411,N_26108,N_26912);
and U29412 (N_29412,N_25433,N_27030);
nand U29413 (N_29413,N_25728,N_26296);
and U29414 (N_29414,N_26967,N_26469);
nand U29415 (N_29415,N_25380,N_25425);
nor U29416 (N_29416,N_27438,N_25346);
or U29417 (N_29417,N_25351,N_25508);
nand U29418 (N_29418,N_26201,N_26098);
nor U29419 (N_29419,N_26278,N_26780);
xnor U29420 (N_29420,N_25346,N_25741);
xnor U29421 (N_29421,N_26469,N_25432);
or U29422 (N_29422,N_27075,N_25392);
xnor U29423 (N_29423,N_27153,N_25145);
xor U29424 (N_29424,N_26087,N_27138);
and U29425 (N_29425,N_25194,N_26746);
and U29426 (N_29426,N_26805,N_26084);
and U29427 (N_29427,N_26119,N_27336);
and U29428 (N_29428,N_26755,N_26156);
nand U29429 (N_29429,N_25771,N_25906);
xor U29430 (N_29430,N_25297,N_26336);
xor U29431 (N_29431,N_27021,N_26540);
xor U29432 (N_29432,N_26002,N_25825);
xnor U29433 (N_29433,N_25960,N_27416);
nor U29434 (N_29434,N_25417,N_27451);
and U29435 (N_29435,N_26465,N_27084);
or U29436 (N_29436,N_25406,N_26279);
nand U29437 (N_29437,N_27379,N_25856);
nand U29438 (N_29438,N_27342,N_25959);
xor U29439 (N_29439,N_27406,N_26707);
nor U29440 (N_29440,N_27493,N_26830);
xnor U29441 (N_29441,N_26448,N_27036);
nor U29442 (N_29442,N_25039,N_25830);
nor U29443 (N_29443,N_27164,N_26235);
nand U29444 (N_29444,N_26071,N_26867);
and U29445 (N_29445,N_25041,N_25472);
and U29446 (N_29446,N_26772,N_26171);
xor U29447 (N_29447,N_25348,N_25800);
and U29448 (N_29448,N_26552,N_27073);
xor U29449 (N_29449,N_27297,N_25796);
xor U29450 (N_29450,N_26152,N_26144);
nand U29451 (N_29451,N_25009,N_26870);
nand U29452 (N_29452,N_25952,N_25196);
nor U29453 (N_29453,N_26034,N_26664);
xnor U29454 (N_29454,N_26057,N_26814);
and U29455 (N_29455,N_26622,N_25680);
nand U29456 (N_29456,N_27164,N_25687);
nand U29457 (N_29457,N_26814,N_25758);
xor U29458 (N_29458,N_25590,N_26589);
and U29459 (N_29459,N_26766,N_25892);
or U29460 (N_29460,N_25755,N_25187);
and U29461 (N_29461,N_26854,N_25314);
xnor U29462 (N_29462,N_25861,N_27428);
nand U29463 (N_29463,N_26772,N_25896);
nand U29464 (N_29464,N_25938,N_27094);
or U29465 (N_29465,N_26492,N_25303);
and U29466 (N_29466,N_25355,N_26846);
xor U29467 (N_29467,N_25094,N_25150);
nor U29468 (N_29468,N_26937,N_26474);
xnor U29469 (N_29469,N_25395,N_25000);
nor U29470 (N_29470,N_26247,N_26831);
nor U29471 (N_29471,N_26014,N_27335);
nor U29472 (N_29472,N_25401,N_26793);
or U29473 (N_29473,N_27338,N_25483);
and U29474 (N_29474,N_26466,N_25868);
or U29475 (N_29475,N_26712,N_26562);
and U29476 (N_29476,N_26694,N_26658);
or U29477 (N_29477,N_26504,N_26672);
nor U29478 (N_29478,N_26635,N_25693);
nor U29479 (N_29479,N_25479,N_25937);
nand U29480 (N_29480,N_25651,N_27076);
nand U29481 (N_29481,N_26699,N_26979);
and U29482 (N_29482,N_26206,N_25919);
or U29483 (N_29483,N_25145,N_25820);
xor U29484 (N_29484,N_25068,N_26621);
xor U29485 (N_29485,N_25260,N_27250);
xor U29486 (N_29486,N_25664,N_27235);
and U29487 (N_29487,N_25157,N_27410);
nor U29488 (N_29488,N_26773,N_25661);
or U29489 (N_29489,N_25002,N_25299);
xor U29490 (N_29490,N_25302,N_25650);
and U29491 (N_29491,N_25228,N_25411);
and U29492 (N_29492,N_26751,N_27086);
xnor U29493 (N_29493,N_25228,N_26230);
nand U29494 (N_29494,N_27116,N_25042);
or U29495 (N_29495,N_25191,N_27031);
nor U29496 (N_29496,N_26390,N_26825);
nand U29497 (N_29497,N_27091,N_27006);
and U29498 (N_29498,N_26882,N_26015);
nand U29499 (N_29499,N_26954,N_26276);
and U29500 (N_29500,N_27267,N_27332);
and U29501 (N_29501,N_26188,N_27433);
nand U29502 (N_29502,N_25143,N_25986);
or U29503 (N_29503,N_25523,N_25088);
nand U29504 (N_29504,N_27070,N_26838);
xor U29505 (N_29505,N_26568,N_26675);
or U29506 (N_29506,N_26006,N_26155);
nor U29507 (N_29507,N_27426,N_26725);
or U29508 (N_29508,N_27441,N_27033);
and U29509 (N_29509,N_26166,N_25587);
nor U29510 (N_29510,N_26926,N_25758);
xnor U29511 (N_29511,N_25048,N_25986);
and U29512 (N_29512,N_25700,N_26206);
nand U29513 (N_29513,N_26026,N_27113);
nand U29514 (N_29514,N_27268,N_26271);
nor U29515 (N_29515,N_25359,N_26380);
or U29516 (N_29516,N_26445,N_25800);
xnor U29517 (N_29517,N_25928,N_27047);
or U29518 (N_29518,N_26611,N_25877);
nor U29519 (N_29519,N_25739,N_25487);
or U29520 (N_29520,N_27155,N_26101);
xor U29521 (N_29521,N_26828,N_26655);
xor U29522 (N_29522,N_26695,N_25567);
xor U29523 (N_29523,N_26076,N_27402);
nor U29524 (N_29524,N_26990,N_26432);
nor U29525 (N_29525,N_25897,N_26727);
xor U29526 (N_29526,N_26898,N_25034);
nand U29527 (N_29527,N_26549,N_26428);
nand U29528 (N_29528,N_25531,N_25315);
and U29529 (N_29529,N_26893,N_25689);
xnor U29530 (N_29530,N_25254,N_27116);
nand U29531 (N_29531,N_26633,N_26669);
and U29532 (N_29532,N_25764,N_25775);
or U29533 (N_29533,N_26022,N_26757);
xor U29534 (N_29534,N_25187,N_25210);
nand U29535 (N_29535,N_26062,N_26501);
nor U29536 (N_29536,N_27237,N_25761);
or U29537 (N_29537,N_25331,N_26686);
nor U29538 (N_29538,N_25683,N_25558);
nand U29539 (N_29539,N_25264,N_25291);
xor U29540 (N_29540,N_25741,N_26367);
xnor U29541 (N_29541,N_27010,N_26833);
xor U29542 (N_29542,N_25360,N_26616);
or U29543 (N_29543,N_25422,N_26861);
or U29544 (N_29544,N_26614,N_25218);
or U29545 (N_29545,N_26105,N_26890);
and U29546 (N_29546,N_26222,N_26096);
or U29547 (N_29547,N_26022,N_27051);
xor U29548 (N_29548,N_25659,N_27418);
nor U29549 (N_29549,N_27253,N_25954);
xnor U29550 (N_29550,N_27225,N_25780);
xnor U29551 (N_29551,N_27041,N_26664);
nor U29552 (N_29552,N_25703,N_25472);
and U29553 (N_29553,N_25280,N_26504);
and U29554 (N_29554,N_25002,N_27207);
xnor U29555 (N_29555,N_25449,N_26761);
nor U29556 (N_29556,N_25722,N_26975);
nor U29557 (N_29557,N_26472,N_26046);
xnor U29558 (N_29558,N_27474,N_26665);
or U29559 (N_29559,N_25145,N_26969);
nand U29560 (N_29560,N_26658,N_27329);
nand U29561 (N_29561,N_25950,N_26677);
xnor U29562 (N_29562,N_27389,N_25839);
or U29563 (N_29563,N_26419,N_27233);
nand U29564 (N_29564,N_27270,N_26822);
xor U29565 (N_29565,N_26999,N_26051);
nand U29566 (N_29566,N_25783,N_26765);
xnor U29567 (N_29567,N_25314,N_26252);
and U29568 (N_29568,N_26924,N_26416);
and U29569 (N_29569,N_25208,N_25937);
nand U29570 (N_29570,N_26359,N_26515);
xnor U29571 (N_29571,N_25721,N_25245);
or U29572 (N_29572,N_25916,N_26326);
or U29573 (N_29573,N_25649,N_26386);
xor U29574 (N_29574,N_25151,N_26646);
nand U29575 (N_29575,N_27148,N_25219);
xor U29576 (N_29576,N_25262,N_27427);
nor U29577 (N_29577,N_26946,N_25381);
nor U29578 (N_29578,N_26109,N_27490);
or U29579 (N_29579,N_25402,N_25039);
nand U29580 (N_29580,N_26150,N_26945);
xor U29581 (N_29581,N_26665,N_25200);
or U29582 (N_29582,N_25225,N_27045);
xor U29583 (N_29583,N_25697,N_25957);
or U29584 (N_29584,N_25526,N_27473);
xnor U29585 (N_29585,N_26785,N_25466);
nor U29586 (N_29586,N_25027,N_25225);
nand U29587 (N_29587,N_27407,N_27433);
nand U29588 (N_29588,N_25814,N_25240);
and U29589 (N_29589,N_26838,N_26832);
and U29590 (N_29590,N_26541,N_27007);
xnor U29591 (N_29591,N_27110,N_27440);
nand U29592 (N_29592,N_26397,N_26624);
or U29593 (N_29593,N_27357,N_25739);
xor U29594 (N_29594,N_25448,N_26482);
xor U29595 (N_29595,N_26859,N_27330);
nor U29596 (N_29596,N_25951,N_26546);
xor U29597 (N_29597,N_25081,N_25621);
and U29598 (N_29598,N_25310,N_27114);
or U29599 (N_29599,N_26163,N_25091);
nor U29600 (N_29600,N_25553,N_25496);
xor U29601 (N_29601,N_25698,N_26721);
xor U29602 (N_29602,N_25605,N_26251);
xnor U29603 (N_29603,N_25492,N_25087);
nor U29604 (N_29604,N_27464,N_25190);
xor U29605 (N_29605,N_27107,N_26994);
and U29606 (N_29606,N_26512,N_25117);
nand U29607 (N_29607,N_26288,N_25683);
and U29608 (N_29608,N_25582,N_26828);
or U29609 (N_29609,N_26149,N_26496);
xnor U29610 (N_29610,N_26164,N_26628);
and U29611 (N_29611,N_26487,N_26773);
and U29612 (N_29612,N_27206,N_27428);
xor U29613 (N_29613,N_27248,N_27300);
nor U29614 (N_29614,N_26804,N_25245);
and U29615 (N_29615,N_26234,N_26087);
nand U29616 (N_29616,N_27367,N_25259);
and U29617 (N_29617,N_25441,N_26741);
and U29618 (N_29618,N_26661,N_26841);
nor U29619 (N_29619,N_26031,N_25232);
and U29620 (N_29620,N_25213,N_26250);
or U29621 (N_29621,N_26722,N_25791);
xnor U29622 (N_29622,N_25251,N_25564);
and U29623 (N_29623,N_25228,N_25410);
nor U29624 (N_29624,N_26257,N_26790);
nor U29625 (N_29625,N_25685,N_25821);
and U29626 (N_29626,N_25607,N_26383);
xor U29627 (N_29627,N_25521,N_25182);
and U29628 (N_29628,N_27243,N_25180);
and U29629 (N_29629,N_26910,N_25822);
and U29630 (N_29630,N_25160,N_27375);
and U29631 (N_29631,N_25742,N_26653);
xor U29632 (N_29632,N_27167,N_26649);
and U29633 (N_29633,N_27382,N_27177);
nand U29634 (N_29634,N_25001,N_26142);
or U29635 (N_29635,N_26391,N_26793);
nand U29636 (N_29636,N_26629,N_26667);
and U29637 (N_29637,N_25562,N_25558);
or U29638 (N_29638,N_26872,N_26275);
xor U29639 (N_29639,N_26150,N_25617);
or U29640 (N_29640,N_27032,N_27193);
xor U29641 (N_29641,N_26324,N_25041);
or U29642 (N_29642,N_26119,N_27415);
or U29643 (N_29643,N_26197,N_25680);
xor U29644 (N_29644,N_25819,N_25653);
xor U29645 (N_29645,N_25046,N_25423);
nor U29646 (N_29646,N_26728,N_25020);
nand U29647 (N_29647,N_25430,N_26814);
and U29648 (N_29648,N_27236,N_25990);
xnor U29649 (N_29649,N_25470,N_27480);
and U29650 (N_29650,N_26258,N_25591);
nand U29651 (N_29651,N_26380,N_26223);
xor U29652 (N_29652,N_25238,N_25858);
or U29653 (N_29653,N_25327,N_25456);
nor U29654 (N_29654,N_26988,N_27069);
nor U29655 (N_29655,N_25373,N_26513);
xnor U29656 (N_29656,N_26920,N_26562);
and U29657 (N_29657,N_26739,N_25869);
nor U29658 (N_29658,N_25102,N_25236);
nand U29659 (N_29659,N_26678,N_25036);
and U29660 (N_29660,N_26196,N_25505);
nor U29661 (N_29661,N_26289,N_25215);
or U29662 (N_29662,N_27409,N_26819);
nor U29663 (N_29663,N_27150,N_25385);
or U29664 (N_29664,N_27080,N_25685);
and U29665 (N_29665,N_27344,N_26652);
or U29666 (N_29666,N_27404,N_25695);
and U29667 (N_29667,N_27392,N_27107);
or U29668 (N_29668,N_26512,N_25330);
nor U29669 (N_29669,N_25401,N_26676);
xnor U29670 (N_29670,N_25080,N_25016);
xnor U29671 (N_29671,N_27059,N_25040);
or U29672 (N_29672,N_26154,N_26600);
nand U29673 (N_29673,N_26409,N_25977);
nand U29674 (N_29674,N_26747,N_26492);
xor U29675 (N_29675,N_26201,N_26770);
and U29676 (N_29676,N_26960,N_25019);
nand U29677 (N_29677,N_27060,N_25147);
and U29678 (N_29678,N_27440,N_27375);
and U29679 (N_29679,N_25682,N_25976);
or U29680 (N_29680,N_25603,N_25917);
xnor U29681 (N_29681,N_25919,N_26766);
nand U29682 (N_29682,N_25468,N_26069);
and U29683 (N_29683,N_25745,N_26798);
and U29684 (N_29684,N_26790,N_26920);
nor U29685 (N_29685,N_26326,N_25779);
nor U29686 (N_29686,N_27299,N_25734);
nor U29687 (N_29687,N_25797,N_26229);
and U29688 (N_29688,N_27229,N_26359);
xnor U29689 (N_29689,N_25756,N_25693);
or U29690 (N_29690,N_26142,N_27382);
or U29691 (N_29691,N_26432,N_27456);
and U29692 (N_29692,N_26258,N_25209);
nand U29693 (N_29693,N_25223,N_26009);
xnor U29694 (N_29694,N_26498,N_25677);
or U29695 (N_29695,N_26272,N_27271);
or U29696 (N_29696,N_25598,N_25743);
or U29697 (N_29697,N_26025,N_27355);
nand U29698 (N_29698,N_27333,N_27414);
xor U29699 (N_29699,N_27015,N_26190);
xor U29700 (N_29700,N_27243,N_25958);
nand U29701 (N_29701,N_26945,N_26145);
nand U29702 (N_29702,N_27390,N_26558);
nor U29703 (N_29703,N_26599,N_25261);
or U29704 (N_29704,N_26329,N_27160);
or U29705 (N_29705,N_27164,N_25164);
nor U29706 (N_29706,N_26556,N_25819);
nor U29707 (N_29707,N_26961,N_27101);
nor U29708 (N_29708,N_26163,N_26949);
xnor U29709 (N_29709,N_26951,N_25011);
and U29710 (N_29710,N_26383,N_27427);
or U29711 (N_29711,N_27139,N_26299);
xor U29712 (N_29712,N_26127,N_25097);
nor U29713 (N_29713,N_27495,N_27463);
nor U29714 (N_29714,N_26096,N_26123);
nor U29715 (N_29715,N_26416,N_25007);
nand U29716 (N_29716,N_27360,N_27422);
and U29717 (N_29717,N_26264,N_27104);
and U29718 (N_29718,N_25829,N_25220);
or U29719 (N_29719,N_25224,N_25398);
nor U29720 (N_29720,N_27355,N_25670);
xnor U29721 (N_29721,N_26154,N_25085);
nand U29722 (N_29722,N_27455,N_26413);
nand U29723 (N_29723,N_27280,N_25713);
and U29724 (N_29724,N_27071,N_25710);
xnor U29725 (N_29725,N_26882,N_26645);
xor U29726 (N_29726,N_25801,N_25360);
or U29727 (N_29727,N_26949,N_25297);
nor U29728 (N_29728,N_25080,N_25059);
xor U29729 (N_29729,N_26094,N_26221);
nor U29730 (N_29730,N_25667,N_26976);
or U29731 (N_29731,N_25921,N_25274);
nor U29732 (N_29732,N_25358,N_27369);
or U29733 (N_29733,N_25390,N_27390);
xnor U29734 (N_29734,N_26901,N_26462);
and U29735 (N_29735,N_25148,N_26306);
xor U29736 (N_29736,N_25948,N_26135);
and U29737 (N_29737,N_26264,N_26792);
nand U29738 (N_29738,N_25004,N_25171);
or U29739 (N_29739,N_25683,N_26930);
nand U29740 (N_29740,N_27249,N_27124);
xor U29741 (N_29741,N_26732,N_27318);
xnor U29742 (N_29742,N_26814,N_26673);
nor U29743 (N_29743,N_27439,N_25197);
nor U29744 (N_29744,N_25613,N_25289);
nor U29745 (N_29745,N_27309,N_25673);
xnor U29746 (N_29746,N_25768,N_26531);
nor U29747 (N_29747,N_26343,N_25566);
nor U29748 (N_29748,N_25053,N_26311);
nand U29749 (N_29749,N_25267,N_26677);
xor U29750 (N_29750,N_25614,N_26564);
xor U29751 (N_29751,N_25177,N_26892);
or U29752 (N_29752,N_27124,N_26763);
or U29753 (N_29753,N_25232,N_26071);
nor U29754 (N_29754,N_25115,N_25232);
xnor U29755 (N_29755,N_27368,N_25693);
and U29756 (N_29756,N_25760,N_26950);
nand U29757 (N_29757,N_25203,N_26999);
or U29758 (N_29758,N_27217,N_27059);
and U29759 (N_29759,N_26656,N_26346);
and U29760 (N_29760,N_26314,N_25070);
nand U29761 (N_29761,N_27161,N_25535);
or U29762 (N_29762,N_25910,N_26934);
and U29763 (N_29763,N_26772,N_26807);
nor U29764 (N_29764,N_27003,N_26650);
nand U29765 (N_29765,N_26534,N_25369);
or U29766 (N_29766,N_26107,N_26856);
nor U29767 (N_29767,N_27186,N_25329);
nand U29768 (N_29768,N_26451,N_25607);
and U29769 (N_29769,N_26600,N_27252);
and U29770 (N_29770,N_27442,N_25077);
and U29771 (N_29771,N_25122,N_25077);
xor U29772 (N_29772,N_27365,N_26262);
nor U29773 (N_29773,N_26502,N_26384);
nand U29774 (N_29774,N_26426,N_26665);
nor U29775 (N_29775,N_26665,N_27320);
xor U29776 (N_29776,N_26533,N_25730);
and U29777 (N_29777,N_27112,N_25586);
and U29778 (N_29778,N_25879,N_25303);
xnor U29779 (N_29779,N_27497,N_26795);
or U29780 (N_29780,N_25076,N_25924);
nand U29781 (N_29781,N_26284,N_25764);
xnor U29782 (N_29782,N_27301,N_27172);
and U29783 (N_29783,N_25214,N_27067);
xor U29784 (N_29784,N_27305,N_27029);
nor U29785 (N_29785,N_25046,N_26556);
nor U29786 (N_29786,N_26502,N_25425);
xnor U29787 (N_29787,N_25394,N_26940);
nor U29788 (N_29788,N_25800,N_27171);
and U29789 (N_29789,N_26694,N_25853);
or U29790 (N_29790,N_25737,N_25583);
nor U29791 (N_29791,N_25194,N_26784);
nor U29792 (N_29792,N_25906,N_26375);
xor U29793 (N_29793,N_25961,N_25489);
xnor U29794 (N_29794,N_26986,N_27149);
xor U29795 (N_29795,N_25248,N_26885);
nor U29796 (N_29796,N_25800,N_26108);
or U29797 (N_29797,N_26544,N_25231);
nor U29798 (N_29798,N_26815,N_26875);
nand U29799 (N_29799,N_25667,N_25393);
and U29800 (N_29800,N_27417,N_26572);
nor U29801 (N_29801,N_27486,N_26069);
xnor U29802 (N_29802,N_25771,N_25281);
xnor U29803 (N_29803,N_27218,N_25556);
and U29804 (N_29804,N_27338,N_27041);
xor U29805 (N_29805,N_26738,N_25052);
nor U29806 (N_29806,N_26488,N_26875);
and U29807 (N_29807,N_25359,N_25318);
xnor U29808 (N_29808,N_25665,N_25998);
nor U29809 (N_29809,N_26977,N_26232);
xnor U29810 (N_29810,N_25928,N_25017);
nor U29811 (N_29811,N_27046,N_26823);
nor U29812 (N_29812,N_25330,N_25186);
xnor U29813 (N_29813,N_27384,N_25630);
nand U29814 (N_29814,N_25414,N_27457);
xnor U29815 (N_29815,N_26533,N_26950);
xor U29816 (N_29816,N_26081,N_25598);
or U29817 (N_29817,N_25472,N_26915);
xnor U29818 (N_29818,N_25508,N_26443);
xor U29819 (N_29819,N_25576,N_26730);
xor U29820 (N_29820,N_25245,N_25427);
or U29821 (N_29821,N_26986,N_25753);
nand U29822 (N_29822,N_25936,N_27106);
or U29823 (N_29823,N_26157,N_27183);
nand U29824 (N_29824,N_26356,N_26955);
nor U29825 (N_29825,N_27487,N_26389);
and U29826 (N_29826,N_25585,N_26055);
or U29827 (N_29827,N_26735,N_26928);
nand U29828 (N_29828,N_26485,N_26972);
or U29829 (N_29829,N_27320,N_26341);
xor U29830 (N_29830,N_26640,N_25640);
nor U29831 (N_29831,N_25326,N_25455);
nor U29832 (N_29832,N_25464,N_26916);
and U29833 (N_29833,N_26432,N_25833);
nand U29834 (N_29834,N_26104,N_26767);
or U29835 (N_29835,N_27338,N_25071);
nor U29836 (N_29836,N_25379,N_26166);
nand U29837 (N_29837,N_26296,N_25955);
nand U29838 (N_29838,N_26889,N_25959);
nor U29839 (N_29839,N_25433,N_27078);
xor U29840 (N_29840,N_27113,N_25199);
xnor U29841 (N_29841,N_26806,N_26985);
or U29842 (N_29842,N_25914,N_26244);
nor U29843 (N_29843,N_26505,N_26332);
or U29844 (N_29844,N_27226,N_26191);
or U29845 (N_29845,N_25407,N_25991);
and U29846 (N_29846,N_25061,N_26422);
and U29847 (N_29847,N_25718,N_26668);
and U29848 (N_29848,N_25185,N_27388);
nand U29849 (N_29849,N_26416,N_25490);
and U29850 (N_29850,N_26203,N_26688);
and U29851 (N_29851,N_26778,N_26386);
or U29852 (N_29852,N_25326,N_25785);
and U29853 (N_29853,N_26989,N_26987);
nor U29854 (N_29854,N_25070,N_25740);
xnor U29855 (N_29855,N_26865,N_25273);
nor U29856 (N_29856,N_25502,N_25270);
xnor U29857 (N_29857,N_26703,N_27371);
nand U29858 (N_29858,N_26432,N_27425);
or U29859 (N_29859,N_27143,N_26459);
nor U29860 (N_29860,N_27184,N_25919);
and U29861 (N_29861,N_25678,N_27069);
or U29862 (N_29862,N_25966,N_26839);
nand U29863 (N_29863,N_25595,N_27484);
and U29864 (N_29864,N_25795,N_27434);
and U29865 (N_29865,N_25370,N_26585);
or U29866 (N_29866,N_26369,N_27469);
xnor U29867 (N_29867,N_25089,N_25979);
and U29868 (N_29868,N_26011,N_26288);
nand U29869 (N_29869,N_27310,N_26274);
xor U29870 (N_29870,N_26430,N_26266);
and U29871 (N_29871,N_26690,N_25291);
nand U29872 (N_29872,N_26920,N_27394);
or U29873 (N_29873,N_26538,N_25357);
xnor U29874 (N_29874,N_26191,N_25016);
nor U29875 (N_29875,N_25866,N_27389);
and U29876 (N_29876,N_26563,N_26333);
xor U29877 (N_29877,N_25106,N_26984);
nor U29878 (N_29878,N_25856,N_25527);
and U29879 (N_29879,N_26651,N_26208);
and U29880 (N_29880,N_25149,N_26117);
and U29881 (N_29881,N_25972,N_25509);
or U29882 (N_29882,N_25011,N_25541);
nor U29883 (N_29883,N_26161,N_25785);
and U29884 (N_29884,N_25271,N_27094);
nand U29885 (N_29885,N_26234,N_27340);
nor U29886 (N_29886,N_27260,N_25980);
nor U29887 (N_29887,N_25493,N_26381);
or U29888 (N_29888,N_25948,N_26501);
and U29889 (N_29889,N_26075,N_26610);
nor U29890 (N_29890,N_25577,N_26135);
or U29891 (N_29891,N_25125,N_25923);
or U29892 (N_29892,N_25004,N_25188);
xnor U29893 (N_29893,N_26947,N_26437);
nand U29894 (N_29894,N_26981,N_26870);
xnor U29895 (N_29895,N_25889,N_25915);
xnor U29896 (N_29896,N_26187,N_25167);
or U29897 (N_29897,N_26034,N_25477);
and U29898 (N_29898,N_25307,N_26268);
nor U29899 (N_29899,N_27106,N_26027);
or U29900 (N_29900,N_25043,N_26235);
xor U29901 (N_29901,N_25541,N_25306);
nor U29902 (N_29902,N_25486,N_27377);
xnor U29903 (N_29903,N_26702,N_25067);
nor U29904 (N_29904,N_27048,N_25372);
and U29905 (N_29905,N_26491,N_25520);
xor U29906 (N_29906,N_26355,N_26281);
xnor U29907 (N_29907,N_27309,N_25660);
and U29908 (N_29908,N_27340,N_26080);
or U29909 (N_29909,N_26582,N_25418);
xnor U29910 (N_29910,N_25204,N_25647);
nand U29911 (N_29911,N_25693,N_25330);
xor U29912 (N_29912,N_25179,N_26472);
and U29913 (N_29913,N_27173,N_26907);
or U29914 (N_29914,N_26887,N_26431);
nor U29915 (N_29915,N_26873,N_27255);
xnor U29916 (N_29916,N_25742,N_25129);
nor U29917 (N_29917,N_25332,N_26902);
and U29918 (N_29918,N_25151,N_25649);
or U29919 (N_29919,N_26811,N_25179);
nand U29920 (N_29920,N_25510,N_27037);
xnor U29921 (N_29921,N_26543,N_26419);
xor U29922 (N_29922,N_27433,N_25130);
or U29923 (N_29923,N_27064,N_25484);
nand U29924 (N_29924,N_26707,N_25773);
and U29925 (N_29925,N_25195,N_25989);
xor U29926 (N_29926,N_27297,N_27095);
nand U29927 (N_29927,N_25391,N_25245);
or U29928 (N_29928,N_25925,N_26985);
nor U29929 (N_29929,N_25249,N_26477);
xnor U29930 (N_29930,N_25044,N_25789);
nand U29931 (N_29931,N_27073,N_26712);
and U29932 (N_29932,N_27470,N_26116);
or U29933 (N_29933,N_25378,N_25551);
nor U29934 (N_29934,N_27114,N_25842);
nor U29935 (N_29935,N_26596,N_25645);
and U29936 (N_29936,N_26667,N_27339);
and U29937 (N_29937,N_26192,N_25635);
nor U29938 (N_29938,N_27005,N_27403);
xor U29939 (N_29939,N_26051,N_26935);
xor U29940 (N_29940,N_25528,N_25620);
or U29941 (N_29941,N_25374,N_25072);
nand U29942 (N_29942,N_25391,N_26088);
nor U29943 (N_29943,N_25349,N_25392);
xor U29944 (N_29944,N_26999,N_25671);
nor U29945 (N_29945,N_27430,N_27091);
nor U29946 (N_29946,N_25508,N_26949);
xnor U29947 (N_29947,N_25749,N_26990);
nand U29948 (N_29948,N_26203,N_25045);
nor U29949 (N_29949,N_26067,N_25597);
and U29950 (N_29950,N_25499,N_25466);
and U29951 (N_29951,N_27269,N_26065);
or U29952 (N_29952,N_27065,N_26085);
nand U29953 (N_29953,N_27499,N_26474);
or U29954 (N_29954,N_26619,N_26927);
nor U29955 (N_29955,N_25605,N_25736);
xnor U29956 (N_29956,N_27261,N_27320);
xnor U29957 (N_29957,N_25622,N_25863);
and U29958 (N_29958,N_26087,N_25816);
nand U29959 (N_29959,N_27489,N_26987);
nand U29960 (N_29960,N_25875,N_25328);
xor U29961 (N_29961,N_26437,N_26513);
xor U29962 (N_29962,N_26979,N_26126);
nand U29963 (N_29963,N_27486,N_26125);
xnor U29964 (N_29964,N_25176,N_25364);
or U29965 (N_29965,N_25158,N_27343);
and U29966 (N_29966,N_25673,N_26891);
nor U29967 (N_29967,N_26368,N_26700);
nand U29968 (N_29968,N_25361,N_25081);
nand U29969 (N_29969,N_27042,N_27107);
and U29970 (N_29970,N_25057,N_26087);
and U29971 (N_29971,N_26659,N_26592);
nand U29972 (N_29972,N_25959,N_26063);
xor U29973 (N_29973,N_26738,N_25317);
and U29974 (N_29974,N_27394,N_25050);
or U29975 (N_29975,N_25027,N_26556);
or U29976 (N_29976,N_25921,N_27235);
and U29977 (N_29977,N_25244,N_26273);
nor U29978 (N_29978,N_25987,N_26987);
and U29979 (N_29979,N_26726,N_25276);
and U29980 (N_29980,N_25965,N_25721);
and U29981 (N_29981,N_26540,N_25709);
or U29982 (N_29982,N_26690,N_25909);
or U29983 (N_29983,N_26770,N_26173);
and U29984 (N_29984,N_26657,N_25138);
and U29985 (N_29985,N_27057,N_27187);
nor U29986 (N_29986,N_26661,N_27409);
or U29987 (N_29987,N_25470,N_25242);
or U29988 (N_29988,N_27014,N_25216);
and U29989 (N_29989,N_25759,N_25800);
nand U29990 (N_29990,N_26830,N_25771);
and U29991 (N_29991,N_26977,N_26426);
and U29992 (N_29992,N_27304,N_26328);
xnor U29993 (N_29993,N_26163,N_26584);
xnor U29994 (N_29994,N_26118,N_25603);
and U29995 (N_29995,N_27145,N_26667);
xor U29996 (N_29996,N_27163,N_26856);
nand U29997 (N_29997,N_27160,N_26076);
nand U29998 (N_29998,N_26093,N_26030);
and U29999 (N_29999,N_26992,N_25609);
nor U30000 (N_30000,N_28666,N_29687);
nor U30001 (N_30001,N_28956,N_29481);
xor U30002 (N_30002,N_29356,N_27627);
xnor U30003 (N_30003,N_29798,N_28331);
nor U30004 (N_30004,N_28382,N_28760);
and U30005 (N_30005,N_27537,N_29061);
or U30006 (N_30006,N_29615,N_29790);
and U30007 (N_30007,N_28966,N_27767);
nor U30008 (N_30008,N_28509,N_27920);
nor U30009 (N_30009,N_27662,N_27727);
or U30010 (N_30010,N_27536,N_27512);
nand U30011 (N_30011,N_29351,N_29906);
nand U30012 (N_30012,N_28819,N_28582);
nor U30013 (N_30013,N_29966,N_28129);
and U30014 (N_30014,N_28820,N_29309);
nor U30015 (N_30015,N_27672,N_29929);
nand U30016 (N_30016,N_29435,N_28886);
nand U30017 (N_30017,N_29197,N_28071);
or U30018 (N_30018,N_28965,N_29415);
nand U30019 (N_30019,N_29577,N_28987);
or U30020 (N_30020,N_29680,N_28437);
nand U30021 (N_30021,N_28789,N_29778);
xnor U30022 (N_30022,N_29525,N_27538);
or U30023 (N_30023,N_29465,N_28799);
xnor U30024 (N_30024,N_29248,N_29177);
and U30025 (N_30025,N_28602,N_29018);
or U30026 (N_30026,N_29382,N_27882);
and U30027 (N_30027,N_29717,N_29972);
nor U30028 (N_30028,N_28366,N_28074);
or U30029 (N_30029,N_28910,N_29802);
or U30030 (N_30030,N_27744,N_27829);
nor U30031 (N_30031,N_28157,N_29064);
xor U30032 (N_30032,N_29576,N_28864);
xnor U30033 (N_30033,N_29488,N_29907);
xnor U30034 (N_30034,N_28455,N_27830);
xnor U30035 (N_30035,N_27603,N_28306);
nand U30036 (N_30036,N_28649,N_27885);
and U30037 (N_30037,N_29119,N_28568);
or U30038 (N_30038,N_27584,N_28988);
and U30039 (N_30039,N_27803,N_29120);
nor U30040 (N_30040,N_29772,N_29083);
nor U30041 (N_30041,N_28131,N_29512);
nand U30042 (N_30042,N_29982,N_28968);
xnor U30043 (N_30043,N_29908,N_29000);
or U30044 (N_30044,N_28749,N_29241);
xnor U30045 (N_30045,N_28177,N_28929);
and U30046 (N_30046,N_28373,N_28462);
xor U30047 (N_30047,N_28089,N_29400);
and U30048 (N_30048,N_28836,N_27894);
nand U30049 (N_30049,N_28942,N_29417);
nand U30050 (N_30050,N_28055,N_29975);
or U30051 (N_30051,N_27625,N_29223);
xor U30052 (N_30052,N_28849,N_28238);
xnor U30053 (N_30053,N_29682,N_29720);
and U30054 (N_30054,N_28931,N_27966);
and U30055 (N_30055,N_29125,N_29602);
nor U30056 (N_30056,N_27516,N_28169);
nor U30057 (N_30057,N_28706,N_29338);
or U30058 (N_30058,N_29865,N_28793);
nor U30059 (N_30059,N_28109,N_29226);
or U30060 (N_30060,N_29864,N_28119);
nor U30061 (N_30061,N_29216,N_29664);
or U30062 (N_30062,N_29314,N_28911);
nand U30063 (N_30063,N_28897,N_29496);
or U30064 (N_30064,N_28404,N_28126);
and U30065 (N_30065,N_28691,N_28673);
and U30066 (N_30066,N_29042,N_29806);
and U30067 (N_30067,N_29339,N_29175);
xnor U30068 (N_30068,N_28435,N_27707);
nand U30069 (N_30069,N_29570,N_28683);
nand U30070 (N_30070,N_29500,N_28241);
and U30071 (N_30071,N_28608,N_29277);
and U30072 (N_30072,N_27589,N_28091);
xnor U30073 (N_30073,N_29058,N_28046);
or U30074 (N_30074,N_29893,N_28226);
nor U30075 (N_30075,N_28719,N_28664);
nor U30076 (N_30076,N_29764,N_28090);
nand U30077 (N_30077,N_28633,N_29821);
nand U30078 (N_30078,N_27757,N_27857);
or U30079 (N_30079,N_28312,N_28040);
xnor U30080 (N_30080,N_27503,N_28518);
xor U30081 (N_30081,N_28287,N_27881);
or U30082 (N_30082,N_27705,N_29200);
and U30083 (N_30083,N_29750,N_28165);
nand U30084 (N_30084,N_29705,N_29921);
xor U30085 (N_30085,N_28184,N_28181);
nand U30086 (N_30086,N_28393,N_27813);
xnor U30087 (N_30087,N_28768,N_29983);
and U30088 (N_30088,N_27559,N_28280);
nor U30089 (N_30089,N_29044,N_29350);
nand U30090 (N_30090,N_28266,N_28646);
xor U30091 (N_30091,N_28637,N_29814);
and U30092 (N_30092,N_28619,N_27545);
and U30093 (N_30093,N_28028,N_29552);
nor U30094 (N_30094,N_28239,N_27546);
or U30095 (N_30095,N_29286,N_27810);
nor U30096 (N_30096,N_28984,N_29089);
or U30097 (N_30097,N_27916,N_29961);
xor U30098 (N_30098,N_28653,N_27549);
and U30099 (N_30099,N_29676,N_29775);
nand U30100 (N_30100,N_29396,N_28363);
nor U30101 (N_30101,N_29546,N_28970);
xor U30102 (N_30102,N_29768,N_28686);
or U30103 (N_30103,N_28511,N_27815);
or U30104 (N_30104,N_28185,N_28422);
and U30105 (N_30105,N_27945,N_28122);
nor U30106 (N_30106,N_27568,N_29548);
or U30107 (N_30107,N_28740,N_28788);
nor U30108 (N_30108,N_28357,N_29914);
nor U30109 (N_30109,N_29431,N_29981);
xnor U30110 (N_30110,N_28172,N_29071);
nor U30111 (N_30111,N_29272,N_28564);
and U30112 (N_30112,N_27930,N_28873);
nand U30113 (N_30113,N_29006,N_27636);
or U30114 (N_30114,N_28595,N_27775);
nor U30115 (N_30115,N_29357,N_29796);
or U30116 (N_30116,N_29078,N_28918);
nor U30117 (N_30117,N_29800,N_28985);
and U30118 (N_30118,N_27939,N_28806);
nand U30119 (N_30119,N_27796,N_29084);
and U30120 (N_30120,N_29183,N_28946);
nor U30121 (N_30121,N_29143,N_29222);
and U30122 (N_30122,N_29569,N_29575);
nor U30123 (N_30123,N_27761,N_28812);
xnor U30124 (N_30124,N_27746,N_27729);
nand U30125 (N_30125,N_28330,N_28412);
or U30126 (N_30126,N_27667,N_28835);
nand U30127 (N_30127,N_28879,N_29180);
and U30128 (N_30128,N_28452,N_29848);
and U30129 (N_30129,N_29059,N_27977);
or U30130 (N_30130,N_28979,N_28097);
nand U30131 (N_30131,N_29360,N_29507);
xnor U30132 (N_30132,N_29746,N_27991);
xnor U30133 (N_30133,N_28187,N_29527);
nor U30134 (N_30134,N_29697,N_29267);
nor U30135 (N_30135,N_28599,N_28207);
xor U30136 (N_30136,N_28853,N_29031);
and U30137 (N_30137,N_28803,N_29532);
and U30138 (N_30138,N_28701,N_29827);
and U30139 (N_30139,N_29699,N_27909);
and U30140 (N_30140,N_27681,N_27583);
and U30141 (N_30141,N_28865,N_28659);
nor U30142 (N_30142,N_29509,N_27755);
and U30143 (N_30143,N_28831,N_29101);
or U30144 (N_30144,N_29539,N_28792);
nand U30145 (N_30145,N_29787,N_29079);
or U30146 (N_30146,N_28240,N_28677);
nor U30147 (N_30147,N_29348,N_28919);
nand U30148 (N_30148,N_27561,N_29232);
and U30149 (N_30149,N_29930,N_28707);
and U30150 (N_30150,N_29766,N_29478);
nand U30151 (N_30151,N_28051,N_29932);
xor U30152 (N_30152,N_29337,N_28903);
nor U30153 (N_30153,N_27782,N_28379);
nor U30154 (N_30154,N_29163,N_28142);
xnor U30155 (N_30155,N_28329,N_29733);
nor U30156 (N_30156,N_28250,N_27696);
xnor U30157 (N_30157,N_29088,N_28874);
nand U30158 (N_30158,N_29178,N_29863);
and U30159 (N_30159,N_29832,N_28496);
xnor U30160 (N_30160,N_28025,N_29898);
or U30161 (N_30161,N_29829,N_29165);
and U30162 (N_30162,N_29938,N_28426);
nand U30163 (N_30163,N_28163,N_28210);
and U30164 (N_30164,N_29943,N_28584);
or U30165 (N_30165,N_29553,N_29991);
nand U30166 (N_30166,N_29156,N_28322);
nor U30167 (N_30167,N_27812,N_28692);
xnor U30168 (N_30168,N_27798,N_28481);
xnor U30169 (N_30169,N_28349,N_28538);
nand U30170 (N_30170,N_27818,N_29645);
nand U30171 (N_30171,N_28112,N_27514);
nor U30172 (N_30172,N_29288,N_29020);
and U30173 (N_30173,N_28394,N_27995);
nand U30174 (N_30174,N_27917,N_28998);
and U30175 (N_30175,N_27821,N_28223);
nor U30176 (N_30176,N_28297,N_27927);
nand U30177 (N_30177,N_27774,N_29955);
nand U30178 (N_30178,N_27621,N_27880);
nand U30179 (N_30179,N_29845,N_28851);
or U30180 (N_30180,N_28283,N_28052);
nand U30181 (N_30181,N_27663,N_29792);
nor U30182 (N_30182,N_29959,N_28606);
xnor U30183 (N_30183,N_28615,N_28704);
nand U30184 (N_30184,N_27527,N_28020);
and U30185 (N_30185,N_29202,N_29106);
nor U30186 (N_30186,N_28004,N_28908);
nor U30187 (N_30187,N_29028,N_28273);
nand U30188 (N_30188,N_28976,N_27724);
nor U30189 (N_30189,N_27997,N_29246);
nand U30190 (N_30190,N_27837,N_27865);
nor U30191 (N_30191,N_29336,N_29536);
xor U30192 (N_30192,N_29451,N_28631);
and U30193 (N_30193,N_29873,N_28450);
nand U30194 (N_30194,N_28365,N_29640);
or U30195 (N_30195,N_28828,N_29940);
nand U30196 (N_30196,N_27982,N_29196);
or U30197 (N_30197,N_28863,N_29504);
nor U30198 (N_30198,N_29540,N_29545);
xor U30199 (N_30199,N_27677,N_28001);
or U30200 (N_30200,N_27553,N_27906);
xor U30201 (N_30201,N_29278,N_28640);
and U30202 (N_30202,N_27780,N_28641);
nor U30203 (N_30203,N_29784,N_27600);
nor U30204 (N_30204,N_28360,N_29926);
or U30205 (N_30205,N_27935,N_27648);
xor U30206 (N_30206,N_28033,N_29249);
or U30207 (N_30207,N_28141,N_29115);
or U30208 (N_30208,N_29203,N_28424);
and U30209 (N_30209,N_28676,N_29153);
nor U30210 (N_30210,N_28500,N_27988);
xnor U30211 (N_30211,N_29148,N_28433);
xor U30212 (N_30212,N_28943,N_28419);
xnor U30213 (N_30213,N_27593,N_28662);
and U30214 (N_30214,N_27522,N_28443);
or U30215 (N_30215,N_29641,N_29100);
or U30216 (N_30216,N_27715,N_27624);
and U30217 (N_30217,N_29783,N_28952);
nor U30218 (N_30218,N_29041,N_28661);
or U30219 (N_30219,N_28274,N_28403);
or U30220 (N_30220,N_29137,N_29639);
nor U30221 (N_30221,N_29953,N_28095);
nor U30222 (N_30222,N_28711,N_29619);
and U30223 (N_30223,N_28871,N_29543);
or U30224 (N_30224,N_29037,N_28242);
or U30225 (N_30225,N_29582,N_27690);
nand U30226 (N_30226,N_29726,N_27855);
nor U30227 (N_30227,N_28688,N_28577);
and U30228 (N_30228,N_29220,N_28024);
xnor U30229 (N_30229,N_27876,N_28983);
or U30230 (N_30230,N_29114,N_28735);
nand U30231 (N_30231,N_27651,N_29367);
nor U30232 (N_30232,N_29996,N_28588);
nor U30233 (N_30233,N_29457,N_28159);
and U30234 (N_30234,N_28405,N_28726);
nor U30235 (N_30235,N_29716,N_27893);
and U30236 (N_30236,N_27858,N_29759);
or U30237 (N_30237,N_27763,N_28473);
nor U30238 (N_30238,N_29070,N_29791);
and U30239 (N_30239,N_29568,N_27776);
xnor U30240 (N_30240,N_27567,N_28124);
nor U30241 (N_30241,N_29774,N_28470);
nor U30242 (N_30242,N_28385,N_27571);
xnor U30243 (N_30243,N_28775,N_29690);
nor U30244 (N_30244,N_28906,N_29564);
nand U30245 (N_30245,N_28939,N_28368);
or U30246 (N_30246,N_29506,N_29852);
or U30247 (N_30247,N_27606,N_28374);
nor U30248 (N_30248,N_27609,N_29069);
or U30249 (N_30249,N_29428,N_28559);
and U30250 (N_30250,N_29743,N_27564);
xnor U30251 (N_30251,N_29316,N_29014);
and U30252 (N_30252,N_29138,N_29741);
xor U30253 (N_30253,N_28591,N_27823);
nor U30254 (N_30254,N_29621,N_29583);
nor U30255 (N_30255,N_29696,N_28940);
xnor U30256 (N_30256,N_28460,N_28060);
xor U30257 (N_30257,N_29811,N_27740);
or U30258 (N_30258,N_28624,N_29096);
nand U30259 (N_30259,N_28202,N_27720);
xor U30260 (N_30260,N_29698,N_28947);
nor U30261 (N_30261,N_29756,N_27628);
nand U30262 (N_30262,N_28010,N_28478);
and U30263 (N_30263,N_28147,N_29198);
or U30264 (N_30264,N_27750,N_29970);
nor U30265 (N_30265,N_27697,N_28698);
nand U30266 (N_30266,N_29007,N_27846);
and U30267 (N_30267,N_28534,N_29067);
nor U30268 (N_30268,N_27731,N_28720);
nor U30269 (N_30269,N_28138,N_28255);
xnor U30270 (N_30270,N_28351,N_27572);
nor U30271 (N_30271,N_29703,N_28769);
nor U30272 (N_30272,N_27862,N_27765);
nor U30273 (N_30273,N_27668,N_28440);
nor U30274 (N_30274,N_28161,N_29477);
nand U30275 (N_30275,N_29313,N_29586);
or U30276 (N_30276,N_29307,N_28042);
nor U30277 (N_30277,N_29857,N_28288);
or U30278 (N_30278,N_29472,N_29954);
nor U30279 (N_30279,N_27869,N_29994);
or U30280 (N_30280,N_29322,N_29389);
and U30281 (N_30281,N_27526,N_27585);
xor U30282 (N_30282,N_28795,N_28798);
nand U30283 (N_30283,N_28220,N_27598);
xor U30284 (N_30284,N_27878,N_29380);
xnor U30285 (N_30285,N_28464,N_29381);
nor U30286 (N_30286,N_28829,N_29474);
xnor U30287 (N_30287,N_29660,N_27695);
nor U30288 (N_30288,N_28684,N_28309);
nand U30289 (N_30289,N_27983,N_27785);
nor U30290 (N_30290,N_27708,N_28291);
nor U30291 (N_30291,N_29779,N_27502);
and U30292 (N_30292,N_28444,N_29134);
and U30293 (N_30293,N_28043,N_28826);
and U30294 (N_30294,N_27847,N_29529);
xor U30295 (N_30295,N_29364,N_29133);
or U30296 (N_30296,N_28376,N_29298);
or U30297 (N_30297,N_27874,N_28638);
or U30298 (N_30298,N_27655,N_29949);
and U30299 (N_30299,N_29468,N_29522);
nor U30300 (N_30300,N_27769,N_27868);
xnor U30301 (N_30301,N_29519,N_28693);
or U30302 (N_30302,N_27670,N_29127);
and U30303 (N_30303,N_28652,N_28019);
nor U30304 (N_30304,N_28409,N_29080);
and U30305 (N_30305,N_29390,N_27658);
nand U30306 (N_30306,N_29378,N_29452);
nor U30307 (N_30307,N_29349,N_29537);
and U30308 (N_30308,N_28813,N_28535);
nor U30309 (N_30309,N_27808,N_29555);
and U30310 (N_30310,N_28108,N_28884);
nor U30311 (N_30311,N_28695,N_28963);
nand U30312 (N_30312,N_29421,N_29928);
nor U30313 (N_30313,N_27726,N_29822);
or U30314 (N_30314,N_27539,N_28816);
or U30315 (N_30315,N_29009,N_28567);
nor U30316 (N_30316,N_29185,N_29934);
nand U30317 (N_30317,N_29654,N_29201);
xor U30318 (N_30318,N_28145,N_29995);
nand U30319 (N_30319,N_29333,N_28318);
xnor U30320 (N_30320,N_27992,N_29151);
or U30321 (N_30321,N_29544,N_28018);
nor U30322 (N_30322,N_28411,N_27659);
xnor U30323 (N_30323,N_29366,N_28400);
and U30324 (N_30324,N_28486,N_29068);
and U30325 (N_30325,N_29590,N_29407);
xnor U30326 (N_30326,N_29793,N_29149);
or U30327 (N_30327,N_28175,N_28182);
nand U30328 (N_30328,N_28517,N_28296);
nor U30329 (N_30329,N_28209,N_27850);
nor U30330 (N_30330,N_29933,N_29235);
nor U30331 (N_30331,N_28503,N_29323);
and U30332 (N_30332,N_29347,N_28032);
xnor U30333 (N_30333,N_29139,N_28468);
nand U30334 (N_30334,N_28949,N_29866);
and U30335 (N_30335,N_29985,N_28315);
nor U30336 (N_30336,N_28362,N_28035);
or U30337 (N_30337,N_28383,N_28326);
nor U30338 (N_30338,N_29283,N_29076);
nor U30339 (N_30339,N_28601,N_28571);
and U30340 (N_30340,N_27678,N_27599);
nor U30341 (N_30341,N_28015,N_28747);
nand U30342 (N_30342,N_28603,N_28003);
xnor U30343 (N_30343,N_28094,N_29057);
nand U30344 (N_30344,N_27840,N_29158);
and U30345 (N_30345,N_29770,N_29160);
nand U30346 (N_30346,N_27899,N_29262);
nor U30347 (N_30347,N_29508,N_28030);
xnor U30348 (N_30348,N_29816,N_28992);
or U30349 (N_30349,N_29871,N_28780);
xor U30350 (N_30350,N_28834,N_29948);
and U30351 (N_30351,N_27519,N_29997);
and U30352 (N_30352,N_27816,N_29335);
xor U30353 (N_30353,N_29442,N_29399);
nor U30354 (N_30354,N_28989,N_29124);
or U30355 (N_30355,N_28777,N_29259);
xnor U30356 (N_30356,N_27657,N_27713);
xor U30357 (N_30357,N_29876,N_28300);
and U30358 (N_30358,N_28974,N_27973);
xnor U30359 (N_30359,N_28512,N_27811);
or U30360 (N_30360,N_28299,N_28805);
or U30361 (N_30361,N_29167,N_29731);
nor U30362 (N_30362,N_28176,N_28390);
nand U30363 (N_30363,N_28047,N_29082);
or U30364 (N_30364,N_28438,N_29825);
xnor U30365 (N_30365,N_27656,N_28017);
or U30366 (N_30366,N_29419,N_29869);
and U30367 (N_30367,N_28621,N_28905);
and U30368 (N_30368,N_28742,N_28204);
xnor U30369 (N_30369,N_29877,N_27569);
or U30370 (N_30370,N_29858,N_28230);
or U30371 (N_30371,N_28817,N_28581);
or U30372 (N_30372,N_29684,N_29651);
nand U30373 (N_30373,N_27711,N_27581);
nand U30374 (N_30374,N_29713,N_28924);
or U30375 (N_30375,N_28002,N_27704);
or U30376 (N_30376,N_29685,N_28941);
nor U30377 (N_30377,N_29980,N_29763);
xnor U30378 (N_30378,N_29300,N_27900);
nor U30379 (N_30379,N_28759,N_29293);
nand U30380 (N_30380,N_28665,N_28578);
nor U30381 (N_30381,N_29195,N_27682);
and U30382 (N_30382,N_29896,N_29861);
nor U30383 (N_30383,N_28079,N_28531);
and U30384 (N_30384,N_27630,N_27528);
and U30385 (N_30385,N_28476,N_29437);
nor U30386 (N_30386,N_28542,N_29686);
or U30387 (N_30387,N_28651,N_29188);
nand U30388 (N_30388,N_29960,N_29179);
nand U30389 (N_30389,N_28099,N_28006);
and U30390 (N_30390,N_28605,N_28823);
or U30391 (N_30391,N_28005,N_29269);
nand U30392 (N_30392,N_29758,N_29438);
nand U30393 (N_30393,N_29661,N_28292);
xor U30394 (N_30394,N_29765,N_29632);
xor U30395 (N_30395,N_29480,N_29986);
nand U30396 (N_30396,N_29150,N_28668);
and U30397 (N_30397,N_27501,N_29181);
xor U30398 (N_30398,N_28731,N_29749);
xnor U30399 (N_30399,N_27518,N_29923);
xor U30400 (N_30400,N_28340,N_27824);
xor U30401 (N_30401,N_27904,N_28703);
nor U30402 (N_30402,N_29393,N_28926);
nand U30403 (N_30403,N_29817,N_29211);
or U30404 (N_30404,N_29636,N_27666);
or U30405 (N_30405,N_29777,N_28549);
nand U30406 (N_30406,N_29190,N_28745);
and U30407 (N_30407,N_28957,N_28990);
and U30408 (N_30408,N_27680,N_29813);
xnor U30409 (N_30409,N_29579,N_27575);
or U30410 (N_30410,N_29842,N_29086);
and U30411 (N_30411,N_28967,N_28958);
nor U30412 (N_30412,N_29332,N_28771);
xnor U30413 (N_30413,N_28894,N_29939);
and U30414 (N_30414,N_29234,N_29571);
or U30415 (N_30415,N_28054,N_29650);
xor U30416 (N_30416,N_28281,N_29268);
xnor U30417 (N_30417,N_27807,N_28537);
nor U30418 (N_30418,N_28544,N_29951);
xnor U30419 (N_30419,N_28876,N_28741);
xor U30420 (N_30420,N_28845,N_27754);
xor U30421 (N_30421,N_29206,N_28574);
or U30422 (N_30422,N_28521,N_29862);
xor U30423 (N_30423,N_28530,N_28449);
or U30424 (N_30424,N_28494,N_28195);
and U30425 (N_30425,N_27962,N_27525);
xor U30426 (N_30426,N_29672,N_28007);
nor U30427 (N_30427,N_29841,N_28062);
nand U30428 (N_30428,N_27948,N_27943);
xnor U30429 (N_30429,N_29662,N_27717);
or U30430 (N_30430,N_29637,N_29767);
xnor U30431 (N_30431,N_27745,N_29285);
nor U30432 (N_30432,N_28136,N_29310);
xor U30433 (N_30433,N_29560,N_28675);
xor U30434 (N_30434,N_28179,N_29567);
nand U30435 (N_30435,N_28493,N_27601);
nand U30436 (N_30436,N_29999,N_29872);
or U30437 (N_30437,N_29912,N_28877);
and U30438 (N_30438,N_29788,N_28259);
or U30439 (N_30439,N_29372,N_29191);
nor U30440 (N_30440,N_28951,N_28102);
xnor U30441 (N_30441,N_28762,N_28474);
or U30442 (N_30442,N_29255,N_29312);
xor U30443 (N_30443,N_29919,N_29172);
or U30444 (N_30444,N_29388,N_29365);
xnor U30445 (N_30445,N_29060,N_29631);
and U30446 (N_30446,N_28682,N_28604);
nand U30447 (N_30447,N_28277,N_27958);
xnor U30448 (N_30448,N_29154,N_29725);
or U30449 (N_30449,N_29706,N_29883);
or U30450 (N_30450,N_29214,N_29225);
or U30451 (N_30451,N_27914,N_28216);
xor U30452 (N_30452,N_28037,N_29168);
xor U30453 (N_30453,N_27620,N_28279);
xnor U30454 (N_30454,N_28014,N_29711);
and U30455 (N_30455,N_28156,N_28272);
nor U30456 (N_30456,N_28846,N_29776);
xnor U30457 (N_30457,N_28858,N_28078);
xor U30458 (N_30458,N_28898,N_27867);
or U30459 (N_30459,N_28458,N_28050);
nor U30460 (N_30460,N_27961,N_29882);
and U30461 (N_30461,N_27779,N_28814);
or U30462 (N_30462,N_29394,N_28971);
nor U30463 (N_30463,N_29528,N_28038);
nand U30464 (N_30464,N_28061,N_28257);
xor U30465 (N_30465,N_27907,N_29353);
nand U30466 (N_30466,N_28441,N_29464);
xor U30467 (N_30467,N_29296,N_29950);
and U30468 (N_30468,N_29977,N_27936);
nand U30469 (N_30469,N_28192,N_28986);
xor U30470 (N_30470,N_28572,N_28372);
nor U30471 (N_30471,N_29847,N_29946);
nand U30472 (N_30472,N_29344,N_28067);
or U30473 (N_30473,N_28150,N_28059);
xnor U30474 (N_30474,N_29771,N_28727);
xnor U30475 (N_30475,N_28492,N_29423);
nor U30476 (N_30476,N_27642,N_27579);
nand U30477 (N_30477,N_28442,N_27739);
nor U30478 (N_30478,N_28151,N_27694);
xnor U30479 (N_30479,N_28513,N_28456);
nor U30480 (N_30480,N_29170,N_27856);
or U30481 (N_30481,N_28679,N_28323);
nor U30482 (N_30482,N_29284,N_29385);
nand U30483 (N_30483,N_28401,N_27998);
nand U30484 (N_30484,N_27712,N_29558);
xnor U30485 (N_30485,N_29701,N_27685);
and U30486 (N_30486,N_28261,N_27901);
nor U30487 (N_30487,N_29547,N_28350);
nor U30488 (N_30488,N_29655,N_28502);
xnor U30489 (N_30489,N_27741,N_27607);
or U30490 (N_30490,N_29988,N_29517);
xor U30491 (N_30491,N_27777,N_28066);
nand U30492 (N_30492,N_27786,N_28774);
xnor U30493 (N_30493,N_28739,N_28495);
nor U30494 (N_30494,N_28128,N_28713);
and U30495 (N_30495,N_28088,N_27849);
and U30496 (N_30496,N_29868,N_28121);
nand U30497 (N_30497,N_27950,N_29294);
and U30498 (N_30498,N_27762,N_29667);
nand U30499 (N_30499,N_29915,N_29092);
nand U30500 (N_30500,N_27535,N_29679);
xor U30501 (N_30501,N_29581,N_29922);
xor U30502 (N_30502,N_29709,N_27912);
xnor U30503 (N_30503,N_28585,N_29473);
nand U30504 (N_30504,N_27587,N_29434);
and U30505 (N_30505,N_29606,N_29623);
xor U30506 (N_30506,N_28840,N_28629);
nand U30507 (N_30507,N_28186,N_27887);
or U30508 (N_30508,N_28541,N_29224);
nand U30509 (N_30509,N_29984,N_28415);
xnor U30510 (N_30510,N_27721,N_29843);
xnor U30511 (N_30511,N_28302,N_29405);
xnor U30512 (N_30512,N_29511,N_28100);
nor U30513 (N_30513,N_29739,N_28252);
or U30514 (N_30514,N_28399,N_28251);
nor U30515 (N_30515,N_27764,N_29665);
xor U30516 (N_30516,N_27646,N_28268);
and U30517 (N_30517,N_28352,N_27698);
xor U30518 (N_30518,N_28790,N_28728);
nor U30519 (N_30519,N_29691,N_28243);
or U30520 (N_30520,N_27831,N_28801);
and U30521 (N_30521,N_27547,N_27889);
or U30522 (N_30522,N_29363,N_28377);
nand U30523 (N_30523,N_28219,N_27753);
nor U30524 (N_30524,N_27938,N_29280);
nor U30525 (N_30525,N_29721,N_28648);
or U30526 (N_30526,N_27954,N_28392);
or U30527 (N_30527,N_29616,N_29688);
nand U30528 (N_30528,N_27919,N_28229);
xnor U30529 (N_30529,N_28276,N_29174);
and U30530 (N_30530,N_28824,N_28237);
and U30531 (N_30531,N_28194,N_28021);
nor U30532 (N_30532,N_29635,N_29622);
or U30533 (N_30533,N_27825,N_28821);
nand U30534 (N_30534,N_27615,N_28627);
and U30535 (N_30535,N_28053,N_28837);
or U30536 (N_30536,N_28700,N_27839);
nand U30537 (N_30537,N_29013,N_27617);
or U30538 (N_30538,N_28166,N_28830);
nor U30539 (N_30539,N_29735,N_29815);
and U30540 (N_30540,N_29913,N_27513);
and U30541 (N_30541,N_29362,N_28134);
or U30542 (N_30542,N_28655,N_28630);
and U30543 (N_30543,N_29094,N_28539);
nor U30544 (N_30544,N_28098,N_28647);
xnor U30545 (N_30545,N_28925,N_28364);
or U30546 (N_30546,N_29081,N_28756);
and U30547 (N_30547,N_28218,N_27692);
xnor U30548 (N_30548,N_27928,N_28154);
or U30549 (N_30549,N_28671,N_27578);
xnor U30550 (N_30550,N_27626,N_29484);
or U30551 (N_30551,N_27911,N_28358);
nand U30552 (N_30552,N_28612,N_28111);
nand U30553 (N_30553,N_28263,N_29231);
nand U30554 (N_30554,N_29990,N_29742);
and U30555 (N_30555,N_28882,N_28575);
and U30556 (N_30556,N_28980,N_28508);
or U30557 (N_30557,N_29486,N_28469);
or U30558 (N_30558,N_29210,N_27709);
xnor U30559 (N_30559,N_29261,N_29016);
or U30560 (N_30560,N_28316,N_28407);
xor U30561 (N_30561,N_28269,N_29745);
xor U30562 (N_30562,N_28106,N_29628);
xor U30563 (N_30563,N_28825,N_28546);
or U30564 (N_30564,N_28155,N_29810);
xor U30565 (N_30565,N_28868,N_28754);
nor U30566 (N_30566,N_29047,N_28716);
nor U30567 (N_30567,N_28170,N_29630);
nand U30568 (N_30568,N_27645,N_27788);
xnor U30569 (N_30569,N_28453,N_29135);
and U30570 (N_30570,N_28623,N_29173);
and U30571 (N_30571,N_28045,N_28841);
or U30572 (N_30572,N_29748,N_29095);
nand U30573 (N_30573,N_28325,N_28650);
nand U30574 (N_30574,N_28211,N_28164);
nor U30575 (N_30575,N_29334,N_28278);
and U30576 (N_30576,N_27934,N_27886);
nand U30577 (N_30577,N_27752,N_28113);
nand U30578 (N_30578,N_28669,N_27960);
and U30579 (N_30579,N_29523,N_27618);
and U30580 (N_30580,N_27594,N_27833);
nand U30581 (N_30581,N_27555,N_27533);
nand U30582 (N_30582,N_29502,N_29140);
xor U30583 (N_30583,N_28936,N_27688);
nand U30584 (N_30584,N_28347,N_28995);
nor U30585 (N_30585,N_28012,N_29171);
or U30586 (N_30586,N_28301,N_28375);
and U30587 (N_30587,N_29874,N_29483);
or U30588 (N_30588,N_29710,N_28674);
nand U30589 (N_30589,N_28809,N_28808);
or U30590 (N_30590,N_28406,N_27730);
and U30591 (N_30591,N_29292,N_28160);
xnor U30592 (N_30592,N_29941,N_27826);
nor U30593 (N_30593,N_28466,N_29392);
nand U30594 (N_30594,N_28132,N_27959);
or U30595 (N_30595,N_29738,N_28439);
nand U30596 (N_30596,N_29925,N_29920);
and U30597 (N_30597,N_29603,N_29780);
nand U30598 (N_30598,N_29964,N_28232);
and U30599 (N_30599,N_28944,N_28758);
xnor U30600 (N_30600,N_27793,N_29329);
or U30601 (N_30601,N_29587,N_28070);
or U30602 (N_30602,N_28738,N_28540);
xnor U30603 (N_30603,N_29531,N_27610);
or U30604 (N_30604,N_29264,N_28872);
and U30605 (N_30605,N_27701,N_27669);
or U30606 (N_30606,N_28663,N_28536);
nor U30607 (N_30607,N_29891,N_29853);
nand U30608 (N_30608,N_28044,N_29681);
or U30609 (N_30609,N_29736,N_29855);
nand U30610 (N_30610,N_27956,N_29595);
nand U30611 (N_30611,N_29391,N_28592);
and U30612 (N_30612,N_27898,N_27964);
nand U30613 (N_30613,N_27993,N_28249);
and U30614 (N_30614,N_28773,N_28173);
nand U30615 (N_30615,N_29971,N_29849);
xor U30616 (N_30616,N_28395,N_29900);
xnor U30617 (N_30617,N_29327,N_28681);
and U30618 (N_30618,N_29518,N_28009);
and U30619 (N_30619,N_28085,N_29136);
or U30620 (N_30620,N_27576,N_29233);
or U30621 (N_30621,N_29755,N_28685);
and U30622 (N_30622,N_28690,N_29707);
and U30623 (N_30623,N_29605,N_29032);
nor U30624 (N_30624,N_28715,N_27902);
and U30625 (N_30625,N_28336,N_29620);
or U30626 (N_30626,N_28850,N_29169);
nand U30627 (N_30627,N_29538,N_29670);
or U30628 (N_30628,N_28432,N_27737);
or U30629 (N_30629,N_29369,N_29422);
or U30630 (N_30630,N_29965,N_27634);
nand U30631 (N_30631,N_28149,N_27732);
nor U30632 (N_30632,N_28483,N_29193);
xnor U30633 (N_30633,N_28144,N_27686);
nand U30634 (N_30634,N_29221,N_29325);
nor U30635 (N_30635,N_29025,N_27932);
xnor U30636 (N_30636,N_28367,N_28431);
and U30637 (N_30637,N_27981,N_29730);
nor U30638 (N_30638,N_29505,N_27957);
nor U30639 (N_30639,N_29888,N_29306);
nor U30640 (N_30640,N_29416,N_27789);
and U30641 (N_30641,N_28786,N_27908);
nand U30642 (N_30642,N_27521,N_29591);
nand U30643 (N_30643,N_28334,N_27652);
and U30644 (N_30644,N_27979,N_27596);
nand U30645 (N_30645,N_27903,N_29732);
and U30646 (N_30646,N_28139,N_28551);
xnor U30647 (N_30647,N_28953,N_27590);
or U30648 (N_30648,N_28497,N_28114);
xnor U30649 (N_30649,N_28420,N_27565);
or U30650 (N_30650,N_29625,N_27994);
or U30651 (N_30651,N_28635,N_28867);
and U30652 (N_30652,N_29901,N_28569);
xor U30653 (N_30653,N_27637,N_29559);
nor U30654 (N_30654,N_29859,N_28454);
xnor U30655 (N_30655,N_29895,N_28341);
xnor U30656 (N_30656,N_29993,N_29549);
or U30657 (N_30657,N_29520,N_29596);
and U30658 (N_30658,N_28314,N_29291);
nor U30659 (N_30659,N_29048,N_28491);
nor U30660 (N_30660,N_27534,N_28954);
nand U30661 (N_30661,N_29475,N_28158);
nor U30662 (N_30662,N_29311,N_28344);
xor U30663 (N_30663,N_28369,N_27921);
nand U30664 (N_30664,N_28446,N_29942);
xnor U30665 (N_30665,N_28729,N_27500);
nor U30666 (N_30666,N_27562,N_29578);
or U30667 (N_30667,N_27586,N_27700);
xnor U30668 (N_30668,N_28275,N_29003);
nor U30669 (N_30669,N_29744,N_29969);
and U30670 (N_30670,N_29879,N_27842);
xnor U30671 (N_30671,N_29458,N_29860);
xor U30672 (N_30672,N_29062,N_27925);
and U30673 (N_30673,N_28135,N_29513);
or U30674 (N_30674,N_29090,N_28782);
or U30675 (N_30675,N_27924,N_27922);
xnor U30676 (N_30676,N_28962,N_29727);
nor U30677 (N_30677,N_28236,N_29131);
nor U30678 (N_30678,N_28861,N_28562);
and U30679 (N_30679,N_29490,N_27822);
or U30680 (N_30680,N_28174,N_28596);
xor U30681 (N_30681,N_27524,N_28196);
and U30682 (N_30682,N_28414,N_28730);
xnor U30683 (N_30683,N_27508,N_27602);
nand U30684 (N_30684,N_28519,N_29851);
nand U30685 (N_30685,N_28235,N_29674);
or U30686 (N_30686,N_29469,N_27890);
nor U30687 (N_30687,N_28593,N_28445);
and U30688 (N_30688,N_29426,N_27517);
xor U30689 (N_30689,N_29015,N_28961);
nand U30690 (N_30690,N_28011,N_27877);
nand U30691 (N_30691,N_29420,N_29005);
xor U30692 (N_30692,N_29958,N_28485);
nor U30693 (N_30693,N_29797,N_29867);
and U30694 (N_30694,N_28346,N_28889);
nor U30695 (N_30695,N_28482,N_28999);
nand U30696 (N_30696,N_28620,N_28463);
nor U30697 (N_30697,N_28048,N_28920);
and U30698 (N_30698,N_28227,N_29075);
xor U30699 (N_30699,N_29352,N_28370);
nand U30700 (N_30700,N_28348,N_29301);
or U30701 (N_30701,N_28110,N_28127);
or U30702 (N_30702,N_28723,N_29276);
or U30703 (N_30703,N_29669,N_28709);
xnor U30704 (N_30704,N_29823,N_27580);
or U30705 (N_30705,N_29342,N_28927);
and U30706 (N_30706,N_28221,N_29979);
and U30707 (N_30707,N_29199,N_29762);
nor U30708 (N_30708,N_28888,N_28023);
nand U30709 (N_30709,N_28959,N_28579);
or U30710 (N_30710,N_28847,N_28644);
nand U30711 (N_30711,N_28610,N_29833);
and U30712 (N_30712,N_28660,N_29753);
and U30713 (N_30713,N_27942,N_27608);
nand U30714 (N_30714,N_27940,N_27591);
and U30715 (N_30715,N_28617,N_28613);
nor U30716 (N_30716,N_28964,N_29065);
and U30717 (N_30717,N_29408,N_27896);
xnor U30718 (N_30718,N_28842,N_29978);
nand U30719 (N_30719,N_27987,N_29495);
or U30720 (N_30720,N_29354,N_27965);
xnor U30721 (N_30721,N_27563,N_29072);
xnor U30722 (N_30722,N_28913,N_28570);
nor U30723 (N_30723,N_28915,N_29427);
xor U30724 (N_30724,N_29021,N_28529);
and U30725 (N_30725,N_28217,N_29963);
nor U30726 (N_30726,N_29466,N_29328);
or U30727 (N_30727,N_29643,N_28561);
xnor U30728 (N_30728,N_28333,N_28548);
xnor U30729 (N_30729,N_29574,N_27641);
and U30730 (N_30730,N_29441,N_27548);
or U30731 (N_30731,N_27592,N_28212);
and U30732 (N_30732,N_28717,N_28712);
nand U30733 (N_30733,N_28791,N_28036);
nor U30734 (N_30734,N_28526,N_28885);
and U30735 (N_30735,N_29395,N_29514);
nor U30736 (N_30736,N_28311,N_29116);
nand U30737 (N_30737,N_29141,N_29789);
or U30738 (N_30738,N_27963,N_29424);
and U30739 (N_30739,N_28228,N_27866);
and U30740 (N_30740,N_29460,N_27978);
xor U30741 (N_30741,N_27632,N_28854);
xnor U30742 (N_30742,N_28565,N_28427);
and U30743 (N_30743,N_28429,N_27716);
nor U30744 (N_30744,N_27560,N_28246);
xnor U30745 (N_30745,N_28072,N_29238);
or U30746 (N_30746,N_28354,N_28289);
and U30747 (N_30747,N_27647,N_28945);
nor U30748 (N_30748,N_29675,N_28862);
nor U30749 (N_30749,N_29737,N_28658);
or U30750 (N_30750,N_28972,N_28794);
xor U30751 (N_30751,N_28811,N_29412);
xnor U30752 (N_30752,N_27639,N_29594);
nor U30753 (N_30753,N_29646,N_28506);
or U30754 (N_30754,N_28068,N_29159);
nand U30755 (N_30755,N_28736,N_28597);
or U30756 (N_30756,N_28528,N_28628);
nor U30757 (N_30757,N_27923,N_29251);
nor U30758 (N_30758,N_29694,N_27506);
nor U30759 (N_30759,N_29281,N_27870);
or U30760 (N_30760,N_27736,N_28208);
nand U30761 (N_30761,N_27554,N_28425);
nor U30762 (N_30762,N_29445,N_28576);
and U30763 (N_30763,N_28721,N_28416);
xor U30764 (N_30764,N_27650,N_29634);
or U30765 (N_30765,N_28815,N_28337);
or U30766 (N_30766,N_27967,N_29718);
and U30767 (N_30767,N_29401,N_28938);
nor U30768 (N_30768,N_28447,N_27891);
and U30769 (N_30769,N_28080,N_29297);
xnor U30770 (N_30770,N_29794,N_29053);
xnor U30771 (N_30771,N_27871,N_29967);
or U30772 (N_30772,N_29228,N_29184);
xor U30773 (N_30773,N_28285,N_29330);
and U30774 (N_30774,N_29611,N_28294);
nand U30775 (N_30775,N_29019,N_28505);
xnor U30776 (N_30776,N_29045,N_28107);
nor U30777 (N_30777,N_28267,N_29618);
nand U30778 (N_30778,N_29722,N_29303);
xor U30779 (N_30779,N_27969,N_27660);
or U30780 (N_30780,N_27541,N_28522);
nand U30781 (N_30781,N_28904,N_27733);
nand U30782 (N_30782,N_27531,N_28258);
xor U30783 (N_30783,N_29245,N_28784);
and U30784 (N_30784,N_29026,N_29533);
xor U30785 (N_30785,N_28191,N_28371);
nor U30786 (N_30786,N_29719,N_29728);
xnor U30787 (N_30787,N_27510,N_28751);
or U30788 (N_30788,N_28625,N_29844);
and U30789 (N_30789,N_28093,N_28993);
nor U30790 (N_30790,N_27542,N_29471);
and U30791 (N_30791,N_27897,N_28857);
or U30792 (N_30792,N_28378,N_28515);
nand U30793 (N_30793,N_28557,N_29087);
nand U30794 (N_30794,N_29444,N_27574);
xor U30795 (N_30795,N_27665,N_29107);
or U30796 (N_30796,N_27687,N_29909);
nor U30797 (N_30797,N_27683,N_27984);
and U30798 (N_30798,N_28844,N_27819);
and U30799 (N_30799,N_28687,N_27806);
xor U30800 (N_30800,N_29840,N_27918);
or U30801 (N_30801,N_28555,N_29142);
nand U30802 (N_30802,N_29319,N_27794);
or U30803 (N_30803,N_29355,N_28320);
or U30804 (N_30804,N_29462,N_27523);
xnor U30805 (N_30805,N_28694,N_28206);
nor U30806 (N_30806,N_29204,N_28123);
nor U30807 (N_30807,N_29769,N_28852);
or U30808 (N_30808,N_29359,N_28991);
xnor U30809 (N_30809,N_28086,N_28818);
xor U30810 (N_30810,N_29447,N_28057);
and U30811 (N_30811,N_29104,N_28678);
and U30812 (N_30812,N_29671,N_28213);
nor U30813 (N_30813,N_28298,N_29243);
nand U30814 (N_30814,N_29270,N_29649);
xor U30815 (N_30815,N_29998,N_28839);
or U30816 (N_30816,N_27772,N_28203);
and U30817 (N_30817,N_29834,N_29491);
or U30818 (N_30818,N_28075,N_28934);
xor U30819 (N_30819,N_29340,N_28656);
nor U30820 (N_30820,N_28188,N_28804);
and U30821 (N_30821,N_29406,N_29207);
and U30822 (N_30822,N_29387,N_29368);
nand U30823 (N_30823,N_27828,N_27756);
and U30824 (N_30824,N_27778,N_28073);
and U30825 (N_30825,N_29689,N_28064);
or U30826 (N_30826,N_27710,N_28645);
nor U30827 (N_30827,N_29250,N_29524);
or U30828 (N_30828,N_29904,N_29237);
and U30829 (N_30829,N_28670,N_28822);
xor U30830 (N_30830,N_28338,N_29952);
xnor U30831 (N_30831,N_28618,N_28843);
nor U30832 (N_30832,N_29786,N_27933);
or U30833 (N_30833,N_29526,N_28750);
and U30834 (N_30834,N_29287,N_29418);
or U30835 (N_30835,N_28118,N_29656);
nor U30836 (N_30836,N_29550,N_27734);
nor U30837 (N_30837,N_28734,N_27629);
nand U30838 (N_30838,N_28525,N_29461);
xnor U30839 (N_30839,N_27781,N_28636);
xor U30840 (N_30840,N_28304,N_27749);
or U30841 (N_30841,N_28859,N_29374);
xnor U30842 (N_30842,N_29487,N_28430);
xor U30843 (N_30843,N_28029,N_27588);
nand U30844 (N_30844,N_29957,N_29838);
nand U30845 (N_30845,N_28264,N_29113);
xnor U30846 (N_30846,N_29884,N_28833);
nand U30847 (N_30847,N_28523,N_27566);
nor U30848 (N_30848,N_29247,N_28245);
and U30849 (N_30849,N_29782,N_29617);
and U30850 (N_30850,N_28262,N_29098);
and U30851 (N_30851,N_28550,N_29652);
nor U30852 (N_30852,N_27573,N_27661);
or U30853 (N_30853,N_28484,N_29887);
xnor U30854 (N_30854,N_28488,N_28955);
nor U30855 (N_30855,N_29229,N_27915);
nand U30856 (N_30856,N_29878,N_28975);
or U30857 (N_30857,N_27895,N_28286);
and U30858 (N_30858,N_29373,N_28937);
and U30859 (N_30859,N_29683,N_29610);
nor U30860 (N_30860,N_28554,N_29052);
nor U30861 (N_30861,N_27723,N_28076);
nor U30862 (N_30862,N_29556,N_29489);
or U30863 (N_30863,N_29804,N_28313);
xor U30864 (N_30864,N_29450,N_27854);
or U30865 (N_30865,N_29118,N_27980);
or U30866 (N_30866,N_29837,N_29693);
and U30867 (N_30867,N_29271,N_28587);
nand U30868 (N_30868,N_29644,N_29256);
xnor U30869 (N_30869,N_29110,N_28973);
nand U30870 (N_30870,N_29105,N_28284);
nor U30871 (N_30871,N_28547,N_28869);
xnor U30872 (N_30872,N_29192,N_27843);
nor U30873 (N_30873,N_27976,N_28104);
or U30874 (N_30874,N_29944,N_28543);
nand U30875 (N_30875,N_29219,N_27505);
or U30876 (N_30876,N_28248,N_29589);
and U30877 (N_30877,N_28922,N_28558);
xnor U30878 (N_30878,N_28039,N_28881);
nor U30879 (N_30879,N_28162,N_28224);
nor U30880 (N_30880,N_27649,N_27638);
nor U30881 (N_30881,N_29604,N_29704);
nor U30882 (N_30882,N_28389,N_28189);
nor U30883 (N_30883,N_29063,N_28848);
and U30884 (N_30884,N_29734,N_29182);
nand U30885 (N_30885,N_27556,N_28421);
and U30886 (N_30886,N_27827,N_29024);
and U30887 (N_30887,N_28680,N_28026);
nor U30888 (N_30888,N_28200,N_28234);
nand U30889 (N_30889,N_27507,N_28499);
or U30890 (N_30890,N_29927,N_28893);
and U30891 (N_30891,N_27892,N_29648);
or U30892 (N_30892,N_28402,N_27614);
or U30893 (N_30893,N_29659,N_29516);
nor U30894 (N_30894,N_27509,N_29515);
or U30895 (N_30895,N_29121,N_28797);
or U30896 (N_30896,N_29023,N_28892);
or U30897 (N_30897,N_29597,N_29807);
nor U30898 (N_30898,N_28785,N_29935);
or U30899 (N_30899,N_28146,N_29724);
nor U30900 (N_30900,N_29304,N_27743);
nand U30901 (N_30901,N_27570,N_29123);
nand U30902 (N_30902,N_28168,N_29551);
xnor U30903 (N_30903,N_28689,N_29077);
and U30904 (N_30904,N_28355,N_28153);
or U30905 (N_30905,N_29155,N_29905);
and U30906 (N_30906,N_29642,N_28084);
and U30907 (N_30907,N_29633,N_29027);
and U30908 (N_30908,N_28418,N_29187);
and U30909 (N_30909,N_28282,N_29638);
nand U30910 (N_30910,N_29557,N_27604);
nand U30911 (N_30911,N_28152,N_29968);
xor U30912 (N_30912,N_27653,N_29386);
or U30913 (N_30913,N_28697,N_29989);
nor U30914 (N_30914,N_28553,N_27996);
nand U30915 (N_30915,N_28233,N_29030);
nor U30916 (N_30916,N_29729,N_28935);
and U30917 (N_30917,N_29761,N_28477);
or U30918 (N_30918,N_29757,N_28932);
xor U30919 (N_30919,N_28718,N_28622);
xor U30920 (N_30920,N_27623,N_29056);
or U30921 (N_30921,N_29535,N_27515);
nand U30922 (N_30922,N_29345,N_29212);
or U30923 (N_30923,N_28324,N_28436);
and U30924 (N_30924,N_29055,N_28883);
and U30925 (N_30925,N_28361,N_27952);
xor U30926 (N_30926,N_28396,N_27759);
or U30927 (N_30927,N_29839,N_28573);
and U30928 (N_30928,N_29702,N_29033);
xnor U30929 (N_30929,N_28353,N_28031);
or U30930 (N_30930,N_28410,N_29485);
nand U30931 (N_30931,N_28307,N_29530);
xnor U30932 (N_30932,N_28832,N_27706);
nor U30933 (N_30933,N_29290,N_29456);
nor U30934 (N_30934,N_28763,N_29446);
nor U30935 (N_30935,N_29274,N_28271);
and U30936 (N_30936,N_27771,N_29049);
xor U30937 (N_30937,N_29561,N_28303);
and U30938 (N_30938,N_29440,N_29453);
xor U30939 (N_30939,N_28016,N_29230);
xnor U30940 (N_30940,N_28253,N_28137);
nor U30941 (N_30941,N_29242,N_28117);
nor U30942 (N_30942,N_28398,N_28487);
xnor U30943 (N_30943,N_29130,N_29145);
nor U30944 (N_30944,N_27845,N_29818);
xnor U30945 (N_30945,N_28566,N_27804);
xnor U30946 (N_30946,N_29812,N_27664);
xor U30947 (N_30947,N_29846,N_27949);
nand U30948 (N_30948,N_29253,N_29593);
or U30949 (N_30949,N_28895,N_29773);
nor U30950 (N_30950,N_28997,N_29346);
and U30951 (N_30951,N_28498,N_27853);
xor U30952 (N_30952,N_28270,N_28860);
or U30953 (N_30953,N_28471,N_28702);
nand U30954 (N_30954,N_28143,N_29341);
or U30955 (N_30955,N_27558,N_28507);
xor U30956 (N_30956,N_27544,N_28247);
and U30957 (N_30957,N_27738,N_27747);
and U30958 (N_30958,N_27792,N_29436);
xor U30959 (N_30959,N_29973,N_27613);
or U30960 (N_30960,N_28981,N_28130);
xor U30961 (N_30961,N_29122,N_28767);
nand U30962 (N_30962,N_29282,N_27770);
nor U30963 (N_30963,N_28265,N_29831);
and U30964 (N_30964,N_28101,N_29409);
and U30965 (N_30965,N_29897,N_27676);
nor U30966 (N_30966,N_28397,N_28609);
nor U30967 (N_30967,N_29035,N_27719);
nand U30968 (N_30968,N_27728,N_29402);
nand U30969 (N_30969,N_29673,N_27971);
and U30970 (N_30970,N_27751,N_28556);
nor U30971 (N_30971,N_28802,N_28148);
and U30972 (N_30972,N_27851,N_29494);
or U30973 (N_30973,N_28746,N_28342);
nor U30974 (N_30974,N_28870,N_29010);
nand U30975 (N_30975,N_29215,N_29146);
nor U30976 (N_30976,N_27859,N_29157);
or U30977 (N_30977,N_28063,N_28428);
nand U30978 (N_30978,N_29493,N_28533);
and U30979 (N_30979,N_28295,N_29708);
xor U30980 (N_30980,N_29987,N_29039);
xnor U30981 (N_30981,N_29308,N_29808);
xor U30982 (N_30982,N_28600,N_29008);
and U30983 (N_30983,N_29541,N_28034);
and U30984 (N_30984,N_28616,N_28260);
and U30985 (N_30985,N_29321,N_29111);
nand U30986 (N_30986,N_29470,N_28912);
nor U30987 (N_30987,N_28133,N_29598);
xnor U30988 (N_30988,N_27684,N_28909);
nand U30989 (N_30989,N_29189,N_27787);
and U30990 (N_30990,N_28027,N_29599);
and U30991 (N_30991,N_28787,N_29022);
or U30992 (N_30992,N_27947,N_28781);
and U30993 (N_30993,N_29700,N_29828);
xnor U30994 (N_30994,N_29370,N_28190);
and U30995 (N_30995,N_28388,N_29074);
and U30996 (N_30996,N_29580,N_29467);
nand U30997 (N_30997,N_27986,N_27832);
nand U30998 (N_30998,N_29799,N_28930);
nor U30999 (N_30999,N_29956,N_29714);
xnor U31000 (N_31000,N_27791,N_28933);
nand U31001 (N_31001,N_29554,N_27543);
xnor U31002 (N_31002,N_27703,N_29692);
nor U31003 (N_31003,N_27953,N_28907);
and U31004 (N_31004,N_27760,N_29752);
nand U31005 (N_31005,N_29331,N_28994);
nand U31006 (N_31006,N_29563,N_29315);
and U31007 (N_31007,N_27852,N_29448);
or U31008 (N_31008,N_28875,N_28887);
nand U31009 (N_31009,N_29613,N_28183);
xnor U31010 (N_31010,N_29257,N_29099);
and U31011 (N_31011,N_29318,N_29894);
nand U31012 (N_31012,N_28761,N_28607);
and U31013 (N_31013,N_29497,N_27689);
nand U31014 (N_31014,N_29910,N_28214);
or U31015 (N_31015,N_29785,N_29361);
nand U31016 (N_31016,N_29162,N_27795);
or U31017 (N_31017,N_29302,N_28391);
nand U31018 (N_31018,N_29432,N_27612);
xnor U31019 (N_31019,N_29108,N_28714);
xor U31020 (N_31020,N_29128,N_28082);
nand U31021 (N_31021,N_27944,N_29492);
xnor U31022 (N_31022,N_27863,N_29585);
or U31023 (N_31023,N_27714,N_29911);
nor U31024 (N_31024,N_28087,N_28590);
xor U31025 (N_31025,N_28978,N_27616);
or U31026 (N_31026,N_29129,N_28880);
nor U31027 (N_31027,N_28583,N_29112);
xor U31028 (N_31028,N_29205,N_29918);
and U31029 (N_31029,N_29411,N_29449);
nand U31030 (N_31030,N_29723,N_29607);
nor U31031 (N_31031,N_29501,N_28475);
nand U31032 (N_31032,N_27550,N_28332);
or U31033 (N_31033,N_28900,N_29002);
and U31034 (N_31034,N_29805,N_29803);
xnor U31035 (N_31035,N_28290,N_28178);
and U31036 (N_31036,N_29413,N_28197);
xor U31037 (N_31037,N_28928,N_28501);
or U31038 (N_31038,N_28766,N_29218);
or U31039 (N_31039,N_28381,N_28724);
xor U31040 (N_31040,N_29668,N_27691);
xnor U31041 (N_31041,N_27758,N_28899);
nor U31042 (N_31042,N_29856,N_28479);
xor U31043 (N_31043,N_28465,N_28757);
nand U31044 (N_31044,N_28733,N_29503);
or U31045 (N_31045,N_28743,N_29880);
and U31046 (N_31046,N_29265,N_29889);
and U31047 (N_31047,N_29208,N_27790);
nor U31048 (N_31048,N_28386,N_28800);
nor U31049 (N_31049,N_28231,N_28725);
xor U31050 (N_31050,N_28105,N_29186);
nor U31051 (N_31051,N_28254,N_29103);
or U31052 (N_31052,N_28459,N_28705);
and U31053 (N_31053,N_27605,N_28356);
nor U31054 (N_31054,N_28744,N_28472);
nand U31055 (N_31055,N_29038,N_29384);
or U31056 (N_31056,N_29903,N_27946);
nor U31057 (N_31057,N_28722,N_28807);
nand U31058 (N_31058,N_29166,N_28205);
nor U31059 (N_31059,N_27557,N_29239);
xor U31060 (N_31060,N_29740,N_28457);
and U31061 (N_31061,N_27679,N_28657);
or U31062 (N_31062,N_29629,N_27640);
xnor U31063 (N_31063,N_29073,N_29295);
nand U31064 (N_31064,N_27884,N_28764);
xnor U31065 (N_31065,N_29624,N_28710);
nor U31066 (N_31066,N_29164,N_27931);
nor U31067 (N_31067,N_29677,N_29463);
nor U31068 (N_31068,N_27635,N_27929);
or U31069 (N_31069,N_29305,N_28732);
and U31070 (N_31070,N_28384,N_27631);
xnor U31071 (N_31071,N_29429,N_28960);
nand U31072 (N_31072,N_28222,N_27999);
or U31073 (N_31073,N_28737,N_29584);
and U31074 (N_31074,N_28077,N_28753);
nand U31075 (N_31075,N_29054,N_27529);
or U31076 (N_31076,N_27722,N_29036);
and U31077 (N_31077,N_28013,N_28708);
or U31078 (N_31078,N_29375,N_28699);
nor U31079 (N_31079,N_28167,N_28917);
nand U31080 (N_31080,N_29657,N_28201);
or U31081 (N_31081,N_28950,N_28982);
and U31082 (N_31082,N_28516,N_28969);
and U31083 (N_31083,N_28783,N_29152);
nor U31084 (N_31084,N_29609,N_29476);
xnor U31085 (N_31085,N_29109,N_29377);
and U31086 (N_31086,N_29011,N_29004);
and U31087 (N_31087,N_29358,N_28256);
or U31088 (N_31088,N_28083,N_27835);
or U31089 (N_31089,N_29937,N_29875);
nor U31090 (N_31090,N_29666,N_28319);
and U31091 (N_31091,N_29263,N_28096);
nor U31092 (N_31092,N_29254,N_28634);
and U31093 (N_31093,N_29244,N_28589);
nor U31094 (N_31094,N_29600,N_28977);
nor U31095 (N_31095,N_28171,N_27673);
nand U31096 (N_31096,N_29102,N_29459);
nor U31097 (N_31097,N_28305,N_29885);
or U31098 (N_31098,N_28527,N_27504);
nor U31099 (N_31099,N_28586,N_29273);
xor U31100 (N_31100,N_27800,N_27817);
nor U31101 (N_31101,N_29801,N_27941);
and U31102 (N_31102,N_29974,N_29826);
nor U31103 (N_31103,N_29326,N_29430);
or U31104 (N_31104,N_27872,N_29835);
xnor U31105 (N_31105,N_29760,N_29614);
and U31106 (N_31106,N_27530,N_28339);
and U31107 (N_31107,N_29398,N_29404);
nand U31108 (N_31108,N_27820,N_27848);
xnor U31109 (N_31109,N_27622,N_28520);
nor U31110 (N_31110,N_27742,N_28225);
nand U31111 (N_31111,N_27860,N_28380);
xnor U31112 (N_31112,N_27913,N_29612);
or U31113 (N_31113,N_29795,N_28611);
and U31114 (N_31114,N_29046,N_28796);
nor U31115 (N_31115,N_29608,N_28120);
and U31116 (N_31116,N_27814,N_29260);
xnor U31117 (N_31117,N_27577,N_27841);
xor U31118 (N_31118,N_28193,N_27844);
nor U31119 (N_31119,N_29161,N_28489);
or U31120 (N_31120,N_28504,N_27955);
nor U31121 (N_31121,N_27802,N_29012);
and U31122 (N_31122,N_29266,N_27883);
and U31123 (N_31123,N_28417,N_27611);
or U31124 (N_31124,N_29899,N_29854);
nand U31125 (N_31125,N_28215,N_29209);
and U31126 (N_31126,N_29034,N_28000);
nor U31127 (N_31127,N_29097,N_29892);
xnor U31128 (N_31128,N_28056,N_27748);
nand U31129 (N_31129,N_29820,N_29001);
and U31130 (N_31130,N_28643,N_27937);
nand U31131 (N_31131,N_28856,N_29534);
or U31132 (N_31132,N_27970,N_29379);
nor U31133 (N_31133,N_28310,N_27552);
nand U31134 (N_31134,N_29712,N_29050);
and U31135 (N_31135,N_29824,N_28510);
xnor U31136 (N_31136,N_29562,N_29443);
and U31137 (N_31137,N_27875,N_28770);
or U31138 (N_31138,N_28293,N_27654);
nand U31139 (N_31139,N_29317,N_28580);
xnor U31140 (N_31140,N_29279,N_29043);
nand U31141 (N_31141,N_29924,N_27951);
xnor U31142 (N_31142,N_28125,N_27532);
nor U31143 (N_31143,N_29936,N_29592);
nor U31144 (N_31144,N_29227,N_29947);
nand U31145 (N_31145,N_27888,N_28103);
xor U31146 (N_31146,N_28065,N_29962);
xor U31147 (N_31147,N_27725,N_27675);
nor U31148 (N_31148,N_28461,N_28092);
nand U31149 (N_31149,N_28896,N_28345);
xnor U31150 (N_31150,N_28594,N_29371);
or U31151 (N_31151,N_28878,N_28654);
nand U31152 (N_31152,N_29091,N_29809);
nor U31153 (N_31153,N_27619,N_29542);
or U31154 (N_31154,N_28827,N_27873);
xor U31155 (N_31155,N_27511,N_29085);
nor U31156 (N_31156,N_28244,N_29573);
and U31157 (N_31157,N_28545,N_28321);
or U31158 (N_31158,N_28448,N_29565);
nor U31159 (N_31159,N_29747,N_28041);
nor U31160 (N_31160,N_29410,N_28639);
and U31161 (N_31161,N_29029,N_28335);
nor U31162 (N_31162,N_29455,N_29236);
xor U31163 (N_31163,N_28343,N_28838);
nor U31164 (N_31164,N_29626,N_29663);
nand U31165 (N_31165,N_27644,N_29454);
nor U31166 (N_31166,N_27861,N_28598);
nand U31167 (N_31167,N_28914,N_28632);
nand U31168 (N_31168,N_27864,N_28642);
nand U31169 (N_31169,N_29658,N_28902);
xor U31170 (N_31170,N_29144,N_27834);
nand U31171 (N_31171,N_29252,N_28891);
and U31172 (N_31172,N_27773,N_29678);
xnor U31173 (N_31173,N_29931,N_29433);
and U31174 (N_31174,N_28069,N_28563);
nor U31175 (N_31175,N_29414,N_29781);
and U31176 (N_31176,N_29754,N_29403);
xor U31177 (N_31177,N_28049,N_27595);
nand U31178 (N_31178,N_28696,N_27910);
or U31179 (N_31179,N_29040,N_29715);
and U31180 (N_31180,N_27990,N_28748);
nand U31181 (N_31181,N_27975,N_29588);
or U31182 (N_31182,N_29258,N_29126);
xnor U31183 (N_31183,N_28308,N_28423);
and U31184 (N_31184,N_27718,N_29830);
xor U31185 (N_31185,N_28008,N_29194);
nor U31186 (N_31186,N_29324,N_29425);
xnor U31187 (N_31187,N_28752,N_29850);
or U31188 (N_31188,N_28866,N_27799);
and U31189 (N_31189,N_29881,N_29498);
nand U31190 (N_31190,N_29653,N_28626);
or U31191 (N_31191,N_28180,N_29343);
nor U31192 (N_31192,N_28776,N_29572);
xnor U31193 (N_31193,N_29093,N_28413);
xor U31194 (N_31194,N_28855,N_28359);
and U31195 (N_31195,N_28387,N_28081);
and U31196 (N_31196,N_27974,N_28116);
nor U31197 (N_31197,N_29902,N_29275);
nand U31198 (N_31198,N_27671,N_29647);
nor U31199 (N_31199,N_29299,N_29147);
or U31200 (N_31200,N_28467,N_28408);
nor U31201 (N_31201,N_27699,N_27768);
nor U31202 (N_31202,N_29213,N_27702);
nor U31203 (N_31203,N_27597,N_27643);
and U31204 (N_31204,N_28115,N_28614);
or U31205 (N_31205,N_28480,N_27972);
nand U31206 (N_31206,N_29510,N_27985);
nor U31207 (N_31207,N_29320,N_28198);
nand U31208 (N_31208,N_29439,N_28434);
nand U31209 (N_31209,N_29376,N_29383);
and U31210 (N_31210,N_29976,N_29695);
and U31211 (N_31211,N_29017,N_29886);
nor U31212 (N_31212,N_27797,N_29051);
nand U31213 (N_31213,N_29117,N_28890);
nor U31214 (N_31214,N_28948,N_27805);
or U31215 (N_31215,N_27540,N_28921);
xnor U31216 (N_31216,N_29917,N_29836);
or U31217 (N_31217,N_29992,N_27968);
and U31218 (N_31218,N_29751,N_28514);
nand U31219 (N_31219,N_28451,N_28532);
or U31220 (N_31220,N_28327,N_28140);
xor U31221 (N_31221,N_27989,N_29601);
nor U31222 (N_31222,N_27838,N_29289);
nor U31223 (N_31223,N_28199,N_29890);
or U31224 (N_31224,N_27693,N_29397);
xor U31225 (N_31225,N_29217,N_29870);
and U31226 (N_31226,N_29482,N_27582);
or U31227 (N_31227,N_29176,N_28772);
and U31228 (N_31228,N_29240,N_27905);
nand U31229 (N_31229,N_28923,N_28317);
and U31230 (N_31230,N_28810,N_27735);
and U31231 (N_31231,N_28916,N_29566);
nand U31232 (N_31232,N_28328,N_28779);
nand U31233 (N_31233,N_27551,N_27633);
nand U31234 (N_31234,N_27809,N_28765);
xnor U31235 (N_31235,N_27783,N_27520);
xnor U31236 (N_31236,N_29066,N_29945);
nand U31237 (N_31237,N_28778,N_28901);
xor U31238 (N_31238,N_27766,N_29499);
nand U31239 (N_31239,N_27801,N_28490);
xnor U31240 (N_31240,N_28755,N_29819);
nand U31241 (N_31241,N_27926,N_29132);
nor U31242 (N_31242,N_27674,N_28667);
nor U31243 (N_31243,N_28560,N_28672);
and U31244 (N_31244,N_28552,N_27836);
nand U31245 (N_31245,N_28996,N_29627);
xnor U31246 (N_31246,N_28524,N_28058);
or U31247 (N_31247,N_27784,N_28022);
and U31248 (N_31248,N_29479,N_29521);
and U31249 (N_31249,N_29916,N_27879);
nand U31250 (N_31250,N_28567,N_28712);
nand U31251 (N_31251,N_29663,N_29143);
and U31252 (N_31252,N_28259,N_29974);
nand U31253 (N_31253,N_28215,N_28692);
nand U31254 (N_31254,N_29421,N_29794);
and U31255 (N_31255,N_29264,N_29312);
or U31256 (N_31256,N_28773,N_28553);
nor U31257 (N_31257,N_29507,N_27579);
and U31258 (N_31258,N_29610,N_29072);
and U31259 (N_31259,N_28380,N_29639);
nor U31260 (N_31260,N_29620,N_27689);
nand U31261 (N_31261,N_29918,N_28249);
nand U31262 (N_31262,N_28639,N_28121);
xnor U31263 (N_31263,N_29371,N_29165);
or U31264 (N_31264,N_27615,N_29517);
or U31265 (N_31265,N_28299,N_29978);
xnor U31266 (N_31266,N_29895,N_28400);
xor U31267 (N_31267,N_29733,N_29268);
nor U31268 (N_31268,N_28722,N_28284);
or U31269 (N_31269,N_28238,N_28969);
or U31270 (N_31270,N_29176,N_28692);
xnor U31271 (N_31271,N_27552,N_28108);
and U31272 (N_31272,N_27532,N_27538);
xor U31273 (N_31273,N_28716,N_28657);
or U31274 (N_31274,N_28005,N_28897);
nand U31275 (N_31275,N_29552,N_28371);
xnor U31276 (N_31276,N_28150,N_29554);
or U31277 (N_31277,N_29232,N_28514);
nand U31278 (N_31278,N_27784,N_28842);
or U31279 (N_31279,N_28828,N_29727);
and U31280 (N_31280,N_29798,N_27930);
nand U31281 (N_31281,N_29880,N_27849);
nor U31282 (N_31282,N_28040,N_29167);
nand U31283 (N_31283,N_28395,N_27643);
nand U31284 (N_31284,N_29923,N_28782);
and U31285 (N_31285,N_28449,N_28267);
and U31286 (N_31286,N_27902,N_28881);
nand U31287 (N_31287,N_29826,N_27847);
xor U31288 (N_31288,N_28806,N_29099);
nand U31289 (N_31289,N_28582,N_28474);
nor U31290 (N_31290,N_28114,N_28449);
xnor U31291 (N_31291,N_27889,N_29069);
or U31292 (N_31292,N_27666,N_27758);
xor U31293 (N_31293,N_29670,N_27551);
and U31294 (N_31294,N_27987,N_28144);
nor U31295 (N_31295,N_29610,N_29116);
nor U31296 (N_31296,N_29857,N_28643);
nor U31297 (N_31297,N_29052,N_28105);
nor U31298 (N_31298,N_28533,N_28960);
or U31299 (N_31299,N_29184,N_28747);
or U31300 (N_31300,N_28677,N_28012);
or U31301 (N_31301,N_29726,N_27761);
nor U31302 (N_31302,N_29657,N_27825);
and U31303 (N_31303,N_28955,N_29337);
xor U31304 (N_31304,N_29721,N_28678);
nand U31305 (N_31305,N_28904,N_28115);
xnor U31306 (N_31306,N_27845,N_29739);
xor U31307 (N_31307,N_29307,N_29353);
and U31308 (N_31308,N_28151,N_29074);
xnor U31309 (N_31309,N_28761,N_29333);
nand U31310 (N_31310,N_29788,N_29993);
xor U31311 (N_31311,N_29419,N_29294);
nor U31312 (N_31312,N_27698,N_28846);
nand U31313 (N_31313,N_28732,N_28527);
xnor U31314 (N_31314,N_28912,N_28032);
xor U31315 (N_31315,N_28276,N_29496);
xor U31316 (N_31316,N_29745,N_29413);
xor U31317 (N_31317,N_27945,N_28756);
nand U31318 (N_31318,N_28052,N_27765);
xor U31319 (N_31319,N_27955,N_28008);
nor U31320 (N_31320,N_27909,N_28266);
or U31321 (N_31321,N_27971,N_29318);
and U31322 (N_31322,N_28856,N_29592);
and U31323 (N_31323,N_27543,N_27717);
nand U31324 (N_31324,N_28629,N_28133);
nor U31325 (N_31325,N_29666,N_29053);
or U31326 (N_31326,N_27940,N_28949);
nand U31327 (N_31327,N_28427,N_29048);
nor U31328 (N_31328,N_27732,N_28109);
xor U31329 (N_31329,N_28470,N_29714);
xnor U31330 (N_31330,N_29830,N_29763);
nor U31331 (N_31331,N_28185,N_29736);
nand U31332 (N_31332,N_29313,N_28252);
xnor U31333 (N_31333,N_28960,N_28695);
and U31334 (N_31334,N_29232,N_29394);
nor U31335 (N_31335,N_28796,N_28205);
or U31336 (N_31336,N_27974,N_29856);
nor U31337 (N_31337,N_29946,N_29103);
nand U31338 (N_31338,N_28546,N_27553);
nor U31339 (N_31339,N_29945,N_28962);
xor U31340 (N_31340,N_29293,N_29879);
nand U31341 (N_31341,N_28546,N_28909);
or U31342 (N_31342,N_27917,N_28863);
nor U31343 (N_31343,N_29735,N_27751);
nor U31344 (N_31344,N_27712,N_27909);
nand U31345 (N_31345,N_27931,N_27506);
xnor U31346 (N_31346,N_28927,N_27762);
nand U31347 (N_31347,N_29074,N_29121);
and U31348 (N_31348,N_28363,N_29340);
or U31349 (N_31349,N_29903,N_29728);
or U31350 (N_31350,N_28474,N_27658);
xnor U31351 (N_31351,N_29068,N_28328);
or U31352 (N_31352,N_27519,N_29332);
or U31353 (N_31353,N_28639,N_27681);
nor U31354 (N_31354,N_28013,N_27835);
or U31355 (N_31355,N_28919,N_29836);
xnor U31356 (N_31356,N_28703,N_28663);
nand U31357 (N_31357,N_28496,N_27957);
xnor U31358 (N_31358,N_28346,N_29657);
and U31359 (N_31359,N_29640,N_28452);
xor U31360 (N_31360,N_28543,N_28385);
nand U31361 (N_31361,N_28962,N_28803);
or U31362 (N_31362,N_28659,N_27540);
nor U31363 (N_31363,N_29699,N_29062);
and U31364 (N_31364,N_28440,N_28653);
or U31365 (N_31365,N_28222,N_29468);
or U31366 (N_31366,N_29117,N_28723);
and U31367 (N_31367,N_27574,N_28587);
xnor U31368 (N_31368,N_29157,N_27788);
or U31369 (N_31369,N_29395,N_28585);
nand U31370 (N_31370,N_28704,N_28337);
xor U31371 (N_31371,N_27749,N_29497);
or U31372 (N_31372,N_28859,N_29420);
nor U31373 (N_31373,N_27776,N_29239);
and U31374 (N_31374,N_29064,N_28725);
nor U31375 (N_31375,N_28091,N_28306);
and U31376 (N_31376,N_28084,N_28692);
and U31377 (N_31377,N_27739,N_29093);
nor U31378 (N_31378,N_27812,N_28942);
or U31379 (N_31379,N_28678,N_29280);
and U31380 (N_31380,N_29558,N_28906);
nand U31381 (N_31381,N_29505,N_29515);
or U31382 (N_31382,N_28853,N_27797);
xnor U31383 (N_31383,N_28565,N_28860);
nor U31384 (N_31384,N_28718,N_28448);
nand U31385 (N_31385,N_29399,N_27742);
nor U31386 (N_31386,N_29539,N_28002);
xnor U31387 (N_31387,N_28599,N_28030);
and U31388 (N_31388,N_28297,N_29304);
xor U31389 (N_31389,N_28775,N_29780);
nand U31390 (N_31390,N_28394,N_28811);
nand U31391 (N_31391,N_29155,N_27962);
and U31392 (N_31392,N_27668,N_28991);
xor U31393 (N_31393,N_29419,N_28909);
nor U31394 (N_31394,N_29234,N_29783);
xor U31395 (N_31395,N_27623,N_29138);
or U31396 (N_31396,N_29080,N_27681);
and U31397 (N_31397,N_27676,N_29962);
xnor U31398 (N_31398,N_27594,N_27538);
xor U31399 (N_31399,N_29521,N_29710);
and U31400 (N_31400,N_29471,N_28416);
nand U31401 (N_31401,N_27595,N_28839);
nor U31402 (N_31402,N_28714,N_27839);
and U31403 (N_31403,N_29138,N_29717);
or U31404 (N_31404,N_29980,N_29940);
nor U31405 (N_31405,N_28767,N_28745);
or U31406 (N_31406,N_28366,N_28468);
or U31407 (N_31407,N_27664,N_27926);
xnor U31408 (N_31408,N_28416,N_28138);
xnor U31409 (N_31409,N_28321,N_29969);
or U31410 (N_31410,N_29052,N_28796);
nor U31411 (N_31411,N_28620,N_28430);
nand U31412 (N_31412,N_27631,N_28083);
xnor U31413 (N_31413,N_29416,N_28447);
and U31414 (N_31414,N_28786,N_27921);
nor U31415 (N_31415,N_28925,N_29154);
and U31416 (N_31416,N_29573,N_27548);
nand U31417 (N_31417,N_28352,N_29467);
xor U31418 (N_31418,N_29545,N_28455);
nand U31419 (N_31419,N_28943,N_28604);
or U31420 (N_31420,N_29904,N_28848);
and U31421 (N_31421,N_28461,N_27639);
or U31422 (N_31422,N_29986,N_29146);
xnor U31423 (N_31423,N_29190,N_29749);
nor U31424 (N_31424,N_29820,N_28981);
xnor U31425 (N_31425,N_28113,N_29816);
and U31426 (N_31426,N_29110,N_28820);
or U31427 (N_31427,N_29432,N_28464);
and U31428 (N_31428,N_27865,N_28625);
nand U31429 (N_31429,N_29262,N_28822);
and U31430 (N_31430,N_27765,N_28465);
or U31431 (N_31431,N_27903,N_27520);
nand U31432 (N_31432,N_28820,N_28010);
and U31433 (N_31433,N_27616,N_28896);
nor U31434 (N_31434,N_28621,N_29752);
and U31435 (N_31435,N_27979,N_28135);
or U31436 (N_31436,N_29388,N_29930);
xnor U31437 (N_31437,N_28795,N_27832);
and U31438 (N_31438,N_29570,N_27817);
xor U31439 (N_31439,N_29444,N_28563);
xor U31440 (N_31440,N_29491,N_28105);
or U31441 (N_31441,N_28412,N_29061);
or U31442 (N_31442,N_29949,N_28662);
and U31443 (N_31443,N_28735,N_27523);
xor U31444 (N_31444,N_28585,N_28534);
nand U31445 (N_31445,N_29415,N_29393);
xor U31446 (N_31446,N_27510,N_28702);
and U31447 (N_31447,N_29192,N_29271);
nor U31448 (N_31448,N_28929,N_28115);
and U31449 (N_31449,N_29655,N_28251);
xor U31450 (N_31450,N_29093,N_29868);
nand U31451 (N_31451,N_29747,N_29491);
or U31452 (N_31452,N_28473,N_28070);
and U31453 (N_31453,N_29524,N_27924);
and U31454 (N_31454,N_29300,N_29373);
nand U31455 (N_31455,N_29538,N_27902);
xnor U31456 (N_31456,N_29387,N_29953);
xor U31457 (N_31457,N_29927,N_29249);
and U31458 (N_31458,N_29083,N_28654);
or U31459 (N_31459,N_28191,N_29716);
nor U31460 (N_31460,N_28510,N_29840);
nand U31461 (N_31461,N_28365,N_28718);
and U31462 (N_31462,N_29360,N_27834);
or U31463 (N_31463,N_29640,N_27641);
or U31464 (N_31464,N_29251,N_28600);
and U31465 (N_31465,N_27523,N_29898);
nor U31466 (N_31466,N_27773,N_28158);
nand U31467 (N_31467,N_29904,N_27881);
xnor U31468 (N_31468,N_29352,N_27859);
and U31469 (N_31469,N_29510,N_28150);
xnor U31470 (N_31470,N_29204,N_28913);
or U31471 (N_31471,N_28579,N_29112);
xnor U31472 (N_31472,N_28218,N_27586);
xnor U31473 (N_31473,N_27650,N_27677);
and U31474 (N_31474,N_28423,N_29586);
and U31475 (N_31475,N_29828,N_29820);
nand U31476 (N_31476,N_28614,N_28052);
xor U31477 (N_31477,N_27936,N_29062);
nor U31478 (N_31478,N_29840,N_29934);
or U31479 (N_31479,N_27644,N_29898);
nand U31480 (N_31480,N_27922,N_29029);
or U31481 (N_31481,N_28145,N_28693);
and U31482 (N_31482,N_29915,N_29380);
nor U31483 (N_31483,N_27576,N_29663);
nor U31484 (N_31484,N_28350,N_28453);
nor U31485 (N_31485,N_29456,N_27952);
nand U31486 (N_31486,N_28708,N_28895);
nor U31487 (N_31487,N_27654,N_28791);
and U31488 (N_31488,N_29312,N_28651);
xnor U31489 (N_31489,N_28462,N_29259);
or U31490 (N_31490,N_29373,N_28530);
nand U31491 (N_31491,N_28323,N_29012);
or U31492 (N_31492,N_27888,N_29825);
and U31493 (N_31493,N_29226,N_29840);
nor U31494 (N_31494,N_28448,N_27712);
or U31495 (N_31495,N_29865,N_28277);
and U31496 (N_31496,N_29965,N_29037);
xor U31497 (N_31497,N_29472,N_28299);
and U31498 (N_31498,N_28419,N_28869);
nor U31499 (N_31499,N_27939,N_29572);
nand U31500 (N_31500,N_27568,N_29274);
or U31501 (N_31501,N_27818,N_27971);
and U31502 (N_31502,N_28181,N_27534);
xor U31503 (N_31503,N_28911,N_29349);
nand U31504 (N_31504,N_27614,N_27514);
or U31505 (N_31505,N_27562,N_27981);
nor U31506 (N_31506,N_27698,N_29019);
nor U31507 (N_31507,N_28661,N_28679);
nand U31508 (N_31508,N_27794,N_29571);
or U31509 (N_31509,N_29334,N_27799);
nand U31510 (N_31510,N_28376,N_27864);
and U31511 (N_31511,N_29793,N_28076);
nor U31512 (N_31512,N_28965,N_27591);
or U31513 (N_31513,N_29901,N_29821);
and U31514 (N_31514,N_29717,N_29178);
and U31515 (N_31515,N_27844,N_28258);
nand U31516 (N_31516,N_29729,N_29086);
or U31517 (N_31517,N_27705,N_29080);
nand U31518 (N_31518,N_27692,N_28986);
or U31519 (N_31519,N_27901,N_29846);
nor U31520 (N_31520,N_28808,N_29081);
xor U31521 (N_31521,N_29151,N_29412);
nand U31522 (N_31522,N_27866,N_29338);
nand U31523 (N_31523,N_28108,N_28266);
xnor U31524 (N_31524,N_28684,N_27806);
and U31525 (N_31525,N_27684,N_29564);
and U31526 (N_31526,N_28689,N_29914);
nand U31527 (N_31527,N_29571,N_29795);
xor U31528 (N_31528,N_29959,N_27990);
nand U31529 (N_31529,N_28409,N_27505);
nor U31530 (N_31530,N_28671,N_29947);
xor U31531 (N_31531,N_29509,N_28884);
nand U31532 (N_31532,N_28867,N_28717);
and U31533 (N_31533,N_29408,N_27597);
or U31534 (N_31534,N_28161,N_27714);
and U31535 (N_31535,N_28588,N_27935);
nand U31536 (N_31536,N_29788,N_28218);
xnor U31537 (N_31537,N_29837,N_27750);
and U31538 (N_31538,N_28018,N_29120);
nand U31539 (N_31539,N_29323,N_29719);
xor U31540 (N_31540,N_28176,N_29034);
or U31541 (N_31541,N_29239,N_28543);
and U31542 (N_31542,N_29188,N_28670);
or U31543 (N_31543,N_27587,N_28674);
or U31544 (N_31544,N_29614,N_29697);
nor U31545 (N_31545,N_29258,N_29482);
nor U31546 (N_31546,N_28636,N_29659);
xnor U31547 (N_31547,N_28733,N_28599);
nor U31548 (N_31548,N_27697,N_29102);
or U31549 (N_31549,N_28705,N_29953);
nor U31550 (N_31550,N_29714,N_28519);
and U31551 (N_31551,N_27717,N_28013);
nor U31552 (N_31552,N_28379,N_27683);
nor U31553 (N_31553,N_28539,N_28381);
or U31554 (N_31554,N_28383,N_28785);
xnor U31555 (N_31555,N_27813,N_27921);
or U31556 (N_31556,N_29708,N_28570);
nand U31557 (N_31557,N_29711,N_29490);
xor U31558 (N_31558,N_29683,N_27911);
nand U31559 (N_31559,N_29578,N_29720);
or U31560 (N_31560,N_29174,N_29894);
and U31561 (N_31561,N_28116,N_27543);
or U31562 (N_31562,N_29919,N_28094);
nand U31563 (N_31563,N_29446,N_28743);
nor U31564 (N_31564,N_27920,N_29655);
nor U31565 (N_31565,N_28835,N_28056);
or U31566 (N_31566,N_29513,N_27872);
nand U31567 (N_31567,N_27820,N_29986);
nand U31568 (N_31568,N_29095,N_28624);
nor U31569 (N_31569,N_28794,N_29351);
nand U31570 (N_31570,N_28766,N_28022);
nor U31571 (N_31571,N_28585,N_28670);
nand U31572 (N_31572,N_28990,N_29180);
nor U31573 (N_31573,N_29632,N_28582);
nand U31574 (N_31574,N_29251,N_29428);
nor U31575 (N_31575,N_29412,N_29877);
nor U31576 (N_31576,N_29493,N_29359);
xor U31577 (N_31577,N_29451,N_28806);
nor U31578 (N_31578,N_29242,N_28670);
nor U31579 (N_31579,N_27686,N_28361);
xor U31580 (N_31580,N_28493,N_29588);
and U31581 (N_31581,N_29285,N_28522);
xnor U31582 (N_31582,N_28841,N_29588);
or U31583 (N_31583,N_27953,N_27975);
nand U31584 (N_31584,N_28432,N_29824);
or U31585 (N_31585,N_29224,N_28373);
xnor U31586 (N_31586,N_27735,N_29136);
nor U31587 (N_31587,N_29544,N_28143);
nor U31588 (N_31588,N_29442,N_27756);
or U31589 (N_31589,N_29260,N_29944);
nor U31590 (N_31590,N_28054,N_29416);
nand U31591 (N_31591,N_29798,N_27622);
xnor U31592 (N_31592,N_29983,N_29239);
nor U31593 (N_31593,N_29018,N_28966);
nor U31594 (N_31594,N_28839,N_29025);
or U31595 (N_31595,N_29976,N_28334);
or U31596 (N_31596,N_29708,N_28712);
xnor U31597 (N_31597,N_28071,N_28524);
xor U31598 (N_31598,N_29576,N_28715);
and U31599 (N_31599,N_27659,N_28618);
or U31600 (N_31600,N_27968,N_29604);
xor U31601 (N_31601,N_27851,N_28372);
or U31602 (N_31602,N_28628,N_29008);
and U31603 (N_31603,N_29452,N_27782);
nor U31604 (N_31604,N_29267,N_28427);
xor U31605 (N_31605,N_28946,N_28261);
nand U31606 (N_31606,N_27649,N_28104);
and U31607 (N_31607,N_29190,N_29408);
xnor U31608 (N_31608,N_27792,N_28066);
and U31609 (N_31609,N_29886,N_29363);
xor U31610 (N_31610,N_28338,N_29706);
nor U31611 (N_31611,N_28574,N_29439);
nand U31612 (N_31612,N_29659,N_29100);
and U31613 (N_31613,N_27519,N_28048);
xnor U31614 (N_31614,N_28289,N_28854);
or U31615 (N_31615,N_28238,N_27552);
xor U31616 (N_31616,N_27846,N_28662);
nand U31617 (N_31617,N_27529,N_29802);
nand U31618 (N_31618,N_29920,N_28572);
or U31619 (N_31619,N_28477,N_29697);
nor U31620 (N_31620,N_28115,N_29198);
xor U31621 (N_31621,N_29204,N_28296);
or U31622 (N_31622,N_28981,N_28756);
nand U31623 (N_31623,N_28394,N_27989);
nor U31624 (N_31624,N_27587,N_29398);
xnor U31625 (N_31625,N_29719,N_29848);
nand U31626 (N_31626,N_28444,N_28620);
and U31627 (N_31627,N_28647,N_28403);
nand U31628 (N_31628,N_27986,N_28511);
nand U31629 (N_31629,N_28428,N_29521);
nor U31630 (N_31630,N_29786,N_27517);
xnor U31631 (N_31631,N_29100,N_28090);
and U31632 (N_31632,N_29133,N_28538);
nand U31633 (N_31633,N_27724,N_28452);
and U31634 (N_31634,N_29065,N_28941);
nor U31635 (N_31635,N_28978,N_27724);
or U31636 (N_31636,N_27923,N_29594);
xor U31637 (N_31637,N_27528,N_28554);
or U31638 (N_31638,N_27510,N_27525);
or U31639 (N_31639,N_29233,N_29416);
nor U31640 (N_31640,N_29305,N_29806);
nor U31641 (N_31641,N_28384,N_29467);
xnor U31642 (N_31642,N_28372,N_29985);
or U31643 (N_31643,N_28517,N_28500);
nand U31644 (N_31644,N_28686,N_28206);
nor U31645 (N_31645,N_29600,N_27840);
nor U31646 (N_31646,N_28994,N_29897);
nor U31647 (N_31647,N_28472,N_29835);
nand U31648 (N_31648,N_28037,N_29579);
and U31649 (N_31649,N_29246,N_29672);
xnor U31650 (N_31650,N_29003,N_29626);
nor U31651 (N_31651,N_28154,N_29201);
xor U31652 (N_31652,N_29789,N_28541);
nand U31653 (N_31653,N_27937,N_29324);
xor U31654 (N_31654,N_27623,N_29045);
nand U31655 (N_31655,N_29661,N_27905);
and U31656 (N_31656,N_27588,N_28039);
and U31657 (N_31657,N_27595,N_28292);
and U31658 (N_31658,N_27612,N_27901);
nor U31659 (N_31659,N_28935,N_29408);
or U31660 (N_31660,N_28321,N_28694);
or U31661 (N_31661,N_29415,N_29734);
nor U31662 (N_31662,N_29002,N_29828);
nor U31663 (N_31663,N_28650,N_28598);
xnor U31664 (N_31664,N_29113,N_28814);
or U31665 (N_31665,N_29713,N_29401);
nor U31666 (N_31666,N_28974,N_29840);
nand U31667 (N_31667,N_29758,N_28880);
nand U31668 (N_31668,N_27840,N_29390);
or U31669 (N_31669,N_28082,N_29980);
xor U31670 (N_31670,N_27669,N_29090);
xor U31671 (N_31671,N_28344,N_28746);
or U31672 (N_31672,N_28899,N_29891);
xor U31673 (N_31673,N_29355,N_29525);
nor U31674 (N_31674,N_28540,N_28683);
xnor U31675 (N_31675,N_28638,N_28113);
nor U31676 (N_31676,N_28497,N_27502);
or U31677 (N_31677,N_28399,N_29336);
or U31678 (N_31678,N_27836,N_27556);
and U31679 (N_31679,N_28082,N_28023);
xor U31680 (N_31680,N_28119,N_29979);
nor U31681 (N_31681,N_28635,N_27727);
and U31682 (N_31682,N_28951,N_28508);
nor U31683 (N_31683,N_28740,N_29204);
or U31684 (N_31684,N_29846,N_28922);
or U31685 (N_31685,N_27607,N_29792);
xnor U31686 (N_31686,N_27844,N_29408);
or U31687 (N_31687,N_29169,N_28959);
nor U31688 (N_31688,N_28014,N_27593);
or U31689 (N_31689,N_29510,N_28075);
nor U31690 (N_31690,N_29512,N_27856);
and U31691 (N_31691,N_28959,N_29047);
or U31692 (N_31692,N_27656,N_28501);
nand U31693 (N_31693,N_28136,N_27804);
xor U31694 (N_31694,N_27873,N_28125);
or U31695 (N_31695,N_27633,N_28052);
or U31696 (N_31696,N_28914,N_27585);
and U31697 (N_31697,N_28005,N_28765);
nor U31698 (N_31698,N_27896,N_29077);
nand U31699 (N_31699,N_27938,N_29761);
nor U31700 (N_31700,N_27897,N_28120);
nand U31701 (N_31701,N_29854,N_28677);
nand U31702 (N_31702,N_28516,N_29163);
xor U31703 (N_31703,N_29783,N_28660);
nor U31704 (N_31704,N_27509,N_29866);
or U31705 (N_31705,N_29031,N_28578);
and U31706 (N_31706,N_27657,N_29806);
or U31707 (N_31707,N_28960,N_27951);
and U31708 (N_31708,N_29987,N_29572);
nor U31709 (N_31709,N_29119,N_29649);
nand U31710 (N_31710,N_28511,N_29003);
or U31711 (N_31711,N_29812,N_28669);
nor U31712 (N_31712,N_29304,N_29024);
and U31713 (N_31713,N_27812,N_27536);
nand U31714 (N_31714,N_28139,N_29267);
xor U31715 (N_31715,N_29806,N_29046);
nand U31716 (N_31716,N_29209,N_27892);
xor U31717 (N_31717,N_27748,N_28821);
or U31718 (N_31718,N_28067,N_27540);
nand U31719 (N_31719,N_28010,N_27738);
or U31720 (N_31720,N_29492,N_29045);
xor U31721 (N_31721,N_28671,N_27725);
xor U31722 (N_31722,N_28808,N_28164);
or U31723 (N_31723,N_29416,N_28124);
or U31724 (N_31724,N_28826,N_29617);
nand U31725 (N_31725,N_28167,N_28102);
xnor U31726 (N_31726,N_28853,N_28354);
nand U31727 (N_31727,N_28656,N_29491);
xor U31728 (N_31728,N_29141,N_29424);
nand U31729 (N_31729,N_28237,N_29050);
nand U31730 (N_31730,N_27684,N_29305);
or U31731 (N_31731,N_29386,N_29902);
or U31732 (N_31732,N_28944,N_28835);
or U31733 (N_31733,N_28518,N_29600);
or U31734 (N_31734,N_28591,N_28545);
nor U31735 (N_31735,N_29599,N_29324);
or U31736 (N_31736,N_29547,N_28524);
nor U31737 (N_31737,N_27795,N_28328);
or U31738 (N_31738,N_27768,N_28766);
nand U31739 (N_31739,N_29836,N_27731);
and U31740 (N_31740,N_28293,N_28509);
or U31741 (N_31741,N_29276,N_28413);
or U31742 (N_31742,N_27992,N_29980);
or U31743 (N_31743,N_29424,N_29888);
nor U31744 (N_31744,N_27834,N_27973);
and U31745 (N_31745,N_28027,N_27860);
xnor U31746 (N_31746,N_29881,N_27547);
or U31747 (N_31747,N_27738,N_27634);
and U31748 (N_31748,N_28582,N_27998);
xnor U31749 (N_31749,N_29638,N_27729);
xor U31750 (N_31750,N_27575,N_29820);
or U31751 (N_31751,N_28470,N_29961);
or U31752 (N_31752,N_29153,N_27602);
or U31753 (N_31753,N_28778,N_29374);
nand U31754 (N_31754,N_28867,N_29980);
nor U31755 (N_31755,N_29282,N_29173);
nor U31756 (N_31756,N_27961,N_27756);
xnor U31757 (N_31757,N_29274,N_28950);
and U31758 (N_31758,N_28583,N_27581);
xnor U31759 (N_31759,N_27680,N_28749);
nand U31760 (N_31760,N_29271,N_29517);
nand U31761 (N_31761,N_28571,N_27761);
and U31762 (N_31762,N_28175,N_28605);
nor U31763 (N_31763,N_29388,N_28135);
nor U31764 (N_31764,N_28333,N_29946);
and U31765 (N_31765,N_29360,N_29058);
or U31766 (N_31766,N_28968,N_28231);
nand U31767 (N_31767,N_27588,N_29326);
nand U31768 (N_31768,N_28277,N_28633);
or U31769 (N_31769,N_27904,N_29753);
or U31770 (N_31770,N_27596,N_29228);
nor U31771 (N_31771,N_28280,N_28835);
or U31772 (N_31772,N_27965,N_27907);
nor U31773 (N_31773,N_27944,N_28654);
and U31774 (N_31774,N_27918,N_28649);
xor U31775 (N_31775,N_28427,N_27843);
and U31776 (N_31776,N_29739,N_29412);
nand U31777 (N_31777,N_29124,N_29467);
nand U31778 (N_31778,N_27623,N_29284);
nand U31779 (N_31779,N_29783,N_29232);
or U31780 (N_31780,N_29263,N_28315);
nand U31781 (N_31781,N_28791,N_27551);
nor U31782 (N_31782,N_28642,N_28219);
nor U31783 (N_31783,N_28807,N_28982);
and U31784 (N_31784,N_28565,N_29334);
and U31785 (N_31785,N_28988,N_29375);
or U31786 (N_31786,N_28903,N_29340);
xor U31787 (N_31787,N_28828,N_28224);
nand U31788 (N_31788,N_29625,N_28383);
and U31789 (N_31789,N_29753,N_28414);
and U31790 (N_31790,N_29229,N_28206);
xnor U31791 (N_31791,N_29189,N_28102);
xnor U31792 (N_31792,N_27595,N_28088);
nor U31793 (N_31793,N_29095,N_29821);
and U31794 (N_31794,N_27622,N_28712);
and U31795 (N_31795,N_28212,N_29271);
nand U31796 (N_31796,N_28564,N_27705);
nand U31797 (N_31797,N_29575,N_29112);
and U31798 (N_31798,N_27590,N_29608);
nand U31799 (N_31799,N_29380,N_29630);
and U31800 (N_31800,N_27663,N_27878);
xor U31801 (N_31801,N_28015,N_29017);
xnor U31802 (N_31802,N_28034,N_29372);
and U31803 (N_31803,N_28051,N_29467);
or U31804 (N_31804,N_28119,N_29573);
nor U31805 (N_31805,N_28144,N_27828);
and U31806 (N_31806,N_28228,N_28981);
nor U31807 (N_31807,N_28861,N_28388);
and U31808 (N_31808,N_28052,N_27829);
or U31809 (N_31809,N_29489,N_27500);
and U31810 (N_31810,N_27786,N_27557);
nor U31811 (N_31811,N_28757,N_28653);
and U31812 (N_31812,N_27921,N_27726);
nor U31813 (N_31813,N_29814,N_29488);
nand U31814 (N_31814,N_29654,N_29111);
nor U31815 (N_31815,N_28562,N_28817);
and U31816 (N_31816,N_27732,N_29859);
and U31817 (N_31817,N_29253,N_28232);
and U31818 (N_31818,N_28427,N_28443);
or U31819 (N_31819,N_29216,N_28962);
nand U31820 (N_31820,N_27792,N_28013);
xor U31821 (N_31821,N_27660,N_29095);
or U31822 (N_31822,N_28269,N_28519);
nand U31823 (N_31823,N_28574,N_29224);
nand U31824 (N_31824,N_29630,N_29426);
nor U31825 (N_31825,N_27632,N_29798);
or U31826 (N_31826,N_28067,N_28724);
nand U31827 (N_31827,N_27715,N_29489);
nand U31828 (N_31828,N_29004,N_29222);
and U31829 (N_31829,N_29127,N_28342);
nor U31830 (N_31830,N_27512,N_27956);
and U31831 (N_31831,N_28739,N_28687);
xor U31832 (N_31832,N_28016,N_29492);
nand U31833 (N_31833,N_29835,N_29817);
nand U31834 (N_31834,N_29560,N_27504);
nor U31835 (N_31835,N_29432,N_28956);
and U31836 (N_31836,N_29891,N_29339);
nand U31837 (N_31837,N_28531,N_29636);
nand U31838 (N_31838,N_27907,N_28405);
or U31839 (N_31839,N_27808,N_28156);
nor U31840 (N_31840,N_28991,N_28605);
or U31841 (N_31841,N_28023,N_28405);
nor U31842 (N_31842,N_27602,N_28039);
nor U31843 (N_31843,N_29135,N_28647);
and U31844 (N_31844,N_29841,N_29552);
nor U31845 (N_31845,N_28402,N_29199);
nand U31846 (N_31846,N_28463,N_29283);
nor U31847 (N_31847,N_29007,N_27695);
or U31848 (N_31848,N_29794,N_29454);
and U31849 (N_31849,N_28329,N_29904);
nor U31850 (N_31850,N_27775,N_28588);
or U31851 (N_31851,N_28897,N_29099);
xor U31852 (N_31852,N_27562,N_28391);
or U31853 (N_31853,N_29421,N_29857);
and U31854 (N_31854,N_29971,N_29741);
nor U31855 (N_31855,N_29750,N_28849);
nand U31856 (N_31856,N_29611,N_28171);
and U31857 (N_31857,N_28425,N_29071);
xnor U31858 (N_31858,N_27663,N_29674);
xor U31859 (N_31859,N_27574,N_27909);
xnor U31860 (N_31860,N_29339,N_29514);
nand U31861 (N_31861,N_27899,N_28468);
nor U31862 (N_31862,N_28242,N_27897);
xor U31863 (N_31863,N_27911,N_28785);
and U31864 (N_31864,N_29244,N_28139);
nor U31865 (N_31865,N_29707,N_28534);
xnor U31866 (N_31866,N_28996,N_27925);
nand U31867 (N_31867,N_29766,N_28901);
nand U31868 (N_31868,N_28156,N_28213);
nor U31869 (N_31869,N_28606,N_28223);
or U31870 (N_31870,N_27878,N_28812);
and U31871 (N_31871,N_28732,N_28820);
or U31872 (N_31872,N_29020,N_29516);
and U31873 (N_31873,N_28293,N_29968);
xnor U31874 (N_31874,N_28150,N_27908);
or U31875 (N_31875,N_29233,N_28458);
or U31876 (N_31876,N_29928,N_28773);
nand U31877 (N_31877,N_27961,N_29055);
and U31878 (N_31878,N_28468,N_28864);
xnor U31879 (N_31879,N_29714,N_28336);
xor U31880 (N_31880,N_27804,N_29793);
nor U31881 (N_31881,N_27919,N_29566);
nand U31882 (N_31882,N_27924,N_28552);
or U31883 (N_31883,N_28821,N_28834);
nor U31884 (N_31884,N_27815,N_29417);
nand U31885 (N_31885,N_29657,N_29892);
nand U31886 (N_31886,N_29605,N_29859);
xor U31887 (N_31887,N_29261,N_28262);
nand U31888 (N_31888,N_28453,N_28346);
or U31889 (N_31889,N_29077,N_28636);
nand U31890 (N_31890,N_29663,N_28362);
and U31891 (N_31891,N_28862,N_28245);
nand U31892 (N_31892,N_29199,N_28796);
and U31893 (N_31893,N_27930,N_27904);
xnor U31894 (N_31894,N_29743,N_29532);
nor U31895 (N_31895,N_29052,N_28249);
nor U31896 (N_31896,N_28451,N_28836);
or U31897 (N_31897,N_28027,N_29911);
or U31898 (N_31898,N_27658,N_28854);
nor U31899 (N_31899,N_28676,N_28281);
nor U31900 (N_31900,N_28693,N_28829);
or U31901 (N_31901,N_28292,N_29065);
nor U31902 (N_31902,N_29313,N_29336);
nor U31903 (N_31903,N_28906,N_28390);
nor U31904 (N_31904,N_29361,N_28894);
or U31905 (N_31905,N_28819,N_29466);
and U31906 (N_31906,N_28020,N_28669);
and U31907 (N_31907,N_29068,N_29103);
and U31908 (N_31908,N_29073,N_29046);
xnor U31909 (N_31909,N_29399,N_28370);
nor U31910 (N_31910,N_28873,N_28626);
nor U31911 (N_31911,N_28350,N_27974);
or U31912 (N_31912,N_29693,N_28808);
or U31913 (N_31913,N_28838,N_28271);
or U31914 (N_31914,N_28592,N_28040);
nor U31915 (N_31915,N_29790,N_29490);
xor U31916 (N_31916,N_27747,N_29419);
and U31917 (N_31917,N_28883,N_28891);
and U31918 (N_31918,N_29499,N_29205);
nand U31919 (N_31919,N_29653,N_28848);
nor U31920 (N_31920,N_28435,N_27721);
nand U31921 (N_31921,N_28645,N_29747);
or U31922 (N_31922,N_29549,N_27606);
xor U31923 (N_31923,N_28002,N_27903);
or U31924 (N_31924,N_28745,N_29604);
xnor U31925 (N_31925,N_29743,N_28433);
and U31926 (N_31926,N_28414,N_28234);
nand U31927 (N_31927,N_28942,N_29937);
nor U31928 (N_31928,N_27640,N_28296);
or U31929 (N_31929,N_29245,N_29714);
xnor U31930 (N_31930,N_29014,N_28291);
and U31931 (N_31931,N_28984,N_28173);
and U31932 (N_31932,N_28525,N_28123);
and U31933 (N_31933,N_28114,N_29479);
nand U31934 (N_31934,N_28819,N_29697);
and U31935 (N_31935,N_28628,N_29312);
xnor U31936 (N_31936,N_29603,N_27690);
nor U31937 (N_31937,N_28776,N_29890);
nor U31938 (N_31938,N_29340,N_27815);
nand U31939 (N_31939,N_27648,N_28590);
xor U31940 (N_31940,N_29998,N_27866);
or U31941 (N_31941,N_29754,N_28772);
xnor U31942 (N_31942,N_28175,N_29589);
xor U31943 (N_31943,N_29487,N_28267);
xor U31944 (N_31944,N_29846,N_28355);
and U31945 (N_31945,N_29360,N_27860);
and U31946 (N_31946,N_27746,N_28688);
and U31947 (N_31947,N_28752,N_27573);
or U31948 (N_31948,N_29890,N_29072);
nand U31949 (N_31949,N_28692,N_29180);
nand U31950 (N_31950,N_27771,N_28664);
nand U31951 (N_31951,N_28130,N_27983);
nand U31952 (N_31952,N_27510,N_29126);
nor U31953 (N_31953,N_27911,N_27969);
or U31954 (N_31954,N_27747,N_29881);
or U31955 (N_31955,N_29144,N_29650);
nand U31956 (N_31956,N_29606,N_29919);
xnor U31957 (N_31957,N_27936,N_29077);
nand U31958 (N_31958,N_27591,N_29813);
nor U31959 (N_31959,N_29672,N_29631);
nor U31960 (N_31960,N_29722,N_29971);
xor U31961 (N_31961,N_28350,N_27599);
or U31962 (N_31962,N_27924,N_27523);
nand U31963 (N_31963,N_29949,N_29012);
xnor U31964 (N_31964,N_28173,N_27627);
nand U31965 (N_31965,N_28305,N_29051);
and U31966 (N_31966,N_27516,N_27986);
nand U31967 (N_31967,N_28822,N_29047);
nand U31968 (N_31968,N_29431,N_28350);
and U31969 (N_31969,N_29035,N_29633);
nand U31970 (N_31970,N_29799,N_28095);
and U31971 (N_31971,N_28822,N_29839);
nor U31972 (N_31972,N_29595,N_28812);
and U31973 (N_31973,N_27538,N_28837);
and U31974 (N_31974,N_28298,N_28549);
xor U31975 (N_31975,N_29213,N_28940);
xor U31976 (N_31976,N_28740,N_28354);
nor U31977 (N_31977,N_27894,N_29440);
or U31978 (N_31978,N_28288,N_29625);
nor U31979 (N_31979,N_29495,N_29475);
nor U31980 (N_31980,N_29537,N_29174);
nor U31981 (N_31981,N_27778,N_27988);
xor U31982 (N_31982,N_28223,N_29928);
and U31983 (N_31983,N_28517,N_29945);
nor U31984 (N_31984,N_29805,N_27605);
nand U31985 (N_31985,N_29422,N_29876);
xnor U31986 (N_31986,N_29600,N_29660);
or U31987 (N_31987,N_29090,N_28345);
and U31988 (N_31988,N_29728,N_28807);
and U31989 (N_31989,N_28904,N_29866);
nand U31990 (N_31990,N_28341,N_29774);
and U31991 (N_31991,N_29865,N_29585);
or U31992 (N_31992,N_29609,N_28054);
nor U31993 (N_31993,N_29241,N_29157);
nor U31994 (N_31994,N_29501,N_29153);
and U31995 (N_31995,N_27605,N_28994);
xnor U31996 (N_31996,N_29257,N_29482);
and U31997 (N_31997,N_28991,N_29966);
or U31998 (N_31998,N_29786,N_29077);
or U31999 (N_31999,N_27956,N_28510);
xor U32000 (N_32000,N_29706,N_28861);
nand U32001 (N_32001,N_29607,N_28079);
nor U32002 (N_32002,N_29761,N_28764);
nand U32003 (N_32003,N_27906,N_28034);
xor U32004 (N_32004,N_28333,N_28558);
nor U32005 (N_32005,N_28493,N_27945);
or U32006 (N_32006,N_29326,N_29046);
nand U32007 (N_32007,N_29393,N_27647);
and U32008 (N_32008,N_29719,N_28465);
nor U32009 (N_32009,N_29117,N_28900);
or U32010 (N_32010,N_28294,N_29652);
and U32011 (N_32011,N_29500,N_29821);
xor U32012 (N_32012,N_29915,N_29173);
nand U32013 (N_32013,N_28999,N_28545);
or U32014 (N_32014,N_28041,N_28149);
nor U32015 (N_32015,N_28041,N_27827);
xnor U32016 (N_32016,N_29175,N_27878);
or U32017 (N_32017,N_27787,N_29774);
or U32018 (N_32018,N_29875,N_29752);
nor U32019 (N_32019,N_29043,N_29398);
and U32020 (N_32020,N_28224,N_29430);
nor U32021 (N_32021,N_28950,N_28292);
xor U32022 (N_32022,N_29248,N_29085);
nand U32023 (N_32023,N_28940,N_28976);
nor U32024 (N_32024,N_27653,N_27776);
xnor U32025 (N_32025,N_29387,N_29435);
xnor U32026 (N_32026,N_28434,N_28117);
xnor U32027 (N_32027,N_27966,N_29015);
nand U32028 (N_32028,N_29397,N_28701);
and U32029 (N_32029,N_28779,N_27888);
nor U32030 (N_32030,N_28152,N_28985);
or U32031 (N_32031,N_29308,N_27708);
nand U32032 (N_32032,N_29474,N_28066);
nor U32033 (N_32033,N_29301,N_27507);
and U32034 (N_32034,N_27687,N_27848);
nand U32035 (N_32035,N_29504,N_28860);
nand U32036 (N_32036,N_28491,N_29689);
or U32037 (N_32037,N_27738,N_29225);
or U32038 (N_32038,N_28734,N_29044);
and U32039 (N_32039,N_27841,N_29131);
xnor U32040 (N_32040,N_28981,N_28667);
xor U32041 (N_32041,N_28146,N_29098);
nor U32042 (N_32042,N_28606,N_27731);
nand U32043 (N_32043,N_28631,N_28292);
or U32044 (N_32044,N_29902,N_27602);
and U32045 (N_32045,N_29492,N_27521);
and U32046 (N_32046,N_28346,N_28994);
xor U32047 (N_32047,N_28898,N_28449);
or U32048 (N_32048,N_27505,N_29039);
and U32049 (N_32049,N_28132,N_29818);
xor U32050 (N_32050,N_27548,N_28685);
or U32051 (N_32051,N_27750,N_28855);
nor U32052 (N_32052,N_28136,N_28668);
xnor U32053 (N_32053,N_28251,N_29871);
and U32054 (N_32054,N_28854,N_29103);
or U32055 (N_32055,N_28433,N_29315);
xor U32056 (N_32056,N_29886,N_27587);
nor U32057 (N_32057,N_28672,N_28047);
and U32058 (N_32058,N_28506,N_27932);
or U32059 (N_32059,N_28438,N_28233);
nor U32060 (N_32060,N_28719,N_27759);
or U32061 (N_32061,N_27512,N_28325);
and U32062 (N_32062,N_29984,N_29639);
and U32063 (N_32063,N_29013,N_29520);
nand U32064 (N_32064,N_29599,N_27712);
nor U32065 (N_32065,N_29720,N_28300);
or U32066 (N_32066,N_27540,N_29410);
and U32067 (N_32067,N_29984,N_28036);
or U32068 (N_32068,N_28157,N_27957);
and U32069 (N_32069,N_29530,N_29434);
nor U32070 (N_32070,N_28623,N_29147);
nor U32071 (N_32071,N_29245,N_29890);
or U32072 (N_32072,N_27571,N_27650);
and U32073 (N_32073,N_27625,N_28790);
xor U32074 (N_32074,N_28380,N_29471);
and U32075 (N_32075,N_28218,N_28023);
nand U32076 (N_32076,N_27632,N_29020);
nand U32077 (N_32077,N_29792,N_28571);
xor U32078 (N_32078,N_28479,N_27732);
nor U32079 (N_32079,N_29316,N_29044);
xor U32080 (N_32080,N_28566,N_27850);
or U32081 (N_32081,N_27810,N_28567);
nor U32082 (N_32082,N_28093,N_27730);
nand U32083 (N_32083,N_28318,N_28293);
xnor U32084 (N_32084,N_29693,N_29185);
or U32085 (N_32085,N_28270,N_27910);
nor U32086 (N_32086,N_28346,N_29727);
xor U32087 (N_32087,N_27950,N_28693);
or U32088 (N_32088,N_29449,N_27716);
or U32089 (N_32089,N_29756,N_28274);
and U32090 (N_32090,N_28691,N_29157);
nor U32091 (N_32091,N_28673,N_29282);
xnor U32092 (N_32092,N_29322,N_28348);
or U32093 (N_32093,N_28893,N_29742);
or U32094 (N_32094,N_29194,N_29518);
nand U32095 (N_32095,N_29189,N_28764);
or U32096 (N_32096,N_28527,N_28436);
or U32097 (N_32097,N_28994,N_27675);
and U32098 (N_32098,N_28788,N_29849);
or U32099 (N_32099,N_27892,N_28694);
xnor U32100 (N_32100,N_29853,N_29907);
nor U32101 (N_32101,N_28601,N_29242);
nor U32102 (N_32102,N_29268,N_29834);
and U32103 (N_32103,N_29973,N_29656);
xor U32104 (N_32104,N_28906,N_29722);
or U32105 (N_32105,N_29788,N_27587);
nand U32106 (N_32106,N_28685,N_28687);
and U32107 (N_32107,N_27905,N_28718);
nor U32108 (N_32108,N_28162,N_27827);
or U32109 (N_32109,N_28926,N_29488);
or U32110 (N_32110,N_27741,N_28041);
or U32111 (N_32111,N_29010,N_28043);
or U32112 (N_32112,N_28472,N_28184);
and U32113 (N_32113,N_28354,N_28051);
xor U32114 (N_32114,N_29366,N_29732);
nand U32115 (N_32115,N_29610,N_28785);
or U32116 (N_32116,N_29853,N_29732);
or U32117 (N_32117,N_28041,N_28585);
and U32118 (N_32118,N_28418,N_28967);
nand U32119 (N_32119,N_29508,N_28279);
nor U32120 (N_32120,N_27832,N_27746);
xor U32121 (N_32121,N_29132,N_28167);
nand U32122 (N_32122,N_29052,N_28925);
nor U32123 (N_32123,N_29143,N_27607);
nor U32124 (N_32124,N_28415,N_27971);
nor U32125 (N_32125,N_28286,N_27558);
nand U32126 (N_32126,N_28329,N_29468);
nor U32127 (N_32127,N_29569,N_28329);
and U32128 (N_32128,N_28131,N_29096);
or U32129 (N_32129,N_29396,N_27645);
nor U32130 (N_32130,N_27761,N_28522);
nand U32131 (N_32131,N_27976,N_29257);
xor U32132 (N_32132,N_28677,N_29066);
xor U32133 (N_32133,N_28596,N_29127);
or U32134 (N_32134,N_28562,N_28700);
or U32135 (N_32135,N_29912,N_29871);
nand U32136 (N_32136,N_29347,N_27926);
nor U32137 (N_32137,N_27803,N_28059);
nor U32138 (N_32138,N_29654,N_29423);
xor U32139 (N_32139,N_27745,N_28724);
nor U32140 (N_32140,N_29346,N_28843);
and U32141 (N_32141,N_28480,N_28793);
nor U32142 (N_32142,N_27917,N_27971);
and U32143 (N_32143,N_28704,N_28360);
or U32144 (N_32144,N_28196,N_29468);
nor U32145 (N_32145,N_28066,N_28818);
nor U32146 (N_32146,N_29686,N_29724);
nor U32147 (N_32147,N_27696,N_28174);
xnor U32148 (N_32148,N_28572,N_28628);
or U32149 (N_32149,N_28718,N_29453);
or U32150 (N_32150,N_29767,N_29148);
and U32151 (N_32151,N_27554,N_27578);
nor U32152 (N_32152,N_29978,N_28724);
nand U32153 (N_32153,N_29120,N_29851);
and U32154 (N_32154,N_29773,N_27842);
xnor U32155 (N_32155,N_27591,N_29880);
xor U32156 (N_32156,N_28698,N_27728);
nor U32157 (N_32157,N_29393,N_27822);
nand U32158 (N_32158,N_27969,N_29977);
or U32159 (N_32159,N_28866,N_28723);
nor U32160 (N_32160,N_27607,N_28070);
nor U32161 (N_32161,N_29015,N_28124);
nor U32162 (N_32162,N_28423,N_29194);
nand U32163 (N_32163,N_29675,N_28340);
or U32164 (N_32164,N_28269,N_28413);
nand U32165 (N_32165,N_28678,N_27641);
or U32166 (N_32166,N_28123,N_27531);
and U32167 (N_32167,N_29550,N_29144);
or U32168 (N_32168,N_27794,N_28883);
and U32169 (N_32169,N_27909,N_29567);
nand U32170 (N_32170,N_28956,N_28681);
nor U32171 (N_32171,N_29921,N_28402);
and U32172 (N_32172,N_28157,N_29267);
nand U32173 (N_32173,N_29976,N_28163);
and U32174 (N_32174,N_29467,N_28797);
nand U32175 (N_32175,N_28353,N_28842);
xnor U32176 (N_32176,N_29317,N_29197);
nand U32177 (N_32177,N_28305,N_28907);
nor U32178 (N_32178,N_29242,N_29936);
xor U32179 (N_32179,N_29123,N_29784);
xnor U32180 (N_32180,N_28718,N_27927);
xor U32181 (N_32181,N_27750,N_28592);
xnor U32182 (N_32182,N_28949,N_28686);
or U32183 (N_32183,N_29689,N_28714);
or U32184 (N_32184,N_27837,N_27683);
nor U32185 (N_32185,N_27682,N_28869);
or U32186 (N_32186,N_29920,N_29486);
or U32187 (N_32187,N_28035,N_28582);
xnor U32188 (N_32188,N_27774,N_29663);
and U32189 (N_32189,N_29060,N_28395);
and U32190 (N_32190,N_28941,N_28581);
nand U32191 (N_32191,N_29601,N_27716);
and U32192 (N_32192,N_27663,N_28695);
xor U32193 (N_32193,N_28327,N_29197);
xnor U32194 (N_32194,N_29661,N_29191);
and U32195 (N_32195,N_28657,N_29181);
and U32196 (N_32196,N_28500,N_28803);
xor U32197 (N_32197,N_29621,N_28915);
nor U32198 (N_32198,N_28091,N_28506);
nand U32199 (N_32199,N_27661,N_28123);
nor U32200 (N_32200,N_27531,N_29779);
and U32201 (N_32201,N_29818,N_27931);
and U32202 (N_32202,N_29041,N_29850);
or U32203 (N_32203,N_29989,N_29936);
xor U32204 (N_32204,N_27637,N_27992);
or U32205 (N_32205,N_29436,N_29999);
and U32206 (N_32206,N_29058,N_28808);
and U32207 (N_32207,N_28442,N_29508);
nand U32208 (N_32208,N_29571,N_27534);
nand U32209 (N_32209,N_29087,N_29529);
nor U32210 (N_32210,N_27875,N_27523);
and U32211 (N_32211,N_29760,N_28159);
nor U32212 (N_32212,N_29603,N_28313);
and U32213 (N_32213,N_28178,N_29963);
nand U32214 (N_32214,N_28670,N_29096);
nor U32215 (N_32215,N_28689,N_27959);
nor U32216 (N_32216,N_28502,N_28198);
or U32217 (N_32217,N_28776,N_27583);
nand U32218 (N_32218,N_28235,N_27757);
xnor U32219 (N_32219,N_28100,N_28002);
xnor U32220 (N_32220,N_28100,N_29317);
and U32221 (N_32221,N_28106,N_27515);
nor U32222 (N_32222,N_29169,N_28848);
or U32223 (N_32223,N_29551,N_28765);
nor U32224 (N_32224,N_29118,N_29487);
nor U32225 (N_32225,N_29555,N_28697);
or U32226 (N_32226,N_27739,N_27578);
xnor U32227 (N_32227,N_27703,N_29587);
or U32228 (N_32228,N_28928,N_28829);
or U32229 (N_32229,N_28323,N_29874);
and U32230 (N_32230,N_28506,N_29193);
xor U32231 (N_32231,N_28063,N_29100);
and U32232 (N_32232,N_29448,N_28153);
nor U32233 (N_32233,N_28229,N_29224);
nand U32234 (N_32234,N_28168,N_28804);
nor U32235 (N_32235,N_29738,N_28970);
xor U32236 (N_32236,N_28542,N_29172);
nor U32237 (N_32237,N_27748,N_28338);
or U32238 (N_32238,N_28718,N_28721);
nor U32239 (N_32239,N_28789,N_27947);
xnor U32240 (N_32240,N_29543,N_29061);
nor U32241 (N_32241,N_29825,N_28051);
or U32242 (N_32242,N_29716,N_29704);
xnor U32243 (N_32243,N_29001,N_29828);
nor U32244 (N_32244,N_28394,N_28042);
nor U32245 (N_32245,N_29174,N_28348);
nand U32246 (N_32246,N_28175,N_28065);
nand U32247 (N_32247,N_28202,N_28629);
or U32248 (N_32248,N_29492,N_27668);
or U32249 (N_32249,N_29944,N_29519);
xor U32250 (N_32250,N_29711,N_29983);
or U32251 (N_32251,N_28384,N_27717);
nand U32252 (N_32252,N_27574,N_29621);
nand U32253 (N_32253,N_28003,N_27590);
nor U32254 (N_32254,N_28986,N_29065);
and U32255 (N_32255,N_29059,N_29630);
xnor U32256 (N_32256,N_29603,N_28450);
or U32257 (N_32257,N_27990,N_29943);
and U32258 (N_32258,N_27674,N_27809);
nand U32259 (N_32259,N_29103,N_28050);
nor U32260 (N_32260,N_28398,N_28730);
and U32261 (N_32261,N_29695,N_29801);
or U32262 (N_32262,N_27690,N_29393);
and U32263 (N_32263,N_29207,N_28813);
or U32264 (N_32264,N_28308,N_29254);
nor U32265 (N_32265,N_27850,N_28725);
or U32266 (N_32266,N_29417,N_28232);
nor U32267 (N_32267,N_27994,N_28057);
nor U32268 (N_32268,N_28265,N_29704);
nor U32269 (N_32269,N_28128,N_28284);
and U32270 (N_32270,N_29089,N_29781);
nor U32271 (N_32271,N_29084,N_28934);
and U32272 (N_32272,N_29970,N_27910);
nand U32273 (N_32273,N_29104,N_29597);
nand U32274 (N_32274,N_28452,N_29407);
and U32275 (N_32275,N_27662,N_28956);
nor U32276 (N_32276,N_28021,N_28878);
xor U32277 (N_32277,N_28646,N_29789);
xnor U32278 (N_32278,N_27588,N_28267);
or U32279 (N_32279,N_29469,N_29786);
nor U32280 (N_32280,N_28090,N_28499);
or U32281 (N_32281,N_28407,N_28514);
nor U32282 (N_32282,N_29643,N_29453);
and U32283 (N_32283,N_28687,N_29810);
xnor U32284 (N_32284,N_27569,N_28939);
or U32285 (N_32285,N_28658,N_29285);
or U32286 (N_32286,N_29048,N_28076);
and U32287 (N_32287,N_28747,N_29959);
nand U32288 (N_32288,N_28626,N_28111);
xnor U32289 (N_32289,N_27844,N_28748);
or U32290 (N_32290,N_29233,N_28007);
nand U32291 (N_32291,N_28089,N_28376);
nand U32292 (N_32292,N_29148,N_28147);
xnor U32293 (N_32293,N_27559,N_29935);
xnor U32294 (N_32294,N_27919,N_27992);
nand U32295 (N_32295,N_28255,N_28356);
or U32296 (N_32296,N_28039,N_27847);
nand U32297 (N_32297,N_28080,N_28024);
nor U32298 (N_32298,N_28935,N_28048);
nand U32299 (N_32299,N_28325,N_28235);
and U32300 (N_32300,N_28281,N_28589);
nand U32301 (N_32301,N_27926,N_29672);
and U32302 (N_32302,N_29238,N_29217);
xor U32303 (N_32303,N_28810,N_28818);
nand U32304 (N_32304,N_28406,N_27548);
nor U32305 (N_32305,N_28808,N_28737);
nand U32306 (N_32306,N_29189,N_27609);
and U32307 (N_32307,N_27884,N_28345);
or U32308 (N_32308,N_27906,N_27755);
xor U32309 (N_32309,N_29764,N_28555);
nand U32310 (N_32310,N_27904,N_29890);
or U32311 (N_32311,N_29700,N_29115);
and U32312 (N_32312,N_28233,N_28643);
nand U32313 (N_32313,N_28668,N_28061);
xnor U32314 (N_32314,N_29792,N_28010);
and U32315 (N_32315,N_29635,N_28438);
xor U32316 (N_32316,N_28255,N_27990);
nor U32317 (N_32317,N_29216,N_28184);
nand U32318 (N_32318,N_29603,N_28922);
or U32319 (N_32319,N_28503,N_28255);
nor U32320 (N_32320,N_28592,N_28645);
and U32321 (N_32321,N_29748,N_29347);
and U32322 (N_32322,N_28516,N_27780);
and U32323 (N_32323,N_28901,N_29086);
and U32324 (N_32324,N_28331,N_29158);
nor U32325 (N_32325,N_28021,N_27768);
nand U32326 (N_32326,N_28076,N_29008);
and U32327 (N_32327,N_27943,N_29143);
nand U32328 (N_32328,N_27791,N_29731);
or U32329 (N_32329,N_29271,N_27546);
nor U32330 (N_32330,N_28764,N_27912);
xor U32331 (N_32331,N_29428,N_28131);
nor U32332 (N_32332,N_28614,N_27530);
and U32333 (N_32333,N_28371,N_27891);
or U32334 (N_32334,N_28212,N_29966);
xnor U32335 (N_32335,N_29541,N_29176);
xnor U32336 (N_32336,N_27923,N_29120);
and U32337 (N_32337,N_28958,N_29918);
or U32338 (N_32338,N_28257,N_29194);
nor U32339 (N_32339,N_28742,N_27510);
and U32340 (N_32340,N_28189,N_28012);
nor U32341 (N_32341,N_29312,N_29550);
nor U32342 (N_32342,N_28090,N_28127);
nor U32343 (N_32343,N_29855,N_28999);
nor U32344 (N_32344,N_28004,N_28524);
xor U32345 (N_32345,N_28240,N_27869);
nand U32346 (N_32346,N_27892,N_28494);
nand U32347 (N_32347,N_28658,N_29991);
nand U32348 (N_32348,N_28078,N_28325);
nor U32349 (N_32349,N_28758,N_28971);
and U32350 (N_32350,N_29891,N_27821);
and U32351 (N_32351,N_28444,N_28690);
nand U32352 (N_32352,N_28188,N_29483);
and U32353 (N_32353,N_29647,N_29633);
and U32354 (N_32354,N_28280,N_29083);
nor U32355 (N_32355,N_29573,N_29366);
or U32356 (N_32356,N_29414,N_28193);
or U32357 (N_32357,N_27712,N_29330);
xnor U32358 (N_32358,N_28640,N_29224);
nand U32359 (N_32359,N_28742,N_27671);
or U32360 (N_32360,N_27741,N_28016);
xor U32361 (N_32361,N_27740,N_27641);
or U32362 (N_32362,N_28843,N_28086);
nand U32363 (N_32363,N_29538,N_29301);
xor U32364 (N_32364,N_29722,N_29820);
xor U32365 (N_32365,N_29471,N_29795);
xnor U32366 (N_32366,N_27561,N_27927);
or U32367 (N_32367,N_28171,N_28862);
and U32368 (N_32368,N_29368,N_29970);
nor U32369 (N_32369,N_29420,N_27628);
xor U32370 (N_32370,N_27878,N_29685);
and U32371 (N_32371,N_29502,N_29889);
xnor U32372 (N_32372,N_29347,N_29195);
or U32373 (N_32373,N_29956,N_29073);
xnor U32374 (N_32374,N_28612,N_29369);
nor U32375 (N_32375,N_28010,N_29727);
nor U32376 (N_32376,N_27943,N_28408);
nand U32377 (N_32377,N_28671,N_28876);
nand U32378 (N_32378,N_29481,N_27527);
nand U32379 (N_32379,N_28126,N_27530);
nor U32380 (N_32380,N_29785,N_27769);
nand U32381 (N_32381,N_29406,N_29617);
nand U32382 (N_32382,N_28587,N_27909);
nor U32383 (N_32383,N_29094,N_28359);
xnor U32384 (N_32384,N_27545,N_28591);
nor U32385 (N_32385,N_27856,N_29392);
xnor U32386 (N_32386,N_28738,N_28731);
nand U32387 (N_32387,N_29064,N_29771);
xor U32388 (N_32388,N_28629,N_27724);
xor U32389 (N_32389,N_29221,N_28285);
or U32390 (N_32390,N_28338,N_29606);
nor U32391 (N_32391,N_29480,N_29418);
nor U32392 (N_32392,N_29845,N_29225);
xor U32393 (N_32393,N_27592,N_27590);
or U32394 (N_32394,N_28636,N_28082);
nand U32395 (N_32395,N_27982,N_27694);
nand U32396 (N_32396,N_29363,N_27846);
nor U32397 (N_32397,N_29227,N_28886);
xor U32398 (N_32398,N_29679,N_28097);
and U32399 (N_32399,N_27787,N_27614);
nand U32400 (N_32400,N_29601,N_27618);
or U32401 (N_32401,N_29026,N_29733);
nor U32402 (N_32402,N_27512,N_29949);
and U32403 (N_32403,N_27942,N_29451);
and U32404 (N_32404,N_28710,N_28470);
and U32405 (N_32405,N_28896,N_28667);
nand U32406 (N_32406,N_28617,N_28367);
nand U32407 (N_32407,N_27860,N_28495);
or U32408 (N_32408,N_29841,N_28327);
nor U32409 (N_32409,N_29747,N_28820);
xor U32410 (N_32410,N_29128,N_28550);
or U32411 (N_32411,N_28414,N_28788);
or U32412 (N_32412,N_27856,N_29089);
nor U32413 (N_32413,N_29706,N_29775);
nand U32414 (N_32414,N_28647,N_28089);
or U32415 (N_32415,N_27571,N_27717);
nor U32416 (N_32416,N_29041,N_27571);
or U32417 (N_32417,N_28312,N_28345);
nand U32418 (N_32418,N_27810,N_28401);
xor U32419 (N_32419,N_29844,N_28418);
nand U32420 (N_32420,N_28740,N_27884);
and U32421 (N_32421,N_29609,N_29063);
and U32422 (N_32422,N_29959,N_28670);
nor U32423 (N_32423,N_29357,N_29024);
xnor U32424 (N_32424,N_29551,N_28821);
and U32425 (N_32425,N_29808,N_29351);
nand U32426 (N_32426,N_29366,N_29029);
nand U32427 (N_32427,N_27900,N_27713);
nor U32428 (N_32428,N_29199,N_27670);
nand U32429 (N_32429,N_28394,N_29375);
and U32430 (N_32430,N_28505,N_27956);
nor U32431 (N_32431,N_29375,N_29557);
xnor U32432 (N_32432,N_29914,N_29820);
and U32433 (N_32433,N_28731,N_29607);
nand U32434 (N_32434,N_29806,N_29584);
xnor U32435 (N_32435,N_29352,N_29465);
nand U32436 (N_32436,N_28653,N_27769);
or U32437 (N_32437,N_28886,N_29983);
xnor U32438 (N_32438,N_29859,N_27571);
or U32439 (N_32439,N_28658,N_29973);
nor U32440 (N_32440,N_28946,N_29319);
or U32441 (N_32441,N_28281,N_28208);
or U32442 (N_32442,N_28159,N_28437);
and U32443 (N_32443,N_27504,N_29470);
nand U32444 (N_32444,N_29625,N_29111);
and U32445 (N_32445,N_29006,N_29930);
nor U32446 (N_32446,N_28115,N_28637);
and U32447 (N_32447,N_28113,N_27813);
nand U32448 (N_32448,N_29439,N_29901);
xnor U32449 (N_32449,N_28484,N_29134);
nand U32450 (N_32450,N_29719,N_29147);
and U32451 (N_32451,N_29791,N_29850);
nand U32452 (N_32452,N_27515,N_29179);
nand U32453 (N_32453,N_29303,N_27701);
nand U32454 (N_32454,N_28492,N_28321);
and U32455 (N_32455,N_29177,N_28671);
or U32456 (N_32456,N_29667,N_29811);
xnor U32457 (N_32457,N_28463,N_27563);
and U32458 (N_32458,N_27568,N_28001);
xor U32459 (N_32459,N_29922,N_29316);
or U32460 (N_32460,N_29106,N_28216);
or U32461 (N_32461,N_27795,N_27718);
and U32462 (N_32462,N_28470,N_29982);
or U32463 (N_32463,N_29340,N_28694);
and U32464 (N_32464,N_27665,N_29168);
nor U32465 (N_32465,N_27519,N_29749);
nand U32466 (N_32466,N_28278,N_28246);
xnor U32467 (N_32467,N_28540,N_29303);
xnor U32468 (N_32468,N_28867,N_28271);
or U32469 (N_32469,N_29742,N_28975);
or U32470 (N_32470,N_27884,N_29213);
and U32471 (N_32471,N_29757,N_27530);
or U32472 (N_32472,N_29907,N_29440);
xor U32473 (N_32473,N_28580,N_28312);
nor U32474 (N_32474,N_29791,N_29137);
or U32475 (N_32475,N_29724,N_28347);
xor U32476 (N_32476,N_29343,N_29181);
nand U32477 (N_32477,N_28917,N_28555);
xor U32478 (N_32478,N_29678,N_27537);
xor U32479 (N_32479,N_28503,N_28657);
nand U32480 (N_32480,N_29049,N_28537);
xor U32481 (N_32481,N_27775,N_28515);
and U32482 (N_32482,N_29734,N_27634);
and U32483 (N_32483,N_27539,N_29328);
nor U32484 (N_32484,N_29823,N_28689);
and U32485 (N_32485,N_28786,N_28646);
and U32486 (N_32486,N_29101,N_28090);
nor U32487 (N_32487,N_29047,N_29355);
xor U32488 (N_32488,N_27786,N_28750);
nor U32489 (N_32489,N_28510,N_28605);
nand U32490 (N_32490,N_27505,N_28632);
xor U32491 (N_32491,N_28300,N_27725);
xor U32492 (N_32492,N_29943,N_29051);
and U32493 (N_32493,N_29402,N_28857);
nor U32494 (N_32494,N_27797,N_28979);
nand U32495 (N_32495,N_29508,N_29790);
xnor U32496 (N_32496,N_29390,N_29139);
and U32497 (N_32497,N_29132,N_28057);
or U32498 (N_32498,N_29493,N_28653);
nand U32499 (N_32499,N_28272,N_29825);
or U32500 (N_32500,N_32185,N_30090);
or U32501 (N_32501,N_30866,N_30905);
nand U32502 (N_32502,N_31558,N_31478);
nand U32503 (N_32503,N_31578,N_31136);
nor U32504 (N_32504,N_31936,N_31041);
xnor U32505 (N_32505,N_32151,N_30276);
xor U32506 (N_32506,N_30924,N_32350);
xnor U32507 (N_32507,N_32163,N_31516);
and U32508 (N_32508,N_31490,N_31570);
nand U32509 (N_32509,N_30889,N_30916);
or U32510 (N_32510,N_31542,N_30001);
or U32511 (N_32511,N_32036,N_31023);
nor U32512 (N_32512,N_30321,N_30672);
xor U32513 (N_32513,N_30060,N_30418);
nand U32514 (N_32514,N_30717,N_31817);
or U32515 (N_32515,N_30368,N_30176);
and U32516 (N_32516,N_31218,N_31195);
and U32517 (N_32517,N_30132,N_31322);
and U32518 (N_32518,N_32331,N_31186);
nand U32519 (N_32519,N_32094,N_30845);
nor U32520 (N_32520,N_32460,N_32464);
and U32521 (N_32521,N_31829,N_32313);
xor U32522 (N_32522,N_32016,N_32011);
xnor U32523 (N_32523,N_31379,N_32021);
xor U32524 (N_32524,N_31224,N_31546);
xnor U32525 (N_32525,N_30912,N_32299);
nor U32526 (N_32526,N_30935,N_30358);
or U32527 (N_32527,N_30265,N_31530);
and U32528 (N_32528,N_31588,N_31622);
xor U32529 (N_32529,N_31400,N_31076);
nor U32530 (N_32530,N_30864,N_30365);
xnor U32531 (N_32531,N_31151,N_31980);
xor U32532 (N_32532,N_31370,N_32069);
nand U32533 (N_32533,N_31914,N_31659);
nand U32534 (N_32534,N_31859,N_30204);
or U32535 (N_32535,N_30434,N_32106);
nand U32536 (N_32536,N_31531,N_30976);
nor U32537 (N_32537,N_31624,N_30712);
nand U32538 (N_32538,N_31437,N_31685);
and U32539 (N_32539,N_31638,N_31392);
xor U32540 (N_32540,N_31726,N_31822);
nand U32541 (N_32541,N_32415,N_30183);
nor U32542 (N_32542,N_31716,N_30240);
or U32543 (N_32543,N_32008,N_30764);
and U32544 (N_32544,N_32167,N_31493);
and U32545 (N_32545,N_30097,N_31368);
xnor U32546 (N_32546,N_30332,N_30068);
xor U32547 (N_32547,N_31335,N_31203);
or U32548 (N_32548,N_30218,N_31728);
or U32549 (N_32549,N_30596,N_30000);
or U32550 (N_32550,N_32043,N_30311);
or U32551 (N_32551,N_31469,N_31489);
and U32552 (N_32552,N_30439,N_30038);
and U32553 (N_32553,N_30887,N_31474);
or U32554 (N_32554,N_30522,N_30566);
or U32555 (N_32555,N_31359,N_30710);
nor U32556 (N_32556,N_31645,N_31727);
and U32557 (N_32557,N_31950,N_31700);
and U32558 (N_32558,N_32403,N_32286);
and U32559 (N_32559,N_31032,N_31197);
and U32560 (N_32560,N_30496,N_31166);
and U32561 (N_32561,N_32079,N_31426);
xor U32562 (N_32562,N_32146,N_31770);
and U32563 (N_32563,N_32120,N_30751);
and U32564 (N_32564,N_30286,N_32044);
or U32565 (N_32565,N_31358,N_31165);
xnor U32566 (N_32566,N_31255,N_30585);
xor U32567 (N_32567,N_30050,N_31154);
xor U32568 (N_32568,N_30174,N_31360);
xor U32569 (N_32569,N_30260,N_31665);
xor U32570 (N_32570,N_30164,N_31124);
xnor U32571 (N_32571,N_30216,N_31177);
nand U32572 (N_32572,N_30476,N_31290);
and U32573 (N_32573,N_31745,N_30033);
and U32574 (N_32574,N_30064,N_32047);
xnor U32575 (N_32575,N_30919,N_31781);
and U32576 (N_32576,N_32272,N_30518);
or U32577 (N_32577,N_32166,N_31621);
nand U32578 (N_32578,N_30115,N_31402);
and U32579 (N_32579,N_30885,N_30709);
nor U32580 (N_32580,N_30612,N_31214);
nor U32581 (N_32581,N_30161,N_30108);
and U32582 (N_32582,N_31088,N_30486);
nand U32583 (N_32583,N_30309,N_31891);
and U32584 (N_32584,N_32294,N_30104);
nand U32585 (N_32585,N_30129,N_30295);
xor U32586 (N_32586,N_31030,N_30150);
and U32587 (N_32587,N_30373,N_32086);
nand U32588 (N_32588,N_32053,N_31742);
or U32589 (N_32589,N_32401,N_30839);
and U32590 (N_32590,N_32127,N_31675);
nand U32591 (N_32591,N_30978,N_30614);
or U32592 (N_32592,N_31539,N_31524);
nor U32593 (N_32593,N_31757,N_32051);
nand U32594 (N_32594,N_31485,N_32027);
nand U32595 (N_32595,N_32372,N_31438);
nand U32596 (N_32596,N_31107,N_32022);
xor U32597 (N_32597,N_31862,N_30966);
nand U32598 (N_32598,N_31086,N_30054);
nand U32599 (N_32599,N_30865,N_32203);
and U32600 (N_32600,N_31634,N_31000);
xnor U32601 (N_32601,N_31673,N_31439);
or U32602 (N_32602,N_30523,N_31432);
xor U32603 (N_32603,N_31674,N_32394);
nand U32604 (N_32604,N_30035,N_30209);
nor U32605 (N_32605,N_32065,N_30472);
xor U32606 (N_32606,N_32380,N_32179);
xnor U32607 (N_32607,N_31344,N_32247);
nand U32608 (N_32608,N_30600,N_31142);
and U32609 (N_32609,N_30473,N_31557);
nand U32610 (N_32610,N_30424,N_30202);
nor U32611 (N_32611,N_30983,N_31187);
nand U32612 (N_32612,N_30113,N_30714);
nand U32613 (N_32613,N_31190,N_31317);
nor U32614 (N_32614,N_30009,N_32335);
and U32615 (N_32615,N_30767,N_30120);
nor U32616 (N_32616,N_30810,N_31475);
xor U32617 (N_32617,N_30993,N_30957);
nand U32618 (N_32618,N_32142,N_31904);
or U32619 (N_32619,N_31461,N_30366);
nand U32620 (N_32620,N_31733,N_30383);
or U32621 (N_32621,N_31605,N_32041);
nor U32622 (N_32622,N_31307,N_31563);
nand U32623 (N_32623,N_31851,N_31927);
nand U32624 (N_32624,N_31212,N_31900);
and U32625 (N_32625,N_32208,N_31794);
or U32626 (N_32626,N_32251,N_30395);
xnor U32627 (N_32627,N_30632,N_30625);
nand U32628 (N_32628,N_31259,N_31408);
nor U32629 (N_32629,N_30055,N_30922);
nor U32630 (N_32630,N_32327,N_31269);
nor U32631 (N_32631,N_32239,N_31574);
nand U32632 (N_32632,N_30788,N_31713);
nand U32633 (N_32633,N_31085,N_30720);
xnor U32634 (N_32634,N_31951,N_30508);
xnor U32635 (N_32635,N_30431,N_31051);
xnor U32636 (N_32636,N_30991,N_31866);
and U32637 (N_32637,N_30151,N_31972);
nor U32638 (N_32638,N_31608,N_30606);
nor U32639 (N_32639,N_31081,N_31689);
nor U32640 (N_32640,N_31620,N_30967);
nand U32641 (N_32641,N_30039,N_31202);
or U32642 (N_32642,N_31281,N_31378);
nand U32643 (N_32643,N_31776,N_31056);
or U32644 (N_32644,N_30323,N_31725);
nor U32645 (N_32645,N_30729,N_32402);
xor U32646 (N_32646,N_31140,N_31057);
and U32647 (N_32647,N_32430,N_31940);
and U32648 (N_32648,N_31007,N_30586);
nand U32649 (N_32649,N_31704,N_30633);
nand U32650 (N_32650,N_31397,N_30812);
nand U32651 (N_32651,N_30313,N_31793);
or U32652 (N_32652,N_31958,N_31048);
xor U32653 (N_32653,N_31006,N_31434);
nand U32654 (N_32654,N_30438,N_30900);
and U32655 (N_32655,N_30381,N_30180);
or U32656 (N_32656,N_30804,N_30364);
and U32657 (N_32657,N_30750,N_32276);
or U32658 (N_32658,N_32024,N_32207);
or U32659 (N_32659,N_30809,N_30584);
nor U32660 (N_32660,N_31897,N_31792);
nand U32661 (N_32661,N_30731,N_31903);
xor U32662 (N_32662,N_30911,N_32152);
nor U32663 (N_32663,N_30948,N_32071);
nand U32664 (N_32664,N_32359,N_31176);
or U32665 (N_32665,N_31134,N_30956);
nor U32666 (N_32666,N_31923,N_30455);
nor U32667 (N_32667,N_31129,N_31816);
xor U32668 (N_32668,N_32366,N_32186);
nor U32669 (N_32669,N_31644,N_32252);
nand U32670 (N_32670,N_30899,N_32305);
and U32671 (N_32671,N_30768,N_30504);
xnor U32672 (N_32672,N_30399,N_30818);
nand U32673 (N_32673,N_30384,N_31948);
nand U32674 (N_32674,N_31744,N_30190);
or U32675 (N_32675,N_30646,N_30917);
and U32676 (N_32676,N_31842,N_31273);
or U32677 (N_32677,N_30601,N_31584);
xnor U32678 (N_32678,N_30668,N_31755);
xnor U32679 (N_32679,N_31931,N_31029);
and U32680 (N_32680,N_31517,N_31435);
xor U32681 (N_32681,N_31099,N_31118);
and U32682 (N_32682,N_30662,N_30985);
nand U32683 (N_32683,N_32153,N_30189);
xnor U32684 (N_32684,N_31483,N_32377);
or U32685 (N_32685,N_30279,N_32360);
nor U32686 (N_32686,N_32499,N_32150);
nor U32687 (N_32687,N_30319,N_30569);
xor U32688 (N_32688,N_31305,N_31836);
and U32689 (N_32689,N_32217,N_31774);
or U32690 (N_32690,N_31497,N_30121);
xor U32691 (N_32691,N_31592,N_30460);
nand U32692 (N_32692,N_30085,N_32479);
and U32693 (N_32693,N_30029,N_31702);
nor U32694 (N_32694,N_30968,N_30241);
nor U32695 (N_32695,N_30023,N_32189);
nor U32696 (N_32696,N_31500,N_31871);
xor U32697 (N_32697,N_32265,N_32116);
nor U32698 (N_32698,N_31921,N_32278);
xor U32699 (N_32699,N_31961,N_30589);
and U32700 (N_32700,N_30172,N_31310);
or U32701 (N_32701,N_31089,N_31430);
or U32702 (N_32702,N_31907,N_31220);
nand U32703 (N_32703,N_31188,N_31382);
nor U32704 (N_32704,N_31441,N_31762);
or U32705 (N_32705,N_31445,N_30410);
or U32706 (N_32706,N_30937,N_30745);
or U32707 (N_32707,N_31298,N_32446);
nor U32708 (N_32708,N_32213,N_30292);
or U32709 (N_32709,N_31328,N_31922);
nand U32710 (N_32710,N_32255,N_31155);
xnor U32711 (N_32711,N_31387,N_30401);
and U32712 (N_32712,N_31686,N_30213);
xor U32713 (N_32713,N_32199,N_30503);
or U32714 (N_32714,N_30275,N_32264);
xnor U32715 (N_32715,N_31103,N_30567);
nand U32716 (N_32716,N_30106,N_30699);
or U32717 (N_32717,N_30941,N_31073);
nor U32718 (N_32718,N_30463,N_30509);
or U32719 (N_32719,N_30031,N_30233);
xor U32720 (N_32720,N_32165,N_30036);
nor U32721 (N_32721,N_31090,N_30010);
and U32722 (N_32722,N_30203,N_31893);
nor U32723 (N_32723,N_31163,N_31204);
nor U32724 (N_32724,N_32450,N_32442);
nor U32725 (N_32725,N_30640,N_32418);
and U32726 (N_32726,N_32145,N_31144);
or U32727 (N_32727,N_30506,N_31607);
nor U32728 (N_32728,N_32381,N_30666);
xor U32729 (N_32729,N_31185,N_30718);
and U32730 (N_32730,N_31617,N_32107);
nor U32731 (N_32731,N_31679,N_31403);
nand U32732 (N_32732,N_30676,N_30101);
xor U32733 (N_32733,N_31106,N_31182);
xor U32734 (N_32734,N_30689,N_32096);
nor U32735 (N_32735,N_30065,N_31910);
xor U32736 (N_32736,N_31208,N_30583);
nand U32737 (N_32737,N_30568,N_32218);
xnor U32738 (N_32738,N_30177,N_30197);
nand U32739 (N_32739,N_32445,N_32438);
nor U32740 (N_32740,N_30784,N_30091);
or U32741 (N_32741,N_30385,N_31348);
nor U32742 (N_32742,N_30477,N_31913);
xnor U32743 (N_32743,N_30843,N_31172);
and U32744 (N_32744,N_31556,N_31612);
and U32745 (N_32745,N_32300,N_31293);
nor U32746 (N_32746,N_31655,N_30847);
nand U32747 (N_32747,N_32470,N_32364);
nand U32748 (N_32748,N_30778,N_30391);
and U32749 (N_32749,N_30524,N_32237);
nand U32750 (N_32750,N_30579,N_30958);
nor U32751 (N_32751,N_31451,N_30988);
or U32752 (N_32752,N_30918,N_30761);
nand U32753 (N_32753,N_32287,N_32469);
nor U32754 (N_32754,N_32405,N_32441);
nor U32755 (N_32755,N_32160,N_31336);
nor U32756 (N_32756,N_31724,N_31362);
or U32757 (N_32757,N_32040,N_31593);
or U32758 (N_32758,N_32088,N_31552);
xor U32759 (N_32759,N_30791,N_30157);
or U32760 (N_32760,N_30474,N_32383);
nand U32761 (N_32761,N_31618,N_32281);
or U32762 (N_32762,N_31960,N_31035);
and U32763 (N_32763,N_31974,N_31941);
and U32764 (N_32764,N_30790,N_31241);
xor U32765 (N_32765,N_30094,N_32156);
and U32766 (N_32766,N_31295,N_30794);
or U32767 (N_32767,N_30015,N_31561);
nand U32768 (N_32768,N_31853,N_32092);
or U32769 (N_32769,N_30757,N_30637);
xor U32770 (N_32770,N_32288,N_31878);
nor U32771 (N_32771,N_30603,N_32333);
nand U32772 (N_32772,N_30874,N_32387);
nor U32773 (N_32773,N_30652,N_32097);
nor U32774 (N_32774,N_30647,N_31161);
or U32775 (N_32775,N_31270,N_31918);
nor U32776 (N_32776,N_32461,N_32173);
or U32777 (N_32777,N_32013,N_30131);
or U32778 (N_32778,N_30975,N_31943);
nand U32779 (N_32779,N_30428,N_32411);
xor U32780 (N_32780,N_32439,N_32001);
xnor U32781 (N_32781,N_30581,N_31016);
nand U32782 (N_32782,N_30012,N_32244);
or U32783 (N_32783,N_31587,N_31882);
or U32784 (N_32784,N_32090,N_32201);
nor U32785 (N_32785,N_31111,N_30738);
xor U32786 (N_32786,N_31779,N_30403);
nand U32787 (N_32787,N_31651,N_31775);
or U32788 (N_32788,N_30682,N_32080);
nand U32789 (N_32789,N_30697,N_30736);
nand U32790 (N_32790,N_31275,N_30374);
xor U32791 (N_32791,N_31534,N_32341);
nor U32792 (N_32792,N_32275,N_32282);
xnor U32793 (N_32793,N_30072,N_30507);
and U32794 (N_32794,N_31283,N_30227);
and U32795 (N_32795,N_30499,N_32225);
nor U32796 (N_32796,N_30946,N_30742);
and U32797 (N_32797,N_30214,N_30427);
and U32798 (N_32798,N_30570,N_32183);
nand U32799 (N_32799,N_31738,N_30136);
nor U32800 (N_32800,N_32374,N_32235);
or U32801 (N_32801,N_31422,N_31070);
nand U32802 (N_32802,N_32444,N_30005);
nand U32803 (N_32803,N_31609,N_32322);
nand U32804 (N_32804,N_30182,N_30206);
nand U32805 (N_32805,N_32228,N_30501);
nor U32806 (N_32806,N_30389,N_30343);
nor U32807 (N_32807,N_31569,N_30327);
nand U32808 (N_32808,N_31394,N_31078);
nor U32809 (N_32809,N_30609,N_31998);
nand U32810 (N_32810,N_31671,N_31205);
xnor U32811 (N_32811,N_30114,N_32240);
and U32812 (N_32812,N_32326,N_30663);
or U32813 (N_32813,N_32370,N_31989);
and U32814 (N_32814,N_30416,N_31374);
or U32815 (N_32815,N_31267,N_31846);
xor U32816 (N_32816,N_31037,N_30133);
and U32817 (N_32817,N_32298,N_31278);
nand U32818 (N_32818,N_31093,N_31223);
and U32819 (N_32819,N_30304,N_32078);
xnor U32820 (N_32820,N_30858,N_31460);
xor U32821 (N_32821,N_30034,N_30653);
nand U32822 (N_32822,N_31573,N_31581);
nor U32823 (N_32823,N_30184,N_30059);
or U32824 (N_32824,N_31855,N_31537);
and U32825 (N_32825,N_30261,N_31019);
and U32826 (N_32826,N_31896,N_30169);
or U32827 (N_32827,N_30667,N_30780);
and U32828 (N_32828,N_31881,N_30686);
or U32829 (N_32829,N_32422,N_31911);
nand U32830 (N_32830,N_30823,N_30397);
nor U32831 (N_32831,N_30215,N_31759);
or U32832 (N_32832,N_32064,N_31292);
nand U32833 (N_32833,N_32279,N_30430);
nor U32834 (N_32834,N_31691,N_30696);
xor U32835 (N_32835,N_30316,N_30145);
or U32836 (N_32836,N_30591,N_30722);
nand U32837 (N_32837,N_30923,N_30003);
nand U32838 (N_32838,N_32123,N_32385);
or U32839 (N_32839,N_32347,N_32081);
nand U32840 (N_32840,N_30974,N_30521);
nor U32841 (N_32841,N_32118,N_30692);
xnor U32842 (N_32842,N_31912,N_30084);
nor U32843 (N_32843,N_32162,N_31004);
xnor U32844 (N_32844,N_31521,N_30868);
xor U32845 (N_32845,N_32436,N_30895);
and U32846 (N_32846,N_30449,N_30724);
or U32847 (N_32847,N_32483,N_30560);
and U32848 (N_32848,N_31338,N_30730);
xor U32849 (N_32849,N_31141,N_32238);
and U32850 (N_32850,N_30677,N_32397);
or U32851 (N_32851,N_30314,N_31981);
nand U32852 (N_32852,N_32109,N_30109);
or U32853 (N_32853,N_30361,N_32306);
and U32854 (N_32854,N_30763,N_30655);
nand U32855 (N_32855,N_31173,N_30456);
nand U32856 (N_32856,N_30540,N_30117);
nand U32857 (N_32857,N_30628,N_31250);
xnor U32858 (N_32858,N_32268,N_31228);
nand U32859 (N_32859,N_30087,N_31311);
nand U32860 (N_32860,N_30402,N_31240);
xor U32861 (N_32861,N_30898,N_32178);
nand U32862 (N_32862,N_30278,N_31063);
or U32863 (N_32863,N_31002,N_31701);
nor U32864 (N_32864,N_30857,N_30777);
and U32865 (N_32865,N_30753,N_30510);
xor U32866 (N_32866,N_31105,N_31590);
or U32867 (N_32867,N_30852,N_30149);
xor U32868 (N_32868,N_31719,N_31528);
nor U32869 (N_32869,N_31681,N_32474);
and U32870 (N_32870,N_31484,N_31211);
nor U32871 (N_32871,N_31800,N_30027);
and U32872 (N_32872,N_32354,N_30681);
xnor U32873 (N_32873,N_30417,N_31347);
or U32874 (N_32874,N_30045,N_32017);
nor U32875 (N_32875,N_32454,N_30860);
nor U32876 (N_32876,N_30746,N_31062);
xnor U32877 (N_32877,N_31879,N_32075);
or U32878 (N_32878,N_30955,N_32262);
nor U32879 (N_32879,N_30467,N_32379);
nor U32880 (N_32880,N_31289,N_32289);
nor U32881 (N_32881,N_30604,N_30495);
xnor U32882 (N_32882,N_30620,N_32158);
nand U32883 (N_32883,N_31251,N_30533);
and U32884 (N_32884,N_32052,N_31135);
xor U32885 (N_32885,N_30719,N_31454);
and U32886 (N_32886,N_31230,N_30158);
and U32887 (N_32887,N_31877,N_31591);
nand U32888 (N_32888,N_30408,N_31840);
nand U32889 (N_32889,N_30312,N_32434);
nand U32890 (N_32890,N_30856,N_32317);
nor U32891 (N_32891,N_31272,N_31463);
nand U32892 (N_32892,N_30817,N_31376);
or U32893 (N_32893,N_30396,N_32465);
xor U32894 (N_32894,N_31935,N_32395);
nand U32895 (N_32895,N_31423,N_31697);
nand U32896 (N_32896,N_31175,N_30191);
xor U32897 (N_32897,N_30485,N_30160);
and U32898 (N_32898,N_31993,N_30073);
or U32899 (N_32899,N_32046,N_32219);
nand U32900 (N_32900,N_32224,N_32074);
nand U32901 (N_32901,N_31352,N_30938);
or U32902 (N_32902,N_30960,N_30882);
xnor U32903 (N_32903,N_31820,N_30369);
xnor U32904 (N_32904,N_31782,N_31477);
or U32905 (N_32905,N_31157,N_30042);
or U32906 (N_32906,N_32202,N_31983);
and U32907 (N_32907,N_32494,N_32025);
or U32908 (N_32908,N_31061,N_31481);
or U32909 (N_32909,N_31649,N_32303);
nand U32910 (N_32910,N_30636,N_32174);
or U32911 (N_32911,N_30269,N_31765);
or U32912 (N_32912,N_31059,N_32113);
nor U32913 (N_32913,N_30290,N_31693);
nand U32914 (N_32914,N_30616,N_31183);
and U32915 (N_32915,N_30116,N_31932);
nor U32916 (N_32916,N_30855,N_32455);
nor U32917 (N_32917,N_30461,N_31244);
nor U32918 (N_32918,N_30685,N_30224);
xnor U32919 (N_32919,N_32037,N_30740);
nor U32920 (N_32920,N_32098,N_31992);
or U32921 (N_32921,N_31424,N_30303);
or U32922 (N_32922,N_31367,N_31327);
nor U32923 (N_32923,N_31633,N_32297);
or U32924 (N_32924,N_31077,N_30139);
nand U32925 (N_32925,N_30657,N_30259);
nand U32926 (N_32926,N_31805,N_31750);
and U32927 (N_32927,N_32263,N_31808);
and U32928 (N_32928,N_32122,N_31375);
nand U32929 (N_32929,N_31857,N_31828);
nand U32930 (N_32930,N_30607,N_30201);
xnor U32931 (N_32931,N_31610,N_31312);
nor U32932 (N_32932,N_31052,N_32009);
or U32933 (N_32933,N_30310,N_30940);
nand U32934 (N_32934,N_30725,N_32332);
or U32935 (N_32935,N_30511,N_31919);
xor U32936 (N_32936,N_31672,N_31296);
nand U32937 (N_32937,N_32191,N_30837);
nand U32938 (N_32938,N_30577,N_32227);
xnor U32939 (N_32939,N_30665,N_30082);
or U32940 (N_32940,N_31880,N_30741);
nand U32941 (N_32941,N_31263,N_31385);
nor U32942 (N_32942,N_31971,N_30272);
xnor U32943 (N_32943,N_31169,N_30230);
and U32944 (N_32944,N_32028,N_30252);
nand U32945 (N_32945,N_31977,N_30088);
nor U32946 (N_32946,N_31227,N_31330);
or U32947 (N_32947,N_31131,N_30462);
nand U32948 (N_32948,N_32030,N_32312);
and U32949 (N_32949,N_31074,N_30929);
and U32950 (N_32950,N_31110,N_32061);
nand U32951 (N_32951,N_31133,N_30043);
or U32952 (N_32952,N_32119,N_30262);
or U32953 (N_32953,N_30013,N_31613);
nand U32954 (N_32954,N_31511,N_30069);
or U32955 (N_32955,N_32443,N_31888);
and U32956 (N_32956,N_31594,N_31149);
nor U32957 (N_32957,N_30972,N_30884);
xor U32958 (N_32958,N_31191,N_30721);
nor U32959 (N_32959,N_31548,N_30380);
and U32960 (N_32960,N_31867,N_30446);
or U32961 (N_32961,N_30238,N_31196);
xnor U32962 (N_32962,N_31410,N_30670);
or U32963 (N_32963,N_32015,N_30249);
and U32964 (N_32964,N_32192,N_30539);
nor U32965 (N_32965,N_31245,N_30836);
nand U32966 (N_32966,N_31146,N_31837);
or U32967 (N_32967,N_30004,N_30824);
nor U32968 (N_32968,N_30076,N_30538);
nor U32969 (N_32969,N_31171,N_30049);
nand U32970 (N_32970,N_31902,N_30305);
xor U32971 (N_32971,N_30664,N_32103);
xor U32972 (N_32972,N_30356,N_30372);
nor U32973 (N_32973,N_30815,N_31095);
or U32974 (N_32974,N_30080,N_32345);
nor U32975 (N_32975,N_31841,N_32110);
nor U32976 (N_32976,N_32414,N_30536);
nand U32977 (N_32977,N_30371,N_31553);
nand U32978 (N_32978,N_31179,N_31568);
or U32979 (N_32979,N_31260,N_32045);
nor U32980 (N_32980,N_31595,N_30808);
and U32981 (N_32981,N_30771,N_31236);
nor U32982 (N_32982,N_30599,N_30329);
and U32983 (N_32983,N_30827,N_30111);
nor U32984 (N_32984,N_31428,N_30246);
and U32985 (N_32985,N_31999,N_30445);
and U32986 (N_32986,N_30914,N_30008);
xnor U32987 (N_32987,N_31010,N_30021);
nor U32988 (N_32988,N_30715,N_30386);
xnor U32989 (N_32989,N_32424,N_31646);
xnor U32990 (N_32990,N_30546,N_32378);
xnor U32991 (N_32991,N_31600,N_30734);
nand U32992 (N_32992,N_31753,N_30353);
or U32993 (N_32993,N_30624,N_30019);
xor U32994 (N_32994,N_32236,N_30561);
nor U32995 (N_32995,N_30095,N_30437);
nand U32996 (N_32996,N_31843,N_31663);
nand U32997 (N_32997,N_32388,N_31339);
nor U32998 (N_32998,N_30271,N_30613);
and U32999 (N_32999,N_30425,N_32121);
nand U33000 (N_33000,N_32133,N_30367);
xor U33001 (N_33001,N_31795,N_31405);
and U33002 (N_33002,N_31318,N_31550);
xnor U33003 (N_33003,N_31100,N_30442);
nor U33004 (N_33004,N_30167,N_30590);
xnor U33005 (N_33005,N_30016,N_31053);
and U33006 (N_33006,N_30679,N_31396);
or U33007 (N_33007,N_32363,N_30322);
and U33008 (N_33008,N_32007,N_31329);
nor U33009 (N_33009,N_30274,N_30317);
and U33010 (N_33010,N_31239,N_32389);
and U33011 (N_33011,N_30291,N_30267);
xor U33012 (N_33012,N_30933,N_32112);
or U33013 (N_33013,N_32196,N_31732);
or U33014 (N_33014,N_30411,N_31213);
nand U33015 (N_33015,N_32168,N_31364);
nand U33016 (N_33016,N_30531,N_32301);
and U33017 (N_33017,N_31758,N_31789);
nand U33018 (N_33018,N_30268,N_31684);
nand U33019 (N_33019,N_30992,N_31409);
nor U33020 (N_33020,N_31268,N_31011);
or U33021 (N_33021,N_31786,N_30925);
and U33022 (N_33022,N_32205,N_31872);
or U33023 (N_33023,N_30649,N_30451);
xnor U33024 (N_33024,N_31308,N_32076);
nand U33025 (N_33025,N_31749,N_30775);
and U33026 (N_33026,N_32246,N_31892);
and U33027 (N_33027,N_30515,N_30762);
nor U33028 (N_33028,N_30705,N_32108);
or U33029 (N_33029,N_32014,N_30025);
or U33030 (N_33030,N_31018,N_31894);
xor U33031 (N_33031,N_31647,N_31968);
and U33032 (N_33032,N_31944,N_30708);
nor U33033 (N_33033,N_30345,N_30330);
nand U33034 (N_33034,N_30118,N_32012);
or U33035 (N_33035,N_30713,N_32492);
xnor U33036 (N_33036,N_31955,N_32373);
or U33037 (N_33037,N_32447,N_31848);
nor U33038 (N_33038,N_30774,N_32056);
and U33039 (N_33039,N_30693,N_31699);
nor U33040 (N_33040,N_31582,N_31519);
xnor U33041 (N_33041,N_30658,N_31503);
nand U33042 (N_33042,N_30936,N_31014);
or U33043 (N_33043,N_30971,N_30654);
nand U33044 (N_33044,N_31544,N_30700);
nand U33045 (N_33045,N_30573,N_31034);
or U33046 (N_33046,N_31670,N_30786);
xor U33047 (N_33047,N_32184,N_31009);
and U33048 (N_33048,N_32077,N_30198);
nor U33049 (N_33049,N_31886,N_31022);
nand U33050 (N_33050,N_31514,N_30079);
nor U33051 (N_33051,N_32497,N_31277);
or U33052 (N_33052,N_31371,N_30393);
nor U33053 (N_33053,N_31884,N_31482);
nand U33054 (N_33054,N_30175,N_30208);
nor U33055 (N_33055,N_31097,N_30754);
and U33056 (N_33056,N_32210,N_31091);
xnor U33057 (N_33057,N_30739,N_31406);
nand U33058 (N_33058,N_31696,N_31012);
xor U33059 (N_33059,N_32136,N_31887);
and U33060 (N_33060,N_31039,N_31160);
nor U33061 (N_33061,N_32468,N_32368);
and U33062 (N_33062,N_30357,N_31126);
and U33063 (N_33063,N_30828,N_32070);
nor U33064 (N_33064,N_31162,N_31873);
nor U33065 (N_33065,N_32139,N_30551);
and U33066 (N_33066,N_30137,N_32230);
xor U33067 (N_33067,N_30687,N_31415);
and U33068 (N_33068,N_31899,N_30660);
xnor U33069 (N_33069,N_31075,N_31564);
or U33070 (N_33070,N_32484,N_31072);
nand U33071 (N_33071,N_30419,N_30146);
nor U33072 (N_33072,N_32131,N_31916);
or U33073 (N_33073,N_31209,N_31604);
xnor U33074 (N_33074,N_30563,N_30211);
and U33075 (N_33075,N_31471,N_32340);
nand U33076 (N_33076,N_32400,N_31082);
or U33077 (N_33077,N_31942,N_31615);
or U33078 (N_33078,N_30789,N_30548);
or U33079 (N_33079,N_30592,N_30491);
or U33080 (N_33080,N_30500,N_31345);
and U33081 (N_33081,N_31810,N_31462);
nor U33082 (N_33082,N_30407,N_32033);
nand U33083 (N_33083,N_30578,N_30338);
and U33084 (N_33084,N_31319,N_30557);
nand U33085 (N_33085,N_32031,N_31321);
and U33086 (N_33086,N_30409,N_31678);
and U33087 (N_33087,N_30289,N_32453);
and U33088 (N_33088,N_32176,N_31928);
nor U33089 (N_33089,N_30973,N_31769);
xnor U33090 (N_33090,N_30061,N_30642);
nor U33091 (N_33091,N_30645,N_31393);
nor U33092 (N_33092,N_30669,N_30597);
or U33093 (N_33093,N_30562,N_30611);
nand U33094 (N_33094,N_31787,N_31596);
xor U33095 (N_33095,N_31933,N_30617);
and U33096 (N_33096,N_31761,N_30420);
or U33097 (N_33097,N_31845,N_31963);
xnor U33098 (N_33098,N_31282,N_30328);
xnor U33099 (N_33099,N_30142,N_31577);
and U33100 (N_33100,N_30627,N_32338);
and U33101 (N_33101,N_30820,N_31987);
or U33102 (N_33102,N_30748,N_32245);
or U33103 (N_33103,N_31953,N_30532);
nand U33104 (N_33104,N_31856,N_30945);
xnor U33105 (N_33105,N_30998,N_31498);
or U33106 (N_33106,N_31698,N_32055);
nor U33107 (N_33107,N_30926,N_30981);
and U33108 (N_33108,N_31949,N_30977);
or U33109 (N_33109,N_30340,N_32362);
or U33110 (N_33110,N_31299,N_31551);
or U33111 (N_33111,N_31473,N_32485);
xor U33112 (N_33112,N_31814,N_30630);
or U33113 (N_33113,N_30758,N_30638);
and U33114 (N_33114,N_31207,N_31984);
nor U33115 (N_33115,N_30352,N_30226);
xor U33116 (N_33116,N_30502,N_32393);
or U33117 (N_33117,N_32318,N_30248);
and U33118 (N_33118,N_30178,N_31003);
xor U33119 (N_33119,N_30986,N_32476);
and U33120 (N_33120,N_32124,N_30285);
and U33121 (N_33121,N_30544,N_32307);
or U33122 (N_33122,N_32324,N_30266);
or U33123 (N_33123,N_31812,N_30838);
or U33124 (N_33124,N_31764,N_31565);
xnor U33125 (N_33125,N_32058,N_32253);
xor U33126 (N_33126,N_31331,N_31501);
and U33127 (N_33127,N_32034,N_31939);
nor U33128 (N_33128,N_32085,N_32198);
and U33129 (N_33129,N_32477,N_30735);
nand U33130 (N_33130,N_32232,N_30331);
xnor U33131 (N_33131,N_30618,N_31771);
or U33132 (N_33132,N_30534,N_30908);
and U33133 (N_33133,N_30853,N_32452);
xnor U33134 (N_33134,N_31337,N_30232);
and U33135 (N_33135,N_30212,N_31286);
nor U33136 (N_33136,N_31831,N_30200);
and U33137 (N_33137,N_31069,N_31145);
and U33138 (N_33138,N_31168,N_31518);
nor U33139 (N_33139,N_32310,N_30805);
or U33140 (N_33140,N_30363,N_31192);
xor U33141 (N_33141,N_30891,N_30772);
and U33142 (N_33142,N_30017,N_31271);
or U33143 (N_33143,N_32410,N_30537);
nand U33144 (N_33144,N_31683,N_32290);
nor U33145 (N_33145,N_30760,N_32093);
and U33146 (N_33146,N_31959,N_31025);
xor U33147 (N_33147,N_31120,N_31125);
nand U33148 (N_33148,N_31013,N_30250);
xnor U33149 (N_33149,N_30675,N_32488);
or U33150 (N_33150,N_32432,N_31143);
and U33151 (N_33151,N_30253,N_30997);
nor U33152 (N_33152,N_31825,N_31087);
nand U33153 (N_33153,N_30849,N_30487);
or U33154 (N_33154,N_31730,N_31815);
or U33155 (N_33155,N_30421,N_31527);
nor U33156 (N_33156,N_30931,N_30123);
nor U33157 (N_33157,N_32068,N_31796);
nor U33158 (N_33158,N_31280,N_30785);
nor U33159 (N_33159,N_30886,N_31046);
or U33160 (N_33160,N_30979,N_30318);
nand U33161 (N_33161,N_30869,N_31449);
xnor U33162 (N_33162,N_31178,N_31803);
nor U33163 (N_33163,N_31112,N_31708);
and U33164 (N_33164,N_31525,N_31391);
nor U33165 (N_33165,N_31996,N_30447);
nor U33166 (N_33166,N_30605,N_32188);
or U33167 (N_33167,N_31252,N_30773);
nand U33168 (N_33168,N_31601,N_30436);
nor U33169 (N_33169,N_31861,N_30904);
nand U33170 (N_33170,N_31353,N_32194);
nor U33171 (N_33171,N_30458,N_31547);
nand U33172 (N_33172,N_31247,N_31917);
nand U33173 (N_33173,N_30479,N_32352);
xnor U33174 (N_33174,N_31249,N_30336);
or U33175 (N_33175,N_31314,N_30078);
nor U33176 (N_33176,N_31806,N_30880);
and U33177 (N_33177,N_31807,N_32293);
nor U33178 (N_33178,N_31834,N_32220);
nor U33179 (N_33179,N_30030,N_30294);
or U33180 (N_33180,N_31874,N_30140);
or U33181 (N_33181,N_30800,N_30930);
or U33182 (N_33182,N_31043,N_31976);
and U33183 (N_33183,N_30492,N_30168);
nand U33184 (N_33184,N_31661,N_32054);
nor U33185 (N_33185,N_32060,N_30454);
xnor U33186 (N_33186,N_30542,N_31811);
nand U33187 (N_33187,N_31079,N_31729);
xor U33188 (N_33188,N_31901,N_30519);
xor U33189 (N_33189,N_32319,N_30947);
and U33190 (N_33190,N_31246,N_31988);
nor U33191 (N_33191,N_31626,N_30711);
xor U33192 (N_33192,N_30728,N_30359);
nand U33193 (N_33193,N_31015,N_31458);
nor U33194 (N_33194,N_31488,N_30576);
or U33195 (N_33195,N_32458,N_30464);
xnor U33196 (N_33196,N_32456,N_31865);
and U33197 (N_33197,N_30545,N_30799);
or U33198 (N_33198,N_31363,N_30489);
nand U33199 (N_33199,N_30680,N_31760);
nor U33200 (N_33200,N_32020,N_31343);
nand U33201 (N_33201,N_31373,N_30337);
nor U33202 (N_33202,N_31468,N_31431);
nand U33203 (N_33203,N_30423,N_30147);
nand U33204 (N_33204,N_30535,N_30565);
nand U33205 (N_33205,N_30987,N_31538);
nor U33206 (N_33206,N_30251,N_31181);
or U33207 (N_33207,N_31258,N_30759);
and U33208 (N_33208,N_32449,N_30498);
xnor U33209 (N_33209,N_32067,N_31668);
and U33210 (N_33210,N_30388,N_32386);
nand U33211 (N_33211,N_31688,N_32157);
nor U33212 (N_33212,N_32311,N_31232);
nor U33213 (N_33213,N_30801,N_30052);
or U33214 (N_33214,N_30130,N_31264);
nand U33215 (N_33215,N_30549,N_31122);
nand U33216 (N_33216,N_31453,N_31257);
and U33217 (N_33217,N_31883,N_32413);
xor U33218 (N_33218,N_32049,N_32280);
or U33219 (N_33219,N_31997,N_31113);
nor U33220 (N_33220,N_31657,N_30089);
nand U33221 (N_33221,N_32149,N_32419);
nor U33222 (N_33222,N_32170,N_30683);
nand U33223 (N_33223,N_31864,N_31938);
nand U33224 (N_33224,N_31711,N_30939);
xor U33225 (N_33225,N_30100,N_30859);
nor U33226 (N_33226,N_31340,N_32091);
and U33227 (N_33227,N_30848,N_30047);
and U33228 (N_33228,N_30194,N_30575);
nand U33229 (N_33229,N_31354,N_31915);
and U33230 (N_33230,N_30870,N_32428);
xnor U33231 (N_33231,N_30006,N_30392);
nor U33232 (N_33232,N_32137,N_32005);
or U33233 (N_33233,N_30264,N_30020);
or U33234 (N_33234,N_31383,N_31598);
and U33235 (N_33235,N_31253,N_31334);
nand U33236 (N_33236,N_32409,N_30127);
nor U33237 (N_33237,N_32029,N_30165);
and U33238 (N_33238,N_30832,N_30125);
and U33239 (N_33239,N_32057,N_31123);
or U33240 (N_33240,N_32003,N_30415);
nand U33241 (N_33241,N_32241,N_31995);
nand U33242 (N_33242,N_30022,N_32346);
and U33243 (N_33243,N_31050,N_32406);
nor U33244 (N_33244,N_30074,N_31715);
and U33245 (N_33245,N_31108,N_31706);
nor U33246 (N_33246,N_30995,N_30107);
and U33247 (N_33247,N_31589,N_30659);
nor U33248 (N_33248,N_31040,N_31114);
nand U33249 (N_33249,N_31116,N_32144);
and U33250 (N_33250,N_31722,N_32334);
nor U33251 (N_33251,N_30781,N_30816);
or U33252 (N_33252,N_30582,N_31184);
and U33253 (N_33253,N_30932,N_32216);
xor U33254 (N_33254,N_31536,N_31890);
nor U33255 (N_33255,N_30883,N_31210);
or U33256 (N_33256,N_32010,N_30806);
and U33257 (N_33257,N_30081,N_31623);
xnor U33258 (N_33258,N_30375,N_32493);
nand U33259 (N_33259,N_30512,N_31198);
nor U33260 (N_33260,N_30915,N_32231);
xnor U33261 (N_33261,N_31237,N_31763);
xnor U33262 (N_33262,N_31905,N_31254);
and U33263 (N_33263,N_31044,N_31773);
and U33264 (N_33264,N_30833,N_32138);
and U33265 (N_33265,N_32425,N_31094);
nand U33266 (N_33266,N_30543,N_31480);
and U33267 (N_33267,N_31486,N_31243);
or U33268 (N_33268,N_31217,N_31830);
or U33269 (N_33269,N_30349,N_32114);
or U33270 (N_33270,N_31576,N_30192);
nand U33271 (N_33271,N_30263,N_32274);
xor U33272 (N_33272,N_31687,N_30547);
nor U33273 (N_33273,N_30527,N_32408);
or U33274 (N_33274,N_31380,N_31783);
xnor U33275 (N_33275,N_32462,N_31751);
or U33276 (N_33276,N_31404,N_31200);
xor U33277 (N_33277,N_30277,N_30608);
and U33278 (N_33278,N_32249,N_30514);
nor U33279 (N_33279,N_30821,N_30651);
xnor U33280 (N_33280,N_30105,N_31138);
or U33281 (N_33281,N_30433,N_31580);
nand U33282 (N_33282,N_32177,N_30484);
or U33283 (N_33283,N_30593,N_30610);
or U33284 (N_33284,N_32296,N_30631);
nand U33285 (N_33285,N_31797,N_30878);
nor U33286 (N_33286,N_32063,N_30643);
and U33287 (N_33287,N_31342,N_31740);
or U33288 (N_33288,N_30469,N_30075);
nor U33289 (N_33289,N_30002,N_32283);
nand U33290 (N_33290,N_32358,N_31602);
xnor U33291 (N_33291,N_32000,N_30378);
nand U33292 (N_33292,N_31316,N_30077);
and U33293 (N_33293,N_31464,N_30698);
or U33294 (N_33294,N_31444,N_31491);
or U33295 (N_33295,N_32256,N_30196);
nor U33296 (N_33296,N_31320,N_31827);
nand U33297 (N_33297,N_31710,N_30255);
or U33298 (N_33298,N_30185,N_30894);
and U33299 (N_33299,N_30171,N_30726);
nand U33300 (N_33300,N_31632,N_31676);
nand U33301 (N_33301,N_31238,N_30024);
nor U33302 (N_33302,N_31813,N_32084);
or U33303 (N_33303,N_31714,N_30098);
nand U33304 (N_33304,N_32050,N_32384);
xor U33305 (N_33305,N_30379,N_30390);
or U33306 (N_33306,N_31068,N_32329);
nor U33307 (N_33307,N_31297,N_30028);
nand U33308 (N_33308,N_31433,N_31466);
and U33309 (N_33309,N_32258,N_31256);
and U33310 (N_33310,N_32435,N_31648);
and U33311 (N_33311,N_32325,N_30732);
xnor U33312 (N_33312,N_30552,N_30598);
nor U33313 (N_33313,N_32260,N_32161);
nand U33314 (N_33314,N_31092,N_31066);
xnor U33315 (N_33315,N_31324,N_30057);
xor U33316 (N_33316,N_30159,N_30901);
and U33317 (N_33317,N_32459,N_30928);
xor U33318 (N_33318,N_30347,N_31677);
and U33319 (N_33319,N_30949,N_30135);
and U33320 (N_33320,N_31164,N_30691);
or U33321 (N_33321,N_30639,N_31024);
nor U33322 (N_33322,N_31513,N_30872);
nor U33323 (N_33323,N_30400,N_32344);
nor U33324 (N_33324,N_32006,N_30444);
or U33325 (N_33325,N_30779,N_30062);
and U33326 (N_33326,N_30656,N_31419);
or U33327 (N_33327,N_32222,N_31174);
nand U33328 (N_33328,N_30221,N_31967);
nand U33329 (N_33329,N_30695,N_31964);
nand U33330 (N_33330,N_31315,N_31889);
xor U33331 (N_33331,N_32062,N_30236);
nand U33332 (N_33332,N_31495,N_30733);
or U33333 (N_33333,N_30962,N_30243);
xor U33334 (N_33334,N_30684,N_30083);
nor U33335 (N_33335,N_30867,N_31291);
nand U33336 (N_33336,N_30051,N_30148);
nand U33337 (N_33337,N_30888,N_32155);
and U33338 (N_33338,N_32356,N_30382);
nand U33339 (N_33339,N_32489,N_31017);
or U33340 (N_33340,N_30776,N_30807);
xor U33341 (N_33341,N_30877,N_31429);
and U33342 (N_33342,N_30994,N_32496);
nand U33343 (N_33343,N_32269,N_30963);
nor U33344 (N_33344,N_31294,N_30270);
nor U33345 (N_33345,N_32355,N_31201);
and U33346 (N_33346,N_32353,N_32481);
xnor U33347 (N_33347,N_31496,N_31954);
or U33348 (N_33348,N_30122,N_31784);
and U33349 (N_33349,N_30326,N_31096);
or U33350 (N_33350,N_31636,N_31985);
or U33351 (N_33351,N_31084,N_30067);
nand U33352 (N_33352,N_31248,N_32234);
xnor U33353 (N_33353,N_30873,N_31416);
or U33354 (N_33354,N_31452,N_32291);
xor U33355 (N_33355,N_31156,N_32154);
xnor U33356 (N_33356,N_31835,N_30861);
nand U33357 (N_33357,N_31033,N_30273);
nor U33358 (N_33358,N_30678,N_32273);
xor U33359 (N_33359,N_30483,N_30044);
and U33360 (N_33360,N_31436,N_30333);
and U33361 (N_33361,N_30927,N_32391);
nand U33362 (N_33362,N_31639,N_30846);
and U33363 (N_33363,N_30952,N_30574);
or U33364 (N_33364,N_30770,N_31660);
and U33365 (N_33365,N_30422,N_30394);
nor U33366 (N_33366,N_30964,N_31945);
and U33367 (N_33367,N_31350,N_32048);
nor U33368 (N_33368,N_30335,N_31398);
nor U33369 (N_33369,N_31332,N_31479);
or U33370 (N_33370,N_30982,N_30959);
xnor U33371 (N_33371,N_30595,N_30453);
xor U33372 (N_33372,N_30793,N_31743);
xor U33373 (N_33373,N_31555,N_31064);
xor U33374 (N_33374,N_31809,N_30320);
nor U33375 (N_33375,N_32019,N_30526);
nor U33376 (N_33376,N_31266,N_30556);
and U33377 (N_33377,N_31418,N_32351);
nand U33378 (N_33378,N_31388,N_31132);
xnor U33379 (N_33379,N_32431,N_31042);
and U33380 (N_33380,N_32169,N_31067);
or U33381 (N_33381,N_31369,N_30513);
nor U33382 (N_33382,N_31898,N_31875);
nor U33383 (N_33383,N_30673,N_31969);
or U33384 (N_33384,N_32004,N_31869);
nor U33385 (N_33385,N_32390,N_31130);
xnor U33386 (N_33386,N_31966,N_31121);
and U33387 (N_33387,N_31788,N_30163);
xor U33388 (N_33388,N_30553,N_32267);
or U33389 (N_33389,N_31115,N_32147);
nand U33390 (N_33390,N_31494,N_30063);
nor U33391 (N_33391,N_30841,N_30706);
nand U33392 (N_33392,N_31222,N_31962);
nand U33393 (N_33393,N_31509,N_31356);
nand U33394 (N_33394,N_31946,N_30629);
xor U33395 (N_33395,N_32382,N_31630);
and U33396 (N_33396,N_32172,N_32320);
nand U33397 (N_33397,N_30302,N_31137);
or U33398 (N_33398,N_30070,N_30119);
and U33399 (N_33399,N_30457,N_31529);
nand U33400 (N_33400,N_31300,N_31206);
and U33401 (N_33401,N_30897,N_30490);
or U33402 (N_33402,N_31520,N_31021);
nand U33403 (N_33403,N_31153,N_31695);
or U33404 (N_33404,N_31080,N_30315);
and U33405 (N_33405,N_31159,N_31990);
or U33406 (N_33406,N_31309,N_31276);
xor U33407 (N_33407,N_31446,N_31189);
and U33408 (N_33408,N_31721,N_31778);
xor U33409 (N_33409,N_31152,N_30749);
and U33410 (N_33410,N_30520,N_32100);
xor U33411 (N_33411,N_32073,N_30284);
nor U33412 (N_33412,N_30210,N_31680);
nor U33413 (N_33413,N_32018,N_31768);
or U33414 (N_33414,N_30432,N_30032);
or U33415 (N_33415,N_31492,N_32463);
nor U33416 (N_33416,N_31818,N_32417);
and U33417 (N_33417,N_30798,N_31355);
nand U33418 (N_33418,N_31055,N_31603);
and U33419 (N_33419,N_30239,N_31139);
nor U33420 (N_33420,N_30041,N_30965);
and U33421 (N_33421,N_31566,N_31723);
and U33422 (N_33422,N_31357,N_30414);
xor U33423 (N_33423,N_30953,N_31279);
and U33424 (N_33424,N_30835,N_31543);
or U33425 (N_33425,N_30505,N_32195);
or U33426 (N_33426,N_30348,N_31885);
xnor U33427 (N_33427,N_32339,N_31720);
xnor U33428 (N_33428,N_32498,N_30283);
xor U33429 (N_33429,N_32277,N_31117);
xor U33430 (N_33430,N_30989,N_32316);
nand U33431 (N_33431,N_31104,N_31098);
and U33432 (N_33432,N_31658,N_31058);
or U33433 (N_33433,N_30141,N_30572);
and U33434 (N_33434,N_30110,N_30093);
nor U33435 (N_33435,N_32143,N_31754);
nand U33436 (N_33436,N_31718,N_30026);
and U33437 (N_33437,N_31667,N_32336);
nand U33438 (N_33438,N_30014,N_30588);
or U33439 (N_33439,N_32148,N_32164);
and U33440 (N_33440,N_32491,N_32471);
nor U33441 (N_33441,N_30377,N_30716);
nor U33442 (N_33442,N_32087,N_31401);
or U33443 (N_33443,N_30622,N_31229);
nand U33444 (N_33444,N_32466,N_31031);
or U33445 (N_33445,N_32369,N_32472);
or U33446 (N_33446,N_30339,N_31459);
and U33447 (N_33447,N_30493,N_30525);
nand U33448 (N_33448,N_31147,N_32314);
or U33449 (N_33449,N_31425,N_30787);
and U33450 (N_33450,N_31512,N_31158);
or U33451 (N_33451,N_30354,N_31694);
or U33452 (N_33452,N_30819,N_30690);
and U33453 (N_33453,N_32072,N_31301);
nand U33454 (N_33454,N_32242,N_32328);
or U33455 (N_33455,N_30346,N_32292);
nand U33456 (N_33456,N_30851,N_31302);
nand U33457 (N_33457,N_32206,N_30893);
nor U33458 (N_33458,N_32407,N_30245);
nor U33459 (N_33459,N_31119,N_32171);
and U33460 (N_33460,N_30155,N_32229);
and U33461 (N_33461,N_30842,N_31506);
nand U33462 (N_33462,N_32099,N_30934);
or U33463 (N_33463,N_30619,N_30452);
and U33464 (N_33464,N_31349,N_31535);
and U33465 (N_33465,N_32095,N_31643);
nand U33466 (N_33466,N_31127,N_32376);
and U33467 (N_33467,N_31233,N_30166);
nand U33468 (N_33468,N_30299,N_30969);
nand U33469 (N_33469,N_32130,N_31844);
or U33470 (N_33470,N_31819,N_30755);
nand U33471 (N_33471,N_32038,N_30441);
nor U33472 (N_33472,N_31824,N_30465);
nand U33473 (N_33473,N_30913,N_31167);
and U33474 (N_33474,N_30890,N_30071);
and U33475 (N_33475,N_31833,N_31148);
or U33476 (N_33476,N_31734,N_32337);
nor U33477 (N_33477,N_31522,N_31386);
nand U33478 (N_33478,N_30990,N_31447);
and U33479 (N_33479,N_32357,N_30792);
and U33480 (N_33480,N_31731,N_32102);
nor U33481 (N_33481,N_30301,N_31717);
nand U33482 (N_33482,N_31170,N_31839);
xnor U33483 (N_33483,N_31641,N_31045);
and U33484 (N_33484,N_31372,N_30406);
xor U33485 (N_33485,N_31389,N_31504);
xnor U33486 (N_33486,N_32248,N_31970);
or U33487 (N_33487,N_32212,N_31930);
nand U33488 (N_33488,N_30482,N_31193);
and U33489 (N_33489,N_32420,N_31823);
and U33490 (N_33490,N_31054,N_32315);
or U33491 (N_33491,N_30470,N_32039);
and U33492 (N_33492,N_32002,N_30822);
nor U33493 (N_33493,N_31791,N_32200);
nand U33494 (N_33494,N_31986,N_30187);
or U33495 (N_33495,N_31395,N_32105);
xnor U33496 (N_33496,N_31442,N_31635);
and U33497 (N_33497,N_31411,N_30297);
and U33498 (N_33498,N_31390,N_31585);
nor U33499 (N_33499,N_32295,N_30723);
nor U33500 (N_33500,N_32437,N_30875);
xnor U33501 (N_33501,N_30707,N_30217);
and U33502 (N_33502,N_31365,N_31586);
nor U33503 (N_33503,N_31756,N_30478);
nor U33504 (N_33504,N_32066,N_31288);
or U33505 (N_33505,N_32495,N_30996);
and U33506 (N_33506,N_32204,N_30086);
or U33507 (N_33507,N_32348,N_32427);
xnor U33508 (N_33508,N_32451,N_32197);
xnor U33509 (N_33509,N_31799,N_32367);
or U33510 (N_33510,N_31838,N_30058);
nand U33511 (N_33511,N_31231,N_31920);
and U33512 (N_33512,N_31606,N_32140);
nor U33513 (N_33513,N_30881,N_30825);
or U33514 (N_33514,N_30688,N_32211);
or U33515 (N_33515,N_30199,N_32126);
or U33516 (N_33516,N_31973,N_31650);
or U33517 (N_33517,N_31027,N_30587);
xnor U33518 (N_33518,N_32396,N_32254);
or U33519 (N_33519,N_30475,N_30942);
nor U33520 (N_33520,N_31508,N_32330);
and U33521 (N_33521,N_32104,N_31654);
nand U33522 (N_33522,N_31690,N_31801);
xor U33523 (N_33523,N_32482,N_31571);
or U33524 (N_33524,N_31952,N_30223);
or U33525 (N_33525,N_32132,N_31631);
nor U33526 (N_33526,N_32250,N_32135);
nand U33527 (N_33527,N_31325,N_30530);
or U33528 (N_33528,N_32181,N_31908);
xor U33529 (N_33529,N_32261,N_31860);
nor U33530 (N_33530,N_30413,N_30341);
xor U33531 (N_33531,N_31421,N_30879);
nand U33532 (N_33532,N_31456,N_32117);
and U33533 (N_33533,N_31507,N_30162);
and U33534 (N_33534,N_31850,N_31752);
and U33535 (N_33535,N_30207,N_30040);
nand U33536 (N_33536,N_30126,N_31487);
nor U33537 (N_33537,N_31399,N_31541);
nand U33538 (N_33538,N_31575,N_31616);
nand U33539 (N_33539,N_31614,N_30306);
nor U33540 (N_33540,N_32321,N_30769);
xor U33541 (N_33541,N_31863,N_30903);
xor U33542 (N_33542,N_32259,N_31979);
nor U33543 (N_33543,N_31026,N_30048);
xnor U33544 (N_33544,N_31619,N_32421);
and U33545 (N_33545,N_32233,N_32223);
or U33546 (N_33546,N_31047,N_32101);
and U33547 (N_33547,N_30342,N_31060);
nand U33548 (N_33548,N_32128,N_30287);
nor U33549 (N_33549,N_31656,N_30494);
nand U33550 (N_33550,N_31150,N_30066);
nand U33551 (N_33551,N_31640,N_31662);
nor U33552 (N_33552,N_30826,N_32214);
and U33553 (N_33553,N_31284,N_30254);
xor U33554 (N_33554,N_31852,N_31199);
and U33555 (N_33555,N_31467,N_30830);
nand U33556 (N_33556,N_31234,N_30743);
or U33557 (N_33557,N_32309,N_30468);
nand U33558 (N_33558,N_30594,N_31472);
nand U33559 (N_33559,N_30803,N_31028);
nand U33560 (N_33560,N_30156,N_31583);
or U33561 (N_33561,N_30844,N_32398);
nand U33562 (N_33562,N_31448,N_30247);
or U33563 (N_33563,N_31101,N_31381);
or U33564 (N_33564,N_32342,N_31049);
nand U33565 (N_33565,N_30951,N_31870);
nor U33566 (N_33566,N_30497,N_30661);
and U33567 (N_33567,N_30143,N_31226);
and U33568 (N_33568,N_31417,N_31377);
nor U33569 (N_33569,N_30242,N_32190);
or U33570 (N_33570,N_32285,N_31407);
and U33571 (N_33571,N_30096,N_30727);
or U33572 (N_33572,N_31532,N_31261);
or U33573 (N_33573,N_32365,N_31826);
nand U33574 (N_33574,N_31265,N_30173);
or U33575 (N_33575,N_32180,N_30950);
xor U33576 (N_33576,N_31326,N_32473);
nand U33577 (N_33577,N_30334,N_30193);
nand U33578 (N_33578,N_31956,N_30559);
nor U33579 (N_33579,N_30862,N_30459);
or U33580 (N_33580,N_31020,N_31560);
or U33581 (N_33581,N_30144,N_30944);
and U33582 (N_33582,N_30634,N_30011);
xnor U33583 (N_33583,N_31748,N_30921);
nand U33584 (N_33584,N_31597,N_31804);
nand U33585 (N_33585,N_31629,N_30644);
xor U33586 (N_33586,N_31262,N_31652);
xnor U33587 (N_33587,N_30674,N_30220);
nor U33588 (N_33588,N_30298,N_31303);
nor U33589 (N_33589,N_30037,N_31628);
nor U33590 (N_33590,N_32487,N_31346);
or U33591 (N_33591,N_30797,N_31924);
nand U33592 (N_33592,N_30701,N_30324);
or U33593 (N_33593,N_32490,N_32083);
xor U33594 (N_33594,N_32270,N_30179);
or U33595 (N_33595,N_30440,N_31412);
nand U33596 (N_33596,N_30829,N_30910);
and U33597 (N_33597,N_30626,N_32035);
or U33598 (N_33598,N_31934,N_30244);
xnor U33599 (N_33599,N_32032,N_30756);
and U33600 (N_33600,N_31777,N_31876);
nor U33601 (N_33601,N_32486,N_32302);
nor U33602 (N_33602,N_31709,N_32209);
xnor U33603 (N_33603,N_30448,N_30704);
or U33604 (N_33604,N_31947,N_32193);
nor U33605 (N_33605,N_31858,N_30615);
xnor U33606 (N_33606,N_32111,N_31929);
nor U33607 (N_33607,N_32215,N_30102);
nor U33608 (N_33608,N_32343,N_30450);
xor U33609 (N_33609,N_30481,N_30355);
xnor U33610 (N_33610,N_30850,N_30906);
or U33611 (N_33611,N_32475,N_30550);
nor U33612 (N_33612,N_31413,N_31476);
xor U33613 (N_33613,N_31925,N_30795);
and U33614 (N_33614,N_30814,N_32134);
xor U33615 (N_33615,N_32361,N_32257);
or U33616 (N_33616,N_31005,N_32423);
or U33617 (N_33617,N_30222,N_31549);
and U33618 (N_33618,N_31502,N_30471);
or U33619 (N_33619,N_32323,N_31994);
or U33620 (N_33620,N_30257,N_31712);
nand U33621 (N_33621,N_30387,N_30186);
and U33622 (N_33622,N_31036,N_32042);
and U33623 (N_33623,N_31798,N_31455);
or U33624 (N_33624,N_32026,N_30225);
nor U33625 (N_33625,N_31572,N_30092);
nand U33626 (N_33626,N_30648,N_30308);
nand U33627 (N_33627,N_31306,N_31772);
nand U33628 (N_33628,N_31767,N_30293);
nor U33629 (N_33629,N_31735,N_30796);
nand U33630 (N_33630,N_31559,N_32392);
xnor U33631 (N_33631,N_31313,N_30876);
and U33632 (N_33632,N_31285,N_31703);
nand U33633 (N_33633,N_31965,N_31747);
or U33634 (N_33634,N_32089,N_31627);
and U33635 (N_33635,N_31957,N_30635);
or U33636 (N_33636,N_30288,N_30623);
or U33637 (N_33637,N_30134,N_32284);
nor U33638 (N_33638,N_31533,N_31065);
nor U33639 (N_33639,N_31854,N_31071);
nor U33640 (N_33640,N_30237,N_31235);
nand U33641 (N_33641,N_30555,N_30154);
nand U33642 (N_33642,N_32115,N_30256);
nor U33643 (N_33643,N_31579,N_31832);
and U33644 (N_33644,N_30195,N_32375);
nand U33645 (N_33645,N_31707,N_30737);
nor U33646 (N_33646,N_31705,N_31653);
nor U33647 (N_33647,N_31515,N_31562);
or U33648 (N_33648,N_31666,N_30641);
or U33649 (N_33649,N_30018,N_31978);
nor U33650 (N_33650,N_31545,N_30671);
nand U33651 (N_33651,N_31128,N_30831);
xor U33652 (N_33652,N_30053,N_31642);
nand U33653 (N_33653,N_32371,N_31287);
and U33654 (N_33654,N_30103,N_30909);
xor U33655 (N_33655,N_30188,N_30056);
or U33656 (N_33656,N_31083,N_32141);
nand U33657 (N_33657,N_31304,N_30124);
or U33658 (N_33658,N_30834,N_30896);
xnor U33659 (N_33659,N_30541,N_30153);
and U33660 (N_33660,N_31599,N_31180);
and U33661 (N_33661,N_30296,N_31008);
nand U33662 (N_33662,N_32349,N_30362);
xor U33663 (N_33663,N_31215,N_30999);
nand U33664 (N_33664,N_30517,N_32187);
xor U33665 (N_33665,N_30571,N_30907);
or U33666 (N_33666,N_30412,N_30744);
xor U33667 (N_33667,N_31991,N_31242);
nor U33668 (N_33668,N_30902,N_32478);
or U33669 (N_33669,N_30235,N_31906);
xnor U33670 (N_33670,N_30128,N_31669);
nor U33671 (N_33671,N_30443,N_31567);
and U33672 (N_33672,N_31505,N_30811);
nor U33673 (N_33673,N_31457,N_30325);
nand U33674 (N_33674,N_31109,N_30181);
nand U33675 (N_33675,N_31937,N_30752);
nor U33676 (N_33676,N_32221,N_31216);
nand U33677 (N_33677,N_31274,N_32448);
nor U33678 (N_33678,N_31692,N_32404);
xor U33679 (N_33679,N_32433,N_31847);
nand U33680 (N_33680,N_32243,N_31470);
xnor U33681 (N_33681,N_31351,N_30350);
nor U33682 (N_33682,N_31465,N_32426);
and U33683 (N_33683,N_30516,N_30112);
nor U33684 (N_33684,N_31637,N_32399);
nand U33685 (N_33685,N_30529,N_30783);
or U33686 (N_33686,N_30398,N_30765);
or U33687 (N_33687,N_30984,N_31333);
or U33688 (N_33688,N_31909,N_31219);
xor U33689 (N_33689,N_30854,N_30426);
nand U33690 (N_33690,N_30943,N_31221);
and U33691 (N_33691,N_31611,N_30961);
nand U33692 (N_33692,N_31499,N_32271);
nor U33693 (N_33693,N_32266,N_30871);
nand U33694 (N_33694,N_30351,N_31384);
xnor U33695 (N_33695,N_30280,N_32125);
xnor U33696 (N_33696,N_30405,N_31926);
or U33697 (N_33697,N_30007,N_31526);
xor U33698 (N_33698,N_31323,N_32082);
and U33699 (N_33699,N_31780,N_32182);
nor U33700 (N_33700,N_31895,N_30360);
or U33701 (N_33701,N_30766,N_30258);
xnor U33702 (N_33702,N_31450,N_32023);
or U33703 (N_33703,N_31102,N_32480);
or U33704 (N_33704,N_32440,N_30488);
and U33705 (N_33705,N_30980,N_31001);
xor U33706 (N_33706,N_31366,N_30307);
and U33707 (N_33707,N_32429,N_32467);
and U33708 (N_33708,N_32304,N_30702);
nor U33709 (N_33709,N_30782,N_30376);
nor U33710 (N_33710,N_30099,N_32412);
and U33711 (N_33711,N_31554,N_30404);
nand U33712 (N_33712,N_31746,N_31737);
xnor U33713 (N_33713,N_31982,N_30480);
nor U33714 (N_33714,N_30863,N_30564);
nand U33715 (N_33715,N_31523,N_30229);
or U33716 (N_33716,N_30152,N_31664);
or U33717 (N_33717,N_30558,N_31194);
nor U33718 (N_33718,N_31510,N_30300);
nor U33719 (N_33719,N_30747,N_31741);
xnor U33720 (N_33720,N_30813,N_31038);
and U33721 (N_33721,N_30138,N_30920);
xnor U33722 (N_33722,N_30703,N_30840);
and U33723 (N_33723,N_32308,N_31420);
and U33724 (N_33724,N_30954,N_32416);
nor U33725 (N_33725,N_30970,N_30205);
nor U33726 (N_33726,N_30554,N_30281);
and U33727 (N_33727,N_30621,N_31849);
or U33728 (N_33728,N_31361,N_32175);
nor U33729 (N_33729,N_31225,N_30370);
or U33730 (N_33730,N_31790,N_30435);
or U33731 (N_33731,N_30650,N_31802);
nand U33732 (N_33732,N_30429,N_31821);
or U33733 (N_33733,N_31682,N_30466);
and U33734 (N_33734,N_31341,N_32159);
nand U33735 (N_33735,N_31975,N_30170);
nor U33736 (N_33736,N_30219,N_30228);
or U33737 (N_33737,N_30892,N_31736);
xor U33738 (N_33738,N_30802,N_30344);
nor U33739 (N_33739,N_32457,N_30046);
nor U33740 (N_33740,N_31440,N_30231);
or U33741 (N_33741,N_31625,N_30694);
and U33742 (N_33742,N_30282,N_31739);
and U33743 (N_33743,N_31868,N_31785);
nor U33744 (N_33744,N_30602,N_32226);
or U33745 (N_33745,N_31427,N_32059);
nor U33746 (N_33746,N_30528,N_32129);
nand U33747 (N_33747,N_30580,N_31414);
nand U33748 (N_33748,N_31540,N_31443);
or U33749 (N_33749,N_30234,N_31766);
nor U33750 (N_33750,N_31725,N_31968);
nor U33751 (N_33751,N_31692,N_30164);
and U33752 (N_33752,N_30909,N_31003);
and U33753 (N_33753,N_30502,N_32387);
and U33754 (N_33754,N_31637,N_31624);
xnor U33755 (N_33755,N_31200,N_31203);
nand U33756 (N_33756,N_31773,N_30983);
xor U33757 (N_33757,N_30880,N_30144);
nor U33758 (N_33758,N_30887,N_32333);
or U33759 (N_33759,N_30251,N_31736);
xor U33760 (N_33760,N_30660,N_31550);
and U33761 (N_33761,N_30443,N_30548);
and U33762 (N_33762,N_32417,N_31852);
xnor U33763 (N_33763,N_31897,N_31424);
or U33764 (N_33764,N_30812,N_31290);
nor U33765 (N_33765,N_31788,N_30285);
nor U33766 (N_33766,N_32110,N_31641);
and U33767 (N_33767,N_30132,N_30000);
xor U33768 (N_33768,N_31153,N_31453);
xnor U33769 (N_33769,N_31111,N_30402);
xor U33770 (N_33770,N_30907,N_32310);
nand U33771 (N_33771,N_31477,N_31484);
nand U33772 (N_33772,N_32360,N_32019);
nand U33773 (N_33773,N_30895,N_31897);
nand U33774 (N_33774,N_30152,N_31869);
xor U33775 (N_33775,N_31073,N_31462);
nand U33776 (N_33776,N_30838,N_31451);
nand U33777 (N_33777,N_31895,N_31068);
nand U33778 (N_33778,N_30089,N_31047);
nand U33779 (N_33779,N_30346,N_31864);
nor U33780 (N_33780,N_31778,N_32119);
xor U33781 (N_33781,N_30657,N_31582);
or U33782 (N_33782,N_31462,N_30260);
xor U33783 (N_33783,N_30978,N_31616);
nand U33784 (N_33784,N_30035,N_30927);
nand U33785 (N_33785,N_30827,N_30239);
nand U33786 (N_33786,N_32338,N_30184);
or U33787 (N_33787,N_30945,N_32272);
or U33788 (N_33788,N_31078,N_30727);
xnor U33789 (N_33789,N_30362,N_30807);
nand U33790 (N_33790,N_30204,N_31349);
or U33791 (N_33791,N_32166,N_30588);
and U33792 (N_33792,N_31632,N_30746);
and U33793 (N_33793,N_31155,N_30560);
nor U33794 (N_33794,N_32302,N_32399);
or U33795 (N_33795,N_31667,N_32473);
and U33796 (N_33796,N_31022,N_30128);
nor U33797 (N_33797,N_30048,N_31232);
nand U33798 (N_33798,N_32451,N_30764);
xnor U33799 (N_33799,N_31648,N_30593);
nor U33800 (N_33800,N_30624,N_31445);
and U33801 (N_33801,N_30571,N_32267);
xnor U33802 (N_33802,N_31608,N_31537);
xor U33803 (N_33803,N_30718,N_31193);
nor U33804 (N_33804,N_31988,N_32317);
xor U33805 (N_33805,N_30092,N_30895);
or U33806 (N_33806,N_32011,N_30743);
and U33807 (N_33807,N_31448,N_31968);
and U33808 (N_33808,N_30598,N_31261);
xnor U33809 (N_33809,N_31144,N_32489);
xor U33810 (N_33810,N_31565,N_30607);
nand U33811 (N_33811,N_31709,N_30484);
xnor U33812 (N_33812,N_32314,N_30004);
nor U33813 (N_33813,N_30558,N_30281);
nand U33814 (N_33814,N_30761,N_31158);
xnor U33815 (N_33815,N_31059,N_30938);
nor U33816 (N_33816,N_30119,N_31228);
nand U33817 (N_33817,N_30872,N_30327);
and U33818 (N_33818,N_32088,N_31197);
nor U33819 (N_33819,N_31563,N_32068);
nor U33820 (N_33820,N_30053,N_32428);
and U33821 (N_33821,N_30283,N_31610);
and U33822 (N_33822,N_31805,N_31085);
nand U33823 (N_33823,N_30149,N_30524);
nand U33824 (N_33824,N_30009,N_31001);
and U33825 (N_33825,N_31668,N_32051);
nor U33826 (N_33826,N_32148,N_31908);
or U33827 (N_33827,N_30590,N_31793);
xnor U33828 (N_33828,N_30133,N_30225);
nand U33829 (N_33829,N_31140,N_30249);
or U33830 (N_33830,N_31815,N_31177);
nand U33831 (N_33831,N_31989,N_30024);
nor U33832 (N_33832,N_31966,N_31551);
nand U33833 (N_33833,N_31421,N_30121);
and U33834 (N_33834,N_30049,N_32430);
and U33835 (N_33835,N_30226,N_32353);
nor U33836 (N_33836,N_31419,N_30131);
xor U33837 (N_33837,N_30453,N_30469);
xor U33838 (N_33838,N_30891,N_31000);
nand U33839 (N_33839,N_30328,N_31643);
xnor U33840 (N_33840,N_32134,N_32012);
nand U33841 (N_33841,N_31278,N_31234);
xor U33842 (N_33842,N_30537,N_30846);
and U33843 (N_33843,N_32336,N_32424);
or U33844 (N_33844,N_31391,N_30790);
nand U33845 (N_33845,N_31666,N_31293);
nand U33846 (N_33846,N_31367,N_30367);
xnor U33847 (N_33847,N_30658,N_30955);
xor U33848 (N_33848,N_30570,N_31934);
and U33849 (N_33849,N_31924,N_31165);
nand U33850 (N_33850,N_30373,N_32406);
nor U33851 (N_33851,N_31744,N_31556);
nand U33852 (N_33852,N_30828,N_30762);
xor U33853 (N_33853,N_32009,N_31980);
or U33854 (N_33854,N_31541,N_30181);
or U33855 (N_33855,N_31015,N_31802);
or U33856 (N_33856,N_32321,N_30336);
xor U33857 (N_33857,N_32138,N_30205);
nand U33858 (N_33858,N_31500,N_32170);
or U33859 (N_33859,N_30143,N_30580);
and U33860 (N_33860,N_30797,N_30683);
xnor U33861 (N_33861,N_30490,N_30583);
nor U33862 (N_33862,N_30700,N_30316);
and U33863 (N_33863,N_31007,N_31730);
nor U33864 (N_33864,N_30798,N_30448);
or U33865 (N_33865,N_30115,N_30135);
or U33866 (N_33866,N_32213,N_31120);
xor U33867 (N_33867,N_32102,N_31915);
or U33868 (N_33868,N_30999,N_31934);
and U33869 (N_33869,N_30187,N_31056);
and U33870 (N_33870,N_30444,N_30524);
or U33871 (N_33871,N_31540,N_32305);
xor U33872 (N_33872,N_32122,N_30916);
nand U33873 (N_33873,N_31443,N_30017);
and U33874 (N_33874,N_30106,N_30317);
nor U33875 (N_33875,N_32280,N_31376);
or U33876 (N_33876,N_31908,N_31329);
and U33877 (N_33877,N_31923,N_31155);
or U33878 (N_33878,N_31774,N_31268);
xnor U33879 (N_33879,N_30998,N_30428);
xnor U33880 (N_33880,N_31708,N_32467);
nand U33881 (N_33881,N_30891,N_30126);
xor U33882 (N_33882,N_30237,N_32238);
and U33883 (N_33883,N_30596,N_32287);
or U33884 (N_33884,N_31878,N_30602);
nor U33885 (N_33885,N_31292,N_32058);
xor U33886 (N_33886,N_32300,N_32126);
xnor U33887 (N_33887,N_30710,N_32248);
nor U33888 (N_33888,N_30940,N_30624);
nand U33889 (N_33889,N_32262,N_30417);
xor U33890 (N_33890,N_30021,N_30948);
or U33891 (N_33891,N_31281,N_32399);
nand U33892 (N_33892,N_31137,N_31658);
nand U33893 (N_33893,N_31324,N_30448);
and U33894 (N_33894,N_31058,N_32463);
or U33895 (N_33895,N_32016,N_31659);
xor U33896 (N_33896,N_30846,N_32462);
or U33897 (N_33897,N_32042,N_31012);
and U33898 (N_33898,N_30651,N_31646);
nor U33899 (N_33899,N_31003,N_31784);
and U33900 (N_33900,N_30536,N_31192);
nand U33901 (N_33901,N_31026,N_30372);
or U33902 (N_33902,N_32264,N_31146);
or U33903 (N_33903,N_31529,N_30403);
and U33904 (N_33904,N_30797,N_32312);
xor U33905 (N_33905,N_32080,N_30745);
or U33906 (N_33906,N_30312,N_31880);
or U33907 (N_33907,N_31105,N_30071);
nand U33908 (N_33908,N_31970,N_31896);
or U33909 (N_33909,N_30765,N_32254);
nand U33910 (N_33910,N_31067,N_31092);
or U33911 (N_33911,N_30365,N_30071);
nand U33912 (N_33912,N_32157,N_31457);
or U33913 (N_33913,N_31341,N_32231);
nand U33914 (N_33914,N_32023,N_30254);
and U33915 (N_33915,N_32041,N_31556);
xnor U33916 (N_33916,N_31108,N_30398);
or U33917 (N_33917,N_31892,N_32166);
and U33918 (N_33918,N_31692,N_31204);
and U33919 (N_33919,N_32030,N_30660);
or U33920 (N_33920,N_31232,N_31052);
or U33921 (N_33921,N_31934,N_30544);
xor U33922 (N_33922,N_32429,N_31966);
xor U33923 (N_33923,N_30867,N_32303);
nor U33924 (N_33924,N_32493,N_31763);
xnor U33925 (N_33925,N_32160,N_32331);
xnor U33926 (N_33926,N_31743,N_30496);
nand U33927 (N_33927,N_32480,N_30160);
xnor U33928 (N_33928,N_30932,N_30202);
and U33929 (N_33929,N_32499,N_31170);
nor U33930 (N_33930,N_30354,N_30056);
nand U33931 (N_33931,N_30098,N_30866);
xor U33932 (N_33932,N_30001,N_31422);
nor U33933 (N_33933,N_30140,N_31222);
xnor U33934 (N_33934,N_30134,N_31147);
or U33935 (N_33935,N_30379,N_31144);
nand U33936 (N_33936,N_32420,N_30557);
xor U33937 (N_33937,N_30626,N_30379);
and U33938 (N_33938,N_32331,N_30358);
xnor U33939 (N_33939,N_30571,N_31371);
and U33940 (N_33940,N_30186,N_30069);
nand U33941 (N_33941,N_31747,N_31767);
or U33942 (N_33942,N_30653,N_32355);
xor U33943 (N_33943,N_31265,N_31090);
xnor U33944 (N_33944,N_31317,N_30892);
and U33945 (N_33945,N_30786,N_30727);
nor U33946 (N_33946,N_31824,N_31393);
and U33947 (N_33947,N_30814,N_31058);
or U33948 (N_33948,N_31766,N_31600);
nor U33949 (N_33949,N_32049,N_31902);
or U33950 (N_33950,N_32051,N_30666);
nor U33951 (N_33951,N_32452,N_30147);
xor U33952 (N_33952,N_30277,N_30025);
nor U33953 (N_33953,N_30884,N_30017);
xor U33954 (N_33954,N_30603,N_32033);
nor U33955 (N_33955,N_30661,N_31712);
or U33956 (N_33956,N_30499,N_30305);
nand U33957 (N_33957,N_32012,N_32285);
or U33958 (N_33958,N_31455,N_30834);
nor U33959 (N_33959,N_30893,N_30625);
or U33960 (N_33960,N_30112,N_31232);
xor U33961 (N_33961,N_30596,N_32227);
nand U33962 (N_33962,N_30091,N_31567);
nor U33963 (N_33963,N_31567,N_30829);
nor U33964 (N_33964,N_30285,N_30500);
nand U33965 (N_33965,N_30143,N_31393);
or U33966 (N_33966,N_31603,N_31544);
and U33967 (N_33967,N_30440,N_31590);
and U33968 (N_33968,N_31622,N_30666);
and U33969 (N_33969,N_32397,N_31087);
and U33970 (N_33970,N_32308,N_31273);
nor U33971 (N_33971,N_30706,N_32106);
and U33972 (N_33972,N_32104,N_30794);
nand U33973 (N_33973,N_31732,N_31772);
nor U33974 (N_33974,N_30359,N_30926);
nand U33975 (N_33975,N_30236,N_30703);
or U33976 (N_33976,N_31797,N_31866);
xor U33977 (N_33977,N_30571,N_31063);
and U33978 (N_33978,N_31696,N_31698);
nor U33979 (N_33979,N_31265,N_30468);
and U33980 (N_33980,N_30893,N_30235);
xnor U33981 (N_33981,N_32456,N_32155);
nand U33982 (N_33982,N_32157,N_30776);
or U33983 (N_33983,N_30173,N_30077);
nor U33984 (N_33984,N_30804,N_30407);
xnor U33985 (N_33985,N_31588,N_31499);
xnor U33986 (N_33986,N_32455,N_31910);
or U33987 (N_33987,N_30477,N_30271);
nor U33988 (N_33988,N_31254,N_30642);
nor U33989 (N_33989,N_30318,N_31657);
and U33990 (N_33990,N_32257,N_31647);
nor U33991 (N_33991,N_30180,N_31871);
or U33992 (N_33992,N_30521,N_32388);
or U33993 (N_33993,N_30257,N_31157);
and U33994 (N_33994,N_31515,N_31149);
or U33995 (N_33995,N_30765,N_32309);
or U33996 (N_33996,N_30509,N_30413);
xnor U33997 (N_33997,N_31109,N_31902);
xor U33998 (N_33998,N_30452,N_30587);
or U33999 (N_33999,N_31333,N_31771);
xor U34000 (N_34000,N_32301,N_32431);
nand U34001 (N_34001,N_30125,N_30036);
nand U34002 (N_34002,N_31467,N_30256);
xor U34003 (N_34003,N_30336,N_31324);
and U34004 (N_34004,N_31584,N_31337);
and U34005 (N_34005,N_31479,N_30410);
nand U34006 (N_34006,N_30102,N_31521);
or U34007 (N_34007,N_31049,N_30837);
xor U34008 (N_34008,N_30824,N_31555);
or U34009 (N_34009,N_31805,N_30011);
xnor U34010 (N_34010,N_30453,N_30050);
nand U34011 (N_34011,N_30590,N_31568);
or U34012 (N_34012,N_30239,N_31731);
and U34013 (N_34013,N_30065,N_32064);
and U34014 (N_34014,N_30156,N_30431);
and U34015 (N_34015,N_31401,N_30409);
or U34016 (N_34016,N_30336,N_31273);
nand U34017 (N_34017,N_30819,N_31555);
nand U34018 (N_34018,N_30540,N_32436);
or U34019 (N_34019,N_30518,N_31375);
xor U34020 (N_34020,N_30632,N_30389);
nor U34021 (N_34021,N_30256,N_31858);
nand U34022 (N_34022,N_30092,N_31181);
nand U34023 (N_34023,N_31342,N_31656);
and U34024 (N_34024,N_30169,N_31341);
nand U34025 (N_34025,N_31485,N_32120);
xor U34026 (N_34026,N_31634,N_31562);
and U34027 (N_34027,N_30155,N_30223);
and U34028 (N_34028,N_32013,N_30239);
or U34029 (N_34029,N_32416,N_30907);
xnor U34030 (N_34030,N_30711,N_31412);
nor U34031 (N_34031,N_32213,N_30769);
nand U34032 (N_34032,N_32447,N_32412);
nand U34033 (N_34033,N_30298,N_30439);
xnor U34034 (N_34034,N_31448,N_31577);
nor U34035 (N_34035,N_31909,N_30304);
or U34036 (N_34036,N_31840,N_30036);
nor U34037 (N_34037,N_30209,N_30737);
or U34038 (N_34038,N_31549,N_31644);
xor U34039 (N_34039,N_30988,N_31899);
nand U34040 (N_34040,N_31831,N_30788);
and U34041 (N_34041,N_32348,N_31833);
nand U34042 (N_34042,N_31987,N_30946);
nand U34043 (N_34043,N_32379,N_30227);
xor U34044 (N_34044,N_31360,N_31721);
and U34045 (N_34045,N_32492,N_31856);
nand U34046 (N_34046,N_30648,N_30080);
xnor U34047 (N_34047,N_30560,N_31052);
nand U34048 (N_34048,N_32089,N_32155);
and U34049 (N_34049,N_30065,N_32125);
and U34050 (N_34050,N_30196,N_31275);
or U34051 (N_34051,N_32403,N_30158);
xor U34052 (N_34052,N_31682,N_30375);
nor U34053 (N_34053,N_31020,N_32007);
or U34054 (N_34054,N_30624,N_32321);
xor U34055 (N_34055,N_30007,N_31400);
xnor U34056 (N_34056,N_30976,N_30737);
or U34057 (N_34057,N_30074,N_31444);
nor U34058 (N_34058,N_31967,N_32495);
or U34059 (N_34059,N_32488,N_30611);
nand U34060 (N_34060,N_31309,N_31607);
and U34061 (N_34061,N_31867,N_30822);
xor U34062 (N_34062,N_30301,N_31279);
xor U34063 (N_34063,N_30229,N_32485);
and U34064 (N_34064,N_31923,N_30736);
and U34065 (N_34065,N_31660,N_30899);
xor U34066 (N_34066,N_30444,N_30379);
nor U34067 (N_34067,N_31146,N_32391);
and U34068 (N_34068,N_30395,N_32463);
and U34069 (N_34069,N_30745,N_30962);
and U34070 (N_34070,N_31573,N_30595);
and U34071 (N_34071,N_30654,N_30000);
or U34072 (N_34072,N_30539,N_31063);
nand U34073 (N_34073,N_30526,N_31619);
or U34074 (N_34074,N_32359,N_31275);
nand U34075 (N_34075,N_32073,N_31922);
nor U34076 (N_34076,N_32318,N_30568);
xnor U34077 (N_34077,N_30323,N_30432);
xnor U34078 (N_34078,N_32298,N_30522);
or U34079 (N_34079,N_30217,N_30977);
nor U34080 (N_34080,N_30906,N_31170);
and U34081 (N_34081,N_30703,N_30408);
xnor U34082 (N_34082,N_30892,N_31109);
nand U34083 (N_34083,N_32009,N_32154);
and U34084 (N_34084,N_30506,N_32221);
nor U34085 (N_34085,N_30827,N_30007);
xnor U34086 (N_34086,N_30891,N_30198);
or U34087 (N_34087,N_30922,N_31813);
and U34088 (N_34088,N_30775,N_30445);
or U34089 (N_34089,N_31963,N_32099);
xor U34090 (N_34090,N_31981,N_30711);
nand U34091 (N_34091,N_31513,N_30195);
and U34092 (N_34092,N_31904,N_30151);
and U34093 (N_34093,N_30016,N_31961);
and U34094 (N_34094,N_30538,N_32179);
or U34095 (N_34095,N_32336,N_31661);
and U34096 (N_34096,N_31093,N_31964);
nand U34097 (N_34097,N_30835,N_30940);
xor U34098 (N_34098,N_30489,N_31105);
nor U34099 (N_34099,N_30380,N_30291);
nor U34100 (N_34100,N_30482,N_32478);
nor U34101 (N_34101,N_31931,N_30058);
xor U34102 (N_34102,N_30498,N_30668);
nand U34103 (N_34103,N_30382,N_30344);
and U34104 (N_34104,N_31685,N_32143);
nand U34105 (N_34105,N_31966,N_31590);
and U34106 (N_34106,N_30299,N_31155);
nand U34107 (N_34107,N_32341,N_30730);
and U34108 (N_34108,N_30521,N_30369);
or U34109 (N_34109,N_31725,N_30179);
xnor U34110 (N_34110,N_30735,N_32145);
and U34111 (N_34111,N_30043,N_31575);
xnor U34112 (N_34112,N_30011,N_31498);
xor U34113 (N_34113,N_31572,N_32182);
and U34114 (N_34114,N_31875,N_30980);
xor U34115 (N_34115,N_31815,N_30355);
and U34116 (N_34116,N_30431,N_32228);
xnor U34117 (N_34117,N_30809,N_30599);
xor U34118 (N_34118,N_30916,N_31634);
nand U34119 (N_34119,N_31084,N_32361);
nor U34120 (N_34120,N_32231,N_31233);
and U34121 (N_34121,N_31734,N_30474);
and U34122 (N_34122,N_30016,N_31316);
nand U34123 (N_34123,N_30816,N_31176);
nor U34124 (N_34124,N_31326,N_31779);
nor U34125 (N_34125,N_30086,N_31561);
nand U34126 (N_34126,N_30151,N_30128);
or U34127 (N_34127,N_31506,N_31667);
and U34128 (N_34128,N_30609,N_31665);
xor U34129 (N_34129,N_31624,N_31765);
nand U34130 (N_34130,N_30780,N_31679);
and U34131 (N_34131,N_32462,N_30096);
or U34132 (N_34132,N_30674,N_30253);
or U34133 (N_34133,N_31866,N_30589);
or U34134 (N_34134,N_31009,N_32291);
nor U34135 (N_34135,N_30534,N_30691);
nor U34136 (N_34136,N_30819,N_31467);
xnor U34137 (N_34137,N_30220,N_30439);
or U34138 (N_34138,N_30021,N_30439);
xnor U34139 (N_34139,N_31464,N_30274);
nand U34140 (N_34140,N_31082,N_31046);
or U34141 (N_34141,N_30485,N_31589);
or U34142 (N_34142,N_30675,N_30854);
xnor U34143 (N_34143,N_30857,N_32464);
nand U34144 (N_34144,N_30796,N_31939);
xor U34145 (N_34145,N_32490,N_31403);
or U34146 (N_34146,N_32388,N_31067);
nand U34147 (N_34147,N_30415,N_30989);
nor U34148 (N_34148,N_32058,N_30472);
nor U34149 (N_34149,N_32243,N_32298);
and U34150 (N_34150,N_31755,N_31500);
and U34151 (N_34151,N_31323,N_32158);
xor U34152 (N_34152,N_30349,N_31540);
nor U34153 (N_34153,N_31940,N_32417);
xnor U34154 (N_34154,N_31306,N_31482);
nand U34155 (N_34155,N_31201,N_31571);
and U34156 (N_34156,N_32243,N_31186);
or U34157 (N_34157,N_32010,N_31418);
xnor U34158 (N_34158,N_32214,N_31023);
xnor U34159 (N_34159,N_30300,N_31162);
and U34160 (N_34160,N_30941,N_31421);
xnor U34161 (N_34161,N_31704,N_31176);
nor U34162 (N_34162,N_31538,N_30183);
and U34163 (N_34163,N_31262,N_30016);
or U34164 (N_34164,N_31453,N_32221);
xor U34165 (N_34165,N_31782,N_30359);
xnor U34166 (N_34166,N_32269,N_31735);
or U34167 (N_34167,N_32405,N_30385);
nand U34168 (N_34168,N_30765,N_30775);
or U34169 (N_34169,N_30258,N_31414);
nor U34170 (N_34170,N_31807,N_32418);
and U34171 (N_34171,N_31820,N_31591);
xor U34172 (N_34172,N_30518,N_31471);
xor U34173 (N_34173,N_30184,N_30562);
and U34174 (N_34174,N_32208,N_31832);
or U34175 (N_34175,N_32279,N_30360);
or U34176 (N_34176,N_31773,N_31154);
nand U34177 (N_34177,N_32154,N_32186);
and U34178 (N_34178,N_30044,N_32085);
xor U34179 (N_34179,N_30457,N_31796);
xor U34180 (N_34180,N_31048,N_30167);
or U34181 (N_34181,N_30392,N_32413);
and U34182 (N_34182,N_32269,N_32445);
and U34183 (N_34183,N_32414,N_31735);
or U34184 (N_34184,N_30165,N_30169);
and U34185 (N_34185,N_30886,N_30610);
or U34186 (N_34186,N_32484,N_30253);
and U34187 (N_34187,N_32328,N_31448);
nor U34188 (N_34188,N_32037,N_32306);
or U34189 (N_34189,N_32170,N_30675);
or U34190 (N_34190,N_32499,N_32302);
nor U34191 (N_34191,N_32437,N_31423);
and U34192 (N_34192,N_30861,N_30772);
xor U34193 (N_34193,N_31608,N_31194);
nor U34194 (N_34194,N_31921,N_32022);
xnor U34195 (N_34195,N_32342,N_31742);
nor U34196 (N_34196,N_30379,N_30073);
nor U34197 (N_34197,N_30574,N_30926);
nand U34198 (N_34198,N_31722,N_31445);
xnor U34199 (N_34199,N_31889,N_31230);
xnor U34200 (N_34200,N_30529,N_30750);
nand U34201 (N_34201,N_32009,N_30343);
and U34202 (N_34202,N_31116,N_30288);
nand U34203 (N_34203,N_30575,N_32463);
nor U34204 (N_34204,N_30177,N_31891);
and U34205 (N_34205,N_30650,N_30701);
xnor U34206 (N_34206,N_31885,N_31730);
nand U34207 (N_34207,N_30956,N_31873);
and U34208 (N_34208,N_30138,N_31730);
or U34209 (N_34209,N_30366,N_31234);
and U34210 (N_34210,N_31979,N_30967);
or U34211 (N_34211,N_32395,N_32252);
nand U34212 (N_34212,N_30933,N_30120);
nand U34213 (N_34213,N_31371,N_31126);
nor U34214 (N_34214,N_32421,N_30342);
or U34215 (N_34215,N_31721,N_30239);
xnor U34216 (N_34216,N_31313,N_31904);
nor U34217 (N_34217,N_30232,N_30798);
nand U34218 (N_34218,N_31265,N_30876);
nor U34219 (N_34219,N_32120,N_31305);
nor U34220 (N_34220,N_31007,N_31835);
xnor U34221 (N_34221,N_30668,N_31748);
or U34222 (N_34222,N_31126,N_31081);
nor U34223 (N_34223,N_30752,N_30980);
xor U34224 (N_34224,N_31039,N_32485);
nor U34225 (N_34225,N_30659,N_32403);
nand U34226 (N_34226,N_30532,N_31118);
and U34227 (N_34227,N_30609,N_30275);
or U34228 (N_34228,N_32486,N_31144);
xor U34229 (N_34229,N_30573,N_30332);
nand U34230 (N_34230,N_30667,N_30886);
xnor U34231 (N_34231,N_31850,N_31278);
and U34232 (N_34232,N_30632,N_31524);
nand U34233 (N_34233,N_31976,N_32469);
xor U34234 (N_34234,N_30086,N_30239);
and U34235 (N_34235,N_30520,N_30518);
xor U34236 (N_34236,N_30708,N_30907);
nor U34237 (N_34237,N_30395,N_32366);
nor U34238 (N_34238,N_30386,N_30124);
xnor U34239 (N_34239,N_31443,N_32426);
or U34240 (N_34240,N_31702,N_32219);
or U34241 (N_34241,N_30264,N_31738);
nand U34242 (N_34242,N_31359,N_30072);
and U34243 (N_34243,N_32159,N_30399);
and U34244 (N_34244,N_32068,N_31596);
or U34245 (N_34245,N_31253,N_31465);
and U34246 (N_34246,N_31762,N_32354);
and U34247 (N_34247,N_30945,N_31637);
xnor U34248 (N_34248,N_31988,N_31632);
or U34249 (N_34249,N_30274,N_31718);
nor U34250 (N_34250,N_32228,N_31352);
and U34251 (N_34251,N_32146,N_31485);
nand U34252 (N_34252,N_30265,N_31256);
and U34253 (N_34253,N_32138,N_31338);
nand U34254 (N_34254,N_32141,N_32410);
nor U34255 (N_34255,N_32289,N_31609);
nor U34256 (N_34256,N_32223,N_30976);
nor U34257 (N_34257,N_30730,N_30173);
and U34258 (N_34258,N_32191,N_31804);
xnor U34259 (N_34259,N_31081,N_31641);
or U34260 (N_34260,N_31081,N_32305);
nor U34261 (N_34261,N_31052,N_31686);
and U34262 (N_34262,N_31913,N_31829);
nor U34263 (N_34263,N_31815,N_31846);
nor U34264 (N_34264,N_30726,N_31113);
nor U34265 (N_34265,N_30336,N_32431);
and U34266 (N_34266,N_31469,N_30141);
and U34267 (N_34267,N_31595,N_31280);
nor U34268 (N_34268,N_31621,N_30625);
or U34269 (N_34269,N_30017,N_31504);
or U34270 (N_34270,N_30534,N_30421);
xor U34271 (N_34271,N_31037,N_30691);
and U34272 (N_34272,N_31613,N_31899);
and U34273 (N_34273,N_31295,N_30507);
xor U34274 (N_34274,N_30354,N_32087);
nor U34275 (N_34275,N_30365,N_32463);
and U34276 (N_34276,N_31500,N_30629);
or U34277 (N_34277,N_31410,N_31087);
and U34278 (N_34278,N_30572,N_31933);
nand U34279 (N_34279,N_30596,N_31238);
xnor U34280 (N_34280,N_31988,N_31890);
or U34281 (N_34281,N_32453,N_30727);
or U34282 (N_34282,N_30633,N_31209);
and U34283 (N_34283,N_31991,N_30757);
xnor U34284 (N_34284,N_31811,N_30284);
nor U34285 (N_34285,N_32188,N_30149);
or U34286 (N_34286,N_31546,N_31070);
nand U34287 (N_34287,N_31418,N_30905);
and U34288 (N_34288,N_30024,N_30737);
xor U34289 (N_34289,N_30971,N_30921);
and U34290 (N_34290,N_32397,N_30918);
and U34291 (N_34291,N_30971,N_30517);
or U34292 (N_34292,N_30935,N_31893);
nand U34293 (N_34293,N_30974,N_31606);
nand U34294 (N_34294,N_32024,N_30342);
nand U34295 (N_34295,N_30972,N_30205);
or U34296 (N_34296,N_31866,N_30896);
or U34297 (N_34297,N_31310,N_31820);
or U34298 (N_34298,N_31957,N_30221);
or U34299 (N_34299,N_30975,N_30346);
nand U34300 (N_34300,N_31431,N_32316);
and U34301 (N_34301,N_32412,N_32166);
nand U34302 (N_34302,N_31534,N_30025);
nand U34303 (N_34303,N_30311,N_30351);
or U34304 (N_34304,N_31584,N_32478);
and U34305 (N_34305,N_30623,N_31386);
nor U34306 (N_34306,N_31227,N_30905);
nor U34307 (N_34307,N_31216,N_30543);
nor U34308 (N_34308,N_30888,N_31044);
xor U34309 (N_34309,N_30435,N_31047);
nand U34310 (N_34310,N_32200,N_30876);
xor U34311 (N_34311,N_31267,N_31776);
or U34312 (N_34312,N_30268,N_30514);
and U34313 (N_34313,N_30524,N_30613);
nor U34314 (N_34314,N_32067,N_30596);
xnor U34315 (N_34315,N_30110,N_30632);
and U34316 (N_34316,N_30801,N_31039);
xor U34317 (N_34317,N_32493,N_30627);
nand U34318 (N_34318,N_32227,N_31120);
xor U34319 (N_34319,N_32150,N_32402);
nor U34320 (N_34320,N_30308,N_31224);
or U34321 (N_34321,N_31481,N_30379);
and U34322 (N_34322,N_30319,N_30775);
nand U34323 (N_34323,N_31971,N_31111);
nor U34324 (N_34324,N_31856,N_32259);
nor U34325 (N_34325,N_31069,N_30493);
and U34326 (N_34326,N_31047,N_31465);
and U34327 (N_34327,N_31710,N_30018);
nand U34328 (N_34328,N_32470,N_30664);
or U34329 (N_34329,N_31101,N_31950);
nand U34330 (N_34330,N_32118,N_32245);
and U34331 (N_34331,N_31080,N_30863);
xor U34332 (N_34332,N_31999,N_31890);
or U34333 (N_34333,N_32430,N_32247);
and U34334 (N_34334,N_31755,N_30100);
nor U34335 (N_34335,N_30597,N_31509);
nor U34336 (N_34336,N_30328,N_32168);
and U34337 (N_34337,N_31522,N_30593);
nand U34338 (N_34338,N_30649,N_30046);
and U34339 (N_34339,N_30552,N_31898);
xor U34340 (N_34340,N_32192,N_31487);
and U34341 (N_34341,N_30213,N_31654);
nor U34342 (N_34342,N_32059,N_31103);
or U34343 (N_34343,N_32421,N_31995);
or U34344 (N_34344,N_31313,N_31315);
and U34345 (N_34345,N_31577,N_31132);
and U34346 (N_34346,N_31708,N_31625);
nor U34347 (N_34347,N_31163,N_30698);
and U34348 (N_34348,N_32337,N_30510);
xnor U34349 (N_34349,N_32446,N_32277);
or U34350 (N_34350,N_30827,N_32097);
and U34351 (N_34351,N_31693,N_32335);
and U34352 (N_34352,N_32159,N_31755);
nand U34353 (N_34353,N_30725,N_31151);
and U34354 (N_34354,N_31632,N_31249);
and U34355 (N_34355,N_31378,N_30564);
and U34356 (N_34356,N_30467,N_30141);
nor U34357 (N_34357,N_30787,N_31972);
or U34358 (N_34358,N_30369,N_30288);
xnor U34359 (N_34359,N_31967,N_32483);
and U34360 (N_34360,N_30215,N_31233);
and U34361 (N_34361,N_30839,N_31089);
nand U34362 (N_34362,N_30790,N_31541);
or U34363 (N_34363,N_32017,N_30693);
and U34364 (N_34364,N_30691,N_31058);
and U34365 (N_34365,N_30792,N_30231);
nor U34366 (N_34366,N_31807,N_31646);
and U34367 (N_34367,N_30664,N_31426);
nand U34368 (N_34368,N_31706,N_30124);
xor U34369 (N_34369,N_30895,N_30146);
nor U34370 (N_34370,N_31147,N_32194);
nor U34371 (N_34371,N_32167,N_32460);
xnor U34372 (N_34372,N_30063,N_30155);
xor U34373 (N_34373,N_31491,N_30323);
or U34374 (N_34374,N_31282,N_30343);
nor U34375 (N_34375,N_32139,N_31417);
nor U34376 (N_34376,N_31231,N_31347);
nand U34377 (N_34377,N_30557,N_31505);
xor U34378 (N_34378,N_32354,N_30650);
xnor U34379 (N_34379,N_31940,N_32057);
nor U34380 (N_34380,N_32346,N_31002);
xor U34381 (N_34381,N_30334,N_32034);
and U34382 (N_34382,N_30835,N_32114);
nor U34383 (N_34383,N_32386,N_32108);
nor U34384 (N_34384,N_30058,N_31371);
xor U34385 (N_34385,N_30060,N_32191);
xor U34386 (N_34386,N_30097,N_30886);
nor U34387 (N_34387,N_31858,N_31746);
and U34388 (N_34388,N_31561,N_30388);
and U34389 (N_34389,N_32224,N_31514);
nor U34390 (N_34390,N_30945,N_31158);
and U34391 (N_34391,N_30863,N_31360);
nand U34392 (N_34392,N_30756,N_31374);
nor U34393 (N_34393,N_30960,N_32318);
nand U34394 (N_34394,N_30408,N_30793);
nor U34395 (N_34395,N_32142,N_31660);
nand U34396 (N_34396,N_32064,N_31431);
or U34397 (N_34397,N_32478,N_30673);
nor U34398 (N_34398,N_30138,N_31263);
nand U34399 (N_34399,N_30646,N_32114);
nand U34400 (N_34400,N_31809,N_31492);
or U34401 (N_34401,N_31505,N_31479);
nand U34402 (N_34402,N_30176,N_31580);
nand U34403 (N_34403,N_32164,N_30600);
or U34404 (N_34404,N_30069,N_31707);
nor U34405 (N_34405,N_30455,N_30299);
and U34406 (N_34406,N_30737,N_30876);
or U34407 (N_34407,N_31410,N_30278);
nand U34408 (N_34408,N_31177,N_31811);
and U34409 (N_34409,N_32099,N_31174);
nor U34410 (N_34410,N_32170,N_30340);
or U34411 (N_34411,N_30567,N_30360);
nor U34412 (N_34412,N_30310,N_32306);
or U34413 (N_34413,N_31959,N_31932);
or U34414 (N_34414,N_30866,N_30911);
nor U34415 (N_34415,N_30808,N_31787);
xnor U34416 (N_34416,N_32073,N_31964);
xnor U34417 (N_34417,N_30272,N_31532);
nand U34418 (N_34418,N_30565,N_31492);
xor U34419 (N_34419,N_31648,N_30125);
or U34420 (N_34420,N_30730,N_30643);
nand U34421 (N_34421,N_31486,N_31449);
or U34422 (N_34422,N_30981,N_30404);
nor U34423 (N_34423,N_30755,N_31398);
and U34424 (N_34424,N_32385,N_31301);
nor U34425 (N_34425,N_32336,N_32213);
and U34426 (N_34426,N_32159,N_31065);
or U34427 (N_34427,N_32383,N_30253);
nor U34428 (N_34428,N_30651,N_31347);
nand U34429 (N_34429,N_31651,N_31159);
nor U34430 (N_34430,N_31350,N_31599);
or U34431 (N_34431,N_32382,N_30552);
nor U34432 (N_34432,N_32187,N_31215);
and U34433 (N_34433,N_31154,N_30328);
xor U34434 (N_34434,N_30238,N_31321);
nor U34435 (N_34435,N_31720,N_32424);
and U34436 (N_34436,N_30169,N_31405);
or U34437 (N_34437,N_31794,N_31626);
xor U34438 (N_34438,N_31334,N_31600);
xnor U34439 (N_34439,N_32354,N_31594);
or U34440 (N_34440,N_32294,N_30877);
or U34441 (N_34441,N_30577,N_31820);
and U34442 (N_34442,N_31200,N_31258);
or U34443 (N_34443,N_31573,N_32116);
nand U34444 (N_34444,N_32228,N_30448);
or U34445 (N_34445,N_32369,N_31444);
xnor U34446 (N_34446,N_31155,N_31651);
nand U34447 (N_34447,N_30274,N_31009);
nand U34448 (N_34448,N_30148,N_30245);
nand U34449 (N_34449,N_31118,N_30628);
nor U34450 (N_34450,N_32474,N_30867);
xor U34451 (N_34451,N_30737,N_30303);
and U34452 (N_34452,N_30726,N_30954);
nand U34453 (N_34453,N_30197,N_30926);
xnor U34454 (N_34454,N_31549,N_31998);
xnor U34455 (N_34455,N_30916,N_31716);
nor U34456 (N_34456,N_30135,N_31250);
and U34457 (N_34457,N_31404,N_32269);
xor U34458 (N_34458,N_31186,N_31596);
xnor U34459 (N_34459,N_32376,N_31067);
nand U34460 (N_34460,N_31468,N_30273);
and U34461 (N_34461,N_30898,N_31969);
and U34462 (N_34462,N_31033,N_31297);
nand U34463 (N_34463,N_30604,N_32254);
nand U34464 (N_34464,N_32094,N_31026);
xnor U34465 (N_34465,N_30984,N_32296);
nor U34466 (N_34466,N_32365,N_31222);
xnor U34467 (N_34467,N_31014,N_30359);
nand U34468 (N_34468,N_32412,N_32315);
and U34469 (N_34469,N_30003,N_32373);
xnor U34470 (N_34470,N_32417,N_31460);
nor U34471 (N_34471,N_30860,N_30770);
xnor U34472 (N_34472,N_30009,N_30991);
xnor U34473 (N_34473,N_30618,N_30640);
xor U34474 (N_34474,N_32271,N_30658);
or U34475 (N_34475,N_32160,N_31898);
xnor U34476 (N_34476,N_32389,N_31189);
xor U34477 (N_34477,N_30786,N_31175);
xnor U34478 (N_34478,N_31055,N_30437);
xor U34479 (N_34479,N_31689,N_30229);
and U34480 (N_34480,N_32290,N_30602);
and U34481 (N_34481,N_30333,N_30286);
and U34482 (N_34482,N_30654,N_30167);
and U34483 (N_34483,N_30854,N_30701);
nor U34484 (N_34484,N_30518,N_30635);
xor U34485 (N_34485,N_31972,N_32155);
nand U34486 (N_34486,N_32345,N_31595);
nor U34487 (N_34487,N_32190,N_30186);
nor U34488 (N_34488,N_30424,N_32210);
xor U34489 (N_34489,N_31224,N_30547);
or U34490 (N_34490,N_32115,N_32319);
xor U34491 (N_34491,N_31614,N_31664);
and U34492 (N_34492,N_30580,N_30185);
and U34493 (N_34493,N_30528,N_30819);
nand U34494 (N_34494,N_31945,N_31408);
xnor U34495 (N_34495,N_31048,N_30976);
nor U34496 (N_34496,N_32368,N_32399);
and U34497 (N_34497,N_30100,N_31068);
or U34498 (N_34498,N_30067,N_31233);
nand U34499 (N_34499,N_32428,N_31201);
nand U34500 (N_34500,N_31242,N_30800);
nand U34501 (N_34501,N_30539,N_30242);
or U34502 (N_34502,N_31647,N_30803);
or U34503 (N_34503,N_30771,N_30547);
or U34504 (N_34504,N_31102,N_30432);
nand U34505 (N_34505,N_31594,N_31043);
and U34506 (N_34506,N_30400,N_31732);
or U34507 (N_34507,N_30321,N_31434);
and U34508 (N_34508,N_32179,N_31227);
or U34509 (N_34509,N_32403,N_31600);
or U34510 (N_34510,N_32066,N_30206);
xnor U34511 (N_34511,N_31496,N_30139);
and U34512 (N_34512,N_30534,N_32403);
nor U34513 (N_34513,N_31608,N_30345);
or U34514 (N_34514,N_32473,N_31887);
and U34515 (N_34515,N_30741,N_31852);
nor U34516 (N_34516,N_30370,N_30202);
and U34517 (N_34517,N_31243,N_30005);
xnor U34518 (N_34518,N_32016,N_32372);
and U34519 (N_34519,N_31802,N_30144);
nor U34520 (N_34520,N_30885,N_32037);
nand U34521 (N_34521,N_30570,N_32127);
and U34522 (N_34522,N_31961,N_31874);
nand U34523 (N_34523,N_30158,N_30594);
nand U34524 (N_34524,N_30090,N_32049);
nor U34525 (N_34525,N_31949,N_32410);
and U34526 (N_34526,N_31607,N_32072);
xor U34527 (N_34527,N_30130,N_30796);
and U34528 (N_34528,N_31788,N_31747);
nor U34529 (N_34529,N_31909,N_31385);
nor U34530 (N_34530,N_30486,N_31216);
or U34531 (N_34531,N_31499,N_30259);
xnor U34532 (N_34532,N_32496,N_31476);
xnor U34533 (N_34533,N_32030,N_31690);
or U34534 (N_34534,N_31129,N_31505);
nand U34535 (N_34535,N_31705,N_31764);
nor U34536 (N_34536,N_31971,N_30379);
or U34537 (N_34537,N_32067,N_30265);
or U34538 (N_34538,N_31108,N_31298);
and U34539 (N_34539,N_30906,N_32242);
or U34540 (N_34540,N_32411,N_30269);
and U34541 (N_34541,N_30421,N_30398);
or U34542 (N_34542,N_30641,N_31359);
and U34543 (N_34543,N_30103,N_32188);
nand U34544 (N_34544,N_31936,N_32465);
nand U34545 (N_34545,N_30871,N_30104);
and U34546 (N_34546,N_32336,N_31154);
nand U34547 (N_34547,N_31731,N_31239);
nor U34548 (N_34548,N_30860,N_30951);
nand U34549 (N_34549,N_30678,N_31203);
and U34550 (N_34550,N_32326,N_31284);
and U34551 (N_34551,N_31713,N_30526);
nand U34552 (N_34552,N_30541,N_30331);
or U34553 (N_34553,N_31207,N_31021);
nand U34554 (N_34554,N_31837,N_31935);
or U34555 (N_34555,N_31021,N_32212);
or U34556 (N_34556,N_32272,N_31150);
and U34557 (N_34557,N_31380,N_30280);
and U34558 (N_34558,N_30457,N_30610);
nor U34559 (N_34559,N_30338,N_32167);
or U34560 (N_34560,N_30231,N_32077);
nor U34561 (N_34561,N_31595,N_31177);
nand U34562 (N_34562,N_31468,N_30780);
xor U34563 (N_34563,N_30257,N_30909);
and U34564 (N_34564,N_30932,N_30229);
xnor U34565 (N_34565,N_31291,N_30308);
xor U34566 (N_34566,N_32349,N_31853);
or U34567 (N_34567,N_32029,N_30373);
nand U34568 (N_34568,N_30384,N_30858);
xnor U34569 (N_34569,N_30785,N_30943);
or U34570 (N_34570,N_30300,N_32175);
nand U34571 (N_34571,N_32317,N_31179);
xor U34572 (N_34572,N_30807,N_31784);
xnor U34573 (N_34573,N_31537,N_30057);
xnor U34574 (N_34574,N_31130,N_30366);
nand U34575 (N_34575,N_31596,N_32385);
or U34576 (N_34576,N_31795,N_31310);
and U34577 (N_34577,N_30244,N_30918);
xnor U34578 (N_34578,N_31205,N_30922);
or U34579 (N_34579,N_30540,N_31588);
nand U34580 (N_34580,N_31153,N_32497);
and U34581 (N_34581,N_31014,N_31096);
nor U34582 (N_34582,N_31291,N_30405);
or U34583 (N_34583,N_30511,N_32379);
and U34584 (N_34584,N_31703,N_30466);
nor U34585 (N_34585,N_30859,N_31730);
xor U34586 (N_34586,N_30951,N_31364);
or U34587 (N_34587,N_32067,N_30058);
nand U34588 (N_34588,N_30818,N_31028);
xnor U34589 (N_34589,N_30679,N_31776);
nor U34590 (N_34590,N_31963,N_32220);
nor U34591 (N_34591,N_30722,N_31335);
xor U34592 (N_34592,N_30386,N_30228);
xor U34593 (N_34593,N_31946,N_31240);
xor U34594 (N_34594,N_30978,N_32248);
xor U34595 (N_34595,N_32279,N_31272);
nand U34596 (N_34596,N_30894,N_32326);
nor U34597 (N_34597,N_31408,N_31210);
xnor U34598 (N_34598,N_32494,N_31479);
nand U34599 (N_34599,N_32092,N_30222);
nand U34600 (N_34600,N_31350,N_31322);
xnor U34601 (N_34601,N_31240,N_32364);
and U34602 (N_34602,N_30510,N_32446);
or U34603 (N_34603,N_30492,N_30385);
nor U34604 (N_34604,N_30470,N_32170);
nand U34605 (N_34605,N_31415,N_32406);
xnor U34606 (N_34606,N_30110,N_31793);
nor U34607 (N_34607,N_31213,N_30867);
xnor U34608 (N_34608,N_31603,N_31820);
nand U34609 (N_34609,N_30244,N_32125);
or U34610 (N_34610,N_30242,N_30531);
nand U34611 (N_34611,N_32354,N_30014);
nand U34612 (N_34612,N_30996,N_32045);
xnor U34613 (N_34613,N_30646,N_30699);
and U34614 (N_34614,N_30537,N_31390);
nor U34615 (N_34615,N_31127,N_30061);
nor U34616 (N_34616,N_32376,N_30486);
and U34617 (N_34617,N_31384,N_30207);
nor U34618 (N_34618,N_30987,N_32341);
and U34619 (N_34619,N_31950,N_32120);
nor U34620 (N_34620,N_31677,N_31042);
xor U34621 (N_34621,N_30413,N_32334);
nand U34622 (N_34622,N_30593,N_32120);
or U34623 (N_34623,N_31668,N_30449);
or U34624 (N_34624,N_31506,N_32376);
xor U34625 (N_34625,N_30524,N_31031);
nor U34626 (N_34626,N_32326,N_30544);
nor U34627 (N_34627,N_30276,N_31817);
and U34628 (N_34628,N_32231,N_31157);
nor U34629 (N_34629,N_30424,N_31780);
or U34630 (N_34630,N_30850,N_30301);
and U34631 (N_34631,N_31517,N_30091);
and U34632 (N_34632,N_31523,N_30445);
and U34633 (N_34633,N_30467,N_31162);
nor U34634 (N_34634,N_31207,N_31700);
xor U34635 (N_34635,N_30881,N_30225);
nand U34636 (N_34636,N_31617,N_31996);
or U34637 (N_34637,N_30412,N_30002);
or U34638 (N_34638,N_30610,N_30165);
or U34639 (N_34639,N_30909,N_30727);
xnor U34640 (N_34640,N_30878,N_31350);
nand U34641 (N_34641,N_30803,N_31721);
xnor U34642 (N_34642,N_30661,N_31997);
nor U34643 (N_34643,N_32059,N_32444);
xor U34644 (N_34644,N_32155,N_32438);
or U34645 (N_34645,N_30395,N_30392);
or U34646 (N_34646,N_30541,N_30547);
and U34647 (N_34647,N_31258,N_31636);
nand U34648 (N_34648,N_30535,N_32087);
nor U34649 (N_34649,N_31290,N_31491);
nand U34650 (N_34650,N_30699,N_31594);
xor U34651 (N_34651,N_32168,N_32109);
or U34652 (N_34652,N_31500,N_30990);
nor U34653 (N_34653,N_30581,N_31458);
nand U34654 (N_34654,N_31670,N_32406);
nor U34655 (N_34655,N_30720,N_32233);
nor U34656 (N_34656,N_31380,N_31890);
and U34657 (N_34657,N_32492,N_30418);
or U34658 (N_34658,N_30496,N_30387);
or U34659 (N_34659,N_30692,N_30812);
or U34660 (N_34660,N_30508,N_31102);
nand U34661 (N_34661,N_30381,N_31379);
or U34662 (N_34662,N_31343,N_30594);
and U34663 (N_34663,N_30740,N_30928);
xor U34664 (N_34664,N_30038,N_30093);
xnor U34665 (N_34665,N_30888,N_32116);
nand U34666 (N_34666,N_31329,N_30285);
nand U34667 (N_34667,N_32028,N_30284);
or U34668 (N_34668,N_32210,N_30549);
nor U34669 (N_34669,N_30688,N_32420);
xnor U34670 (N_34670,N_32184,N_31350);
nor U34671 (N_34671,N_31512,N_31373);
nand U34672 (N_34672,N_31719,N_31834);
nor U34673 (N_34673,N_31593,N_30925);
nand U34674 (N_34674,N_32082,N_32157);
xnor U34675 (N_34675,N_32035,N_30749);
and U34676 (N_34676,N_31424,N_30044);
nor U34677 (N_34677,N_31635,N_30991);
and U34678 (N_34678,N_32257,N_32099);
nand U34679 (N_34679,N_30615,N_31181);
nand U34680 (N_34680,N_30511,N_32124);
nor U34681 (N_34681,N_32187,N_30178);
xor U34682 (N_34682,N_30875,N_30670);
nand U34683 (N_34683,N_30269,N_31737);
and U34684 (N_34684,N_30755,N_31020);
xor U34685 (N_34685,N_31094,N_31891);
nor U34686 (N_34686,N_30280,N_30733);
or U34687 (N_34687,N_31986,N_32010);
and U34688 (N_34688,N_31824,N_31941);
nor U34689 (N_34689,N_30237,N_30800);
or U34690 (N_34690,N_30082,N_30705);
nor U34691 (N_34691,N_32119,N_32323);
and U34692 (N_34692,N_31888,N_31087);
or U34693 (N_34693,N_30424,N_32422);
xor U34694 (N_34694,N_30802,N_30561);
xnor U34695 (N_34695,N_31722,N_30863);
or U34696 (N_34696,N_30260,N_31906);
or U34697 (N_34697,N_31518,N_31403);
nor U34698 (N_34698,N_31626,N_31286);
xor U34699 (N_34699,N_32051,N_32299);
xnor U34700 (N_34700,N_30653,N_30820);
xor U34701 (N_34701,N_30054,N_30943);
xor U34702 (N_34702,N_32327,N_30596);
xor U34703 (N_34703,N_32361,N_31264);
or U34704 (N_34704,N_30693,N_31323);
or U34705 (N_34705,N_30433,N_31041);
xnor U34706 (N_34706,N_30313,N_31620);
nand U34707 (N_34707,N_30870,N_31482);
nand U34708 (N_34708,N_31714,N_32462);
xor U34709 (N_34709,N_30798,N_32295);
and U34710 (N_34710,N_30879,N_30398);
xor U34711 (N_34711,N_32007,N_30831);
nand U34712 (N_34712,N_31669,N_31933);
xnor U34713 (N_34713,N_30357,N_31206);
and U34714 (N_34714,N_30964,N_31838);
nand U34715 (N_34715,N_31223,N_30254);
nor U34716 (N_34716,N_30186,N_31348);
or U34717 (N_34717,N_31666,N_32362);
and U34718 (N_34718,N_31509,N_32033);
and U34719 (N_34719,N_32005,N_31181);
xnor U34720 (N_34720,N_31938,N_30052);
xor U34721 (N_34721,N_32155,N_31958);
xnor U34722 (N_34722,N_31995,N_30038);
and U34723 (N_34723,N_30866,N_32145);
and U34724 (N_34724,N_30320,N_30021);
nand U34725 (N_34725,N_31692,N_30465);
or U34726 (N_34726,N_30879,N_30015);
and U34727 (N_34727,N_31006,N_30889);
and U34728 (N_34728,N_32239,N_32059);
nand U34729 (N_34729,N_30583,N_30250);
nand U34730 (N_34730,N_31437,N_30810);
and U34731 (N_34731,N_31684,N_32083);
and U34732 (N_34732,N_32154,N_32407);
nor U34733 (N_34733,N_32357,N_30901);
or U34734 (N_34734,N_32313,N_30229);
nand U34735 (N_34735,N_32413,N_31144);
and U34736 (N_34736,N_30050,N_30335);
xor U34737 (N_34737,N_31403,N_31915);
nand U34738 (N_34738,N_31465,N_32438);
nor U34739 (N_34739,N_30906,N_31799);
and U34740 (N_34740,N_32003,N_30831);
and U34741 (N_34741,N_30974,N_31910);
nand U34742 (N_34742,N_32144,N_32062);
or U34743 (N_34743,N_32415,N_30405);
xor U34744 (N_34744,N_30408,N_32461);
nor U34745 (N_34745,N_31825,N_30999);
nand U34746 (N_34746,N_32271,N_32341);
xor U34747 (N_34747,N_30474,N_32349);
nor U34748 (N_34748,N_31702,N_32267);
and U34749 (N_34749,N_31967,N_30132);
nand U34750 (N_34750,N_30829,N_32003);
or U34751 (N_34751,N_31622,N_30484);
nand U34752 (N_34752,N_31340,N_31122);
or U34753 (N_34753,N_30461,N_32325);
nor U34754 (N_34754,N_31421,N_31847);
or U34755 (N_34755,N_31292,N_31402);
xor U34756 (N_34756,N_31821,N_32392);
or U34757 (N_34757,N_32084,N_31024);
nand U34758 (N_34758,N_30353,N_31177);
xor U34759 (N_34759,N_31814,N_30877);
xnor U34760 (N_34760,N_30360,N_32487);
and U34761 (N_34761,N_31797,N_32014);
nand U34762 (N_34762,N_30108,N_32327);
or U34763 (N_34763,N_31263,N_31373);
or U34764 (N_34764,N_30667,N_30844);
or U34765 (N_34765,N_31946,N_31829);
or U34766 (N_34766,N_31054,N_30101);
and U34767 (N_34767,N_30680,N_32495);
or U34768 (N_34768,N_30609,N_31994);
nand U34769 (N_34769,N_31940,N_30193);
nor U34770 (N_34770,N_32332,N_30220);
or U34771 (N_34771,N_32357,N_32118);
or U34772 (N_34772,N_31709,N_31495);
nand U34773 (N_34773,N_30784,N_31848);
or U34774 (N_34774,N_30774,N_31776);
or U34775 (N_34775,N_30453,N_31590);
or U34776 (N_34776,N_30085,N_30154);
nand U34777 (N_34777,N_31929,N_32273);
or U34778 (N_34778,N_30130,N_30066);
and U34779 (N_34779,N_31359,N_30742);
or U34780 (N_34780,N_30574,N_31849);
nor U34781 (N_34781,N_31468,N_30286);
xor U34782 (N_34782,N_32302,N_32083);
or U34783 (N_34783,N_30253,N_30639);
and U34784 (N_34784,N_31974,N_31561);
nand U34785 (N_34785,N_30088,N_30524);
xor U34786 (N_34786,N_31948,N_31617);
nor U34787 (N_34787,N_31662,N_31161);
nor U34788 (N_34788,N_31449,N_31493);
xnor U34789 (N_34789,N_32007,N_30092);
nand U34790 (N_34790,N_31707,N_31351);
xor U34791 (N_34791,N_31244,N_31486);
xnor U34792 (N_34792,N_31793,N_30170);
xnor U34793 (N_34793,N_32012,N_31831);
or U34794 (N_34794,N_30106,N_31217);
nor U34795 (N_34795,N_31123,N_30502);
or U34796 (N_34796,N_32191,N_30224);
nor U34797 (N_34797,N_32048,N_31356);
nand U34798 (N_34798,N_31736,N_30104);
nor U34799 (N_34799,N_32026,N_30623);
or U34800 (N_34800,N_30540,N_32401);
xnor U34801 (N_34801,N_31437,N_32458);
and U34802 (N_34802,N_32336,N_32342);
and U34803 (N_34803,N_30720,N_30182);
xor U34804 (N_34804,N_31966,N_31710);
xnor U34805 (N_34805,N_31254,N_32349);
or U34806 (N_34806,N_31552,N_32192);
nor U34807 (N_34807,N_30565,N_30000);
nor U34808 (N_34808,N_30706,N_31254);
or U34809 (N_34809,N_30186,N_30271);
and U34810 (N_34810,N_30223,N_31456);
nor U34811 (N_34811,N_31708,N_31540);
xnor U34812 (N_34812,N_31714,N_31156);
nand U34813 (N_34813,N_31744,N_30991);
nor U34814 (N_34814,N_31085,N_31049);
and U34815 (N_34815,N_31595,N_32209);
nor U34816 (N_34816,N_31809,N_30413);
nor U34817 (N_34817,N_30718,N_32180);
xor U34818 (N_34818,N_30945,N_31255);
xnor U34819 (N_34819,N_32150,N_32233);
or U34820 (N_34820,N_30673,N_31371);
nor U34821 (N_34821,N_31796,N_32496);
nor U34822 (N_34822,N_30706,N_31189);
and U34823 (N_34823,N_32489,N_30996);
xnor U34824 (N_34824,N_30781,N_31678);
nand U34825 (N_34825,N_32446,N_30208);
and U34826 (N_34826,N_32195,N_31732);
or U34827 (N_34827,N_30866,N_32162);
xnor U34828 (N_34828,N_31837,N_32009);
xnor U34829 (N_34829,N_30037,N_30628);
or U34830 (N_34830,N_30863,N_32221);
xnor U34831 (N_34831,N_31725,N_30151);
or U34832 (N_34832,N_30016,N_31694);
xor U34833 (N_34833,N_31997,N_30889);
and U34834 (N_34834,N_32278,N_30487);
xor U34835 (N_34835,N_30645,N_30944);
or U34836 (N_34836,N_31776,N_31790);
nor U34837 (N_34837,N_30001,N_31276);
and U34838 (N_34838,N_30482,N_30208);
or U34839 (N_34839,N_31490,N_30438);
nor U34840 (N_34840,N_30567,N_32006);
or U34841 (N_34841,N_31783,N_30262);
nor U34842 (N_34842,N_32440,N_32072);
nand U34843 (N_34843,N_32489,N_31181);
nand U34844 (N_34844,N_31892,N_31906);
nand U34845 (N_34845,N_31542,N_30018);
nor U34846 (N_34846,N_31498,N_31394);
nor U34847 (N_34847,N_30827,N_30244);
xnor U34848 (N_34848,N_31686,N_31288);
nor U34849 (N_34849,N_30788,N_30497);
or U34850 (N_34850,N_31841,N_30683);
nor U34851 (N_34851,N_30834,N_30516);
nor U34852 (N_34852,N_30233,N_31330);
nand U34853 (N_34853,N_30906,N_31728);
or U34854 (N_34854,N_31494,N_31394);
xnor U34855 (N_34855,N_31609,N_31073);
nor U34856 (N_34856,N_30695,N_30054);
xor U34857 (N_34857,N_30167,N_30041);
xnor U34858 (N_34858,N_31801,N_31617);
nand U34859 (N_34859,N_30823,N_30941);
nor U34860 (N_34860,N_31195,N_30583);
and U34861 (N_34861,N_30437,N_31235);
or U34862 (N_34862,N_31319,N_30641);
xnor U34863 (N_34863,N_31095,N_32289);
xnor U34864 (N_34864,N_31594,N_31918);
xnor U34865 (N_34865,N_31900,N_31429);
and U34866 (N_34866,N_32123,N_30779);
and U34867 (N_34867,N_32305,N_31441);
and U34868 (N_34868,N_31252,N_30601);
and U34869 (N_34869,N_30276,N_31680);
nand U34870 (N_34870,N_32168,N_30294);
nand U34871 (N_34871,N_31583,N_31349);
xnor U34872 (N_34872,N_31998,N_30156);
or U34873 (N_34873,N_30855,N_30691);
or U34874 (N_34874,N_30880,N_31551);
or U34875 (N_34875,N_31296,N_32364);
or U34876 (N_34876,N_30016,N_30260);
or U34877 (N_34877,N_30205,N_31554);
nand U34878 (N_34878,N_30588,N_30328);
nor U34879 (N_34879,N_32315,N_30026);
xnor U34880 (N_34880,N_30630,N_30560);
and U34881 (N_34881,N_31915,N_30207);
nor U34882 (N_34882,N_31613,N_32444);
or U34883 (N_34883,N_30766,N_32428);
or U34884 (N_34884,N_30301,N_31196);
xor U34885 (N_34885,N_31663,N_31937);
and U34886 (N_34886,N_32221,N_32068);
nor U34887 (N_34887,N_30901,N_30644);
xnor U34888 (N_34888,N_31869,N_31698);
and U34889 (N_34889,N_32317,N_32164);
or U34890 (N_34890,N_30721,N_30832);
nor U34891 (N_34891,N_31639,N_31446);
nand U34892 (N_34892,N_32050,N_32070);
nand U34893 (N_34893,N_30698,N_31451);
or U34894 (N_34894,N_30772,N_31047);
nand U34895 (N_34895,N_30508,N_32291);
or U34896 (N_34896,N_32485,N_32428);
nor U34897 (N_34897,N_30615,N_31206);
xor U34898 (N_34898,N_32176,N_32206);
nor U34899 (N_34899,N_31925,N_30245);
nand U34900 (N_34900,N_30277,N_32294);
and U34901 (N_34901,N_30847,N_30579);
nand U34902 (N_34902,N_32373,N_31031);
or U34903 (N_34903,N_30392,N_32404);
or U34904 (N_34904,N_31953,N_32212);
nor U34905 (N_34905,N_30457,N_31551);
and U34906 (N_34906,N_31930,N_31371);
nand U34907 (N_34907,N_30309,N_30143);
nor U34908 (N_34908,N_30126,N_30635);
nand U34909 (N_34909,N_30015,N_30207);
and U34910 (N_34910,N_30053,N_31873);
or U34911 (N_34911,N_31364,N_32440);
nor U34912 (N_34912,N_31369,N_31990);
nor U34913 (N_34913,N_31389,N_30532);
xor U34914 (N_34914,N_30046,N_32201);
nor U34915 (N_34915,N_30898,N_30626);
xnor U34916 (N_34916,N_31649,N_32391);
and U34917 (N_34917,N_32473,N_32456);
nor U34918 (N_34918,N_30271,N_31443);
and U34919 (N_34919,N_32308,N_30300);
or U34920 (N_34920,N_30729,N_30298);
and U34921 (N_34921,N_30207,N_30017);
or U34922 (N_34922,N_30955,N_31164);
and U34923 (N_34923,N_30626,N_30518);
nand U34924 (N_34924,N_31114,N_32103);
or U34925 (N_34925,N_30486,N_30023);
and U34926 (N_34926,N_30192,N_31453);
or U34927 (N_34927,N_32038,N_31426);
or U34928 (N_34928,N_31911,N_30715);
nor U34929 (N_34929,N_30256,N_32276);
and U34930 (N_34930,N_32005,N_30058);
or U34931 (N_34931,N_31381,N_30827);
xnor U34932 (N_34932,N_32185,N_30950);
xor U34933 (N_34933,N_30727,N_30726);
and U34934 (N_34934,N_32013,N_31867);
xnor U34935 (N_34935,N_30098,N_30506);
and U34936 (N_34936,N_31895,N_30907);
or U34937 (N_34937,N_32489,N_30145);
and U34938 (N_34938,N_30888,N_31488);
nor U34939 (N_34939,N_32006,N_31351);
nor U34940 (N_34940,N_32021,N_30750);
xnor U34941 (N_34941,N_30149,N_30426);
xnor U34942 (N_34942,N_30828,N_31548);
xnor U34943 (N_34943,N_31195,N_31296);
and U34944 (N_34944,N_31346,N_32083);
nand U34945 (N_34945,N_30165,N_31329);
xnor U34946 (N_34946,N_31776,N_30510);
or U34947 (N_34947,N_30171,N_31117);
and U34948 (N_34948,N_31457,N_30857);
xor U34949 (N_34949,N_32215,N_31259);
or U34950 (N_34950,N_30477,N_32110);
xor U34951 (N_34951,N_31791,N_31643);
nor U34952 (N_34952,N_32327,N_32082);
and U34953 (N_34953,N_30871,N_31602);
nor U34954 (N_34954,N_31299,N_32285);
nor U34955 (N_34955,N_31442,N_32252);
and U34956 (N_34956,N_30178,N_30452);
nor U34957 (N_34957,N_30929,N_30234);
xor U34958 (N_34958,N_31878,N_31468);
nor U34959 (N_34959,N_31476,N_30059);
or U34960 (N_34960,N_31767,N_31953);
nor U34961 (N_34961,N_30449,N_30222);
or U34962 (N_34962,N_31267,N_30340);
and U34963 (N_34963,N_30366,N_30332);
or U34964 (N_34964,N_31347,N_30052);
nand U34965 (N_34965,N_32234,N_30441);
nand U34966 (N_34966,N_30763,N_30028);
or U34967 (N_34967,N_32290,N_30707);
or U34968 (N_34968,N_31076,N_32147);
and U34969 (N_34969,N_31373,N_30398);
nor U34970 (N_34970,N_30106,N_30032);
nand U34971 (N_34971,N_31285,N_32037);
xor U34972 (N_34972,N_30647,N_30164);
xor U34973 (N_34973,N_30374,N_30760);
nor U34974 (N_34974,N_32266,N_31572);
and U34975 (N_34975,N_32084,N_31177);
and U34976 (N_34976,N_31041,N_30852);
or U34977 (N_34977,N_31290,N_31845);
nand U34978 (N_34978,N_30552,N_31200);
xor U34979 (N_34979,N_30464,N_30203);
nor U34980 (N_34980,N_30566,N_30575);
nor U34981 (N_34981,N_32300,N_32163);
or U34982 (N_34982,N_32375,N_31933);
nand U34983 (N_34983,N_31281,N_31369);
or U34984 (N_34984,N_30372,N_31576);
nor U34985 (N_34985,N_32417,N_31466);
or U34986 (N_34986,N_31947,N_32407);
xnor U34987 (N_34987,N_32139,N_32453);
xnor U34988 (N_34988,N_30410,N_30042);
nand U34989 (N_34989,N_31485,N_30632);
and U34990 (N_34990,N_32231,N_30119);
or U34991 (N_34991,N_30123,N_32479);
nor U34992 (N_34992,N_31595,N_32449);
xnor U34993 (N_34993,N_32494,N_32131);
nor U34994 (N_34994,N_31184,N_30103);
nand U34995 (N_34995,N_31277,N_31365);
xor U34996 (N_34996,N_30859,N_31265);
or U34997 (N_34997,N_32496,N_30671);
or U34998 (N_34998,N_31768,N_30621);
nor U34999 (N_34999,N_30618,N_30735);
nand U35000 (N_35000,N_32543,N_33987);
nand U35001 (N_35001,N_33612,N_33756);
and U35002 (N_35002,N_33947,N_34812);
xor U35003 (N_35003,N_34224,N_34593);
and U35004 (N_35004,N_34785,N_32584);
nand U35005 (N_35005,N_33480,N_34118);
and U35006 (N_35006,N_34390,N_33727);
nor U35007 (N_35007,N_34730,N_33151);
nand U35008 (N_35008,N_33616,N_33690);
xnor U35009 (N_35009,N_33767,N_33092);
nor U35010 (N_35010,N_33447,N_34635);
xor U35011 (N_35011,N_33420,N_33649);
xnor U35012 (N_35012,N_33923,N_33744);
or U35013 (N_35013,N_34962,N_34333);
or U35014 (N_35014,N_32866,N_33951);
and U35015 (N_35015,N_34692,N_32669);
nand U35016 (N_35016,N_32536,N_34285);
and U35017 (N_35017,N_34819,N_33816);
xnor U35018 (N_35018,N_33541,N_34493);
nor U35019 (N_35019,N_34013,N_34765);
nor U35020 (N_35020,N_34791,N_33419);
or U35021 (N_35021,N_34180,N_33027);
and U35022 (N_35022,N_34469,N_33320);
nand U35023 (N_35023,N_33554,N_33812);
and U35024 (N_35024,N_34039,N_33835);
and U35025 (N_35025,N_33721,N_34214);
nor U35026 (N_35026,N_33709,N_34426);
nor U35027 (N_35027,N_33280,N_34682);
and U35028 (N_35028,N_34746,N_33393);
nand U35029 (N_35029,N_34826,N_33982);
nand U35030 (N_35030,N_33441,N_34919);
or U35031 (N_35031,N_32708,N_32966);
nor U35032 (N_35032,N_33518,N_34782);
nand U35033 (N_35033,N_32995,N_32632);
and U35034 (N_35034,N_33636,N_34632);
and U35035 (N_35035,N_33907,N_34450);
nor U35036 (N_35036,N_32733,N_32820);
and U35037 (N_35037,N_33196,N_34492);
nor U35038 (N_35038,N_34095,N_34773);
nor U35039 (N_35039,N_33378,N_33657);
nand U35040 (N_35040,N_33400,N_34953);
xnor U35041 (N_35041,N_34136,N_33857);
nand U35042 (N_35042,N_33736,N_34551);
or U35043 (N_35043,N_34975,N_34293);
nand U35044 (N_35044,N_33183,N_34689);
and U35045 (N_35045,N_32519,N_33574);
nor U35046 (N_35046,N_33549,N_32975);
xor U35047 (N_35047,N_34631,N_34092);
nand U35048 (N_35048,N_32715,N_34575);
or U35049 (N_35049,N_34318,N_33137);
or U35050 (N_35050,N_32647,N_34900);
nor U35051 (N_35051,N_32904,N_34604);
and U35052 (N_35052,N_33954,N_34438);
nor U35053 (N_35053,N_34662,N_33846);
nand U35054 (N_35054,N_33314,N_33429);
nand U35055 (N_35055,N_33012,N_34643);
nand U35056 (N_35056,N_32730,N_34331);
xnor U35057 (N_35057,N_32711,N_34183);
or U35058 (N_35058,N_34208,N_34741);
and U35059 (N_35059,N_34146,N_34673);
and U35060 (N_35060,N_33208,N_33459);
xnor U35061 (N_35061,N_32668,N_32795);
nor U35062 (N_35062,N_34994,N_32874);
or U35063 (N_35063,N_34802,N_33868);
xor U35064 (N_35064,N_33808,N_34622);
xor U35065 (N_35065,N_34553,N_32852);
or U35066 (N_35066,N_34442,N_32681);
or U35067 (N_35067,N_33089,N_33482);
xor U35068 (N_35068,N_33953,N_34577);
or U35069 (N_35069,N_33837,N_32687);
or U35070 (N_35070,N_32801,N_34102);
and U35071 (N_35071,N_33638,N_33057);
and U35072 (N_35072,N_32812,N_32593);
nand U35073 (N_35073,N_34235,N_33859);
or U35074 (N_35074,N_34656,N_33567);
nor U35075 (N_35075,N_33527,N_34592);
nor U35076 (N_35076,N_34532,N_33855);
and U35077 (N_35077,N_33038,N_32685);
nor U35078 (N_35078,N_33738,N_34565);
nor U35079 (N_35079,N_34211,N_33087);
or U35080 (N_35080,N_34361,N_32809);
or U35081 (N_35081,N_33271,N_32581);
nand U35082 (N_35082,N_34941,N_33720);
nand U35083 (N_35083,N_33064,N_34357);
nand U35084 (N_35084,N_34713,N_33002);
and U35085 (N_35085,N_32684,N_33413);
nor U35086 (N_35086,N_33747,N_33559);
or U35087 (N_35087,N_32773,N_34836);
nand U35088 (N_35088,N_32533,N_33056);
xnor U35089 (N_35089,N_32744,N_34248);
or U35090 (N_35090,N_33160,N_33509);
and U35091 (N_35091,N_34083,N_34174);
xnor U35092 (N_35092,N_32695,N_33239);
xnor U35093 (N_35093,N_33798,N_32784);
and U35094 (N_35094,N_33524,N_34723);
nand U35095 (N_35095,N_34720,N_33202);
nor U35096 (N_35096,N_34396,N_33123);
nor U35097 (N_35097,N_34987,N_32527);
nand U35098 (N_35098,N_34144,N_33799);
xnor U35099 (N_35099,N_34311,N_33753);
or U35100 (N_35100,N_33237,N_33935);
xnor U35101 (N_35101,N_33316,N_34574);
or U35102 (N_35102,N_34959,N_32909);
or U35103 (N_35103,N_34230,N_33508);
xor U35104 (N_35104,N_33504,N_33981);
or U35105 (N_35105,N_34965,N_33725);
xor U35106 (N_35106,N_33354,N_34718);
nand U35107 (N_35107,N_32511,N_33689);
or U35108 (N_35108,N_34456,N_34536);
or U35109 (N_35109,N_34849,N_33368);
nor U35110 (N_35110,N_34704,N_34940);
xor U35111 (N_35111,N_33888,N_33604);
xor U35112 (N_35112,N_34087,N_34885);
and U35113 (N_35113,N_33333,N_33204);
and U35114 (N_35114,N_34863,N_32549);
and U35115 (N_35115,N_33172,N_33005);
xor U35116 (N_35116,N_32792,N_33807);
or U35117 (N_35117,N_34925,N_34217);
xor U35118 (N_35118,N_32580,N_34984);
xor U35119 (N_35119,N_33860,N_33464);
nand U35120 (N_35120,N_34666,N_33376);
or U35121 (N_35121,N_34362,N_33742);
or U35122 (N_35122,N_34758,N_34249);
nor U35123 (N_35123,N_34529,N_34800);
xnor U35124 (N_35124,N_33884,N_33593);
nor U35125 (N_35125,N_33676,N_33283);
xor U35126 (N_35126,N_32918,N_34937);
or U35127 (N_35127,N_32919,N_34322);
nand U35128 (N_35128,N_33372,N_32845);
and U35129 (N_35129,N_32888,N_33922);
nor U35130 (N_35130,N_32547,N_34088);
nand U35131 (N_35131,N_34245,N_33406);
xnor U35132 (N_35132,N_33847,N_34910);
nor U35133 (N_35133,N_34147,N_33820);
xor U35134 (N_35134,N_33402,N_34848);
nand U35135 (N_35135,N_32528,N_34295);
xnor U35136 (N_35136,N_34058,N_34290);
nor U35137 (N_35137,N_33531,N_33957);
xnor U35138 (N_35138,N_34204,N_34124);
nand U35139 (N_35139,N_34268,N_33295);
xnor U35140 (N_35140,N_33519,N_34015);
or U35141 (N_35141,N_33737,N_32651);
or U35142 (N_35142,N_32885,N_33805);
xnor U35143 (N_35143,N_33457,N_33181);
and U35144 (N_35144,N_33887,N_34133);
and U35145 (N_35145,N_32783,N_33018);
and U35146 (N_35146,N_34415,N_34363);
nor U35147 (N_35147,N_33908,N_33249);
or U35148 (N_35148,N_34379,N_32623);
nand U35149 (N_35149,N_34862,N_33793);
and U35150 (N_35150,N_33227,N_32871);
nor U35151 (N_35151,N_33153,N_34184);
nand U35152 (N_35152,N_34664,N_33770);
xor U35153 (N_35153,N_32825,N_33804);
xor U35154 (N_35154,N_34710,N_33111);
nor U35155 (N_35155,N_34513,N_33124);
or U35156 (N_35156,N_34467,N_32940);
xnor U35157 (N_35157,N_33363,N_33833);
and U35158 (N_35158,N_33155,N_33041);
and U35159 (N_35159,N_33296,N_33886);
xor U35160 (N_35160,N_34423,N_34961);
or U35161 (N_35161,N_34639,N_32564);
nor U35162 (N_35162,N_34891,N_34884);
and U35163 (N_35163,N_33544,N_32794);
nand U35164 (N_35164,N_33061,N_33517);
or U35165 (N_35165,N_34296,N_34756);
xor U35166 (N_35166,N_32804,N_34552);
and U35167 (N_35167,N_33337,N_33060);
xor U35168 (N_35168,N_34271,N_34827);
or U35169 (N_35169,N_34353,N_34135);
xor U35170 (N_35170,N_32810,N_34657);
and U35171 (N_35171,N_33199,N_34914);
nor U35172 (N_35172,N_33562,N_34864);
and U35173 (N_35173,N_32726,N_34612);
xor U35174 (N_35174,N_34138,N_33017);
xor U35175 (N_35175,N_33465,N_33302);
nand U35176 (N_35176,N_32611,N_33255);
and U35177 (N_35177,N_33339,N_33161);
or U35178 (N_35178,N_34518,N_32878);
or U35179 (N_35179,N_32709,N_33543);
xnor U35180 (N_35180,N_33881,N_32513);
xor U35181 (N_35181,N_33022,N_32501);
and U35182 (N_35182,N_33252,N_34549);
and U35183 (N_35183,N_33547,N_33775);
and U35184 (N_35184,N_33150,N_33746);
and U35185 (N_35185,N_34276,N_33421);
and U35186 (N_35186,N_34070,N_34610);
and U35187 (N_35187,N_32544,N_34150);
nor U35188 (N_35188,N_33462,N_34957);
or U35189 (N_35189,N_34561,N_34403);
and U35190 (N_35190,N_33755,N_32911);
or U35191 (N_35191,N_32831,N_34227);
and U35192 (N_35192,N_32616,N_34752);
or U35193 (N_35193,N_34137,N_34619);
or U35194 (N_35194,N_34648,N_33872);
nand U35195 (N_35195,N_34808,N_33079);
xor U35196 (N_35196,N_34834,N_33620);
and U35197 (N_35197,N_34097,N_32900);
and U35198 (N_35198,N_34428,N_33307);
nor U35199 (N_35199,N_34743,N_33588);
or U35200 (N_35200,N_34901,N_32968);
and U35201 (N_35201,N_32816,N_34742);
xor U35202 (N_35202,N_33810,N_32908);
nor U35203 (N_35203,N_33502,N_33309);
xor U35204 (N_35204,N_34120,N_33630);
nor U35205 (N_35205,N_34778,N_34371);
nand U35206 (N_35206,N_32659,N_33545);
or U35207 (N_35207,N_33900,N_33511);
or U35208 (N_35208,N_34906,N_34392);
nor U35209 (N_35209,N_33093,N_33594);
and U35210 (N_35210,N_34308,N_32850);
and U35211 (N_35211,N_34062,N_33539);
xor U35212 (N_35212,N_32673,N_32741);
xor U35213 (N_35213,N_34907,N_32987);
xnor U35214 (N_35214,N_34236,N_33234);
and U35215 (N_35215,N_33282,N_34745);
and U35216 (N_35216,N_32592,N_33156);
nor U35217 (N_35217,N_34942,N_33285);
or U35218 (N_35218,N_34776,N_33577);
or U35219 (N_35219,N_34929,N_32525);
nor U35220 (N_35220,N_33455,N_33563);
and U35221 (N_35221,N_32742,N_34094);
and U35222 (N_35222,N_33780,N_33047);
and U35223 (N_35223,N_32808,N_32548);
and U35224 (N_35224,N_34559,N_33409);
or U35225 (N_35225,N_32759,N_34568);
or U35226 (N_35226,N_33965,N_32969);
nand U35227 (N_35227,N_33351,N_32563);
and U35228 (N_35228,N_34668,N_34048);
nor U35229 (N_35229,N_33347,N_34508);
nor U35230 (N_35230,N_32999,N_34177);
nand U35231 (N_35231,N_34916,N_34754);
or U35232 (N_35232,N_34455,N_33814);
nor U35233 (N_35233,N_33090,N_33401);
and U35234 (N_35234,N_34524,N_34626);
nor U35235 (N_35235,N_32596,N_33381);
xnor U35236 (N_35236,N_33412,N_33197);
and U35237 (N_35237,N_32614,N_33146);
or U35238 (N_35238,N_33829,N_34496);
nor U35239 (N_35239,N_33203,N_33792);
or U35240 (N_35240,N_34020,N_32841);
or U35241 (N_35241,N_33344,N_33443);
xor U35242 (N_35242,N_32806,N_33450);
xnor U35243 (N_35243,N_34878,N_32587);
and U35244 (N_35244,N_33077,N_33743);
nor U35245 (N_35245,N_34859,N_34918);
nor U35246 (N_35246,N_34931,N_34380);
and U35247 (N_35247,N_32601,N_34465);
xnor U35248 (N_35248,N_33879,N_34867);
nor U35249 (N_35249,N_34797,N_34328);
nor U35250 (N_35250,N_34176,N_34952);
xor U35251 (N_35251,N_34820,N_34943);
nor U35252 (N_35252,N_33537,N_34385);
xor U35253 (N_35253,N_32579,N_34044);
xor U35254 (N_35254,N_33542,N_32644);
xnor U35255 (N_35255,N_33745,N_32504);
and U35256 (N_35256,N_32722,N_32857);
and U35257 (N_35257,N_34468,N_34521);
nand U35258 (N_35258,N_32760,N_33417);
or U35259 (N_35259,N_34163,N_33610);
and U35260 (N_35260,N_34696,N_34882);
and U35261 (N_35261,N_32824,N_32849);
xnor U35262 (N_35262,N_34375,N_34072);
nor U35263 (N_35263,N_33867,N_34338);
xor U35264 (N_35264,N_32858,N_34016);
and U35265 (N_35265,N_34181,N_34169);
or U35266 (N_35266,N_33374,N_33717);
xor U35267 (N_35267,N_33882,N_34125);
xnor U35268 (N_35268,N_33692,N_34410);
and U35269 (N_35269,N_34772,N_33176);
nand U35270 (N_35270,N_34935,N_33434);
or U35271 (N_35271,N_32807,N_34527);
xor U35272 (N_35272,N_33048,N_34924);
or U35273 (N_35273,N_34413,N_34414);
nand U35274 (N_35274,N_33473,N_33582);
xor U35275 (N_35275,N_32833,N_34749);
nand U35276 (N_35276,N_34425,N_34241);
xor U35277 (N_35277,N_34434,N_32901);
nor U35278 (N_35278,N_33201,N_34326);
nand U35279 (N_35279,N_33139,N_32518);
nor U35280 (N_35280,N_32646,N_33754);
or U35281 (N_35281,N_33325,N_33110);
or U35282 (N_35282,N_34903,N_34126);
nor U35283 (N_35283,N_32855,N_32671);
and U35284 (N_35284,N_34578,N_32972);
nand U35285 (N_35285,N_33468,N_32713);
or U35286 (N_35286,N_34708,N_34621);
or U35287 (N_35287,N_34860,N_34011);
nand U35288 (N_35288,N_34499,N_33033);
nand U35289 (N_35289,N_34277,N_34106);
xor U35290 (N_35290,N_33532,N_34437);
nand U35291 (N_35291,N_33379,N_34764);
xnor U35292 (N_35292,N_33865,N_33335);
and U35293 (N_35293,N_34793,N_34075);
xnor U35294 (N_35294,N_33983,N_34642);
or U35295 (N_35295,N_33758,N_33261);
nand U35296 (N_35296,N_33587,N_32771);
and U35297 (N_35297,N_32949,N_33605);
nand U35298 (N_35298,N_33192,N_33822);
xor U35299 (N_35299,N_34402,N_34400);
nand U35300 (N_35300,N_33693,N_33037);
or U35301 (N_35301,N_34654,N_34037);
and U35302 (N_35302,N_34922,N_33100);
nand U35303 (N_35303,N_32943,N_33084);
nor U35304 (N_35304,N_33315,N_32750);
and U35305 (N_35305,N_34003,N_33205);
xor U35306 (N_35306,N_32802,N_33677);
nor U35307 (N_35307,N_32755,N_33575);
or U35308 (N_35308,N_32923,N_34395);
nor U35309 (N_35309,N_34387,N_34525);
xnor U35310 (N_35310,N_34783,N_32590);
xnor U35311 (N_35311,N_33453,N_33890);
or U35312 (N_35312,N_34556,N_32512);
nor U35313 (N_35313,N_34669,N_33704);
and U35314 (N_35314,N_34355,N_32641);
or U35315 (N_35315,N_32546,N_34405);
and U35316 (N_35316,N_34875,N_34844);
and U35317 (N_35317,N_34085,N_34790);
nand U35318 (N_35318,N_32690,N_32656);
and U35319 (N_35319,N_34634,N_33903);
and U35320 (N_35320,N_34131,N_32682);
nand U35321 (N_35321,N_32558,N_33422);
nor U35322 (N_35322,N_34339,N_34832);
or U35323 (N_35323,N_33842,N_33134);
nand U35324 (N_35324,N_32840,N_33186);
and U35325 (N_35325,N_33643,N_32848);
xnor U35326 (N_35326,N_33169,N_33926);
xor U35327 (N_35327,N_32550,N_32844);
nand U35328 (N_35328,N_33287,N_33757);
nand U35329 (N_35329,N_32936,N_33278);
and U35330 (N_35330,N_34300,N_34411);
nand U35331 (N_35331,N_32986,N_34000);
xnor U35332 (N_35332,N_34596,N_34307);
nand U35333 (N_35333,N_34107,N_33556);
xnor U35334 (N_35334,N_32775,N_33941);
xnor U35335 (N_35335,N_34419,N_34917);
nor U35336 (N_35336,N_32798,N_34650);
nor U35337 (N_35337,N_33839,N_34841);
nor U35338 (N_35338,N_33942,N_33963);
xor U35339 (N_35339,N_34737,N_33584);
or U35340 (N_35340,N_33332,N_32612);
and U35341 (N_35341,N_34356,N_33003);
xor U35342 (N_35342,N_33385,N_32891);
xor U35343 (N_35343,N_33329,N_33218);
or U35344 (N_35344,N_34829,N_32754);
xnor U35345 (N_35345,N_32572,N_34550);
xnor U35346 (N_35346,N_33581,N_32516);
nand U35347 (N_35347,N_33991,N_33066);
xor U35348 (N_35348,N_33711,N_34047);
and U35349 (N_35349,N_34201,N_34658);
xnor U35350 (N_35350,N_33439,N_33485);
nand U35351 (N_35351,N_34341,N_34698);
xor U35352 (N_35352,N_33722,N_33328);
nand U35353 (N_35353,N_34024,N_34872);
nor U35354 (N_35354,N_34580,N_33708);
nor U35355 (N_35355,N_34449,N_32799);
nor U35356 (N_35356,N_33533,N_33477);
and U35357 (N_35357,N_33794,N_34284);
or U35358 (N_35358,N_34771,N_34694);
and U35359 (N_35359,N_34190,N_34576);
nor U35360 (N_35360,N_34343,N_34850);
and U35361 (N_35361,N_34351,N_33850);
nor U35362 (N_35362,N_34494,N_33784);
nor U35363 (N_35363,N_34420,N_34287);
nor U35364 (N_35364,N_34195,N_34971);
nand U35365 (N_35365,N_33592,N_34223);
nand U35366 (N_35366,N_34546,N_32836);
or U35367 (N_35367,N_32663,N_33341);
and U35368 (N_35368,N_34686,N_32745);
nand U35369 (N_35369,N_34096,N_34555);
xnor U35370 (N_35370,N_34335,N_33553);
nor U35371 (N_35371,N_34346,N_32915);
nor U35372 (N_35372,N_33896,N_32961);
nor U35373 (N_35373,N_33613,N_33040);
nor U35374 (N_35374,N_34286,N_33586);
xnor U35375 (N_35375,N_34207,N_34851);
nor U35376 (N_35376,N_33976,N_34022);
nand U35377 (N_35377,N_32560,N_33245);
and U35378 (N_35378,N_33128,N_33086);
and U35379 (N_35379,N_34283,N_32971);
and U35380 (N_35380,N_33028,N_34558);
nor U35381 (N_35381,N_33702,N_33055);
xnor U35382 (N_35382,N_34623,N_34388);
or U35383 (N_35383,N_32886,N_33371);
xor U35384 (N_35384,N_32657,N_32507);
xnor U35385 (N_35385,N_34655,N_33801);
and U35386 (N_35386,N_34842,N_32822);
nand U35387 (N_35387,N_33580,N_34838);
xor U35388 (N_35388,N_34101,N_33566);
nor U35389 (N_35389,N_34570,N_34792);
or U35390 (N_35390,N_32867,N_33108);
nand U35391 (N_35391,N_34263,N_34889);
and U35392 (N_35392,N_33797,N_34435);
nand U35393 (N_35393,N_32991,N_34534);
nor U35394 (N_35394,N_32959,N_34923);
xor U35395 (N_35395,N_32894,N_34583);
nor U35396 (N_35396,N_32803,N_34944);
nor U35397 (N_35397,N_33251,N_32985);
nand U35398 (N_35398,N_33551,N_33733);
or U35399 (N_35399,N_34004,N_33818);
and U35400 (N_35400,N_32903,N_33946);
nor U35401 (N_35401,N_33019,N_33046);
nor U35402 (N_35402,N_32719,N_33607);
or U35403 (N_35403,N_33790,N_34025);
and U35404 (N_35404,N_33303,N_32994);
or U35405 (N_35405,N_34113,N_33682);
nand U35406 (N_35406,N_34242,N_32984);
and U35407 (N_35407,N_34065,N_34701);
nand U35408 (N_35408,N_33270,N_34352);
and U35409 (N_35409,N_33555,N_32703);
xnor U35410 (N_35410,N_34837,N_33752);
nor U35411 (N_35411,N_32620,N_33297);
nor U35412 (N_35412,N_34288,N_34430);
and U35413 (N_35413,N_32977,N_33403);
nor U35414 (N_35414,N_33065,N_34168);
and U35415 (N_35415,N_32557,N_34519);
and U35416 (N_35416,N_34421,N_32860);
and U35417 (N_35417,N_32683,N_34014);
nand U35418 (N_35418,N_34833,N_32735);
nor U35419 (N_35419,N_33015,N_34377);
nor U35420 (N_35420,N_34299,N_33564);
xor U35421 (N_35421,N_33802,N_33663);
xor U35422 (N_35422,N_33821,N_33114);
and U35423 (N_35423,N_33599,N_32628);
nor U35424 (N_35424,N_33490,N_33650);
nand U35425 (N_35425,N_33062,N_33841);
and U35426 (N_35426,N_33990,N_34109);
or U35427 (N_35427,N_32594,N_33985);
xnor U35428 (N_35428,N_32751,N_33217);
nor U35429 (N_35429,N_32956,N_32827);
xor U35430 (N_35430,N_33284,N_33945);
or U35431 (N_35431,N_33142,N_33505);
and U35432 (N_35432,N_32505,N_32770);
and U35433 (N_35433,N_34151,N_33874);
nor U35434 (N_35434,N_33254,N_34074);
nor U35435 (N_35435,N_34409,N_34404);
nand U35436 (N_35436,N_33052,N_34012);
or U35437 (N_35437,N_33195,N_33349);
and U35438 (N_35438,N_32736,N_34384);
and U35439 (N_35439,N_34117,N_33917);
nor U35440 (N_35440,N_33471,N_33370);
nor U35441 (N_35441,N_34165,N_34312);
nand U35442 (N_35442,N_33398,N_33645);
xnor U35443 (N_35443,N_34586,N_32658);
nand U35444 (N_35444,N_33474,N_34157);
nand U35445 (N_35445,N_34569,N_34440);
xor U35446 (N_35446,N_32929,N_33431);
nor U35447 (N_35447,N_34946,N_33083);
nand U35448 (N_35448,N_34482,N_32749);
nor U35449 (N_35449,N_33984,N_33665);
nand U35450 (N_35450,N_33259,N_34951);
nand U35451 (N_35451,N_33488,N_33165);
or U35452 (N_35452,N_33740,N_33885);
nand U35453 (N_35453,N_34266,N_34533);
and U35454 (N_35454,N_33796,N_33787);
or U35455 (N_35455,N_33646,N_32763);
or U35456 (N_35456,N_32960,N_33904);
nand U35457 (N_35457,N_34269,N_34986);
or U35458 (N_35458,N_34877,N_33236);
xor U35459 (N_35459,N_33762,N_33826);
and U35460 (N_35460,N_32837,N_34050);
nand U35461 (N_35461,N_34777,N_32704);
and U35462 (N_35462,N_33448,N_33695);
and U35463 (N_35463,N_34049,N_34178);
nor U35464 (N_35464,N_33751,N_33813);
nor U35465 (N_35465,N_33373,N_34142);
xor U35466 (N_35466,N_33020,N_34342);
nand U35467 (N_35467,N_33127,N_32851);
xor U35468 (N_35468,N_33375,N_33070);
or U35469 (N_35469,N_34607,N_34606);
nor U35470 (N_35470,N_34077,N_33739);
xnor U35471 (N_35471,N_33726,N_34683);
nand U35472 (N_35472,N_33454,N_33873);
and U35473 (N_35473,N_33633,N_33013);
xor U35474 (N_35474,N_34590,N_33444);
or U35475 (N_35475,N_32935,N_33388);
xor U35476 (N_35476,N_34869,N_32514);
nor U35477 (N_35477,N_34264,N_34824);
xor U35478 (N_35478,N_34954,N_34731);
and U35479 (N_35479,N_32978,N_32648);
nor U35480 (N_35480,N_34712,N_34498);
nor U35481 (N_35481,N_33932,N_33656);
nand U35482 (N_35482,N_33483,N_33452);
or U35483 (N_35483,N_33119,N_32898);
xnor U35484 (N_35484,N_33618,N_33121);
nor U35485 (N_35485,N_34093,N_32666);
and U35486 (N_35486,N_33357,N_33906);
and U35487 (N_35487,N_33456,N_32702);
nor U35488 (N_35488,N_32869,N_33306);
nor U35489 (N_35489,N_33988,N_34677);
and U35490 (N_35490,N_33267,N_33809);
nand U35491 (N_35491,N_34002,N_32665);
or U35492 (N_35492,N_33094,N_32862);
nand U35493 (N_35493,N_34625,N_34649);
xnor U35494 (N_35494,N_33819,N_34843);
nor U35495 (N_35495,N_32714,N_33715);
nand U35496 (N_35496,N_33623,N_33597);
nor U35497 (N_35497,N_34376,N_33617);
or U35498 (N_35498,N_33530,N_33570);
xor U35499 (N_35499,N_32649,N_34818);
xnor U35500 (N_35500,N_33823,N_32538);
xor U35501 (N_35501,N_34279,N_34857);
nor U35502 (N_35502,N_33185,N_33749);
or U35503 (N_35503,N_33310,N_32652);
nand U35504 (N_35504,N_34018,N_32895);
or U35505 (N_35505,N_33608,N_33159);
and U35506 (N_35506,N_32785,N_32796);
nand U35507 (N_35507,N_34391,N_32688);
or U35508 (N_35508,N_32757,N_33230);
and U35509 (N_35509,N_34509,N_33894);
or U35510 (N_35510,N_34210,N_33870);
nor U35511 (N_35511,N_34640,N_34246);
and U35512 (N_35512,N_34458,N_33324);
nor U35513 (N_35513,N_32815,N_32737);
or U35514 (N_35514,N_34399,N_33774);
nor U35515 (N_35515,N_32502,N_34603);
and U35516 (N_35516,N_33243,N_34528);
nand U35517 (N_35517,N_33552,N_33523);
xor U35518 (N_35518,N_33590,N_34389);
nor U35519 (N_35519,N_34397,N_33782);
and U35520 (N_35520,N_33858,N_33975);
nor U35521 (N_35521,N_33394,N_34383);
or U35522 (N_35522,N_32916,N_34477);
and U35523 (N_35523,N_34721,N_34681);
xor U35524 (N_35524,N_32675,N_33615);
nand U35525 (N_35525,N_32982,N_33415);
xnor U35526 (N_35526,N_34256,N_34968);
nor U35527 (N_35527,N_34966,N_34502);
nand U35528 (N_35528,N_34665,N_34334);
or U35529 (N_35529,N_34491,N_32619);
xnor U35530 (N_35530,N_34958,N_34108);
nor U35531 (N_35531,N_33661,N_33977);
or U35532 (N_35532,N_34511,N_33182);
and U35533 (N_35533,N_33117,N_33891);
or U35534 (N_35534,N_32571,N_34781);
xor U35535 (N_35535,N_32654,N_32776);
xnor U35536 (N_35536,N_34503,N_33694);
nand U35537 (N_35537,N_34364,N_34129);
nand U35538 (N_35538,N_33898,N_32965);
xor U35539 (N_35539,N_33944,N_32930);
and U35540 (N_35540,N_33034,N_33440);
xor U35541 (N_35541,N_33036,N_33853);
nand U35542 (N_35542,N_32613,N_34200);
and U35543 (N_35543,N_32630,N_34080);
xnor U35544 (N_35544,N_33276,N_34160);
and U35545 (N_35545,N_32637,N_34398);
xor U35546 (N_35546,N_33174,N_33322);
nor U35547 (N_35547,N_34651,N_33154);
nand U35548 (N_35548,N_33622,N_34436);
or U35549 (N_35549,N_34111,N_34732);
xor U35550 (N_35550,N_32650,N_34751);
and U35551 (N_35551,N_34715,N_34019);
and U35552 (N_35552,N_34368,N_33219);
nor U35553 (N_35553,N_34078,N_33830);
nor U35554 (N_35554,N_33152,N_34254);
or U35555 (N_35555,N_34716,N_33528);
or U35556 (N_35556,N_34194,N_34691);
nand U35557 (N_35557,N_34401,N_34641);
or U35558 (N_35558,N_33075,N_34463);
or U35559 (N_35559,N_33178,N_34432);
and U35560 (N_35560,N_32786,N_33286);
and U35561 (N_35561,N_33148,N_34325);
xor U35562 (N_35562,N_33274,N_34809);
and U35563 (N_35563,N_32555,N_32552);
nor U35564 (N_35564,N_33180,N_33225);
xnor U35565 (N_35565,N_34609,N_33968);
nor U35566 (N_35566,N_33058,N_34270);
or U35567 (N_35567,N_34260,N_33603);
xnor U35568 (N_35568,N_32781,N_32554);
nor U35569 (N_35569,N_33294,N_33425);
and U35570 (N_35570,N_33250,N_32933);
xnor U35571 (N_35571,N_34676,N_34199);
nor U35572 (N_35572,N_34960,N_34497);
nand U35573 (N_35573,N_34327,N_34316);
and U35574 (N_35574,N_34945,N_33861);
xnor U35575 (N_35575,N_33700,N_33418);
and U35576 (N_35576,N_34562,N_33660);
nor U35577 (N_35577,N_33840,N_34707);
or U35578 (N_35578,N_32928,N_32541);
nor U35579 (N_35579,N_32913,N_33091);
and U35580 (N_35580,N_32747,N_34608);
or U35581 (N_35581,N_34936,N_34212);
nor U35582 (N_35582,N_34349,N_32832);
nor U35583 (N_35583,N_33632,N_33844);
and U35584 (N_35584,N_34989,N_34171);
xnor U35585 (N_35585,N_34472,N_33191);
and U35586 (N_35586,N_32899,N_32876);
xnor U35587 (N_35587,N_34871,N_34309);
xnor U35588 (N_35588,N_34367,N_34693);
or U35589 (N_35589,N_34744,N_33115);
nor U35590 (N_35590,N_33761,N_32789);
xnor U35591 (N_35591,N_33606,N_32939);
xnor U35592 (N_35592,N_33503,N_32606);
nor U35593 (N_35593,N_33773,N_34620);
nand U35594 (N_35594,N_34273,N_33331);
xor U35595 (N_35595,N_33827,N_34059);
nor U35596 (N_35596,N_32535,N_33129);
nand U35597 (N_35597,N_33081,N_33011);
or U35598 (N_35598,N_33952,N_32615);
nand U35599 (N_35599,N_32946,N_34557);
and U35600 (N_35600,N_33486,N_33889);
or U35601 (N_35601,N_34795,N_34881);
nor U35602 (N_35602,N_34955,N_34733);
xnor U35603 (N_35603,N_32998,N_32964);
xnor U35604 (N_35604,N_33914,N_34815);
nor U35605 (N_35605,N_33659,N_32568);
nor U35606 (N_35606,N_34089,N_34816);
or U35607 (N_35607,N_34821,N_33334);
nor U35608 (N_35608,N_32604,N_34998);
or U35609 (N_35609,N_32676,N_32952);
nor U35610 (N_35610,N_33458,N_33101);
xor U35611 (N_35611,N_34582,N_34251);
or U35612 (N_35612,N_34759,N_33292);
and U35613 (N_35613,N_34173,N_33362);
xor U35614 (N_35614,N_33004,N_32950);
nand U35615 (N_35615,N_33263,N_33030);
or U35616 (N_35616,N_33481,N_32642);
nor U35617 (N_35617,N_34218,N_34225);
xnor U35618 (N_35618,N_33122,N_34140);
and U35619 (N_35619,N_34810,N_32847);
nand U35620 (N_35620,N_34238,N_32853);
nand U35621 (N_35621,N_34674,N_34688);
nor U35622 (N_35622,N_32609,N_33573);
nand U35623 (N_35623,N_32578,N_34205);
xor U35624 (N_35624,N_34563,N_32569);
nand U35625 (N_35625,N_34735,N_33614);
xor U35626 (N_35626,N_32990,N_33288);
xor U35627 (N_35627,N_33212,N_33538);
and U35628 (N_35628,N_33684,N_32842);
nand U35629 (N_35629,N_33701,N_34624);
nor U35630 (N_35630,N_33383,N_32721);
xor U35631 (N_35631,N_34567,N_33764);
xnor U35632 (N_35632,N_34149,N_33585);
and U35633 (N_35633,N_34544,N_32532);
xor U35634 (N_35634,N_32545,N_34947);
nor U35635 (N_35635,N_32953,N_33731);
or U35636 (N_35636,N_33014,N_34179);
or U35637 (N_35637,N_32556,N_33506);
nor U35638 (N_35638,N_34636,N_33231);
or U35639 (N_35639,N_34706,N_33007);
and U35640 (N_35640,N_32826,N_34993);
nand U35641 (N_35641,N_34537,N_32838);
nand U35642 (N_35642,N_33460,N_33512);
xnor U35643 (N_35643,N_34480,N_34856);
nand U35644 (N_35644,N_34192,N_34679);
or U35645 (N_35645,N_34393,N_34719);
or U35646 (N_35646,N_33931,N_32729);
or U35647 (N_35647,N_33596,N_34868);
and U35648 (N_35648,N_33327,N_33010);
nor U35649 (N_35649,N_33849,N_32618);
xnor U35650 (N_35650,N_33705,N_33340);
xor U35651 (N_35651,N_32778,N_32640);
nand U35652 (N_35652,N_33862,N_33238);
nand U35653 (N_35653,N_33042,N_34250);
nor U35654 (N_35654,N_33550,N_33085);
or U35655 (N_35655,N_33193,N_32963);
nand U35656 (N_35656,N_33546,N_33994);
xor U35657 (N_35657,N_33190,N_32526);
and U35658 (N_35658,N_33760,N_32882);
or U35659 (N_35659,N_34905,N_34365);
or U35660 (N_35660,N_34897,N_32748);
xor U35661 (N_35661,N_33662,N_34587);
xor U35662 (N_35662,N_33765,N_34110);
nor U35663 (N_35663,N_33063,N_34675);
xor U35664 (N_35664,N_33125,N_33845);
nor U35665 (N_35665,N_33936,N_33832);
nand U35666 (N_35666,N_32787,N_33921);
and U35667 (N_35667,N_33318,N_34010);
nand U35668 (N_35668,N_33326,N_33168);
nor U35669 (N_35669,N_34134,N_32780);
xnor U35670 (N_35670,N_33366,N_33031);
nand U35671 (N_35671,N_33244,N_33143);
nand U35672 (N_35672,N_32740,N_32700);
nand U35673 (N_35673,N_34081,N_32680);
xnor U35674 (N_35674,N_33097,N_32997);
xor U35675 (N_35675,N_33668,N_32884);
xor U35676 (N_35676,N_32914,N_33300);
nand U35677 (N_35677,N_34301,N_34645);
nand U35678 (N_35678,N_34382,N_34193);
xor U35679 (N_35679,N_34835,N_32725);
nor U35680 (N_35680,N_34441,N_34028);
or U35681 (N_35681,N_34774,N_33639);
and U35682 (N_35682,N_34017,N_34007);
nand U35683 (N_35683,N_33445,N_33910);
and U35684 (N_35684,N_33427,N_34289);
or U35685 (N_35685,N_33177,N_34446);
or U35686 (N_35686,N_33515,N_34813);
nand U35687 (N_35687,N_34886,N_32765);
xor U35688 (N_35688,N_33836,N_33653);
nand U35689 (N_35689,N_33025,N_34504);
xnor U35690 (N_35690,N_33304,N_33913);
and U35691 (N_35691,N_32660,N_33644);
xor U35692 (N_35692,N_34920,N_32967);
nor U35693 (N_35693,N_33257,N_32877);
or U35694 (N_35694,N_34542,N_33494);
or U35695 (N_35695,N_33786,N_34071);
nor U35696 (N_35696,N_33391,N_34416);
and U35697 (N_35697,N_32542,N_34158);
and U35698 (N_35698,N_32664,N_32992);
or U35699 (N_35699,N_32979,N_33685);
and U35700 (N_35700,N_33206,N_33966);
and U35701 (N_35701,N_34229,N_32790);
xor U35702 (N_35702,N_32839,N_33927);
or U35703 (N_35703,N_34161,N_33716);
nand U35704 (N_35704,N_34883,N_33838);
nor U35705 (N_35705,N_33500,N_33962);
nand U35706 (N_35706,N_32638,N_33435);
and U35707 (N_35707,N_32818,N_34767);
xor U35708 (N_35708,N_32724,N_34262);
and U35709 (N_35709,N_34417,N_34073);
and U35710 (N_35710,N_33598,N_32868);
nor U35711 (N_35711,N_32944,N_33045);
xor U35712 (N_35712,N_34671,N_34443);
nor U35713 (N_35713,N_33173,N_34757);
and U35714 (N_35714,N_33338,N_33803);
or U35715 (N_35715,N_34272,N_33771);
and U35716 (N_35716,N_33116,N_34323);
nor U35717 (N_35717,N_33625,N_33130);
and U35718 (N_35718,N_33795,N_34069);
nand U35719 (N_35719,N_34873,N_33469);
or U35720 (N_35720,N_32521,N_33364);
and U35721 (N_35721,N_34526,N_33258);
or U35722 (N_35722,N_33912,N_34775);
or U35723 (N_35723,N_33126,N_34155);
or U35724 (N_35724,N_34303,N_32927);
nor U35725 (N_35725,N_32575,N_33595);
and U35726 (N_35726,N_32567,N_34275);
nand U35727 (N_35727,N_34659,N_33713);
nand U35728 (N_35728,N_33902,N_34535);
or U35729 (N_35729,N_33750,N_33414);
xnor U35730 (N_35730,N_32861,N_33967);
or U35731 (N_35731,N_33671,N_33557);
nor U35732 (N_35732,N_32880,N_33536);
nor U35733 (N_35733,N_34890,N_33478);
nand U35734 (N_35734,N_32821,N_34203);
nand U35735 (N_35735,N_33825,N_34350);
xor U35736 (N_35736,N_34830,N_32811);
nand U35737 (N_35737,N_33848,N_34514);
nand U35738 (N_35738,N_33076,N_32834);
xor U35739 (N_35739,N_33175,N_34992);
xnor U35740 (N_35740,N_34475,N_32716);
nor U35741 (N_35741,N_34663,N_34999);
nor U35742 (N_35742,N_34079,N_34647);
or U35743 (N_35743,N_33266,N_34315);
or U35744 (N_35744,N_33843,N_34033);
or U35745 (N_35745,N_32989,N_34466);
and U35746 (N_35746,N_34870,N_32537);
nand U35747 (N_35747,N_34801,N_34973);
nand U35748 (N_35748,N_33078,N_34548);
xor U35749 (N_35749,N_33883,N_32621);
nor U35750 (N_35750,N_34154,N_33112);
nand U35751 (N_35751,N_34566,N_33470);
nand U35752 (N_35752,N_34473,N_32672);
or U35753 (N_35753,N_34141,N_32777);
xnor U35754 (N_35754,N_33410,N_34485);
and U35755 (N_35755,N_32693,N_33067);
nor U35756 (N_35756,N_32947,N_32823);
nand U35757 (N_35757,N_34516,N_32980);
nor U35758 (N_35758,N_33628,N_33735);
and U35759 (N_35759,N_32756,N_34406);
and U35760 (N_35760,N_34988,N_32910);
and U35761 (N_35761,N_32955,N_33144);
xnor U35762 (N_35762,N_32689,N_34766);
nand U35763 (N_35763,N_34579,N_32662);
and U35764 (N_35764,N_33522,N_32697);
nand U35765 (N_35765,N_34633,N_34036);
nor U35766 (N_35766,N_34344,N_34298);
nor U35767 (N_35767,N_34220,N_32889);
nand U35768 (N_35768,N_33909,N_32973);
nand U35769 (N_35769,N_34023,N_34755);
or U35770 (N_35770,N_34814,N_33817);
and U35771 (N_35771,N_33396,N_33996);
or U35772 (N_35772,N_33937,N_33389);
and U35773 (N_35773,N_33355,N_33140);
nor U35774 (N_35774,N_33673,N_33980);
and U35775 (N_35775,N_32976,N_32573);
and U35776 (N_35776,N_33424,N_34175);
xor U35777 (N_35777,N_34156,N_33714);
nand U35778 (N_35778,N_33938,N_32864);
nand U35779 (N_35779,N_34471,N_33105);
and U35780 (N_35780,N_34613,N_34660);
nand U35781 (N_35781,N_32524,N_34370);
and U35782 (N_35782,N_33228,N_34690);
nor U35783 (N_35783,N_32902,N_34152);
and U35784 (N_35784,N_33997,N_34063);
nand U35785 (N_35785,N_32925,N_33430);
and U35786 (N_35786,N_33686,N_33233);
xnor U35787 (N_35787,N_34317,N_34614);
and U35788 (N_35788,N_33961,N_33674);
nor U35789 (N_35789,N_32595,N_32679);
and U35790 (N_35790,N_34452,N_32752);
and U35791 (N_35791,N_33971,N_32941);
or U35792 (N_35792,N_34052,N_33411);
and U35793 (N_35793,N_34939,N_34483);
xor U35794 (N_35794,N_33899,N_32863);
and U35795 (N_35795,N_34554,N_34372);
or U35796 (N_35796,N_34068,N_33157);
nor U35797 (N_35797,N_34505,N_34709);
nor U35798 (N_35798,N_32893,N_34433);
nor U35799 (N_35799,N_34572,N_33815);
nand U35800 (N_35800,N_33188,N_33216);
xor U35801 (N_35801,N_33687,N_32942);
nand U35802 (N_35802,N_34930,N_32872);
nor U35803 (N_35803,N_33719,N_34571);
nor U35804 (N_35804,N_34366,N_33451);
and U35805 (N_35805,N_34407,N_33972);
or U35806 (N_35806,N_34605,N_33214);
xor U35807 (N_35807,N_34933,N_33647);
xor U35808 (N_35808,N_34064,N_34462);
or U35809 (N_35809,N_34853,N_34803);
nand U35810 (N_35810,N_34386,N_34615);
and U35811 (N_35811,N_33568,N_33346);
nand U35812 (N_35812,N_33436,N_32772);
nand U35813 (N_35813,N_33995,N_33426);
nor U35814 (N_35814,N_34244,N_34009);
nand U35815 (N_35815,N_32846,N_34799);
xnor U35816 (N_35816,N_34543,N_33920);
or U35817 (N_35817,N_32510,N_33405);
or U35818 (N_35818,N_33352,N_33776);
nand U35819 (N_35819,N_33107,N_33395);
nand U35820 (N_35820,N_33911,N_34119);
nor U35821 (N_35821,N_33382,N_34447);
nor U35822 (N_35822,N_33611,N_34345);
and U35823 (N_35823,N_33082,N_33950);
nor U35824 (N_35824,N_34806,N_34280);
and U35825 (N_35825,N_34976,N_32540);
nand U35826 (N_35826,N_34530,N_32608);
or U35827 (N_35827,N_32500,N_33806);
and U35828 (N_35828,N_33969,N_33232);
xor U35829 (N_35829,N_34148,N_32635);
xor U35830 (N_35830,N_33785,N_34750);
nand U35831 (N_35831,N_32957,N_32817);
nor U35832 (N_35832,N_32686,N_34661);
nand U35833 (N_35833,N_34261,N_34159);
and U35834 (N_35834,N_32530,N_34045);
xnor U35835 (N_35835,N_33583,N_34040);
or U35836 (N_35836,N_34038,N_34740);
and U35837 (N_35837,N_34310,N_34700);
nand U35838 (N_35838,N_34358,N_34589);
nor U35839 (N_35839,N_33008,N_33029);
or U35840 (N_35840,N_34523,N_32626);
and U35841 (N_35841,N_34247,N_34928);
xnor U35842 (N_35842,N_34336,N_33949);
nand U35843 (N_35843,N_34240,N_34451);
or U35844 (N_35844,N_32732,N_33724);
xor U35845 (N_35845,N_33472,N_33959);
and U35846 (N_35846,N_32958,N_32962);
and U35847 (N_35847,N_33466,N_33279);
xor U35848 (N_35848,N_34116,N_34035);
xor U35849 (N_35849,N_32782,N_34274);
and U35850 (N_35850,N_34100,N_32865);
and U35851 (N_35851,N_32996,N_33728);
and U35852 (N_35852,N_34726,N_33016);
nand U35853 (N_35853,N_34738,N_34314);
or U35854 (N_35854,N_34164,N_34685);
xor U35855 (N_35855,N_34823,N_33247);
and U35856 (N_35856,N_33438,N_33367);
nand U35857 (N_35857,N_33602,N_32843);
nand U35858 (N_35858,N_32945,N_33145);
xor U35859 (N_35859,N_34703,N_33299);
or U35860 (N_35860,N_34488,N_32890);
and U35861 (N_35861,N_33384,N_33664);
xnor U35862 (N_35862,N_33893,N_34969);
and U35863 (N_35863,N_33289,N_33824);
or U35864 (N_35864,N_32954,N_33095);
nand U35865 (N_35865,N_32710,N_33359);
nor U35866 (N_35866,N_33487,N_34980);
nand U35867 (N_35867,N_32970,N_34001);
nand U35868 (N_35868,N_33308,N_34560);
xnor U35869 (N_35869,N_34112,N_33133);
and U35870 (N_35870,N_34874,N_34876);
nor U35871 (N_35871,N_34974,N_32634);
or U35872 (N_35872,N_33723,N_32503);
nor U35873 (N_35873,N_32677,N_34320);
or U35874 (N_35874,N_34162,N_32583);
or U35875 (N_35875,N_34760,N_32892);
xor U35876 (N_35876,N_34305,N_33621);
and U35877 (N_35877,N_33207,N_33834);
xnor U35878 (N_35878,N_34644,N_32718);
nand U35879 (N_35879,N_34854,N_33073);
or U35880 (N_35880,N_33905,N_34979);
xnor U35881 (N_35881,N_32561,N_32758);
and U35882 (N_35882,N_34122,N_34747);
xnor U35883 (N_35883,N_34132,N_34748);
nand U35884 (N_35884,N_33651,N_33697);
and U35885 (N_35885,N_33319,N_33940);
nor U35886 (N_35886,N_34484,N_34982);
and U35887 (N_35887,N_32586,N_33691);
and U35888 (N_35888,N_32791,N_34182);
nor U35889 (N_35889,N_34500,N_33565);
or U35890 (N_35890,N_32529,N_34490);
nor U35891 (N_35891,N_33273,N_34239);
nand U35892 (N_35892,N_34510,N_33009);
nand U35893 (N_35893,N_34232,N_32907);
or U35894 (N_35894,N_34055,N_33189);
xnor U35895 (N_35895,N_32643,N_34950);
xor U35896 (N_35896,N_34029,N_32582);
and U35897 (N_35897,N_33779,N_33526);
and U35898 (N_35898,N_34418,N_34359);
xor U35899 (N_35899,N_33162,N_33680);
or U35900 (N_35900,N_32515,N_34506);
xnor U35901 (N_35901,N_33312,N_34329);
nor U35902 (N_35902,N_33591,N_34828);
xnor U35903 (N_35903,N_33072,N_32706);
nor U35904 (N_35904,N_33006,N_32610);
and U35905 (N_35905,N_34429,N_34292);
or U35906 (N_35906,N_33712,N_32988);
xnor U35907 (N_35907,N_34172,N_33298);
and U35908 (N_35908,N_32698,N_34304);
and U35909 (N_35909,N_34259,N_32655);
xor U35910 (N_35910,N_34866,N_33730);
or U35911 (N_35911,N_33514,N_34904);
and U35912 (N_35912,N_33262,N_34825);
and U35913 (N_35913,N_33548,N_32551);
and U35914 (N_35914,N_34354,N_32938);
and U35915 (N_35915,N_33499,N_33933);
or U35916 (N_35916,N_34460,N_33672);
nor U35917 (N_35917,N_34595,N_33561);
nand U35918 (N_35918,N_34638,N_34769);
and U35919 (N_35919,N_33305,N_32670);
xnor U35920 (N_35920,N_32797,N_33313);
nand U35921 (N_35921,N_33109,N_34369);
xor U35922 (N_35922,N_32559,N_33069);
nor U35923 (N_35923,N_34474,N_33901);
nand U35924 (N_35924,N_33222,N_34728);
and U35925 (N_35925,N_32743,N_34470);
or U35926 (N_35926,N_34054,N_34032);
and U35927 (N_35927,N_34486,N_33993);
or U35928 (N_35928,N_33120,N_34967);
nand U35929 (N_35929,N_34896,N_34234);
nand U35930 (N_35930,N_32576,N_32779);
xnor U35931 (N_35931,N_32522,N_34573);
nor U35932 (N_35932,N_34233,N_33521);
or U35933 (N_35933,N_33866,N_33992);
nand U35934 (N_35934,N_32667,N_32993);
nand U35935 (N_35935,N_33609,N_33492);
or U35936 (N_35936,N_33600,N_34787);
nand U35937 (N_35937,N_33878,N_33851);
or U35938 (N_35938,N_32600,N_34822);
xnor U35939 (N_35939,N_34902,N_34887);
and U35940 (N_35940,N_32624,N_33135);
nor U35941 (N_35941,N_34637,N_33493);
or U35942 (N_35942,N_34213,N_33442);
or U35943 (N_35943,N_32631,N_33654);
and U35944 (N_35944,N_33929,N_33897);
nor U35945 (N_35945,N_34459,N_33675);
or U35946 (N_35946,N_32605,N_33928);
xnor U35947 (N_35947,N_34932,N_33211);
or U35948 (N_35948,N_33345,N_34056);
nor U35949 (N_35949,N_33640,N_34564);
nor U35950 (N_35950,N_34629,N_34893);
or U35951 (N_35951,N_32585,N_34739);
and U35952 (N_35952,N_32897,N_34427);
xnor U35953 (N_35953,N_32717,N_33919);
xor U35954 (N_35954,N_33679,N_32983);
xnor U35955 (N_35955,N_34130,N_33433);
and U35956 (N_35956,N_32951,N_34911);
or U35957 (N_35957,N_33163,N_34057);
or U35958 (N_35958,N_34031,N_33678);
nor U35959 (N_35959,N_33024,N_34865);
xor U35960 (N_35960,N_34997,N_33229);
xor U35961 (N_35961,N_34915,N_32633);
or U35962 (N_35962,N_33223,N_33220);
xnor U35963 (N_35963,N_34898,N_33437);
nor U35964 (N_35964,N_33423,N_34522);
nor U35965 (N_35965,N_33916,N_34360);
or U35966 (N_35966,N_32788,N_32924);
nor U35967 (N_35967,N_33670,N_34330);
and U35968 (N_35968,N_34337,N_33275);
nand U35969 (N_35969,N_34699,N_33164);
nor U35970 (N_35970,N_34880,N_33253);
nand U35971 (N_35971,N_34127,N_32705);
xnor U35972 (N_35972,N_33789,N_34489);
nand U35973 (N_35973,N_33635,N_33141);
and U35974 (N_35974,N_33147,N_34221);
nor U35975 (N_35975,N_33655,N_32870);
or U35976 (N_35976,N_33934,N_34253);
nor U35977 (N_35977,N_33221,N_33788);
or U35978 (N_35978,N_32701,N_32574);
and U35979 (N_35979,N_34257,N_32562);
nand U35980 (N_35980,N_33209,N_34695);
or U35981 (N_35981,N_32692,N_33576);
nor U35982 (N_35982,N_32828,N_34066);
and U35983 (N_35983,N_33560,N_34067);
nand U35984 (N_35984,N_32859,N_32974);
xor U35985 (N_35985,N_34216,N_33291);
or U35986 (N_35986,N_33021,N_33852);
nand U35987 (N_35987,N_34340,N_33387);
or U35988 (N_35988,N_33106,N_32738);
xnor U35989 (N_35989,N_32570,N_34378);
and U35990 (N_35990,N_34302,N_34373);
nand U35991 (N_35991,N_34652,N_33863);
or U35992 (N_35992,N_34839,N_34476);
nand U35993 (N_35993,N_34927,N_32800);
and U35994 (N_35994,N_34798,N_33408);
nor U35995 (N_35995,N_32720,N_33876);
and U35996 (N_35996,N_33540,N_34684);
nand U35997 (N_35997,N_33210,N_33529);
xor U35998 (N_35998,N_32639,N_34042);
nand U35999 (N_35999,N_34678,N_34332);
and U36000 (N_36000,N_34727,N_34584);
or U36001 (N_36001,N_34581,N_34237);
and U36002 (N_36002,N_33103,N_32517);
or U36003 (N_36003,N_34805,N_33132);
and U36004 (N_36004,N_32830,N_34616);
or U36005 (N_36005,N_34005,N_33783);
xnor U36006 (N_36006,N_33293,N_33558);
nand U36007 (N_36007,N_34099,N_34243);
or U36008 (N_36008,N_33958,N_33397);
nand U36009 (N_36009,N_33489,N_33924);
or U36010 (N_36010,N_34324,N_32707);
or U36011 (N_36011,N_33948,N_34278);
and U36012 (N_36012,N_33989,N_33360);
nand U36013 (N_36013,N_33467,N_34702);
xnor U36014 (N_36014,N_32565,N_33601);
nor U36015 (N_36015,N_33943,N_34840);
xnor U36016 (N_36016,N_33392,N_34098);
or U36017 (N_36017,N_33696,N_33707);
and U36018 (N_36018,N_33918,N_33272);
nor U36019 (N_36019,N_34722,N_33380);
xnor U36020 (N_36020,N_34972,N_34714);
xor U36021 (N_36021,N_34934,N_33811);
and U36022 (N_36022,N_33892,N_32764);
and U36023 (N_36023,N_33449,N_33688);
xor U36024 (N_36024,N_34990,N_33875);
nor U36025 (N_36025,N_33149,N_32607);
xor U36026 (N_36026,N_32912,N_34439);
xor U36027 (N_36027,N_33698,N_33496);
nor U36028 (N_36028,N_33999,N_32887);
and U36029 (N_36029,N_33428,N_34770);
nor U36030 (N_36030,N_34780,N_34600);
nand U36031 (N_36031,N_34412,N_34588);
nand U36032 (N_36032,N_34478,N_33706);
nand U36033 (N_36033,N_34949,N_34348);
nand U36034 (N_36034,N_32599,N_33497);
nor U36035 (N_36035,N_33658,N_33198);
xor U36036 (N_36036,N_34186,N_34265);
or U36037 (N_36037,N_34167,N_33104);
nor U36038 (N_36038,N_33051,N_34082);
nand U36039 (N_36039,N_32508,N_34894);
nor U36040 (N_36040,N_34938,N_34628);
nor U36041 (N_36041,N_33343,N_34956);
nand U36042 (N_36042,N_34601,N_32883);
xnor U36043 (N_36043,N_33356,N_32534);
nand U36044 (N_36044,N_34105,N_34858);
xor U36045 (N_36045,N_33032,N_34855);
nand U36046 (N_36046,N_34453,N_32917);
nand U36047 (N_36047,N_34991,N_33053);
nor U36048 (N_36048,N_34779,N_33880);
and U36049 (N_36049,N_32622,N_34255);
nand U36050 (N_36050,N_32553,N_33939);
nand U36051 (N_36051,N_34090,N_32873);
nand U36052 (N_36052,N_34762,N_34291);
and U36053 (N_36053,N_33342,N_33404);
and U36054 (N_36054,N_33498,N_33096);
nand U36055 (N_36055,N_33734,N_32819);
xnor U36056 (N_36056,N_33915,N_33699);
nor U36057 (N_36057,N_33301,N_34381);
and U36058 (N_36058,N_34892,N_34187);
or U36059 (N_36059,N_32881,N_33358);
and U36060 (N_36060,N_34043,N_34487);
nand U36061 (N_36061,N_34734,N_33516);
nor U36062 (N_36062,N_34191,N_33446);
or U36063 (N_36063,N_33399,N_34258);
or U36064 (N_36064,N_32767,N_34481);
nand U36065 (N_36065,N_34086,N_34448);
nor U36066 (N_36066,N_34541,N_34899);
nor U36067 (N_36067,N_34852,N_33167);
nor U36068 (N_36068,N_34804,N_34545);
nand U36069 (N_36069,N_34139,N_32731);
xor U36070 (N_36070,N_33039,N_33641);
or U36071 (N_36071,N_32981,N_32805);
xnor U36072 (N_36072,N_34206,N_33507);
nand U36073 (N_36073,N_32509,N_34422);
xor U36074 (N_36074,N_33930,N_33323);
and U36075 (N_36075,N_34784,N_33059);
nor U36076 (N_36076,N_33759,N_34517);
and U36077 (N_36077,N_34170,N_32766);
nand U36078 (N_36078,N_34921,N_33772);
nor U36079 (N_36079,N_34051,N_33369);
xor U36080 (N_36080,N_34926,N_32769);
or U36081 (N_36081,N_34531,N_34672);
nor U36082 (N_36082,N_33184,N_32728);
xnor U36083 (N_36083,N_34680,N_34444);
nor U36084 (N_36084,N_34598,N_34321);
nand U36085 (N_36085,N_33200,N_32921);
and U36086 (N_36086,N_33330,N_32627);
or U36087 (N_36087,N_33461,N_33365);
and U36088 (N_36088,N_33321,N_34845);
nor U36089 (N_36089,N_34985,N_33998);
and U36090 (N_36090,N_33044,N_34978);
nor U36091 (N_36091,N_32674,N_32625);
nand U36092 (N_36092,N_34807,N_33179);
nor U36093 (N_36093,N_33956,N_34602);
and U36094 (N_36094,N_34888,N_32629);
nor U36095 (N_36095,N_34021,N_33978);
nand U36096 (N_36096,N_34008,N_33484);
or U36097 (N_36097,N_33246,N_34027);
nand U36098 (N_36098,N_34599,N_33703);
xor U36099 (N_36099,N_34030,N_34977);
or U36100 (N_36100,N_34197,N_34908);
nand U36101 (N_36101,N_34128,N_34981);
and U36102 (N_36102,N_33513,N_33187);
or U36103 (N_36103,N_33050,N_33973);
or U36104 (N_36104,N_33974,N_34115);
and U36105 (N_36105,N_34313,N_34053);
nor U36106 (N_36106,N_33629,N_34879);
and U36107 (N_36107,N_34041,N_33281);
nor U36108 (N_36108,N_34846,N_34084);
nand U36109 (N_36109,N_33170,N_34319);
xor U36110 (N_36110,N_33000,N_34711);
nand U36111 (N_36111,N_34145,N_33416);
xnor U36112 (N_36112,N_32598,N_33619);
or U36113 (N_36113,N_33001,N_33256);
or U36114 (N_36114,N_33264,N_34222);
nor U36115 (N_36115,N_34753,N_32856);
or U36116 (N_36116,N_32948,N_33235);
or U36117 (N_36117,N_33241,N_32753);
nand U36118 (N_36118,N_34061,N_33777);
and U36119 (N_36119,N_33074,N_32636);
nand U36120 (N_36120,N_32813,N_34611);
xor U36121 (N_36121,N_32577,N_32591);
or U36122 (N_36122,N_34547,N_34591);
nand U36123 (N_36123,N_33741,N_33681);
nor U36124 (N_36124,N_33350,N_32539);
nand U36125 (N_36125,N_32829,N_34034);
nand U36126 (N_36126,N_32566,N_33240);
xnor U36127 (N_36127,N_33791,N_33386);
nor U36128 (N_36128,N_33265,N_34667);
nor U36129 (N_36129,N_34912,N_34761);
nand U36130 (N_36130,N_33652,N_33669);
nand U36131 (N_36131,N_33491,N_32531);
or U36132 (N_36132,N_34281,N_34597);
and U36133 (N_36133,N_34202,N_33637);
and U36134 (N_36134,N_33748,N_34646);
nor U36135 (N_36135,N_34501,N_34226);
nor U36136 (N_36136,N_33054,N_34431);
xor U36137 (N_36137,N_34267,N_32691);
xnor U36138 (N_36138,N_34970,N_32653);
nor U36139 (N_36139,N_33348,N_33224);
and U36140 (N_36140,N_33831,N_34445);
xnor U36141 (N_36141,N_33136,N_33361);
or U36142 (N_36142,N_34653,N_33080);
and U36143 (N_36143,N_33589,N_34143);
nand U36144 (N_36144,N_33520,N_33624);
nand U36145 (N_36145,N_33336,N_33864);
nand U36146 (N_36146,N_32723,N_34996);
or U36147 (N_36147,N_34763,N_33534);
nor U36148 (N_36148,N_34786,N_33277);
and U36149 (N_36149,N_34114,N_33778);
xnor U36150 (N_36150,N_34103,N_34796);
nand U36151 (N_36151,N_33666,N_33158);
nor U36152 (N_36152,N_34347,N_34394);
and U36153 (N_36153,N_33579,N_33099);
or U36154 (N_36154,N_34909,N_32835);
and U36155 (N_36155,N_34948,N_32694);
and U36156 (N_36156,N_33710,N_32520);
xnor U36157 (N_36157,N_34861,N_34408);
xor U36158 (N_36158,N_34076,N_33854);
nor U36159 (N_36159,N_34831,N_34687);
nand U36160 (N_36160,N_33525,N_33495);
nand U36161 (N_36161,N_32727,N_32793);
xnor U36162 (N_36162,N_32603,N_33353);
nand U36163 (N_36163,N_32712,N_34539);
nand U36164 (N_36164,N_32589,N_32937);
nand U36165 (N_36165,N_33113,N_34294);
xnor U36166 (N_36166,N_32761,N_33569);
and U36167 (N_36167,N_33260,N_33925);
xnor U36168 (N_36168,N_34768,N_33631);
and U36169 (N_36169,N_33226,N_33732);
and U36170 (N_36170,N_34121,N_34520);
or U36171 (N_36171,N_33667,N_33895);
and U36172 (N_36172,N_32926,N_32774);
nand U36173 (N_36173,N_33800,N_34198);
and U36174 (N_36174,N_33626,N_33102);
nand U36175 (N_36175,N_34188,N_33871);
and U36176 (N_36176,N_34983,N_34196);
and U36177 (N_36177,N_34697,N_34123);
nor U36178 (N_36178,N_34913,N_34964);
xnor U36179 (N_36179,N_33432,N_33098);
or U36180 (N_36180,N_33068,N_34374);
xnor U36181 (N_36181,N_34895,N_33049);
nand U36182 (N_36182,N_33571,N_33986);
or U36183 (N_36183,N_34963,N_33377);
or U36184 (N_36184,N_32696,N_33026);
nand U36185 (N_36185,N_33856,N_34618);
xor U36186 (N_36186,N_32734,N_32617);
xnor U36187 (N_36187,N_32602,N_33964);
nand U36188 (N_36188,N_32523,N_32678);
nand U36189 (N_36189,N_33869,N_33572);
nand U36190 (N_36190,N_32854,N_34540);
and U36191 (N_36191,N_33035,N_32875);
nor U36192 (N_36192,N_34789,N_33269);
xor U36193 (N_36193,N_33763,N_32931);
nor U36194 (N_36194,N_33979,N_34297);
xor U36195 (N_36195,N_34515,N_34594);
and U36196 (N_36196,N_32922,N_33194);
xnor U36197 (N_36197,N_33071,N_34185);
xor U36198 (N_36198,N_34454,N_32506);
nor U36199 (N_36199,N_33642,N_34046);
xor U36200 (N_36200,N_34811,N_34670);
or U36201 (N_36201,N_32932,N_34026);
nand U36202 (N_36202,N_34209,N_34231);
and U36203 (N_36203,N_33138,N_34512);
nor U36204 (N_36204,N_33768,N_32814);
nand U36205 (N_36205,N_33479,N_32645);
and U36206 (N_36206,N_34724,N_33501);
and U36207 (N_36207,N_33510,N_34794);
nor U36208 (N_36208,N_33242,N_34995);
xor U36209 (N_36209,N_34729,N_32699);
and U36210 (N_36210,N_33023,N_34153);
nor U36211 (N_36211,N_33769,N_33475);
or U36212 (N_36212,N_33407,N_34538);
nor U36213 (N_36213,N_34091,N_34630);
and U36214 (N_36214,N_34457,N_33088);
nand U36215 (N_36215,N_33215,N_34461);
xnor U36216 (N_36216,N_34166,N_34705);
xor U36217 (N_36217,N_33627,N_32920);
xnor U36218 (N_36218,N_34215,N_33118);
nor U36219 (N_36219,N_33213,N_33476);
nand U36220 (N_36220,N_33828,N_33535);
nor U36221 (N_36221,N_33955,N_34464);
xnor U36222 (N_36222,N_34717,N_32588);
and U36223 (N_36223,N_33268,N_34006);
xnor U36224 (N_36224,N_33729,N_34228);
or U36225 (N_36225,N_34306,N_32896);
xnor U36226 (N_36226,N_32661,N_32905);
nor U36227 (N_36227,N_34252,N_33311);
nor U36228 (N_36228,N_33683,N_33043);
nand U36229 (N_36229,N_33781,N_34282);
and U36230 (N_36230,N_34507,N_32739);
xnor U36231 (N_36231,N_33718,N_32879);
xor U36232 (N_36232,N_32597,N_32906);
xnor U36233 (N_36233,N_33578,N_34817);
nand U36234 (N_36234,N_34617,N_34585);
xnor U36235 (N_36235,N_33648,N_34788);
nand U36236 (N_36236,N_33248,N_33317);
and U36237 (N_36237,N_33290,N_34060);
nor U36238 (N_36238,N_34736,N_32762);
or U36239 (N_36239,N_33171,N_33634);
xnor U36240 (N_36240,N_34104,N_34627);
nor U36241 (N_36241,N_33877,N_33766);
or U36242 (N_36242,N_33390,N_34189);
or U36243 (N_36243,N_34219,N_34424);
or U36244 (N_36244,N_34479,N_34847);
nand U36245 (N_36245,N_32746,N_33960);
nor U36246 (N_36246,N_33463,N_33131);
nand U36247 (N_36247,N_32768,N_34495);
nor U36248 (N_36248,N_34725,N_33970);
nand U36249 (N_36249,N_32934,N_33166);
xnor U36250 (N_36250,N_32704,N_32746);
nor U36251 (N_36251,N_33044,N_34082);
nor U36252 (N_36252,N_32966,N_32635);
or U36253 (N_36253,N_33516,N_34470);
or U36254 (N_36254,N_33792,N_33218);
and U36255 (N_36255,N_33313,N_34424);
nor U36256 (N_36256,N_34186,N_34884);
nand U36257 (N_36257,N_33708,N_33096);
xnor U36258 (N_36258,N_33499,N_32674);
nand U36259 (N_36259,N_34879,N_32970);
or U36260 (N_36260,N_33050,N_33832);
nor U36261 (N_36261,N_33766,N_33922);
and U36262 (N_36262,N_34707,N_32809);
xnor U36263 (N_36263,N_32678,N_34783);
nor U36264 (N_36264,N_33155,N_34244);
and U36265 (N_36265,N_34296,N_32940);
xnor U36266 (N_36266,N_32708,N_34647);
nand U36267 (N_36267,N_33266,N_33983);
xnor U36268 (N_36268,N_33523,N_32919);
and U36269 (N_36269,N_34775,N_34701);
nand U36270 (N_36270,N_32934,N_33351);
and U36271 (N_36271,N_33505,N_33071);
and U36272 (N_36272,N_34772,N_34832);
and U36273 (N_36273,N_34410,N_34604);
nand U36274 (N_36274,N_33025,N_33063);
xnor U36275 (N_36275,N_34369,N_32668);
or U36276 (N_36276,N_32749,N_34721);
nor U36277 (N_36277,N_32686,N_33781);
nor U36278 (N_36278,N_32626,N_32911);
and U36279 (N_36279,N_34623,N_32761);
and U36280 (N_36280,N_33917,N_34940);
nor U36281 (N_36281,N_32907,N_34670);
nor U36282 (N_36282,N_34450,N_32599);
nor U36283 (N_36283,N_32740,N_33635);
nand U36284 (N_36284,N_34019,N_34630);
nand U36285 (N_36285,N_34212,N_34708);
xor U36286 (N_36286,N_33933,N_33676);
and U36287 (N_36287,N_34645,N_33760);
xnor U36288 (N_36288,N_33075,N_32617);
nor U36289 (N_36289,N_33871,N_32780);
or U36290 (N_36290,N_33897,N_34329);
nand U36291 (N_36291,N_33112,N_34171);
nand U36292 (N_36292,N_33197,N_33931);
xnor U36293 (N_36293,N_33363,N_34308);
or U36294 (N_36294,N_34601,N_33120);
and U36295 (N_36295,N_34826,N_34042);
nand U36296 (N_36296,N_33297,N_33213);
xor U36297 (N_36297,N_34845,N_34310);
xor U36298 (N_36298,N_32704,N_34021);
xor U36299 (N_36299,N_33167,N_32838);
and U36300 (N_36300,N_34719,N_32668);
or U36301 (N_36301,N_33970,N_34142);
nand U36302 (N_36302,N_34438,N_33046);
or U36303 (N_36303,N_32861,N_33134);
nand U36304 (N_36304,N_34908,N_34837);
nand U36305 (N_36305,N_33684,N_33851);
and U36306 (N_36306,N_33208,N_33915);
nand U36307 (N_36307,N_32509,N_34953);
nor U36308 (N_36308,N_34471,N_34925);
or U36309 (N_36309,N_32741,N_32852);
nand U36310 (N_36310,N_32544,N_34825);
and U36311 (N_36311,N_32612,N_32656);
nand U36312 (N_36312,N_34999,N_34640);
nor U36313 (N_36313,N_34291,N_33346);
nand U36314 (N_36314,N_34868,N_34813);
and U36315 (N_36315,N_34739,N_34936);
xnor U36316 (N_36316,N_33994,N_34405);
or U36317 (N_36317,N_34056,N_32772);
nand U36318 (N_36318,N_32809,N_32754);
and U36319 (N_36319,N_34984,N_34645);
nand U36320 (N_36320,N_33821,N_32912);
nor U36321 (N_36321,N_32627,N_34888);
or U36322 (N_36322,N_33841,N_33515);
nand U36323 (N_36323,N_34503,N_32585);
and U36324 (N_36324,N_33596,N_34159);
nand U36325 (N_36325,N_34008,N_34531);
or U36326 (N_36326,N_32727,N_32893);
nand U36327 (N_36327,N_33900,N_34858);
xnor U36328 (N_36328,N_33512,N_34873);
nor U36329 (N_36329,N_34196,N_34074);
nand U36330 (N_36330,N_33524,N_33651);
and U36331 (N_36331,N_34237,N_34569);
or U36332 (N_36332,N_33644,N_34853);
xnor U36333 (N_36333,N_33627,N_33650);
or U36334 (N_36334,N_33355,N_33044);
and U36335 (N_36335,N_34543,N_32714);
nor U36336 (N_36336,N_33967,N_33340);
or U36337 (N_36337,N_34429,N_33301);
or U36338 (N_36338,N_34842,N_34120);
nand U36339 (N_36339,N_32946,N_33521);
nand U36340 (N_36340,N_34200,N_32630);
nand U36341 (N_36341,N_33554,N_33393);
or U36342 (N_36342,N_33441,N_33129);
and U36343 (N_36343,N_33444,N_33681);
xor U36344 (N_36344,N_32857,N_34004);
or U36345 (N_36345,N_33690,N_34264);
or U36346 (N_36346,N_33187,N_33782);
and U36347 (N_36347,N_33474,N_33116);
xor U36348 (N_36348,N_34382,N_33870);
nand U36349 (N_36349,N_33590,N_33711);
nand U36350 (N_36350,N_34033,N_34745);
xor U36351 (N_36351,N_32895,N_34554);
and U36352 (N_36352,N_34930,N_34305);
nor U36353 (N_36353,N_34594,N_33171);
and U36354 (N_36354,N_34096,N_34454);
nand U36355 (N_36355,N_34604,N_33060);
and U36356 (N_36356,N_33595,N_33628);
nor U36357 (N_36357,N_34790,N_34569);
nor U36358 (N_36358,N_33214,N_33452);
and U36359 (N_36359,N_33757,N_33709);
nor U36360 (N_36360,N_34111,N_32747);
or U36361 (N_36361,N_33816,N_33746);
xor U36362 (N_36362,N_32706,N_33202);
xnor U36363 (N_36363,N_33592,N_32585);
nand U36364 (N_36364,N_32522,N_34290);
and U36365 (N_36365,N_33396,N_34290);
or U36366 (N_36366,N_33590,N_33596);
nor U36367 (N_36367,N_34330,N_34389);
nor U36368 (N_36368,N_34422,N_34694);
nor U36369 (N_36369,N_32910,N_34049);
and U36370 (N_36370,N_32541,N_33500);
or U36371 (N_36371,N_32915,N_32777);
xor U36372 (N_36372,N_32761,N_32675);
nor U36373 (N_36373,N_33228,N_34132);
and U36374 (N_36374,N_34350,N_32798);
xnor U36375 (N_36375,N_34943,N_34883);
or U36376 (N_36376,N_33443,N_34517);
xnor U36377 (N_36377,N_33138,N_33405);
nor U36378 (N_36378,N_34816,N_33182);
xor U36379 (N_36379,N_33565,N_32954);
nor U36380 (N_36380,N_33940,N_33866);
xnor U36381 (N_36381,N_33080,N_34607);
nand U36382 (N_36382,N_33356,N_33049);
nor U36383 (N_36383,N_34422,N_33295);
xnor U36384 (N_36384,N_34433,N_33436);
xnor U36385 (N_36385,N_34736,N_34439);
or U36386 (N_36386,N_34391,N_32623);
or U36387 (N_36387,N_33364,N_34712);
xnor U36388 (N_36388,N_33312,N_33115);
nand U36389 (N_36389,N_34307,N_34699);
nand U36390 (N_36390,N_32562,N_33033);
nand U36391 (N_36391,N_33178,N_33692);
nand U36392 (N_36392,N_33071,N_34806);
xor U36393 (N_36393,N_33478,N_32926);
nor U36394 (N_36394,N_34844,N_33000);
nor U36395 (N_36395,N_32632,N_34449);
or U36396 (N_36396,N_33187,N_33330);
and U36397 (N_36397,N_33487,N_33576);
and U36398 (N_36398,N_33093,N_32749);
xor U36399 (N_36399,N_33153,N_32913);
nor U36400 (N_36400,N_32786,N_34084);
nand U36401 (N_36401,N_33304,N_33219);
nor U36402 (N_36402,N_32676,N_33124);
nand U36403 (N_36403,N_34512,N_33960);
and U36404 (N_36404,N_33086,N_34124);
and U36405 (N_36405,N_32923,N_33901);
and U36406 (N_36406,N_34067,N_34727);
nor U36407 (N_36407,N_32652,N_32890);
nor U36408 (N_36408,N_33328,N_33256);
nand U36409 (N_36409,N_33259,N_34535);
xnor U36410 (N_36410,N_33461,N_34480);
xor U36411 (N_36411,N_34938,N_33530);
xor U36412 (N_36412,N_32510,N_32790);
nor U36413 (N_36413,N_32683,N_33126);
and U36414 (N_36414,N_33369,N_33997);
nor U36415 (N_36415,N_33526,N_34873);
xor U36416 (N_36416,N_32661,N_33501);
nor U36417 (N_36417,N_32592,N_33511);
nor U36418 (N_36418,N_34784,N_32500);
and U36419 (N_36419,N_34583,N_32988);
nand U36420 (N_36420,N_34879,N_34680);
nor U36421 (N_36421,N_33378,N_33863);
or U36422 (N_36422,N_32579,N_34160);
nor U36423 (N_36423,N_33338,N_34161);
nor U36424 (N_36424,N_32639,N_34624);
nand U36425 (N_36425,N_34147,N_33926);
nor U36426 (N_36426,N_34939,N_34550);
nor U36427 (N_36427,N_34633,N_33081);
nand U36428 (N_36428,N_34477,N_33480);
and U36429 (N_36429,N_33651,N_34979);
and U36430 (N_36430,N_34756,N_34134);
or U36431 (N_36431,N_34667,N_33736);
xor U36432 (N_36432,N_33534,N_33821);
nor U36433 (N_36433,N_33382,N_34210);
nor U36434 (N_36434,N_33306,N_33105);
nand U36435 (N_36435,N_32659,N_33784);
and U36436 (N_36436,N_32917,N_32883);
nor U36437 (N_36437,N_32976,N_33265);
or U36438 (N_36438,N_34198,N_33901);
and U36439 (N_36439,N_32624,N_32874);
nand U36440 (N_36440,N_33509,N_32855);
nand U36441 (N_36441,N_32996,N_33137);
xnor U36442 (N_36442,N_33675,N_32625);
and U36443 (N_36443,N_33374,N_33184);
or U36444 (N_36444,N_32569,N_33711);
nor U36445 (N_36445,N_34591,N_33664);
nand U36446 (N_36446,N_34631,N_32765);
nor U36447 (N_36447,N_33716,N_33744);
nor U36448 (N_36448,N_32939,N_33203);
and U36449 (N_36449,N_33063,N_34826);
or U36450 (N_36450,N_32664,N_32634);
or U36451 (N_36451,N_33925,N_34749);
and U36452 (N_36452,N_34444,N_34405);
nand U36453 (N_36453,N_34857,N_33911);
or U36454 (N_36454,N_32788,N_33741);
xor U36455 (N_36455,N_33083,N_32755);
xor U36456 (N_36456,N_32682,N_34188);
nor U36457 (N_36457,N_34344,N_32557);
or U36458 (N_36458,N_32736,N_33139);
nor U36459 (N_36459,N_33542,N_32925);
and U36460 (N_36460,N_34497,N_34736);
nand U36461 (N_36461,N_34850,N_34821);
nor U36462 (N_36462,N_33372,N_32921);
and U36463 (N_36463,N_33302,N_34688);
and U36464 (N_36464,N_34753,N_34212);
and U36465 (N_36465,N_33877,N_34860);
nand U36466 (N_36466,N_34879,N_33037);
and U36467 (N_36467,N_34767,N_33870);
nor U36468 (N_36468,N_34297,N_34562);
or U36469 (N_36469,N_33264,N_32521);
and U36470 (N_36470,N_33906,N_34228);
nand U36471 (N_36471,N_33047,N_33410);
nand U36472 (N_36472,N_34777,N_33087);
or U36473 (N_36473,N_32751,N_32707);
nor U36474 (N_36474,N_34392,N_33715);
or U36475 (N_36475,N_33279,N_32654);
or U36476 (N_36476,N_33183,N_34610);
nand U36477 (N_36477,N_33575,N_33128);
or U36478 (N_36478,N_33090,N_33099);
and U36479 (N_36479,N_32968,N_33060);
nand U36480 (N_36480,N_33051,N_33337);
nor U36481 (N_36481,N_33423,N_33794);
xor U36482 (N_36482,N_33589,N_34678);
xor U36483 (N_36483,N_32736,N_33902);
and U36484 (N_36484,N_33553,N_34300);
or U36485 (N_36485,N_32794,N_32744);
and U36486 (N_36486,N_32695,N_34482);
nor U36487 (N_36487,N_33297,N_33692);
xnor U36488 (N_36488,N_32502,N_34912);
and U36489 (N_36489,N_33596,N_34292);
xor U36490 (N_36490,N_33394,N_33843);
or U36491 (N_36491,N_32593,N_34369);
nor U36492 (N_36492,N_34325,N_33428);
and U36493 (N_36493,N_34753,N_33041);
and U36494 (N_36494,N_34864,N_34134);
nand U36495 (N_36495,N_33017,N_32728);
nor U36496 (N_36496,N_33582,N_33857);
nor U36497 (N_36497,N_34353,N_32915);
nor U36498 (N_36498,N_33766,N_33204);
and U36499 (N_36499,N_33149,N_34564);
nor U36500 (N_36500,N_32781,N_32697);
nand U36501 (N_36501,N_34078,N_34537);
or U36502 (N_36502,N_33459,N_32505);
or U36503 (N_36503,N_33731,N_33949);
nand U36504 (N_36504,N_32626,N_34067);
xor U36505 (N_36505,N_33423,N_33718);
nor U36506 (N_36506,N_32963,N_33937);
xnor U36507 (N_36507,N_33720,N_32664);
nor U36508 (N_36508,N_32534,N_33673);
nor U36509 (N_36509,N_34739,N_34974);
and U36510 (N_36510,N_32639,N_33416);
xnor U36511 (N_36511,N_34035,N_33485);
nand U36512 (N_36512,N_34407,N_32801);
nor U36513 (N_36513,N_32512,N_34083);
xor U36514 (N_36514,N_34864,N_34924);
xor U36515 (N_36515,N_34425,N_33782);
and U36516 (N_36516,N_33396,N_32570);
or U36517 (N_36517,N_33001,N_32706);
xnor U36518 (N_36518,N_34269,N_32700);
nand U36519 (N_36519,N_33051,N_32910);
nor U36520 (N_36520,N_33341,N_32798);
and U36521 (N_36521,N_33112,N_33644);
or U36522 (N_36522,N_33463,N_33010);
xor U36523 (N_36523,N_32593,N_34587);
and U36524 (N_36524,N_34187,N_33171);
nor U36525 (N_36525,N_34794,N_33588);
nor U36526 (N_36526,N_32907,N_33867);
and U36527 (N_36527,N_33883,N_32655);
nand U36528 (N_36528,N_34708,N_34126);
nand U36529 (N_36529,N_34296,N_33646);
and U36530 (N_36530,N_32657,N_32539);
nor U36531 (N_36531,N_33688,N_34334);
nor U36532 (N_36532,N_33168,N_34642);
xor U36533 (N_36533,N_32600,N_32535);
and U36534 (N_36534,N_33315,N_33641);
nor U36535 (N_36535,N_33295,N_33260);
or U36536 (N_36536,N_34900,N_34495);
nor U36537 (N_36537,N_33491,N_33175);
nand U36538 (N_36538,N_32814,N_33206);
xnor U36539 (N_36539,N_34467,N_33852);
and U36540 (N_36540,N_33420,N_34614);
and U36541 (N_36541,N_33421,N_32586);
nor U36542 (N_36542,N_32693,N_32805);
nand U36543 (N_36543,N_34245,N_32505);
nand U36544 (N_36544,N_34729,N_34885);
nor U36545 (N_36545,N_34538,N_32710);
or U36546 (N_36546,N_33407,N_33651);
nor U36547 (N_36547,N_34950,N_33581);
nor U36548 (N_36548,N_33856,N_33651);
or U36549 (N_36549,N_33695,N_32732);
or U36550 (N_36550,N_33326,N_33341);
nand U36551 (N_36551,N_33533,N_33879);
and U36552 (N_36552,N_33513,N_34397);
or U36553 (N_36553,N_34319,N_33222);
or U36554 (N_36554,N_33070,N_33825);
nand U36555 (N_36555,N_33479,N_32632);
or U36556 (N_36556,N_34629,N_34286);
nand U36557 (N_36557,N_33711,N_32944);
nand U36558 (N_36558,N_33654,N_32803);
xnor U36559 (N_36559,N_34051,N_33796);
and U36560 (N_36560,N_33880,N_33609);
and U36561 (N_36561,N_34167,N_33222);
and U36562 (N_36562,N_34394,N_33743);
or U36563 (N_36563,N_34661,N_34785);
and U36564 (N_36564,N_32914,N_34381);
xnor U36565 (N_36565,N_33468,N_33155);
xnor U36566 (N_36566,N_32809,N_32854);
nand U36567 (N_36567,N_33382,N_34468);
xnor U36568 (N_36568,N_33711,N_32903);
nand U36569 (N_36569,N_32640,N_32975);
nand U36570 (N_36570,N_32605,N_34158);
xor U36571 (N_36571,N_33728,N_33103);
nor U36572 (N_36572,N_34386,N_33829);
nor U36573 (N_36573,N_33924,N_34221);
or U36574 (N_36574,N_34012,N_34471);
nand U36575 (N_36575,N_33884,N_33706);
xor U36576 (N_36576,N_33312,N_33154);
and U36577 (N_36577,N_32922,N_33152);
or U36578 (N_36578,N_33432,N_34789);
xnor U36579 (N_36579,N_34739,N_34503);
xnor U36580 (N_36580,N_33662,N_33488);
nand U36581 (N_36581,N_32619,N_34162);
xnor U36582 (N_36582,N_33911,N_33954);
and U36583 (N_36583,N_32547,N_32796);
nand U36584 (N_36584,N_32734,N_32632);
nand U36585 (N_36585,N_33097,N_32609);
and U36586 (N_36586,N_33393,N_34264);
nand U36587 (N_36587,N_32592,N_32856);
nor U36588 (N_36588,N_32629,N_34932);
xor U36589 (N_36589,N_34496,N_32866);
nand U36590 (N_36590,N_34850,N_33635);
nor U36591 (N_36591,N_33820,N_32732);
xnor U36592 (N_36592,N_32511,N_34650);
xor U36593 (N_36593,N_32688,N_34113);
and U36594 (N_36594,N_32555,N_34447);
or U36595 (N_36595,N_33321,N_33428);
nand U36596 (N_36596,N_33199,N_32580);
or U36597 (N_36597,N_32706,N_34781);
nor U36598 (N_36598,N_34379,N_33793);
xor U36599 (N_36599,N_34537,N_34243);
or U36600 (N_36600,N_33834,N_34067);
and U36601 (N_36601,N_32649,N_32800);
or U36602 (N_36602,N_33479,N_34704);
xnor U36603 (N_36603,N_34022,N_32569);
and U36604 (N_36604,N_33252,N_34130);
and U36605 (N_36605,N_34098,N_34120);
nor U36606 (N_36606,N_34852,N_33268);
nand U36607 (N_36607,N_34525,N_34199);
nor U36608 (N_36608,N_33733,N_33717);
and U36609 (N_36609,N_33820,N_34097);
or U36610 (N_36610,N_32533,N_34460);
or U36611 (N_36611,N_34140,N_34833);
nand U36612 (N_36612,N_33027,N_33942);
xnor U36613 (N_36613,N_33333,N_33041);
or U36614 (N_36614,N_34120,N_34976);
xnor U36615 (N_36615,N_34166,N_33932);
and U36616 (N_36616,N_34277,N_32707);
nand U36617 (N_36617,N_34666,N_33945);
xor U36618 (N_36618,N_33138,N_34546);
nand U36619 (N_36619,N_33591,N_34228);
or U36620 (N_36620,N_33539,N_33772);
and U36621 (N_36621,N_33578,N_34854);
and U36622 (N_36622,N_33530,N_32617);
and U36623 (N_36623,N_32714,N_32964);
or U36624 (N_36624,N_33486,N_34577);
nand U36625 (N_36625,N_33508,N_34039);
nand U36626 (N_36626,N_33705,N_34528);
nand U36627 (N_36627,N_33821,N_34254);
and U36628 (N_36628,N_34507,N_34552);
and U36629 (N_36629,N_34582,N_33548);
nand U36630 (N_36630,N_32702,N_33823);
nor U36631 (N_36631,N_34909,N_33953);
nor U36632 (N_36632,N_33185,N_34884);
nor U36633 (N_36633,N_33803,N_34985);
xor U36634 (N_36634,N_33750,N_33749);
and U36635 (N_36635,N_33033,N_32802);
nor U36636 (N_36636,N_33915,N_33414);
nor U36637 (N_36637,N_34176,N_34923);
xnor U36638 (N_36638,N_33663,N_32703);
nor U36639 (N_36639,N_33161,N_34399);
nor U36640 (N_36640,N_33268,N_34473);
and U36641 (N_36641,N_34592,N_33456);
nand U36642 (N_36642,N_33961,N_33598);
nand U36643 (N_36643,N_33428,N_32884);
nor U36644 (N_36644,N_34984,N_33115);
and U36645 (N_36645,N_33402,N_34493);
xor U36646 (N_36646,N_32656,N_34215);
and U36647 (N_36647,N_32789,N_34910);
nor U36648 (N_36648,N_34266,N_33171);
and U36649 (N_36649,N_32691,N_34661);
or U36650 (N_36650,N_33939,N_32563);
and U36651 (N_36651,N_32593,N_33776);
nor U36652 (N_36652,N_32532,N_33378);
or U36653 (N_36653,N_33199,N_34422);
nor U36654 (N_36654,N_32644,N_33256);
and U36655 (N_36655,N_33416,N_34798);
and U36656 (N_36656,N_34237,N_33869);
xnor U36657 (N_36657,N_34201,N_34128);
nand U36658 (N_36658,N_32688,N_32984);
nand U36659 (N_36659,N_34873,N_32685);
or U36660 (N_36660,N_34674,N_32586);
nor U36661 (N_36661,N_33847,N_33121);
and U36662 (N_36662,N_34099,N_34130);
xnor U36663 (N_36663,N_34465,N_32851);
nand U36664 (N_36664,N_33156,N_33943);
nand U36665 (N_36665,N_34150,N_32731);
xor U36666 (N_36666,N_34586,N_33895);
or U36667 (N_36667,N_32990,N_33150);
nand U36668 (N_36668,N_33080,N_33529);
xor U36669 (N_36669,N_34669,N_34254);
nor U36670 (N_36670,N_33760,N_34752);
nand U36671 (N_36671,N_34018,N_33484);
xor U36672 (N_36672,N_33280,N_32577);
and U36673 (N_36673,N_34838,N_34996);
and U36674 (N_36674,N_32979,N_32517);
xnor U36675 (N_36675,N_34309,N_33083);
nor U36676 (N_36676,N_32626,N_34881);
nor U36677 (N_36677,N_33667,N_33725);
and U36678 (N_36678,N_33266,N_32634);
nand U36679 (N_36679,N_33779,N_33879);
or U36680 (N_36680,N_33974,N_34296);
nand U36681 (N_36681,N_34994,N_32501);
and U36682 (N_36682,N_33443,N_32733);
or U36683 (N_36683,N_33633,N_33369);
xor U36684 (N_36684,N_33754,N_32843);
xnor U36685 (N_36685,N_33438,N_33047);
and U36686 (N_36686,N_34477,N_33563);
nand U36687 (N_36687,N_34279,N_34818);
or U36688 (N_36688,N_33092,N_33121);
nor U36689 (N_36689,N_34796,N_33720);
xnor U36690 (N_36690,N_34901,N_34872);
xor U36691 (N_36691,N_33756,N_32598);
or U36692 (N_36692,N_33240,N_34367);
and U36693 (N_36693,N_34437,N_34979);
nor U36694 (N_36694,N_33869,N_32605);
or U36695 (N_36695,N_32844,N_33515);
xor U36696 (N_36696,N_32902,N_32678);
and U36697 (N_36697,N_33390,N_33336);
and U36698 (N_36698,N_32526,N_33455);
xor U36699 (N_36699,N_33888,N_34476);
nand U36700 (N_36700,N_33577,N_33683);
nand U36701 (N_36701,N_32765,N_34399);
xnor U36702 (N_36702,N_32830,N_33485);
xnor U36703 (N_36703,N_33250,N_34851);
and U36704 (N_36704,N_33813,N_33495);
xnor U36705 (N_36705,N_33711,N_34824);
and U36706 (N_36706,N_33189,N_33806);
xor U36707 (N_36707,N_34068,N_34467);
or U36708 (N_36708,N_34141,N_33406);
nand U36709 (N_36709,N_34978,N_32927);
nand U36710 (N_36710,N_34684,N_34932);
nor U36711 (N_36711,N_34324,N_33895);
xnor U36712 (N_36712,N_32663,N_33733);
and U36713 (N_36713,N_34086,N_33062);
xor U36714 (N_36714,N_33515,N_34548);
xor U36715 (N_36715,N_34010,N_34363);
or U36716 (N_36716,N_34173,N_32738);
and U36717 (N_36717,N_33065,N_34978);
and U36718 (N_36718,N_33402,N_34996);
nand U36719 (N_36719,N_33817,N_32718);
xor U36720 (N_36720,N_34373,N_34951);
xor U36721 (N_36721,N_34921,N_33348);
and U36722 (N_36722,N_34060,N_32756);
xor U36723 (N_36723,N_33401,N_34107);
xor U36724 (N_36724,N_33160,N_34129);
nor U36725 (N_36725,N_33016,N_34038);
and U36726 (N_36726,N_32735,N_34877);
and U36727 (N_36727,N_34146,N_32999);
nor U36728 (N_36728,N_34072,N_32825);
xnor U36729 (N_36729,N_33346,N_33795);
nand U36730 (N_36730,N_34177,N_33726);
or U36731 (N_36731,N_33952,N_33134);
and U36732 (N_36732,N_32641,N_34778);
or U36733 (N_36733,N_32564,N_34409);
and U36734 (N_36734,N_33444,N_32837);
nor U36735 (N_36735,N_34420,N_34802);
or U36736 (N_36736,N_34376,N_33010);
or U36737 (N_36737,N_32822,N_34362);
and U36738 (N_36738,N_33129,N_34896);
and U36739 (N_36739,N_33271,N_32769);
nand U36740 (N_36740,N_34664,N_34063);
nand U36741 (N_36741,N_32948,N_34000);
or U36742 (N_36742,N_32792,N_34594);
xor U36743 (N_36743,N_34367,N_33284);
or U36744 (N_36744,N_34389,N_34314);
nor U36745 (N_36745,N_34961,N_33719);
nor U36746 (N_36746,N_33421,N_33186);
xor U36747 (N_36747,N_33948,N_34347);
and U36748 (N_36748,N_33438,N_34030);
and U36749 (N_36749,N_34422,N_34778);
nor U36750 (N_36750,N_33520,N_32990);
nor U36751 (N_36751,N_34936,N_32718);
xnor U36752 (N_36752,N_33674,N_34509);
nand U36753 (N_36753,N_32532,N_33356);
nand U36754 (N_36754,N_33843,N_34238);
or U36755 (N_36755,N_32897,N_33554);
or U36756 (N_36756,N_33405,N_34190);
and U36757 (N_36757,N_34079,N_33805);
or U36758 (N_36758,N_33653,N_34062);
nor U36759 (N_36759,N_33687,N_34322);
nand U36760 (N_36760,N_34160,N_32761);
and U36761 (N_36761,N_34121,N_33499);
xor U36762 (N_36762,N_32842,N_33804);
nor U36763 (N_36763,N_33895,N_34482);
and U36764 (N_36764,N_32624,N_32608);
and U36765 (N_36765,N_33203,N_34635);
xnor U36766 (N_36766,N_34638,N_33025);
and U36767 (N_36767,N_34777,N_34334);
nor U36768 (N_36768,N_33295,N_34366);
nor U36769 (N_36769,N_33362,N_34086);
xnor U36770 (N_36770,N_34095,N_33163);
nor U36771 (N_36771,N_33743,N_34870);
nor U36772 (N_36772,N_32877,N_34342);
and U36773 (N_36773,N_32655,N_33789);
xor U36774 (N_36774,N_32994,N_33985);
and U36775 (N_36775,N_32623,N_34076);
xor U36776 (N_36776,N_33442,N_32832);
and U36777 (N_36777,N_33005,N_34668);
and U36778 (N_36778,N_34583,N_34414);
nor U36779 (N_36779,N_34932,N_33265);
nor U36780 (N_36780,N_33542,N_33451);
nor U36781 (N_36781,N_33414,N_34610);
or U36782 (N_36782,N_33139,N_32540);
nand U36783 (N_36783,N_33095,N_34383);
nand U36784 (N_36784,N_33066,N_33955);
and U36785 (N_36785,N_33838,N_34929);
or U36786 (N_36786,N_32912,N_32839);
nor U36787 (N_36787,N_34614,N_33340);
nand U36788 (N_36788,N_32871,N_32710);
xor U36789 (N_36789,N_33308,N_33110);
xor U36790 (N_36790,N_34611,N_33523);
nor U36791 (N_36791,N_34424,N_34294);
xor U36792 (N_36792,N_33263,N_34522);
nor U36793 (N_36793,N_32780,N_34527);
and U36794 (N_36794,N_34768,N_33308);
xnor U36795 (N_36795,N_33158,N_33239);
nand U36796 (N_36796,N_33970,N_33418);
or U36797 (N_36797,N_32565,N_33830);
xnor U36798 (N_36798,N_34579,N_33273);
xnor U36799 (N_36799,N_34533,N_34486);
or U36800 (N_36800,N_34802,N_33905);
or U36801 (N_36801,N_32929,N_34791);
xor U36802 (N_36802,N_34223,N_34916);
nor U36803 (N_36803,N_32874,N_34577);
or U36804 (N_36804,N_33449,N_33379);
or U36805 (N_36805,N_32575,N_33392);
or U36806 (N_36806,N_32595,N_33499);
nand U36807 (N_36807,N_32558,N_33129);
nand U36808 (N_36808,N_33646,N_33424);
or U36809 (N_36809,N_34444,N_34459);
or U36810 (N_36810,N_33404,N_34980);
nand U36811 (N_36811,N_34599,N_33327);
xor U36812 (N_36812,N_34207,N_33543);
or U36813 (N_36813,N_33792,N_33912);
or U36814 (N_36814,N_34063,N_32822);
nand U36815 (N_36815,N_33413,N_33491);
nor U36816 (N_36816,N_34764,N_33800);
and U36817 (N_36817,N_33316,N_33677);
or U36818 (N_36818,N_33975,N_33241);
or U36819 (N_36819,N_33709,N_34414);
or U36820 (N_36820,N_34298,N_34293);
nand U36821 (N_36821,N_32638,N_32865);
nor U36822 (N_36822,N_33166,N_34652);
nor U36823 (N_36823,N_32671,N_32583);
nor U36824 (N_36824,N_32783,N_33156);
and U36825 (N_36825,N_33249,N_33291);
and U36826 (N_36826,N_34261,N_34202);
and U36827 (N_36827,N_34299,N_34149);
nor U36828 (N_36828,N_32560,N_32657);
nand U36829 (N_36829,N_33329,N_32584);
and U36830 (N_36830,N_32965,N_33454);
and U36831 (N_36831,N_32998,N_32530);
nor U36832 (N_36832,N_34761,N_32597);
nor U36833 (N_36833,N_34072,N_32949);
nand U36834 (N_36834,N_34434,N_34207);
xor U36835 (N_36835,N_32903,N_33083);
nor U36836 (N_36836,N_33316,N_33620);
and U36837 (N_36837,N_34125,N_34424);
nand U36838 (N_36838,N_34827,N_33100);
xnor U36839 (N_36839,N_32959,N_34906);
or U36840 (N_36840,N_33821,N_33372);
and U36841 (N_36841,N_32937,N_34723);
xor U36842 (N_36842,N_32605,N_32744);
or U36843 (N_36843,N_33738,N_33556);
nor U36844 (N_36844,N_34881,N_34092);
nor U36845 (N_36845,N_33239,N_32933);
nor U36846 (N_36846,N_34872,N_34074);
nor U36847 (N_36847,N_33117,N_33780);
and U36848 (N_36848,N_33381,N_34774);
and U36849 (N_36849,N_32801,N_32817);
and U36850 (N_36850,N_34161,N_33140);
or U36851 (N_36851,N_34893,N_34134);
nor U36852 (N_36852,N_32687,N_33653);
nor U36853 (N_36853,N_34515,N_33609);
and U36854 (N_36854,N_32764,N_34563);
and U36855 (N_36855,N_33593,N_34003);
nand U36856 (N_36856,N_32660,N_33964);
xnor U36857 (N_36857,N_34412,N_34903);
nand U36858 (N_36858,N_33460,N_34479);
and U36859 (N_36859,N_34792,N_33676);
nor U36860 (N_36860,N_32762,N_34948);
nor U36861 (N_36861,N_34669,N_33649);
nand U36862 (N_36862,N_34978,N_34933);
xor U36863 (N_36863,N_34130,N_33638);
and U36864 (N_36864,N_33619,N_33171);
nor U36865 (N_36865,N_33473,N_33030);
nor U36866 (N_36866,N_34204,N_34529);
xnor U36867 (N_36867,N_34732,N_33548);
xnor U36868 (N_36868,N_33648,N_32950);
and U36869 (N_36869,N_32927,N_34666);
xnor U36870 (N_36870,N_33399,N_33649);
nor U36871 (N_36871,N_34723,N_33876);
nand U36872 (N_36872,N_34698,N_32930);
and U36873 (N_36873,N_34437,N_34285);
nand U36874 (N_36874,N_32567,N_34774);
or U36875 (N_36875,N_34393,N_32562);
xor U36876 (N_36876,N_33546,N_33039);
and U36877 (N_36877,N_34534,N_33591);
and U36878 (N_36878,N_33809,N_33333);
nor U36879 (N_36879,N_32636,N_33865);
nand U36880 (N_36880,N_33748,N_34319);
nor U36881 (N_36881,N_34859,N_32973);
nor U36882 (N_36882,N_34173,N_32771);
nand U36883 (N_36883,N_33645,N_32611);
nor U36884 (N_36884,N_32978,N_34215);
nor U36885 (N_36885,N_34518,N_32602);
nand U36886 (N_36886,N_33809,N_34739);
nor U36887 (N_36887,N_34367,N_34507);
nand U36888 (N_36888,N_33670,N_33153);
or U36889 (N_36889,N_34710,N_34676);
xor U36890 (N_36890,N_32870,N_34891);
nor U36891 (N_36891,N_32856,N_33474);
and U36892 (N_36892,N_33889,N_32783);
or U36893 (N_36893,N_34725,N_34219);
or U36894 (N_36894,N_33484,N_33538);
and U36895 (N_36895,N_32784,N_33880);
nand U36896 (N_36896,N_33554,N_33253);
and U36897 (N_36897,N_33846,N_34520);
or U36898 (N_36898,N_32800,N_34494);
nor U36899 (N_36899,N_33302,N_33317);
and U36900 (N_36900,N_33663,N_33602);
and U36901 (N_36901,N_34688,N_33328);
and U36902 (N_36902,N_33822,N_33120);
or U36903 (N_36903,N_33072,N_33633);
and U36904 (N_36904,N_34254,N_34020);
nand U36905 (N_36905,N_34598,N_32564);
xnor U36906 (N_36906,N_34522,N_32937);
nand U36907 (N_36907,N_32605,N_33535);
xor U36908 (N_36908,N_33146,N_33218);
and U36909 (N_36909,N_33225,N_34158);
xnor U36910 (N_36910,N_34673,N_33978);
or U36911 (N_36911,N_33971,N_32751);
and U36912 (N_36912,N_33015,N_34018);
nand U36913 (N_36913,N_34829,N_33489);
xnor U36914 (N_36914,N_33410,N_33966);
or U36915 (N_36915,N_32610,N_34901);
nor U36916 (N_36916,N_32907,N_32560);
nand U36917 (N_36917,N_32976,N_33733);
and U36918 (N_36918,N_33146,N_33162);
nand U36919 (N_36919,N_32563,N_34888);
or U36920 (N_36920,N_34333,N_33545);
or U36921 (N_36921,N_33037,N_34761);
xor U36922 (N_36922,N_33188,N_34633);
or U36923 (N_36923,N_32561,N_33118);
nand U36924 (N_36924,N_33812,N_34143);
nor U36925 (N_36925,N_33017,N_34355);
xor U36926 (N_36926,N_33923,N_33320);
and U36927 (N_36927,N_34470,N_33024);
xnor U36928 (N_36928,N_34038,N_33765);
nor U36929 (N_36929,N_33500,N_33310);
xnor U36930 (N_36930,N_34159,N_34373);
nor U36931 (N_36931,N_32545,N_34480);
nand U36932 (N_36932,N_33886,N_32988);
and U36933 (N_36933,N_33469,N_32668);
nand U36934 (N_36934,N_33489,N_33431);
xor U36935 (N_36935,N_32509,N_33231);
nor U36936 (N_36936,N_34753,N_34248);
xor U36937 (N_36937,N_33041,N_34010);
nand U36938 (N_36938,N_32934,N_34706);
and U36939 (N_36939,N_33515,N_32596);
or U36940 (N_36940,N_34083,N_33576);
or U36941 (N_36941,N_33001,N_32588);
xnor U36942 (N_36942,N_34987,N_34719);
or U36943 (N_36943,N_32781,N_33216);
or U36944 (N_36944,N_33143,N_33491);
xnor U36945 (N_36945,N_34506,N_34801);
nand U36946 (N_36946,N_33284,N_33390);
nand U36947 (N_36947,N_34948,N_34490);
or U36948 (N_36948,N_33195,N_32953);
nor U36949 (N_36949,N_33441,N_32944);
or U36950 (N_36950,N_32694,N_32831);
xor U36951 (N_36951,N_33246,N_34593);
and U36952 (N_36952,N_33020,N_33466);
or U36953 (N_36953,N_34586,N_34296);
nand U36954 (N_36954,N_34811,N_33840);
or U36955 (N_36955,N_33934,N_32528);
or U36956 (N_36956,N_33421,N_33058);
nand U36957 (N_36957,N_33816,N_33907);
nand U36958 (N_36958,N_33201,N_33956);
xnor U36959 (N_36959,N_34076,N_34408);
nand U36960 (N_36960,N_32647,N_34321);
nor U36961 (N_36961,N_33203,N_34557);
nor U36962 (N_36962,N_34901,N_33067);
nand U36963 (N_36963,N_34145,N_34360);
nand U36964 (N_36964,N_33412,N_32582);
nand U36965 (N_36965,N_33887,N_34939);
nor U36966 (N_36966,N_32570,N_33938);
xor U36967 (N_36967,N_34189,N_34638);
nor U36968 (N_36968,N_34129,N_34784);
nand U36969 (N_36969,N_33270,N_34232);
or U36970 (N_36970,N_32853,N_34881);
or U36971 (N_36971,N_33842,N_34603);
xnor U36972 (N_36972,N_33992,N_34498);
nand U36973 (N_36973,N_33202,N_32764);
xor U36974 (N_36974,N_33932,N_32659);
nand U36975 (N_36975,N_33986,N_33036);
or U36976 (N_36976,N_34110,N_33496);
and U36977 (N_36977,N_33764,N_33908);
nor U36978 (N_36978,N_34913,N_33345);
nor U36979 (N_36979,N_34871,N_34569);
and U36980 (N_36980,N_34580,N_33169);
and U36981 (N_36981,N_34010,N_33638);
and U36982 (N_36982,N_33195,N_33569);
or U36983 (N_36983,N_33561,N_32967);
xnor U36984 (N_36984,N_32630,N_33364);
nor U36985 (N_36985,N_33517,N_34205);
or U36986 (N_36986,N_34951,N_32595);
xor U36987 (N_36987,N_33477,N_32660);
xnor U36988 (N_36988,N_32885,N_34198);
or U36989 (N_36989,N_34923,N_33075);
nor U36990 (N_36990,N_33009,N_33419);
nand U36991 (N_36991,N_34651,N_33314);
or U36992 (N_36992,N_33643,N_34036);
nor U36993 (N_36993,N_34307,N_33606);
or U36994 (N_36994,N_33021,N_34538);
and U36995 (N_36995,N_33833,N_33791);
and U36996 (N_36996,N_34742,N_33310);
xor U36997 (N_36997,N_34100,N_32745);
xor U36998 (N_36998,N_33902,N_34810);
nand U36999 (N_36999,N_34496,N_32856);
xnor U37000 (N_37000,N_34789,N_34143);
and U37001 (N_37001,N_33308,N_33868);
xor U37002 (N_37002,N_33399,N_33312);
and U37003 (N_37003,N_34529,N_34861);
or U37004 (N_37004,N_32964,N_33350);
nand U37005 (N_37005,N_34462,N_34305);
nor U37006 (N_37006,N_33779,N_34916);
or U37007 (N_37007,N_33366,N_33519);
nor U37008 (N_37008,N_33352,N_33405);
or U37009 (N_37009,N_34416,N_34137);
nand U37010 (N_37010,N_33729,N_34872);
nor U37011 (N_37011,N_34741,N_34121);
nor U37012 (N_37012,N_33283,N_33208);
nand U37013 (N_37013,N_34456,N_34381);
xor U37014 (N_37014,N_32883,N_33730);
xor U37015 (N_37015,N_34028,N_34351);
nand U37016 (N_37016,N_32572,N_34564);
xnor U37017 (N_37017,N_34139,N_32550);
and U37018 (N_37018,N_34139,N_32558);
nor U37019 (N_37019,N_34417,N_32580);
nand U37020 (N_37020,N_34987,N_34371);
and U37021 (N_37021,N_33387,N_34040);
xor U37022 (N_37022,N_32638,N_33988);
nor U37023 (N_37023,N_34959,N_32914);
and U37024 (N_37024,N_34718,N_34257);
nor U37025 (N_37025,N_33896,N_32917);
nand U37026 (N_37026,N_34186,N_33211);
and U37027 (N_37027,N_34877,N_32986);
nand U37028 (N_37028,N_33037,N_33374);
nor U37029 (N_37029,N_34289,N_33305);
xnor U37030 (N_37030,N_34435,N_33427);
nor U37031 (N_37031,N_34738,N_32731);
nor U37032 (N_37032,N_33393,N_32673);
nor U37033 (N_37033,N_32810,N_33224);
nand U37034 (N_37034,N_33355,N_34043);
and U37035 (N_37035,N_32752,N_33674);
or U37036 (N_37036,N_33218,N_34880);
or U37037 (N_37037,N_34622,N_33086);
xnor U37038 (N_37038,N_34980,N_33287);
nor U37039 (N_37039,N_33655,N_33170);
nand U37040 (N_37040,N_34053,N_32892);
or U37041 (N_37041,N_34083,N_33685);
nand U37042 (N_37042,N_34914,N_34083);
and U37043 (N_37043,N_33006,N_34198);
xnor U37044 (N_37044,N_33453,N_33713);
or U37045 (N_37045,N_33537,N_34750);
nand U37046 (N_37046,N_32500,N_34566);
nor U37047 (N_37047,N_34362,N_34281);
nand U37048 (N_37048,N_33801,N_33154);
nor U37049 (N_37049,N_34570,N_32983);
and U37050 (N_37050,N_33207,N_34970);
xor U37051 (N_37051,N_34516,N_33116);
xor U37052 (N_37052,N_34398,N_32712);
xnor U37053 (N_37053,N_33553,N_34253);
xor U37054 (N_37054,N_32938,N_34254);
nand U37055 (N_37055,N_33972,N_32765);
nand U37056 (N_37056,N_33689,N_32649);
xnor U37057 (N_37057,N_34194,N_34853);
or U37058 (N_37058,N_34680,N_34685);
and U37059 (N_37059,N_33513,N_34070);
and U37060 (N_37060,N_33396,N_34335);
or U37061 (N_37061,N_32987,N_34405);
nor U37062 (N_37062,N_33081,N_34833);
xor U37063 (N_37063,N_33120,N_32511);
xor U37064 (N_37064,N_34112,N_34665);
nor U37065 (N_37065,N_33636,N_34599);
nor U37066 (N_37066,N_32852,N_34005);
or U37067 (N_37067,N_32741,N_33737);
and U37068 (N_37068,N_34709,N_33848);
nor U37069 (N_37069,N_33510,N_32527);
or U37070 (N_37070,N_33054,N_33285);
nor U37071 (N_37071,N_34632,N_34771);
or U37072 (N_37072,N_34380,N_34376);
nand U37073 (N_37073,N_32960,N_33433);
nand U37074 (N_37074,N_33682,N_32727);
and U37075 (N_37075,N_33067,N_34975);
nand U37076 (N_37076,N_32641,N_33709);
xnor U37077 (N_37077,N_33157,N_32983);
xor U37078 (N_37078,N_34623,N_32537);
nor U37079 (N_37079,N_34264,N_33225);
nand U37080 (N_37080,N_32991,N_34205);
xor U37081 (N_37081,N_33860,N_34529);
and U37082 (N_37082,N_33156,N_34058);
nand U37083 (N_37083,N_34766,N_33477);
xor U37084 (N_37084,N_34937,N_32903);
and U37085 (N_37085,N_32597,N_32905);
nand U37086 (N_37086,N_33854,N_34554);
nand U37087 (N_37087,N_34748,N_33302);
and U37088 (N_37088,N_33387,N_34152);
or U37089 (N_37089,N_33433,N_32609);
nand U37090 (N_37090,N_33658,N_34796);
or U37091 (N_37091,N_34873,N_34054);
nand U37092 (N_37092,N_33767,N_33105);
xnor U37093 (N_37093,N_34147,N_33961);
or U37094 (N_37094,N_32950,N_33899);
nor U37095 (N_37095,N_33869,N_33720);
nand U37096 (N_37096,N_34610,N_32665);
or U37097 (N_37097,N_33852,N_33453);
nand U37098 (N_37098,N_32535,N_33724);
nor U37099 (N_37099,N_34874,N_32719);
xor U37100 (N_37100,N_33659,N_32992);
xor U37101 (N_37101,N_33910,N_33671);
xor U37102 (N_37102,N_33756,N_32702);
nor U37103 (N_37103,N_33793,N_34473);
or U37104 (N_37104,N_34930,N_33429);
nor U37105 (N_37105,N_34436,N_33342);
and U37106 (N_37106,N_34273,N_34242);
or U37107 (N_37107,N_34621,N_34248);
xnor U37108 (N_37108,N_33071,N_34196);
xor U37109 (N_37109,N_34583,N_32591);
xor U37110 (N_37110,N_34100,N_34096);
or U37111 (N_37111,N_33211,N_34633);
or U37112 (N_37112,N_32579,N_32966);
or U37113 (N_37113,N_33398,N_33200);
nand U37114 (N_37114,N_33262,N_34553);
and U37115 (N_37115,N_33505,N_33501);
nor U37116 (N_37116,N_34021,N_33627);
xor U37117 (N_37117,N_32733,N_33756);
nor U37118 (N_37118,N_34482,N_34225);
and U37119 (N_37119,N_32998,N_33569);
xor U37120 (N_37120,N_34808,N_34612);
nor U37121 (N_37121,N_34757,N_34674);
nand U37122 (N_37122,N_34416,N_32993);
nor U37123 (N_37123,N_33935,N_34135);
nand U37124 (N_37124,N_33583,N_32720);
and U37125 (N_37125,N_33950,N_34130);
and U37126 (N_37126,N_34471,N_32707);
nor U37127 (N_37127,N_34798,N_32817);
xor U37128 (N_37128,N_34380,N_32526);
and U37129 (N_37129,N_32638,N_34507);
nor U37130 (N_37130,N_32528,N_34102);
or U37131 (N_37131,N_33243,N_32994);
and U37132 (N_37132,N_34628,N_33267);
nor U37133 (N_37133,N_34049,N_34088);
and U37134 (N_37134,N_34746,N_33477);
nand U37135 (N_37135,N_34247,N_33749);
nor U37136 (N_37136,N_33533,N_33764);
or U37137 (N_37137,N_33583,N_33999);
xnor U37138 (N_37138,N_33001,N_34038);
xnor U37139 (N_37139,N_33486,N_34936);
xor U37140 (N_37140,N_34552,N_34572);
nand U37141 (N_37141,N_34726,N_34624);
and U37142 (N_37142,N_32703,N_33505);
xnor U37143 (N_37143,N_34852,N_33799);
xnor U37144 (N_37144,N_33928,N_34678);
nand U37145 (N_37145,N_34468,N_32697);
or U37146 (N_37146,N_34076,N_34804);
and U37147 (N_37147,N_33806,N_32992);
nand U37148 (N_37148,N_34826,N_33351);
nand U37149 (N_37149,N_34592,N_34975);
and U37150 (N_37150,N_34138,N_34879);
xnor U37151 (N_37151,N_33322,N_34548);
xor U37152 (N_37152,N_34461,N_33348);
nand U37153 (N_37153,N_34313,N_33264);
nor U37154 (N_37154,N_34335,N_34607);
and U37155 (N_37155,N_34329,N_34616);
or U37156 (N_37156,N_34764,N_33003);
or U37157 (N_37157,N_32862,N_34411);
nand U37158 (N_37158,N_34424,N_34781);
and U37159 (N_37159,N_32957,N_33937);
xnor U37160 (N_37160,N_34990,N_32992);
nor U37161 (N_37161,N_34833,N_34142);
and U37162 (N_37162,N_33822,N_34456);
xnor U37163 (N_37163,N_33039,N_34661);
or U37164 (N_37164,N_33794,N_33643);
xor U37165 (N_37165,N_33829,N_32925);
xnor U37166 (N_37166,N_33059,N_32908);
or U37167 (N_37167,N_33049,N_32572);
and U37168 (N_37168,N_34003,N_32524);
nor U37169 (N_37169,N_34574,N_33852);
or U37170 (N_37170,N_34343,N_33161);
xnor U37171 (N_37171,N_32955,N_32717);
or U37172 (N_37172,N_34614,N_34590);
xor U37173 (N_37173,N_32841,N_34487);
nor U37174 (N_37174,N_32778,N_34687);
or U37175 (N_37175,N_33265,N_33234);
xnor U37176 (N_37176,N_34769,N_33229);
xnor U37177 (N_37177,N_33330,N_34053);
nand U37178 (N_37178,N_33208,N_34990);
nand U37179 (N_37179,N_33283,N_33509);
xor U37180 (N_37180,N_32703,N_34274);
or U37181 (N_37181,N_32675,N_34839);
or U37182 (N_37182,N_33120,N_33186);
or U37183 (N_37183,N_34022,N_34099);
and U37184 (N_37184,N_32785,N_34825);
nand U37185 (N_37185,N_32893,N_33581);
nand U37186 (N_37186,N_34784,N_33570);
xnor U37187 (N_37187,N_34327,N_34962);
and U37188 (N_37188,N_33796,N_34634);
nor U37189 (N_37189,N_34836,N_32944);
or U37190 (N_37190,N_33661,N_34786);
or U37191 (N_37191,N_34912,N_33621);
xnor U37192 (N_37192,N_32714,N_33314);
xnor U37193 (N_37193,N_33490,N_33344);
xnor U37194 (N_37194,N_32551,N_33638);
xor U37195 (N_37195,N_34321,N_32899);
nor U37196 (N_37196,N_34447,N_34149);
or U37197 (N_37197,N_34637,N_34108);
xnor U37198 (N_37198,N_33029,N_33770);
and U37199 (N_37199,N_33714,N_32651);
nor U37200 (N_37200,N_32820,N_32595);
nor U37201 (N_37201,N_32638,N_34758);
nand U37202 (N_37202,N_33382,N_33623);
nand U37203 (N_37203,N_33738,N_32504);
xnor U37204 (N_37204,N_32616,N_33620);
or U37205 (N_37205,N_34308,N_34568);
xor U37206 (N_37206,N_33574,N_33016);
nor U37207 (N_37207,N_33145,N_32926);
nor U37208 (N_37208,N_34823,N_34870);
xnor U37209 (N_37209,N_34365,N_33910);
or U37210 (N_37210,N_32959,N_34528);
xnor U37211 (N_37211,N_34536,N_33946);
and U37212 (N_37212,N_32547,N_34774);
nand U37213 (N_37213,N_34925,N_34965);
nor U37214 (N_37214,N_34803,N_32640);
xor U37215 (N_37215,N_34899,N_32593);
nor U37216 (N_37216,N_32819,N_33951);
nand U37217 (N_37217,N_34615,N_33304);
nor U37218 (N_37218,N_32646,N_32730);
xnor U37219 (N_37219,N_32908,N_34008);
nand U37220 (N_37220,N_32811,N_32851);
nor U37221 (N_37221,N_33025,N_32748);
nand U37222 (N_37222,N_33702,N_32596);
and U37223 (N_37223,N_34935,N_33499);
xnor U37224 (N_37224,N_34567,N_33043);
nand U37225 (N_37225,N_34034,N_33091);
nand U37226 (N_37226,N_34869,N_34126);
nand U37227 (N_37227,N_33958,N_34158);
and U37228 (N_37228,N_32990,N_34677);
and U37229 (N_37229,N_33289,N_32841);
nor U37230 (N_37230,N_34063,N_32775);
nor U37231 (N_37231,N_33885,N_33870);
nand U37232 (N_37232,N_33212,N_34093);
or U37233 (N_37233,N_34297,N_33908);
nand U37234 (N_37234,N_34808,N_33375);
nand U37235 (N_37235,N_34079,N_34375);
nor U37236 (N_37236,N_34212,N_34858);
or U37237 (N_37237,N_33782,N_34005);
nor U37238 (N_37238,N_33263,N_33879);
or U37239 (N_37239,N_34470,N_33120);
or U37240 (N_37240,N_33029,N_33053);
or U37241 (N_37241,N_33443,N_33434);
xor U37242 (N_37242,N_34824,N_32882);
nor U37243 (N_37243,N_34158,N_32512);
or U37244 (N_37244,N_34956,N_34326);
and U37245 (N_37245,N_33004,N_34826);
xnor U37246 (N_37246,N_34007,N_34149);
or U37247 (N_37247,N_33910,N_34588);
nand U37248 (N_37248,N_32874,N_32728);
xnor U37249 (N_37249,N_32730,N_34813);
xnor U37250 (N_37250,N_33449,N_34737);
nand U37251 (N_37251,N_33834,N_34810);
xor U37252 (N_37252,N_33351,N_33505);
nor U37253 (N_37253,N_32743,N_32910);
or U37254 (N_37254,N_34484,N_33070);
xnor U37255 (N_37255,N_33868,N_32589);
nor U37256 (N_37256,N_34184,N_34839);
xnor U37257 (N_37257,N_32665,N_34980);
xor U37258 (N_37258,N_32635,N_33993);
nor U37259 (N_37259,N_34963,N_33657);
or U37260 (N_37260,N_34850,N_33589);
xnor U37261 (N_37261,N_34063,N_34142);
and U37262 (N_37262,N_34511,N_34273);
and U37263 (N_37263,N_34375,N_34625);
nor U37264 (N_37264,N_33816,N_32846);
nand U37265 (N_37265,N_34196,N_34454);
and U37266 (N_37266,N_34975,N_33074);
nor U37267 (N_37267,N_34003,N_32644);
nor U37268 (N_37268,N_34189,N_32742);
and U37269 (N_37269,N_33440,N_33904);
nand U37270 (N_37270,N_32729,N_34215);
and U37271 (N_37271,N_32590,N_32557);
and U37272 (N_37272,N_33437,N_32532);
and U37273 (N_37273,N_33287,N_33799);
nand U37274 (N_37274,N_32826,N_34051);
nand U37275 (N_37275,N_32575,N_33351);
nand U37276 (N_37276,N_32990,N_32874);
nor U37277 (N_37277,N_33155,N_33090);
or U37278 (N_37278,N_32661,N_34969);
xor U37279 (N_37279,N_34112,N_33701);
xnor U37280 (N_37280,N_33180,N_34624);
nand U37281 (N_37281,N_34721,N_34034);
xor U37282 (N_37282,N_34101,N_34402);
and U37283 (N_37283,N_33134,N_34048);
or U37284 (N_37284,N_33282,N_34591);
xor U37285 (N_37285,N_33079,N_34099);
xnor U37286 (N_37286,N_33970,N_33457);
nand U37287 (N_37287,N_32962,N_33181);
nand U37288 (N_37288,N_33648,N_34393);
nor U37289 (N_37289,N_33769,N_33293);
or U37290 (N_37290,N_34862,N_34930);
nor U37291 (N_37291,N_33332,N_33166);
and U37292 (N_37292,N_34226,N_34276);
nor U37293 (N_37293,N_33378,N_32885);
and U37294 (N_37294,N_33759,N_34058);
or U37295 (N_37295,N_34107,N_33488);
nor U37296 (N_37296,N_33053,N_34094);
nand U37297 (N_37297,N_34141,N_33429);
nand U37298 (N_37298,N_33556,N_33405);
nand U37299 (N_37299,N_34549,N_32521);
nand U37300 (N_37300,N_34757,N_33034);
nor U37301 (N_37301,N_32934,N_34070);
nand U37302 (N_37302,N_34308,N_33950);
xnor U37303 (N_37303,N_32778,N_34348);
nand U37304 (N_37304,N_33447,N_32908);
nand U37305 (N_37305,N_33129,N_33259);
or U37306 (N_37306,N_34360,N_33340);
or U37307 (N_37307,N_33359,N_32539);
nor U37308 (N_37308,N_33901,N_33405);
and U37309 (N_37309,N_33404,N_33934);
and U37310 (N_37310,N_34291,N_33334);
and U37311 (N_37311,N_34959,N_33853);
nand U37312 (N_37312,N_34668,N_34590);
nand U37313 (N_37313,N_32997,N_33113);
xor U37314 (N_37314,N_34537,N_33484);
or U37315 (N_37315,N_33947,N_34763);
and U37316 (N_37316,N_33235,N_33586);
or U37317 (N_37317,N_32999,N_33751);
nand U37318 (N_37318,N_34442,N_32735);
xnor U37319 (N_37319,N_34125,N_33713);
nor U37320 (N_37320,N_34666,N_32647);
or U37321 (N_37321,N_33504,N_34195);
nand U37322 (N_37322,N_33815,N_32964);
or U37323 (N_37323,N_33540,N_34573);
nand U37324 (N_37324,N_33604,N_34736);
and U37325 (N_37325,N_33935,N_33312);
nor U37326 (N_37326,N_34223,N_34879);
xnor U37327 (N_37327,N_34780,N_33868);
or U37328 (N_37328,N_33374,N_33095);
and U37329 (N_37329,N_32593,N_34160);
nand U37330 (N_37330,N_34179,N_32807);
nand U37331 (N_37331,N_33147,N_34042);
nor U37332 (N_37332,N_33601,N_34812);
nand U37333 (N_37333,N_32690,N_32897);
and U37334 (N_37334,N_33633,N_34102);
nor U37335 (N_37335,N_34572,N_32970);
or U37336 (N_37336,N_34709,N_33539);
xor U37337 (N_37337,N_33043,N_34222);
xor U37338 (N_37338,N_34802,N_34660);
nor U37339 (N_37339,N_34228,N_33004);
xnor U37340 (N_37340,N_33051,N_34042);
or U37341 (N_37341,N_34172,N_32850);
nor U37342 (N_37342,N_34671,N_33830);
nand U37343 (N_37343,N_32716,N_33460);
and U37344 (N_37344,N_33270,N_34546);
nor U37345 (N_37345,N_33315,N_33608);
and U37346 (N_37346,N_33666,N_33052);
xnor U37347 (N_37347,N_34527,N_34864);
nand U37348 (N_37348,N_32974,N_32648);
or U37349 (N_37349,N_32991,N_34638);
xnor U37350 (N_37350,N_34519,N_33551);
or U37351 (N_37351,N_33834,N_33838);
xor U37352 (N_37352,N_34517,N_32823);
nor U37353 (N_37353,N_34533,N_34031);
nor U37354 (N_37354,N_33586,N_33206);
nand U37355 (N_37355,N_32955,N_34175);
and U37356 (N_37356,N_34505,N_33136);
xor U37357 (N_37357,N_33418,N_33373);
and U37358 (N_37358,N_33654,N_33872);
or U37359 (N_37359,N_34793,N_32609);
nor U37360 (N_37360,N_33228,N_34907);
or U37361 (N_37361,N_32504,N_34670);
or U37362 (N_37362,N_33833,N_34928);
and U37363 (N_37363,N_33584,N_33789);
nand U37364 (N_37364,N_32813,N_33862);
nor U37365 (N_37365,N_32683,N_32937);
xor U37366 (N_37366,N_33574,N_34417);
xor U37367 (N_37367,N_34456,N_34859);
nand U37368 (N_37368,N_32937,N_32612);
nor U37369 (N_37369,N_34565,N_33848);
nand U37370 (N_37370,N_32821,N_34834);
nor U37371 (N_37371,N_34802,N_32679);
and U37372 (N_37372,N_34877,N_32501);
or U37373 (N_37373,N_34268,N_33320);
xnor U37374 (N_37374,N_33484,N_34105);
nand U37375 (N_37375,N_34781,N_34092);
nand U37376 (N_37376,N_34203,N_32697);
and U37377 (N_37377,N_33323,N_33937);
or U37378 (N_37378,N_34052,N_34057);
nor U37379 (N_37379,N_34794,N_33377);
nor U37380 (N_37380,N_33294,N_33274);
xor U37381 (N_37381,N_34467,N_33405);
xnor U37382 (N_37382,N_34382,N_32972);
xor U37383 (N_37383,N_34070,N_33609);
nand U37384 (N_37384,N_32916,N_33940);
nor U37385 (N_37385,N_33924,N_34695);
or U37386 (N_37386,N_32886,N_33598);
and U37387 (N_37387,N_33889,N_32790);
and U37388 (N_37388,N_33925,N_34246);
nand U37389 (N_37389,N_33594,N_33094);
xnor U37390 (N_37390,N_34489,N_32821);
and U37391 (N_37391,N_33244,N_33235);
xor U37392 (N_37392,N_34970,N_32907);
nand U37393 (N_37393,N_34394,N_34121);
nor U37394 (N_37394,N_34969,N_33636);
and U37395 (N_37395,N_32597,N_34767);
nor U37396 (N_37396,N_33941,N_34778);
nor U37397 (N_37397,N_33286,N_32520);
nor U37398 (N_37398,N_32836,N_33806);
nor U37399 (N_37399,N_32772,N_33994);
xor U37400 (N_37400,N_34095,N_34125);
and U37401 (N_37401,N_33551,N_34933);
nand U37402 (N_37402,N_33175,N_33402);
or U37403 (N_37403,N_33405,N_33411);
nor U37404 (N_37404,N_33249,N_34563);
nor U37405 (N_37405,N_32521,N_32576);
xnor U37406 (N_37406,N_34523,N_33273);
or U37407 (N_37407,N_34187,N_33135);
nor U37408 (N_37408,N_33751,N_34264);
nor U37409 (N_37409,N_33078,N_33999);
or U37410 (N_37410,N_33755,N_34324);
or U37411 (N_37411,N_32722,N_32702);
nor U37412 (N_37412,N_32614,N_33030);
or U37413 (N_37413,N_34603,N_34775);
nand U37414 (N_37414,N_32929,N_32775);
and U37415 (N_37415,N_34926,N_32958);
nor U37416 (N_37416,N_33304,N_34971);
and U37417 (N_37417,N_33251,N_34033);
or U37418 (N_37418,N_32863,N_34579);
or U37419 (N_37419,N_34152,N_33760);
xor U37420 (N_37420,N_34305,N_34028);
and U37421 (N_37421,N_33251,N_33592);
or U37422 (N_37422,N_34082,N_32890);
or U37423 (N_37423,N_33834,N_33357);
nand U37424 (N_37424,N_32767,N_34013);
nand U37425 (N_37425,N_33230,N_33660);
and U37426 (N_37426,N_34719,N_33897);
nor U37427 (N_37427,N_34909,N_34572);
nor U37428 (N_37428,N_34147,N_34491);
xnor U37429 (N_37429,N_33842,N_32613);
nor U37430 (N_37430,N_34536,N_33227);
nand U37431 (N_37431,N_34130,N_33733);
and U37432 (N_37432,N_32864,N_32870);
nor U37433 (N_37433,N_34292,N_34155);
nand U37434 (N_37434,N_32564,N_33230);
xor U37435 (N_37435,N_32911,N_33724);
xnor U37436 (N_37436,N_32947,N_34351);
or U37437 (N_37437,N_33453,N_34666);
nor U37438 (N_37438,N_34029,N_33459);
nor U37439 (N_37439,N_34412,N_33641);
nand U37440 (N_37440,N_32636,N_34175);
or U37441 (N_37441,N_33720,N_32654);
or U37442 (N_37442,N_33752,N_34030);
and U37443 (N_37443,N_33551,N_34401);
and U37444 (N_37444,N_34954,N_32792);
or U37445 (N_37445,N_32758,N_32501);
xor U37446 (N_37446,N_33333,N_32844);
nor U37447 (N_37447,N_34320,N_33256);
and U37448 (N_37448,N_32729,N_33458);
or U37449 (N_37449,N_33407,N_34905);
nand U37450 (N_37450,N_33074,N_33322);
xor U37451 (N_37451,N_33110,N_32826);
or U37452 (N_37452,N_32856,N_34712);
and U37453 (N_37453,N_33783,N_34942);
nand U37454 (N_37454,N_32630,N_32687);
or U37455 (N_37455,N_33588,N_32620);
and U37456 (N_37456,N_33463,N_32502);
or U37457 (N_37457,N_34818,N_34912);
nand U37458 (N_37458,N_34278,N_34619);
nor U37459 (N_37459,N_32827,N_32846);
nand U37460 (N_37460,N_33487,N_33829);
xor U37461 (N_37461,N_32575,N_33723);
nor U37462 (N_37462,N_33247,N_33093);
nand U37463 (N_37463,N_34893,N_34832);
nor U37464 (N_37464,N_34082,N_33806);
xor U37465 (N_37465,N_33341,N_34183);
or U37466 (N_37466,N_33082,N_33349);
nor U37467 (N_37467,N_33299,N_34271);
nor U37468 (N_37468,N_32657,N_33546);
xor U37469 (N_37469,N_33079,N_34983);
or U37470 (N_37470,N_34992,N_34318);
xor U37471 (N_37471,N_32753,N_33283);
or U37472 (N_37472,N_33490,N_34987);
nor U37473 (N_37473,N_33214,N_34454);
xor U37474 (N_37474,N_32768,N_32575);
or U37475 (N_37475,N_33064,N_32645);
nor U37476 (N_37476,N_34464,N_32664);
xnor U37477 (N_37477,N_34874,N_33809);
nor U37478 (N_37478,N_33980,N_32859);
and U37479 (N_37479,N_33168,N_33930);
nand U37480 (N_37480,N_34444,N_34969);
nand U37481 (N_37481,N_34214,N_33526);
nand U37482 (N_37482,N_34321,N_34185);
nor U37483 (N_37483,N_34084,N_34699);
nand U37484 (N_37484,N_32992,N_34977);
nand U37485 (N_37485,N_33026,N_33731);
xnor U37486 (N_37486,N_32638,N_33916);
xor U37487 (N_37487,N_32766,N_34635);
or U37488 (N_37488,N_33005,N_33753);
nor U37489 (N_37489,N_34801,N_32658);
nand U37490 (N_37490,N_34759,N_34282);
nand U37491 (N_37491,N_32575,N_33101);
or U37492 (N_37492,N_33506,N_34225);
xnor U37493 (N_37493,N_33425,N_34449);
nand U37494 (N_37494,N_34755,N_32575);
nor U37495 (N_37495,N_34394,N_33000);
and U37496 (N_37496,N_34139,N_33339);
nor U37497 (N_37497,N_32525,N_33716);
nand U37498 (N_37498,N_33431,N_33688);
nor U37499 (N_37499,N_33990,N_34592);
nor U37500 (N_37500,N_37496,N_36249);
nor U37501 (N_37501,N_35768,N_35548);
nand U37502 (N_37502,N_36111,N_36237);
nor U37503 (N_37503,N_35975,N_35816);
xor U37504 (N_37504,N_36986,N_35019);
nand U37505 (N_37505,N_35554,N_35000);
xnor U37506 (N_37506,N_35306,N_35905);
and U37507 (N_37507,N_36978,N_35557);
or U37508 (N_37508,N_36674,N_36288);
nor U37509 (N_37509,N_35998,N_36607);
nand U37510 (N_37510,N_35967,N_37464);
nand U37511 (N_37511,N_37322,N_37288);
nand U37512 (N_37512,N_35500,N_35224);
nand U37513 (N_37513,N_37492,N_36903);
or U37514 (N_37514,N_37209,N_35239);
or U37515 (N_37515,N_36523,N_36490);
xnor U37516 (N_37516,N_35441,N_35493);
or U37517 (N_37517,N_35787,N_35217);
xor U37518 (N_37518,N_35249,N_36301);
or U37519 (N_37519,N_36478,N_35052);
and U37520 (N_37520,N_36166,N_35489);
nand U37521 (N_37521,N_36621,N_36259);
or U37522 (N_37522,N_35755,N_36026);
xnor U37523 (N_37523,N_37271,N_36744);
xnor U37524 (N_37524,N_36436,N_36873);
nor U37525 (N_37525,N_37179,N_35439);
xor U37526 (N_37526,N_35319,N_36729);
or U37527 (N_37527,N_37443,N_35640);
nand U37528 (N_37528,N_35522,N_35234);
nand U37529 (N_37529,N_35890,N_36278);
nor U37530 (N_37530,N_37174,N_35783);
nand U37531 (N_37531,N_35729,N_35564);
nand U37532 (N_37532,N_37212,N_35464);
nand U37533 (N_37533,N_37335,N_35925);
nor U37534 (N_37534,N_36118,N_35681);
xnor U37535 (N_37535,N_35386,N_36567);
and U37536 (N_37536,N_35460,N_35115);
and U37537 (N_37537,N_36002,N_36746);
nand U37538 (N_37538,N_35773,N_35305);
nand U37539 (N_37539,N_36518,N_36416);
nor U37540 (N_37540,N_36352,N_36481);
nor U37541 (N_37541,N_37205,N_36181);
nor U37542 (N_37542,N_35825,N_35374);
nor U37543 (N_37543,N_35997,N_36138);
or U37544 (N_37544,N_35670,N_35603);
nand U37545 (N_37545,N_36265,N_36940);
and U37546 (N_37546,N_36504,N_36022);
xnor U37547 (N_37547,N_35119,N_36457);
or U37548 (N_37548,N_35340,N_36546);
or U37549 (N_37549,N_37094,N_36205);
nor U37550 (N_37550,N_36686,N_35186);
nand U37551 (N_37551,N_36858,N_37272);
and U37552 (N_37552,N_36362,N_36805);
nand U37553 (N_37553,N_35085,N_36335);
nor U37554 (N_37554,N_36437,N_37059);
nand U37555 (N_37555,N_35308,N_35533);
and U37556 (N_37556,N_36829,N_35206);
nand U37557 (N_37557,N_36284,N_37268);
and U37558 (N_37558,N_36139,N_37008);
and U37559 (N_37559,N_35553,N_37308);
nand U37560 (N_37560,N_36326,N_36492);
xnor U37561 (N_37561,N_35722,N_36286);
or U37562 (N_37562,N_35760,N_35710);
and U37563 (N_37563,N_36250,N_35274);
nor U37564 (N_37564,N_37186,N_35034);
nand U37565 (N_37565,N_36705,N_35289);
xor U37566 (N_37566,N_35209,N_36754);
xnor U37567 (N_37567,N_37111,N_36402);
xnor U37568 (N_37568,N_35262,N_37331);
nor U37569 (N_37569,N_35611,N_35094);
nand U37570 (N_37570,N_36506,N_36146);
nand U37571 (N_37571,N_37064,N_36390);
xor U37572 (N_37572,N_35994,N_35245);
nand U37573 (N_37573,N_37448,N_35802);
xnor U37574 (N_37574,N_37227,N_35941);
nand U37575 (N_37575,N_35327,N_35425);
nor U37576 (N_37576,N_36882,N_35932);
nor U37577 (N_37577,N_35972,N_35738);
nand U37578 (N_37578,N_36564,N_36984);
nor U37579 (N_37579,N_36083,N_35510);
xor U37580 (N_37580,N_35951,N_36130);
or U37581 (N_37581,N_36399,N_35259);
nor U37582 (N_37582,N_35476,N_35384);
nand U37583 (N_37583,N_35665,N_36015);
xnor U37584 (N_37584,N_36602,N_36531);
xnor U37585 (N_37585,N_36660,N_35704);
nand U37586 (N_37586,N_35799,N_37267);
nand U37587 (N_37587,N_35463,N_37010);
xor U37588 (N_37588,N_35069,N_36274);
nor U37589 (N_37589,N_36944,N_37396);
and U37590 (N_37590,N_36217,N_37489);
xor U37591 (N_37591,N_35931,N_35814);
and U37592 (N_37592,N_35287,N_35562);
and U37593 (N_37593,N_35108,N_37152);
xor U37594 (N_37594,N_37126,N_36792);
or U37595 (N_37595,N_35937,N_36959);
xnor U37596 (N_37596,N_35604,N_36300);
or U37597 (N_37597,N_36615,N_36895);
nand U37598 (N_37598,N_35162,N_35201);
nor U37599 (N_37599,N_36669,N_36706);
xor U37600 (N_37600,N_37370,N_37219);
nor U37601 (N_37601,N_36779,N_36039);
nor U37602 (N_37602,N_35626,N_36807);
nand U37603 (N_37603,N_35938,N_36994);
and U37604 (N_37604,N_35839,N_35467);
or U37605 (N_37605,N_35101,N_36899);
xor U37606 (N_37606,N_37021,N_36804);
xor U37607 (N_37607,N_35283,N_36117);
xnor U37608 (N_37608,N_35494,N_36846);
and U37609 (N_37609,N_36368,N_37254);
and U37610 (N_37610,N_37098,N_37442);
xnor U37611 (N_37611,N_36195,N_36879);
xnor U37612 (N_37612,N_36939,N_35204);
nor U37613 (N_37613,N_35215,N_35674);
or U37614 (N_37614,N_36637,N_35195);
xnor U37615 (N_37615,N_35978,N_35643);
nand U37616 (N_37616,N_36539,N_36965);
xor U37617 (N_37617,N_36517,N_36623);
nor U37618 (N_37618,N_36422,N_35541);
nor U37619 (N_37619,N_35855,N_37298);
and U37620 (N_37620,N_36107,N_35586);
nand U37621 (N_37621,N_35468,N_35584);
and U37622 (N_37622,N_36868,N_36734);
xnor U37623 (N_37623,N_36737,N_37208);
nand U37624 (N_37624,N_37218,N_36787);
nor U37625 (N_37625,N_36699,N_35521);
and U37626 (N_37626,N_37201,N_35841);
xnor U37627 (N_37627,N_36296,N_37407);
or U37628 (N_37628,N_37257,N_37194);
xnor U37629 (N_37629,N_37433,N_37223);
xor U37630 (N_37630,N_36200,N_35632);
and U37631 (N_37631,N_36604,N_36397);
or U37632 (N_37632,N_36678,N_36247);
and U37633 (N_37633,N_37488,N_37099);
and U37634 (N_37634,N_37157,N_36507);
and U37635 (N_37635,N_35648,N_35082);
or U37636 (N_37636,N_37334,N_36912);
nor U37637 (N_37637,N_35796,N_36332);
or U37638 (N_37638,N_37414,N_35976);
and U37639 (N_37639,N_36781,N_35096);
nand U37640 (N_37640,N_35743,N_36204);
and U37641 (N_37641,N_36854,N_36459);
or U37642 (N_37642,N_37222,N_35326);
xnor U37643 (N_37643,N_35328,N_35285);
or U37644 (N_37644,N_37214,N_35155);
xor U37645 (N_37645,N_35711,N_37112);
and U37646 (N_37646,N_37124,N_35072);
nor U37647 (N_37647,N_36682,N_35465);
xor U37648 (N_37648,N_37460,N_36981);
xor U37649 (N_37649,N_35068,N_35291);
nor U37650 (N_37650,N_37350,N_37483);
nor U37651 (N_37651,N_35039,N_36593);
and U37652 (N_37652,N_35697,N_36442);
xnor U37653 (N_37653,N_35213,N_35872);
nand U37654 (N_37654,N_36580,N_36486);
nor U37655 (N_37655,N_37203,N_35583);
or U37656 (N_37656,N_36864,N_35636);
xor U37657 (N_37657,N_36998,N_36400);
or U37658 (N_37658,N_36659,N_35875);
and U37659 (N_37659,N_35853,N_35620);
nand U37660 (N_37660,N_37012,N_36140);
xor U37661 (N_37661,N_37360,N_35448);
nand U37662 (N_37662,N_36426,N_36095);
xor U37663 (N_37663,N_35590,N_37255);
nand U37664 (N_37664,N_35293,N_36796);
or U37665 (N_37665,N_36584,N_36281);
nand U37666 (N_37666,N_35246,N_35680);
nor U37667 (N_37667,N_35232,N_35255);
nand U37668 (N_37668,N_35982,N_37088);
or U37669 (N_37669,N_36811,N_36413);
xor U37670 (N_37670,N_37326,N_37056);
and U37671 (N_37671,N_37463,N_36215);
or U37672 (N_37672,N_35278,N_36232);
and U37673 (N_37673,N_36894,N_35803);
xor U37674 (N_37674,N_36255,N_36411);
nor U37675 (N_37675,N_36968,N_37379);
or U37676 (N_37676,N_35701,N_36641);
xnor U37677 (N_37677,N_36340,N_36740);
nor U37678 (N_37678,N_35668,N_35145);
or U37679 (N_37679,N_35296,N_37232);
xnor U37680 (N_37680,N_36155,N_36901);
or U37681 (N_37681,N_36387,N_36679);
nand U37682 (N_37682,N_36950,N_36677);
or U37683 (N_37683,N_36603,N_35402);
nor U37684 (N_37684,N_37235,N_36048);
and U37685 (N_37685,N_35826,N_35093);
xor U37686 (N_37686,N_35721,N_36435);
xnor U37687 (N_37687,N_37458,N_35807);
or U37688 (N_37688,N_36353,N_35102);
nand U37689 (N_37689,N_35926,N_36720);
or U37690 (N_37690,N_36521,N_37491);
nor U37691 (N_37691,N_36810,N_35970);
or U37692 (N_37692,N_37459,N_35824);
and U37693 (N_37693,N_35180,N_36407);
nor U37694 (N_37694,N_36318,N_35786);
or U37695 (N_37695,N_35672,N_36363);
and U37696 (N_37696,N_35687,N_35200);
nand U37697 (N_37697,N_35227,N_35619);
nor U37698 (N_37698,N_35138,N_37180);
and U37699 (N_37699,N_35651,N_35910);
nor U37700 (N_37700,N_37085,N_35950);
or U37701 (N_37701,N_35149,N_36624);
nor U37702 (N_37702,N_35889,N_36150);
xnor U37703 (N_37703,N_35833,N_37382);
or U37704 (N_37704,N_36384,N_36925);
nor U37705 (N_37705,N_35673,N_36474);
and U37706 (N_37706,N_37402,N_36548);
or U37707 (N_37707,N_35112,N_36020);
or U37708 (N_37708,N_35746,N_37013);
xnor U37709 (N_37709,N_37487,N_36691);
xnor U37710 (N_37710,N_36410,N_36820);
or U37711 (N_37711,N_36105,N_36742);
and U37712 (N_37712,N_36997,N_36631);
and U37713 (N_37713,N_36844,N_37340);
and U37714 (N_37714,N_35018,N_36446);
nor U37715 (N_37715,N_36601,N_36109);
and U37716 (N_37716,N_36099,N_37125);
or U37717 (N_37717,N_36738,N_35633);
and U37718 (N_37718,N_36656,N_35136);
or U37719 (N_37719,N_36769,N_35003);
and U37720 (N_37720,N_36955,N_36424);
nand U37721 (N_37721,N_36739,N_35405);
xor U37722 (N_37722,N_35295,N_35453);
and U37723 (N_37723,N_36954,N_36665);
nand U37724 (N_37724,N_35426,N_36951);
xor U37725 (N_37725,N_36916,N_36645);
nand U37726 (N_37726,N_35081,N_36075);
and U37727 (N_37727,N_35895,N_36917);
and U37728 (N_37728,N_36159,N_37033);
or U37729 (N_37729,N_36432,N_36135);
nand U37730 (N_37730,N_35505,N_37310);
or U37731 (N_37731,N_36927,N_36524);
or U37732 (N_37732,N_36772,N_37348);
nor U37733 (N_37733,N_37327,N_36224);
or U37734 (N_37734,N_35432,N_37357);
or U37735 (N_37735,N_36897,N_36412);
xnor U37736 (N_37736,N_35264,N_36240);
nand U37737 (N_37737,N_36789,N_37371);
and U37738 (N_37738,N_37049,N_36559);
and U37739 (N_37739,N_35689,N_36822);
nor U37740 (N_37740,N_35258,N_36845);
nand U37741 (N_37741,N_36110,N_35908);
nand U37742 (N_37742,N_36186,N_36377);
xnor U37743 (N_37743,N_35776,N_35912);
or U37744 (N_37744,N_36608,N_36651);
or U37745 (N_37745,N_36067,N_35471);
xor U37746 (N_37746,N_36272,N_35116);
nand U37747 (N_37747,N_36134,N_36439);
or U37748 (N_37748,N_36992,N_35804);
and U37749 (N_37749,N_36694,N_36719);
xnor U37750 (N_37750,N_35190,N_36800);
nand U37751 (N_37751,N_36444,N_35167);
nand U37752 (N_37752,N_37103,N_35621);
nand U37753 (N_37753,N_35860,N_37373);
xnor U37754 (N_37754,N_36017,N_36576);
nor U37755 (N_37755,N_35172,N_35806);
nor U37756 (N_37756,N_37044,N_35161);
and U37757 (N_37757,N_36733,N_35133);
nor U37758 (N_37758,N_36736,N_36730);
and U37759 (N_37759,N_35867,N_36196);
or U37760 (N_37760,N_36834,N_37072);
xor U37761 (N_37761,N_35380,N_35131);
xor U37762 (N_37762,N_35748,N_35605);
nand U37763 (N_37763,N_35399,N_36023);
nand U37764 (N_37764,N_36308,N_36752);
xor U37765 (N_37765,N_35477,N_35488);
nor U37766 (N_37766,N_35430,N_36935);
nand U37767 (N_37767,N_36154,N_35304);
nand U37768 (N_37768,N_35171,N_36741);
or U37769 (N_37769,N_35040,N_35914);
or U37770 (N_37770,N_35623,N_37333);
and U37771 (N_37771,N_37274,N_36386);
nor U37772 (N_37772,N_37145,N_35515);
nand U37773 (N_37773,N_37282,N_36497);
nand U37774 (N_37774,N_36261,N_36409);
and U37775 (N_37775,N_35222,N_35442);
nand U37776 (N_37776,N_36883,N_36188);
xnor U37777 (N_37777,N_37493,N_36723);
xor U37778 (N_37778,N_36070,N_35717);
or U37779 (N_37779,N_35595,N_35363);
or U37780 (N_37780,N_35892,N_35745);
xnor U37781 (N_37781,N_36589,N_36922);
nand U37782 (N_37782,N_35501,N_36743);
nor U37783 (N_37783,N_35986,N_35290);
or U37784 (N_37784,N_36192,N_35723);
and U37785 (N_37785,N_37106,N_35598);
nor U37786 (N_37786,N_35028,N_36010);
nor U37787 (N_37787,N_35742,N_36536);
xor U37788 (N_37788,N_35736,N_35236);
or U37789 (N_37789,N_37116,N_36859);
or U37790 (N_37790,N_36086,N_35545);
nor U37791 (N_37791,N_36722,N_36228);
nor U37792 (N_37792,N_36392,N_37473);
xor U37793 (N_37793,N_35381,N_35820);
xnor U37794 (N_37794,N_37262,N_35434);
xnor U37795 (N_37795,N_36221,N_35411);
or U37796 (N_37796,N_35220,N_36141);
nor U37797 (N_37797,N_35568,N_36183);
nor U37798 (N_37798,N_35791,N_35303);
nand U37799 (N_37799,N_37482,N_37143);
nand U37800 (N_37800,N_36482,N_35177);
nand U37801 (N_37801,N_37184,N_35563);
xnor U37802 (N_37802,N_36838,N_37418);
or U37803 (N_37803,N_35531,N_35832);
and U37804 (N_37804,N_35676,N_36885);
xnor U37805 (N_37805,N_35342,N_36690);
xor U37806 (N_37806,N_36891,N_37095);
nand U37807 (N_37807,N_36463,N_37265);
and U37808 (N_37808,N_35995,N_35005);
nor U37809 (N_37809,N_35141,N_35387);
nor U37810 (N_37810,N_35606,N_35764);
nor U37811 (N_37811,N_36967,N_35961);
and U37812 (N_37812,N_36191,N_36069);
xor U37813 (N_37813,N_35030,N_35397);
nand U37814 (N_37814,N_36330,N_36214);
xnor U37815 (N_37815,N_35840,N_35341);
nand U37816 (N_37816,N_37189,N_37229);
nand U37817 (N_37817,N_36571,N_36535);
nor U37818 (N_37818,N_37449,N_37122);
xor U37819 (N_37819,N_35747,N_36003);
or U37820 (N_37820,N_36000,N_35608);
xor U37821 (N_37821,N_36904,N_36013);
and U37822 (N_37822,N_36465,N_35933);
nor U37823 (N_37823,N_36197,N_35631);
nor U37824 (N_37824,N_36600,N_35237);
nand U37825 (N_37825,N_35302,N_35404);
or U37826 (N_37826,N_36294,N_37197);
xor U37827 (N_37827,N_37119,N_35659);
nor U37828 (N_37828,N_37381,N_35029);
and U37829 (N_37829,N_37062,N_37450);
and U37830 (N_37830,N_36709,N_35315);
nor U37831 (N_37831,N_36454,N_35944);
xnor U37832 (N_37832,N_35197,N_36434);
and U37833 (N_37833,N_35045,N_36458);
nor U37834 (N_37834,N_35990,N_36848);
xor U37835 (N_37835,N_35428,N_35777);
xor U37836 (N_37836,N_35076,N_36046);
nor U37837 (N_37837,N_36452,N_35412);
nor U37838 (N_37838,N_35333,N_37244);
and U37839 (N_37839,N_37127,N_35491);
or U37840 (N_37840,N_37477,N_35187);
nand U37841 (N_37841,N_35216,N_37250);
nand U37842 (N_37842,N_35396,N_36327);
or U37843 (N_37843,N_37387,N_35312);
and U37844 (N_37844,N_37071,N_37213);
nand U37845 (N_37845,N_36703,N_37380);
nand U37846 (N_37846,N_35055,N_35298);
and U37847 (N_37847,N_36563,N_36761);
nor U37848 (N_37848,N_35241,N_36053);
or U37849 (N_37849,N_35727,N_36648);
and U37850 (N_37850,N_36448,N_37037);
and U37851 (N_37851,N_35750,N_37048);
xor U37852 (N_37852,N_35856,N_36666);
nor U37853 (N_37853,N_37343,N_35366);
and U37854 (N_37854,N_36892,N_36290);
and U37855 (N_37855,N_35146,N_36587);
or U37856 (N_37856,N_37299,N_35886);
or U37857 (N_37857,N_35212,N_37234);
and U37858 (N_37858,N_36812,N_36136);
or U37859 (N_37859,N_35225,N_35939);
and U37860 (N_37860,N_36728,N_35725);
nand U37861 (N_37861,N_35771,N_35592);
xnor U37862 (N_37862,N_35269,N_35898);
nand U37863 (N_37863,N_36835,N_35999);
nand U37864 (N_37864,N_37353,N_36661);
nand U37865 (N_37865,N_35831,N_37083);
and U37866 (N_37866,N_35165,N_35079);
or U37867 (N_37867,N_37027,N_36170);
xor U37868 (N_37868,N_35379,N_36760);
nand U37869 (N_37869,N_36203,N_36842);
nor U37870 (N_37870,N_35752,N_37165);
and U37871 (N_37871,N_35194,N_36374);
nand U37872 (N_37872,N_35140,N_36008);
and U37873 (N_37873,N_35210,N_35123);
nor U37874 (N_37874,N_36404,N_36151);
or U37875 (N_37875,N_37225,N_35472);
and U37876 (N_37876,N_36907,N_36208);
and U37877 (N_37877,N_36716,N_35885);
and U37878 (N_37878,N_35694,N_37046);
xnor U37879 (N_37879,N_35547,N_36317);
xor U37880 (N_37880,N_37242,N_36189);
or U37881 (N_37881,N_37276,N_36642);
or U37882 (N_37882,N_35654,N_35125);
xor U37883 (N_37883,N_36532,N_36244);
nand U37884 (N_37884,N_37080,N_35556);
xor U37885 (N_37885,N_36906,N_36216);
nor U37886 (N_37886,N_36771,N_35208);
or U37887 (N_37887,N_35569,N_36647);
and U37888 (N_37888,N_35642,N_37376);
nand U37889 (N_37889,N_35969,N_35966);
and U37890 (N_37890,N_35699,N_35487);
xor U37891 (N_37891,N_37063,N_36933);
nand U37892 (N_37892,N_35486,N_35709);
or U37893 (N_37893,N_35946,N_35953);
and U37894 (N_37894,N_37199,N_36630);
nand U37895 (N_37895,N_35575,N_35767);
xnor U37896 (N_37896,N_36227,N_36996);
or U37897 (N_37897,N_35974,N_35713);
nor U37898 (N_37898,N_37023,N_35202);
and U37899 (N_37899,N_37097,N_36103);
nand U37900 (N_37900,N_35257,N_35135);
nand U37901 (N_37901,N_35139,N_36349);
nand U37902 (N_37902,N_36878,N_35887);
or U37903 (N_37903,N_36322,N_35148);
and U37904 (N_37904,N_36391,N_36824);
nor U37905 (N_37905,N_36610,N_36383);
and U37906 (N_37906,N_36094,N_36639);
xor U37907 (N_37907,N_36757,N_36849);
xor U37908 (N_37908,N_37216,N_35027);
nand U37909 (N_37909,N_35002,N_36114);
and U37910 (N_37910,N_36263,N_35421);
and U37911 (N_37911,N_36865,N_37035);
nand U37912 (N_37912,N_35331,N_36484);
or U37913 (N_37913,N_36818,N_36886);
and U37914 (N_37914,N_37009,N_36928);
nand U37915 (N_37915,N_35958,N_35936);
nor U37916 (N_37916,N_36670,N_36974);
xor U37917 (N_37917,N_36125,N_35025);
or U37918 (N_37918,N_35830,N_35026);
and U37919 (N_37919,N_37193,N_36074);
and U37920 (N_37920,N_35928,N_36606);
nand U37921 (N_37921,N_36766,N_35391);
nor U37922 (N_37922,N_36050,N_37055);
and U37923 (N_37923,N_35706,N_37025);
nor U37924 (N_37924,N_35378,N_35074);
and U37925 (N_37925,N_37345,N_37332);
nand U37926 (N_37926,N_36543,N_36596);
or U37927 (N_37927,N_37156,N_37260);
xnor U37928 (N_37928,N_35567,N_37153);
xor U37929 (N_37929,N_36793,N_36293);
or U37930 (N_37930,N_37256,N_37398);
or U37931 (N_37931,N_35024,N_35001);
xnor U37932 (N_37932,N_36202,N_35716);
xnor U37933 (N_37933,N_36063,N_36096);
xnor U37934 (N_37934,N_36356,N_37224);
or U37935 (N_37935,N_36934,N_37317);
nor U37936 (N_37936,N_36776,N_37040);
nand U37937 (N_37937,N_35991,N_35032);
nand U37938 (N_37938,N_37129,N_35354);
and U37939 (N_37939,N_36887,N_35438);
xnor U37940 (N_37940,N_36080,N_37200);
nand U37941 (N_37941,N_35517,N_37454);
and U37942 (N_37942,N_35666,N_35900);
nand U37943 (N_37943,N_36176,N_37211);
and U37944 (N_37944,N_36488,N_37365);
nand U37945 (N_37945,N_36747,N_37470);
xor U37946 (N_37946,N_36632,N_36866);
xnor U37947 (N_37947,N_37230,N_36342);
nand U37948 (N_37948,N_36305,N_36541);
nand U37949 (N_37949,N_35451,N_35169);
xnor U37950 (N_37950,N_37022,N_35347);
nand U37951 (N_37951,N_35252,N_35573);
xnor U37952 (N_37952,N_35006,N_35693);
and U37953 (N_37953,N_35016,N_35552);
xnor U37954 (N_37954,N_35506,N_36473);
nand U37955 (N_37955,N_36408,N_36280);
or U37956 (N_37956,N_37485,N_37187);
nand U37957 (N_37957,N_37196,N_37384);
nand U37958 (N_37958,N_35981,N_37057);
nor U37959 (N_37959,N_36282,N_35250);
xnor U37960 (N_37960,N_36334,N_36267);
xnor U37961 (N_37961,N_36311,N_36403);
nor U37962 (N_37962,N_36447,N_37270);
and U37963 (N_37963,N_37385,N_36929);
nor U37964 (N_37964,N_35033,N_36262);
nor U37965 (N_37965,N_36756,N_35427);
or U37966 (N_37966,N_36554,N_35737);
and U37967 (N_37967,N_35330,N_37302);
or U37968 (N_37968,N_35546,N_36643);
xnor U37969 (N_37969,N_35514,N_36428);
nor U37970 (N_37970,N_36037,N_35530);
nor U37971 (N_37971,N_36087,N_37413);
xnor U37972 (N_37972,N_35795,N_36019);
and U37973 (N_37973,N_35821,N_36801);
or U37974 (N_37974,N_35770,N_37294);
and U37975 (N_37975,N_36084,N_37425);
xnor U37976 (N_37976,N_37053,N_36235);
xor U37977 (N_37977,N_36876,N_36908);
or U37978 (N_37978,N_36758,N_36178);
and U37979 (N_37979,N_37002,N_36931);
nand U37980 (N_37980,N_36027,N_36668);
nand U37981 (N_37981,N_37362,N_35857);
nand U37982 (N_37982,N_36863,N_37195);
nand U37983 (N_37983,N_36123,N_36085);
and U37984 (N_37984,N_35062,N_36045);
and U37985 (N_37985,N_36382,N_36809);
and U37986 (N_37986,N_36595,N_36106);
xnor U37987 (N_37987,N_37364,N_36348);
or U37988 (N_37988,N_36370,N_35192);
and U37989 (N_37989,N_37176,N_36120);
and U37990 (N_37990,N_37281,N_36585);
nor U37991 (N_37991,N_36076,N_36609);
and U37992 (N_37992,N_36806,N_37206);
nand U37993 (N_37993,N_35398,N_35454);
nand U37994 (N_37994,N_37436,N_36827);
or U37995 (N_37995,N_37006,N_37163);
nand U37996 (N_37996,N_36129,N_37043);
and U37997 (N_37997,N_37139,N_35863);
xnor U37998 (N_37998,N_35596,N_36636);
nand U37999 (N_37999,N_35248,N_35372);
and U38000 (N_38000,N_35406,N_37160);
nand U38001 (N_38001,N_35587,N_35324);
or U38002 (N_38002,N_35789,N_36770);
and U38003 (N_38003,N_36896,N_36773);
and U38004 (N_38004,N_35475,N_35849);
or U38005 (N_38005,N_35763,N_37007);
nor U38006 (N_38006,N_35544,N_36116);
and U38007 (N_38007,N_35351,N_36358);
and U38008 (N_38008,N_36206,N_35338);
nand U38009 (N_38009,N_37166,N_36018);
xnor U38010 (N_38010,N_35637,N_35943);
xnor U38011 (N_38011,N_35408,N_35686);
or U38012 (N_38012,N_35124,N_35504);
xnor U38013 (N_38013,N_35616,N_37476);
nor U38014 (N_38014,N_37456,N_35979);
nor U38015 (N_38015,N_36881,N_35678);
or U38016 (N_38016,N_35915,N_35602);
xnor U38017 (N_38017,N_36920,N_36969);
or U38018 (N_38018,N_36574,N_35004);
nor U38019 (N_38019,N_36266,N_35403);
nand U38020 (N_38020,N_35349,N_36938);
and U38021 (N_38021,N_37231,N_35419);
or U38022 (N_38022,N_36629,N_35909);
nand U38023 (N_38023,N_36350,N_37484);
nor U38024 (N_38024,N_36791,N_37393);
xor U38025 (N_38025,N_36419,N_35088);
and U38026 (N_38026,N_36777,N_36292);
and U38027 (N_38027,N_35513,N_36544);
nor U38028 (N_38028,N_36376,N_35253);
xor U38029 (N_38029,N_35535,N_35624);
or U38030 (N_38030,N_36952,N_35479);
nand U38031 (N_38031,N_35866,N_35658);
xor U38032 (N_38032,N_35320,N_35732);
and U38033 (N_38033,N_35843,N_36652);
nand U38034 (N_38034,N_35221,N_37445);
nand U38035 (N_38035,N_35566,N_35435);
nor U38036 (N_38036,N_35525,N_35041);
and U38037 (N_38037,N_36364,N_36983);
or U38038 (N_38038,N_35189,N_35675);
nand U38039 (N_38039,N_36790,N_36471);
nand U38040 (N_38040,N_35766,N_36926);
xor U38041 (N_38041,N_37494,N_35474);
nor U38042 (N_38042,N_37421,N_35509);
and U38043 (N_38043,N_35357,N_35720);
nor U38044 (N_38044,N_35835,N_36689);
nand U38045 (N_38045,N_35641,N_35854);
nor U38046 (N_38046,N_35645,N_36487);
or U38047 (N_38047,N_35228,N_36852);
or U38048 (N_38048,N_36681,N_35873);
nor U38049 (N_38049,N_36993,N_37427);
and U38050 (N_38050,N_36001,N_35878);
or U38051 (N_38051,N_37319,N_37401);
xor U38052 (N_38052,N_36683,N_35382);
nor U38053 (N_38053,N_36143,N_36222);
nor U38054 (N_38054,N_36461,N_35907);
xnor U38055 (N_38055,N_35884,N_35497);
nor U38056 (N_38056,N_36970,N_37457);
or U38057 (N_38057,N_35218,N_35980);
xnor U38058 (N_38058,N_37123,N_37301);
or U38059 (N_38059,N_36612,N_36236);
nor U38060 (N_38060,N_36401,N_36287);
or U38061 (N_38061,N_35917,N_37296);
nand U38062 (N_38062,N_35507,N_36367);
nand U38063 (N_38063,N_36855,N_35173);
and U38064 (N_38064,N_35698,N_37161);
nor U38065 (N_38065,N_36870,N_37204);
and U38066 (N_38066,N_35238,N_35150);
xor U38067 (N_38067,N_36165,N_37344);
or U38068 (N_38068,N_35811,N_36638);
xor U38069 (N_38069,N_37029,N_35580);
nor U38070 (N_38070,N_35576,N_36102);
or U38071 (N_38071,N_36260,N_35930);
xnor U38072 (N_38072,N_36121,N_35762);
xnor U38073 (N_38073,N_36128,N_35417);
nand U38074 (N_38074,N_36242,N_35483);
nor U38075 (N_38075,N_37453,N_35056);
xnor U38076 (N_38076,N_35663,N_36514);
nor U38077 (N_38077,N_36888,N_35176);
and U38078 (N_38078,N_36936,N_36774);
and U38079 (N_38079,N_36628,N_37293);
and U38080 (N_38080,N_36527,N_36957);
nand U38081 (N_38081,N_35700,N_36275);
or U38082 (N_38082,N_36126,N_35695);
xnor U38083 (N_38083,N_35277,N_36451);
xor U38084 (N_38084,N_35896,N_35231);
xnor U38085 (N_38085,N_36007,N_35271);
xor U38086 (N_38086,N_36088,N_35057);
or U38087 (N_38087,N_35667,N_35809);
nor U38088 (N_38088,N_36066,N_37202);
nand U38089 (N_38089,N_35865,N_36988);
nand U38090 (N_38090,N_35682,N_37409);
xnor U38091 (N_38091,N_35549,N_36579);
nand U38092 (N_38092,N_36243,N_37278);
or U38093 (N_38093,N_37415,N_37304);
or U38094 (N_38094,N_37283,N_35929);
or U38095 (N_38095,N_36470,N_37297);
xor U38096 (N_38096,N_35949,N_36753);
or U38097 (N_38097,N_35539,N_35375);
or U38098 (N_38098,N_36064,N_35394);
and U38099 (N_38099,N_35368,N_37287);
xor U38100 (N_38100,N_36594,N_37366);
nor U38101 (N_38101,N_35733,N_36592);
or U38102 (N_38102,N_36059,N_36707);
or U38103 (N_38103,N_35235,N_36839);
xnor U38104 (N_38104,N_35871,N_35174);
and U38105 (N_38105,N_36687,N_35266);
nand U38106 (N_38106,N_35600,N_36372);
xor U38107 (N_38107,N_35134,N_36826);
nor U38108 (N_38108,N_36815,N_36646);
nor U38109 (N_38109,N_36483,N_37091);
nor U38110 (N_38110,N_36101,N_35661);
nor U38111 (N_38111,N_36538,N_36418);
and U38112 (N_38112,N_35317,N_35449);
nor U38113 (N_38113,N_35367,N_36953);
nand U38114 (N_38114,N_37423,N_36254);
xor U38115 (N_38115,N_35012,N_37076);
and U38116 (N_38116,N_35143,N_37431);
or U38117 (N_38117,N_35356,N_37068);
nand U38118 (N_38118,N_35407,N_36172);
xnor U38119 (N_38119,N_35389,N_36314);
or U38120 (N_38120,N_36464,N_35325);
nor U38121 (N_38121,N_36338,N_36175);
or U38122 (N_38122,N_37104,N_37164);
and U38123 (N_38123,N_35793,N_37236);
xnor U38124 (N_38124,N_35061,N_36561);
and U38125 (N_38125,N_36241,N_35744);
xor U38126 (N_38126,N_37383,N_36995);
and U38127 (N_38127,N_36378,N_37003);
or U38128 (N_38128,N_35188,N_37065);
xor U38129 (N_38129,N_35316,N_35690);
nor U38130 (N_38130,N_36914,N_36547);
or U38131 (N_38131,N_35498,N_35207);
xor U38132 (N_38132,N_35343,N_35309);
nand U38133 (N_38133,N_36077,N_37252);
and U38134 (N_38134,N_36566,N_36964);
xor U38135 (N_38135,N_36861,N_35132);
or U38136 (N_38136,N_36583,N_37183);
nand U38137 (N_38137,N_36655,N_35550);
xor U38138 (N_38138,N_37277,N_36044);
nand U38139 (N_38139,N_36999,N_36313);
nand U38140 (N_38140,N_35650,N_35741);
xor U38141 (N_38141,N_36910,N_35617);
or U38142 (N_38142,N_36441,N_37079);
nor U38143 (N_38143,N_35753,N_37279);
nand U38144 (N_38144,N_37391,N_37318);
nand U38145 (N_38145,N_35036,N_36526);
nand U38146 (N_38146,N_36732,N_37378);
or U38147 (N_38147,N_35612,N_36725);
nor U38148 (N_38148,N_35754,N_35899);
xnor U38149 (N_38149,N_35392,N_36230);
nor U38150 (N_38150,N_35916,N_35555);
xnor U38151 (N_38151,N_36704,N_37311);
or U38152 (N_38152,N_36918,N_36671);
nand U38153 (N_38153,N_36012,N_35339);
and U38154 (N_38154,N_35655,N_35536);
or U38155 (N_38155,N_36032,N_37110);
or U38156 (N_38156,N_37352,N_37226);
nor U38157 (N_38157,N_36598,N_36341);
nand U38158 (N_38158,N_35263,N_37490);
xor U38159 (N_38159,N_36331,N_35964);
xnor U38160 (N_38160,N_35757,N_36345);
xor U38161 (N_38161,N_37320,N_36745);
nor U38162 (N_38162,N_36160,N_35719);
xor U38163 (N_38163,N_36971,N_35395);
nand U38164 (N_38164,N_35869,N_37359);
nand U38165 (N_38165,N_36911,N_36718);
nor U38166 (N_38166,N_35838,N_35254);
nor U38167 (N_38167,N_35481,N_36194);
xnor U38168 (N_38168,N_37042,N_35798);
or U38169 (N_38169,N_35073,N_36626);
xnor U38170 (N_38170,N_37439,N_35561);
nand U38171 (N_38171,N_36218,N_36238);
nor U38172 (N_38172,N_35223,N_35075);
or U38173 (N_38173,N_36025,N_36147);
nand U38174 (N_38174,N_35084,N_37486);
nand U38175 (N_38175,N_35708,N_37135);
or U38176 (N_38176,N_37130,N_37093);
nand U38177 (N_38177,N_35850,N_37404);
or U38178 (N_38178,N_37465,N_36856);
and U38179 (N_38179,N_36127,N_35362);
nor U38180 (N_38180,N_36289,N_35307);
nor U38181 (N_38181,N_37285,N_35524);
and U38182 (N_38182,N_37167,N_36054);
or U38183 (N_38183,N_36450,N_36057);
xnor U38184 (N_38184,N_35265,N_35952);
and U38185 (N_38185,N_35461,N_37475);
xor U38186 (N_38186,N_35518,N_35823);
nand U38187 (N_38187,N_37480,N_37084);
xnor U38188 (N_38188,N_35336,N_35103);
nand U38189 (N_38189,N_36058,N_37253);
and U38190 (N_38190,N_36445,N_35170);
xor U38191 (N_38191,N_35610,N_35657);
nor U38192 (N_38192,N_35211,N_36987);
or U38193 (N_38193,N_35240,N_37141);
nand U38194 (N_38194,N_35859,N_35098);
nor U38195 (N_38195,N_35182,N_36947);
and U38196 (N_38196,N_36041,N_36542);
nand U38197 (N_38197,N_36190,N_35009);
xnor U38198 (N_38198,N_35469,N_35870);
and U38199 (N_38199,N_37032,N_36717);
xor U38200 (N_38200,N_36803,N_36937);
and U38201 (N_38201,N_35519,N_37246);
nand U38202 (N_38202,N_37498,N_37158);
nor U38203 (N_38203,N_36271,N_36062);
and U38204 (N_38204,N_36201,N_35913);
nor U38205 (N_38205,N_37309,N_35836);
xor U38206 (N_38206,N_36466,N_36385);
nand U38207 (N_38207,N_35321,N_35348);
nand U38208 (N_38208,N_36537,N_35893);
nand U38209 (N_38209,N_37389,N_35163);
nand U38210 (N_38210,N_36344,N_36562);
xnor U38211 (N_38211,N_35268,N_37051);
nand U38212 (N_38212,N_36328,N_37307);
and U38213 (N_38213,N_36220,N_36872);
nand U38214 (N_38214,N_36347,N_35989);
nand U38215 (N_38215,N_35364,N_36590);
nand U38216 (N_38216,N_36239,N_35297);
and U38217 (N_38217,N_36823,N_35198);
or U38218 (N_38218,N_36476,N_36510);
xnor U38219 (N_38219,N_36869,N_35627);
or U38220 (N_38220,N_35542,N_35543);
nor U38221 (N_38221,N_36821,N_36676);
nand U38222 (N_38222,N_36389,N_35647);
and U38223 (N_38223,N_36591,N_36209);
and U38224 (N_38224,N_37146,N_36989);
nand U38225 (N_38225,N_36991,N_35848);
and U38226 (N_38226,N_36393,N_35778);
xor U38227 (N_38227,N_35118,N_36520);
and U38228 (N_38228,N_36680,N_37109);
nand U38229 (N_38229,N_37263,N_36700);
nand U38230 (N_38230,N_35275,N_36479);
xnor U38231 (N_38231,N_36775,N_35021);
xnor U38232 (N_38232,N_35099,N_37437);
nand U38233 (N_38233,N_36078,N_36082);
xnor U38234 (N_38234,N_36831,N_36167);
nand U38235 (N_38235,N_35156,N_37411);
and U38236 (N_38236,N_35677,N_35609);
xnor U38237 (N_38237,N_37147,N_35436);
and U38238 (N_38238,N_35314,N_35388);
or U38239 (N_38239,N_35080,N_35361);
nand U38240 (N_38240,N_36113,N_35323);
nand U38241 (N_38241,N_36455,N_36945);
nand U38242 (N_38242,N_36494,N_36814);
xnor U38243 (N_38243,N_35058,N_36093);
nor U38244 (N_38244,N_35644,N_35921);
nor U38245 (N_38245,N_36213,N_37451);
or U38246 (N_38246,N_37169,N_36297);
nor U38247 (N_38247,N_36702,N_35815);
nand U38248 (N_38248,N_35983,N_36371);
or U38249 (N_38249,N_37447,N_36550);
xor U38250 (N_38250,N_35183,N_36560);
xor U38251 (N_38251,N_36816,N_36068);
and U38252 (N_38252,N_35817,N_36357);
or U38253 (N_38253,N_36724,N_36168);
or U38254 (N_38254,N_36004,N_35558);
nor U38255 (N_38255,N_35199,N_35782);
and U38256 (N_38256,N_37324,N_36540);
or U38257 (N_38257,N_35581,N_36778);
or U38258 (N_38258,N_35154,N_37392);
xor U38259 (N_38259,N_36420,N_35496);
nor U38260 (N_38260,N_36030,N_35560);
nor U38261 (N_38261,N_35511,N_36749);
nand U38262 (N_38262,N_36708,N_36851);
or U38263 (N_38263,N_36588,N_36599);
nand U38264 (N_38264,N_36198,N_36475);
or U38265 (N_38265,N_37400,N_37172);
xnor U38266 (N_38266,N_36875,N_37354);
and U38267 (N_38267,N_35462,N_36233);
nand U38268 (N_38268,N_35409,N_35168);
or U38269 (N_38269,N_36611,N_35400);
or U38270 (N_38270,N_35774,N_37269);
or U38271 (N_38271,N_35691,N_35819);
and U38272 (N_38272,N_36443,N_37245);
nor U38273 (N_38273,N_35484,N_35385);
xnor U38274 (N_38274,N_36161,N_35346);
nor U38275 (N_38275,N_36505,N_35470);
and U38276 (N_38276,N_36137,N_37154);
and U38277 (N_38277,N_36351,N_35064);
nand U38278 (N_38278,N_35178,N_36512);
or U38279 (N_38279,N_36038,N_37441);
or U38280 (N_38280,N_36759,N_36693);
and U38281 (N_38281,N_36529,N_36649);
or U38282 (N_38282,N_36162,N_37394);
nor U38283 (N_38283,N_37036,N_36379);
nand U38284 (N_38284,N_37058,N_36813);
and U38285 (N_38285,N_36456,N_35358);
xnor U38286 (N_38286,N_36616,N_37170);
or U38287 (N_38287,N_35107,N_37117);
nor U38288 (N_38288,N_35715,N_35864);
or U38289 (N_38289,N_35646,N_36575);
xnor U38290 (N_38290,N_36223,N_36158);
or U38291 (N_38291,N_35047,N_35726);
nand U38292 (N_38292,N_35284,N_36277);
xor U38293 (N_38293,N_36193,N_35512);
or U38294 (N_38294,N_37372,N_37039);
nand U38295 (N_38295,N_37248,N_37323);
nor U38296 (N_38296,N_36860,N_37495);
nor U38297 (N_38297,N_37406,N_37466);
xnor U38298 (N_38298,N_36765,N_35273);
and U38299 (N_38299,N_36199,N_37120);
nor U38300 (N_38300,N_35355,N_35046);
nor U38301 (N_38301,N_36684,N_37177);
nand U38302 (N_38302,N_36902,N_35490);
or U38303 (N_38303,N_37300,N_36605);
and U38304 (N_38304,N_36555,N_36306);
nand U38305 (N_38305,N_36692,N_36572);
and U38306 (N_38306,N_35193,N_36453);
nand U38307 (N_38307,N_35585,N_35401);
or U38308 (N_38308,N_36315,N_36782);
and U38309 (N_38309,N_36415,N_37247);
nor U38310 (N_38310,N_36100,N_36909);
or U38311 (N_38311,N_35157,N_37136);
nor U38312 (N_38312,N_35260,N_37171);
nor U38313 (N_38313,N_37090,N_35444);
and U38314 (N_38314,N_35851,N_35794);
nand U38315 (N_38315,N_36047,N_35756);
nand U38316 (N_38316,N_35551,N_35153);
nand U38317 (N_38317,N_36179,N_37243);
and U38318 (N_38318,N_35054,N_36697);
xnor U38319 (N_38319,N_36979,N_35114);
xor U38320 (N_38320,N_35482,N_35344);
xor U38321 (N_38321,N_37266,N_36319);
nor U38322 (N_38322,N_37258,N_35993);
or U38323 (N_38323,N_36956,N_35294);
or U38324 (N_38324,N_35458,N_36874);
and U38325 (N_38325,N_35089,N_37198);
xor U38326 (N_38326,N_35455,N_37325);
xnor U38327 (N_38327,N_37089,N_36405);
or U38328 (N_38328,N_35130,N_36480);
and U38329 (N_38329,N_37306,N_36712);
nand U38330 (N_38330,N_37070,N_35111);
xnor U38331 (N_38331,N_36496,N_36304);
or U38332 (N_38332,N_37292,N_36090);
nand U38333 (N_38333,N_36884,N_35888);
or U38334 (N_38334,N_35718,N_36229);
or U38335 (N_38335,N_37026,N_37468);
xnor U38336 (N_38336,N_36534,N_36156);
and U38337 (N_38337,N_36152,N_36614);
nor U38338 (N_38338,N_35393,N_35311);
or U38339 (N_38339,N_36688,N_35159);
nor U38340 (N_38340,N_37312,N_36283);
and U38341 (N_38341,N_35142,N_35662);
xor U38342 (N_38342,N_36169,N_35653);
nor U38343 (N_38343,N_37397,N_36508);
xnor U38344 (N_38344,N_36963,N_35414);
nand U38345 (N_38345,N_37367,N_37430);
and U38346 (N_38346,N_36354,N_35582);
xnor U38347 (N_38347,N_37429,N_35920);
nor U38348 (N_38348,N_36921,N_37069);
and U38349 (N_38349,N_37497,N_36731);
nand U38350 (N_38350,N_35988,N_35613);
or U38351 (N_38351,N_36253,N_36568);
nand U38352 (N_38352,N_35485,N_36366);
and U38353 (N_38353,N_36091,N_35158);
xor U38354 (N_38354,N_36079,N_36569);
nand U38355 (N_38355,N_35818,N_37017);
or U38356 (N_38356,N_36635,N_37041);
xor U38357 (N_38357,N_36667,N_36960);
nor U38358 (N_38358,N_37128,N_35911);
nor U38359 (N_38359,N_36962,N_35352);
nor U38360 (N_38360,N_35031,N_36701);
nand U38361 (N_38361,N_35985,N_37005);
or U38362 (N_38362,N_35973,N_35160);
or U38363 (N_38363,N_35957,N_35127);
or U38364 (N_38364,N_37001,N_37233);
nand U38365 (N_38365,N_36619,N_35313);
or U38366 (N_38366,N_36880,N_36977);
or U38367 (N_38367,N_36395,N_37355);
nand U38368 (N_38368,N_35322,N_37356);
nand U38369 (N_38369,N_35365,N_37024);
or U38370 (N_38370,N_35113,N_36381);
and U38371 (N_38371,N_35904,N_35203);
or U38372 (N_38372,N_36525,N_35923);
nand U38373 (N_38373,N_35882,N_37132);
or U38374 (N_38374,N_35759,N_35874);
and U38375 (N_38375,N_35128,N_37151);
nand U38376 (N_38376,N_36180,N_35630);
or U38377 (N_38377,N_35332,N_37314);
xor U38378 (N_38378,N_37031,N_35800);
nand U38379 (N_38379,N_37249,N_37369);
nor U38380 (N_38380,N_36509,N_36421);
xnor U38381 (N_38381,N_36545,N_36843);
nor U38382 (N_38382,N_36133,N_37461);
nor U38383 (N_38383,N_35299,N_35429);
nand U38384 (N_38384,N_36163,N_37455);
and U38385 (N_38385,N_36620,N_37328);
or U38386 (N_38386,N_35191,N_37499);
nor U38387 (N_38387,N_36794,N_37479);
and U38388 (N_38388,N_35591,N_36295);
or U38389 (N_38389,N_36943,N_35868);
and U38390 (N_38390,N_36597,N_36557);
nand U38391 (N_38391,N_36153,N_35960);
nand U38392 (N_38392,N_36726,N_37075);
nor U38393 (N_38393,N_36573,N_35109);
or U38394 (N_38394,N_36658,N_36941);
nand U38395 (N_38395,N_37133,N_37181);
nor U38396 (N_38396,N_37215,N_35963);
or U38397 (N_38397,N_35959,N_37138);
or U38398 (N_38398,N_36052,N_36503);
xor U38399 (N_38399,N_37432,N_35593);
xnor U38400 (N_38400,N_36177,N_35452);
nand U38401 (N_38401,N_36312,N_36031);
xor U38402 (N_38402,N_36361,N_37148);
xnor U38403 (N_38403,N_35377,N_37388);
nand U38404 (N_38404,N_35924,N_37363);
and U38405 (N_38405,N_36040,N_37346);
nor U38406 (N_38406,N_36014,N_37067);
and U38407 (N_38407,N_37289,N_36710);
xor U38408 (N_38408,N_37412,N_35520);
or U38409 (N_38409,N_36124,N_35705);
nand U38410 (N_38410,N_35784,N_35965);
and U38411 (N_38411,N_36104,N_35570);
and U38412 (N_38412,N_35376,N_37462);
nor U38413 (N_38413,N_36558,N_36795);
nand U38414 (N_38414,N_36375,N_37426);
and U38415 (N_38415,N_37159,N_36406);
or U38416 (N_38416,N_36515,N_35527);
and U38417 (N_38417,N_35184,N_36462);
nor U38418 (N_38418,N_36501,N_36913);
or U38419 (N_38419,N_36122,N_35565);
nor U38420 (N_38420,N_36915,N_35649);
nand U38421 (N_38421,N_35282,N_35861);
xor U38422 (N_38422,N_36005,N_35063);
xor U38423 (N_38423,N_36673,N_35013);
nand U38424 (N_38424,N_36252,N_35740);
nor U38425 (N_38425,N_37074,N_35629);
or U38426 (N_38426,N_35105,N_35842);
and U38427 (N_38427,N_35137,N_35730);
nand U38428 (N_38428,N_36867,N_35707);
nand U38429 (N_38429,N_35122,N_35758);
or U38430 (N_38430,N_37092,N_35879);
and U38431 (N_38431,N_35226,N_35383);
xnor U38432 (N_38432,N_35805,N_35792);
or U38433 (N_38433,N_36808,N_36522);
xnor U38434 (N_38434,N_37155,N_35256);
nand U38435 (N_38435,N_36073,N_35903);
xor U38436 (N_38436,N_35780,N_35812);
nor U38437 (N_38437,N_35447,N_36131);
and U38438 (N_38438,N_35270,N_36797);
nor U38439 (N_38439,N_36817,N_36650);
nand U38440 (N_38440,N_36946,N_36245);
xor U38441 (N_38441,N_35844,N_36570);
and U38442 (N_38442,N_36043,N_37000);
nor U38443 (N_38443,N_37472,N_35059);
nor U38444 (N_38444,N_36853,N_37030);
xnor U38445 (N_38445,N_37142,N_36586);
and U38446 (N_38446,N_37336,N_36033);
xor U38447 (N_38447,N_35671,N_36036);
or U38448 (N_38448,N_37440,N_36898);
nor U38449 (N_38449,N_36119,N_35664);
nand U38450 (N_38450,N_37286,N_35456);
or U38451 (N_38451,N_37228,N_35267);
or U38452 (N_38452,N_35984,N_35751);
or U38453 (N_38453,N_36565,N_35656);
xnor U38454 (N_38454,N_35373,N_37358);
or U38455 (N_38455,N_36751,N_35696);
nand U38456 (N_38456,N_36491,N_35529);
and U38457 (N_38457,N_36890,N_35020);
or U38458 (N_38458,N_36625,N_35739);
nand U38459 (N_38459,N_35614,N_36640);
nor U38460 (N_38460,N_37390,N_37321);
nand U38461 (N_38461,N_35440,N_36388);
xnor U38462 (N_38462,N_35051,N_37330);
and U38463 (N_38463,N_36145,N_36857);
nor U38464 (N_38464,N_35714,N_37337);
and U38465 (N_38465,N_35466,N_35037);
and U38466 (N_38466,N_35523,N_35219);
nand U38467 (N_38467,N_36980,N_36763);
or U38468 (N_38468,N_35360,N_36449);
and U38469 (N_38469,N_37207,N_37419);
nand U38470 (N_38470,N_36949,N_35091);
nand U38471 (N_38471,N_35790,N_37467);
or U38472 (N_38472,N_35955,N_37038);
xor U38473 (N_38473,N_35420,N_35813);
xor U38474 (N_38474,N_36750,N_36174);
nor U38475 (N_38475,N_35422,N_35734);
nand U38476 (N_38476,N_37435,N_36958);
nor U38477 (N_38477,N_35922,N_36654);
xnor U38478 (N_38478,N_36627,N_36664);
nand U38479 (N_38479,N_37238,N_35007);
or U38480 (N_38480,N_35144,N_36662);
nand U38481 (N_38481,N_35279,N_36336);
xnor U38482 (N_38482,N_36035,N_35100);
or U38483 (N_38483,N_35060,N_36499);
nor U38484 (N_38484,N_36500,N_35996);
or U38485 (N_38485,N_37210,N_36764);
nand U38486 (N_38486,N_36768,N_37078);
xnor U38487 (N_38487,N_35940,N_35247);
nor U38488 (N_38488,N_35272,N_35242);
or U38489 (N_38489,N_37178,N_36905);
nand U38490 (N_38490,N_35092,N_35473);
xor U38491 (N_38491,N_37107,N_37052);
nor U38492 (N_38492,N_37341,N_35345);
nor U38493 (N_38493,N_36302,N_35684);
or U38494 (N_38494,N_36269,N_36427);
nor U38495 (N_38495,N_36144,N_35588);
and U38496 (N_38496,N_35660,N_36990);
or U38497 (N_38497,N_35810,N_35229);
xnor U38498 (N_38498,N_35431,N_36185);
xor U38499 (N_38499,N_35288,N_37349);
or U38500 (N_38500,N_35369,N_36577);
xor U38501 (N_38501,N_36173,N_35540);
or U38502 (N_38502,N_36184,N_37061);
and U38503 (N_38503,N_35281,N_35902);
or U38504 (N_38504,N_35334,N_36425);
nand U38505 (N_38505,N_36072,N_37315);
xor U38506 (N_38506,N_36467,N_37377);
or U38507 (N_38507,N_36298,N_37149);
nand U38508 (N_38508,N_36715,N_35087);
or U38509 (N_38509,N_37375,N_37096);
nor U38510 (N_38510,N_36329,N_35797);
xor U38511 (N_38511,N_35968,N_37185);
xor U38512 (N_38512,N_36948,N_35589);
or U38513 (N_38513,N_36713,N_36325);
or U38514 (N_38514,N_36533,N_37416);
or U38515 (N_38515,N_36234,N_37162);
xnor U38516 (N_38516,N_35977,N_37060);
nand U38517 (N_38517,N_36553,N_36398);
nor U38518 (N_38518,N_36337,N_35971);
xor U38519 (N_38519,N_36006,N_37438);
and U38520 (N_38520,N_37237,N_36355);
nor U38521 (N_38521,N_37361,N_37134);
nor U38522 (N_38522,N_37113,N_36042);
and U38523 (N_38523,N_35166,N_35532);
and U38524 (N_38524,N_35934,N_36477);
and U38525 (N_38525,N_37020,N_36021);
nor U38526 (N_38526,N_36698,N_36893);
nor U38527 (N_38527,N_37368,N_36011);
nor U38528 (N_38528,N_36832,N_36226);
nor U38529 (N_38529,N_36617,N_35038);
or U38530 (N_38530,N_35067,N_36973);
and U38531 (N_38531,N_35423,N_36644);
nand U38532 (N_38532,N_37081,N_36551);
and U38533 (N_38533,N_37291,N_36672);
nand U38534 (N_38534,N_37424,N_36613);
nor U38535 (N_38535,N_37474,N_37399);
nor U38536 (N_38536,N_35775,N_36365);
and U38537 (N_38537,N_37131,N_35607);
or U38538 (N_38538,N_35992,N_35008);
nand U38539 (N_38539,N_36394,N_35276);
nor U38540 (N_38540,N_35014,N_35071);
nor U38541 (N_38541,N_35735,N_36985);
or U38542 (N_38542,N_35599,N_36786);
and U38543 (N_38543,N_35577,N_36976);
xor U38544 (N_38544,N_35876,N_35370);
and U38545 (N_38545,N_36663,N_35538);
or U38546 (N_38546,N_36633,N_36417);
xnor U38547 (N_38547,N_36171,N_35919);
nor U38548 (N_38548,N_36489,N_36346);
nor U38549 (N_38549,N_36634,N_36309);
xor U38550 (N_38550,N_35731,N_35635);
nand U38551 (N_38551,N_35023,N_35769);
xnor U38552 (N_38552,N_37408,N_36513);
or U38553 (N_38553,N_37108,N_37273);
xor U38554 (N_38554,N_35110,N_35846);
or U38555 (N_38555,N_37114,N_37420);
nor U38556 (N_38556,N_36149,N_37105);
or U38557 (N_38557,N_36164,N_37221);
nor U38558 (N_38558,N_36798,N_37073);
nor U38559 (N_38559,N_36339,N_36653);
or U38560 (N_38560,N_37347,N_35845);
xor U38561 (N_38561,N_37338,N_35822);
nor U38562 (N_38562,N_35702,N_36511);
xor U38563 (N_38563,N_36472,N_35077);
or U38564 (N_38564,N_36930,N_35918);
and U38565 (N_38565,N_36108,N_35104);
xnor U38566 (N_38566,N_35862,N_35151);
xnor U38567 (N_38567,N_37140,N_37428);
nand U38568 (N_38568,N_35010,N_35495);
nand U38569 (N_38569,N_36112,N_35418);
and U38570 (N_38570,N_35243,N_36009);
nand U38571 (N_38571,N_36248,N_36225);
nand U38572 (N_38572,N_35230,N_37481);
nand U38573 (N_38573,N_36440,N_36380);
xor U38574 (N_38574,N_35526,N_36258);
and U38575 (N_38575,N_36219,N_36029);
nor U38576 (N_38576,N_36071,N_37192);
nor U38577 (N_38577,N_35492,N_35147);
nor U38578 (N_38578,N_35433,N_35120);
nand U38579 (N_38579,N_36211,N_36695);
or U38580 (N_38580,N_35121,N_36055);
nand U38581 (N_38581,N_36785,N_35669);
or U38582 (N_38582,N_35233,N_35446);
nor U38583 (N_38583,N_36307,N_36502);
nor U38584 (N_38584,N_36830,N_37100);
or U38585 (N_38585,N_35634,N_35906);
nor U38586 (N_38586,N_37175,N_37054);
or U38587 (N_38587,N_35049,N_37469);
or U38588 (N_38588,N_37240,N_37339);
and U38589 (N_38589,N_36320,N_36285);
and U38590 (N_38590,N_36469,N_35280);
nand U38591 (N_38591,N_35827,N_35129);
and U38592 (N_38592,N_37295,N_35772);
nand U38593 (N_38593,N_36097,N_35179);
or U38594 (N_38594,N_36182,N_37403);
nor U38595 (N_38595,N_35478,N_36433);
nand U38596 (N_38596,N_36900,N_36714);
or U38597 (N_38597,N_35574,N_36841);
nor U38598 (N_38598,N_35765,N_35353);
and U38599 (N_38599,N_37251,N_36098);
xnor U38600 (N_38600,N_35808,N_36618);
nor U38601 (N_38601,N_35251,N_35891);
and U38602 (N_38602,N_35301,N_37045);
nor U38603 (N_38603,N_36034,N_36430);
xnor U38604 (N_38604,N_36802,N_35622);
and U38605 (N_38605,N_36942,N_35502);
nor U38606 (N_38606,N_35685,N_35829);
nor U38607 (N_38607,N_37115,N_36528);
nand U38608 (N_38608,N_36982,N_35424);
nand U38609 (N_38609,N_35779,N_36833);
xnor U38610 (N_38610,N_36549,N_35078);
or U38611 (N_38611,N_37182,N_36210);
xor U38612 (N_38612,N_36157,N_35371);
nand U38613 (N_38613,N_35300,N_35942);
xor U38614 (N_38614,N_37217,N_35390);
nor U38615 (N_38615,N_36316,N_36685);
nor U38616 (N_38616,N_35945,N_37018);
or U38617 (N_38617,N_35688,N_37284);
xnor U38618 (N_38618,N_36092,N_36369);
and U38619 (N_38619,N_35335,N_36578);
and U38620 (N_38620,N_36556,N_36498);
or U38621 (N_38621,N_37446,N_37434);
and U38622 (N_38622,N_36333,N_35459);
or U38623 (N_38623,N_35956,N_36061);
nor U38624 (N_38624,N_37342,N_35749);
nand U38625 (N_38625,N_36431,N_35152);
or U38626 (N_38626,N_37303,N_37014);
or U38627 (N_38627,N_37417,N_36089);
or U38628 (N_38628,N_36919,N_36552);
nor U38629 (N_38629,N_35987,N_35450);
xor U38630 (N_38630,N_36438,N_36429);
and U38631 (N_38631,N_36060,N_37386);
nor U38632 (N_38632,N_36051,N_35534);
or U38633 (N_38633,N_35410,N_36414);
or U38634 (N_38634,N_36493,N_36273);
or U38635 (N_38635,N_36767,N_37280);
and U38636 (N_38636,N_36783,N_37191);
xor U38637 (N_38637,N_35628,N_36321);
nand U38638 (N_38638,N_36755,N_37478);
nor U38639 (N_38639,N_35480,N_36343);
and U38640 (N_38640,N_36711,N_37239);
xnor U38641 (N_38641,N_35126,N_35801);
or U38642 (N_38642,N_37077,N_37190);
nor U38643 (N_38643,N_35050,N_36780);
nand U38644 (N_38644,N_36696,N_37290);
and U38645 (N_38645,N_37066,N_36056);
nor U38646 (N_38646,N_36251,N_35724);
xor U38647 (N_38647,N_36212,N_37444);
nor U38648 (N_38648,N_35416,N_36966);
nand U38649 (N_38649,N_36932,N_35728);
xor U38650 (N_38650,N_36721,N_36877);
or U38651 (N_38651,N_35437,N_35962);
nor U38652 (N_38652,N_35894,N_35053);
and U38653 (N_38653,N_36324,N_35703);
or U38654 (N_38654,N_36622,N_36291);
and U38655 (N_38655,N_35877,N_35881);
or U38656 (N_38656,N_37471,N_37118);
and U38657 (N_38657,N_36727,N_35847);
nand U38658 (N_38658,N_36657,N_36961);
xnor U38659 (N_38659,N_36279,N_37261);
xor U38660 (N_38660,N_36582,N_35516);
nand U38661 (N_38661,N_35572,N_35837);
and U38662 (N_38662,N_35083,N_35086);
nand U38663 (N_38663,N_36024,N_36468);
xnor U38664 (N_38664,N_35413,N_37452);
xor U38665 (N_38665,N_35095,N_35579);
nor U38666 (N_38666,N_36016,N_35828);
xnor U38667 (N_38667,N_36246,N_35638);
nor U38668 (N_38668,N_36270,N_35594);
nor U38669 (N_38669,N_37264,N_36323);
nand U38670 (N_38670,N_37034,N_37220);
xor U38671 (N_38671,N_35292,N_35559);
nor U38672 (N_38672,N_36360,N_35597);
or U38673 (N_38673,N_35852,N_36819);
or U38674 (N_38674,N_36303,N_35185);
nor U38675 (N_38675,N_36187,N_35761);
and U38676 (N_38676,N_35615,N_35781);
nand U38677 (N_38677,N_35901,N_36837);
or U38678 (N_38678,N_36581,N_36359);
nand U38679 (N_38679,N_36975,N_36268);
nand U38680 (N_38680,N_35897,N_35359);
and U38681 (N_38681,N_37188,N_36485);
and U38682 (N_38682,N_36825,N_35205);
or U38683 (N_38683,N_35683,N_36850);
and U38684 (N_38684,N_35090,N_35443);
nand U38685 (N_38685,N_35097,N_36784);
nor U38686 (N_38686,N_35954,N_36276);
or U38687 (N_38687,N_37275,N_35181);
nor U38688 (N_38688,N_35022,N_36516);
nand U38689 (N_38689,N_37102,N_37316);
or U38690 (N_38690,N_37241,N_35042);
nand U38691 (N_38691,N_35261,N_35035);
xor U38692 (N_38692,N_37395,N_37050);
nand U38693 (N_38693,N_37016,N_35017);
or U38694 (N_38694,N_36028,N_36495);
or U38695 (N_38695,N_35499,N_35883);
and U38696 (N_38696,N_35639,N_35310);
and U38697 (N_38697,N_35834,N_35571);
and U38698 (N_38698,N_35329,N_35117);
xnor U38699 (N_38699,N_37086,N_35065);
and U38700 (N_38700,N_36519,N_35601);
nor U38701 (N_38701,N_35927,N_37028);
and U38702 (N_38702,N_35652,N_35537);
nor U38703 (N_38703,N_37101,N_36788);
xor U38704 (N_38704,N_37087,N_37173);
and U38705 (N_38705,N_35044,N_37121);
and U38706 (N_38706,N_35164,N_35350);
or U38707 (N_38707,N_35528,N_36840);
and U38708 (N_38708,N_36207,N_35712);
or U38709 (N_38709,N_36299,N_37137);
and U38710 (N_38710,N_36373,N_36132);
xnor U38711 (N_38711,N_36264,N_35445);
nand U38712 (N_38712,N_37004,N_37410);
nor U38713 (N_38713,N_35011,N_35415);
or U38714 (N_38714,N_36972,N_36924);
and U38715 (N_38715,N_37422,N_37144);
nand U38716 (N_38716,N_37168,N_36231);
nand U38717 (N_38717,N_35948,N_36923);
xor U38718 (N_38718,N_37150,N_35286);
xnor U38719 (N_38719,N_36675,N_35788);
and U38720 (N_38720,N_36828,N_35175);
and U38721 (N_38721,N_35625,N_37011);
nor U38722 (N_38722,N_37047,N_36871);
or U38723 (N_38723,N_35337,N_37351);
nor U38724 (N_38724,N_35935,N_36762);
xor U38725 (N_38725,N_35244,N_36862);
and U38726 (N_38726,N_36847,N_36748);
or U38727 (N_38727,N_36836,N_36460);
xor U38728 (N_38728,N_35043,N_35457);
xnor U38729 (N_38729,N_37313,N_36256);
nand U38730 (N_38730,N_37329,N_36799);
nand U38731 (N_38731,N_35508,N_35947);
nand U38732 (N_38732,N_37259,N_36530);
nor U38733 (N_38733,N_36049,N_36081);
xor U38734 (N_38734,N_35015,N_35066);
nand U38735 (N_38735,N_36310,N_37015);
nand U38736 (N_38736,N_35318,N_35858);
xor U38737 (N_38737,N_35679,N_36396);
xnor U38738 (N_38738,N_36257,N_36115);
or U38739 (N_38739,N_36148,N_35618);
nor U38740 (N_38740,N_35880,N_35578);
or U38741 (N_38741,N_37019,N_35106);
nor U38742 (N_38742,N_36423,N_35503);
nand U38743 (N_38743,N_35048,N_37305);
xnor U38744 (N_38744,N_35070,N_35785);
and U38745 (N_38745,N_36065,N_37405);
or U38746 (N_38746,N_35214,N_37082);
or U38747 (N_38747,N_35692,N_36735);
and U38748 (N_38748,N_36889,N_36142);
nand U38749 (N_38749,N_37374,N_35196);
and U38750 (N_38750,N_36083,N_36798);
or U38751 (N_38751,N_36479,N_37202);
and U38752 (N_38752,N_35190,N_35620);
nor U38753 (N_38753,N_35466,N_35524);
nor U38754 (N_38754,N_36711,N_35296);
nor U38755 (N_38755,N_37446,N_35016);
xor U38756 (N_38756,N_37122,N_35079);
or U38757 (N_38757,N_35830,N_35154);
nor U38758 (N_38758,N_37313,N_36441);
nand U38759 (N_38759,N_36905,N_36450);
or U38760 (N_38760,N_36211,N_36017);
or U38761 (N_38761,N_36289,N_35092);
xor U38762 (N_38762,N_35227,N_35752);
xor U38763 (N_38763,N_36947,N_37215);
and U38764 (N_38764,N_36437,N_35999);
xnor U38765 (N_38765,N_36273,N_36149);
nor U38766 (N_38766,N_36980,N_36266);
nand U38767 (N_38767,N_36278,N_35795);
xnor U38768 (N_38768,N_37297,N_37067);
and U38769 (N_38769,N_36288,N_35857);
xor U38770 (N_38770,N_35929,N_35996);
nand U38771 (N_38771,N_35069,N_35317);
nor U38772 (N_38772,N_35160,N_35689);
nor U38773 (N_38773,N_36325,N_35885);
and U38774 (N_38774,N_35807,N_35485);
and U38775 (N_38775,N_37027,N_36194);
and U38776 (N_38776,N_37497,N_35977);
xor U38777 (N_38777,N_35156,N_35109);
or U38778 (N_38778,N_35821,N_37478);
xor U38779 (N_38779,N_35130,N_36780);
nand U38780 (N_38780,N_35061,N_36808);
nor U38781 (N_38781,N_35569,N_35386);
xnor U38782 (N_38782,N_35185,N_35715);
and U38783 (N_38783,N_36150,N_36829);
and U38784 (N_38784,N_35234,N_36193);
and U38785 (N_38785,N_37256,N_37464);
or U38786 (N_38786,N_36527,N_36280);
and U38787 (N_38787,N_37282,N_36307);
xor U38788 (N_38788,N_37474,N_37055);
xnor U38789 (N_38789,N_35629,N_35789);
nand U38790 (N_38790,N_36426,N_35097);
nor U38791 (N_38791,N_35326,N_35562);
nand U38792 (N_38792,N_35271,N_36968);
xnor U38793 (N_38793,N_37165,N_37096);
nor U38794 (N_38794,N_36698,N_36155);
nor U38795 (N_38795,N_37129,N_35798);
or U38796 (N_38796,N_36935,N_36571);
and U38797 (N_38797,N_35559,N_36463);
xor U38798 (N_38798,N_36354,N_35782);
and U38799 (N_38799,N_35825,N_36606);
or U38800 (N_38800,N_35786,N_36630);
or U38801 (N_38801,N_35045,N_36153);
and U38802 (N_38802,N_37381,N_37278);
and U38803 (N_38803,N_36208,N_35555);
and U38804 (N_38804,N_36234,N_37240);
or U38805 (N_38805,N_37089,N_36366);
or U38806 (N_38806,N_37218,N_35532);
nor U38807 (N_38807,N_37343,N_35542);
xnor U38808 (N_38808,N_35484,N_36471);
nand U38809 (N_38809,N_36921,N_35861);
nor U38810 (N_38810,N_37052,N_35731);
xnor U38811 (N_38811,N_36123,N_35126);
xnor U38812 (N_38812,N_36334,N_36911);
xor U38813 (N_38813,N_37358,N_35775);
nor U38814 (N_38814,N_35677,N_36461);
nor U38815 (N_38815,N_35256,N_35510);
nand U38816 (N_38816,N_37043,N_35904);
nor U38817 (N_38817,N_35739,N_37426);
nand U38818 (N_38818,N_36549,N_35124);
xnor U38819 (N_38819,N_35123,N_35272);
nor U38820 (N_38820,N_36357,N_36706);
and U38821 (N_38821,N_35554,N_36604);
and U38822 (N_38822,N_36611,N_36758);
xor U38823 (N_38823,N_36437,N_35727);
nand U38824 (N_38824,N_37290,N_35636);
xor U38825 (N_38825,N_37342,N_36400);
nand U38826 (N_38826,N_35564,N_35353);
and U38827 (N_38827,N_36657,N_35611);
xnor U38828 (N_38828,N_37250,N_37207);
or U38829 (N_38829,N_35876,N_35634);
xor U38830 (N_38830,N_35482,N_36464);
nand U38831 (N_38831,N_36421,N_35013);
nor U38832 (N_38832,N_35597,N_35410);
nor U38833 (N_38833,N_35557,N_36877);
xnor U38834 (N_38834,N_37344,N_35114);
nor U38835 (N_38835,N_35476,N_37108);
or U38836 (N_38836,N_37463,N_35444);
nand U38837 (N_38837,N_35260,N_36881);
and U38838 (N_38838,N_36367,N_35496);
or U38839 (N_38839,N_37170,N_36379);
nand U38840 (N_38840,N_37213,N_37174);
nand U38841 (N_38841,N_36644,N_35244);
nor U38842 (N_38842,N_37137,N_35813);
nor U38843 (N_38843,N_36646,N_36270);
nand U38844 (N_38844,N_36502,N_35780);
nor U38845 (N_38845,N_35422,N_36118);
xnor U38846 (N_38846,N_37427,N_37453);
or U38847 (N_38847,N_36603,N_36557);
nor U38848 (N_38848,N_36447,N_36670);
nand U38849 (N_38849,N_37248,N_36399);
nand U38850 (N_38850,N_35101,N_36447);
nand U38851 (N_38851,N_37305,N_35184);
xor U38852 (N_38852,N_37032,N_37266);
xnor U38853 (N_38853,N_35624,N_35958);
nand U38854 (N_38854,N_36957,N_35623);
or U38855 (N_38855,N_36421,N_35264);
nand U38856 (N_38856,N_35899,N_36492);
nor U38857 (N_38857,N_36874,N_36088);
xor U38858 (N_38858,N_35596,N_35903);
or U38859 (N_38859,N_35037,N_35565);
nor U38860 (N_38860,N_35361,N_36553);
nand U38861 (N_38861,N_36843,N_36372);
and U38862 (N_38862,N_35397,N_37146);
nor U38863 (N_38863,N_36386,N_35379);
nand U38864 (N_38864,N_36045,N_37466);
or U38865 (N_38865,N_37395,N_36069);
and U38866 (N_38866,N_37188,N_35116);
or U38867 (N_38867,N_35755,N_36297);
xnor U38868 (N_38868,N_35989,N_37165);
or U38869 (N_38869,N_36441,N_36341);
nor U38870 (N_38870,N_35479,N_35652);
xor U38871 (N_38871,N_37004,N_36335);
or U38872 (N_38872,N_35908,N_35817);
xnor U38873 (N_38873,N_36492,N_37305);
xnor U38874 (N_38874,N_35789,N_35782);
nand U38875 (N_38875,N_36603,N_37280);
or U38876 (N_38876,N_35382,N_37097);
nand U38877 (N_38877,N_36954,N_36410);
nand U38878 (N_38878,N_36643,N_36633);
or U38879 (N_38879,N_37187,N_36502);
xnor U38880 (N_38880,N_37429,N_35188);
or U38881 (N_38881,N_36790,N_35141);
or U38882 (N_38882,N_35299,N_35961);
xor U38883 (N_38883,N_35725,N_37343);
nand U38884 (N_38884,N_35985,N_35257);
xor U38885 (N_38885,N_37005,N_36490);
nand U38886 (N_38886,N_36738,N_35031);
xor U38887 (N_38887,N_35444,N_36205);
nor U38888 (N_38888,N_35078,N_35847);
nor U38889 (N_38889,N_35587,N_37248);
xnor U38890 (N_38890,N_35542,N_37159);
or U38891 (N_38891,N_36043,N_37282);
or U38892 (N_38892,N_36869,N_36119);
xor U38893 (N_38893,N_37308,N_35881);
or U38894 (N_38894,N_36993,N_35054);
or U38895 (N_38895,N_36276,N_36838);
and U38896 (N_38896,N_36458,N_36522);
or U38897 (N_38897,N_37457,N_36163);
nor U38898 (N_38898,N_36950,N_37422);
and U38899 (N_38899,N_37124,N_36624);
nand U38900 (N_38900,N_35460,N_36344);
and U38901 (N_38901,N_37128,N_35428);
nand U38902 (N_38902,N_35451,N_35799);
nor U38903 (N_38903,N_35779,N_36402);
or U38904 (N_38904,N_36466,N_35219);
xnor U38905 (N_38905,N_36588,N_37232);
nor U38906 (N_38906,N_35440,N_37154);
nand U38907 (N_38907,N_37142,N_36798);
and U38908 (N_38908,N_35948,N_35861);
nand U38909 (N_38909,N_35668,N_36910);
or U38910 (N_38910,N_35066,N_36357);
nor U38911 (N_38911,N_36737,N_35276);
nor U38912 (N_38912,N_37418,N_37330);
xor U38913 (N_38913,N_36818,N_35962);
xor U38914 (N_38914,N_36685,N_36225);
or U38915 (N_38915,N_35251,N_35589);
xor U38916 (N_38916,N_36558,N_35530);
and U38917 (N_38917,N_36913,N_37314);
nor U38918 (N_38918,N_35758,N_37393);
xor U38919 (N_38919,N_35128,N_35556);
xor U38920 (N_38920,N_35084,N_37075);
nor U38921 (N_38921,N_35130,N_36693);
nand U38922 (N_38922,N_37286,N_35597);
nor U38923 (N_38923,N_35020,N_36767);
or U38924 (N_38924,N_35979,N_36807);
nand U38925 (N_38925,N_36231,N_35444);
and U38926 (N_38926,N_37346,N_36597);
xor U38927 (N_38927,N_36678,N_35089);
or U38928 (N_38928,N_36724,N_35234);
and U38929 (N_38929,N_36193,N_35298);
nand U38930 (N_38930,N_37014,N_35848);
xor U38931 (N_38931,N_35310,N_35483);
xor U38932 (N_38932,N_37238,N_35358);
and U38933 (N_38933,N_35770,N_36947);
and U38934 (N_38934,N_37188,N_36599);
nand U38935 (N_38935,N_37165,N_35119);
or U38936 (N_38936,N_37089,N_36048);
nand U38937 (N_38937,N_35779,N_37212);
or U38938 (N_38938,N_35172,N_36362);
and U38939 (N_38939,N_37173,N_36412);
and U38940 (N_38940,N_36125,N_37207);
and U38941 (N_38941,N_35478,N_35471);
nor U38942 (N_38942,N_36088,N_37291);
or U38943 (N_38943,N_36094,N_35717);
nand U38944 (N_38944,N_36591,N_35071);
nor U38945 (N_38945,N_36348,N_35254);
and U38946 (N_38946,N_36409,N_36766);
nand U38947 (N_38947,N_36938,N_36896);
nor U38948 (N_38948,N_37361,N_37042);
xnor U38949 (N_38949,N_37477,N_36654);
nand U38950 (N_38950,N_35633,N_35398);
and U38951 (N_38951,N_37396,N_36602);
nand U38952 (N_38952,N_36011,N_35810);
and U38953 (N_38953,N_36243,N_37445);
and U38954 (N_38954,N_35035,N_37003);
nand U38955 (N_38955,N_35926,N_35584);
or U38956 (N_38956,N_36279,N_37198);
nand U38957 (N_38957,N_37179,N_36170);
or U38958 (N_38958,N_36436,N_35726);
or U38959 (N_38959,N_35330,N_35303);
or U38960 (N_38960,N_35830,N_35393);
nor U38961 (N_38961,N_37146,N_36530);
nand U38962 (N_38962,N_37292,N_35434);
xnor U38963 (N_38963,N_37207,N_37296);
and U38964 (N_38964,N_35391,N_36605);
xnor U38965 (N_38965,N_37100,N_36997);
or U38966 (N_38966,N_35707,N_35852);
xor U38967 (N_38967,N_36629,N_35849);
nor U38968 (N_38968,N_35128,N_36976);
or U38969 (N_38969,N_37287,N_36705);
xnor U38970 (N_38970,N_36291,N_35293);
nand U38971 (N_38971,N_35385,N_35912);
nor U38972 (N_38972,N_36663,N_35705);
nand U38973 (N_38973,N_35618,N_36002);
nor U38974 (N_38974,N_36389,N_36965);
nand U38975 (N_38975,N_36721,N_37349);
and U38976 (N_38976,N_36433,N_36513);
or U38977 (N_38977,N_36071,N_35588);
xor U38978 (N_38978,N_36173,N_36274);
nand U38979 (N_38979,N_35851,N_35655);
nor U38980 (N_38980,N_35579,N_35470);
xor U38981 (N_38981,N_36298,N_36256);
nor U38982 (N_38982,N_35278,N_35771);
nand U38983 (N_38983,N_36992,N_35348);
nand U38984 (N_38984,N_37104,N_36759);
nor U38985 (N_38985,N_37117,N_36428);
nand U38986 (N_38986,N_35086,N_36764);
nand U38987 (N_38987,N_35576,N_35921);
or U38988 (N_38988,N_35376,N_37343);
nor U38989 (N_38989,N_35485,N_35270);
nand U38990 (N_38990,N_35380,N_35873);
or U38991 (N_38991,N_36860,N_36823);
and U38992 (N_38992,N_36764,N_37398);
and U38993 (N_38993,N_36881,N_36191);
or U38994 (N_38994,N_35018,N_36779);
nor U38995 (N_38995,N_35412,N_36435);
and U38996 (N_38996,N_36698,N_37284);
nor U38997 (N_38997,N_36253,N_36663);
xor U38998 (N_38998,N_36075,N_36429);
xnor U38999 (N_38999,N_36916,N_37380);
nor U39000 (N_39000,N_37307,N_36234);
xnor U39001 (N_39001,N_36164,N_37207);
and U39002 (N_39002,N_36323,N_36893);
and U39003 (N_39003,N_35925,N_37082);
or U39004 (N_39004,N_36201,N_36021);
nand U39005 (N_39005,N_35908,N_36893);
or U39006 (N_39006,N_35230,N_36083);
or U39007 (N_39007,N_36530,N_35100);
nand U39008 (N_39008,N_35486,N_37344);
xnor U39009 (N_39009,N_35891,N_36508);
xor U39010 (N_39010,N_36218,N_35619);
nor U39011 (N_39011,N_36235,N_37288);
xnor U39012 (N_39012,N_35077,N_35648);
nand U39013 (N_39013,N_37078,N_37104);
xor U39014 (N_39014,N_36149,N_35528);
nand U39015 (N_39015,N_36132,N_37428);
and U39016 (N_39016,N_36533,N_35555);
nor U39017 (N_39017,N_36951,N_36578);
and U39018 (N_39018,N_36049,N_37493);
nor U39019 (N_39019,N_36145,N_35080);
nor U39020 (N_39020,N_36732,N_37131);
or U39021 (N_39021,N_36963,N_36722);
nand U39022 (N_39022,N_36011,N_35693);
or U39023 (N_39023,N_35906,N_36707);
nor U39024 (N_39024,N_36026,N_35221);
or U39025 (N_39025,N_36363,N_35466);
and U39026 (N_39026,N_35150,N_35323);
and U39027 (N_39027,N_36573,N_37243);
xnor U39028 (N_39028,N_36560,N_36417);
xnor U39029 (N_39029,N_35464,N_36408);
and U39030 (N_39030,N_37000,N_36817);
or U39031 (N_39031,N_37361,N_35137);
and U39032 (N_39032,N_36648,N_36730);
or U39033 (N_39033,N_37355,N_36826);
xor U39034 (N_39034,N_37494,N_37390);
or U39035 (N_39035,N_36441,N_37350);
xor U39036 (N_39036,N_36767,N_35850);
or U39037 (N_39037,N_37234,N_36525);
nand U39038 (N_39038,N_36539,N_35601);
xor U39039 (N_39039,N_37452,N_37327);
and U39040 (N_39040,N_36658,N_35745);
and U39041 (N_39041,N_35210,N_37303);
nor U39042 (N_39042,N_35237,N_36283);
or U39043 (N_39043,N_36767,N_35758);
nand U39044 (N_39044,N_35929,N_35661);
xor U39045 (N_39045,N_37134,N_35757);
and U39046 (N_39046,N_37109,N_36864);
xnor U39047 (N_39047,N_36615,N_36065);
nand U39048 (N_39048,N_35859,N_36205);
or U39049 (N_39049,N_35274,N_35101);
xor U39050 (N_39050,N_37060,N_36114);
and U39051 (N_39051,N_35262,N_35552);
or U39052 (N_39052,N_35121,N_36577);
or U39053 (N_39053,N_35894,N_35652);
and U39054 (N_39054,N_36850,N_37033);
and U39055 (N_39055,N_35372,N_35148);
or U39056 (N_39056,N_36856,N_36449);
xor U39057 (N_39057,N_36350,N_37026);
or U39058 (N_39058,N_35920,N_37356);
and U39059 (N_39059,N_35525,N_35951);
nor U39060 (N_39060,N_35838,N_35813);
and U39061 (N_39061,N_36788,N_35833);
nor U39062 (N_39062,N_36430,N_36108);
and U39063 (N_39063,N_36074,N_37316);
nor U39064 (N_39064,N_36001,N_35721);
or U39065 (N_39065,N_37207,N_35857);
nand U39066 (N_39066,N_35959,N_35367);
xor U39067 (N_39067,N_37229,N_37495);
nand U39068 (N_39068,N_37274,N_36727);
xnor U39069 (N_39069,N_35222,N_35580);
xor U39070 (N_39070,N_35353,N_36884);
nor U39071 (N_39071,N_37354,N_36227);
and U39072 (N_39072,N_35742,N_36258);
nor U39073 (N_39073,N_36236,N_35393);
nand U39074 (N_39074,N_36060,N_37492);
or U39075 (N_39075,N_35072,N_36858);
nor U39076 (N_39076,N_35391,N_35614);
nand U39077 (N_39077,N_36052,N_36056);
or U39078 (N_39078,N_35601,N_35321);
nor U39079 (N_39079,N_35000,N_35673);
and U39080 (N_39080,N_36099,N_35234);
nor U39081 (N_39081,N_36852,N_37117);
xnor U39082 (N_39082,N_36305,N_36986);
or U39083 (N_39083,N_36662,N_36567);
or U39084 (N_39084,N_35178,N_36043);
xor U39085 (N_39085,N_36919,N_36306);
and U39086 (N_39086,N_37288,N_37344);
nor U39087 (N_39087,N_35672,N_36777);
xor U39088 (N_39088,N_36070,N_36718);
xnor U39089 (N_39089,N_37202,N_36469);
xnor U39090 (N_39090,N_35782,N_36783);
nand U39091 (N_39091,N_37147,N_35729);
xor U39092 (N_39092,N_36371,N_35072);
xnor U39093 (N_39093,N_37332,N_35237);
nor U39094 (N_39094,N_36436,N_36278);
or U39095 (N_39095,N_37389,N_35165);
or U39096 (N_39096,N_35522,N_35351);
nand U39097 (N_39097,N_35897,N_36134);
or U39098 (N_39098,N_35686,N_35627);
nor U39099 (N_39099,N_36268,N_36169);
nor U39100 (N_39100,N_36675,N_36705);
or U39101 (N_39101,N_36607,N_35581);
or U39102 (N_39102,N_35990,N_36102);
nand U39103 (N_39103,N_36259,N_35324);
nor U39104 (N_39104,N_36451,N_36641);
xor U39105 (N_39105,N_37300,N_35158);
nand U39106 (N_39106,N_35093,N_35632);
xnor U39107 (N_39107,N_35049,N_35970);
nor U39108 (N_39108,N_37485,N_35277);
xnor U39109 (N_39109,N_36331,N_35521);
or U39110 (N_39110,N_37208,N_35891);
xnor U39111 (N_39111,N_36945,N_36907);
xnor U39112 (N_39112,N_35302,N_36771);
nand U39113 (N_39113,N_36378,N_36267);
nor U39114 (N_39114,N_36860,N_36154);
or U39115 (N_39115,N_35385,N_36482);
nor U39116 (N_39116,N_36906,N_35748);
nor U39117 (N_39117,N_35096,N_37368);
nor U39118 (N_39118,N_35030,N_37421);
or U39119 (N_39119,N_37467,N_36623);
and U39120 (N_39120,N_37354,N_37431);
nand U39121 (N_39121,N_37069,N_35915);
nor U39122 (N_39122,N_35224,N_36020);
xor U39123 (N_39123,N_36244,N_35536);
or U39124 (N_39124,N_36355,N_36597);
nor U39125 (N_39125,N_35833,N_37499);
xnor U39126 (N_39126,N_35548,N_36322);
and U39127 (N_39127,N_36578,N_37266);
or U39128 (N_39128,N_35083,N_36507);
nand U39129 (N_39129,N_35744,N_37458);
xnor U39130 (N_39130,N_35869,N_37323);
or U39131 (N_39131,N_36711,N_37102);
nand U39132 (N_39132,N_35594,N_36219);
nand U39133 (N_39133,N_35431,N_35714);
or U39134 (N_39134,N_35463,N_35813);
nor U39135 (N_39135,N_36546,N_36843);
xor U39136 (N_39136,N_35794,N_36035);
and U39137 (N_39137,N_36505,N_35811);
and U39138 (N_39138,N_35667,N_36098);
xnor U39139 (N_39139,N_36804,N_36260);
xnor U39140 (N_39140,N_35088,N_35557);
and U39141 (N_39141,N_35065,N_36867);
or U39142 (N_39142,N_37303,N_36785);
and U39143 (N_39143,N_35660,N_36282);
xnor U39144 (N_39144,N_36962,N_35074);
nor U39145 (N_39145,N_35908,N_37305);
nand U39146 (N_39146,N_36693,N_35728);
nor U39147 (N_39147,N_37381,N_36211);
nor U39148 (N_39148,N_36191,N_36833);
or U39149 (N_39149,N_36713,N_36657);
nor U39150 (N_39150,N_37394,N_35391);
xor U39151 (N_39151,N_36083,N_36917);
nand U39152 (N_39152,N_37430,N_36102);
xor U39153 (N_39153,N_36175,N_36800);
xnor U39154 (N_39154,N_37008,N_37060);
and U39155 (N_39155,N_36876,N_35097);
xnor U39156 (N_39156,N_35178,N_36198);
or U39157 (N_39157,N_36003,N_37342);
nor U39158 (N_39158,N_35423,N_35710);
xor U39159 (N_39159,N_36297,N_35317);
nand U39160 (N_39160,N_37223,N_36030);
xor U39161 (N_39161,N_35472,N_36008);
nor U39162 (N_39162,N_36940,N_36966);
nand U39163 (N_39163,N_36209,N_36557);
and U39164 (N_39164,N_37465,N_37125);
or U39165 (N_39165,N_36941,N_36664);
xnor U39166 (N_39166,N_36151,N_36380);
xnor U39167 (N_39167,N_35325,N_37025);
nor U39168 (N_39168,N_36374,N_36373);
nand U39169 (N_39169,N_36640,N_35172);
nand U39170 (N_39170,N_35603,N_35922);
nor U39171 (N_39171,N_35251,N_36806);
nand U39172 (N_39172,N_36421,N_35474);
and U39173 (N_39173,N_37151,N_36594);
xor U39174 (N_39174,N_36708,N_35809);
nor U39175 (N_39175,N_35188,N_37141);
or U39176 (N_39176,N_36631,N_36617);
and U39177 (N_39177,N_36940,N_35460);
and U39178 (N_39178,N_36305,N_35599);
xor U39179 (N_39179,N_35868,N_35667);
nand U39180 (N_39180,N_35179,N_36545);
nand U39181 (N_39181,N_35008,N_36946);
xnor U39182 (N_39182,N_36286,N_35636);
and U39183 (N_39183,N_37216,N_35180);
and U39184 (N_39184,N_37132,N_36003);
or U39185 (N_39185,N_35563,N_36365);
nand U39186 (N_39186,N_37357,N_36811);
nand U39187 (N_39187,N_37348,N_36764);
and U39188 (N_39188,N_36847,N_36053);
and U39189 (N_39189,N_36426,N_35437);
nor U39190 (N_39190,N_35003,N_35046);
nand U39191 (N_39191,N_35033,N_35467);
or U39192 (N_39192,N_36379,N_37220);
nand U39193 (N_39193,N_36336,N_36023);
nor U39194 (N_39194,N_35541,N_35390);
xnor U39195 (N_39195,N_35180,N_36793);
nand U39196 (N_39196,N_36865,N_36697);
or U39197 (N_39197,N_36466,N_35892);
nand U39198 (N_39198,N_37426,N_36236);
nand U39199 (N_39199,N_35720,N_36801);
nand U39200 (N_39200,N_35720,N_36441);
and U39201 (N_39201,N_36255,N_35768);
or U39202 (N_39202,N_35668,N_37177);
xnor U39203 (N_39203,N_37075,N_36480);
and U39204 (N_39204,N_37112,N_35033);
nand U39205 (N_39205,N_35442,N_37208);
or U39206 (N_39206,N_36250,N_35325);
nor U39207 (N_39207,N_37493,N_36868);
and U39208 (N_39208,N_36876,N_35597);
nand U39209 (N_39209,N_37082,N_37399);
and U39210 (N_39210,N_35521,N_36007);
or U39211 (N_39211,N_35434,N_36160);
nor U39212 (N_39212,N_35571,N_36506);
nand U39213 (N_39213,N_36856,N_35994);
nor U39214 (N_39214,N_36542,N_37467);
xnor U39215 (N_39215,N_37189,N_36984);
xnor U39216 (N_39216,N_36876,N_36168);
and U39217 (N_39217,N_36278,N_37382);
nor U39218 (N_39218,N_36413,N_35663);
or U39219 (N_39219,N_35062,N_36875);
or U39220 (N_39220,N_35919,N_35051);
and U39221 (N_39221,N_35988,N_35157);
nand U39222 (N_39222,N_37138,N_37160);
or U39223 (N_39223,N_35864,N_35388);
and U39224 (N_39224,N_36252,N_36716);
xor U39225 (N_39225,N_36906,N_35030);
nand U39226 (N_39226,N_35687,N_35928);
and U39227 (N_39227,N_35875,N_36161);
nor U39228 (N_39228,N_36126,N_35060);
or U39229 (N_39229,N_36969,N_35437);
or U39230 (N_39230,N_37181,N_35824);
or U39231 (N_39231,N_35035,N_37321);
and U39232 (N_39232,N_35956,N_35762);
or U39233 (N_39233,N_37087,N_35471);
xnor U39234 (N_39234,N_35326,N_36305);
or U39235 (N_39235,N_35240,N_35412);
and U39236 (N_39236,N_36961,N_35038);
nor U39237 (N_39237,N_36729,N_37347);
xor U39238 (N_39238,N_37112,N_35861);
or U39239 (N_39239,N_36465,N_37179);
xor U39240 (N_39240,N_35790,N_37439);
and U39241 (N_39241,N_36237,N_36835);
nand U39242 (N_39242,N_35402,N_36580);
or U39243 (N_39243,N_35254,N_36248);
nand U39244 (N_39244,N_36256,N_36260);
or U39245 (N_39245,N_35993,N_35223);
xor U39246 (N_39246,N_35638,N_35687);
nor U39247 (N_39247,N_37083,N_35585);
and U39248 (N_39248,N_35007,N_35985);
nand U39249 (N_39249,N_37071,N_35718);
and U39250 (N_39250,N_36280,N_36752);
or U39251 (N_39251,N_37172,N_36317);
nand U39252 (N_39252,N_36819,N_37111);
xnor U39253 (N_39253,N_37297,N_37090);
or U39254 (N_39254,N_37492,N_37283);
nor U39255 (N_39255,N_36386,N_35706);
nand U39256 (N_39256,N_35517,N_36745);
xor U39257 (N_39257,N_36418,N_35352);
nor U39258 (N_39258,N_36693,N_35439);
xnor U39259 (N_39259,N_36296,N_35714);
nand U39260 (N_39260,N_35680,N_35945);
nand U39261 (N_39261,N_35869,N_36076);
xnor U39262 (N_39262,N_36566,N_36571);
xnor U39263 (N_39263,N_36040,N_37115);
nor U39264 (N_39264,N_36808,N_36287);
and U39265 (N_39265,N_35680,N_35353);
and U39266 (N_39266,N_35607,N_36949);
nor U39267 (N_39267,N_37142,N_35472);
and U39268 (N_39268,N_36408,N_36345);
nor U39269 (N_39269,N_37036,N_35088);
nor U39270 (N_39270,N_37235,N_36856);
xnor U39271 (N_39271,N_36307,N_36587);
or U39272 (N_39272,N_36284,N_35377);
nor U39273 (N_39273,N_36807,N_36687);
or U39274 (N_39274,N_35080,N_37114);
and U39275 (N_39275,N_37373,N_36272);
and U39276 (N_39276,N_36445,N_35611);
nand U39277 (N_39277,N_35272,N_36285);
or U39278 (N_39278,N_37035,N_35694);
and U39279 (N_39279,N_35387,N_37359);
xor U39280 (N_39280,N_36183,N_37318);
nand U39281 (N_39281,N_35995,N_36847);
and U39282 (N_39282,N_37137,N_36814);
xnor U39283 (N_39283,N_36863,N_36794);
xnor U39284 (N_39284,N_36285,N_35023);
xor U39285 (N_39285,N_36717,N_36016);
nand U39286 (N_39286,N_35386,N_35498);
and U39287 (N_39287,N_36878,N_35179);
nand U39288 (N_39288,N_37202,N_36020);
xnor U39289 (N_39289,N_36670,N_35036);
or U39290 (N_39290,N_36669,N_37005);
and U39291 (N_39291,N_35794,N_36703);
and U39292 (N_39292,N_37278,N_35287);
nor U39293 (N_39293,N_35040,N_36363);
nand U39294 (N_39294,N_36068,N_35101);
and U39295 (N_39295,N_35244,N_36104);
nor U39296 (N_39296,N_35185,N_35066);
nor U39297 (N_39297,N_36184,N_36389);
xor U39298 (N_39298,N_36354,N_37232);
nand U39299 (N_39299,N_35904,N_36004);
xor U39300 (N_39300,N_36186,N_37340);
and U39301 (N_39301,N_37230,N_36095);
xnor U39302 (N_39302,N_35724,N_35271);
or U39303 (N_39303,N_35073,N_35899);
nor U39304 (N_39304,N_35288,N_35465);
nor U39305 (N_39305,N_36145,N_36471);
nand U39306 (N_39306,N_35980,N_35483);
nand U39307 (N_39307,N_35479,N_35331);
and U39308 (N_39308,N_36034,N_36483);
or U39309 (N_39309,N_36767,N_36921);
or U39310 (N_39310,N_36956,N_36282);
xor U39311 (N_39311,N_35222,N_35489);
nor U39312 (N_39312,N_36401,N_36786);
or U39313 (N_39313,N_37293,N_36862);
or U39314 (N_39314,N_37102,N_36219);
or U39315 (N_39315,N_36293,N_35054);
or U39316 (N_39316,N_35683,N_35135);
and U39317 (N_39317,N_35807,N_36068);
xnor U39318 (N_39318,N_36811,N_35687);
nor U39319 (N_39319,N_35673,N_36184);
nor U39320 (N_39320,N_35091,N_35363);
and U39321 (N_39321,N_36282,N_35846);
nor U39322 (N_39322,N_36872,N_36907);
and U39323 (N_39323,N_36756,N_35888);
nand U39324 (N_39324,N_35368,N_37188);
nand U39325 (N_39325,N_35800,N_37052);
and U39326 (N_39326,N_36097,N_36171);
xnor U39327 (N_39327,N_37148,N_36185);
nand U39328 (N_39328,N_36701,N_37415);
nor U39329 (N_39329,N_36329,N_35015);
nor U39330 (N_39330,N_37246,N_35243);
and U39331 (N_39331,N_35385,N_37241);
xor U39332 (N_39332,N_36087,N_36960);
xor U39333 (N_39333,N_35112,N_35035);
nand U39334 (N_39334,N_35226,N_37035);
nor U39335 (N_39335,N_35741,N_35192);
xnor U39336 (N_39336,N_35936,N_36134);
or U39337 (N_39337,N_36854,N_36183);
and U39338 (N_39338,N_36336,N_37355);
and U39339 (N_39339,N_37123,N_35109);
nor U39340 (N_39340,N_36234,N_36931);
and U39341 (N_39341,N_35076,N_35504);
or U39342 (N_39342,N_35046,N_36724);
nand U39343 (N_39343,N_37244,N_37436);
and U39344 (N_39344,N_35806,N_37445);
nor U39345 (N_39345,N_35515,N_35724);
and U39346 (N_39346,N_35240,N_35858);
nand U39347 (N_39347,N_36148,N_35377);
and U39348 (N_39348,N_35467,N_36086);
or U39349 (N_39349,N_35299,N_36639);
xor U39350 (N_39350,N_35964,N_36563);
xnor U39351 (N_39351,N_35031,N_37378);
or U39352 (N_39352,N_35008,N_35785);
xor U39353 (N_39353,N_35217,N_36752);
xor U39354 (N_39354,N_35565,N_36516);
nor U39355 (N_39355,N_37256,N_35312);
nand U39356 (N_39356,N_37384,N_36969);
nor U39357 (N_39357,N_36826,N_36392);
nor U39358 (N_39358,N_37319,N_35299);
and U39359 (N_39359,N_36237,N_36893);
xor U39360 (N_39360,N_35028,N_36039);
nor U39361 (N_39361,N_37236,N_36091);
nand U39362 (N_39362,N_37012,N_36169);
and U39363 (N_39363,N_37005,N_35162);
nand U39364 (N_39364,N_36813,N_36106);
nor U39365 (N_39365,N_36025,N_35173);
or U39366 (N_39366,N_35566,N_36531);
xor U39367 (N_39367,N_35783,N_36114);
or U39368 (N_39368,N_36877,N_36650);
and U39369 (N_39369,N_35404,N_35685);
or U39370 (N_39370,N_35131,N_36032);
nand U39371 (N_39371,N_35780,N_36171);
nor U39372 (N_39372,N_35411,N_35368);
or U39373 (N_39373,N_36357,N_36978);
nand U39374 (N_39374,N_36835,N_35797);
and U39375 (N_39375,N_35611,N_37422);
xor U39376 (N_39376,N_35870,N_36179);
or U39377 (N_39377,N_36496,N_36692);
nor U39378 (N_39378,N_37238,N_37315);
nand U39379 (N_39379,N_37169,N_35265);
xor U39380 (N_39380,N_36230,N_36808);
or U39381 (N_39381,N_36640,N_37186);
and U39382 (N_39382,N_36767,N_35011);
nand U39383 (N_39383,N_35234,N_37167);
and U39384 (N_39384,N_37477,N_35635);
or U39385 (N_39385,N_36352,N_37439);
nand U39386 (N_39386,N_37091,N_37119);
xnor U39387 (N_39387,N_36496,N_35600);
and U39388 (N_39388,N_36396,N_36603);
nor U39389 (N_39389,N_36839,N_35207);
and U39390 (N_39390,N_36625,N_37033);
nor U39391 (N_39391,N_37322,N_35639);
and U39392 (N_39392,N_36446,N_37329);
xnor U39393 (N_39393,N_37139,N_35830);
nor U39394 (N_39394,N_36560,N_35625);
nor U39395 (N_39395,N_35827,N_35882);
nand U39396 (N_39396,N_35839,N_36139);
and U39397 (N_39397,N_37448,N_36159);
and U39398 (N_39398,N_36069,N_37047);
or U39399 (N_39399,N_37100,N_35842);
xor U39400 (N_39400,N_36544,N_36603);
nand U39401 (N_39401,N_36398,N_37384);
or U39402 (N_39402,N_35142,N_37173);
xnor U39403 (N_39403,N_36806,N_36254);
nand U39404 (N_39404,N_35665,N_36595);
or U39405 (N_39405,N_35194,N_36979);
xnor U39406 (N_39406,N_36264,N_36559);
nand U39407 (N_39407,N_36507,N_37162);
and U39408 (N_39408,N_35440,N_35075);
xor U39409 (N_39409,N_35018,N_36605);
or U39410 (N_39410,N_35743,N_35547);
or U39411 (N_39411,N_36709,N_36199);
nand U39412 (N_39412,N_36658,N_36839);
or U39413 (N_39413,N_36720,N_36214);
nand U39414 (N_39414,N_37298,N_36600);
and U39415 (N_39415,N_35388,N_35575);
nand U39416 (N_39416,N_35240,N_36791);
xor U39417 (N_39417,N_35899,N_35105);
or U39418 (N_39418,N_36191,N_36486);
nor U39419 (N_39419,N_35652,N_35270);
xor U39420 (N_39420,N_36882,N_35840);
or U39421 (N_39421,N_36747,N_37041);
nand U39422 (N_39422,N_36743,N_35928);
nor U39423 (N_39423,N_36744,N_36519);
or U39424 (N_39424,N_36027,N_36279);
or U39425 (N_39425,N_35561,N_35296);
nand U39426 (N_39426,N_35116,N_35682);
nand U39427 (N_39427,N_35941,N_36287);
nand U39428 (N_39428,N_36698,N_37109);
and U39429 (N_39429,N_35452,N_35685);
nand U39430 (N_39430,N_37156,N_35961);
nand U39431 (N_39431,N_35674,N_35070);
or U39432 (N_39432,N_36346,N_35906);
nor U39433 (N_39433,N_37188,N_35389);
nand U39434 (N_39434,N_37014,N_35944);
and U39435 (N_39435,N_35114,N_37003);
and U39436 (N_39436,N_36245,N_35338);
or U39437 (N_39437,N_35577,N_37182);
nand U39438 (N_39438,N_36545,N_35566);
or U39439 (N_39439,N_35554,N_35216);
or U39440 (N_39440,N_37289,N_37310);
and U39441 (N_39441,N_37059,N_35875);
nor U39442 (N_39442,N_36992,N_37133);
nor U39443 (N_39443,N_35105,N_35233);
or U39444 (N_39444,N_36325,N_36283);
nand U39445 (N_39445,N_36629,N_36188);
nor U39446 (N_39446,N_35155,N_36110);
and U39447 (N_39447,N_35879,N_37414);
xnor U39448 (N_39448,N_36411,N_37249);
or U39449 (N_39449,N_36763,N_37073);
xnor U39450 (N_39450,N_35197,N_35478);
nor U39451 (N_39451,N_35245,N_35959);
and U39452 (N_39452,N_35481,N_37022);
nor U39453 (N_39453,N_36466,N_35847);
nand U39454 (N_39454,N_36298,N_35320);
xnor U39455 (N_39455,N_37166,N_35644);
and U39456 (N_39456,N_36761,N_36188);
xnor U39457 (N_39457,N_35524,N_35188);
nand U39458 (N_39458,N_37158,N_37157);
nor U39459 (N_39459,N_36763,N_35928);
nand U39460 (N_39460,N_36548,N_37048);
or U39461 (N_39461,N_36200,N_35258);
nor U39462 (N_39462,N_35773,N_37398);
nor U39463 (N_39463,N_36185,N_36194);
xor U39464 (N_39464,N_35773,N_36396);
or U39465 (N_39465,N_35041,N_36146);
and U39466 (N_39466,N_35994,N_36932);
nand U39467 (N_39467,N_36000,N_36424);
or U39468 (N_39468,N_37496,N_35184);
and U39469 (N_39469,N_37086,N_36744);
or U39470 (N_39470,N_35298,N_36632);
nor U39471 (N_39471,N_35167,N_37093);
xor U39472 (N_39472,N_36010,N_37161);
and U39473 (N_39473,N_36341,N_35799);
nand U39474 (N_39474,N_36193,N_37372);
and U39475 (N_39475,N_35855,N_36204);
and U39476 (N_39476,N_35391,N_36949);
and U39477 (N_39477,N_36380,N_35598);
or U39478 (N_39478,N_36728,N_35231);
nor U39479 (N_39479,N_35960,N_35636);
nor U39480 (N_39480,N_35220,N_36888);
and U39481 (N_39481,N_36435,N_35415);
or U39482 (N_39482,N_36622,N_36480);
nand U39483 (N_39483,N_36802,N_35935);
nor U39484 (N_39484,N_36708,N_36478);
and U39485 (N_39485,N_35411,N_36017);
nand U39486 (N_39486,N_36745,N_37166);
xor U39487 (N_39487,N_37356,N_35222);
nand U39488 (N_39488,N_35267,N_36535);
or U39489 (N_39489,N_37072,N_36192);
or U39490 (N_39490,N_36384,N_37173);
nor U39491 (N_39491,N_36986,N_35842);
and U39492 (N_39492,N_36632,N_36152);
nand U39493 (N_39493,N_35974,N_36465);
xnor U39494 (N_39494,N_37330,N_35585);
nor U39495 (N_39495,N_35481,N_35505);
or U39496 (N_39496,N_35364,N_35041);
or U39497 (N_39497,N_36878,N_35484);
or U39498 (N_39498,N_36155,N_35785);
nor U39499 (N_39499,N_35446,N_35834);
xor U39500 (N_39500,N_35255,N_35665);
or U39501 (N_39501,N_36097,N_36292);
xnor U39502 (N_39502,N_35300,N_36583);
nor U39503 (N_39503,N_35178,N_35688);
nand U39504 (N_39504,N_36035,N_35089);
xnor U39505 (N_39505,N_36770,N_36637);
nor U39506 (N_39506,N_35216,N_37097);
or U39507 (N_39507,N_35643,N_36253);
and U39508 (N_39508,N_36070,N_36683);
nand U39509 (N_39509,N_35423,N_37423);
nand U39510 (N_39510,N_35500,N_37403);
nor U39511 (N_39511,N_35013,N_35655);
nor U39512 (N_39512,N_35032,N_35940);
nor U39513 (N_39513,N_36529,N_35343);
xor U39514 (N_39514,N_37229,N_37113);
nor U39515 (N_39515,N_35872,N_37262);
nor U39516 (N_39516,N_36007,N_37227);
nand U39517 (N_39517,N_35501,N_37109);
and U39518 (N_39518,N_37486,N_36343);
nand U39519 (N_39519,N_36964,N_35097);
or U39520 (N_39520,N_35293,N_37266);
nor U39521 (N_39521,N_36639,N_35910);
nor U39522 (N_39522,N_36366,N_36764);
xnor U39523 (N_39523,N_36272,N_37178);
or U39524 (N_39524,N_37432,N_35003);
nand U39525 (N_39525,N_36509,N_35699);
xnor U39526 (N_39526,N_36143,N_35200);
or U39527 (N_39527,N_35750,N_36749);
xor U39528 (N_39528,N_35036,N_35204);
or U39529 (N_39529,N_36941,N_37117);
xor U39530 (N_39530,N_36682,N_36507);
nor U39531 (N_39531,N_37331,N_36330);
nor U39532 (N_39532,N_36534,N_35297);
nor U39533 (N_39533,N_37241,N_35496);
or U39534 (N_39534,N_37460,N_36252);
xnor U39535 (N_39535,N_36003,N_36983);
and U39536 (N_39536,N_36536,N_35735);
nor U39537 (N_39537,N_37206,N_37184);
and U39538 (N_39538,N_36569,N_37295);
and U39539 (N_39539,N_35317,N_35716);
nand U39540 (N_39540,N_35631,N_36621);
or U39541 (N_39541,N_37418,N_36216);
nand U39542 (N_39542,N_35655,N_35726);
nor U39543 (N_39543,N_35258,N_35513);
or U39544 (N_39544,N_35066,N_35599);
nor U39545 (N_39545,N_36300,N_37024);
nor U39546 (N_39546,N_35392,N_37257);
and U39547 (N_39547,N_37007,N_36058);
nor U39548 (N_39548,N_36086,N_37231);
or U39549 (N_39549,N_35690,N_35682);
or U39550 (N_39550,N_35227,N_37127);
nor U39551 (N_39551,N_35052,N_37415);
xor U39552 (N_39552,N_35084,N_35715);
xnor U39553 (N_39553,N_37466,N_35957);
and U39554 (N_39554,N_36801,N_36401);
or U39555 (N_39555,N_35693,N_37067);
nor U39556 (N_39556,N_35551,N_36101);
nand U39557 (N_39557,N_35195,N_37474);
nand U39558 (N_39558,N_35230,N_35876);
nor U39559 (N_39559,N_36281,N_35128);
nor U39560 (N_39560,N_36771,N_35930);
xnor U39561 (N_39561,N_36746,N_36921);
xnor U39562 (N_39562,N_36233,N_37383);
nand U39563 (N_39563,N_36486,N_36164);
nor U39564 (N_39564,N_36180,N_36120);
xnor U39565 (N_39565,N_36594,N_35901);
xnor U39566 (N_39566,N_35038,N_37408);
and U39567 (N_39567,N_36938,N_36684);
xor U39568 (N_39568,N_36792,N_35073);
nor U39569 (N_39569,N_36507,N_35113);
nor U39570 (N_39570,N_36300,N_35901);
nor U39571 (N_39571,N_37204,N_35492);
or U39572 (N_39572,N_36583,N_36981);
or U39573 (N_39573,N_35849,N_35162);
and U39574 (N_39574,N_35223,N_36898);
or U39575 (N_39575,N_35237,N_36289);
nand U39576 (N_39576,N_37296,N_36499);
xnor U39577 (N_39577,N_37260,N_35992);
nor U39578 (N_39578,N_36406,N_36641);
and U39579 (N_39579,N_35999,N_36580);
and U39580 (N_39580,N_35434,N_36146);
and U39581 (N_39581,N_35755,N_35103);
nor U39582 (N_39582,N_35862,N_37433);
nand U39583 (N_39583,N_35120,N_37363);
or U39584 (N_39584,N_36181,N_35191);
and U39585 (N_39585,N_36101,N_36815);
xor U39586 (N_39586,N_35498,N_36795);
and U39587 (N_39587,N_37189,N_36878);
xor U39588 (N_39588,N_37419,N_35810);
nand U39589 (N_39589,N_35584,N_35496);
xor U39590 (N_39590,N_37129,N_35260);
nor U39591 (N_39591,N_36193,N_36674);
and U39592 (N_39592,N_36801,N_35025);
nand U39593 (N_39593,N_37409,N_37273);
nor U39594 (N_39594,N_36157,N_36785);
and U39595 (N_39595,N_37331,N_36572);
xnor U39596 (N_39596,N_35296,N_36285);
or U39597 (N_39597,N_37173,N_36657);
xor U39598 (N_39598,N_37006,N_35678);
or U39599 (N_39599,N_36129,N_36847);
xnor U39600 (N_39600,N_35605,N_35681);
nor U39601 (N_39601,N_36205,N_36725);
and U39602 (N_39602,N_35059,N_37112);
nand U39603 (N_39603,N_36850,N_35998);
and U39604 (N_39604,N_35297,N_37356);
and U39605 (N_39605,N_35135,N_35214);
nor U39606 (N_39606,N_36864,N_35147);
and U39607 (N_39607,N_35894,N_36515);
and U39608 (N_39608,N_36145,N_35172);
and U39609 (N_39609,N_37223,N_35024);
and U39610 (N_39610,N_37250,N_35321);
and U39611 (N_39611,N_37403,N_36917);
and U39612 (N_39612,N_35071,N_35424);
nand U39613 (N_39613,N_36969,N_36060);
xnor U39614 (N_39614,N_36986,N_36031);
or U39615 (N_39615,N_37158,N_36096);
nand U39616 (N_39616,N_35316,N_35921);
nor U39617 (N_39617,N_36244,N_36396);
and U39618 (N_39618,N_36476,N_36604);
nor U39619 (N_39619,N_35924,N_36265);
nand U39620 (N_39620,N_36811,N_37268);
xor U39621 (N_39621,N_36707,N_35902);
or U39622 (N_39622,N_35658,N_36529);
xor U39623 (N_39623,N_35574,N_35212);
nand U39624 (N_39624,N_35955,N_35427);
or U39625 (N_39625,N_36819,N_36761);
nor U39626 (N_39626,N_35540,N_36384);
xor U39627 (N_39627,N_36845,N_36517);
xnor U39628 (N_39628,N_35870,N_37243);
or U39629 (N_39629,N_36172,N_35578);
and U39630 (N_39630,N_36026,N_35135);
or U39631 (N_39631,N_36567,N_37296);
and U39632 (N_39632,N_37445,N_35647);
nand U39633 (N_39633,N_37150,N_36929);
or U39634 (N_39634,N_37257,N_37067);
and U39635 (N_39635,N_36156,N_36254);
or U39636 (N_39636,N_37418,N_35274);
xnor U39637 (N_39637,N_36336,N_35618);
nor U39638 (N_39638,N_36396,N_36010);
nand U39639 (N_39639,N_36559,N_35601);
nand U39640 (N_39640,N_35627,N_37025);
nor U39641 (N_39641,N_36869,N_35203);
nor U39642 (N_39642,N_37167,N_36281);
nand U39643 (N_39643,N_36443,N_35801);
nor U39644 (N_39644,N_36180,N_35307);
xor U39645 (N_39645,N_37176,N_35324);
nand U39646 (N_39646,N_36065,N_35992);
or U39647 (N_39647,N_37245,N_37109);
nand U39648 (N_39648,N_36781,N_36827);
nor U39649 (N_39649,N_36276,N_37469);
and U39650 (N_39650,N_37112,N_37043);
nor U39651 (N_39651,N_36578,N_37241);
nand U39652 (N_39652,N_35667,N_35046);
or U39653 (N_39653,N_36071,N_36527);
and U39654 (N_39654,N_36078,N_37332);
and U39655 (N_39655,N_36960,N_37058);
nor U39656 (N_39656,N_35047,N_36142);
xnor U39657 (N_39657,N_35942,N_36021);
xnor U39658 (N_39658,N_35398,N_35325);
and U39659 (N_39659,N_36765,N_36898);
nand U39660 (N_39660,N_35696,N_36834);
and U39661 (N_39661,N_35313,N_37034);
xor U39662 (N_39662,N_36990,N_36383);
nor U39663 (N_39663,N_36683,N_35222);
xor U39664 (N_39664,N_35486,N_35464);
xor U39665 (N_39665,N_35525,N_35813);
xor U39666 (N_39666,N_36970,N_36466);
xor U39667 (N_39667,N_35783,N_37477);
nor U39668 (N_39668,N_35390,N_35141);
or U39669 (N_39669,N_37328,N_35401);
and U39670 (N_39670,N_35099,N_35238);
nand U39671 (N_39671,N_35901,N_36428);
xor U39672 (N_39672,N_37191,N_36395);
or U39673 (N_39673,N_37256,N_37166);
or U39674 (N_39674,N_36664,N_37122);
nor U39675 (N_39675,N_35975,N_37387);
or U39676 (N_39676,N_37091,N_36212);
nor U39677 (N_39677,N_36455,N_36381);
and U39678 (N_39678,N_35945,N_35022);
nand U39679 (N_39679,N_35414,N_37073);
and U39680 (N_39680,N_35877,N_35164);
or U39681 (N_39681,N_36311,N_36039);
xor U39682 (N_39682,N_35232,N_35214);
and U39683 (N_39683,N_35328,N_36033);
and U39684 (N_39684,N_35499,N_35623);
or U39685 (N_39685,N_36931,N_35400);
xnor U39686 (N_39686,N_37369,N_35800);
or U39687 (N_39687,N_35615,N_36765);
xnor U39688 (N_39688,N_35034,N_36162);
xnor U39689 (N_39689,N_35328,N_35624);
or U39690 (N_39690,N_36769,N_35984);
and U39691 (N_39691,N_36275,N_36873);
nor U39692 (N_39692,N_35658,N_35239);
and U39693 (N_39693,N_36849,N_35460);
nor U39694 (N_39694,N_35160,N_37185);
xor U39695 (N_39695,N_36565,N_37279);
nand U39696 (N_39696,N_35287,N_35614);
and U39697 (N_39697,N_35234,N_37276);
and U39698 (N_39698,N_35194,N_36518);
and U39699 (N_39699,N_35009,N_36358);
or U39700 (N_39700,N_36219,N_36482);
nor U39701 (N_39701,N_35238,N_35373);
or U39702 (N_39702,N_36896,N_37323);
nor U39703 (N_39703,N_36083,N_36484);
or U39704 (N_39704,N_36645,N_35378);
or U39705 (N_39705,N_35160,N_35281);
and U39706 (N_39706,N_35366,N_35664);
nor U39707 (N_39707,N_35450,N_36047);
xnor U39708 (N_39708,N_36814,N_36101);
xnor U39709 (N_39709,N_37079,N_35283);
or U39710 (N_39710,N_37047,N_36946);
nand U39711 (N_39711,N_35937,N_37080);
nand U39712 (N_39712,N_36355,N_36959);
xor U39713 (N_39713,N_35428,N_36423);
nand U39714 (N_39714,N_35631,N_36160);
or U39715 (N_39715,N_36011,N_35627);
or U39716 (N_39716,N_35292,N_36508);
xor U39717 (N_39717,N_37041,N_36216);
or U39718 (N_39718,N_35861,N_35521);
xnor U39719 (N_39719,N_35568,N_36043);
nand U39720 (N_39720,N_37146,N_35817);
nand U39721 (N_39721,N_35044,N_36593);
xnor U39722 (N_39722,N_37221,N_37318);
xor U39723 (N_39723,N_35973,N_36292);
xnor U39724 (N_39724,N_35959,N_35794);
and U39725 (N_39725,N_35540,N_37371);
or U39726 (N_39726,N_36715,N_37176);
nor U39727 (N_39727,N_36445,N_36972);
xnor U39728 (N_39728,N_36767,N_35289);
nor U39729 (N_39729,N_36819,N_37492);
and U39730 (N_39730,N_35740,N_37025);
nand U39731 (N_39731,N_35592,N_35269);
or U39732 (N_39732,N_35143,N_35935);
nand U39733 (N_39733,N_36630,N_35783);
and U39734 (N_39734,N_36977,N_36935);
and U39735 (N_39735,N_36375,N_35626);
xor U39736 (N_39736,N_35417,N_35462);
nand U39737 (N_39737,N_36852,N_35174);
nor U39738 (N_39738,N_36083,N_35164);
or U39739 (N_39739,N_36464,N_35955);
nor U39740 (N_39740,N_36659,N_36812);
nor U39741 (N_39741,N_35251,N_36896);
nand U39742 (N_39742,N_35317,N_35433);
and U39743 (N_39743,N_35712,N_36655);
nand U39744 (N_39744,N_37213,N_36735);
and U39745 (N_39745,N_37396,N_35329);
and U39746 (N_39746,N_36270,N_36597);
and U39747 (N_39747,N_36057,N_36342);
or U39748 (N_39748,N_36517,N_36914);
nand U39749 (N_39749,N_35155,N_37255);
or U39750 (N_39750,N_36666,N_37025);
xnor U39751 (N_39751,N_35551,N_36184);
and U39752 (N_39752,N_37088,N_36779);
xor U39753 (N_39753,N_35080,N_37307);
nor U39754 (N_39754,N_37492,N_37458);
nand U39755 (N_39755,N_35905,N_36568);
nor U39756 (N_39756,N_36639,N_36012);
nor U39757 (N_39757,N_35859,N_35086);
and U39758 (N_39758,N_35022,N_37346);
or U39759 (N_39759,N_37416,N_36328);
or U39760 (N_39760,N_36665,N_37190);
and U39761 (N_39761,N_36318,N_35934);
nand U39762 (N_39762,N_37102,N_36520);
nand U39763 (N_39763,N_35071,N_35242);
xor U39764 (N_39764,N_35941,N_37176);
xnor U39765 (N_39765,N_36269,N_37314);
xor U39766 (N_39766,N_35251,N_36378);
xor U39767 (N_39767,N_35942,N_36705);
xor U39768 (N_39768,N_35931,N_35790);
nor U39769 (N_39769,N_35373,N_35388);
nor U39770 (N_39770,N_37145,N_37481);
nand U39771 (N_39771,N_36880,N_35039);
xnor U39772 (N_39772,N_37016,N_37067);
xor U39773 (N_39773,N_35277,N_36642);
nor U39774 (N_39774,N_36527,N_35405);
or U39775 (N_39775,N_37176,N_35257);
or U39776 (N_39776,N_36923,N_37107);
nand U39777 (N_39777,N_36040,N_37343);
xor U39778 (N_39778,N_37409,N_35152);
nand U39779 (N_39779,N_36177,N_37029);
nand U39780 (N_39780,N_37209,N_37255);
xor U39781 (N_39781,N_36611,N_35427);
nor U39782 (N_39782,N_37053,N_36666);
nor U39783 (N_39783,N_35942,N_35026);
nand U39784 (N_39784,N_37076,N_35774);
and U39785 (N_39785,N_37125,N_36153);
and U39786 (N_39786,N_35135,N_36170);
nand U39787 (N_39787,N_37269,N_35210);
and U39788 (N_39788,N_37075,N_35559);
or U39789 (N_39789,N_36173,N_36950);
nor U39790 (N_39790,N_36795,N_37499);
nor U39791 (N_39791,N_35757,N_37288);
and U39792 (N_39792,N_35342,N_35844);
nand U39793 (N_39793,N_37445,N_35283);
and U39794 (N_39794,N_37464,N_36271);
xor U39795 (N_39795,N_36117,N_37489);
and U39796 (N_39796,N_36231,N_36854);
nand U39797 (N_39797,N_37264,N_36801);
or U39798 (N_39798,N_36833,N_36016);
xnor U39799 (N_39799,N_36079,N_37208);
and U39800 (N_39800,N_37027,N_36345);
nor U39801 (N_39801,N_35515,N_37050);
nor U39802 (N_39802,N_36430,N_35846);
xor U39803 (N_39803,N_37336,N_37040);
nand U39804 (N_39804,N_35022,N_35854);
xnor U39805 (N_39805,N_35044,N_36419);
xnor U39806 (N_39806,N_35289,N_35002);
or U39807 (N_39807,N_36072,N_36498);
or U39808 (N_39808,N_37190,N_35197);
nor U39809 (N_39809,N_37170,N_35351);
or U39810 (N_39810,N_35578,N_37114);
nor U39811 (N_39811,N_35169,N_35355);
or U39812 (N_39812,N_37040,N_36933);
and U39813 (N_39813,N_37141,N_37459);
or U39814 (N_39814,N_36878,N_37014);
xnor U39815 (N_39815,N_36961,N_35985);
and U39816 (N_39816,N_35880,N_37115);
nand U39817 (N_39817,N_35397,N_35323);
nor U39818 (N_39818,N_35231,N_35761);
nand U39819 (N_39819,N_37473,N_35071);
xor U39820 (N_39820,N_36691,N_36730);
and U39821 (N_39821,N_36170,N_35102);
or U39822 (N_39822,N_37247,N_35344);
and U39823 (N_39823,N_35390,N_37153);
nand U39824 (N_39824,N_36498,N_36754);
or U39825 (N_39825,N_36573,N_36399);
and U39826 (N_39826,N_35029,N_36340);
xnor U39827 (N_39827,N_37122,N_35768);
nor U39828 (N_39828,N_37391,N_35570);
nand U39829 (N_39829,N_37011,N_36483);
nand U39830 (N_39830,N_35178,N_36938);
xnor U39831 (N_39831,N_35361,N_36539);
xnor U39832 (N_39832,N_36387,N_36994);
xor U39833 (N_39833,N_37287,N_36240);
nand U39834 (N_39834,N_35880,N_36208);
and U39835 (N_39835,N_36458,N_35658);
nor U39836 (N_39836,N_36650,N_37271);
and U39837 (N_39837,N_36588,N_35897);
or U39838 (N_39838,N_35635,N_36941);
nor U39839 (N_39839,N_35649,N_36372);
xnor U39840 (N_39840,N_35045,N_36164);
nor U39841 (N_39841,N_37030,N_35460);
nand U39842 (N_39842,N_37114,N_35728);
or U39843 (N_39843,N_35238,N_37357);
nor U39844 (N_39844,N_35642,N_37459);
xnor U39845 (N_39845,N_35626,N_36031);
or U39846 (N_39846,N_36661,N_35069);
and U39847 (N_39847,N_36889,N_35421);
xnor U39848 (N_39848,N_37438,N_35038);
or U39849 (N_39849,N_37302,N_35383);
nand U39850 (N_39850,N_35261,N_35102);
nor U39851 (N_39851,N_35323,N_36721);
nor U39852 (N_39852,N_36588,N_35403);
nand U39853 (N_39853,N_36418,N_35589);
xor U39854 (N_39854,N_37102,N_36079);
and U39855 (N_39855,N_36070,N_35935);
xnor U39856 (N_39856,N_36854,N_36803);
nor U39857 (N_39857,N_35835,N_37207);
nand U39858 (N_39858,N_36944,N_35504);
nand U39859 (N_39859,N_36359,N_35692);
nand U39860 (N_39860,N_36231,N_37055);
and U39861 (N_39861,N_36126,N_35159);
or U39862 (N_39862,N_36120,N_36252);
xnor U39863 (N_39863,N_37076,N_36529);
and U39864 (N_39864,N_35959,N_35746);
nor U39865 (N_39865,N_35194,N_35505);
xnor U39866 (N_39866,N_36332,N_36962);
nor U39867 (N_39867,N_35015,N_36336);
or U39868 (N_39868,N_35361,N_35514);
nand U39869 (N_39869,N_36518,N_35997);
and U39870 (N_39870,N_37425,N_35100);
nand U39871 (N_39871,N_37463,N_36991);
nand U39872 (N_39872,N_35296,N_36060);
nand U39873 (N_39873,N_36689,N_37260);
nand U39874 (N_39874,N_37164,N_36036);
and U39875 (N_39875,N_36169,N_35595);
and U39876 (N_39876,N_36540,N_36251);
xnor U39877 (N_39877,N_35343,N_36687);
or U39878 (N_39878,N_35758,N_36936);
nor U39879 (N_39879,N_36906,N_35743);
nand U39880 (N_39880,N_37412,N_37368);
nand U39881 (N_39881,N_36033,N_35026);
xor U39882 (N_39882,N_36074,N_35998);
and U39883 (N_39883,N_35818,N_36122);
nand U39884 (N_39884,N_36825,N_36847);
nor U39885 (N_39885,N_35251,N_36303);
nand U39886 (N_39886,N_35108,N_35919);
or U39887 (N_39887,N_37457,N_35417);
nand U39888 (N_39888,N_36624,N_37348);
or U39889 (N_39889,N_36695,N_35881);
or U39890 (N_39890,N_36718,N_35451);
nand U39891 (N_39891,N_35591,N_35666);
xor U39892 (N_39892,N_35081,N_36659);
nand U39893 (N_39893,N_37049,N_36962);
nand U39894 (N_39894,N_35803,N_36912);
or U39895 (N_39895,N_37103,N_36253);
nor U39896 (N_39896,N_36197,N_36147);
xnor U39897 (N_39897,N_36982,N_35470);
nor U39898 (N_39898,N_35632,N_36254);
or U39899 (N_39899,N_35534,N_36964);
or U39900 (N_39900,N_35653,N_35499);
and U39901 (N_39901,N_35375,N_35345);
xor U39902 (N_39902,N_36486,N_37194);
nor U39903 (N_39903,N_36212,N_35872);
nand U39904 (N_39904,N_36036,N_35122);
nand U39905 (N_39905,N_35111,N_36744);
or U39906 (N_39906,N_36583,N_35129);
nand U39907 (N_39907,N_36874,N_35504);
or U39908 (N_39908,N_35519,N_36652);
nor U39909 (N_39909,N_37380,N_35478);
and U39910 (N_39910,N_35827,N_37478);
nor U39911 (N_39911,N_36219,N_35511);
or U39912 (N_39912,N_37093,N_37351);
nand U39913 (N_39913,N_36302,N_35331);
nor U39914 (N_39914,N_35444,N_37284);
xor U39915 (N_39915,N_35163,N_37011);
nand U39916 (N_39916,N_35204,N_36805);
or U39917 (N_39917,N_35211,N_37415);
xnor U39918 (N_39918,N_35727,N_35233);
nor U39919 (N_39919,N_36172,N_35330);
nand U39920 (N_39920,N_35933,N_36938);
and U39921 (N_39921,N_36328,N_35332);
nand U39922 (N_39922,N_37452,N_37329);
nor U39923 (N_39923,N_35891,N_37446);
or U39924 (N_39924,N_36098,N_36661);
or U39925 (N_39925,N_35274,N_35382);
and U39926 (N_39926,N_36686,N_37386);
and U39927 (N_39927,N_37326,N_35597);
or U39928 (N_39928,N_35708,N_35661);
or U39929 (N_39929,N_36093,N_35573);
xor U39930 (N_39930,N_35155,N_37290);
or U39931 (N_39931,N_37475,N_35449);
nor U39932 (N_39932,N_36313,N_37216);
xor U39933 (N_39933,N_35212,N_36534);
nor U39934 (N_39934,N_36555,N_37438);
and U39935 (N_39935,N_35283,N_35931);
nand U39936 (N_39936,N_36666,N_37454);
and U39937 (N_39937,N_37060,N_35374);
xor U39938 (N_39938,N_37123,N_37312);
nand U39939 (N_39939,N_35819,N_35425);
and U39940 (N_39940,N_35355,N_36299);
nand U39941 (N_39941,N_37193,N_37062);
xnor U39942 (N_39942,N_37015,N_35036);
or U39943 (N_39943,N_35258,N_36024);
or U39944 (N_39944,N_35874,N_35612);
xnor U39945 (N_39945,N_37330,N_37228);
and U39946 (N_39946,N_35563,N_35143);
or U39947 (N_39947,N_36251,N_35564);
xnor U39948 (N_39948,N_35619,N_36573);
and U39949 (N_39949,N_35167,N_35154);
or U39950 (N_39950,N_36243,N_35784);
xor U39951 (N_39951,N_37107,N_36413);
or U39952 (N_39952,N_35056,N_35378);
nand U39953 (N_39953,N_36365,N_36285);
and U39954 (N_39954,N_36659,N_35163);
nor U39955 (N_39955,N_36705,N_35851);
and U39956 (N_39956,N_35659,N_36986);
or U39957 (N_39957,N_36666,N_35541);
nand U39958 (N_39958,N_35776,N_35724);
or U39959 (N_39959,N_35439,N_36815);
nand U39960 (N_39960,N_35838,N_35859);
nor U39961 (N_39961,N_36602,N_36472);
xnor U39962 (N_39962,N_36121,N_36474);
or U39963 (N_39963,N_35718,N_35183);
or U39964 (N_39964,N_35492,N_35830);
nand U39965 (N_39965,N_37205,N_35740);
nand U39966 (N_39966,N_37162,N_36173);
xor U39967 (N_39967,N_35165,N_37121);
nand U39968 (N_39968,N_35914,N_37420);
xnor U39969 (N_39969,N_35901,N_36830);
nand U39970 (N_39970,N_36420,N_37357);
and U39971 (N_39971,N_35576,N_36268);
and U39972 (N_39972,N_36289,N_35004);
or U39973 (N_39973,N_35481,N_35746);
xnor U39974 (N_39974,N_36200,N_36793);
nand U39975 (N_39975,N_36864,N_36331);
nor U39976 (N_39976,N_35359,N_37351);
and U39977 (N_39977,N_35352,N_37322);
or U39978 (N_39978,N_35235,N_37030);
and U39979 (N_39979,N_35733,N_36309);
and U39980 (N_39980,N_36278,N_36946);
or U39981 (N_39981,N_35017,N_35849);
xor U39982 (N_39982,N_35001,N_37105);
and U39983 (N_39983,N_37180,N_35469);
or U39984 (N_39984,N_35415,N_37440);
xnor U39985 (N_39985,N_35537,N_37483);
xnor U39986 (N_39986,N_35472,N_37299);
or U39987 (N_39987,N_36427,N_36588);
and U39988 (N_39988,N_35956,N_35601);
xor U39989 (N_39989,N_37383,N_37142);
and U39990 (N_39990,N_36853,N_36924);
and U39991 (N_39991,N_37338,N_37333);
nand U39992 (N_39992,N_36990,N_35541);
xor U39993 (N_39993,N_35547,N_36084);
and U39994 (N_39994,N_35083,N_36649);
xnor U39995 (N_39995,N_35249,N_36087);
and U39996 (N_39996,N_35026,N_37287);
nand U39997 (N_39997,N_35826,N_36382);
xor U39998 (N_39998,N_36075,N_35719);
nand U39999 (N_39999,N_35821,N_35151);
and U40000 (N_40000,N_38966,N_38193);
xor U40001 (N_40001,N_37815,N_38080);
or U40002 (N_40002,N_38187,N_38663);
nand U40003 (N_40003,N_38765,N_38030);
nand U40004 (N_40004,N_38308,N_38880);
and U40005 (N_40005,N_39133,N_37677);
nand U40006 (N_40006,N_38550,N_39011);
nor U40007 (N_40007,N_38725,N_39813);
nand U40008 (N_40008,N_38428,N_39985);
nand U40009 (N_40009,N_39948,N_38841);
or U40010 (N_40010,N_39470,N_39931);
or U40011 (N_40011,N_37638,N_39201);
or U40012 (N_40012,N_38331,N_37977);
or U40013 (N_40013,N_37981,N_38120);
nor U40014 (N_40014,N_38695,N_38934);
nor U40015 (N_40015,N_38319,N_38954);
and U40016 (N_40016,N_37788,N_38038);
and U40017 (N_40017,N_38090,N_38026);
or U40018 (N_40018,N_38031,N_38562);
nand U40019 (N_40019,N_39112,N_37812);
or U40020 (N_40020,N_39146,N_37530);
or U40021 (N_40021,N_37560,N_39473);
and U40022 (N_40022,N_39387,N_38497);
xor U40023 (N_40023,N_37880,N_39062);
nor U40024 (N_40024,N_38449,N_37776);
nor U40025 (N_40025,N_39632,N_38226);
xnor U40026 (N_40026,N_39800,N_37564);
nor U40027 (N_40027,N_39194,N_38472);
xor U40028 (N_40028,N_37970,N_39132);
or U40029 (N_40029,N_39452,N_39450);
nor U40030 (N_40030,N_39501,N_37831);
xor U40031 (N_40031,N_37646,N_39270);
or U40032 (N_40032,N_39301,N_38404);
or U40033 (N_40033,N_38859,N_38672);
xor U40034 (N_40034,N_38526,N_39822);
and U40035 (N_40035,N_39268,N_38718);
or U40036 (N_40036,N_37605,N_38864);
nor U40037 (N_40037,N_38680,N_38789);
xnor U40038 (N_40038,N_39588,N_39811);
nor U40039 (N_40039,N_38877,N_37935);
nand U40040 (N_40040,N_38250,N_37541);
and U40041 (N_40041,N_38588,N_37660);
xnor U40042 (N_40042,N_39593,N_39430);
and U40043 (N_40043,N_38816,N_38557);
and U40044 (N_40044,N_39656,N_39866);
nor U40045 (N_40045,N_39373,N_38612);
nor U40046 (N_40046,N_38028,N_38796);
or U40047 (N_40047,N_39255,N_39644);
or U40048 (N_40048,N_37549,N_39873);
nand U40049 (N_40049,N_38502,N_38742);
xor U40050 (N_40050,N_39143,N_39190);
and U40051 (N_40051,N_39758,N_38848);
or U40052 (N_40052,N_38068,N_38256);
xnor U40053 (N_40053,N_37714,N_37681);
or U40054 (N_40054,N_38884,N_38128);
nand U40055 (N_40055,N_38721,N_39668);
nor U40056 (N_40056,N_37552,N_37915);
nor U40057 (N_40057,N_39429,N_39377);
xor U40058 (N_40058,N_38434,N_39486);
nor U40059 (N_40059,N_37958,N_38282);
xnor U40060 (N_40060,N_38362,N_39551);
nand U40061 (N_40061,N_39085,N_38854);
nor U40062 (N_40062,N_38437,N_39174);
and U40063 (N_40063,N_38813,N_38543);
nand U40064 (N_40064,N_38525,N_37898);
or U40065 (N_40065,N_38286,N_37548);
nand U40066 (N_40066,N_39565,N_38961);
nor U40067 (N_40067,N_39530,N_39349);
nand U40068 (N_40068,N_39363,N_37697);
and U40069 (N_40069,N_39582,N_38211);
xor U40070 (N_40070,N_39111,N_39331);
nand U40071 (N_40071,N_39084,N_38145);
and U40072 (N_40072,N_39015,N_38444);
nor U40073 (N_40073,N_37851,N_39445);
nand U40074 (N_40074,N_38684,N_37645);
nand U40075 (N_40075,N_38316,N_38084);
or U40076 (N_40076,N_39858,N_39649);
and U40077 (N_40077,N_38986,N_38755);
nor U40078 (N_40078,N_38743,N_39952);
or U40079 (N_40079,N_37874,N_39755);
nor U40080 (N_40080,N_37855,N_37668);
or U40081 (N_40081,N_39449,N_38981);
nor U40082 (N_40082,N_38803,N_38845);
nor U40083 (N_40083,N_37844,N_39026);
nor U40084 (N_40084,N_37911,N_38091);
and U40085 (N_40085,N_38441,N_38804);
nand U40086 (N_40086,N_38691,N_39369);
xnor U40087 (N_40087,N_39716,N_37651);
nor U40088 (N_40088,N_39217,N_38369);
or U40089 (N_40089,N_38868,N_39919);
nand U40090 (N_40090,N_39825,N_37773);
xnor U40091 (N_40091,N_38486,N_38227);
or U40092 (N_40092,N_37910,N_39667);
xor U40093 (N_40093,N_38446,N_39202);
and U40094 (N_40094,N_38558,N_38930);
and U40095 (N_40095,N_39471,N_39506);
and U40096 (N_40096,N_39910,N_39786);
or U40097 (N_40097,N_39722,N_38949);
or U40098 (N_40098,N_38552,N_38243);
nand U40099 (N_40099,N_37975,N_39809);
and U40100 (N_40100,N_38733,N_37886);
or U40101 (N_40101,N_39864,N_38730);
nand U40102 (N_40102,N_38759,N_37985);
or U40103 (N_40103,N_38198,N_38665);
nor U40104 (N_40104,N_38312,N_37571);
nand U40105 (N_40105,N_37700,N_37518);
and U40106 (N_40106,N_38073,N_37639);
xor U40107 (N_40107,N_39730,N_39658);
and U40108 (N_40108,N_39521,N_39454);
or U40109 (N_40109,N_39078,N_38216);
xor U40110 (N_40110,N_39797,N_38777);
nand U40111 (N_40111,N_39226,N_38944);
xnor U40112 (N_40112,N_38361,N_38522);
and U40113 (N_40113,N_38277,N_39974);
nand U40114 (N_40114,N_39317,N_38548);
nor U40115 (N_40115,N_39478,N_38290);
nor U40116 (N_40116,N_38248,N_39806);
or U40117 (N_40117,N_39046,N_38594);
nor U40118 (N_40118,N_39199,N_37903);
and U40119 (N_40119,N_38592,N_38159);
xor U40120 (N_40120,N_39737,N_38137);
xor U40121 (N_40121,N_39433,N_39110);
and U40122 (N_40122,N_38870,N_37912);
or U40123 (N_40123,N_38093,N_38438);
nand U40124 (N_40124,N_38027,N_38927);
nor U40125 (N_40125,N_38426,N_39292);
and U40126 (N_40126,N_38055,N_38058);
nor U40127 (N_40127,N_39150,N_37735);
nand U40128 (N_40128,N_39930,N_37828);
and U40129 (N_40129,N_39118,N_39594);
and U40130 (N_40130,N_39256,N_38790);
or U40131 (N_40131,N_39945,N_39224);
xnor U40132 (N_40132,N_39036,N_37547);
and U40133 (N_40133,N_38200,N_39872);
and U40134 (N_40134,N_38009,N_38156);
or U40135 (N_40135,N_38511,N_39954);
xor U40136 (N_40136,N_39814,N_37826);
or U40137 (N_40137,N_39849,N_38303);
nor U40138 (N_40138,N_39720,N_37967);
and U40139 (N_40139,N_37705,N_37909);
nand U40140 (N_40140,N_39051,N_38571);
xor U40141 (N_40141,N_38240,N_39525);
nand U40142 (N_40142,N_39340,N_37959);
and U40143 (N_40143,N_39789,N_39048);
nor U40144 (N_40144,N_37919,N_38297);
xor U40145 (N_40145,N_39949,N_38197);
nor U40146 (N_40146,N_39993,N_39803);
nor U40147 (N_40147,N_37782,N_39659);
nor U40148 (N_40148,N_37615,N_37606);
and U40149 (N_40149,N_38766,N_39288);
or U40150 (N_40150,N_39299,N_37557);
xnor U40151 (N_40151,N_38910,N_38062);
or U40152 (N_40152,N_39953,N_39172);
nor U40153 (N_40153,N_38300,N_39741);
or U40154 (N_40154,N_37708,N_37576);
xor U40155 (N_40155,N_38131,N_38991);
nor U40156 (N_40156,N_38064,N_37839);
and U40157 (N_40157,N_39714,N_37584);
nand U40158 (N_40158,N_38349,N_37781);
nand U40159 (N_40159,N_38095,N_38056);
or U40160 (N_40160,N_39176,N_37768);
nand U40161 (N_40161,N_39425,N_37974);
and U40162 (N_40162,N_39390,N_39164);
nor U40163 (N_40163,N_37670,N_39087);
or U40164 (N_40164,N_39337,N_38631);
and U40165 (N_40165,N_38077,N_39837);
nor U40166 (N_40166,N_38435,N_38540);
nor U40167 (N_40167,N_39098,N_39041);
xnor U40168 (N_40168,N_38587,N_39443);
nor U40169 (N_40169,N_38632,N_38768);
or U40170 (N_40170,N_38236,N_38683);
xnor U40171 (N_40171,N_39281,N_37783);
nor U40172 (N_40172,N_37846,N_38810);
and U40173 (N_40173,N_39155,N_38351);
xor U40174 (N_40174,N_38454,N_39596);
nand U40175 (N_40175,N_39855,N_37620);
nand U40176 (N_40176,N_38639,N_38638);
xor U40177 (N_40177,N_37743,N_38387);
and U40178 (N_40178,N_38829,N_38542);
and U40179 (N_40179,N_38086,N_37722);
nand U40180 (N_40180,N_37956,N_39918);
xor U40181 (N_40181,N_39505,N_37515);
nand U40182 (N_40182,N_39453,N_38179);
xor U40183 (N_40183,N_37951,N_39264);
or U40184 (N_40184,N_38258,N_38229);
or U40185 (N_40185,N_37635,N_37865);
or U40186 (N_40186,N_39988,N_39345);
nor U40187 (N_40187,N_37613,N_38141);
nor U40188 (N_40188,N_38218,N_37751);
nor U40189 (N_40189,N_39093,N_37770);
nand U40190 (N_40190,N_39076,N_39014);
nor U40191 (N_40191,N_38190,N_38895);
xor U40192 (N_40192,N_38136,N_39397);
and U40193 (N_40193,N_38726,N_38151);
and U40194 (N_40194,N_38922,N_38067);
xnor U40195 (N_40195,N_39116,N_39294);
or U40196 (N_40196,N_39859,N_38414);
nor U40197 (N_40197,N_39964,N_38205);
or U40198 (N_40198,N_39332,N_38046);
or U40199 (N_40199,N_39179,N_38563);
nor U40200 (N_40200,N_38906,N_38042);
or U40201 (N_40201,N_38310,N_38840);
and U40202 (N_40202,N_39485,N_39065);
nand U40203 (N_40203,N_38629,N_38701);
or U40204 (N_40204,N_38931,N_38161);
nand U40205 (N_40205,N_39560,N_38005);
nor U40206 (N_40206,N_39392,N_39831);
xnor U40207 (N_40207,N_37795,N_38115);
or U40208 (N_40208,N_38057,N_38590);
nand U40209 (N_40209,N_38037,N_37827);
xor U40210 (N_40210,N_39262,N_38419);
and U40211 (N_40211,N_38196,N_38717);
xnor U40212 (N_40212,N_38346,N_38760);
nand U40213 (N_40213,N_37664,N_38424);
or U40214 (N_40214,N_37942,N_39295);
xor U40215 (N_40215,N_39599,N_38500);
nor U40216 (N_40216,N_39017,N_39423);
xnor U40217 (N_40217,N_38280,N_39100);
nor U40218 (N_40218,N_38012,N_37682);
or U40219 (N_40219,N_38754,N_38289);
and U40220 (N_40220,N_38283,N_37864);
and U40221 (N_40221,N_38516,N_37612);
and U40222 (N_40222,N_39689,N_38427);
and U40223 (N_40223,N_37940,N_38202);
xor U40224 (N_40224,N_39520,N_38463);
or U40225 (N_40225,N_37995,N_37580);
xor U40226 (N_40226,N_39258,N_38208);
nor U40227 (N_40227,N_38342,N_39489);
or U40228 (N_40228,N_39372,N_38998);
and U40229 (N_40229,N_38819,N_37748);
or U40230 (N_40230,N_37927,N_37938);
nand U40231 (N_40231,N_39400,N_37845);
nand U40232 (N_40232,N_39573,N_38549);
nor U40233 (N_40233,N_39223,N_39043);
nor U40234 (N_40234,N_39068,N_38014);
or U40235 (N_40235,N_37508,N_39677);
nand U40236 (N_40236,N_37583,N_39214);
nor U40237 (N_40237,N_39526,N_38882);
xor U40238 (N_40238,N_37930,N_37542);
nor U40239 (N_40239,N_37969,N_38116);
nand U40240 (N_40240,N_39519,N_38538);
and U40241 (N_40241,N_38839,N_38178);
nor U40242 (N_40242,N_39069,N_37799);
xnor U40243 (N_40243,N_37961,N_39330);
and U40244 (N_40244,N_37752,N_38809);
and U40245 (N_40245,N_38255,N_38953);
nor U40246 (N_40246,N_39769,N_37611);
nand U40247 (N_40247,N_38746,N_38078);
and U40248 (N_40248,N_38583,N_39399);
nor U40249 (N_40249,N_39559,N_39481);
nand U40250 (N_40250,N_39220,N_37652);
nand U40251 (N_40251,N_37698,N_38339);
xnor U40252 (N_40252,N_38469,N_38398);
nand U40253 (N_40253,N_39420,N_39876);
and U40254 (N_40254,N_37578,N_38475);
and U40255 (N_40255,N_39005,N_38386);
or U40256 (N_40256,N_39760,N_37767);
or U40257 (N_40257,N_39042,N_38977);
and U40258 (N_40258,N_39427,N_39549);
nor U40259 (N_40259,N_38158,N_38626);
xor U40260 (N_40260,N_39839,N_38415);
or U40261 (N_40261,N_38654,N_38293);
and U40262 (N_40262,N_37889,N_37528);
or U40263 (N_40263,N_37993,N_38020);
or U40264 (N_40264,N_38407,N_39793);
nand U40265 (N_40265,N_39894,N_39911);
xor U40266 (N_40266,N_39216,N_37872);
nand U40267 (N_40267,N_37502,N_39302);
and U40268 (N_40268,N_38430,N_39462);
nor U40269 (N_40269,N_38709,N_39616);
nand U40270 (N_40270,N_38843,N_39564);
and U40271 (N_40271,N_39165,N_38281);
nand U40272 (N_40272,N_39991,N_39885);
or U40273 (N_40273,N_39824,N_37892);
xor U40274 (N_40274,N_37617,N_39973);
and U40275 (N_40275,N_39263,N_37610);
or U40276 (N_40276,N_37805,N_39448);
nand U40277 (N_40277,N_37600,N_39867);
and U40278 (N_40278,N_39021,N_38969);
nand U40279 (N_40279,N_39468,N_39718);
nand U40280 (N_40280,N_38506,N_39185);
nor U40281 (N_40281,N_39339,N_37521);
nand U40282 (N_40282,N_39039,N_37833);
or U40283 (N_40283,N_39682,N_39290);
nand U40284 (N_40284,N_39635,N_39099);
and U40285 (N_40285,N_38276,N_38180);
nand U40286 (N_40286,N_39619,N_39200);
nand U40287 (N_40287,N_38114,N_38504);
or U40288 (N_40288,N_38007,N_39447);
and U40289 (N_40289,N_39354,N_37627);
xnor U40290 (N_40290,N_38181,N_39283);
nand U40291 (N_40291,N_39536,N_37894);
or U40292 (N_40292,N_39804,N_38872);
nor U40293 (N_40293,N_39514,N_39298);
nor U40294 (N_40294,N_39972,N_39035);
nor U40295 (N_40295,N_38044,N_39749);
nand U40296 (N_40296,N_39842,N_39388);
and U40297 (N_40297,N_39827,N_38745);
or U40298 (N_40298,N_37775,N_39856);
and U40299 (N_40299,N_38821,N_38261);
nor U40300 (N_40300,N_39456,N_38923);
nand U40301 (N_40301,N_37738,N_37699);
or U40302 (N_40302,N_39013,N_37726);
and U40303 (N_40303,N_38466,N_37569);
nor U40304 (N_40304,N_39002,N_37591);
or U40305 (N_40305,N_38455,N_38940);
nand U40306 (N_40306,N_39484,N_38828);
xnor U40307 (N_40307,N_38264,N_37684);
and U40308 (N_40308,N_38917,N_39517);
and U40309 (N_40309,N_39927,N_38971);
or U40310 (N_40310,N_38621,N_38384);
xor U40311 (N_40311,N_38397,N_39543);
nor U40312 (N_40312,N_37721,N_37717);
xor U40313 (N_40313,N_37992,N_39413);
xnor U40314 (N_40314,N_39810,N_39757);
nor U40315 (N_40315,N_37533,N_38499);
nand U40316 (N_40316,N_37785,N_38017);
and U40317 (N_40317,N_38560,N_38204);
or U40318 (N_40318,N_37729,N_39605);
or U40319 (N_40319,N_37741,N_39625);
nand U40320 (N_40320,N_38757,N_37663);
xnor U40321 (N_40321,N_39670,N_39844);
nor U40322 (N_40322,N_39113,N_38262);
or U40323 (N_40323,N_38222,N_37968);
nor U40324 (N_40324,N_38727,N_38527);
and U40325 (N_40325,N_37650,N_38119);
and U40326 (N_40326,N_39197,N_37554);
xnor U40327 (N_40327,N_39572,N_38168);
or U40328 (N_40328,N_39004,N_38436);
xnor U40329 (N_40329,N_38174,N_39904);
nand U40330 (N_40330,N_39271,N_39790);
xnor U40331 (N_40331,N_38659,N_38324);
or U40332 (N_40332,N_39016,N_38879);
xnor U40333 (N_40333,N_39034,N_39406);
nand U40334 (N_40334,N_39905,N_39325);
xor U40335 (N_40335,N_39812,N_39037);
or U40336 (N_40336,N_37900,N_39728);
nor U40337 (N_40337,N_39799,N_38322);
nor U40338 (N_40338,N_39296,N_39578);
nor U40339 (N_40339,N_39030,N_37863);
or U40340 (N_40340,N_38022,N_39279);
or U40341 (N_40341,N_38495,N_38690);
or U40342 (N_40342,N_39943,N_39207);
or U40343 (N_40343,N_39845,N_37858);
nand U40344 (N_40344,N_39879,N_39784);
nor U40345 (N_40345,N_39242,N_39322);
nand U40346 (N_40346,N_37631,N_38914);
and U40347 (N_40347,N_38474,N_38140);
and U40348 (N_40348,N_39696,N_38780);
nand U40349 (N_40349,N_38154,N_38983);
nand U40350 (N_40350,N_38894,N_38199);
xnor U40351 (N_40351,N_38967,N_39744);
and U40352 (N_40352,N_39297,N_39986);
or U40353 (N_40353,N_39464,N_38947);
or U40354 (N_40354,N_39571,N_37672);
nor U40355 (N_40355,N_37575,N_37511);
xnor U40356 (N_40356,N_38788,N_39699);
nand U40357 (N_40357,N_39958,N_39055);
nand U40358 (N_40358,N_38539,N_38869);
nand U40359 (N_40359,N_37739,N_38805);
and U40360 (N_40360,N_37922,N_37715);
xnor U40361 (N_40361,N_38175,N_38360);
or U40362 (N_40362,N_38697,N_39208);
xor U40363 (N_40363,N_37566,N_38596);
or U40364 (N_40364,N_38729,N_39114);
nor U40365 (N_40365,N_38837,N_39691);
nor U40366 (N_40366,N_39678,N_38274);
or U40367 (N_40367,N_38406,N_38555);
or U40368 (N_40368,N_37811,N_39982);
nor U40369 (N_40369,N_39333,N_37932);
xor U40370 (N_40370,N_39173,N_37939);
nor U40371 (N_40371,N_37997,N_39712);
xor U40372 (N_40372,N_38832,N_38429);
xnor U40373 (N_40373,N_38041,N_38108);
xor U40374 (N_40374,N_38318,N_37669);
xor U40375 (N_40375,N_38439,N_37506);
or U40376 (N_40376,N_39874,N_39494);
and U40377 (N_40377,N_38992,N_38660);
xor U40378 (N_40378,N_37861,N_39541);
nand U40379 (N_40379,N_39282,N_39159);
or U40380 (N_40380,N_39142,N_38333);
nand U40381 (N_40381,N_38442,N_39683);
nand U40382 (N_40382,N_37559,N_39555);
nand U40383 (N_40383,N_38850,N_38946);
nand U40384 (N_40384,N_38160,N_38185);
and U40385 (N_40385,N_37551,N_39311);
or U40386 (N_40386,N_37963,N_39773);
or U40387 (N_40387,N_39259,N_39818);
and U40388 (N_40388,N_37821,N_38388);
nand U40389 (N_40389,N_39556,N_37572);
nor U40390 (N_40390,N_37960,N_39685);
xor U40391 (N_40391,N_37840,N_39426);
nor U40392 (N_40392,N_37707,N_38123);
nor U40393 (N_40393,N_38155,N_38738);
xor U40394 (N_40394,N_38862,N_38634);
nand U40395 (N_40395,N_38317,N_37834);
or U40396 (N_40396,N_38004,N_38509);
or U40397 (N_40397,N_39975,N_39067);
nand U40398 (N_40398,N_39167,N_39291);
nor U40399 (N_40399,N_38589,N_39396);
and U40400 (N_40400,N_38938,N_39774);
nand U40401 (N_40401,N_37998,N_39892);
xor U40402 (N_40402,N_39626,N_39407);
and U40403 (N_40403,N_38929,N_38827);
xor U40404 (N_40404,N_38065,N_37570);
nor U40405 (N_40405,N_39653,N_39908);
xor U40406 (N_40406,N_38347,N_38959);
nor U40407 (N_40407,N_37984,N_37562);
or U40408 (N_40408,N_37792,N_39671);
xor U40409 (N_40409,N_39843,N_38416);
xor U40410 (N_40410,N_39580,N_39126);
nor U40411 (N_40411,N_39779,N_38023);
or U40412 (N_40412,N_37686,N_39591);
nand U40413 (N_40413,N_39545,N_39680);
nand U40414 (N_40414,N_38620,N_39431);
nor U40415 (N_40415,N_39511,N_39168);
xnor U40416 (N_40416,N_38521,N_37585);
xnor U40417 (N_40417,N_37577,N_39655);
nor U40418 (N_40418,N_37803,N_38547);
or U40419 (N_40419,N_39980,N_39568);
or U40420 (N_40420,N_38075,N_38450);
or U40421 (N_40421,N_39480,N_39969);
nand U40422 (N_40422,N_39976,N_37885);
nor U40423 (N_40423,N_38678,N_38348);
nor U40424 (N_40424,N_39601,N_38195);
nand U40425 (N_40425,N_37593,N_37822);
nor U40426 (N_40426,N_39375,N_39257);
xnor U40427 (N_40427,N_39412,N_38996);
and U40428 (N_40428,N_39492,N_37778);
and U40429 (N_40429,N_38842,N_39024);
xnor U40430 (N_40430,N_37901,N_38926);
xor U40431 (N_40431,N_39537,N_39630);
and U40432 (N_40432,N_38873,N_38941);
and U40433 (N_40433,N_39515,N_38792);
and U40434 (N_40434,N_39393,N_38565);
or U40435 (N_40435,N_39692,N_38006);
nor U40436 (N_40436,N_38537,N_39830);
nand U40437 (N_40437,N_38097,N_39293);
or U40438 (N_40438,N_39459,N_39542);
nor U40439 (N_40439,N_39726,N_39891);
and U40440 (N_40440,N_38591,N_39472);
nand U40441 (N_40441,N_39977,N_38071);
xor U40442 (N_40442,N_37766,N_37671);
and U40443 (N_40443,N_39368,N_38273);
or U40444 (N_40444,N_38482,N_38722);
and U40445 (N_40445,N_39328,N_38890);
or U40446 (N_40446,N_39237,N_38488);
nor U40447 (N_40447,N_39847,N_38799);
xnor U40448 (N_40448,N_38682,N_38036);
nor U40449 (N_40449,N_37973,N_39346);
nor U40450 (N_40450,N_39877,N_38148);
or U40451 (N_40451,N_38149,N_37854);
or U40452 (N_40452,N_38272,N_38355);
or U40453 (N_40453,N_39808,N_38650);
or U40454 (N_40454,N_38478,N_39437);
or U40455 (N_40455,N_39360,N_39404);
nand U40456 (N_40456,N_39736,N_39086);
nand U40457 (N_40457,N_37829,N_38876);
and U40458 (N_40458,N_38896,N_39990);
or U40459 (N_40459,N_39687,N_38315);
nand U40460 (N_40460,N_39315,N_39401);
or U40461 (N_40461,N_37825,N_39451);
xor U40462 (N_40462,N_38207,N_38514);
or U40463 (N_40463,N_38616,N_39706);
and U40464 (N_40464,N_38242,N_39182);
or U40465 (N_40465,N_37820,N_37500);
xor U40466 (N_40466,N_38040,N_38921);
or U40467 (N_40467,N_37666,N_39836);
nand U40468 (N_40468,N_38100,N_39355);
or U40469 (N_40469,N_38422,N_39651);
or U40470 (N_40470,N_38301,N_39917);
xnor U40471 (N_40471,N_39731,N_39902);
or U40472 (N_40472,N_39603,N_37730);
or U40473 (N_40473,N_39092,N_37579);
or U40474 (N_40474,N_38231,N_38213);
or U40475 (N_40475,N_38418,N_39018);
or U40476 (N_40476,N_38479,N_37962);
nand U40477 (N_40477,N_39000,N_38993);
nor U40478 (N_40478,N_38192,N_37765);
nand U40479 (N_40479,N_38076,N_38666);
nand U40480 (N_40480,N_38963,N_39131);
nor U40481 (N_40481,N_39432,N_38358);
and U40482 (N_40482,N_38445,N_37544);
and U40483 (N_40483,N_38948,N_39045);
and U40484 (N_40484,N_39265,N_37946);
nor U40485 (N_40485,N_37887,N_38244);
or U40486 (N_40486,N_39648,N_38054);
nor U40487 (N_40487,N_38985,N_38477);
xor U40488 (N_40488,N_38332,N_39356);
or U40489 (N_40489,N_38999,N_38844);
nor U40490 (N_40490,N_39935,N_39495);
nand U40491 (N_40491,N_39781,N_37644);
xor U40492 (N_40492,N_39970,N_37988);
xor U40493 (N_40493,N_38210,N_39912);
nand U40494 (N_40494,N_38942,N_38913);
and U40495 (N_40495,N_39796,N_38003);
xor U40496 (N_40496,N_37870,N_38846);
and U40497 (N_40497,N_38602,N_38888);
or U40498 (N_40498,N_38390,N_38249);
xor U40499 (N_40499,N_38364,N_37704);
nor U40500 (N_40500,N_39240,N_39175);
nand U40501 (N_40501,N_38642,N_38716);
nand U40502 (N_40502,N_39965,N_37687);
or U40503 (N_40503,N_38126,N_37505);
or U40504 (N_40504,N_37760,N_39888);
nand U40505 (N_40505,N_39933,N_37649);
nand U40506 (N_40506,N_38545,N_37929);
nor U40507 (N_40507,N_39149,N_38919);
nand U40508 (N_40508,N_38124,N_37640);
nor U40509 (N_40509,N_37745,N_39598);
nand U40510 (N_40510,N_38183,N_38807);
nand U40511 (N_40511,N_39612,N_38412);
and U40512 (N_40512,N_37527,N_39665);
and U40513 (N_40513,N_39664,N_38970);
nor U40514 (N_40514,N_39469,N_38391);
or U40515 (N_40515,N_38604,N_38652);
and U40516 (N_40516,N_37690,N_37794);
and U40517 (N_40517,N_39535,N_38704);
xor U40518 (N_40518,N_39466,N_38579);
or U40519 (N_40519,N_38483,N_39195);
and U40520 (N_40520,N_38370,N_39415);
xor U40521 (N_40521,N_39052,N_39579);
or U40522 (N_40522,N_39887,N_39157);
nor U40523 (N_40523,N_39906,N_38597);
nand U40524 (N_40524,N_37891,N_39666);
nor U40525 (N_40525,N_39130,N_39033);
nand U40526 (N_40526,N_37808,N_37513);
xnor U40527 (N_40527,N_37604,N_37667);
nand U40528 (N_40528,N_37656,N_38772);
nor U40529 (N_40529,N_37876,N_38496);
or U40530 (N_40530,N_38354,N_39787);
and U40531 (N_40531,N_39688,N_38671);
nor U40532 (N_40532,N_39499,N_39896);
and U40533 (N_40533,N_38974,N_38668);
and U40534 (N_40534,N_37737,N_39442);
xnor U40535 (N_40535,N_37804,N_38791);
xnor U40536 (N_40536,N_38689,N_39721);
nor U40537 (N_40537,N_38260,N_38367);
nand U40538 (N_40538,N_39324,N_37586);
xor U40539 (N_40539,N_37727,N_38498);
and U40540 (N_40540,N_38637,N_37675);
nand U40541 (N_40541,N_37629,N_37835);
nor U40542 (N_40542,N_37525,N_39516);
nor U40543 (N_40543,N_38608,N_38601);
xor U40544 (N_40544,N_37653,N_38595);
or U40545 (N_40545,N_39614,N_38157);
nor U40546 (N_40546,N_39631,N_39627);
nor U40547 (N_40547,N_37563,N_37916);
xnor U40548 (N_40548,N_38172,N_37618);
nand U40549 (N_40549,N_39090,N_38889);
and U40550 (N_40550,N_38973,N_38139);
nand U40551 (N_40551,N_37581,N_39539);
xnor U40552 (N_40552,N_38756,N_37934);
nor U40553 (N_40553,N_38950,N_39502);
or U40554 (N_40554,N_37628,N_39956);
nand U40555 (N_40555,N_38164,N_38566);
and U40556 (N_40556,N_39329,N_38203);
nor U40557 (N_40557,N_38133,N_38624);
and U40558 (N_40558,N_39221,N_39082);
xnor U40559 (N_40559,N_39161,N_38951);
and U40560 (N_40560,N_38059,N_38377);
nor U40561 (N_40561,N_39403,N_39457);
or U40562 (N_40562,N_38693,N_39049);
nand U40563 (N_40563,N_39006,N_39771);
or U40564 (N_40564,N_38893,N_38885);
nand U40565 (N_40565,N_39075,N_38978);
nand U40566 (N_40566,N_39621,N_38575);
and U40567 (N_40567,N_37702,N_38117);
xnor U40568 (N_40568,N_39487,N_38865);
or U40569 (N_40569,N_38206,N_38866);
nor U40570 (N_40570,N_37990,N_39848);
nand U40571 (N_40571,N_39788,N_38531);
and U40572 (N_40572,N_38875,N_37925);
nand U40573 (N_40573,N_39681,N_37661);
nor U40574 (N_40574,N_39646,N_38423);
and U40575 (N_40575,N_37524,N_39597);
or U40576 (N_40576,N_39124,N_39761);
or U40577 (N_40577,N_38935,N_38008);
nor U40578 (N_40578,N_38784,N_37734);
nor U40579 (N_40579,N_38177,N_39352);
xor U40580 (N_40580,N_37510,N_38630);
nor U40581 (N_40581,N_38018,N_38299);
nor U40582 (N_40582,N_38662,N_38501);
xnor U40583 (N_40583,N_39639,N_39669);
nand U40584 (N_40584,N_39235,N_39613);
xnor U40585 (N_40585,N_39709,N_38257);
and U40586 (N_40586,N_38787,N_39316);
nor U40587 (N_40587,N_39838,N_37802);
nand U40588 (N_40588,N_39698,N_38909);
nor U40589 (N_40589,N_38976,N_39141);
or U40590 (N_40590,N_38001,N_37567);
xnor U40591 (N_40591,N_39107,N_38473);
xnor U40592 (N_40592,N_39273,N_37693);
or U40593 (N_40593,N_39674,N_38465);
nand U40594 (N_40594,N_39476,N_38763);
and U40595 (N_40595,N_39009,N_37800);
xor U40596 (N_40596,N_39828,N_39225);
xnor U40597 (N_40597,N_39554,N_39899);
nor U40598 (N_40598,N_38793,N_39586);
or U40599 (N_40599,N_38623,N_38962);
nor U40600 (N_40600,N_37582,N_38307);
nor U40601 (N_40601,N_39012,N_39756);
nor U40602 (N_40602,N_38874,N_37540);
nor U40603 (N_40603,N_39144,N_38268);
xnor U40604 (N_40604,N_37888,N_39490);
nand U40605 (N_40605,N_38752,N_37561);
nor U40606 (N_40606,N_39743,N_39077);
nand U40607 (N_40607,N_39604,N_38344);
xnor U40608 (N_40608,N_39768,N_39941);
xnor U40609 (N_40609,N_39102,N_38901);
nor U40610 (N_40610,N_38338,N_39351);
nand U40611 (N_40611,N_39694,N_38674);
nor U40612 (N_40612,N_39615,N_37837);
xnor U40613 (N_40613,N_38852,N_38241);
nor U40614 (N_40614,N_37665,N_39629);
nor U40615 (N_40615,N_37847,N_38366);
nand U40616 (N_40616,N_38103,N_39101);
and U40617 (N_40617,N_39230,N_39684);
nand U40618 (N_40618,N_39548,N_38083);
and U40619 (N_40619,N_38425,N_39512);
and U40620 (N_40620,N_39703,N_39538);
nand U40621 (N_40621,N_38087,N_39080);
xnor U40622 (N_40622,N_39984,N_37823);
or U40623 (N_40623,N_38585,N_39850);
nor U40624 (N_40624,N_38806,N_39286);
nand U40625 (N_40625,N_38239,N_39567);
and U40626 (N_40626,N_38771,N_37780);
and U40627 (N_40627,N_37556,N_39483);
or U40628 (N_40628,N_39576,N_39570);
xnor U40629 (N_40629,N_37873,N_38170);
xnor U40630 (N_40630,N_37662,N_39384);
nand U40631 (N_40631,N_37869,N_38556);
and U40632 (N_40632,N_37905,N_38109);
xor U40633 (N_40633,N_38066,N_37592);
nand U40634 (N_40634,N_37750,N_38853);
and U40635 (N_40635,N_39921,N_39503);
and U40636 (N_40636,N_37816,N_37602);
xor U40637 (N_40637,N_38052,N_39177);
or U40638 (N_40638,N_38024,N_39767);
xnor U40639 (N_40639,N_39777,N_39819);
xnor U40640 (N_40640,N_38201,N_38861);
xor U40641 (N_40641,N_39909,N_38676);
nand U40642 (N_40642,N_38858,N_37798);
and U40643 (N_40643,N_38340,N_37852);
or U40644 (N_40644,N_39782,N_38653);
xor U40645 (N_40645,N_39261,N_38188);
and U40646 (N_40646,N_39600,N_37924);
nor U40647 (N_40647,N_39934,N_39826);
or U40648 (N_40648,N_38728,N_38774);
or U40649 (N_40649,N_39898,N_38411);
nand U40650 (N_40650,N_39196,N_38800);
xnor U40651 (N_40651,N_37949,N_38902);
nand U40652 (N_40652,N_37657,N_38233);
or U40653 (N_40653,N_37877,N_38153);
and U40654 (N_40654,N_39620,N_38831);
or U40655 (N_40655,N_37917,N_39441);
and U40656 (N_40656,N_38764,N_39191);
nor U40657 (N_40657,N_37691,N_38708);
and U40658 (N_40658,N_39379,N_38053);
and U40659 (N_40659,N_39791,N_37814);
or U40660 (N_40660,N_37991,N_38060);
nand U40661 (N_40661,N_39121,N_38673);
nor U40662 (N_40662,N_39183,N_39314);
or U40663 (N_40663,N_39319,N_37926);
xor U40664 (N_40664,N_39966,N_37849);
or U40665 (N_40665,N_39359,N_38968);
xnor U40666 (N_40666,N_39835,N_39001);
and U40667 (N_40667,N_38171,N_38389);
or U40668 (N_40668,N_37860,N_39374);
or U40669 (N_40669,N_38420,N_39947);
and U40670 (N_40670,N_38468,N_39852);
and U40671 (N_40671,N_37862,N_38452);
xor U40672 (N_40672,N_38494,N_38972);
or U40673 (N_40673,N_37830,N_39211);
or U40674 (N_40674,N_39186,N_38373);
and U40675 (N_40675,N_39061,N_38070);
or U40676 (N_40676,N_38851,N_39139);
nand U40677 (N_40677,N_37550,N_37711);
and U40678 (N_40678,N_38649,N_38838);
nand U40679 (N_40679,N_39239,N_39122);
nor U40680 (N_40680,N_39097,N_38021);
and U40681 (N_40681,N_39890,N_38002);
or U40682 (N_40682,N_38263,N_38685);
or U40683 (N_40683,N_38321,N_39550);
and U40684 (N_40684,N_37740,N_38641);
or U40685 (N_40685,N_39128,N_37999);
or U40686 (N_40686,N_39785,N_39341);
xnor U40687 (N_40687,N_38737,N_38491);
and U40688 (N_40688,N_39944,N_39929);
or U40689 (N_40689,N_39676,N_39170);
xor U40690 (N_40690,N_38686,N_38104);
xnor U40691 (N_40691,N_39675,N_38916);
nand U40692 (N_40692,N_37810,N_38167);
nand U40693 (N_40693,N_38997,N_38292);
nand U40694 (N_40694,N_39458,N_38015);
or U40695 (N_40695,N_38019,N_39533);
nor U40696 (N_40696,N_37777,N_38904);
nand U40697 (N_40697,N_38618,N_37643);
or U40698 (N_40698,N_39343,N_38920);
or U40699 (N_40699,N_37982,N_37531);
or U40700 (N_40700,N_39253,N_37758);
nand U40701 (N_40701,N_39753,N_38814);
xor U40702 (N_40702,N_38029,N_39507);
and U40703 (N_40703,N_39951,N_38069);
nand U40704 (N_40704,N_38747,N_37539);
xor U40705 (N_40705,N_39702,N_38072);
nand U40706 (N_40706,N_39926,N_39245);
nor U40707 (N_40707,N_37733,N_39020);
and U40708 (N_40708,N_38580,N_37553);
xor U40709 (N_40709,N_38232,N_37526);
and U40710 (N_40710,N_39320,N_39125);
nand U40711 (N_40711,N_38955,N_37692);
and U40712 (N_40712,N_38325,N_38363);
nand U40713 (N_40713,N_38731,N_37971);
xnor U40714 (N_40714,N_37616,N_39732);
or U40715 (N_40715,N_39792,N_39050);
or U40716 (N_40716,N_38467,N_38696);
nand U40717 (N_40717,N_39634,N_37546);
xnor U40718 (N_40718,N_37920,N_39040);
and U40719 (N_40719,N_38856,N_38860);
or U40720 (N_40720,N_38907,N_38311);
or U40721 (N_40721,N_37728,N_39544);
nand U40722 (N_40722,N_39461,N_39247);
and U40723 (N_40723,N_39334,N_37674);
or U40724 (N_40724,N_39750,N_39344);
xnor U40725 (N_40725,N_39558,N_39193);
and U40726 (N_40726,N_39327,N_38960);
or U40727 (N_40727,N_39189,N_38306);
and U40728 (N_40728,N_38457,N_38573);
and U40729 (N_40729,N_37824,N_39417);
nand U40730 (N_40730,N_39058,N_38459);
xnor U40731 (N_40731,N_39747,N_38484);
xor U40732 (N_40732,N_38648,N_37545);
nand U40733 (N_40733,N_38234,N_39971);
xor U40734 (N_40734,N_38925,N_39234);
and U40735 (N_40735,N_37857,N_37819);
or U40736 (N_40736,N_39089,N_37609);
and U40737 (N_40737,N_39336,N_38769);
nor U40738 (N_40738,N_37807,N_38110);
xor U40739 (N_40739,N_39105,N_38287);
xnor U40740 (N_40740,N_38818,N_38470);
xor U40741 (N_40741,N_37923,N_38735);
and U40742 (N_40742,N_39562,N_38461);
nand U40743 (N_40743,N_38392,N_37517);
and U40744 (N_40744,N_38033,N_39897);
xor U40745 (N_40745,N_37658,N_38561);
or U40746 (N_40746,N_37573,N_39611);
or U40747 (N_40747,N_38162,N_39738);
nor U40748 (N_40748,N_38801,N_38371);
or U40749 (N_40749,N_37952,N_39595);
and U40750 (N_40750,N_39701,N_39807);
or U40751 (N_40751,N_38891,N_38039);
xnor U40752 (N_40752,N_38254,N_37709);
or U40753 (N_40753,N_39531,N_38609);
and U40754 (N_40754,N_39120,N_38614);
nor U40755 (N_40755,N_37838,N_38235);
and U40756 (N_40756,N_38221,N_39188);
xor U40757 (N_40757,N_39059,N_38267);
nand U40758 (N_40758,N_38867,N_39056);
nor U40759 (N_40759,N_38279,N_38980);
or U40760 (N_40760,N_39802,N_39252);
or U40761 (N_40761,N_38523,N_39742);
xor U40762 (N_40762,N_39552,N_39623);
xor U40763 (N_40763,N_38352,N_39633);
or U40764 (N_40764,N_39673,N_39957);
nor U40765 (N_40765,N_39805,N_37621);
nor U40766 (N_40766,N_39711,N_37626);
xnor U40767 (N_40767,N_37941,N_37537);
nor U40768 (N_40768,N_37676,N_39038);
xor U40769 (N_40769,N_37630,N_37996);
and U40770 (N_40770,N_39776,N_38253);
nor U40771 (N_40771,N_38237,N_39679);
xnor U40772 (N_40772,N_38823,N_39243);
or U40773 (N_40773,N_38045,N_38503);
nor U40774 (N_40774,N_38421,N_39860);
nand U40775 (N_40775,N_39660,N_39717);
xor U40776 (N_40776,N_37742,N_37522);
or U40777 (N_40777,N_38309,N_39072);
xor U40778 (N_40778,N_37866,N_39402);
nor U40779 (N_40779,N_39959,N_37588);
or U40780 (N_40780,N_38781,N_39088);
and U40781 (N_40781,N_38625,N_39119);
xor U40782 (N_40782,N_38939,N_39524);
xnor U40783 (N_40783,N_38834,N_38471);
nand U40784 (N_40784,N_38505,N_37789);
nor U40785 (N_40785,N_39795,N_38385);
nand U40786 (N_40786,N_38912,N_37599);
or U40787 (N_40787,N_39607,N_38169);
or U40788 (N_40788,N_39924,N_38987);
xor U40789 (N_40789,N_38176,N_39884);
nor U40790 (N_40790,N_38656,N_39725);
nor U40791 (N_40791,N_38758,N_37703);
and U40792 (N_40792,N_38817,N_38786);
and U40793 (N_40793,N_39916,N_37907);
nand U40794 (N_40794,N_37764,N_37753);
and U40795 (N_40795,N_39409,N_39960);
and U40796 (N_40796,N_39385,N_37624);
nand U40797 (N_40797,N_38713,N_39923);
or U40798 (N_40798,N_39723,N_39383);
nor U40799 (N_40799,N_37817,N_39135);
nor U40800 (N_40800,N_39523,N_39386);
and U40801 (N_40801,N_38863,N_39816);
nor U40802 (N_40802,N_39063,N_37937);
or U40803 (N_40803,N_38719,N_39287);
nor U40804 (N_40804,N_38089,N_38378);
nand U40805 (N_40805,N_38228,N_37921);
and U40806 (N_40806,N_39637,N_39233);
nand U40807 (N_40807,N_39109,N_38753);
or U40808 (N_40808,N_38000,N_39759);
nand U40809 (N_40809,N_39215,N_39236);
xor U40810 (N_40810,N_39203,N_39928);
nor U40811 (N_40811,N_39348,N_38508);
and U40812 (N_40812,N_38661,N_38129);
nor U40813 (N_40813,N_37879,N_37754);
nand U40814 (N_40814,N_38881,N_37689);
xnor U40815 (N_40815,N_39868,N_38336);
nor U40816 (N_40816,N_39103,N_39312);
nor U40817 (N_40817,N_39740,N_38581);
and U40818 (N_40818,N_37787,N_38855);
nand U40819 (N_40819,N_38394,N_38622);
nand U40820 (N_40820,N_37659,N_39187);
nand U40821 (N_40821,N_39347,N_39123);
nand U40822 (N_40822,N_38783,N_38739);
nand U40823 (N_40823,N_37771,N_38892);
xnor U40824 (N_40824,N_38401,N_39436);
xor U40825 (N_40825,N_39152,N_38298);
and U40826 (N_40826,N_39326,N_38432);
nor U40827 (N_40827,N_38762,N_39053);
nand U40828 (N_40828,N_39475,N_37637);
or U40829 (N_40829,N_39137,N_39274);
nand U40830 (N_40830,N_38365,N_39411);
or U40831 (N_40831,N_39996,N_38294);
or U40832 (N_40832,N_37945,N_37772);
xnor U40833 (N_40833,N_38826,N_38462);
nand U40834 (N_40834,N_37853,N_38532);
nor U40835 (N_40835,N_39434,N_39946);
and U40836 (N_40836,N_38605,N_39047);
nor U40837 (N_40837,N_37529,N_39663);
and U40838 (N_40838,N_39060,N_39395);
nor U40839 (N_40839,N_39249,N_39840);
nor U40840 (N_40840,N_38048,N_38480);
and U40841 (N_40841,N_39863,N_37683);
xnor U40842 (N_40842,N_39285,N_39460);
nand U40843 (N_40843,N_39968,N_38493);
xor U40844 (N_40844,N_37913,N_39222);
xnor U40845 (N_40845,N_37976,N_39932);
and U40846 (N_40846,N_38607,N_39127);
or U40847 (N_40847,N_38278,N_39267);
nor U40848 (N_40848,N_39398,N_38271);
nand U40849 (N_40849,N_38460,N_38165);
nor U40850 (N_40850,N_38518,N_38928);
nor U40851 (N_40851,N_37928,N_38356);
nor U40852 (N_40852,N_38275,N_37636);
and U40853 (N_40853,N_39134,N_39861);
xor U40854 (N_40854,N_39727,N_37906);
nor U40855 (N_40855,N_38105,N_39248);
or U40856 (N_40856,N_37598,N_37881);
nor U40857 (N_40857,N_38409,N_39376);
and U40858 (N_40858,N_39066,N_39751);
xor U40859 (N_40859,N_39871,N_38900);
nand U40860 (N_40860,N_37614,N_39820);
nand U40861 (N_40861,N_39232,N_38871);
and U40862 (N_40862,N_38326,N_38353);
nand U40863 (N_40863,N_38132,N_39380);
nand U40864 (N_40864,N_39151,N_37955);
or U40865 (N_40865,N_38524,N_39705);
or U40866 (N_40866,N_39895,N_39266);
or U40867 (N_40867,N_38628,N_38937);
and U40868 (N_40868,N_37694,N_38464);
and U40869 (N_40869,N_37520,N_39695);
and U40870 (N_40870,N_37713,N_39662);
xnor U40871 (N_40871,N_38447,N_38824);
xor U40872 (N_40872,N_38035,N_37868);
and U40873 (N_40873,N_38010,N_39504);
and U40874 (N_40874,N_39783,N_39229);
or U40875 (N_40875,N_37809,N_39023);
or U40876 (N_40876,N_39697,N_38043);
and U40877 (N_40877,N_38530,N_38720);
or U40878 (N_40878,N_39463,N_37596);
nand U40879 (N_40879,N_37987,N_38700);
xnor U40880 (N_40880,N_38918,N_38507);
xnor U40881 (N_40881,N_38705,N_37535);
nand U40882 (N_40882,N_38142,N_37503);
and U40883 (N_40883,N_39823,N_37914);
or U40884 (N_40884,N_39735,N_38924);
or U40885 (N_40885,N_38382,N_39522);
nand U40886 (N_40886,N_37565,N_39907);
and U40887 (N_40887,N_38712,N_38094);
nor U40888 (N_40888,N_38711,N_39154);
nand U40889 (N_40889,N_39238,N_38578);
nand U40890 (N_40890,N_37757,N_39998);
nand U40891 (N_40891,N_39618,N_39693);
nor U40892 (N_40892,N_38574,N_39465);
nand U40893 (N_40893,N_39700,N_38643);
nor U40894 (N_40894,N_39569,N_37832);
and U40895 (N_40895,N_39745,N_39019);
or U40896 (N_40896,N_38911,N_38776);
or U40897 (N_40897,N_38265,N_38403);
nor U40898 (N_40898,N_38586,N_39335);
and U40899 (N_40899,N_38329,N_38615);
nand U40900 (N_40900,N_39638,N_39198);
nor U40901 (N_40901,N_37601,N_38147);
nand U40902 (N_40902,N_37972,N_39219);
nor U40903 (N_40903,N_39228,N_37878);
or U40904 (N_40904,N_37989,N_39162);
xor U40905 (N_40905,N_38553,N_38945);
nand U40906 (N_40906,N_39081,N_37897);
nand U40907 (N_40907,N_39479,N_39881);
nor U40908 (N_40908,N_38112,N_39833);
nor U40909 (N_40909,N_39622,N_39624);
nor U40910 (N_40910,N_38443,N_38811);
or U40911 (N_40911,N_39416,N_38182);
nor U40912 (N_40912,N_39983,N_39936);
and U40913 (N_40913,N_38399,N_37983);
or U40914 (N_40914,N_38677,N_39563);
nor U40915 (N_40915,N_39883,N_38886);
and U40916 (N_40916,N_39305,N_38225);
xnor U40917 (N_40917,N_37568,N_39746);
nand U40918 (N_40918,N_39733,N_37597);
nor U40919 (N_40919,N_39027,N_37813);
or U40920 (N_40920,N_38050,N_39801);
and U40921 (N_40921,N_38808,N_37936);
xor U40922 (N_40922,N_39961,N_39497);
nor U40923 (N_40923,N_39889,N_39184);
and U40924 (N_40924,N_39764,N_37790);
nand U40925 (N_40925,N_39995,N_37801);
or U40926 (N_40926,N_39962,N_37642);
nand U40927 (N_40927,N_37978,N_38107);
or U40928 (N_40928,N_39350,N_38593);
or U40929 (N_40929,N_38687,N_39754);
or U40930 (N_40930,N_37523,N_37543);
and U40931 (N_40931,N_39584,N_39277);
or U40932 (N_40932,N_39748,N_39708);
xnor U40933 (N_40933,N_38651,N_38825);
nand U40934 (N_40934,N_37836,N_37818);
nand U40935 (N_40935,N_39602,N_38598);
and U40936 (N_40936,N_39438,N_38088);
or U40937 (N_40937,N_39498,N_39886);
or U40938 (N_40938,N_39643,N_38584);
or U40939 (N_40939,N_39493,N_39421);
nand U40940 (N_40940,N_38952,N_38770);
nand U40941 (N_40941,N_39424,N_39364);
or U40942 (N_40942,N_39158,N_39491);
or U40943 (N_40943,N_38698,N_39734);
nor U40944 (N_40944,N_37695,N_38102);
and U40945 (N_40945,N_39870,N_38979);
xnor U40946 (N_40946,N_38989,N_38313);
nor U40947 (N_40947,N_38350,N_38529);
and U40948 (N_40948,N_39496,N_38191);
nand U40949 (N_40949,N_38957,N_39878);
or U40950 (N_40950,N_38212,N_38688);
or U40951 (N_40951,N_37883,N_38304);
xnor U40952 (N_40952,N_37769,N_38375);
and U40953 (N_40953,N_37867,N_39209);
nor U40954 (N_40954,N_38707,N_38767);
nor U40955 (N_40955,N_38633,N_38251);
or U40956 (N_40956,N_39419,N_39762);
or U40957 (N_40957,N_39003,N_38617);
or U40958 (N_40958,N_38013,N_38744);
or U40959 (N_40959,N_37841,N_38343);
nand U40960 (N_40960,N_39321,N_38291);
and U40961 (N_40961,N_38544,N_38440);
nand U40962 (N_40962,N_37647,N_39382);
xor U40963 (N_40963,N_38223,N_39367);
or U40964 (N_40964,N_39640,N_39981);
nand U40965 (N_40965,N_39008,N_39474);
xnor U40966 (N_40966,N_39577,N_38302);
or U40967 (N_40967,N_39378,N_38099);
or U40968 (N_40968,N_39444,N_38699);
nor U40969 (N_40969,N_38635,N_38259);
nor U40970 (N_40970,N_38288,N_37933);
or U40971 (N_40971,N_38572,N_38238);
nand U40972 (N_40972,N_39628,N_39204);
and U40973 (N_40973,N_37761,N_39815);
and U40974 (N_40974,N_38736,N_38096);
xor U40975 (N_40975,N_38381,N_39213);
xor U40976 (N_40976,N_37679,N_38138);
nor U40977 (N_40977,N_39145,N_39313);
xnor U40978 (N_40978,N_38857,N_39532);
and U40979 (N_40979,N_39950,N_38230);
nand U40980 (N_40980,N_38383,N_38554);
or U40981 (N_40981,N_38541,N_37896);
nor U40982 (N_40982,N_38453,N_38376);
and U40983 (N_40983,N_38245,N_37654);
nor U40984 (N_40984,N_39227,N_38732);
xor U40985 (N_40985,N_38943,N_39587);
xor U40986 (N_40986,N_38476,N_37723);
or U40987 (N_40987,N_38079,N_38640);
xnor U40988 (N_40988,N_37718,N_39647);
nand U40989 (N_40989,N_37688,N_37514);
nor U40990 (N_40990,N_39318,N_39608);
or U40991 (N_40991,N_38675,N_38681);
xor U40992 (N_40992,N_39254,N_38956);
or U40993 (N_40993,N_39999,N_39500);
nand U40994 (N_40994,N_37724,N_39854);
or U40995 (N_40995,N_37607,N_39903);
xor U40996 (N_40996,N_38915,N_39212);
or U40997 (N_40997,N_37536,N_39713);
nand U40998 (N_40998,N_37747,N_38011);
nor U40999 (N_40999,N_38994,N_37895);
or U41000 (N_41000,N_38433,N_37986);
nand U41001 (N_41001,N_38334,N_37595);
xor U41002 (N_41002,N_38341,N_38849);
xor U41003 (N_41003,N_37762,N_37587);
and U41004 (N_41004,N_38209,N_38305);
or U41005 (N_41005,N_37710,N_39817);
nor U41006 (N_41006,N_39138,N_37756);
and U41007 (N_41007,N_39394,N_37648);
and U41008 (N_41008,N_38644,N_38219);
nor U41009 (N_41009,N_38568,N_38489);
and U41010 (N_41010,N_39370,N_38152);
xnor U41011 (N_41011,N_39661,N_39590);
nor U41012 (N_41012,N_39467,N_39942);
nor U41013 (N_41013,N_38820,N_39914);
nand U41014 (N_41014,N_37884,N_39022);
nor U41015 (N_41015,N_39652,N_38337);
nor U41016 (N_41016,N_39592,N_38448);
nand U41017 (N_41017,N_37890,N_38520);
and U41018 (N_41018,N_39414,N_39435);
nand U41019 (N_41019,N_37979,N_39171);
nand U41020 (N_41020,N_39794,N_38706);
and U41021 (N_41021,N_38481,N_37685);
nand U41022 (N_41022,N_38402,N_38487);
or U41023 (N_41023,N_39657,N_38186);
nand U41024 (N_41024,N_37793,N_38797);
or U41025 (N_41025,N_38408,N_38379);
and U41026 (N_41026,N_37634,N_37779);
nand U41027 (N_41027,N_39156,N_39832);
or U41028 (N_41028,N_39408,N_39278);
or U41029 (N_41029,N_38134,N_37953);
xnor U41030 (N_41030,N_37850,N_39284);
or U41031 (N_41031,N_39251,N_38984);
xnor U41032 (N_41032,N_38761,N_39362);
and U41033 (N_41033,N_39869,N_38679);
xor U41034 (N_41034,N_38569,N_39178);
and U41035 (N_41035,N_37603,N_39967);
nor U41036 (N_41036,N_38515,N_37507);
xor U41037 (N_41037,N_38782,N_38374);
and U41038 (N_41038,N_38092,N_37678);
nor U41039 (N_41039,N_39729,N_38269);
nand U41040 (N_41040,N_38567,N_39920);
nor U41041 (N_41041,N_38270,N_39583);
nand U41042 (N_41042,N_37882,N_39610);
and U41043 (N_41043,N_38995,N_37712);
or U41044 (N_41044,N_39851,N_38135);
xnor U41045 (N_41045,N_39250,N_39104);
nand U41046 (N_41046,N_38646,N_37786);
or U41047 (N_41047,N_38551,N_38130);
xnor U41048 (N_41048,N_39455,N_38431);
xnor U41049 (N_41049,N_38405,N_38658);
nor U41050 (N_41050,N_37856,N_38664);
nor U41051 (N_41051,N_39589,N_37918);
nand U41052 (N_41052,N_38750,N_39862);
xor U41053 (N_41053,N_38246,N_39880);
xor U41054 (N_41054,N_38667,N_37680);
nor U41055 (N_41055,N_39829,N_39218);
nand U41056 (N_41056,N_37622,N_38636);
xor U41057 (N_41057,N_38703,N_38417);
xnor U41058 (N_41058,N_38830,N_37594);
or U41059 (N_41059,N_39508,N_38016);
xnor U41060 (N_41060,N_39477,N_38047);
nand U41061 (N_41061,N_39381,N_39690);
or U41062 (N_41062,N_39260,N_39246);
xnor U41063 (N_41063,N_38380,N_37731);
or U41064 (N_41064,N_38903,N_38144);
and U41065 (N_41065,N_37512,N_37736);
and U41066 (N_41066,N_39358,N_38534);
nand U41067 (N_41067,N_38284,N_38715);
or U41068 (N_41068,N_38314,N_39857);
or U41069 (N_41069,N_38163,N_39488);
or U41070 (N_41070,N_39509,N_37719);
nand U41071 (N_41071,N_38899,N_39798);
nand U41072 (N_41072,N_39901,N_39241);
nand U41073 (N_41073,N_38328,N_38936);
or U41074 (N_41074,N_37943,N_38410);
nor U41075 (N_41075,N_37716,N_39117);
and U41076 (N_41076,N_39724,N_38694);
and U41077 (N_41077,N_38194,N_38081);
or U41078 (N_41078,N_37964,N_38647);
or U41079 (N_41079,N_38025,N_38669);
nand U41080 (N_41080,N_39645,N_37746);
nor U41081 (N_41081,N_39269,N_38166);
nor U41082 (N_41082,N_39136,N_39853);
nor U41083 (N_41083,N_39900,N_39553);
xnor U41084 (N_41084,N_38619,N_37655);
nand U41085 (N_41085,N_39306,N_39992);
or U41086 (N_41086,N_37796,N_37720);
or U41087 (N_41087,N_39025,N_37555);
or U41088 (N_41088,N_37791,N_39095);
xor U41089 (N_41089,N_37519,N_37501);
xor U41090 (N_41090,N_39391,N_37966);
and U41091 (N_41091,N_38815,N_38908);
xor U41092 (N_41092,N_38285,N_39366);
nor U41093 (N_41093,N_39310,N_39546);
and U41094 (N_41094,N_37696,N_38878);
xnor U41095 (N_41095,N_39180,N_39915);
xor U41096 (N_41096,N_39752,N_39989);
xor U41097 (N_41097,N_39153,N_39192);
and U41098 (N_41098,N_39922,N_38143);
and U41099 (N_41099,N_38610,N_39482);
and U41100 (N_41100,N_39510,N_37732);
xor U41101 (N_41101,N_39739,N_39865);
or U41102 (N_41102,N_39581,N_39913);
and U41103 (N_41103,N_39071,N_37908);
and U41104 (N_41104,N_39528,N_38564);
nand U41105 (N_41105,N_38118,N_38582);
and U41106 (N_41106,N_39780,N_39686);
and U41107 (N_41107,N_39994,N_39361);
nor U41108 (N_41108,N_39834,N_39308);
and U41109 (N_41109,N_37590,N_38217);
nor U41110 (N_41110,N_38295,N_39704);
nor U41111 (N_41111,N_38127,N_38513);
nand U41112 (N_41112,N_38812,N_38085);
xnor U41113 (N_41113,N_39079,N_38749);
xor U41114 (N_41114,N_38320,N_39428);
or U41115 (N_41115,N_38220,N_38032);
and U41116 (N_41116,N_39987,N_38599);
xor U41117 (N_41117,N_38528,N_37574);
nor U41118 (N_41118,N_38330,N_39106);
or U41119 (N_41119,N_38372,N_38490);
or U41120 (N_41120,N_39309,N_39654);
and U41121 (N_41121,N_39938,N_38327);
or U41122 (N_41122,N_39534,N_38345);
and U41123 (N_41123,N_38627,N_39719);
or U41124 (N_41124,N_38822,N_38393);
nand U41125 (N_41125,N_37893,N_38723);
nand U41126 (N_41126,N_38510,N_38082);
nor U41127 (N_41127,N_38833,N_39094);
and U41128 (N_41128,N_39940,N_38794);
or U41129 (N_41129,N_37948,N_38778);
and U41130 (N_41130,N_39875,N_38775);
and U41131 (N_41131,N_39073,N_39440);
or U41132 (N_41132,N_39275,N_38603);
or U41133 (N_41133,N_38266,N_39636);
nor U41134 (N_41134,N_38559,N_38655);
and U41135 (N_41135,N_39300,N_39585);
nand U41136 (N_41136,N_39707,N_38296);
and U41137 (N_41137,N_38702,N_38335);
xor U41138 (N_41138,N_38357,N_39304);
nand U41139 (N_41139,N_37859,N_39418);
xnor U41140 (N_41140,N_38247,N_37763);
and U41141 (N_41141,N_38883,N_37504);
xor U41142 (N_41142,N_39181,N_39342);
nor U41143 (N_41143,N_38751,N_38982);
or U41144 (N_41144,N_38456,N_38670);
and U41145 (N_41145,N_37902,N_39955);
xnor U41146 (N_41146,N_37706,N_37755);
xor U41147 (N_41147,N_38546,N_38074);
or U41148 (N_41148,N_38485,N_39070);
nor U41149 (N_41149,N_39763,N_39371);
and U41150 (N_41150,N_39893,N_38905);
nor U41151 (N_41151,N_38519,N_38887);
or U41152 (N_41152,N_39518,N_38413);
nor U41153 (N_41153,N_39289,N_38359);
nand U41154 (N_41154,N_39513,N_38214);
nor U41155 (N_41155,N_39446,N_39169);
nor U41156 (N_41156,N_38975,N_39997);
or U41157 (N_41157,N_37558,N_39566);
nand U41158 (N_41158,N_39029,N_38034);
and U41159 (N_41159,N_38150,N_39244);
nand U41160 (N_41160,N_37875,N_38184);
xor U41161 (N_41161,N_39091,N_37625);
and U41162 (N_41162,N_38958,N_39672);
and U41163 (N_41163,N_38710,N_39963);
nand U41164 (N_41164,N_37641,N_39410);
nand U41165 (N_41165,N_39778,N_39766);
nor U41166 (N_41166,N_38451,N_38492);
nand U41167 (N_41167,N_38773,N_38692);
nand U41168 (N_41168,N_38101,N_38111);
nor U41169 (N_41169,N_38125,N_38988);
or U41170 (N_41170,N_39606,N_38512);
and U41171 (N_41171,N_38122,N_39074);
nor U41172 (N_41172,N_38724,N_37950);
nand U41173 (N_41173,N_37965,N_38836);
or U41174 (N_41174,N_37632,N_38714);
nand U41175 (N_41175,N_39166,N_38224);
nor U41176 (N_41176,N_37749,N_39054);
nor U41177 (N_41177,N_39276,N_38577);
nor U41178 (N_41178,N_39979,N_38098);
xor U41179 (N_41179,N_39557,N_37623);
nor U41180 (N_41180,N_37784,N_39710);
nor U41181 (N_41181,N_38933,N_39307);
xor U41182 (N_41182,N_38611,N_39129);
nor U41183 (N_41183,N_38106,N_38146);
and U41184 (N_41184,N_38657,N_38798);
xnor U41185 (N_41185,N_39140,N_39160);
xnor U41186 (N_41186,N_37931,N_39650);
nand U41187 (N_41187,N_38847,N_38535);
or U41188 (N_41188,N_38802,N_37619);
and U41189 (N_41189,N_37947,N_37534);
nand U41190 (N_41190,N_37899,N_39925);
or U41191 (N_41191,N_37954,N_39083);
nor U41192 (N_41192,N_38049,N_37673);
xnor U41193 (N_41193,N_38740,N_39846);
or U41194 (N_41194,N_37538,N_39280);
nand U41195 (N_41195,N_39032,N_37633);
or U41196 (N_41196,N_38368,N_37842);
or U41197 (N_41197,N_37774,N_38323);
nand U41198 (N_41198,N_37516,N_39096);
nor U41199 (N_41199,N_39108,N_39365);
xor U41200 (N_41200,N_37980,N_38898);
nand U41201 (N_41201,N_37701,N_38964);
xor U41202 (N_41202,N_38734,N_39527);
or U41203 (N_41203,N_38835,N_37848);
and U41204 (N_41204,N_37944,N_38063);
nand U41205 (N_41205,N_38536,N_38121);
or U41206 (N_41206,N_38458,N_39028);
or U41207 (N_41207,N_39439,N_39422);
nand U41208 (N_41208,N_38741,N_39978);
nand U41209 (N_41209,N_39357,N_38606);
xnor U41210 (N_41210,N_39303,N_37608);
xor U41211 (N_41211,N_39405,N_38533);
nor U41212 (N_41212,N_38400,N_38779);
nand U41213 (N_41213,N_37797,N_39353);
or U41214 (N_41214,N_39210,N_37957);
and U41215 (N_41215,N_38570,N_39007);
or U41216 (N_41216,N_39547,N_39882);
and U41217 (N_41217,N_38932,N_39765);
nor U41218 (N_41218,N_39575,N_38897);
and U41219 (N_41219,N_38189,N_37871);
nor U41220 (N_41220,N_39609,N_39389);
or U41221 (N_41221,N_39147,N_38645);
xnor U41222 (N_41222,N_39775,N_38613);
xor U41223 (N_41223,N_39821,N_37994);
and U41224 (N_41224,N_39561,N_38215);
nor U41225 (N_41225,N_39772,N_39031);
nand U41226 (N_41226,N_39064,N_39010);
or U41227 (N_41227,N_37759,N_39338);
nand U41228 (N_41228,N_38396,N_37806);
nor U41229 (N_41229,N_37843,N_39617);
and U41230 (N_41230,N_38576,N_39148);
xor U41231 (N_41231,N_39529,N_38748);
and U41232 (N_41232,N_39323,N_37509);
and U41233 (N_41233,N_38990,N_39206);
or U41234 (N_41234,N_38785,N_39163);
nand U41235 (N_41235,N_39540,N_39574);
or U41236 (N_41236,N_37904,N_39115);
nand U41237 (N_41237,N_38395,N_38051);
xnor U41238 (N_41238,N_39841,N_38965);
nor U41239 (N_41239,N_37744,N_39715);
xor U41240 (N_41240,N_39272,N_39641);
nand U41241 (N_41241,N_39044,N_37589);
and U41242 (N_41242,N_37532,N_39231);
or U41243 (N_41243,N_38795,N_39205);
nand U41244 (N_41244,N_38061,N_38113);
or U41245 (N_41245,N_37725,N_39939);
and U41246 (N_41246,N_39937,N_39057);
nor U41247 (N_41247,N_39642,N_38173);
nand U41248 (N_41248,N_38252,N_38517);
xnor U41249 (N_41249,N_38600,N_39770);
nor U41250 (N_41250,N_38194,N_38182);
nor U41251 (N_41251,N_39859,N_39772);
xor U41252 (N_41252,N_37900,N_39448);
nor U41253 (N_41253,N_38689,N_39240);
nor U41254 (N_41254,N_38443,N_37945);
nor U41255 (N_41255,N_38269,N_37669);
nand U41256 (N_41256,N_39721,N_39379);
and U41257 (N_41257,N_38974,N_37755);
nand U41258 (N_41258,N_38739,N_38659);
and U41259 (N_41259,N_38324,N_37678);
or U41260 (N_41260,N_39190,N_38384);
nand U41261 (N_41261,N_39428,N_39319);
or U41262 (N_41262,N_38112,N_38124);
and U41263 (N_41263,N_38565,N_38472);
or U41264 (N_41264,N_37513,N_37587);
xor U41265 (N_41265,N_37556,N_38292);
nor U41266 (N_41266,N_39959,N_39177);
xor U41267 (N_41267,N_39081,N_39771);
and U41268 (N_41268,N_38884,N_37896);
and U41269 (N_41269,N_38949,N_38693);
or U41270 (N_41270,N_39623,N_39266);
nand U41271 (N_41271,N_39074,N_39850);
or U41272 (N_41272,N_38289,N_37677);
nor U41273 (N_41273,N_37836,N_38586);
nor U41274 (N_41274,N_38648,N_39346);
nand U41275 (N_41275,N_38307,N_38358);
xor U41276 (N_41276,N_39562,N_38718);
nand U41277 (N_41277,N_39004,N_37613);
nor U41278 (N_41278,N_37609,N_39285);
nand U41279 (N_41279,N_39807,N_39136);
xor U41280 (N_41280,N_39374,N_37551);
nand U41281 (N_41281,N_39590,N_39014);
xnor U41282 (N_41282,N_39565,N_38753);
nor U41283 (N_41283,N_38304,N_37800);
and U41284 (N_41284,N_39414,N_38674);
xor U41285 (N_41285,N_37503,N_38671);
or U41286 (N_41286,N_37863,N_37856);
or U41287 (N_41287,N_39520,N_39994);
and U41288 (N_41288,N_39207,N_38290);
and U41289 (N_41289,N_39634,N_37747);
or U41290 (N_41290,N_38106,N_38060);
xnor U41291 (N_41291,N_38291,N_38687);
or U41292 (N_41292,N_39181,N_38299);
and U41293 (N_41293,N_39171,N_37833);
xor U41294 (N_41294,N_38014,N_37500);
xor U41295 (N_41295,N_38898,N_39539);
and U41296 (N_41296,N_37545,N_39461);
and U41297 (N_41297,N_37942,N_39656);
nor U41298 (N_41298,N_38103,N_38468);
nand U41299 (N_41299,N_38533,N_38452);
xor U41300 (N_41300,N_38280,N_39234);
and U41301 (N_41301,N_39127,N_38011);
xor U41302 (N_41302,N_38078,N_37784);
xor U41303 (N_41303,N_38248,N_37719);
nand U41304 (N_41304,N_39943,N_37765);
and U41305 (N_41305,N_38925,N_38600);
and U41306 (N_41306,N_39644,N_39016);
and U41307 (N_41307,N_39354,N_38953);
or U41308 (N_41308,N_39902,N_38370);
or U41309 (N_41309,N_39319,N_38878);
nor U41310 (N_41310,N_38489,N_38277);
or U41311 (N_41311,N_37839,N_38170);
nand U41312 (N_41312,N_39299,N_38937);
or U41313 (N_41313,N_38886,N_39364);
nor U41314 (N_41314,N_38274,N_38282);
or U41315 (N_41315,N_39371,N_39477);
nand U41316 (N_41316,N_37950,N_39362);
and U41317 (N_41317,N_39675,N_38100);
nand U41318 (N_41318,N_39909,N_38021);
nand U41319 (N_41319,N_38875,N_38018);
xor U41320 (N_41320,N_38503,N_39066);
nor U41321 (N_41321,N_39988,N_39965);
or U41322 (N_41322,N_38322,N_38514);
xor U41323 (N_41323,N_39838,N_39750);
nand U41324 (N_41324,N_39135,N_39283);
nor U41325 (N_41325,N_38964,N_38124);
xnor U41326 (N_41326,N_37890,N_38352);
nor U41327 (N_41327,N_38278,N_39971);
xor U41328 (N_41328,N_39196,N_39150);
nor U41329 (N_41329,N_38308,N_39343);
nand U41330 (N_41330,N_39780,N_37820);
or U41331 (N_41331,N_38060,N_39645);
and U41332 (N_41332,N_39846,N_39722);
and U41333 (N_41333,N_38170,N_39567);
nand U41334 (N_41334,N_37998,N_38339);
or U41335 (N_41335,N_38201,N_38907);
nor U41336 (N_41336,N_39873,N_39586);
nor U41337 (N_41337,N_38898,N_38538);
nand U41338 (N_41338,N_39866,N_39663);
nor U41339 (N_41339,N_38673,N_38304);
nand U41340 (N_41340,N_39545,N_38731);
and U41341 (N_41341,N_39363,N_38862);
nor U41342 (N_41342,N_38732,N_39877);
nor U41343 (N_41343,N_37913,N_39095);
nor U41344 (N_41344,N_38974,N_37838);
or U41345 (N_41345,N_39801,N_38912);
and U41346 (N_41346,N_38875,N_38093);
xor U41347 (N_41347,N_38497,N_37520);
nand U41348 (N_41348,N_37860,N_38258);
or U41349 (N_41349,N_39560,N_37520);
and U41350 (N_41350,N_38032,N_39167);
xnor U41351 (N_41351,N_37566,N_37675);
and U41352 (N_41352,N_39452,N_38994);
and U41353 (N_41353,N_38655,N_38197);
nand U41354 (N_41354,N_39963,N_37501);
or U41355 (N_41355,N_38104,N_39525);
xor U41356 (N_41356,N_38435,N_38664);
and U41357 (N_41357,N_38109,N_39078);
or U41358 (N_41358,N_39425,N_39756);
nand U41359 (N_41359,N_38644,N_38066);
and U41360 (N_41360,N_38614,N_38506);
or U41361 (N_41361,N_39001,N_39372);
xnor U41362 (N_41362,N_39675,N_37930);
nor U41363 (N_41363,N_38680,N_39717);
xor U41364 (N_41364,N_38297,N_39697);
xnor U41365 (N_41365,N_39188,N_39584);
nand U41366 (N_41366,N_39108,N_38161);
xnor U41367 (N_41367,N_38468,N_38144);
and U41368 (N_41368,N_38115,N_38726);
nor U41369 (N_41369,N_38040,N_38256);
nand U41370 (N_41370,N_38591,N_38261);
xnor U41371 (N_41371,N_38001,N_38488);
nor U41372 (N_41372,N_39200,N_37703);
nand U41373 (N_41373,N_39730,N_39193);
xnor U41374 (N_41374,N_38338,N_38459);
nand U41375 (N_41375,N_39049,N_39643);
or U41376 (N_41376,N_37733,N_38915);
xor U41377 (N_41377,N_39444,N_39744);
or U41378 (N_41378,N_39233,N_39434);
or U41379 (N_41379,N_37993,N_38532);
nand U41380 (N_41380,N_37651,N_38191);
or U41381 (N_41381,N_39477,N_39933);
nor U41382 (N_41382,N_37743,N_38698);
or U41383 (N_41383,N_37848,N_37525);
or U41384 (N_41384,N_39840,N_38377);
nor U41385 (N_41385,N_38212,N_39214);
xor U41386 (N_41386,N_38282,N_39401);
xor U41387 (N_41387,N_39640,N_38900);
nand U41388 (N_41388,N_37795,N_39760);
xnor U41389 (N_41389,N_39113,N_38033);
or U41390 (N_41390,N_39283,N_39180);
nor U41391 (N_41391,N_38842,N_37706);
nor U41392 (N_41392,N_39481,N_38186);
nand U41393 (N_41393,N_39997,N_38814);
and U41394 (N_41394,N_39463,N_39574);
xnor U41395 (N_41395,N_38934,N_39145);
xnor U41396 (N_41396,N_38726,N_38058);
and U41397 (N_41397,N_39749,N_38119);
xor U41398 (N_41398,N_37617,N_38523);
and U41399 (N_41399,N_38731,N_39609);
or U41400 (N_41400,N_39994,N_37632);
nor U41401 (N_41401,N_37903,N_38074);
nand U41402 (N_41402,N_37686,N_37761);
nor U41403 (N_41403,N_38350,N_39721);
xnor U41404 (N_41404,N_38651,N_37502);
xor U41405 (N_41405,N_38665,N_38532);
nand U41406 (N_41406,N_39002,N_39756);
xor U41407 (N_41407,N_38447,N_38594);
xor U41408 (N_41408,N_38136,N_37902);
nor U41409 (N_41409,N_38227,N_39251);
nand U41410 (N_41410,N_38408,N_39337);
nand U41411 (N_41411,N_38647,N_38222);
xor U41412 (N_41412,N_39722,N_37717);
nor U41413 (N_41413,N_38337,N_37555);
nand U41414 (N_41414,N_37946,N_39235);
nand U41415 (N_41415,N_38224,N_38176);
nand U41416 (N_41416,N_38056,N_39073);
nor U41417 (N_41417,N_37898,N_37646);
or U41418 (N_41418,N_39469,N_37775);
xor U41419 (N_41419,N_38625,N_39214);
and U41420 (N_41420,N_37729,N_37509);
xnor U41421 (N_41421,N_38473,N_39306);
or U41422 (N_41422,N_38547,N_37745);
or U41423 (N_41423,N_37524,N_38594);
or U41424 (N_41424,N_37613,N_38712);
and U41425 (N_41425,N_38068,N_39313);
or U41426 (N_41426,N_37996,N_39029);
nand U41427 (N_41427,N_38284,N_37803);
xnor U41428 (N_41428,N_38700,N_37563);
xor U41429 (N_41429,N_39229,N_39441);
and U41430 (N_41430,N_39841,N_38600);
nor U41431 (N_41431,N_38120,N_39789);
xor U41432 (N_41432,N_38200,N_37747);
xnor U41433 (N_41433,N_37855,N_39761);
and U41434 (N_41434,N_39847,N_39227);
nand U41435 (N_41435,N_39544,N_39430);
xnor U41436 (N_41436,N_38751,N_39688);
nand U41437 (N_41437,N_38963,N_38848);
or U41438 (N_41438,N_39473,N_38334);
and U41439 (N_41439,N_37633,N_37832);
nor U41440 (N_41440,N_37958,N_38778);
or U41441 (N_41441,N_39197,N_39982);
or U41442 (N_41442,N_39332,N_38361);
and U41443 (N_41443,N_38966,N_39483);
nand U41444 (N_41444,N_38214,N_38595);
nand U41445 (N_41445,N_38645,N_39253);
nand U41446 (N_41446,N_39391,N_39791);
nor U41447 (N_41447,N_39903,N_38795);
nor U41448 (N_41448,N_39781,N_39611);
or U41449 (N_41449,N_39732,N_38218);
or U41450 (N_41450,N_38843,N_38226);
nor U41451 (N_41451,N_38307,N_38331);
or U41452 (N_41452,N_38536,N_38107);
nor U41453 (N_41453,N_38013,N_37657);
xnor U41454 (N_41454,N_38761,N_37718);
nor U41455 (N_41455,N_38622,N_39155);
nor U41456 (N_41456,N_37727,N_39283);
and U41457 (N_41457,N_39278,N_39455);
nor U41458 (N_41458,N_37663,N_39969);
xnor U41459 (N_41459,N_39758,N_37973);
xnor U41460 (N_41460,N_38424,N_37630);
nor U41461 (N_41461,N_39598,N_38138);
xnor U41462 (N_41462,N_39280,N_39816);
or U41463 (N_41463,N_39374,N_39526);
xor U41464 (N_41464,N_37736,N_38738);
and U41465 (N_41465,N_37831,N_38055);
nor U41466 (N_41466,N_37672,N_39315);
nand U41467 (N_41467,N_38294,N_39990);
and U41468 (N_41468,N_38899,N_39944);
xnor U41469 (N_41469,N_37771,N_39306);
nor U41470 (N_41470,N_39639,N_39315);
and U41471 (N_41471,N_38741,N_37903);
or U41472 (N_41472,N_38415,N_37645);
xor U41473 (N_41473,N_38981,N_39841);
nor U41474 (N_41474,N_39239,N_39614);
nor U41475 (N_41475,N_38758,N_38766);
xor U41476 (N_41476,N_38236,N_37880);
nand U41477 (N_41477,N_39887,N_38267);
nand U41478 (N_41478,N_37646,N_37870);
nand U41479 (N_41479,N_39618,N_39086);
or U41480 (N_41480,N_39926,N_39296);
nor U41481 (N_41481,N_39487,N_39724);
and U41482 (N_41482,N_38099,N_37584);
and U41483 (N_41483,N_38726,N_38307);
and U41484 (N_41484,N_39086,N_38587);
nor U41485 (N_41485,N_38225,N_38714);
or U41486 (N_41486,N_38112,N_39540);
or U41487 (N_41487,N_38036,N_39555);
nor U41488 (N_41488,N_39160,N_37880);
xor U41489 (N_41489,N_39201,N_39718);
xor U41490 (N_41490,N_39597,N_37915);
nor U41491 (N_41491,N_39904,N_39970);
xor U41492 (N_41492,N_39280,N_37918);
nand U41493 (N_41493,N_39813,N_39329);
nor U41494 (N_41494,N_39220,N_39938);
or U41495 (N_41495,N_38076,N_39205);
and U41496 (N_41496,N_37976,N_38986);
nor U41497 (N_41497,N_39386,N_39465);
and U41498 (N_41498,N_39630,N_38106);
and U41499 (N_41499,N_38271,N_38925);
nand U41500 (N_41500,N_38987,N_39240);
nor U41501 (N_41501,N_39472,N_39153);
or U41502 (N_41502,N_38624,N_39663);
and U41503 (N_41503,N_38775,N_39021);
nor U41504 (N_41504,N_38809,N_39447);
xnor U41505 (N_41505,N_39746,N_38207);
or U41506 (N_41506,N_38298,N_39580);
or U41507 (N_41507,N_37569,N_39367);
and U41508 (N_41508,N_39046,N_37806);
xnor U41509 (N_41509,N_39683,N_38109);
or U41510 (N_41510,N_37943,N_38196);
nand U41511 (N_41511,N_38247,N_39345);
or U41512 (N_41512,N_39546,N_37596);
or U41513 (N_41513,N_38316,N_39381);
nor U41514 (N_41514,N_38870,N_39765);
or U41515 (N_41515,N_39447,N_39437);
nor U41516 (N_41516,N_38701,N_39131);
and U41517 (N_41517,N_37609,N_38528);
xnor U41518 (N_41518,N_37663,N_39975);
nor U41519 (N_41519,N_37904,N_39271);
or U41520 (N_41520,N_38916,N_39682);
nor U41521 (N_41521,N_39980,N_38963);
and U41522 (N_41522,N_39934,N_37814);
and U41523 (N_41523,N_38653,N_37768);
and U41524 (N_41524,N_39400,N_39991);
or U41525 (N_41525,N_38905,N_37764);
nand U41526 (N_41526,N_38987,N_38272);
xor U41527 (N_41527,N_39885,N_38479);
nand U41528 (N_41528,N_37933,N_38250);
nor U41529 (N_41529,N_37506,N_39223);
xnor U41530 (N_41530,N_37714,N_39326);
nand U41531 (N_41531,N_39654,N_38335);
nand U41532 (N_41532,N_39326,N_39408);
nand U41533 (N_41533,N_39304,N_38087);
nand U41534 (N_41534,N_37504,N_39517);
nand U41535 (N_41535,N_37558,N_39221);
and U41536 (N_41536,N_39628,N_38777);
or U41537 (N_41537,N_38393,N_37847);
and U41538 (N_41538,N_39024,N_39163);
xor U41539 (N_41539,N_37721,N_39296);
nor U41540 (N_41540,N_38898,N_37613);
and U41541 (N_41541,N_38936,N_38429);
nand U41542 (N_41542,N_37782,N_39633);
nor U41543 (N_41543,N_37658,N_37722);
and U41544 (N_41544,N_37681,N_38719);
or U41545 (N_41545,N_38981,N_37712);
or U41546 (N_41546,N_39891,N_39363);
nor U41547 (N_41547,N_39856,N_38270);
and U41548 (N_41548,N_38031,N_37816);
xnor U41549 (N_41549,N_37576,N_37819);
and U41550 (N_41550,N_39342,N_37906);
or U41551 (N_41551,N_38893,N_38431);
or U41552 (N_41552,N_39583,N_37675);
and U41553 (N_41553,N_38230,N_39425);
and U41554 (N_41554,N_39957,N_38243);
and U41555 (N_41555,N_38136,N_39053);
nor U41556 (N_41556,N_37937,N_38014);
and U41557 (N_41557,N_38297,N_38302);
nor U41558 (N_41558,N_39263,N_37997);
nand U41559 (N_41559,N_37904,N_38322);
and U41560 (N_41560,N_39549,N_39365);
nor U41561 (N_41561,N_38686,N_39424);
and U41562 (N_41562,N_37770,N_37556);
nor U41563 (N_41563,N_39575,N_38623);
nor U41564 (N_41564,N_39533,N_39993);
nor U41565 (N_41565,N_39649,N_38330);
xnor U41566 (N_41566,N_38347,N_37789);
and U41567 (N_41567,N_38949,N_38818);
nor U41568 (N_41568,N_39549,N_37510);
nand U41569 (N_41569,N_38429,N_38956);
nand U41570 (N_41570,N_39180,N_38532);
or U41571 (N_41571,N_39454,N_39345);
or U41572 (N_41572,N_38207,N_38559);
nand U41573 (N_41573,N_39905,N_38980);
xnor U41574 (N_41574,N_37873,N_38625);
nor U41575 (N_41575,N_38118,N_39803);
and U41576 (N_41576,N_38656,N_39239);
nand U41577 (N_41577,N_37823,N_38965);
or U41578 (N_41578,N_39859,N_38145);
xor U41579 (N_41579,N_39767,N_39270);
or U41580 (N_41580,N_38906,N_39220);
xnor U41581 (N_41581,N_38825,N_39967);
nor U41582 (N_41582,N_39875,N_39587);
xnor U41583 (N_41583,N_39309,N_39018);
nor U41584 (N_41584,N_38233,N_37530);
or U41585 (N_41585,N_38201,N_38264);
nand U41586 (N_41586,N_38659,N_38899);
xor U41587 (N_41587,N_39083,N_38515);
xnor U41588 (N_41588,N_38739,N_38931);
nor U41589 (N_41589,N_37857,N_39963);
xor U41590 (N_41590,N_39283,N_38819);
and U41591 (N_41591,N_37963,N_39141);
and U41592 (N_41592,N_39412,N_38792);
nand U41593 (N_41593,N_39946,N_39687);
and U41594 (N_41594,N_38819,N_37571);
xor U41595 (N_41595,N_39151,N_38683);
and U41596 (N_41596,N_38053,N_37519);
nand U41597 (N_41597,N_39126,N_38023);
nor U41598 (N_41598,N_39567,N_37925);
xor U41599 (N_41599,N_38720,N_38251);
or U41600 (N_41600,N_38891,N_38555);
nor U41601 (N_41601,N_38944,N_37596);
xnor U41602 (N_41602,N_38151,N_38168);
nand U41603 (N_41603,N_39216,N_39479);
and U41604 (N_41604,N_38040,N_39560);
xnor U41605 (N_41605,N_38844,N_38278);
xnor U41606 (N_41606,N_39205,N_37788);
and U41607 (N_41607,N_37857,N_39893);
nand U41608 (N_41608,N_39795,N_38689);
nor U41609 (N_41609,N_39392,N_39404);
and U41610 (N_41610,N_37603,N_39096);
xnor U41611 (N_41611,N_39869,N_37763);
nand U41612 (N_41612,N_39625,N_39573);
xor U41613 (N_41613,N_37614,N_39834);
and U41614 (N_41614,N_39165,N_38030);
nor U41615 (N_41615,N_39593,N_39592);
and U41616 (N_41616,N_37891,N_38410);
nand U41617 (N_41617,N_39543,N_39427);
nor U41618 (N_41618,N_37573,N_39718);
xor U41619 (N_41619,N_38218,N_39417);
nor U41620 (N_41620,N_39669,N_39881);
nand U41621 (N_41621,N_37503,N_38752);
xor U41622 (N_41622,N_38993,N_38289);
and U41623 (N_41623,N_39107,N_39222);
nand U41624 (N_41624,N_38707,N_39524);
nand U41625 (N_41625,N_37642,N_37760);
and U41626 (N_41626,N_39027,N_38586);
or U41627 (N_41627,N_38879,N_37794);
nand U41628 (N_41628,N_39223,N_39993);
nand U41629 (N_41629,N_38498,N_38127);
xor U41630 (N_41630,N_37849,N_38889);
or U41631 (N_41631,N_38642,N_37550);
xor U41632 (N_41632,N_37832,N_37733);
and U41633 (N_41633,N_38605,N_38130);
nand U41634 (N_41634,N_39394,N_38612);
and U41635 (N_41635,N_39925,N_38311);
or U41636 (N_41636,N_37557,N_39884);
or U41637 (N_41637,N_39552,N_38821);
and U41638 (N_41638,N_39754,N_38898);
xor U41639 (N_41639,N_37535,N_37603);
or U41640 (N_41640,N_39945,N_38934);
and U41641 (N_41641,N_39765,N_39490);
xor U41642 (N_41642,N_39106,N_37548);
and U41643 (N_41643,N_38378,N_39321);
and U41644 (N_41644,N_39680,N_39702);
or U41645 (N_41645,N_38981,N_39411);
nand U41646 (N_41646,N_37850,N_38758);
nand U41647 (N_41647,N_38049,N_37870);
xnor U41648 (N_41648,N_37676,N_37841);
nor U41649 (N_41649,N_38040,N_37828);
xnor U41650 (N_41650,N_39391,N_39021);
and U41651 (N_41651,N_37663,N_39106);
xnor U41652 (N_41652,N_39908,N_37719);
nand U41653 (N_41653,N_38524,N_37863);
or U41654 (N_41654,N_38940,N_37620);
and U41655 (N_41655,N_39101,N_37671);
or U41656 (N_41656,N_39292,N_39895);
and U41657 (N_41657,N_38102,N_39416);
xor U41658 (N_41658,N_38462,N_38264);
or U41659 (N_41659,N_39980,N_37834);
xnor U41660 (N_41660,N_37996,N_39891);
nor U41661 (N_41661,N_39501,N_38290);
nand U41662 (N_41662,N_38907,N_38826);
nand U41663 (N_41663,N_39047,N_39206);
xor U41664 (N_41664,N_39741,N_37691);
nand U41665 (N_41665,N_38109,N_38494);
and U41666 (N_41666,N_37505,N_38175);
or U41667 (N_41667,N_39047,N_37951);
xor U41668 (N_41668,N_37976,N_39971);
or U41669 (N_41669,N_39960,N_38485);
nor U41670 (N_41670,N_37935,N_39573);
xor U41671 (N_41671,N_38923,N_38398);
or U41672 (N_41672,N_39091,N_39392);
and U41673 (N_41673,N_39995,N_37944);
and U41674 (N_41674,N_39514,N_38459);
nand U41675 (N_41675,N_38383,N_39656);
or U41676 (N_41676,N_39202,N_37773);
xor U41677 (N_41677,N_38047,N_39059);
or U41678 (N_41678,N_38465,N_39630);
nand U41679 (N_41679,N_38744,N_39980);
or U41680 (N_41680,N_38303,N_39876);
and U41681 (N_41681,N_38651,N_37851);
nor U41682 (N_41682,N_39691,N_38973);
or U41683 (N_41683,N_37785,N_38319);
xor U41684 (N_41684,N_38098,N_38183);
xor U41685 (N_41685,N_38069,N_39651);
and U41686 (N_41686,N_38734,N_39432);
nand U41687 (N_41687,N_38048,N_38115);
and U41688 (N_41688,N_39734,N_39485);
nand U41689 (N_41689,N_38667,N_39618);
nor U41690 (N_41690,N_38437,N_38414);
nor U41691 (N_41691,N_37867,N_37668);
and U41692 (N_41692,N_39801,N_38808);
nand U41693 (N_41693,N_38852,N_37784);
nand U41694 (N_41694,N_38307,N_37736);
xnor U41695 (N_41695,N_39780,N_38197);
nor U41696 (N_41696,N_38645,N_37805);
nand U41697 (N_41697,N_39216,N_37567);
or U41698 (N_41698,N_39233,N_39964);
nand U41699 (N_41699,N_37648,N_38652);
and U41700 (N_41700,N_39516,N_39527);
nand U41701 (N_41701,N_38341,N_37781);
nand U41702 (N_41702,N_38311,N_37904);
and U41703 (N_41703,N_39510,N_37871);
xnor U41704 (N_41704,N_38468,N_38415);
nor U41705 (N_41705,N_39747,N_37567);
nor U41706 (N_41706,N_39618,N_39182);
nor U41707 (N_41707,N_39401,N_39279);
xor U41708 (N_41708,N_38619,N_38194);
nand U41709 (N_41709,N_37592,N_37734);
or U41710 (N_41710,N_39250,N_39526);
and U41711 (N_41711,N_37502,N_37670);
nor U41712 (N_41712,N_38375,N_38525);
or U41713 (N_41713,N_37834,N_37581);
and U41714 (N_41714,N_39951,N_38878);
or U41715 (N_41715,N_38181,N_39360);
xor U41716 (N_41716,N_39941,N_38718);
and U41717 (N_41717,N_38707,N_38050);
and U41718 (N_41718,N_38351,N_39595);
nand U41719 (N_41719,N_39221,N_39967);
or U41720 (N_41720,N_39690,N_39126);
xor U41721 (N_41721,N_37816,N_39518);
or U41722 (N_41722,N_39543,N_37994);
xor U41723 (N_41723,N_38403,N_38431);
and U41724 (N_41724,N_37689,N_37888);
or U41725 (N_41725,N_37605,N_37637);
nand U41726 (N_41726,N_38345,N_38304);
nor U41727 (N_41727,N_39219,N_39744);
nand U41728 (N_41728,N_37778,N_39388);
xnor U41729 (N_41729,N_38423,N_39311);
nor U41730 (N_41730,N_39521,N_39194);
nor U41731 (N_41731,N_38156,N_37544);
xnor U41732 (N_41732,N_39079,N_37965);
nand U41733 (N_41733,N_38760,N_39247);
xor U41734 (N_41734,N_39680,N_39065);
nor U41735 (N_41735,N_39398,N_37694);
and U41736 (N_41736,N_39887,N_37834);
or U41737 (N_41737,N_39548,N_39229);
nor U41738 (N_41738,N_38048,N_39206);
nand U41739 (N_41739,N_38383,N_38288);
nor U41740 (N_41740,N_37687,N_37829);
nor U41741 (N_41741,N_38929,N_37890);
and U41742 (N_41742,N_38978,N_37689);
nand U41743 (N_41743,N_39415,N_39618);
nand U41744 (N_41744,N_38146,N_38777);
or U41745 (N_41745,N_39106,N_39968);
xnor U41746 (N_41746,N_37980,N_38417);
and U41747 (N_41747,N_39120,N_38613);
nor U41748 (N_41748,N_39117,N_39100);
or U41749 (N_41749,N_37789,N_38823);
and U41750 (N_41750,N_37902,N_38949);
nor U41751 (N_41751,N_39434,N_38639);
xnor U41752 (N_41752,N_38945,N_38348);
or U41753 (N_41753,N_38537,N_39316);
xnor U41754 (N_41754,N_38543,N_38395);
xnor U41755 (N_41755,N_38531,N_37895);
xor U41756 (N_41756,N_38982,N_38836);
nor U41757 (N_41757,N_38661,N_38788);
or U41758 (N_41758,N_37884,N_37983);
nor U41759 (N_41759,N_37905,N_39338);
xor U41760 (N_41760,N_38460,N_39063);
and U41761 (N_41761,N_39917,N_39008);
or U41762 (N_41762,N_38343,N_37640);
nand U41763 (N_41763,N_39212,N_37851);
xor U41764 (N_41764,N_39904,N_37848);
nand U41765 (N_41765,N_39492,N_38200);
nand U41766 (N_41766,N_37992,N_37611);
nor U41767 (N_41767,N_38216,N_38916);
nor U41768 (N_41768,N_38352,N_38335);
nand U41769 (N_41769,N_39216,N_38438);
nor U41770 (N_41770,N_39346,N_38233);
or U41771 (N_41771,N_39214,N_38231);
or U41772 (N_41772,N_39710,N_39464);
nor U41773 (N_41773,N_39016,N_39325);
nand U41774 (N_41774,N_39631,N_37919);
nand U41775 (N_41775,N_37628,N_38186);
xnor U41776 (N_41776,N_39477,N_37841);
nand U41777 (N_41777,N_38513,N_39379);
nor U41778 (N_41778,N_38172,N_38888);
nand U41779 (N_41779,N_38708,N_38022);
nand U41780 (N_41780,N_39025,N_38797);
nand U41781 (N_41781,N_38281,N_39941);
nor U41782 (N_41782,N_39304,N_37794);
nor U41783 (N_41783,N_39259,N_38217);
or U41784 (N_41784,N_39626,N_39677);
nand U41785 (N_41785,N_38168,N_39205);
or U41786 (N_41786,N_39557,N_38937);
nand U41787 (N_41787,N_39785,N_39230);
nor U41788 (N_41788,N_39477,N_38686);
nor U41789 (N_41789,N_38140,N_38825);
or U41790 (N_41790,N_38081,N_37791);
and U41791 (N_41791,N_37636,N_39024);
nand U41792 (N_41792,N_38448,N_39550);
xor U41793 (N_41793,N_39202,N_39595);
xnor U41794 (N_41794,N_38512,N_38339);
nor U41795 (N_41795,N_39065,N_39894);
nor U41796 (N_41796,N_39006,N_38868);
or U41797 (N_41797,N_38238,N_38659);
and U41798 (N_41798,N_38095,N_38885);
nor U41799 (N_41799,N_39592,N_38032);
nor U41800 (N_41800,N_39281,N_37708);
nor U41801 (N_41801,N_38157,N_39918);
nor U41802 (N_41802,N_38402,N_38644);
nand U41803 (N_41803,N_39148,N_37777);
or U41804 (N_41804,N_39363,N_37901);
xor U41805 (N_41805,N_38503,N_39023);
nor U41806 (N_41806,N_38158,N_39375);
nor U41807 (N_41807,N_38126,N_39138);
xor U41808 (N_41808,N_38433,N_37794);
or U41809 (N_41809,N_39180,N_38189);
nor U41810 (N_41810,N_38848,N_38571);
or U41811 (N_41811,N_38193,N_39875);
and U41812 (N_41812,N_39710,N_39430);
or U41813 (N_41813,N_37765,N_38311);
nor U41814 (N_41814,N_39320,N_39437);
nor U41815 (N_41815,N_39399,N_38782);
and U41816 (N_41816,N_37650,N_38207);
nand U41817 (N_41817,N_37976,N_39050);
or U41818 (N_41818,N_39446,N_39849);
xor U41819 (N_41819,N_38401,N_39064);
and U41820 (N_41820,N_39487,N_38377);
nor U41821 (N_41821,N_38517,N_39736);
xor U41822 (N_41822,N_39225,N_37923);
xnor U41823 (N_41823,N_39467,N_38325);
nand U41824 (N_41824,N_39924,N_38374);
or U41825 (N_41825,N_38371,N_38587);
and U41826 (N_41826,N_39526,N_37538);
nor U41827 (N_41827,N_39954,N_39337);
nand U41828 (N_41828,N_39230,N_39593);
nor U41829 (N_41829,N_38574,N_38097);
nor U41830 (N_41830,N_37718,N_38987);
nand U41831 (N_41831,N_39537,N_37568);
nand U41832 (N_41832,N_38734,N_38927);
xnor U41833 (N_41833,N_38368,N_38692);
nand U41834 (N_41834,N_38337,N_39085);
and U41835 (N_41835,N_39212,N_38704);
and U41836 (N_41836,N_37810,N_38343);
or U41837 (N_41837,N_39309,N_37618);
nand U41838 (N_41838,N_39502,N_39792);
nand U41839 (N_41839,N_38341,N_37520);
xnor U41840 (N_41840,N_39913,N_37855);
and U41841 (N_41841,N_38770,N_39651);
nand U41842 (N_41842,N_37872,N_38922);
nand U41843 (N_41843,N_39750,N_37800);
nand U41844 (N_41844,N_38780,N_39956);
or U41845 (N_41845,N_39692,N_39749);
or U41846 (N_41846,N_37908,N_39619);
and U41847 (N_41847,N_39182,N_38661);
and U41848 (N_41848,N_38081,N_37926);
nand U41849 (N_41849,N_38605,N_38088);
nand U41850 (N_41850,N_39256,N_38961);
xor U41851 (N_41851,N_38889,N_39940);
or U41852 (N_41852,N_39067,N_39246);
xor U41853 (N_41853,N_39422,N_39652);
and U41854 (N_41854,N_38270,N_38941);
xnor U41855 (N_41855,N_38994,N_37674);
nand U41856 (N_41856,N_39660,N_38191);
nand U41857 (N_41857,N_39008,N_39461);
xnor U41858 (N_41858,N_38601,N_39581);
nand U41859 (N_41859,N_37837,N_39573);
nand U41860 (N_41860,N_39072,N_37630);
and U41861 (N_41861,N_38625,N_38634);
xnor U41862 (N_41862,N_38682,N_38139);
and U41863 (N_41863,N_38317,N_39209);
nor U41864 (N_41864,N_39255,N_37681);
nand U41865 (N_41865,N_38425,N_39144);
and U41866 (N_41866,N_38042,N_38684);
nor U41867 (N_41867,N_38614,N_37768);
xnor U41868 (N_41868,N_37901,N_39126);
and U41869 (N_41869,N_39082,N_37799);
xor U41870 (N_41870,N_39685,N_39617);
nor U41871 (N_41871,N_38969,N_38032);
or U41872 (N_41872,N_37979,N_39475);
or U41873 (N_41873,N_38598,N_39405);
nor U41874 (N_41874,N_39161,N_37529);
nand U41875 (N_41875,N_37795,N_39304);
or U41876 (N_41876,N_37609,N_39024);
or U41877 (N_41877,N_37901,N_39099);
or U41878 (N_41878,N_38341,N_39645);
nor U41879 (N_41879,N_39888,N_38193);
nand U41880 (N_41880,N_37991,N_37545);
nor U41881 (N_41881,N_38424,N_37815);
or U41882 (N_41882,N_39792,N_39755);
nor U41883 (N_41883,N_37506,N_39015);
nand U41884 (N_41884,N_38642,N_38637);
nor U41885 (N_41885,N_39797,N_38821);
nor U41886 (N_41886,N_38565,N_38627);
xor U41887 (N_41887,N_37679,N_39097);
xor U41888 (N_41888,N_38728,N_39163);
nor U41889 (N_41889,N_37606,N_39500);
or U41890 (N_41890,N_37803,N_38582);
xnor U41891 (N_41891,N_38912,N_39755);
or U41892 (N_41892,N_39437,N_38181);
and U41893 (N_41893,N_39505,N_38474);
and U41894 (N_41894,N_37994,N_37934);
or U41895 (N_41895,N_39478,N_38858);
nor U41896 (N_41896,N_39155,N_38183);
or U41897 (N_41897,N_37588,N_39318);
xor U41898 (N_41898,N_39510,N_39421);
and U41899 (N_41899,N_39808,N_39900);
or U41900 (N_41900,N_38604,N_38623);
and U41901 (N_41901,N_37735,N_39552);
nand U41902 (N_41902,N_38088,N_38249);
xor U41903 (N_41903,N_39794,N_38750);
nor U41904 (N_41904,N_39281,N_38387);
nand U41905 (N_41905,N_38245,N_39005);
or U41906 (N_41906,N_39204,N_38590);
xor U41907 (N_41907,N_39336,N_38332);
nor U41908 (N_41908,N_38338,N_38687);
nand U41909 (N_41909,N_38655,N_37563);
or U41910 (N_41910,N_39748,N_37740);
nor U41911 (N_41911,N_38861,N_39918);
nand U41912 (N_41912,N_37862,N_38122);
and U41913 (N_41913,N_39337,N_38930);
nor U41914 (N_41914,N_37525,N_39016);
and U41915 (N_41915,N_39508,N_37870);
or U41916 (N_41916,N_39410,N_38165);
nor U41917 (N_41917,N_37743,N_38471);
xor U41918 (N_41918,N_38280,N_39721);
nand U41919 (N_41919,N_38896,N_38984);
nand U41920 (N_41920,N_39809,N_37663);
or U41921 (N_41921,N_38140,N_39385);
and U41922 (N_41922,N_39440,N_39050);
and U41923 (N_41923,N_39645,N_39029);
nand U41924 (N_41924,N_38913,N_38430);
and U41925 (N_41925,N_38478,N_38290);
nor U41926 (N_41926,N_38108,N_39177);
nor U41927 (N_41927,N_38948,N_39425);
nor U41928 (N_41928,N_39829,N_38685);
nand U41929 (N_41929,N_37685,N_38905);
nand U41930 (N_41930,N_37892,N_38118);
xor U41931 (N_41931,N_38964,N_37667);
xnor U41932 (N_41932,N_38946,N_37907);
or U41933 (N_41933,N_38567,N_39072);
and U41934 (N_41934,N_37713,N_38836);
and U41935 (N_41935,N_39474,N_37903);
and U41936 (N_41936,N_39484,N_38663);
nor U41937 (N_41937,N_37818,N_39139);
and U41938 (N_41938,N_39405,N_39972);
nand U41939 (N_41939,N_39738,N_39914);
nor U41940 (N_41940,N_38806,N_38743);
nor U41941 (N_41941,N_37830,N_39174);
nand U41942 (N_41942,N_37581,N_38396);
nor U41943 (N_41943,N_38838,N_37869);
nand U41944 (N_41944,N_37551,N_38472);
nor U41945 (N_41945,N_39563,N_39974);
or U41946 (N_41946,N_37739,N_38491);
and U41947 (N_41947,N_39157,N_38494);
xor U41948 (N_41948,N_39370,N_39494);
nor U41949 (N_41949,N_39986,N_38625);
nor U41950 (N_41950,N_39756,N_37508);
or U41951 (N_41951,N_39145,N_39660);
or U41952 (N_41952,N_39110,N_37870);
and U41953 (N_41953,N_39468,N_39827);
or U41954 (N_41954,N_38753,N_39416);
xor U41955 (N_41955,N_39076,N_39357);
nand U41956 (N_41956,N_39285,N_38989);
and U41957 (N_41957,N_37745,N_37652);
and U41958 (N_41958,N_38363,N_39674);
and U41959 (N_41959,N_37981,N_38646);
or U41960 (N_41960,N_39144,N_38120);
or U41961 (N_41961,N_37868,N_37826);
nor U41962 (N_41962,N_37511,N_39693);
xnor U41963 (N_41963,N_39125,N_37828);
and U41964 (N_41964,N_37814,N_39794);
and U41965 (N_41965,N_39299,N_39339);
nand U41966 (N_41966,N_38667,N_38802);
or U41967 (N_41967,N_38753,N_37532);
nand U41968 (N_41968,N_39592,N_38344);
and U41969 (N_41969,N_39859,N_39075);
nand U41970 (N_41970,N_39296,N_38377);
nand U41971 (N_41971,N_38187,N_37720);
nand U41972 (N_41972,N_39582,N_39229);
nand U41973 (N_41973,N_38543,N_39319);
nand U41974 (N_41974,N_38979,N_38915);
nor U41975 (N_41975,N_37762,N_39694);
and U41976 (N_41976,N_38656,N_39372);
or U41977 (N_41977,N_38677,N_39287);
or U41978 (N_41978,N_39844,N_39817);
nand U41979 (N_41979,N_38848,N_37748);
nor U41980 (N_41980,N_37911,N_38585);
xor U41981 (N_41981,N_39466,N_39683);
nor U41982 (N_41982,N_39618,N_38369);
nor U41983 (N_41983,N_37610,N_38758);
and U41984 (N_41984,N_38288,N_38374);
nor U41985 (N_41985,N_38510,N_38595);
nand U41986 (N_41986,N_39490,N_39340);
or U41987 (N_41987,N_38754,N_37581);
or U41988 (N_41988,N_38314,N_38176);
or U41989 (N_41989,N_38714,N_37855);
nand U41990 (N_41990,N_38696,N_39876);
or U41991 (N_41991,N_37694,N_37978);
or U41992 (N_41992,N_38021,N_38920);
or U41993 (N_41993,N_39625,N_39859);
xnor U41994 (N_41994,N_37790,N_39735);
nor U41995 (N_41995,N_39482,N_37965);
or U41996 (N_41996,N_38067,N_38239);
nor U41997 (N_41997,N_39761,N_38385);
and U41998 (N_41998,N_37952,N_39457);
or U41999 (N_41999,N_39933,N_38850);
and U42000 (N_42000,N_39198,N_38518);
nand U42001 (N_42001,N_37630,N_38736);
or U42002 (N_42002,N_38635,N_39022);
nand U42003 (N_42003,N_38677,N_39208);
or U42004 (N_42004,N_39610,N_39122);
and U42005 (N_42005,N_38737,N_38662);
nand U42006 (N_42006,N_39738,N_37680);
xor U42007 (N_42007,N_37637,N_38052);
nor U42008 (N_42008,N_39178,N_38851);
or U42009 (N_42009,N_38021,N_37561);
nand U42010 (N_42010,N_39333,N_38446);
xnor U42011 (N_42011,N_38019,N_38058);
xor U42012 (N_42012,N_38007,N_39835);
xnor U42013 (N_42013,N_39810,N_39216);
xor U42014 (N_42014,N_39488,N_39654);
and U42015 (N_42015,N_38158,N_38141);
xnor U42016 (N_42016,N_38855,N_39625);
or U42017 (N_42017,N_39094,N_38682);
nor U42018 (N_42018,N_38549,N_37587);
and U42019 (N_42019,N_39764,N_37963);
and U42020 (N_42020,N_39570,N_37812);
or U42021 (N_42021,N_38418,N_37999);
nor U42022 (N_42022,N_38267,N_38654);
xnor U42023 (N_42023,N_37692,N_38793);
nor U42024 (N_42024,N_39572,N_39433);
xor U42025 (N_42025,N_39969,N_39029);
nand U42026 (N_42026,N_39752,N_38192);
nand U42027 (N_42027,N_38226,N_38172);
and U42028 (N_42028,N_38054,N_38585);
xnor U42029 (N_42029,N_39680,N_37671);
or U42030 (N_42030,N_38545,N_39475);
and U42031 (N_42031,N_39204,N_39342);
or U42032 (N_42032,N_38165,N_38237);
or U42033 (N_42033,N_38724,N_37960);
or U42034 (N_42034,N_38747,N_37715);
nand U42035 (N_42035,N_39993,N_39538);
nor U42036 (N_42036,N_38332,N_38002);
nor U42037 (N_42037,N_39378,N_38906);
or U42038 (N_42038,N_39972,N_38850);
or U42039 (N_42039,N_39576,N_37733);
nor U42040 (N_42040,N_39583,N_39890);
nor U42041 (N_42041,N_37543,N_37869);
nand U42042 (N_42042,N_39288,N_39121);
xnor U42043 (N_42043,N_38339,N_38801);
nand U42044 (N_42044,N_38538,N_38891);
nor U42045 (N_42045,N_38186,N_38477);
nor U42046 (N_42046,N_38112,N_38501);
and U42047 (N_42047,N_38091,N_37695);
nor U42048 (N_42048,N_39673,N_39729);
xor U42049 (N_42049,N_39986,N_38489);
xnor U42050 (N_42050,N_39911,N_39541);
nor U42051 (N_42051,N_38376,N_38884);
or U42052 (N_42052,N_38139,N_38868);
nor U42053 (N_42053,N_37605,N_39756);
nor U42054 (N_42054,N_39878,N_39924);
nor U42055 (N_42055,N_39056,N_37602);
nand U42056 (N_42056,N_39064,N_38160);
xnor U42057 (N_42057,N_39700,N_39606);
xor U42058 (N_42058,N_39337,N_38153);
nor U42059 (N_42059,N_37560,N_39401);
nand U42060 (N_42060,N_39013,N_37967);
nand U42061 (N_42061,N_39253,N_39700);
xnor U42062 (N_42062,N_37951,N_39727);
and U42063 (N_42063,N_39365,N_38135);
nor U42064 (N_42064,N_39257,N_39969);
nand U42065 (N_42065,N_38228,N_39620);
and U42066 (N_42066,N_39398,N_39893);
or U42067 (N_42067,N_38765,N_37809);
and U42068 (N_42068,N_37798,N_39090);
and U42069 (N_42069,N_39962,N_38718);
nand U42070 (N_42070,N_37580,N_37516);
xor U42071 (N_42071,N_38282,N_39538);
and U42072 (N_42072,N_39071,N_38426);
xnor U42073 (N_42073,N_39867,N_39720);
nor U42074 (N_42074,N_39147,N_38848);
nand U42075 (N_42075,N_37838,N_38650);
nand U42076 (N_42076,N_38830,N_39071);
or U42077 (N_42077,N_37640,N_39628);
nand U42078 (N_42078,N_38807,N_39956);
and U42079 (N_42079,N_38459,N_39870);
nand U42080 (N_42080,N_38640,N_38609);
nor U42081 (N_42081,N_38312,N_39679);
xnor U42082 (N_42082,N_39312,N_39972);
nor U42083 (N_42083,N_37990,N_38551);
xnor U42084 (N_42084,N_39216,N_39750);
and U42085 (N_42085,N_38155,N_39285);
nor U42086 (N_42086,N_39114,N_38303);
xor U42087 (N_42087,N_39822,N_39794);
or U42088 (N_42088,N_38338,N_38053);
nor U42089 (N_42089,N_38818,N_38620);
xnor U42090 (N_42090,N_39879,N_39719);
nand U42091 (N_42091,N_39159,N_38258);
nand U42092 (N_42092,N_39316,N_37785);
or U42093 (N_42093,N_38041,N_38289);
nor U42094 (N_42094,N_39399,N_39968);
or U42095 (N_42095,N_38547,N_37863);
xnor U42096 (N_42096,N_37553,N_37502);
and U42097 (N_42097,N_37706,N_39507);
or U42098 (N_42098,N_38484,N_38127);
or U42099 (N_42099,N_39970,N_39206);
nand U42100 (N_42100,N_38079,N_38200);
and U42101 (N_42101,N_39314,N_38592);
nor U42102 (N_42102,N_37878,N_39289);
nor U42103 (N_42103,N_39818,N_37794);
nor U42104 (N_42104,N_37846,N_38014);
nand U42105 (N_42105,N_39169,N_38401);
or U42106 (N_42106,N_39563,N_39105);
nand U42107 (N_42107,N_39806,N_38837);
nand U42108 (N_42108,N_38354,N_39576);
nor U42109 (N_42109,N_39352,N_37884);
nor U42110 (N_42110,N_38962,N_38253);
and U42111 (N_42111,N_39730,N_38721);
and U42112 (N_42112,N_37551,N_39317);
or U42113 (N_42113,N_38663,N_39573);
xnor U42114 (N_42114,N_39930,N_38558);
xnor U42115 (N_42115,N_39764,N_38974);
xnor U42116 (N_42116,N_39332,N_39287);
xnor U42117 (N_42117,N_39637,N_37880);
nand U42118 (N_42118,N_38765,N_38528);
xor U42119 (N_42119,N_39365,N_39264);
xor U42120 (N_42120,N_38805,N_39365);
or U42121 (N_42121,N_38102,N_39388);
nor U42122 (N_42122,N_38426,N_39964);
nor U42123 (N_42123,N_37837,N_37589);
or U42124 (N_42124,N_39583,N_39117);
xnor U42125 (N_42125,N_38885,N_38695);
nand U42126 (N_42126,N_39536,N_37543);
xnor U42127 (N_42127,N_39711,N_38238);
and U42128 (N_42128,N_39749,N_38210);
and U42129 (N_42129,N_37622,N_39179);
or U42130 (N_42130,N_39933,N_37947);
xnor U42131 (N_42131,N_38883,N_38577);
nand U42132 (N_42132,N_39695,N_38598);
nor U42133 (N_42133,N_38387,N_37620);
nor U42134 (N_42134,N_37646,N_39334);
nor U42135 (N_42135,N_39340,N_38225);
and U42136 (N_42136,N_38561,N_38241);
nand U42137 (N_42137,N_39285,N_37776);
xor U42138 (N_42138,N_38702,N_37611);
xnor U42139 (N_42139,N_37875,N_39973);
nor U42140 (N_42140,N_39768,N_38854);
nor U42141 (N_42141,N_39393,N_38653);
and U42142 (N_42142,N_38213,N_37729);
and U42143 (N_42143,N_39135,N_37906);
or U42144 (N_42144,N_38234,N_37926);
nand U42145 (N_42145,N_39519,N_37929);
xor U42146 (N_42146,N_37580,N_37897);
and U42147 (N_42147,N_38640,N_38304);
xnor U42148 (N_42148,N_38747,N_38174);
nand U42149 (N_42149,N_39751,N_37894);
or U42150 (N_42150,N_38309,N_39586);
nand U42151 (N_42151,N_38972,N_37537);
nand U42152 (N_42152,N_38806,N_38202);
or U42153 (N_42153,N_39281,N_39801);
and U42154 (N_42154,N_37869,N_38585);
xor U42155 (N_42155,N_39944,N_38777);
nand U42156 (N_42156,N_38683,N_38285);
or U42157 (N_42157,N_39543,N_38421);
and U42158 (N_42158,N_39307,N_37678);
xor U42159 (N_42159,N_38798,N_38629);
nor U42160 (N_42160,N_39291,N_38285);
nand U42161 (N_42161,N_38914,N_39592);
xor U42162 (N_42162,N_37991,N_39049);
or U42163 (N_42163,N_39577,N_39026);
nand U42164 (N_42164,N_39152,N_38319);
nor U42165 (N_42165,N_39730,N_39898);
nand U42166 (N_42166,N_37890,N_38399);
and U42167 (N_42167,N_39485,N_37859);
nor U42168 (N_42168,N_38023,N_37598);
and U42169 (N_42169,N_37667,N_37595);
and U42170 (N_42170,N_38465,N_39439);
or U42171 (N_42171,N_39153,N_38291);
or U42172 (N_42172,N_37839,N_39471);
nand U42173 (N_42173,N_39147,N_38397);
and U42174 (N_42174,N_39174,N_39875);
or U42175 (N_42175,N_39456,N_38532);
nand U42176 (N_42176,N_37562,N_37914);
or U42177 (N_42177,N_39332,N_37609);
nor U42178 (N_42178,N_39406,N_37868);
or U42179 (N_42179,N_39052,N_38364);
nor U42180 (N_42180,N_38666,N_39883);
or U42181 (N_42181,N_39254,N_39625);
or U42182 (N_42182,N_39907,N_39985);
xor U42183 (N_42183,N_39269,N_38959);
nor U42184 (N_42184,N_39029,N_39244);
nand U42185 (N_42185,N_38325,N_38683);
xnor U42186 (N_42186,N_38443,N_38353);
xnor U42187 (N_42187,N_39001,N_38379);
nand U42188 (N_42188,N_37740,N_37731);
nor U42189 (N_42189,N_39100,N_39867);
nand U42190 (N_42190,N_39492,N_39958);
nor U42191 (N_42191,N_38182,N_38708);
and U42192 (N_42192,N_38343,N_38374);
or U42193 (N_42193,N_38566,N_38516);
and U42194 (N_42194,N_38079,N_38247);
and U42195 (N_42195,N_37913,N_38683);
nor U42196 (N_42196,N_37518,N_39176);
and U42197 (N_42197,N_37695,N_38313);
and U42198 (N_42198,N_38357,N_38966);
or U42199 (N_42199,N_39581,N_38266);
and U42200 (N_42200,N_38895,N_38871);
nor U42201 (N_42201,N_39395,N_39387);
nand U42202 (N_42202,N_38726,N_37690);
and U42203 (N_42203,N_39404,N_39370);
and U42204 (N_42204,N_38255,N_39244);
or U42205 (N_42205,N_38705,N_39076);
and U42206 (N_42206,N_39367,N_38933);
or U42207 (N_42207,N_38093,N_38865);
nand U42208 (N_42208,N_38156,N_39584);
nand U42209 (N_42209,N_38110,N_38089);
and U42210 (N_42210,N_37517,N_38521);
nand U42211 (N_42211,N_38642,N_37706);
or U42212 (N_42212,N_39034,N_38459);
xnor U42213 (N_42213,N_38053,N_38775);
or U42214 (N_42214,N_37779,N_39499);
and U42215 (N_42215,N_38302,N_38803);
nor U42216 (N_42216,N_38641,N_38934);
and U42217 (N_42217,N_38423,N_38517);
xnor U42218 (N_42218,N_39335,N_38894);
nand U42219 (N_42219,N_38294,N_38997);
xnor U42220 (N_42220,N_38397,N_38945);
xor U42221 (N_42221,N_38123,N_39946);
nand U42222 (N_42222,N_39367,N_39180);
nand U42223 (N_42223,N_39536,N_37835);
or U42224 (N_42224,N_38193,N_39699);
xor U42225 (N_42225,N_37567,N_37822);
nor U42226 (N_42226,N_39423,N_38731);
xor U42227 (N_42227,N_39350,N_37954);
nor U42228 (N_42228,N_37856,N_39278);
nor U42229 (N_42229,N_39876,N_38577);
nor U42230 (N_42230,N_39530,N_39565);
xnor U42231 (N_42231,N_39667,N_37890);
xor U42232 (N_42232,N_39025,N_38373);
and U42233 (N_42233,N_38434,N_39700);
xor U42234 (N_42234,N_39386,N_39871);
nand U42235 (N_42235,N_39285,N_39054);
xor U42236 (N_42236,N_39059,N_39750);
nand U42237 (N_42237,N_39471,N_39973);
and U42238 (N_42238,N_38071,N_38309);
nor U42239 (N_42239,N_37783,N_37754);
nor U42240 (N_42240,N_39103,N_38765);
and U42241 (N_42241,N_39871,N_39676);
and U42242 (N_42242,N_38000,N_37588);
nand U42243 (N_42243,N_38945,N_38754);
nand U42244 (N_42244,N_38991,N_39731);
nand U42245 (N_42245,N_39449,N_39523);
or U42246 (N_42246,N_38814,N_38901);
xor U42247 (N_42247,N_39039,N_37674);
or U42248 (N_42248,N_39219,N_39280);
nor U42249 (N_42249,N_39002,N_37779);
and U42250 (N_42250,N_39197,N_38484);
or U42251 (N_42251,N_37780,N_38931);
nor U42252 (N_42252,N_37867,N_37701);
nand U42253 (N_42253,N_38182,N_37565);
and U42254 (N_42254,N_38494,N_38375);
or U42255 (N_42255,N_38382,N_39417);
nand U42256 (N_42256,N_37808,N_38654);
or U42257 (N_42257,N_38861,N_39058);
and U42258 (N_42258,N_37656,N_39761);
nand U42259 (N_42259,N_37764,N_38362);
nor U42260 (N_42260,N_39713,N_39998);
nand U42261 (N_42261,N_39700,N_39740);
nor U42262 (N_42262,N_39352,N_38250);
xor U42263 (N_42263,N_37891,N_37751);
nor U42264 (N_42264,N_39083,N_38849);
nand U42265 (N_42265,N_39688,N_38887);
xor U42266 (N_42266,N_37698,N_39621);
nor U42267 (N_42267,N_39598,N_37816);
and U42268 (N_42268,N_39137,N_38865);
xor U42269 (N_42269,N_39480,N_38231);
or U42270 (N_42270,N_39827,N_38773);
nand U42271 (N_42271,N_38753,N_37593);
or U42272 (N_42272,N_38928,N_37988);
and U42273 (N_42273,N_37612,N_39500);
and U42274 (N_42274,N_38286,N_39189);
nand U42275 (N_42275,N_37996,N_38252);
and U42276 (N_42276,N_38902,N_39212);
and U42277 (N_42277,N_37915,N_37505);
nand U42278 (N_42278,N_38039,N_37647);
or U42279 (N_42279,N_38489,N_38892);
xnor U42280 (N_42280,N_38518,N_39739);
xor U42281 (N_42281,N_39171,N_37543);
xor U42282 (N_42282,N_38377,N_39145);
xnor U42283 (N_42283,N_37690,N_37682);
or U42284 (N_42284,N_38338,N_38626);
xor U42285 (N_42285,N_39969,N_38689);
nand U42286 (N_42286,N_39444,N_39735);
nor U42287 (N_42287,N_38043,N_37819);
xnor U42288 (N_42288,N_39408,N_39690);
nor U42289 (N_42289,N_38148,N_39633);
nand U42290 (N_42290,N_38475,N_38159);
or U42291 (N_42291,N_39556,N_38282);
or U42292 (N_42292,N_38249,N_39250);
nor U42293 (N_42293,N_39305,N_37724);
or U42294 (N_42294,N_38115,N_39671);
or U42295 (N_42295,N_38813,N_39638);
nor U42296 (N_42296,N_37922,N_39207);
nand U42297 (N_42297,N_39146,N_39904);
and U42298 (N_42298,N_37550,N_37779);
or U42299 (N_42299,N_39783,N_39533);
or U42300 (N_42300,N_37935,N_37893);
nand U42301 (N_42301,N_38859,N_39993);
and U42302 (N_42302,N_38592,N_39382);
nand U42303 (N_42303,N_39389,N_39533);
nor U42304 (N_42304,N_39750,N_37995);
nand U42305 (N_42305,N_38436,N_39134);
or U42306 (N_42306,N_39755,N_37573);
and U42307 (N_42307,N_38078,N_39606);
xor U42308 (N_42308,N_39353,N_38223);
xnor U42309 (N_42309,N_38723,N_39515);
nor U42310 (N_42310,N_39552,N_37694);
nor U42311 (N_42311,N_39318,N_39389);
and U42312 (N_42312,N_39439,N_39062);
xor U42313 (N_42313,N_39807,N_38360);
nand U42314 (N_42314,N_38304,N_39367);
or U42315 (N_42315,N_38583,N_38615);
nand U42316 (N_42316,N_39414,N_39706);
or U42317 (N_42317,N_39073,N_39769);
nor U42318 (N_42318,N_37812,N_38536);
and U42319 (N_42319,N_37646,N_37770);
nand U42320 (N_42320,N_37642,N_39436);
and U42321 (N_42321,N_39485,N_39980);
or U42322 (N_42322,N_37868,N_37824);
nand U42323 (N_42323,N_38226,N_38570);
and U42324 (N_42324,N_37743,N_39379);
nand U42325 (N_42325,N_37903,N_39874);
and U42326 (N_42326,N_39510,N_38261);
nand U42327 (N_42327,N_39862,N_38311);
and U42328 (N_42328,N_38219,N_39887);
nor U42329 (N_42329,N_37604,N_37503);
nor U42330 (N_42330,N_37671,N_38693);
xor U42331 (N_42331,N_39778,N_38716);
nand U42332 (N_42332,N_39411,N_37818);
or U42333 (N_42333,N_37566,N_39301);
xor U42334 (N_42334,N_39359,N_38641);
and U42335 (N_42335,N_39280,N_39010);
and U42336 (N_42336,N_39999,N_39918);
xnor U42337 (N_42337,N_39479,N_39258);
and U42338 (N_42338,N_38295,N_39036);
and U42339 (N_42339,N_37564,N_39631);
nand U42340 (N_42340,N_39143,N_39932);
nor U42341 (N_42341,N_37929,N_39059);
nor U42342 (N_42342,N_38288,N_38997);
or U42343 (N_42343,N_39135,N_39086);
xor U42344 (N_42344,N_38331,N_39983);
xnor U42345 (N_42345,N_38282,N_38836);
or U42346 (N_42346,N_39928,N_39937);
or U42347 (N_42347,N_38604,N_38238);
and U42348 (N_42348,N_38785,N_39645);
xor U42349 (N_42349,N_38971,N_38999);
nand U42350 (N_42350,N_39452,N_38406);
xor U42351 (N_42351,N_38590,N_38768);
nand U42352 (N_42352,N_37792,N_38691);
xor U42353 (N_42353,N_39651,N_38969);
or U42354 (N_42354,N_38898,N_37510);
or U42355 (N_42355,N_38361,N_39256);
or U42356 (N_42356,N_38466,N_38825);
xor U42357 (N_42357,N_39224,N_39320);
xor U42358 (N_42358,N_38807,N_38193);
nor U42359 (N_42359,N_38682,N_39222);
and U42360 (N_42360,N_37595,N_38965);
nand U42361 (N_42361,N_38931,N_38066);
xnor U42362 (N_42362,N_39969,N_39680);
nand U42363 (N_42363,N_37540,N_38670);
and U42364 (N_42364,N_38708,N_38498);
nor U42365 (N_42365,N_38078,N_39644);
or U42366 (N_42366,N_37658,N_37998);
nand U42367 (N_42367,N_38287,N_38410);
nand U42368 (N_42368,N_39769,N_39135);
and U42369 (N_42369,N_37528,N_39300);
xnor U42370 (N_42370,N_39565,N_39860);
nor U42371 (N_42371,N_37774,N_39121);
nand U42372 (N_42372,N_38025,N_38697);
nor U42373 (N_42373,N_37750,N_37978);
xnor U42374 (N_42374,N_39277,N_38975);
and U42375 (N_42375,N_39557,N_38083);
nor U42376 (N_42376,N_38816,N_39586);
or U42377 (N_42377,N_39083,N_38562);
nor U42378 (N_42378,N_37676,N_39093);
nand U42379 (N_42379,N_39128,N_38140);
or U42380 (N_42380,N_39416,N_39213);
nor U42381 (N_42381,N_38842,N_38927);
or U42382 (N_42382,N_38727,N_37755);
and U42383 (N_42383,N_39549,N_38178);
xor U42384 (N_42384,N_39646,N_39817);
or U42385 (N_42385,N_38936,N_38588);
nor U42386 (N_42386,N_37507,N_38836);
nand U42387 (N_42387,N_37640,N_37692);
or U42388 (N_42388,N_39755,N_39708);
or U42389 (N_42389,N_37831,N_38071);
nor U42390 (N_42390,N_38074,N_38888);
and U42391 (N_42391,N_38988,N_38650);
and U42392 (N_42392,N_39636,N_39712);
xor U42393 (N_42393,N_38535,N_39149);
nand U42394 (N_42394,N_38795,N_38592);
xnor U42395 (N_42395,N_38204,N_38215);
or U42396 (N_42396,N_38702,N_39275);
or U42397 (N_42397,N_38328,N_38134);
xor U42398 (N_42398,N_39785,N_38293);
nor U42399 (N_42399,N_38136,N_39599);
or U42400 (N_42400,N_39255,N_38052);
xor U42401 (N_42401,N_37964,N_38769);
nand U42402 (N_42402,N_38113,N_38358);
nand U42403 (N_42403,N_38948,N_39898);
and U42404 (N_42404,N_39036,N_39394);
or U42405 (N_42405,N_39261,N_38902);
nand U42406 (N_42406,N_37641,N_39598);
or U42407 (N_42407,N_38002,N_38690);
or U42408 (N_42408,N_38035,N_37881);
or U42409 (N_42409,N_37742,N_38210);
xnor U42410 (N_42410,N_39210,N_37988);
nand U42411 (N_42411,N_37648,N_38623);
nand U42412 (N_42412,N_39766,N_38061);
nand U42413 (N_42413,N_37740,N_39923);
nor U42414 (N_42414,N_38273,N_38546);
xor U42415 (N_42415,N_39363,N_39128);
nand U42416 (N_42416,N_38441,N_39373);
nand U42417 (N_42417,N_38022,N_38928);
nor U42418 (N_42418,N_38205,N_39891);
and U42419 (N_42419,N_37918,N_39110);
nor U42420 (N_42420,N_39259,N_38128);
nand U42421 (N_42421,N_38441,N_37682);
and U42422 (N_42422,N_39413,N_37950);
nor U42423 (N_42423,N_37850,N_39809);
xor U42424 (N_42424,N_39447,N_39073);
nor U42425 (N_42425,N_39630,N_39878);
nand U42426 (N_42426,N_39285,N_39616);
and U42427 (N_42427,N_39507,N_39625);
nor U42428 (N_42428,N_37785,N_37930);
or U42429 (N_42429,N_38669,N_38798);
xor U42430 (N_42430,N_38791,N_37758);
or U42431 (N_42431,N_38542,N_38977);
and U42432 (N_42432,N_37801,N_37933);
or U42433 (N_42433,N_38938,N_39389);
nand U42434 (N_42434,N_37986,N_38412);
nor U42435 (N_42435,N_38269,N_39563);
or U42436 (N_42436,N_39668,N_37898);
and U42437 (N_42437,N_39575,N_38698);
nor U42438 (N_42438,N_38080,N_38872);
and U42439 (N_42439,N_38701,N_38888);
nor U42440 (N_42440,N_37649,N_39768);
nor U42441 (N_42441,N_38487,N_39407);
and U42442 (N_42442,N_37750,N_37885);
and U42443 (N_42443,N_38594,N_38487);
xor U42444 (N_42444,N_38699,N_38237);
nand U42445 (N_42445,N_39217,N_39948);
xor U42446 (N_42446,N_39761,N_39883);
xor U42447 (N_42447,N_38133,N_38543);
nor U42448 (N_42448,N_37968,N_39234);
or U42449 (N_42449,N_38549,N_39892);
and U42450 (N_42450,N_38518,N_38967);
nor U42451 (N_42451,N_38458,N_38082);
nor U42452 (N_42452,N_38693,N_39019);
and U42453 (N_42453,N_38942,N_38237);
or U42454 (N_42454,N_38155,N_38012);
nand U42455 (N_42455,N_38636,N_39958);
or U42456 (N_42456,N_37668,N_39942);
or U42457 (N_42457,N_38778,N_39831);
nor U42458 (N_42458,N_37679,N_39830);
or U42459 (N_42459,N_38444,N_39224);
and U42460 (N_42460,N_39128,N_37683);
nand U42461 (N_42461,N_38997,N_38055);
nand U42462 (N_42462,N_39600,N_39991);
and U42463 (N_42463,N_38824,N_38730);
nor U42464 (N_42464,N_39119,N_38146);
nor U42465 (N_42465,N_37988,N_38612);
xor U42466 (N_42466,N_37649,N_39879);
and U42467 (N_42467,N_38819,N_38855);
and U42468 (N_42468,N_38943,N_39218);
or U42469 (N_42469,N_38342,N_37791);
xor U42470 (N_42470,N_39422,N_37524);
or U42471 (N_42471,N_38896,N_39366);
nand U42472 (N_42472,N_37672,N_37946);
nand U42473 (N_42473,N_39544,N_38203);
or U42474 (N_42474,N_38552,N_38491);
nand U42475 (N_42475,N_38897,N_38069);
and U42476 (N_42476,N_38622,N_38662);
or U42477 (N_42477,N_38007,N_39191);
or U42478 (N_42478,N_38115,N_39500);
xor U42479 (N_42479,N_39554,N_38026);
xnor U42480 (N_42480,N_37744,N_38412);
or U42481 (N_42481,N_38479,N_38276);
and U42482 (N_42482,N_38281,N_38658);
nor U42483 (N_42483,N_37935,N_39963);
and U42484 (N_42484,N_39249,N_37986);
or U42485 (N_42485,N_38554,N_38638);
and U42486 (N_42486,N_39955,N_38575);
nor U42487 (N_42487,N_37737,N_38235);
nor U42488 (N_42488,N_38370,N_38712);
nor U42489 (N_42489,N_39375,N_37555);
and U42490 (N_42490,N_37984,N_39469);
or U42491 (N_42491,N_38772,N_37635);
and U42492 (N_42492,N_39167,N_38246);
nand U42493 (N_42493,N_37635,N_37850);
and U42494 (N_42494,N_37874,N_39710);
or U42495 (N_42495,N_39631,N_39157);
or U42496 (N_42496,N_39727,N_38411);
or U42497 (N_42497,N_39728,N_37843);
and U42498 (N_42498,N_37588,N_39679);
or U42499 (N_42499,N_39008,N_39634);
or U42500 (N_42500,N_41123,N_41674);
nand U42501 (N_42501,N_42283,N_40582);
xor U42502 (N_42502,N_40424,N_40905);
or U42503 (N_42503,N_40332,N_40246);
xor U42504 (N_42504,N_40363,N_40537);
xnor U42505 (N_42505,N_42093,N_41653);
nor U42506 (N_42506,N_40245,N_41370);
nor U42507 (N_42507,N_40543,N_40214);
nand U42508 (N_42508,N_42121,N_40063);
nor U42509 (N_42509,N_40681,N_41752);
and U42510 (N_42510,N_40888,N_42169);
or U42511 (N_42511,N_41871,N_40460);
nor U42512 (N_42512,N_42278,N_41881);
and U42513 (N_42513,N_41529,N_40461);
nor U42514 (N_42514,N_40873,N_41096);
and U42515 (N_42515,N_41775,N_41533);
or U42516 (N_42516,N_42461,N_41641);
and U42517 (N_42517,N_42444,N_41099);
and U42518 (N_42518,N_40694,N_41421);
and U42519 (N_42519,N_40539,N_41458);
nor U42520 (N_42520,N_41578,N_41877);
or U42521 (N_42521,N_40816,N_40528);
xor U42522 (N_42522,N_40978,N_41713);
and U42523 (N_42523,N_40630,N_40941);
nand U42524 (N_42524,N_41730,N_40493);
and U42525 (N_42525,N_40326,N_41728);
and U42526 (N_42526,N_42078,N_41587);
nor U42527 (N_42527,N_42231,N_40285);
xor U42528 (N_42528,N_40558,N_40810);
nand U42529 (N_42529,N_40282,N_40385);
nand U42530 (N_42530,N_40331,N_41467);
and U42531 (N_42531,N_40463,N_42383);
nor U42532 (N_42532,N_40125,N_41814);
and U42533 (N_42533,N_40456,N_40360);
and U42534 (N_42534,N_40447,N_42467);
nand U42535 (N_42535,N_42295,N_40945);
or U42536 (N_42536,N_41361,N_40754);
and U42537 (N_42537,N_41279,N_41299);
and U42538 (N_42538,N_41124,N_42447);
or U42539 (N_42539,N_40176,N_40114);
xnor U42540 (N_42540,N_42016,N_40614);
or U42541 (N_42541,N_41495,N_41816);
nand U42542 (N_42542,N_40751,N_40504);
and U42543 (N_42543,N_40172,N_42191);
and U42544 (N_42544,N_40159,N_40092);
and U42545 (N_42545,N_40773,N_41548);
or U42546 (N_42546,N_41913,N_42087);
nand U42547 (N_42547,N_42276,N_40429);
nor U42548 (N_42548,N_41621,N_42303);
nand U42549 (N_42549,N_40716,N_41072);
nand U42550 (N_42550,N_41874,N_40970);
xnor U42551 (N_42551,N_41318,N_41635);
or U42552 (N_42552,N_42466,N_41089);
nor U42553 (N_42553,N_42242,N_41900);
and U42554 (N_42554,N_41356,N_42199);
and U42555 (N_42555,N_41040,N_40604);
and U42556 (N_42556,N_42109,N_40319);
and U42557 (N_42557,N_42437,N_41032);
and U42558 (N_42558,N_41451,N_41748);
nor U42559 (N_42559,N_41504,N_40184);
nand U42560 (N_42560,N_40964,N_41494);
nor U42561 (N_42561,N_40309,N_40966);
or U42562 (N_42562,N_40141,N_41935);
xor U42563 (N_42563,N_41273,N_41563);
or U42564 (N_42564,N_42042,N_40281);
xor U42565 (N_42565,N_41159,N_41717);
nor U42566 (N_42566,N_42334,N_40173);
xor U42567 (N_42567,N_42309,N_41559);
nor U42568 (N_42568,N_40288,N_41114);
or U42569 (N_42569,N_41378,N_40106);
nand U42570 (N_42570,N_41425,N_41836);
xnor U42571 (N_42571,N_40554,N_41064);
and U42572 (N_42572,N_42223,N_42014);
xor U42573 (N_42573,N_40984,N_40157);
and U42574 (N_42574,N_41339,N_41917);
nor U42575 (N_42575,N_41245,N_41920);
or U42576 (N_42576,N_42054,N_41868);
nor U42577 (N_42577,N_40564,N_41510);
or U42578 (N_42578,N_41837,N_41979);
nor U42579 (N_42579,N_41586,N_42055);
and U42580 (N_42580,N_40737,N_41798);
and U42581 (N_42581,N_40919,N_41244);
nor U42582 (N_42582,N_40110,N_41945);
nor U42583 (N_42583,N_40771,N_40840);
and U42584 (N_42584,N_41139,N_41033);
nor U42585 (N_42585,N_40165,N_42480);
xnor U42586 (N_42586,N_40766,N_41895);
nor U42587 (N_42587,N_40629,N_42038);
or U42588 (N_42588,N_40039,N_40312);
or U42589 (N_42589,N_40739,N_41854);
and U42590 (N_42590,N_41324,N_40591);
xnor U42591 (N_42591,N_41531,N_42454);
nand U42592 (N_42592,N_42413,N_40512);
nor U42593 (N_42593,N_40408,N_42060);
xor U42594 (N_42594,N_41859,N_41046);
nand U42595 (N_42595,N_41289,N_41109);
and U42596 (N_42596,N_41851,N_41455);
nand U42597 (N_42597,N_41779,N_40889);
nor U42598 (N_42598,N_42187,N_41232);
and U42599 (N_42599,N_41841,N_42089);
or U42600 (N_42600,N_42498,N_41843);
and U42601 (N_42601,N_42373,N_41155);
or U42602 (N_42602,N_40803,N_41661);
xor U42603 (N_42603,N_40894,N_41119);
nand U42604 (N_42604,N_40896,N_42327);
or U42605 (N_42605,N_41902,N_41024);
and U42606 (N_42606,N_40683,N_42182);
and U42607 (N_42607,N_42420,N_40358);
or U42608 (N_42608,N_40191,N_40817);
and U42609 (N_42609,N_41600,N_42185);
nand U42610 (N_42610,N_40823,N_42439);
xor U42611 (N_42611,N_41879,N_41258);
nand U42612 (N_42612,N_41118,N_41625);
and U42613 (N_42613,N_40797,N_41508);
and U42614 (N_42614,N_42357,N_41190);
nor U42615 (N_42615,N_42022,N_40928);
nand U42616 (N_42616,N_40248,N_42219);
or U42617 (N_42617,N_41929,N_41822);
or U42618 (N_42618,N_40085,N_42393);
xnor U42619 (N_42619,N_41426,N_41380);
xor U42620 (N_42620,N_40433,N_41283);
xnor U42621 (N_42621,N_42266,N_42114);
nand U42622 (N_42622,N_41715,N_41084);
nor U42623 (N_42623,N_40301,N_41825);
nor U42624 (N_42624,N_41227,N_41857);
and U42625 (N_42625,N_41626,N_41000);
or U42626 (N_42626,N_40047,N_40858);
nand U42627 (N_42627,N_41523,N_40814);
or U42628 (N_42628,N_40428,N_42059);
nor U42629 (N_42629,N_42139,N_42064);
nand U42630 (N_42630,N_41400,N_41177);
or U42631 (N_42631,N_41321,N_42364);
xnor U42632 (N_42632,N_41937,N_40801);
and U42633 (N_42633,N_41699,N_41434);
nor U42634 (N_42634,N_41517,N_42485);
xor U42635 (N_42635,N_42049,N_41127);
nor U42636 (N_42636,N_41703,N_41628);
or U42637 (N_42637,N_41320,N_40013);
or U42638 (N_42638,N_42484,N_41027);
xor U42639 (N_42639,N_42183,N_40393);
nor U42640 (N_42640,N_42288,N_42062);
xor U42641 (N_42641,N_41242,N_41154);
and U42642 (N_42642,N_40208,N_42149);
xor U42643 (N_42643,N_41296,N_41212);
nor U42644 (N_42644,N_40418,N_40649);
nor U42645 (N_42645,N_40497,N_40035);
nor U42646 (N_42646,N_40343,N_40618);
nor U42647 (N_42647,N_40202,N_41169);
nor U42648 (N_42648,N_41844,N_40796);
or U42649 (N_42649,N_40811,N_42493);
and U42650 (N_42650,N_41813,N_40259);
nor U42651 (N_42651,N_40071,N_40325);
nand U42652 (N_42652,N_41444,N_41146);
and U42653 (N_42653,N_40425,N_41145);
and U42654 (N_42654,N_41860,N_40726);
nor U42655 (N_42655,N_41465,N_40160);
and U42656 (N_42656,N_40608,N_42116);
xor U42657 (N_42657,N_41041,N_40718);
nand U42658 (N_42658,N_40728,N_40451);
and U42659 (N_42659,N_40083,N_41233);
or U42660 (N_42660,N_40074,N_42048);
and U42661 (N_42661,N_41330,N_42353);
or U42662 (N_42662,N_42255,N_40401);
or U42663 (N_42663,N_40741,N_41838);
xnor U42664 (N_42664,N_40854,N_40107);
and U42665 (N_42665,N_42287,N_41654);
or U42666 (N_42666,N_42072,N_40606);
nor U42667 (N_42667,N_40507,N_40989);
and U42668 (N_42668,N_41098,N_41058);
nand U42669 (N_42669,N_40375,N_41256);
nor U42670 (N_42670,N_41484,N_40471);
xnor U42671 (N_42671,N_40122,N_40480);
xnor U42672 (N_42672,N_41776,N_40836);
and U42673 (N_42673,N_40943,N_42172);
nor U42674 (N_42674,N_41669,N_41107);
and U42675 (N_42675,N_41565,N_40475);
xor U42676 (N_42676,N_42227,N_41409);
or U42677 (N_42677,N_41360,N_41391);
xor U42678 (N_42678,N_41012,N_41452);
or U42679 (N_42679,N_40581,N_41202);
xnor U42680 (N_42680,N_41521,N_40339);
and U42681 (N_42681,N_40825,N_40464);
and U42682 (N_42682,N_41062,N_41846);
or U42683 (N_42683,N_41090,N_41315);
or U42684 (N_42684,N_41785,N_40559);
nand U42685 (N_42685,N_41938,N_41608);
or U42686 (N_42686,N_40243,N_40225);
xnor U42687 (N_42687,N_41787,N_41973);
nand U42688 (N_42688,N_40844,N_42312);
and U42689 (N_42689,N_42339,N_40257);
nand U42690 (N_42690,N_42319,N_42264);
xnor U42691 (N_42691,N_40570,N_42488);
or U42692 (N_42692,N_40598,N_41778);
nor U42693 (N_42693,N_40027,N_41926);
and U42694 (N_42694,N_41863,N_41542);
nor U42695 (N_42695,N_41166,N_40620);
or U42696 (N_42696,N_42145,N_41821);
or U42697 (N_42697,N_41094,N_40364);
nor U42698 (N_42698,N_40426,N_41055);
xor U42699 (N_42699,N_41566,N_41848);
or U42700 (N_42700,N_40177,N_41709);
nand U42701 (N_42701,N_40183,N_40891);
nor U42702 (N_42702,N_40546,N_40699);
and U42703 (N_42703,N_40111,N_41589);
xnor U42704 (N_42704,N_40879,N_40166);
xor U42705 (N_42705,N_40832,N_41053);
nand U42706 (N_42706,N_42051,N_42425);
xnor U42707 (N_42707,N_41039,N_41942);
nor U42708 (N_42708,N_41708,N_41035);
nor U42709 (N_42709,N_40899,N_40254);
nand U42710 (N_42710,N_41304,N_40065);
or U42711 (N_42711,N_41671,N_42030);
xnor U42712 (N_42712,N_40109,N_42019);
nor U42713 (N_42713,N_41718,N_41535);
and U42714 (N_42714,N_40732,N_41250);
nand U42715 (N_42715,N_41948,N_41052);
nor U42716 (N_42716,N_41178,N_41684);
nor U42717 (N_42717,N_42052,N_40575);
or U42718 (N_42718,N_41372,N_42232);
and U42719 (N_42719,N_41137,N_40032);
and U42720 (N_42720,N_42245,N_42193);
nand U42721 (N_42721,N_42099,N_42027);
xor U42722 (N_42722,N_41382,N_42321);
nor U42723 (N_42723,N_42256,N_42167);
xnor U42724 (N_42724,N_41911,N_41316);
and U42725 (N_42725,N_40959,N_41716);
or U42726 (N_42726,N_40508,N_41476);
xnor U42727 (N_42727,N_40410,N_40453);
or U42728 (N_42728,N_41422,N_40596);
nand U42729 (N_42729,N_41644,N_40200);
nor U42730 (N_42730,N_41440,N_40361);
nor U42731 (N_42731,N_42147,N_41679);
and U42732 (N_42732,N_40302,N_42065);
nor U42733 (N_42733,N_41348,N_41922);
nand U42734 (N_42734,N_40234,N_41077);
nand U42735 (N_42735,N_42229,N_40968);
xnor U42736 (N_42736,N_41101,N_42270);
nor U42737 (N_42737,N_40824,N_41855);
nor U42738 (N_42738,N_42369,N_41925);
xor U42739 (N_42739,N_40226,N_41095);
or U42740 (N_42740,N_42472,N_41369);
and U42741 (N_42741,N_41683,N_41038);
nor U42742 (N_42742,N_41007,N_40684);
xor U42743 (N_42743,N_42214,N_42403);
nor U42744 (N_42744,N_40270,N_42047);
xor U42745 (N_42745,N_40344,N_41737);
nor U42746 (N_42746,N_41078,N_42128);
nand U42747 (N_42747,N_41598,N_41261);
and U42748 (N_42748,N_40218,N_41065);
and U42749 (N_42749,N_40932,N_42363);
and U42750 (N_42750,N_40272,N_40357);
or U42751 (N_42751,N_41694,N_41964);
nand U42752 (N_42752,N_42127,N_40164);
or U42753 (N_42753,N_42098,N_41350);
nor U42754 (N_42754,N_40223,N_41477);
and U42755 (N_42755,N_41710,N_40756);
and U42756 (N_42756,N_41128,N_40204);
nor U42757 (N_42757,N_40096,N_41284);
or U42758 (N_42758,N_41489,N_40443);
nand U42759 (N_42759,N_41750,N_40403);
or U42760 (N_42760,N_40067,N_41918);
xor U42761 (N_42761,N_40755,N_40887);
xnor U42762 (N_42762,N_41497,N_41329);
xnor U42763 (N_42763,N_42448,N_42143);
nand U42764 (N_42764,N_41796,N_41777);
xnor U42765 (N_42765,N_41930,N_41005);
and U42766 (N_42766,N_41097,N_41376);
or U42767 (N_42767,N_40567,N_40793);
nor U42768 (N_42768,N_41470,N_42310);
nand U42769 (N_42769,N_40579,N_41905);
or U42770 (N_42770,N_41211,N_42251);
nand U42771 (N_42771,N_41664,N_41558);
xnor U42772 (N_42772,N_40278,N_42379);
xor U42773 (N_42773,N_41503,N_40522);
nand U42774 (N_42774,N_42160,N_42152);
xor U42775 (N_42775,N_42213,N_41173);
and U42776 (N_42776,N_40830,N_42120);
and U42777 (N_42777,N_40438,N_40822);
and U42778 (N_42778,N_40616,N_42424);
nor U42779 (N_42779,N_40053,N_42071);
nand U42780 (N_42780,N_40648,N_40264);
nand U42781 (N_42781,N_42279,N_41165);
nand U42782 (N_42782,N_41524,N_40473);
xnor U42783 (N_42783,N_42090,N_41666);
xnor U42784 (N_42784,N_41959,N_41840);
nand U42785 (N_42785,N_42208,N_41619);
xnor U42786 (N_42786,N_40483,N_42240);
nor U42787 (N_42787,N_40631,N_40008);
nor U42788 (N_42788,N_42415,N_40249);
and U42789 (N_42789,N_42431,N_41347);
and U42790 (N_42790,N_41552,N_40229);
and U42791 (N_42791,N_40232,N_41665);
nand U42792 (N_42792,N_40623,N_40486);
xnor U42793 (N_42793,N_41714,N_40267);
nand U42794 (N_42794,N_41014,N_40593);
nor U42795 (N_42795,N_42377,N_40153);
xor U42796 (N_42796,N_41519,N_40667);
xor U42797 (N_42797,N_40777,N_40014);
nand U42798 (N_42798,N_41474,N_41682);
or U42799 (N_42799,N_40380,N_40055);
nor U42800 (N_42800,N_42076,N_41952);
or U42801 (N_42801,N_42165,N_42181);
nand U42802 (N_42802,N_40911,N_40127);
and U42803 (N_42803,N_41867,N_42384);
nor U42804 (N_42804,N_42487,N_40406);
nor U42805 (N_42805,N_42380,N_42492);
nor U42806 (N_42806,N_42083,N_42180);
nand U42807 (N_42807,N_41130,N_40637);
nand U42808 (N_42808,N_40626,N_40409);
xnor U42809 (N_42809,N_41463,N_42402);
and U42810 (N_42810,N_40452,N_40506);
or U42811 (N_42811,N_40691,N_41026);
nand U42812 (N_42812,N_42331,N_41656);
and U42813 (N_42813,N_42088,N_42164);
nor U42814 (N_42814,N_40304,N_41511);
xor U42815 (N_42815,N_40359,N_41646);
or U42816 (N_42816,N_40072,N_42226);
and U42817 (N_42817,N_41736,N_42138);
nor U42818 (N_42818,N_41645,N_40277);
nor U42819 (N_42819,N_40383,N_40875);
nand U42820 (N_42820,N_40330,N_40790);
nand U42821 (N_42821,N_41006,N_41357);
nand U42822 (N_42822,N_41488,N_40569);
and U42823 (N_42823,N_40449,N_41575);
nand U42824 (N_42824,N_42391,N_40155);
nor U42825 (N_42825,N_41527,N_42299);
or U42826 (N_42826,N_41622,N_40839);
xor U42827 (N_42827,N_41904,N_42296);
or U42828 (N_42828,N_42095,N_40088);
and U42829 (N_42829,N_40525,N_40396);
and U42830 (N_42830,N_41428,N_40747);
nor U42831 (N_42831,N_40856,N_42176);
or U42832 (N_42832,N_40075,N_42246);
nand U42833 (N_42833,N_40702,N_41176);
and U42834 (N_42834,N_41997,N_40435);
or U42835 (N_42835,N_41305,N_40617);
nand U42836 (N_42836,N_40759,N_41201);
xor U42837 (N_42837,N_41291,N_40763);
and U42838 (N_42838,N_41649,N_40199);
and U42839 (N_42839,N_40073,N_41195);
nor U42840 (N_42840,N_40413,N_41398);
or U42841 (N_42841,N_40016,N_41856);
and U42842 (N_42842,N_40472,N_41104);
and U42843 (N_42843,N_42489,N_41249);
or U42844 (N_42844,N_41416,N_40952);
xor U42845 (N_42845,N_40397,N_41267);
or U42846 (N_42846,N_42024,N_41804);
nand U42847 (N_42847,N_40962,N_41269);
xnor U42848 (N_42848,N_40542,N_41358);
or U42849 (N_42849,N_41810,N_41915);
xor U42850 (N_42850,N_42222,N_41274);
nand U42851 (N_42851,N_41082,N_41023);
and U42852 (N_42852,N_41429,N_40284);
nand U42853 (N_42853,N_41262,N_41652);
nand U42854 (N_42854,N_42221,N_40927);
or U42855 (N_42855,N_40263,N_41206);
nor U42856 (N_42856,N_40156,N_40185);
and U42857 (N_42857,N_40697,N_42247);
and U42858 (N_42858,N_40686,N_41762);
nor U42859 (N_42859,N_41725,N_40026);
nor U42860 (N_42860,N_40576,N_41158);
nand U42861 (N_42861,N_41323,N_41138);
nand U42862 (N_42862,N_40171,N_41751);
nand U42863 (N_42863,N_40010,N_41362);
xnor U42864 (N_42864,N_41368,N_40897);
nor U42865 (N_42865,N_40354,N_40336);
or U42866 (N_42866,N_40914,N_40130);
nand U42867 (N_42867,N_42112,N_42486);
or U42868 (N_42868,N_41120,N_41886);
or U42869 (N_42869,N_41912,N_40863);
or U42870 (N_42870,N_41883,N_40216);
nor U42871 (N_42871,N_42441,N_41592);
and U42872 (N_42872,N_40224,N_40124);
xor U42873 (N_42873,N_40242,N_42274);
or U42874 (N_42874,N_41793,N_40024);
nand U42875 (N_42875,N_40398,N_41819);
nor U42876 (N_42876,N_41236,N_42244);
and U42877 (N_42877,N_41208,N_40174);
nand U42878 (N_42878,N_40807,N_41235);
and U42879 (N_42879,N_40213,N_40091);
and U42880 (N_42880,N_41835,N_42053);
and U42881 (N_42881,N_41093,N_40640);
and U42882 (N_42882,N_41591,N_40033);
nor U42883 (N_42883,N_41438,N_40087);
and U42884 (N_42884,N_40484,N_41932);
xnor U42885 (N_42885,N_40862,N_40561);
and U42886 (N_42886,N_41733,N_41204);
and U42887 (N_42887,N_41260,N_41583);
nor U42888 (N_42888,N_41083,N_42471);
nand U42889 (N_42889,N_40972,N_41353);
nand U42890 (N_42890,N_41086,N_40289);
or U42891 (N_42891,N_41971,N_40338);
nand U42892 (N_42892,N_40253,N_40780);
xnor U42893 (N_42893,N_41462,N_42355);
or U42894 (N_42894,N_42032,N_40168);
nand U42895 (N_42895,N_40538,N_40735);
nand U42896 (N_42896,N_40740,N_42204);
xor U42897 (N_42897,N_40712,N_40210);
xnor U42898 (N_42898,N_40280,N_40916);
or U42899 (N_42899,N_41282,N_41771);
xnor U42900 (N_42900,N_41188,N_41799);
nand U42901 (N_42901,N_41486,N_42146);
and U42902 (N_42902,N_40139,N_40520);
and U42903 (N_42903,N_40511,N_42455);
and U42904 (N_42904,N_41543,N_40900);
nor U42905 (N_42905,N_41346,N_41601);
or U42906 (N_42906,N_41693,N_41336);
nand U42907 (N_42907,N_40909,N_40745);
nor U42908 (N_42908,N_41056,N_41593);
nor U42909 (N_42909,N_41695,N_41116);
and U42910 (N_42910,N_41496,N_41588);
nor U42911 (N_42911,N_40679,N_41167);
and U42912 (N_42912,N_41958,N_40209);
xor U42913 (N_42913,N_41092,N_42034);
nor U42914 (N_42914,N_40791,N_40379);
and U42915 (N_42915,N_40995,N_41248);
nand U42916 (N_42916,N_42201,N_40706);
or U42917 (N_42917,N_42217,N_41757);
nand U42918 (N_42918,N_40673,N_42236);
or U42919 (N_42919,N_40201,N_40835);
and U42920 (N_42920,N_41240,N_40300);
or U42921 (N_42921,N_41896,N_42328);
xnor U42922 (N_42922,N_42170,N_41744);
nor U42923 (N_42923,N_41220,N_40761);
or U42924 (N_42924,N_41512,N_40847);
and U42925 (N_42925,N_41224,N_40827);
nand U42926 (N_42926,N_41374,N_40513);
nor U42927 (N_42927,N_40306,N_41383);
nand U42928 (N_42928,N_41557,N_40350);
or U42929 (N_42929,N_40536,N_42066);
or U42930 (N_42930,N_40400,N_42365);
xnor U42931 (N_42931,N_41332,N_42297);
and U42932 (N_42932,N_41605,N_40235);
nand U42933 (N_42933,N_41272,N_42130);
and U42934 (N_42934,N_41739,N_42011);
nand U42935 (N_42935,N_40316,N_40434);
or U42936 (N_42936,N_42496,N_41824);
and U42937 (N_42937,N_42440,N_42341);
or U42938 (N_42938,N_40977,N_40685);
or U42939 (N_42939,N_41327,N_42238);
and U42940 (N_42940,N_40432,N_41156);
nand U42941 (N_42941,N_42207,N_41492);
nor U42942 (N_42942,N_41532,N_40238);
nand U42943 (N_42943,N_41987,N_41670);
nor U42944 (N_42944,N_41658,N_42458);
and U42945 (N_42945,N_41050,N_42330);
nand U42946 (N_42946,N_42451,N_41899);
nand U42947 (N_42947,N_42122,N_40329);
nor U42948 (N_42948,N_42432,N_41160);
nor U42949 (N_42949,N_40126,N_40644);
nor U42950 (N_42950,N_40314,N_41680);
nand U42951 (N_42951,N_40178,N_41916);
or U42952 (N_42952,N_40129,N_40152);
xor U42953 (N_42953,N_41355,N_40069);
nand U42954 (N_42954,N_40872,N_42253);
and U42955 (N_42955,N_42366,N_41264);
xnor U42956 (N_42956,N_41268,N_40866);
and U42957 (N_42957,N_41554,N_42301);
xnor U42958 (N_42958,N_41044,N_41157);
xor U42959 (N_42959,N_42332,N_40700);
and U42960 (N_42960,N_41872,N_40005);
nor U42961 (N_42961,N_40381,N_40588);
nand U42962 (N_42962,N_41759,N_41317);
or U42963 (N_42963,N_41756,N_40369);
nand U42964 (N_42964,N_40104,N_40923);
nand U42965 (N_42965,N_40275,N_40386);
xnor U42966 (N_42966,N_40946,N_40081);
and U42967 (N_42967,N_40999,N_40247);
nor U42968 (N_42968,N_41610,N_41878);
or U42969 (N_42969,N_42061,N_41547);
nor U42970 (N_42970,N_40056,N_40222);
xor U42971 (N_42971,N_41216,N_41414);
or U42972 (N_42972,N_41833,N_40310);
and U42973 (N_42973,N_42449,N_42004);
or U42974 (N_42974,N_42017,N_40994);
or U42975 (N_42975,N_40274,N_41121);
nand U42976 (N_42976,N_41795,N_40098);
and U42977 (N_42977,N_41638,N_40136);
and U42978 (N_42978,N_42411,N_40529);
and U42979 (N_42979,N_42422,N_41627);
xnor U42980 (N_42980,N_41140,N_40041);
or U42981 (N_42981,N_41515,N_40327);
nor U42982 (N_42982,N_41403,N_40391);
xnor U42983 (N_42983,N_41681,N_40286);
or U42984 (N_42984,N_40594,N_41633);
nand U42985 (N_42985,N_40592,N_41830);
and U42986 (N_42986,N_40474,N_42329);
and U42987 (N_42987,N_40351,N_40421);
or U42988 (N_42988,N_40342,N_40965);
xor U42989 (N_42989,N_41424,N_40599);
xor U42990 (N_42990,N_40782,N_41657);
nor U42991 (N_42991,N_41069,N_42342);
and U42992 (N_42992,N_41051,N_40636);
nand U42993 (N_42993,N_42478,N_41433);
nor U42994 (N_42994,N_41105,N_41970);
xnor U42995 (N_42995,N_40799,N_41031);
nand U42996 (N_42996,N_42442,N_41483);
nand U42997 (N_42997,N_41528,N_41004);
nor U42998 (N_42998,N_41300,N_41161);
and U42999 (N_42999,N_40059,N_41667);
and U43000 (N_43000,N_40298,N_42389);
xnor U43001 (N_43001,N_40635,N_40920);
and U43002 (N_43002,N_40979,N_40258);
and U43003 (N_43003,N_42346,N_40672);
nor U43004 (N_43004,N_41615,N_40244);
nand U43005 (N_43005,N_40105,N_42300);
nand U43006 (N_43006,N_40240,N_40004);
and U43007 (N_43007,N_40347,N_40487);
nor U43008 (N_43008,N_41991,N_40052);
or U43009 (N_43009,N_42345,N_41115);
nand U43010 (N_43010,N_41676,N_40785);
xnor U43011 (N_43011,N_41271,N_41436);
and U43012 (N_43012,N_42473,N_40647);
and U43013 (N_43013,N_41561,N_40731);
nand U43014 (N_43014,N_41662,N_41191);
nand U43015 (N_43015,N_40662,N_40677);
or U43016 (N_43016,N_42446,N_42243);
nor U43017 (N_43017,N_41581,N_41947);
nor U43018 (N_43018,N_41839,N_40519);
and U43019 (N_43019,N_40813,N_40885);
xor U43020 (N_43020,N_42323,N_41394);
and U43021 (N_43021,N_41919,N_41473);
xnor U43022 (N_43022,N_42018,N_42317);
nor U43023 (N_43023,N_41013,N_40880);
and U43024 (N_43024,N_42436,N_40402);
xnor U43025 (N_43025,N_42494,N_40044);
and U43026 (N_43026,N_40193,N_40730);
and U43027 (N_43027,N_41509,N_40633);
and U43028 (N_43028,N_40874,N_41789);
nor U43029 (N_43029,N_40861,N_41067);
and U43030 (N_43030,N_40211,N_41659);
and U43031 (N_43031,N_41199,N_40265);
or U43032 (N_43032,N_41534,N_41168);
xnor U43033 (N_43033,N_41122,N_41387);
xor U43034 (N_43034,N_40057,N_40076);
nor U43035 (N_43035,N_42307,N_41914);
xnor U43036 (N_43036,N_42406,N_42400);
and U43037 (N_43037,N_42189,N_40646);
xor U43038 (N_43038,N_41826,N_40061);
nand U43039 (N_43039,N_41502,N_40212);
nor U43040 (N_43040,N_42387,N_41147);
xnor U43041 (N_43041,N_41927,N_40145);
nor U43042 (N_43042,N_40976,N_42198);
nand U43043 (N_43043,N_40757,N_42316);
nand U43044 (N_43044,N_40585,N_41349);
xnor U43045 (N_43045,N_41786,N_41745);
and U43046 (N_43046,N_40195,N_41999);
and U43047 (N_43047,N_40333,N_41892);
and U43048 (N_43048,N_41590,N_40855);
xnor U43049 (N_43049,N_40427,N_40668);
xor U43050 (N_43050,N_40315,N_41344);
nand U43051 (N_43051,N_40659,N_41481);
nand U43052 (N_43052,N_40196,N_42007);
xnor U43053 (N_43053,N_41729,N_41549);
nand U43054 (N_43054,N_41246,N_41325);
xnor U43055 (N_43055,N_41228,N_40786);
xnor U43056 (N_43056,N_42465,N_40940);
nor U43057 (N_43057,N_41998,N_41407);
nand U43058 (N_43058,N_40846,N_40382);
nor U43059 (N_43059,N_41252,N_41686);
nand U43060 (N_43060,N_40675,N_41110);
and U43061 (N_43061,N_41364,N_40587);
nor U43062 (N_43062,N_41435,N_40415);
xnor U43063 (N_43063,N_42118,N_41969);
and U43064 (N_43064,N_41614,N_42315);
or U43065 (N_43065,N_40121,N_40030);
nand U43066 (N_43066,N_40025,N_41408);
nand U43067 (N_43067,N_41449,N_41701);
and U43068 (N_43068,N_41331,N_41573);
or U43069 (N_43069,N_41726,N_40666);
and U43070 (N_43070,N_40837,N_41102);
or U43071 (N_43071,N_41263,N_41849);
nand U43072 (N_43072,N_40925,N_40828);
nor U43073 (N_43073,N_41112,N_41982);
nor U43074 (N_43074,N_41420,N_41042);
nand U43075 (N_43075,N_41990,N_42368);
and U43076 (N_43076,N_40148,N_40643);
and U43077 (N_43077,N_42335,N_40356);
or U43078 (N_43078,N_40902,N_41545);
nor U43079 (N_43079,N_41980,N_40607);
nand U43080 (N_43080,N_41672,N_41864);
nand U43081 (N_43081,N_41399,N_41150);
nand U43082 (N_43082,N_40046,N_40038);
nor U43083 (N_43083,N_41774,N_40910);
or U43084 (N_43084,N_40501,N_41311);
or U43085 (N_43085,N_41749,N_41957);
and U43086 (N_43086,N_42009,N_41392);
nor U43087 (N_43087,N_41266,N_40957);
xnor U43088 (N_43088,N_42237,N_41108);
xnor U43089 (N_43089,N_42302,N_40938);
nand U43090 (N_43090,N_40578,N_40707);
xnor U43091 (N_43091,N_41479,N_41412);
xor U43092 (N_43092,N_41063,N_40366);
or U43093 (N_43093,N_40708,N_42044);
or U43094 (N_43094,N_42468,N_41210);
nand U43095 (N_43095,N_41555,N_41020);
nor U43096 (N_43096,N_40573,N_41319);
and U43097 (N_43097,N_40290,N_42381);
xor U43098 (N_43098,N_40491,N_41976);
and U43099 (N_43099,N_41572,N_40003);
xnor U43100 (N_43100,N_40857,N_41769);
nor U43101 (N_43101,N_42233,N_40348);
nor U43102 (N_43102,N_40086,N_40414);
xnor U43103 (N_43103,N_40181,N_41427);
or U43104 (N_43104,N_40792,N_40661);
and U43105 (N_43105,N_40568,N_40743);
nand U43106 (N_43106,N_41933,N_41943);
or U43107 (N_43107,N_41490,N_41576);
nor U43108 (N_43108,N_40665,N_40973);
and U43109 (N_43109,N_40192,N_41359);
and U43110 (N_43110,N_40605,N_40251);
and U43111 (N_43111,N_40169,N_41743);
and U43112 (N_43112,N_42041,N_40521);
and U43113 (N_43113,N_41522,N_41500);
xor U43114 (N_43114,N_40996,N_40906);
or U43115 (N_43115,N_40012,N_41363);
and U43116 (N_43116,N_40527,N_40749);
nor U43117 (N_43117,N_41237,N_41673);
or U43118 (N_43118,N_41003,N_41487);
nor U43119 (N_43119,N_41560,N_41338);
or U43120 (N_43120,N_42161,N_42291);
nor U43121 (N_43121,N_40942,N_40859);
or U43122 (N_43122,N_41540,N_41450);
or U43123 (N_43123,N_42386,N_41910);
nand U43124 (N_43124,N_42350,N_40458);
xor U43125 (N_43125,N_41472,N_41617);
and U43126 (N_43126,N_42006,N_40313);
and U43127 (N_43127,N_40307,N_40006);
nand U43128 (N_43128,N_40346,N_40419);
nor U43129 (N_43129,N_40645,N_42397);
nor U43130 (N_43130,N_42070,N_41594);
nand U43131 (N_43131,N_41788,N_41008);
xnor U43132 (N_43132,N_41755,N_40935);
or U43133 (N_43133,N_42028,N_42125);
and U43134 (N_43134,N_42271,N_40465);
nand U43135 (N_43135,N_41406,N_42037);
and U43136 (N_43136,N_41596,N_40054);
and U43137 (N_43137,N_41314,N_40710);
xnor U43138 (N_43138,N_41845,N_40405);
nand U43139 (N_43139,N_41043,N_42086);
or U43140 (N_43140,N_41194,N_40496);
and U43141 (N_43141,N_41965,N_41829);
or U43142 (N_43142,N_40353,N_42096);
or U43143 (N_43143,N_40266,N_40577);
xnor U43144 (N_43144,N_41047,N_42094);
or U43145 (N_43145,N_40744,N_40028);
and U43146 (N_43146,N_41939,N_40101);
or U43147 (N_43147,N_40116,N_42285);
xor U43148 (N_43148,N_41075,N_41828);
xnor U43149 (N_43149,N_40058,N_41782);
or U43150 (N_43150,N_41341,N_41908);
nand U43151 (N_43151,N_42102,N_41852);
or U43152 (N_43152,N_40279,N_41126);
xnor U43153 (N_43153,N_41797,N_40231);
nand U43154 (N_43154,N_41187,N_40963);
xnor U43155 (N_43155,N_41525,N_40108);
nor U43156 (N_43156,N_41758,N_40709);
xor U43157 (N_43157,N_41197,N_42354);
nor U43158 (N_43158,N_40851,N_40628);
nand U43159 (N_43159,N_41071,N_41536);
and U43160 (N_43160,N_41171,N_40770);
nand U43161 (N_43161,N_41270,N_42258);
nor U43162 (N_43162,N_40221,N_41891);
nand U43163 (N_43163,N_40748,N_41802);
nand U43164 (N_43164,N_42367,N_42029);
nand U43165 (N_43165,N_41921,N_40283);
or U43166 (N_43166,N_40634,N_41518);
nor U43167 (N_43167,N_40510,N_41876);
or U43168 (N_43168,N_40954,N_41516);
nor U43169 (N_43169,N_40600,N_41901);
nand U43170 (N_43170,N_40753,N_40560);
nor U43171 (N_43171,N_42033,N_40143);
nand U43172 (N_43172,N_41636,N_42103);
nand U43173 (N_43173,N_42067,N_41898);
xor U43174 (N_43174,N_40034,N_40769);
or U43175 (N_43175,N_40239,N_41688);
xnor U43176 (N_43176,N_42259,N_41309);
xor U43177 (N_43177,N_41151,N_41574);
xnor U43178 (N_43178,N_41229,N_40454);
xor U43179 (N_43179,N_40514,N_40215);
or U43180 (N_43180,N_40574,N_40660);
and U43181 (N_43181,N_41081,N_40650);
nor U43182 (N_43182,N_40768,N_41162);
or U43183 (N_43183,N_42340,N_41257);
nor U43184 (N_43184,N_40924,N_41866);
and U43185 (N_43185,N_41460,N_41491);
or U43186 (N_43186,N_41754,N_42252);
xor U43187 (N_43187,N_42490,N_40377);
or U43188 (N_43188,N_40602,N_41815);
nor U43189 (N_43189,N_41618,N_40981);
xor U43190 (N_43190,N_41553,N_41584);
and U43191 (N_43191,N_41609,N_40831);
and U43192 (N_43192,N_41506,N_40137);
nor U43193 (N_43193,N_41893,N_41307);
and U43194 (N_43194,N_41247,N_40865);
or U43195 (N_43195,N_40256,N_40079);
or U43196 (N_43196,N_41597,N_41367);
or U43197 (N_43197,N_41457,N_42284);
and U43198 (N_43198,N_42031,N_42421);
nor U43199 (N_43199,N_41800,N_40042);
nand U43200 (N_43200,N_41214,N_40120);
xnor U43201 (N_43201,N_41882,N_41738);
nand U43202 (N_43202,N_41390,N_41526);
or U43203 (N_43203,N_40490,N_40890);
xor U43204 (N_43204,N_41741,N_42001);
nor U43205 (N_43205,N_41996,N_41066);
nor U43206 (N_43206,N_40262,N_40701);
nand U43207 (N_43207,N_40982,N_41085);
xnor U43208 (N_43208,N_40291,N_42435);
xnor U43209 (N_43209,N_40980,N_41953);
xor U43210 (N_43210,N_41189,N_42101);
xnor U43211 (N_43211,N_42158,N_42476);
or U43212 (N_43212,N_40448,N_42280);
nand U43213 (N_43213,N_40161,N_40680);
nor U43214 (N_43214,N_40705,N_42050);
nand U43215 (N_43215,N_40808,N_40656);
and U43216 (N_43216,N_41808,N_42378);
xor U43217 (N_43217,N_41983,N_40719);
nor U43218 (N_43218,N_40671,N_40115);
nor U43219 (N_43219,N_41731,N_40062);
nor U43220 (N_43220,N_40131,N_41687);
nor U43221 (N_43221,N_41773,N_41087);
and U43222 (N_43222,N_41021,N_42450);
or U43223 (N_43223,N_41960,N_41478);
or U43224 (N_43224,N_41612,N_40615);
or U43225 (N_43225,N_42129,N_42123);
and U43226 (N_43226,N_41538,N_41221);
or U43227 (N_43227,N_41595,N_41764);
xnor U43228 (N_43228,N_40595,N_40717);
and U43229 (N_43229,N_40918,N_40812);
nor U43230 (N_43230,N_40020,N_42000);
xor U43231 (N_43231,N_41303,N_40788);
nor U43232 (N_43232,N_40392,N_41706);
or U43233 (N_43233,N_41962,N_41972);
or U43234 (N_43234,N_41234,N_41501);
nor U43235 (N_43235,N_42282,N_41278);
or U43236 (N_43236,N_41446,N_41869);
or U43237 (N_43237,N_41780,N_40276);
or U43238 (N_43238,N_40001,N_40252);
nand U43239 (N_43239,N_41034,N_41445);
nor U43240 (N_43240,N_42460,N_41397);
and U43241 (N_43241,N_40913,N_41599);
nor U43242 (N_43242,N_42399,N_40470);
nand U43243 (N_43243,N_41513,N_40746);
nand U43244 (N_43244,N_40303,N_40819);
nor U43245 (N_43245,N_40436,N_41766);
nand U43246 (N_43246,N_41880,N_41135);
and U43247 (N_43247,N_40881,N_42230);
nand U43248 (N_43248,N_40688,N_40557);
nand U43249 (N_43249,N_41482,N_42073);
xnor U43250 (N_43250,N_40084,N_40118);
nor U43251 (N_43251,N_41809,N_40586);
nand U43252 (N_43252,N_41281,N_40269);
nor U43253 (N_43253,N_42275,N_42443);
and U43254 (N_43254,N_42156,N_42002);
or U43255 (N_43255,N_41616,N_40841);
and U43256 (N_43256,N_40154,N_40829);
and U43257 (N_43257,N_41724,N_40362);
nor U43258 (N_43258,N_41923,N_41459);
xor U43259 (N_43259,N_41909,N_40795);
or U43260 (N_43260,N_42108,N_41411);
nor U43261 (N_43261,N_42388,N_41277);
nor U43262 (N_43262,N_40388,N_41298);
xor U43263 (N_43263,N_41772,N_42200);
nand U43264 (N_43264,N_41678,N_41286);
and U43265 (N_43265,N_40815,N_40230);
xnor U43266 (N_43266,N_40917,N_42483);
or U43267 (N_43267,N_40022,N_40517);
nor U43268 (N_43268,N_40187,N_41373);
or U43269 (N_43269,N_40676,N_40860);
nor U43270 (N_43270,N_40117,N_42314);
nand U43271 (N_43271,N_40322,N_42190);
nor U43272 (N_43272,N_40190,N_41310);
nor U43273 (N_43273,N_40467,N_42133);
or U43274 (N_43274,N_40450,N_40412);
nor U43275 (N_43275,N_42404,N_42209);
nor U43276 (N_43276,N_41696,N_42464);
xor U43277 (N_43277,N_40198,N_40934);
xnor U43278 (N_43278,N_42405,N_41520);
xor U43279 (N_43279,N_40713,N_41009);
or U43280 (N_43280,N_40162,N_41550);
nor U43281 (N_43281,N_42141,N_42410);
nand U43282 (N_43282,N_40149,N_40352);
or U43283 (N_43283,N_42412,N_42254);
or U43284 (N_43284,N_42263,N_42045);
and U43285 (N_43285,N_40476,N_41253);
and U43286 (N_43286,N_40371,N_41181);
or U43287 (N_43287,N_41530,N_40534);
and U43288 (N_43288,N_41213,N_42469);
nor U43289 (N_43289,N_40535,N_40430);
and U43290 (N_43290,N_40948,N_40031);
nor U43291 (N_43291,N_41760,N_41265);
nand U43292 (N_43292,N_42218,N_40724);
and U43293 (N_43293,N_42104,N_40509);
and U43294 (N_43294,N_42394,N_41389);
nor U43295 (N_43295,N_42457,N_42092);
and U43296 (N_43296,N_40674,N_42281);
nor U43297 (N_43297,N_42322,N_41820);
and U43298 (N_43298,N_40268,N_41230);
or U43299 (N_43299,N_41418,N_42268);
or U43300 (N_43300,N_41215,N_40992);
xor U43301 (N_43301,N_41606,N_40261);
or U43302 (N_43302,N_41639,N_40103);
nor U43303 (N_43303,N_41430,N_42115);
or U43304 (N_43304,N_42290,N_41136);
nand U43305 (N_43305,N_40203,N_40090);
nand U43306 (N_43306,N_40372,N_42126);
or U43307 (N_43307,N_40128,N_40915);
xnor U43308 (N_43308,N_40624,N_40734);
and U43309 (N_43309,N_40655,N_41651);
nand U43310 (N_43310,N_41702,N_40205);
nor U43311 (N_43311,N_40341,N_40933);
nor U43312 (N_43312,N_42456,N_40112);
or U43313 (N_43313,N_41238,N_40877);
nor U43314 (N_43314,N_40985,N_41727);
xor U43315 (N_43315,N_41017,N_41806);
nor U43316 (N_43316,N_41906,N_42482);
or U43317 (N_43317,N_41951,N_40113);
or U43318 (N_43318,N_42241,N_41057);
and U43319 (N_43319,N_42385,N_42091);
and U43320 (N_43320,N_41203,N_42151);
and U43321 (N_43321,N_40144,N_40818);
nor U43322 (N_43322,N_42056,N_41001);
or U43323 (N_43323,N_41631,N_40255);
nor U43324 (N_43324,N_40625,N_42398);
nor U43325 (N_43325,N_40787,N_41328);
or U43326 (N_43326,N_40019,N_42186);
xor U43327 (N_43327,N_40953,N_41448);
and U43328 (N_43328,N_41405,N_42491);
and U43329 (N_43329,N_41995,N_41163);
xor U43330 (N_43330,N_40197,N_42111);
and U43331 (N_43331,N_41541,N_40869);
nand U43332 (N_43332,N_41946,N_41170);
nand U43333 (N_43333,N_42058,N_41453);
or U43334 (N_43334,N_41393,N_40956);
and U43335 (N_43335,N_42148,N_42359);
nor U43336 (N_43336,N_40018,N_40455);
xor U43337 (N_43337,N_40219,N_40871);
or U43338 (N_43338,N_40930,N_40834);
and U43339 (N_43339,N_40439,N_41241);
xor U43340 (N_43340,N_40077,N_42477);
xor U43341 (N_43341,N_40775,N_40884);
xor U43342 (N_43342,N_42239,N_40097);
nor U43343 (N_43343,N_40533,N_42039);
xnor U43344 (N_43344,N_41698,N_42257);
or U43345 (N_43345,N_40563,N_40498);
or U43346 (N_43346,N_40642,N_41054);
nand U43347 (N_43347,N_41288,N_42344);
or U43348 (N_43348,N_42175,N_40373);
and U43349 (N_43349,N_41753,N_41768);
nand U43350 (N_43350,N_40798,N_41184);
and U43351 (N_43351,N_42433,N_40597);
nand U43352 (N_43352,N_41292,N_42154);
nor U43353 (N_43353,N_41700,N_40524);
xor U43354 (N_43354,N_41847,N_41604);
or U43355 (N_43355,N_40947,N_41335);
xnor U43356 (N_43356,N_41931,N_41507);
xnor U43357 (N_43357,N_41375,N_40423);
nor U43358 (N_43358,N_40868,N_41961);
nor U43359 (N_43359,N_41388,N_41569);
nand U43360 (N_43360,N_41432,N_40967);
or U43361 (N_43361,N_42106,N_41734);
and U43362 (N_43362,N_40715,N_42216);
nor U43363 (N_43363,N_40903,N_40936);
and U43364 (N_43364,N_40789,N_41015);
and U43365 (N_43365,N_41968,N_41805);
and U43366 (N_43366,N_42015,N_42084);
xor U43367 (N_43367,N_41924,N_40912);
nand U43368 (N_43368,N_41469,N_40068);
or U43369 (N_43369,N_40809,N_40664);
nor U43370 (N_43370,N_42304,N_41722);
and U43371 (N_43371,N_41306,N_41765);
and U43372 (N_43372,N_40800,N_42409);
nand U43373 (N_43373,N_40340,N_40904);
nand U43374 (N_43374,N_40997,N_42046);
nand U43375 (N_43375,N_40961,N_40011);
nor U43376 (N_43376,N_40589,N_41129);
and U43377 (N_43377,N_41275,N_41402);
nor U43378 (N_43378,N_40390,N_40457);
or U43379 (N_43379,N_41967,N_40750);
and U43380 (N_43380,N_41290,N_41989);
nand U43381 (N_43381,N_42075,N_41345);
or U43382 (N_43382,N_40337,N_41301);
or U43383 (N_43383,N_40742,N_42206);
nor U43384 (N_43384,N_41179,N_41539);
nor U43385 (N_43385,N_41611,N_42375);
or U43386 (N_43386,N_40552,N_42459);
nand U43387 (N_43387,N_40958,N_40207);
nor U43388 (N_43388,N_41144,N_41812);
and U43389 (N_43389,N_41384,N_42438);
xnor U43390 (N_43390,N_42035,N_40553);
nor U43391 (N_43391,N_42261,N_40163);
nor U43392 (N_43392,N_41148,N_41624);
nand U43393 (N_43393,N_40036,N_41419);
nor U43394 (N_43394,N_40652,N_40545);
and U43395 (N_43395,N_41551,N_42308);
or U43396 (N_43396,N_41562,N_40532);
nand U43397 (N_43397,N_40722,N_40931);
nand U43398 (N_43398,N_40293,N_40431);
nand U43399 (N_43399,N_42429,N_42430);
or U43400 (N_43400,N_40612,N_40653);
and U43401 (N_43401,N_40774,N_41888);
xor U43402 (N_43402,N_42192,N_41705);
and U43403 (N_43403,N_41480,N_40541);
xnor U43404 (N_43404,N_40395,N_40898);
xnor U43405 (N_43405,N_40601,N_41048);
or U43406 (N_43406,N_41763,N_42396);
and U43407 (N_43407,N_41732,N_40622);
nor U43408 (N_43408,N_42351,N_42277);
nand U43409 (N_43409,N_41784,N_42177);
nand U43410 (N_43410,N_41862,N_40138);
nand U43411 (N_43411,N_41985,N_40260);
xnor U43412 (N_43412,N_41196,N_40002);
nor U43413 (N_43413,N_40690,N_40882);
nor U43414 (N_43414,N_40937,N_40974);
nand U43415 (N_43415,N_41354,N_40370);
or U43416 (N_43416,N_41343,N_40170);
nor U43417 (N_43417,N_41742,N_40477);
and U43418 (N_43418,N_40853,N_40764);
or U43419 (N_43419,N_40023,N_41984);
and U43420 (N_43420,N_42153,N_42020);
or U43421 (N_43421,N_40733,N_40804);
and U43422 (N_43422,N_42497,N_41475);
and U43423 (N_43423,N_41125,N_40015);
or U43424 (N_43424,N_41132,N_42352);
nand U43425 (N_43425,N_40220,N_40609);
or U43426 (N_43426,N_40848,N_40583);
and U43427 (N_43427,N_40048,N_41875);
nor U43428 (N_43428,N_40488,N_41333);
xor U43429 (N_43429,N_41295,N_42068);
nand U43430 (N_43430,N_41537,N_42358);
nand U43431 (N_43431,N_40772,N_40689);
nor U43432 (N_43432,N_41907,N_41655);
nand U43433 (N_43433,N_41239,N_40000);
nand U43434 (N_43434,N_40499,N_40040);
xnor U43435 (N_43435,N_40893,N_40029);
nor U43436 (N_43436,N_41111,N_40540);
or U43437 (N_43437,N_42294,N_42372);
nand U43438 (N_43438,N_41746,N_42361);
or U43439 (N_43439,N_40794,N_42318);
xor U43440 (N_43440,N_41936,N_41294);
or U43441 (N_43441,N_41218,N_41832);
nand U43442 (N_43442,N_40349,N_41823);
xor U43443 (N_43443,N_42100,N_42224);
nand U43444 (N_43444,N_41297,N_41807);
nand U43445 (N_43445,N_41966,N_41255);
nor U43446 (N_43446,N_41704,N_40548);
or U43447 (N_43447,N_40551,N_40721);
and U43448 (N_43448,N_40526,N_42134);
nand U43449 (N_43449,N_40147,N_40781);
and U43450 (N_43450,N_40627,N_42196);
nand U43451 (N_43451,N_41711,N_41884);
and U43452 (N_43452,N_40939,N_42474);
nor U43453 (N_43453,N_42043,N_41192);
and U43454 (N_43454,N_41865,N_41801);
and U43455 (N_43455,N_40621,N_40611);
xor U43456 (N_43456,N_41842,N_40845);
xnor U43457 (N_43457,N_42113,N_42097);
nor U43458 (N_43458,N_41415,N_40696);
nor U43459 (N_43459,N_41934,N_42371);
nor U43460 (N_43460,N_40901,N_41029);
nor U43461 (N_43461,N_41834,N_41954);
nor U43462 (N_43462,N_40151,N_40670);
and U43463 (N_43463,N_40878,N_40523);
nand U43464 (N_43464,N_41049,N_42136);
or U43465 (N_43465,N_40292,N_40440);
nand U43466 (N_43466,N_40489,N_40404);
nor U43467 (N_43467,N_40287,N_41060);
nand U43468 (N_43468,N_42427,N_40368);
xnor U43469 (N_43469,N_41141,N_41308);
nand U43470 (N_43470,N_40478,N_40132);
nor U43471 (N_43471,N_41461,N_40955);
xor U43472 (N_43472,N_42159,N_42401);
xor U43473 (N_43473,N_40021,N_41721);
and U43474 (N_43474,N_42144,N_40987);
or U43475 (N_43475,N_40641,N_40321);
nor U43476 (N_43476,N_42077,N_41499);
and U43477 (N_43477,N_40378,N_40736);
and U43478 (N_43478,N_42225,N_41259);
and U43479 (N_43479,N_40250,N_41174);
nor U43480 (N_43480,N_41091,N_40094);
and U43481 (N_43481,N_40565,N_40562);
xnor U43482 (N_43482,N_40571,N_42445);
nand U43483 (N_43483,N_40544,N_40444);
and U43484 (N_43484,N_42036,N_40446);
nor U43485 (N_43485,N_41439,N_41185);
nor U43486 (N_43486,N_41885,N_40045);
or U43487 (N_43487,N_40693,N_41342);
nand U43488 (N_43488,N_41442,N_42179);
xnor U43489 (N_43489,N_40870,N_41226);
xnor U43490 (N_43490,N_41992,N_40466);
nand U43491 (N_43491,N_41607,N_40070);
nor U43492 (N_43492,N_40502,N_41723);
nor U43493 (N_43493,N_40294,N_40064);
and U43494 (N_43494,N_41117,N_41994);
or U43495 (N_43495,N_42184,N_42292);
or U43496 (N_43496,N_40323,N_40037);
xor U43497 (N_43497,N_40308,N_41571);
and U43498 (N_43498,N_41334,N_42390);
or U43499 (N_43499,N_42140,N_41735);
or U43500 (N_43500,N_40678,N_41395);
nor U43501 (N_43501,N_41685,N_42021);
xor U43502 (N_43502,N_40271,N_41149);
and U43503 (N_43503,N_40459,N_41811);
and U43504 (N_43504,N_40806,N_40311);
nor U43505 (N_43505,N_41988,N_40367);
nand U43506 (N_43506,N_40335,N_40765);
or U43507 (N_43507,N_41103,N_42462);
xnor U43508 (N_43508,N_41831,N_41164);
and U43509 (N_43509,N_40556,N_41193);
or U43510 (N_43510,N_40133,N_42215);
nand U43511 (N_43511,N_41689,N_40669);
nand U43512 (N_43512,N_40971,N_40420);
nor U43513 (N_43513,N_41632,N_42205);
and U43514 (N_43514,N_41142,N_40990);
xor U43515 (N_43515,N_40566,N_40711);
or U43516 (N_43516,N_41544,N_40066);
or U43517 (N_43517,N_42135,N_41385);
xor U43518 (N_43518,N_40993,N_40485);
and U43519 (N_43519,N_42171,N_40907);
nand U43520 (N_43520,N_40227,N_41712);
nor U43521 (N_43521,N_40206,N_40555);
nand U43522 (N_43522,N_41890,N_41949);
nand U43523 (N_43523,N_42005,N_41505);
nor U43524 (N_43524,N_41514,N_42010);
xor U43525 (N_43525,N_40194,N_40758);
and U43526 (N_43526,N_42311,N_41697);
nor U43527 (N_43527,N_40345,N_41903);
nor U43528 (N_43528,N_40394,N_41817);
and U43529 (N_43529,N_42426,N_40500);
xnor U43530 (N_43530,N_40549,N_40407);
xor U43531 (N_43531,N_40462,N_41352);
or U43532 (N_43532,N_40049,N_41016);
or U43533 (N_43533,N_41648,N_41761);
or U43534 (N_43534,N_42026,N_41861);
nand U43535 (N_43535,N_40704,N_40007);
and U43536 (N_43536,N_40228,N_41396);
or U43537 (N_43537,N_40852,N_42040);
xnor U43538 (N_43538,N_41577,N_40998);
nand U43539 (N_43539,N_40417,N_40784);
nand U43540 (N_43540,N_41570,N_42262);
nor U43541 (N_43541,N_42142,N_41580);
nor U43542 (N_43542,N_41404,N_42418);
and U43543 (N_43543,N_41276,N_40723);
xnor U43544 (N_43544,N_40838,N_42417);
nand U43545 (N_43545,N_42376,N_41205);
nand U43546 (N_43546,N_41993,N_40687);
xnor U43547 (N_43547,N_40580,N_42349);
nor U43548 (N_43548,N_40017,N_40820);
nand U43549 (N_43549,N_40080,N_41381);
or U43550 (N_43550,N_42298,N_40515);
nor U43551 (N_43551,N_40482,N_41113);
or U43552 (N_43552,N_42265,N_42362);
xnor U43553 (N_43553,N_42269,N_40297);
or U43554 (N_43554,N_42481,N_41377);
nor U43555 (N_43555,N_41302,N_41794);
or U43556 (N_43556,N_42343,N_40099);
nand U43557 (N_43557,N_41243,N_40779);
nor U43558 (N_43558,N_40590,N_40422);
and U43559 (N_43559,N_41133,N_41207);
nor U43560 (N_43560,N_40776,N_40365);
or U43561 (N_43561,N_40043,N_41172);
nor U43562 (N_43562,N_40503,N_42150);
xnor U43563 (N_43563,N_41131,N_41219);
nor U43564 (N_43564,N_41963,N_41579);
nand U43565 (N_43565,N_40355,N_42212);
nor U43566 (N_43566,N_42434,N_41827);
xnor U43567 (N_43567,N_40188,N_40089);
and U43568 (N_43568,N_41351,N_40638);
xor U43569 (N_43569,N_41074,N_41944);
nor U43570 (N_43570,N_40682,N_41950);
or U43571 (N_43571,N_40833,N_42419);
or U43572 (N_43572,N_42211,N_42414);
xor U43573 (N_43573,N_42013,N_42124);
or U43574 (N_43574,N_41200,N_41251);
nor U43575 (N_43575,N_41740,N_41894);
xor U43576 (N_43576,N_40180,N_41582);
xnor U43577 (N_43577,N_41792,N_40657);
and U43578 (N_43578,N_41401,N_41642);
nor U43579 (N_43579,N_40142,N_42475);
nand U43580 (N_43580,N_42423,N_41546);
and U43581 (N_43581,N_40100,N_41853);
nor U43582 (N_43582,N_41285,N_42107);
nand U43583 (N_43583,N_40495,N_40140);
nor U43584 (N_43584,N_42117,N_42132);
xnor U43585 (N_43585,N_41366,N_42110);
nor U43586 (N_43586,N_41019,N_40986);
nand U43587 (N_43587,N_40135,N_40060);
nor U43588 (N_43588,N_40387,N_41978);
and U43589 (N_43589,N_40505,N_42012);
xor U43590 (N_43590,N_40720,N_41977);
xnor U43591 (N_43591,N_42069,N_40328);
nor U43592 (N_43592,N_41152,N_41322);
nor U43593 (N_43593,N_42347,N_41603);
xnor U43594 (N_43594,N_42338,N_41143);
nand U43595 (N_43595,N_40481,N_41326);
xnor U43596 (N_43596,N_40236,N_42210);
xnor U43597 (N_43597,N_41783,N_41002);
and U43598 (N_43598,N_40572,N_41280);
nor U43599 (N_43599,N_41423,N_42293);
nor U43600 (N_43600,N_41940,N_41818);
nand U43601 (N_43601,N_40411,N_40698);
nor U43602 (N_43602,N_42320,N_40805);
xnor U43603 (N_43603,N_40783,N_41209);
xnor U43604 (N_43604,N_40658,N_41312);
nor U43605 (N_43605,N_40802,N_40095);
or U43606 (N_43606,N_40217,N_42360);
xor U43607 (N_43607,N_41720,N_40437);
xnor U43608 (N_43608,N_40078,N_41630);
xnor U43609 (N_43609,N_40729,N_40603);
nand U43610 (N_43610,N_40692,N_42495);
and U43611 (N_43611,N_41018,N_41620);
or U43612 (N_43612,N_42063,N_42228);
nand U43613 (N_43613,N_41153,N_41955);
and U43614 (N_43614,N_41677,N_42194);
or U43615 (N_43615,N_41287,N_41956);
nand U43616 (N_43616,N_41365,N_41431);
xor U43617 (N_43617,N_40695,N_40102);
xnor U43618 (N_43618,N_42248,N_42289);
or U43619 (N_43619,N_40445,N_42131);
xnor U43620 (N_43620,N_42336,N_40727);
xor U43621 (N_43621,N_42166,N_41293);
nand U43622 (N_43622,N_41371,N_40241);
or U43623 (N_43623,N_41634,N_42470);
xnor U43624 (N_43624,N_41928,N_40969);
nand U43625 (N_43625,N_41088,N_42155);
and U43626 (N_43626,N_42428,N_40051);
nand U43627 (N_43627,N_40237,N_42057);
and U43628 (N_43628,N_40123,N_41025);
or U43629 (N_43629,N_40399,N_41623);
xor U43630 (N_43630,N_40843,N_40584);
nand U43631 (N_43631,N_40950,N_42324);
xor U43632 (N_43632,N_41254,N_40550);
or U43633 (N_43633,N_41707,N_41803);
nand U43634 (N_43634,N_41337,N_40175);
nor U43635 (N_43635,N_42080,N_42081);
nor U43636 (N_43636,N_41182,N_40416);
nor U43637 (N_43637,N_42326,N_40082);
and U43638 (N_43638,N_41059,N_41747);
nand U43639 (N_43639,N_40760,N_40610);
xnor U43640 (N_43640,N_40295,N_42025);
nand U43641 (N_43641,N_40849,N_41556);
xor U43642 (N_43642,N_40469,N_41850);
and U43643 (N_43643,N_41471,N_42085);
nand U43644 (N_43644,N_40960,N_41975);
or U43645 (N_43645,N_41217,N_41313);
nor U43646 (N_43646,N_42325,N_40389);
or U43647 (N_43647,N_42305,N_40922);
nand U43648 (N_43648,N_41079,N_41791);
or U43649 (N_43649,N_40895,N_40703);
or U43650 (N_43650,N_41070,N_42079);
nand U43651 (N_43651,N_42074,N_40093);
or U43652 (N_43652,N_40179,N_40944);
nand U43653 (N_43653,N_40883,N_40778);
or U43654 (N_43654,N_42203,N_42260);
nand U43655 (N_43655,N_42374,N_40299);
xor U43656 (N_43656,N_40663,N_41602);
nor U43657 (N_43657,N_41568,N_40442);
or U43658 (N_43658,N_41887,N_41456);
and U43659 (N_43659,N_42188,N_40479);
nor U43660 (N_43660,N_40134,N_42453);
nor U43661 (N_43661,N_40494,N_40119);
nand U43662 (N_43662,N_40050,N_42499);
and U43663 (N_43663,N_41030,N_40850);
nor U43664 (N_43664,N_42082,N_42286);
nor U43665 (N_43665,N_42337,N_40725);
nor U43666 (N_43666,N_42348,N_41498);
nor U43667 (N_43667,N_41231,N_41870);
and U43668 (N_43668,N_41466,N_41441);
or U43669 (N_43669,N_40921,N_41889);
or U43670 (N_43670,N_40767,N_42234);
nor U43671 (N_43671,N_40492,N_42273);
nor U43672 (N_43672,N_41981,N_41037);
and U43673 (N_43673,N_40632,N_42119);
xor U43674 (N_43674,N_40983,N_42105);
nor U43675 (N_43675,N_42202,N_40334);
xor U43676 (N_43676,N_41340,N_40384);
nand U43677 (N_43677,N_42463,N_40233);
and U43678 (N_43678,N_40892,N_40146);
xnor U43679 (N_43679,N_42162,N_42382);
xor U43680 (N_43680,N_41660,N_40613);
xnor U43681 (N_43681,N_40273,N_40518);
and U43682 (N_43682,N_40908,N_41379);
and U43683 (N_43683,N_41028,N_41010);
or U43684 (N_43684,N_40189,N_40752);
nand U43685 (N_43685,N_42197,N_40929);
or U43686 (N_43686,N_40186,N_41647);
xnor U43687 (N_43687,N_41100,N_42220);
nor U43688 (N_43688,N_42173,N_42408);
xnor U43689 (N_43689,N_41454,N_40324);
nand U43690 (N_43690,N_42416,N_42370);
nand U43691 (N_43691,N_40158,N_40876);
or U43692 (N_43692,N_41585,N_41036);
nor U43693 (N_43693,N_40009,N_40468);
and U43694 (N_43694,N_40150,N_42168);
and U43695 (N_43695,N_40441,N_42157);
nand U43696 (N_43696,N_41106,N_41437);
nor U43697 (N_43697,N_41663,N_41629);
nand U43698 (N_43698,N_41767,N_41134);
nor U43699 (N_43699,N_41781,N_41464);
xnor U43700 (N_43700,N_42137,N_42008);
and U43701 (N_43701,N_41225,N_41417);
nor U43702 (N_43702,N_41080,N_41613);
xnor U43703 (N_43703,N_40951,N_42195);
nand U43704 (N_43704,N_40821,N_40318);
and U43705 (N_43705,N_42249,N_40738);
nand U43706 (N_43706,N_40639,N_40374);
and U43707 (N_43707,N_41974,N_41386);
xor U43708 (N_43708,N_41447,N_41468);
xor U43709 (N_43709,N_42272,N_41643);
xor U43710 (N_43710,N_41011,N_40826);
and U43711 (N_43711,N_40317,N_42407);
xor U43712 (N_43712,N_42392,N_42174);
or U43713 (N_43713,N_41068,N_42178);
and U43714 (N_43714,N_40714,N_41413);
or U43715 (N_43715,N_41986,N_42306);
nand U43716 (N_43716,N_40867,N_42023);
xor U43717 (N_43717,N_40531,N_41443);
and U43718 (N_43718,N_40762,N_40975);
xnor U43719 (N_43719,N_42163,N_41873);
nor U43720 (N_43720,N_41222,N_40320);
nor U43721 (N_43721,N_40886,N_41790);
or U43722 (N_43722,N_41198,N_42356);
nor U43723 (N_43723,N_41076,N_41223);
nor U43724 (N_43724,N_41897,N_40926);
xor U43725 (N_43725,N_41175,N_40305);
nand U43726 (N_43726,N_42479,N_40182);
xor U43727 (N_43727,N_42235,N_41690);
and U43728 (N_43728,N_41073,N_41640);
nand U43729 (N_43729,N_41045,N_42267);
nand U43730 (N_43730,N_40864,N_40654);
nor U43731 (N_43731,N_41941,N_40167);
and U43732 (N_43732,N_41719,N_40988);
nand U43733 (N_43733,N_41567,N_42313);
nand U43734 (N_43734,N_41485,N_40619);
nor U43735 (N_43735,N_41186,N_40530);
nand U43736 (N_43736,N_41564,N_41691);
nand U43737 (N_43737,N_40842,N_41061);
xnor U43738 (N_43738,N_42333,N_41668);
xor U43739 (N_43739,N_42250,N_42003);
and U43740 (N_43740,N_41493,N_41637);
and U43741 (N_43741,N_40991,N_41675);
or U43742 (N_43742,N_41858,N_41410);
nand U43743 (N_43743,N_40376,N_42452);
or U43744 (N_43744,N_40651,N_41650);
nor U43745 (N_43745,N_41770,N_42395);
or U43746 (N_43746,N_41022,N_40949);
nor U43747 (N_43747,N_41180,N_40547);
nand U43748 (N_43748,N_41692,N_40296);
or U43749 (N_43749,N_40516,N_41183);
nor U43750 (N_43750,N_42316,N_40156);
xnor U43751 (N_43751,N_42228,N_42128);
or U43752 (N_43752,N_41828,N_41819);
nor U43753 (N_43753,N_40814,N_42459);
and U43754 (N_43754,N_40749,N_40846);
or U43755 (N_43755,N_40593,N_41987);
xor U43756 (N_43756,N_40261,N_42170);
and U43757 (N_43757,N_40425,N_40486);
or U43758 (N_43758,N_40156,N_40793);
xor U43759 (N_43759,N_42470,N_40946);
xnor U43760 (N_43760,N_41045,N_42087);
and U43761 (N_43761,N_42270,N_40919);
nand U43762 (N_43762,N_40540,N_40703);
xnor U43763 (N_43763,N_40338,N_41264);
nor U43764 (N_43764,N_41607,N_40326);
or U43765 (N_43765,N_40956,N_40451);
xor U43766 (N_43766,N_40997,N_41350);
and U43767 (N_43767,N_41270,N_41957);
xnor U43768 (N_43768,N_41163,N_42357);
and U43769 (N_43769,N_40057,N_40226);
and U43770 (N_43770,N_42101,N_42225);
xor U43771 (N_43771,N_41026,N_41178);
or U43772 (N_43772,N_40742,N_41454);
nand U43773 (N_43773,N_41323,N_42214);
xnor U43774 (N_43774,N_40023,N_41628);
and U43775 (N_43775,N_41445,N_42112);
xnor U43776 (N_43776,N_41672,N_41255);
and U43777 (N_43777,N_42164,N_40810);
nor U43778 (N_43778,N_41437,N_40292);
and U43779 (N_43779,N_40846,N_41071);
nor U43780 (N_43780,N_40149,N_40439);
nand U43781 (N_43781,N_40767,N_42463);
nor U43782 (N_43782,N_40388,N_41309);
and U43783 (N_43783,N_40524,N_41240);
nor U43784 (N_43784,N_40183,N_41260);
nand U43785 (N_43785,N_42399,N_42329);
nand U43786 (N_43786,N_42460,N_42436);
nor U43787 (N_43787,N_42489,N_41001);
nand U43788 (N_43788,N_41501,N_41499);
nor U43789 (N_43789,N_41498,N_40687);
xor U43790 (N_43790,N_40165,N_40769);
nor U43791 (N_43791,N_40851,N_40859);
and U43792 (N_43792,N_41127,N_41253);
nand U43793 (N_43793,N_41969,N_41084);
and U43794 (N_43794,N_42301,N_41331);
and U43795 (N_43795,N_40199,N_42421);
nand U43796 (N_43796,N_41457,N_40077);
xnor U43797 (N_43797,N_41903,N_42412);
xor U43798 (N_43798,N_40665,N_41315);
xnor U43799 (N_43799,N_41955,N_41903);
nand U43800 (N_43800,N_40732,N_40907);
nand U43801 (N_43801,N_42399,N_41651);
nor U43802 (N_43802,N_41508,N_41105);
nand U43803 (N_43803,N_41277,N_40801);
nor U43804 (N_43804,N_42021,N_40540);
xnor U43805 (N_43805,N_41423,N_41712);
xor U43806 (N_43806,N_41247,N_41317);
xnor U43807 (N_43807,N_40835,N_40627);
or U43808 (N_43808,N_42160,N_40177);
or U43809 (N_43809,N_40452,N_40746);
nand U43810 (N_43810,N_40301,N_40551);
and U43811 (N_43811,N_40505,N_41195);
nand U43812 (N_43812,N_40587,N_40096);
xnor U43813 (N_43813,N_42045,N_42115);
nand U43814 (N_43814,N_40887,N_42278);
nand U43815 (N_43815,N_41829,N_42348);
or U43816 (N_43816,N_41655,N_40706);
nor U43817 (N_43817,N_42373,N_40101);
nand U43818 (N_43818,N_40412,N_40049);
and U43819 (N_43819,N_41516,N_40056);
or U43820 (N_43820,N_41151,N_40083);
nand U43821 (N_43821,N_40894,N_40567);
or U43822 (N_43822,N_42472,N_42077);
nor U43823 (N_43823,N_40454,N_40251);
and U43824 (N_43824,N_42404,N_42315);
and U43825 (N_43825,N_41828,N_41156);
xor U43826 (N_43826,N_41217,N_42085);
nor U43827 (N_43827,N_41886,N_41576);
xnor U43828 (N_43828,N_40375,N_40608);
xnor U43829 (N_43829,N_41598,N_40515);
nor U43830 (N_43830,N_40578,N_42484);
xnor U43831 (N_43831,N_40031,N_40083);
nand U43832 (N_43832,N_40335,N_42437);
or U43833 (N_43833,N_40282,N_41607);
and U43834 (N_43834,N_40636,N_42088);
nor U43835 (N_43835,N_42412,N_41405);
nand U43836 (N_43836,N_40344,N_41714);
and U43837 (N_43837,N_42494,N_42053);
and U43838 (N_43838,N_40410,N_42491);
or U43839 (N_43839,N_40788,N_40151);
nand U43840 (N_43840,N_42234,N_42094);
or U43841 (N_43841,N_41932,N_41901);
nor U43842 (N_43842,N_42371,N_41129);
xnor U43843 (N_43843,N_41646,N_41150);
nor U43844 (N_43844,N_40807,N_40156);
xor U43845 (N_43845,N_42494,N_42329);
nand U43846 (N_43846,N_41051,N_40047);
nand U43847 (N_43847,N_40110,N_40797);
and U43848 (N_43848,N_40118,N_40417);
xnor U43849 (N_43849,N_42460,N_40554);
nand U43850 (N_43850,N_41755,N_42000);
nor U43851 (N_43851,N_40716,N_40960);
or U43852 (N_43852,N_41146,N_42229);
nor U43853 (N_43853,N_40512,N_40908);
or U43854 (N_43854,N_40735,N_41399);
xor U43855 (N_43855,N_41745,N_40395);
nor U43856 (N_43856,N_41037,N_41027);
and U43857 (N_43857,N_40124,N_40954);
nand U43858 (N_43858,N_40090,N_41425);
nor U43859 (N_43859,N_40289,N_42376);
nor U43860 (N_43860,N_41103,N_41916);
or U43861 (N_43861,N_40614,N_40850);
xor U43862 (N_43862,N_42167,N_42354);
and U43863 (N_43863,N_41833,N_40250);
or U43864 (N_43864,N_40694,N_40254);
nor U43865 (N_43865,N_41690,N_40456);
xor U43866 (N_43866,N_40700,N_41022);
xor U43867 (N_43867,N_41669,N_41545);
or U43868 (N_43868,N_41130,N_42078);
or U43869 (N_43869,N_40830,N_41260);
nor U43870 (N_43870,N_40685,N_41818);
nor U43871 (N_43871,N_42392,N_41760);
or U43872 (N_43872,N_40750,N_40842);
nand U43873 (N_43873,N_40278,N_40523);
xor U43874 (N_43874,N_40384,N_40599);
or U43875 (N_43875,N_42054,N_40573);
xnor U43876 (N_43876,N_42304,N_41280);
nand U43877 (N_43877,N_40865,N_41908);
nor U43878 (N_43878,N_41778,N_41808);
nor U43879 (N_43879,N_42255,N_42415);
and U43880 (N_43880,N_42213,N_41093);
and U43881 (N_43881,N_41150,N_42363);
nor U43882 (N_43882,N_40619,N_40023);
nand U43883 (N_43883,N_42243,N_42437);
or U43884 (N_43884,N_42484,N_41963);
nand U43885 (N_43885,N_42021,N_40972);
and U43886 (N_43886,N_42290,N_42318);
or U43887 (N_43887,N_41371,N_42397);
xor U43888 (N_43888,N_42012,N_42163);
and U43889 (N_43889,N_40102,N_41109);
xor U43890 (N_43890,N_42282,N_41363);
xor U43891 (N_43891,N_41184,N_41719);
nor U43892 (N_43892,N_40243,N_41712);
nor U43893 (N_43893,N_41851,N_42284);
xor U43894 (N_43894,N_41636,N_41409);
xor U43895 (N_43895,N_40766,N_40242);
xor U43896 (N_43896,N_42052,N_41556);
or U43897 (N_43897,N_41097,N_40925);
nor U43898 (N_43898,N_40540,N_41078);
nor U43899 (N_43899,N_40484,N_40663);
nor U43900 (N_43900,N_41429,N_40782);
xor U43901 (N_43901,N_40852,N_41047);
and U43902 (N_43902,N_40544,N_42442);
xnor U43903 (N_43903,N_41476,N_42095);
or U43904 (N_43904,N_41523,N_42170);
nor U43905 (N_43905,N_41684,N_41349);
or U43906 (N_43906,N_40088,N_41331);
nor U43907 (N_43907,N_40223,N_40664);
or U43908 (N_43908,N_41329,N_41528);
and U43909 (N_43909,N_41715,N_41196);
and U43910 (N_43910,N_41009,N_41836);
nand U43911 (N_43911,N_42393,N_40121);
and U43912 (N_43912,N_42391,N_41180);
xor U43913 (N_43913,N_42016,N_41647);
or U43914 (N_43914,N_41961,N_41845);
nor U43915 (N_43915,N_41152,N_40144);
xnor U43916 (N_43916,N_40296,N_41734);
xnor U43917 (N_43917,N_40504,N_41067);
and U43918 (N_43918,N_41817,N_40587);
and U43919 (N_43919,N_41236,N_40390);
nand U43920 (N_43920,N_42004,N_40547);
or U43921 (N_43921,N_40392,N_40924);
nand U43922 (N_43922,N_41672,N_41248);
and U43923 (N_43923,N_40470,N_41098);
nor U43924 (N_43924,N_40172,N_40130);
and U43925 (N_43925,N_40321,N_40491);
nor U43926 (N_43926,N_41962,N_41493);
nor U43927 (N_43927,N_40423,N_42133);
nand U43928 (N_43928,N_41039,N_41703);
nand U43929 (N_43929,N_41613,N_41610);
or U43930 (N_43930,N_40243,N_42207);
nor U43931 (N_43931,N_42053,N_41703);
and U43932 (N_43932,N_40304,N_41850);
or U43933 (N_43933,N_40549,N_42383);
and U43934 (N_43934,N_40465,N_42304);
nand U43935 (N_43935,N_41498,N_40800);
nor U43936 (N_43936,N_40191,N_42168);
nand U43937 (N_43937,N_41292,N_41595);
nand U43938 (N_43938,N_40107,N_42408);
and U43939 (N_43939,N_40584,N_40917);
and U43940 (N_43940,N_41763,N_42229);
nor U43941 (N_43941,N_41151,N_42116);
nor U43942 (N_43942,N_41364,N_41014);
nand U43943 (N_43943,N_41044,N_40958);
xnor U43944 (N_43944,N_41668,N_40326);
nor U43945 (N_43945,N_40276,N_40439);
or U43946 (N_43946,N_40487,N_41059);
xor U43947 (N_43947,N_40716,N_41116);
nand U43948 (N_43948,N_41848,N_40856);
nor U43949 (N_43949,N_41168,N_42370);
xnor U43950 (N_43950,N_40480,N_40420);
or U43951 (N_43951,N_40312,N_40390);
nand U43952 (N_43952,N_40862,N_40764);
or U43953 (N_43953,N_40601,N_42496);
nand U43954 (N_43954,N_40937,N_40065);
nor U43955 (N_43955,N_40132,N_41312);
nand U43956 (N_43956,N_41825,N_42087);
or U43957 (N_43957,N_40023,N_40966);
xor U43958 (N_43958,N_42426,N_41552);
and U43959 (N_43959,N_42223,N_42376);
and U43960 (N_43960,N_41967,N_40496);
nand U43961 (N_43961,N_42067,N_41433);
xor U43962 (N_43962,N_40561,N_40774);
xnor U43963 (N_43963,N_42042,N_40245);
xor U43964 (N_43964,N_42033,N_42225);
or U43965 (N_43965,N_40963,N_40264);
nand U43966 (N_43966,N_41682,N_41351);
and U43967 (N_43967,N_41658,N_42151);
nor U43968 (N_43968,N_42169,N_41366);
nand U43969 (N_43969,N_40644,N_40374);
nand U43970 (N_43970,N_41761,N_41617);
and U43971 (N_43971,N_41978,N_41250);
or U43972 (N_43972,N_40643,N_41328);
and U43973 (N_43973,N_40131,N_40614);
xnor U43974 (N_43974,N_41147,N_41715);
and U43975 (N_43975,N_41479,N_42273);
xor U43976 (N_43976,N_41094,N_40481);
and U43977 (N_43977,N_41303,N_40750);
nand U43978 (N_43978,N_42445,N_40327);
xnor U43979 (N_43979,N_41910,N_42430);
nor U43980 (N_43980,N_41296,N_41049);
and U43981 (N_43981,N_41439,N_42177);
or U43982 (N_43982,N_40889,N_40805);
nor U43983 (N_43983,N_40605,N_42474);
nand U43984 (N_43984,N_40039,N_40997);
nor U43985 (N_43985,N_40984,N_41808);
nand U43986 (N_43986,N_41394,N_41663);
xor U43987 (N_43987,N_41527,N_41319);
nand U43988 (N_43988,N_40012,N_41009);
nand U43989 (N_43989,N_41062,N_42401);
or U43990 (N_43990,N_40641,N_41003);
nand U43991 (N_43991,N_41793,N_41445);
or U43992 (N_43992,N_41629,N_41408);
nor U43993 (N_43993,N_42444,N_41667);
nor U43994 (N_43994,N_41418,N_41907);
or U43995 (N_43995,N_41186,N_40332);
xnor U43996 (N_43996,N_40080,N_42066);
nand U43997 (N_43997,N_40655,N_42278);
nand U43998 (N_43998,N_42183,N_42134);
nor U43999 (N_43999,N_41777,N_41823);
or U44000 (N_44000,N_42035,N_41462);
xnor U44001 (N_44001,N_40445,N_40503);
xnor U44002 (N_44002,N_42065,N_41801);
xor U44003 (N_44003,N_40696,N_41849);
and U44004 (N_44004,N_41075,N_41523);
nor U44005 (N_44005,N_41082,N_41883);
nor U44006 (N_44006,N_41523,N_41427);
and U44007 (N_44007,N_41306,N_40568);
nand U44008 (N_44008,N_41977,N_41741);
nand U44009 (N_44009,N_40774,N_41409);
xnor U44010 (N_44010,N_41247,N_41451);
nand U44011 (N_44011,N_41318,N_42014);
or U44012 (N_44012,N_40438,N_42170);
nand U44013 (N_44013,N_41700,N_40082);
nand U44014 (N_44014,N_42091,N_41018);
nand U44015 (N_44015,N_40069,N_41972);
nor U44016 (N_44016,N_42121,N_41370);
xor U44017 (N_44017,N_40910,N_40030);
nand U44018 (N_44018,N_41885,N_42126);
nor U44019 (N_44019,N_40298,N_40338);
or U44020 (N_44020,N_41750,N_40063);
nor U44021 (N_44021,N_42206,N_41369);
nand U44022 (N_44022,N_42450,N_41660);
and U44023 (N_44023,N_40977,N_41493);
nor U44024 (N_44024,N_41280,N_42401);
or U44025 (N_44025,N_42413,N_40100);
and U44026 (N_44026,N_41782,N_42070);
or U44027 (N_44027,N_41329,N_40949);
xnor U44028 (N_44028,N_40491,N_40123);
xnor U44029 (N_44029,N_42174,N_42037);
and U44030 (N_44030,N_41745,N_41475);
and U44031 (N_44031,N_41187,N_40317);
and U44032 (N_44032,N_41387,N_41527);
or U44033 (N_44033,N_41869,N_40969);
or U44034 (N_44034,N_42141,N_42032);
or U44035 (N_44035,N_41901,N_41573);
nand U44036 (N_44036,N_41539,N_41965);
xor U44037 (N_44037,N_41799,N_40578);
xor U44038 (N_44038,N_41814,N_41011);
nand U44039 (N_44039,N_41946,N_42217);
nor U44040 (N_44040,N_41000,N_40093);
xnor U44041 (N_44041,N_42461,N_42110);
or U44042 (N_44042,N_40808,N_41146);
nor U44043 (N_44043,N_41372,N_40932);
nand U44044 (N_44044,N_40797,N_41647);
or U44045 (N_44045,N_40482,N_40845);
or U44046 (N_44046,N_40711,N_40096);
nand U44047 (N_44047,N_41521,N_40623);
and U44048 (N_44048,N_41424,N_40223);
or U44049 (N_44049,N_41953,N_40222);
or U44050 (N_44050,N_41329,N_40369);
nor U44051 (N_44051,N_41555,N_41910);
nor U44052 (N_44052,N_41815,N_40661);
nor U44053 (N_44053,N_40108,N_41267);
or U44054 (N_44054,N_40723,N_42187);
nor U44055 (N_44055,N_42021,N_40065);
nand U44056 (N_44056,N_40520,N_41634);
nand U44057 (N_44057,N_40041,N_42412);
nand U44058 (N_44058,N_40969,N_41876);
nor U44059 (N_44059,N_42195,N_42337);
nand U44060 (N_44060,N_41346,N_40062);
nor U44061 (N_44061,N_41555,N_42307);
xor U44062 (N_44062,N_40628,N_40967);
and U44063 (N_44063,N_40362,N_41153);
or U44064 (N_44064,N_41244,N_41527);
nor U44065 (N_44065,N_41805,N_40594);
xnor U44066 (N_44066,N_40874,N_41551);
xnor U44067 (N_44067,N_41670,N_41460);
nand U44068 (N_44068,N_40854,N_41157);
nor U44069 (N_44069,N_41246,N_41403);
and U44070 (N_44070,N_40672,N_40612);
nand U44071 (N_44071,N_40739,N_40448);
nor U44072 (N_44072,N_42057,N_42027);
nand U44073 (N_44073,N_41305,N_42281);
and U44074 (N_44074,N_42182,N_41633);
xor U44075 (N_44075,N_42416,N_40589);
xnor U44076 (N_44076,N_41708,N_41424);
or U44077 (N_44077,N_40577,N_40660);
nor U44078 (N_44078,N_41177,N_40124);
or U44079 (N_44079,N_40778,N_40364);
nand U44080 (N_44080,N_40387,N_41840);
nand U44081 (N_44081,N_40682,N_40159);
or U44082 (N_44082,N_40488,N_40689);
or U44083 (N_44083,N_41362,N_41732);
nor U44084 (N_44084,N_40504,N_40743);
and U44085 (N_44085,N_41671,N_41014);
and U44086 (N_44086,N_41191,N_40085);
and U44087 (N_44087,N_42286,N_40986);
nor U44088 (N_44088,N_42347,N_41374);
nand U44089 (N_44089,N_40567,N_41657);
xnor U44090 (N_44090,N_40222,N_40751);
xor U44091 (N_44091,N_41162,N_40984);
nor U44092 (N_44092,N_40243,N_41158);
xnor U44093 (N_44093,N_40643,N_42035);
or U44094 (N_44094,N_40376,N_40313);
nor U44095 (N_44095,N_40403,N_41473);
nor U44096 (N_44096,N_41295,N_41449);
nor U44097 (N_44097,N_40876,N_41886);
nand U44098 (N_44098,N_41470,N_42096);
nor U44099 (N_44099,N_42278,N_40805);
or U44100 (N_44100,N_40746,N_42328);
nand U44101 (N_44101,N_41242,N_40945);
xnor U44102 (N_44102,N_41862,N_40647);
nor U44103 (N_44103,N_40346,N_41122);
and U44104 (N_44104,N_41048,N_42204);
xor U44105 (N_44105,N_42428,N_40288);
xnor U44106 (N_44106,N_41265,N_40164);
nor U44107 (N_44107,N_40524,N_40940);
xnor U44108 (N_44108,N_42435,N_41361);
nor U44109 (N_44109,N_41102,N_41934);
and U44110 (N_44110,N_42195,N_41300);
xor U44111 (N_44111,N_42414,N_41479);
nor U44112 (N_44112,N_40870,N_41588);
nor U44113 (N_44113,N_42449,N_42226);
nand U44114 (N_44114,N_41176,N_41749);
and U44115 (N_44115,N_41815,N_42299);
and U44116 (N_44116,N_40201,N_41923);
or U44117 (N_44117,N_40976,N_40933);
xnor U44118 (N_44118,N_40311,N_41057);
and U44119 (N_44119,N_41671,N_41429);
nand U44120 (N_44120,N_41538,N_42463);
nor U44121 (N_44121,N_40928,N_41021);
nor U44122 (N_44122,N_41463,N_41483);
nor U44123 (N_44123,N_40884,N_40318);
xnor U44124 (N_44124,N_41710,N_41678);
and U44125 (N_44125,N_42429,N_42175);
xnor U44126 (N_44126,N_42349,N_41539);
nor U44127 (N_44127,N_40506,N_41394);
and U44128 (N_44128,N_41655,N_42113);
or U44129 (N_44129,N_42113,N_42018);
nand U44130 (N_44130,N_41177,N_41833);
nand U44131 (N_44131,N_42275,N_42184);
nor U44132 (N_44132,N_40839,N_42060);
or U44133 (N_44133,N_41978,N_40787);
or U44134 (N_44134,N_42234,N_40759);
nor U44135 (N_44135,N_41688,N_42399);
xnor U44136 (N_44136,N_41886,N_41042);
or U44137 (N_44137,N_40541,N_41156);
nand U44138 (N_44138,N_40928,N_40743);
or U44139 (N_44139,N_40315,N_41982);
or U44140 (N_44140,N_41788,N_40471);
or U44141 (N_44141,N_41055,N_41109);
nor U44142 (N_44142,N_42088,N_41038);
nor U44143 (N_44143,N_41016,N_41014);
and U44144 (N_44144,N_40571,N_42143);
or U44145 (N_44145,N_41532,N_41761);
xor U44146 (N_44146,N_40230,N_42233);
xor U44147 (N_44147,N_40504,N_42407);
xnor U44148 (N_44148,N_41996,N_41030);
and U44149 (N_44149,N_41068,N_40052);
or U44150 (N_44150,N_41843,N_41662);
or U44151 (N_44151,N_40058,N_40281);
nor U44152 (N_44152,N_40417,N_41284);
or U44153 (N_44153,N_41125,N_40855);
nor U44154 (N_44154,N_41941,N_41534);
and U44155 (N_44155,N_40873,N_41912);
xor U44156 (N_44156,N_40556,N_40455);
or U44157 (N_44157,N_40635,N_40768);
and U44158 (N_44158,N_40790,N_41881);
nand U44159 (N_44159,N_42478,N_41041);
and U44160 (N_44160,N_41399,N_41560);
or U44161 (N_44161,N_41753,N_41473);
or U44162 (N_44162,N_40121,N_40103);
nand U44163 (N_44163,N_42345,N_40105);
or U44164 (N_44164,N_41775,N_40109);
nand U44165 (N_44165,N_41667,N_41403);
and U44166 (N_44166,N_41769,N_41584);
or U44167 (N_44167,N_40217,N_40473);
and U44168 (N_44168,N_41344,N_40941);
and U44169 (N_44169,N_41112,N_40638);
and U44170 (N_44170,N_40819,N_40729);
xor U44171 (N_44171,N_41679,N_41761);
nor U44172 (N_44172,N_41584,N_40068);
xor U44173 (N_44173,N_40211,N_40823);
nand U44174 (N_44174,N_41385,N_40003);
and U44175 (N_44175,N_41619,N_40099);
nand U44176 (N_44176,N_40010,N_41294);
nand U44177 (N_44177,N_40675,N_41834);
xor U44178 (N_44178,N_41613,N_41466);
xor U44179 (N_44179,N_40394,N_40830);
nand U44180 (N_44180,N_42485,N_42151);
and U44181 (N_44181,N_40608,N_40903);
or U44182 (N_44182,N_42291,N_42133);
or U44183 (N_44183,N_42050,N_40852);
nor U44184 (N_44184,N_41099,N_41080);
xor U44185 (N_44185,N_40017,N_41201);
and U44186 (N_44186,N_40027,N_40546);
or U44187 (N_44187,N_41950,N_41934);
or U44188 (N_44188,N_40737,N_42308);
and U44189 (N_44189,N_41610,N_42268);
and U44190 (N_44190,N_42248,N_41655);
and U44191 (N_44191,N_40673,N_41404);
nor U44192 (N_44192,N_40143,N_41748);
and U44193 (N_44193,N_42327,N_41657);
xor U44194 (N_44194,N_42231,N_42148);
or U44195 (N_44195,N_41677,N_41651);
or U44196 (N_44196,N_42109,N_42187);
nand U44197 (N_44197,N_40132,N_40789);
nor U44198 (N_44198,N_40700,N_42032);
xor U44199 (N_44199,N_41401,N_40578);
and U44200 (N_44200,N_41819,N_41724);
or U44201 (N_44201,N_42264,N_40286);
or U44202 (N_44202,N_40061,N_41227);
xor U44203 (N_44203,N_40542,N_40258);
and U44204 (N_44204,N_40242,N_40932);
and U44205 (N_44205,N_40808,N_42047);
or U44206 (N_44206,N_40799,N_41818);
xnor U44207 (N_44207,N_42167,N_41680);
xnor U44208 (N_44208,N_41402,N_41631);
and U44209 (N_44209,N_40155,N_40540);
nor U44210 (N_44210,N_41924,N_40837);
nor U44211 (N_44211,N_40110,N_41443);
and U44212 (N_44212,N_41828,N_40370);
xnor U44213 (N_44213,N_41060,N_40817);
nand U44214 (N_44214,N_40605,N_40442);
xnor U44215 (N_44215,N_40486,N_41001);
and U44216 (N_44216,N_42036,N_41623);
or U44217 (N_44217,N_40113,N_41029);
or U44218 (N_44218,N_41385,N_41076);
or U44219 (N_44219,N_40080,N_41453);
xnor U44220 (N_44220,N_40257,N_42089);
or U44221 (N_44221,N_41613,N_41416);
xnor U44222 (N_44222,N_41339,N_41089);
nand U44223 (N_44223,N_41683,N_40944);
and U44224 (N_44224,N_40826,N_42495);
or U44225 (N_44225,N_40261,N_42066);
nor U44226 (N_44226,N_41185,N_40389);
nand U44227 (N_44227,N_42117,N_40888);
or U44228 (N_44228,N_40537,N_41769);
and U44229 (N_44229,N_42376,N_41487);
nor U44230 (N_44230,N_42246,N_41504);
and U44231 (N_44231,N_40186,N_41690);
nor U44232 (N_44232,N_42367,N_40101);
or U44233 (N_44233,N_42207,N_40505);
nor U44234 (N_44234,N_40063,N_40684);
xnor U44235 (N_44235,N_42200,N_41755);
and U44236 (N_44236,N_40323,N_41396);
or U44237 (N_44237,N_41244,N_40942);
and U44238 (N_44238,N_40307,N_41991);
nand U44239 (N_44239,N_41610,N_40185);
and U44240 (N_44240,N_40074,N_41018);
or U44241 (N_44241,N_41217,N_41557);
and U44242 (N_44242,N_42240,N_41461);
and U44243 (N_44243,N_40190,N_41996);
and U44244 (N_44244,N_42290,N_40750);
nor U44245 (N_44245,N_40446,N_40379);
xnor U44246 (N_44246,N_41278,N_40152);
or U44247 (N_44247,N_40877,N_41285);
and U44248 (N_44248,N_42328,N_42489);
or U44249 (N_44249,N_40272,N_41440);
xor U44250 (N_44250,N_42138,N_40581);
and U44251 (N_44251,N_41161,N_40192);
nand U44252 (N_44252,N_42216,N_41155);
or U44253 (N_44253,N_41263,N_40271);
nand U44254 (N_44254,N_40806,N_40918);
nor U44255 (N_44255,N_40969,N_41006);
nand U44256 (N_44256,N_40510,N_40432);
nor U44257 (N_44257,N_42260,N_41221);
or U44258 (N_44258,N_42348,N_41717);
nand U44259 (N_44259,N_40663,N_40976);
or U44260 (N_44260,N_40433,N_42083);
nand U44261 (N_44261,N_41925,N_41733);
xnor U44262 (N_44262,N_41618,N_41745);
nand U44263 (N_44263,N_40178,N_40078);
nand U44264 (N_44264,N_40495,N_40808);
and U44265 (N_44265,N_42150,N_40289);
nand U44266 (N_44266,N_40357,N_40517);
nor U44267 (N_44267,N_41531,N_40137);
or U44268 (N_44268,N_40591,N_41651);
or U44269 (N_44269,N_40571,N_41109);
nor U44270 (N_44270,N_42018,N_42371);
xor U44271 (N_44271,N_41081,N_40147);
nor U44272 (N_44272,N_40299,N_41636);
nand U44273 (N_44273,N_42427,N_41709);
nand U44274 (N_44274,N_40863,N_40858);
nand U44275 (N_44275,N_40989,N_42139);
nor U44276 (N_44276,N_41536,N_40874);
or U44277 (N_44277,N_40264,N_40775);
xnor U44278 (N_44278,N_42204,N_42158);
nor U44279 (N_44279,N_42135,N_42088);
nor U44280 (N_44280,N_40293,N_41372);
or U44281 (N_44281,N_41068,N_40452);
or U44282 (N_44282,N_41310,N_40399);
or U44283 (N_44283,N_41738,N_40464);
xor U44284 (N_44284,N_40506,N_40063);
nor U44285 (N_44285,N_41124,N_40226);
nor U44286 (N_44286,N_41323,N_41677);
and U44287 (N_44287,N_40629,N_40476);
nor U44288 (N_44288,N_42234,N_40394);
nor U44289 (N_44289,N_41879,N_41082);
or U44290 (N_44290,N_41699,N_40221);
and U44291 (N_44291,N_41279,N_41930);
and U44292 (N_44292,N_40421,N_40357);
nand U44293 (N_44293,N_40482,N_41572);
or U44294 (N_44294,N_41274,N_42308);
and U44295 (N_44295,N_40309,N_40460);
nor U44296 (N_44296,N_40277,N_41111);
nor U44297 (N_44297,N_42190,N_40539);
xor U44298 (N_44298,N_41029,N_40381);
nand U44299 (N_44299,N_42207,N_40009);
and U44300 (N_44300,N_40802,N_40725);
xor U44301 (N_44301,N_41260,N_41205);
nor U44302 (N_44302,N_41459,N_41783);
and U44303 (N_44303,N_41647,N_40264);
nand U44304 (N_44304,N_41603,N_42210);
nor U44305 (N_44305,N_42276,N_40988);
xnor U44306 (N_44306,N_40534,N_41519);
or U44307 (N_44307,N_41124,N_40645);
and U44308 (N_44308,N_40722,N_41902);
nand U44309 (N_44309,N_41726,N_42415);
nor U44310 (N_44310,N_41113,N_41296);
nor U44311 (N_44311,N_40646,N_42369);
nor U44312 (N_44312,N_42318,N_40419);
and U44313 (N_44313,N_41530,N_41856);
nand U44314 (N_44314,N_40357,N_40834);
xor U44315 (N_44315,N_42101,N_41485);
or U44316 (N_44316,N_40388,N_41604);
and U44317 (N_44317,N_42363,N_41616);
and U44318 (N_44318,N_40967,N_41634);
or U44319 (N_44319,N_41304,N_40117);
and U44320 (N_44320,N_40108,N_41269);
nand U44321 (N_44321,N_40566,N_42216);
or U44322 (N_44322,N_42267,N_42407);
nor U44323 (N_44323,N_41105,N_40859);
or U44324 (N_44324,N_41979,N_41486);
or U44325 (N_44325,N_41299,N_41684);
nor U44326 (N_44326,N_40376,N_41540);
nand U44327 (N_44327,N_42249,N_40030);
xor U44328 (N_44328,N_41021,N_40026);
or U44329 (N_44329,N_40594,N_40189);
or U44330 (N_44330,N_41448,N_41341);
nand U44331 (N_44331,N_41393,N_41906);
nor U44332 (N_44332,N_40616,N_40021);
nand U44333 (N_44333,N_42143,N_40000);
nor U44334 (N_44334,N_41364,N_40438);
xor U44335 (N_44335,N_40389,N_41198);
nand U44336 (N_44336,N_41417,N_40500);
nor U44337 (N_44337,N_40027,N_41947);
and U44338 (N_44338,N_41749,N_41713);
xnor U44339 (N_44339,N_41577,N_40324);
and U44340 (N_44340,N_41878,N_41985);
or U44341 (N_44341,N_40093,N_40977);
and U44342 (N_44342,N_41286,N_40357);
nand U44343 (N_44343,N_42028,N_40002);
nand U44344 (N_44344,N_41556,N_40559);
and U44345 (N_44345,N_40037,N_41654);
xor U44346 (N_44346,N_41823,N_40629);
or U44347 (N_44347,N_41937,N_40566);
nor U44348 (N_44348,N_41096,N_40599);
or U44349 (N_44349,N_42302,N_40898);
nor U44350 (N_44350,N_40931,N_40988);
xor U44351 (N_44351,N_41822,N_40129);
and U44352 (N_44352,N_40389,N_41581);
nor U44353 (N_44353,N_41650,N_42062);
nand U44354 (N_44354,N_41216,N_40989);
xor U44355 (N_44355,N_40659,N_40544);
nor U44356 (N_44356,N_40177,N_40857);
nand U44357 (N_44357,N_41732,N_42189);
nor U44358 (N_44358,N_42071,N_40419);
xor U44359 (N_44359,N_41477,N_40958);
xor U44360 (N_44360,N_40939,N_40316);
nor U44361 (N_44361,N_41004,N_40228);
or U44362 (N_44362,N_40609,N_42232);
nor U44363 (N_44363,N_41332,N_41092);
xnor U44364 (N_44364,N_41293,N_41386);
nand U44365 (N_44365,N_42035,N_41999);
xnor U44366 (N_44366,N_40343,N_41491);
xnor U44367 (N_44367,N_41536,N_41797);
or U44368 (N_44368,N_40740,N_40559);
nand U44369 (N_44369,N_42150,N_40701);
or U44370 (N_44370,N_41933,N_41122);
nor U44371 (N_44371,N_40900,N_42356);
nand U44372 (N_44372,N_40753,N_41364);
nor U44373 (N_44373,N_42104,N_42153);
nor U44374 (N_44374,N_40550,N_41510);
nand U44375 (N_44375,N_42422,N_41343);
and U44376 (N_44376,N_42224,N_40929);
or U44377 (N_44377,N_41158,N_41529);
nor U44378 (N_44378,N_41901,N_41643);
and U44379 (N_44379,N_41486,N_40667);
nand U44380 (N_44380,N_41341,N_41902);
xnor U44381 (N_44381,N_40912,N_41892);
nor U44382 (N_44382,N_41866,N_40141);
or U44383 (N_44383,N_41948,N_40555);
or U44384 (N_44384,N_40685,N_40954);
nand U44385 (N_44385,N_41988,N_41341);
xor U44386 (N_44386,N_42119,N_40441);
xnor U44387 (N_44387,N_41640,N_42229);
nand U44388 (N_44388,N_40479,N_41698);
xor U44389 (N_44389,N_40462,N_40854);
nand U44390 (N_44390,N_41546,N_42432);
or U44391 (N_44391,N_40373,N_41986);
or U44392 (N_44392,N_40747,N_41296);
nor U44393 (N_44393,N_40836,N_40475);
nand U44394 (N_44394,N_40004,N_41694);
or U44395 (N_44395,N_41265,N_40740);
xnor U44396 (N_44396,N_42103,N_42260);
nand U44397 (N_44397,N_40180,N_40069);
nor U44398 (N_44398,N_41928,N_40970);
and U44399 (N_44399,N_41348,N_41717);
nand U44400 (N_44400,N_42265,N_40416);
or U44401 (N_44401,N_41484,N_42092);
or U44402 (N_44402,N_40889,N_40750);
xor U44403 (N_44403,N_41587,N_40942);
and U44404 (N_44404,N_42193,N_41837);
xor U44405 (N_44405,N_42331,N_40073);
xor U44406 (N_44406,N_40855,N_42121);
and U44407 (N_44407,N_41635,N_41101);
or U44408 (N_44408,N_40145,N_41837);
nand U44409 (N_44409,N_40448,N_41275);
nor U44410 (N_44410,N_40585,N_40609);
nor U44411 (N_44411,N_41903,N_40721);
nand U44412 (N_44412,N_41311,N_41666);
nand U44413 (N_44413,N_40183,N_42296);
nand U44414 (N_44414,N_41127,N_40994);
and U44415 (N_44415,N_40987,N_41283);
nor U44416 (N_44416,N_40030,N_41432);
nor U44417 (N_44417,N_40928,N_40887);
nand U44418 (N_44418,N_41783,N_40674);
nor U44419 (N_44419,N_41573,N_40221);
nand U44420 (N_44420,N_41926,N_40777);
nor U44421 (N_44421,N_41541,N_40300);
nor U44422 (N_44422,N_41290,N_41853);
nor U44423 (N_44423,N_41042,N_41942);
or U44424 (N_44424,N_40574,N_40334);
or U44425 (N_44425,N_40038,N_40655);
xnor U44426 (N_44426,N_40761,N_42438);
and U44427 (N_44427,N_42421,N_40352);
nand U44428 (N_44428,N_42313,N_41509);
xor U44429 (N_44429,N_40785,N_41108);
nand U44430 (N_44430,N_40494,N_40236);
or U44431 (N_44431,N_42141,N_41299);
nor U44432 (N_44432,N_41352,N_42351);
nand U44433 (N_44433,N_41423,N_40394);
xor U44434 (N_44434,N_40227,N_41496);
and U44435 (N_44435,N_42211,N_41258);
and U44436 (N_44436,N_40617,N_40874);
and U44437 (N_44437,N_40225,N_42084);
nor U44438 (N_44438,N_40628,N_42003);
xor U44439 (N_44439,N_41739,N_41442);
and U44440 (N_44440,N_42450,N_42115);
nand U44441 (N_44441,N_40496,N_40984);
xnor U44442 (N_44442,N_41578,N_41588);
and U44443 (N_44443,N_41043,N_40745);
nand U44444 (N_44444,N_42178,N_42458);
xnor U44445 (N_44445,N_40322,N_41323);
and U44446 (N_44446,N_40693,N_41794);
nor U44447 (N_44447,N_40562,N_42427);
and U44448 (N_44448,N_40038,N_41380);
nor U44449 (N_44449,N_41964,N_40175);
xnor U44450 (N_44450,N_41838,N_42294);
nor U44451 (N_44451,N_41036,N_42411);
xor U44452 (N_44452,N_42148,N_41273);
nor U44453 (N_44453,N_42383,N_42075);
or U44454 (N_44454,N_40756,N_42256);
and U44455 (N_44455,N_40392,N_40420);
nor U44456 (N_44456,N_42157,N_41892);
nand U44457 (N_44457,N_40162,N_40308);
nand U44458 (N_44458,N_40202,N_42444);
or U44459 (N_44459,N_41749,N_42222);
xor U44460 (N_44460,N_41803,N_41168);
nand U44461 (N_44461,N_40539,N_42377);
xnor U44462 (N_44462,N_42226,N_40696);
nor U44463 (N_44463,N_40225,N_40626);
or U44464 (N_44464,N_40847,N_40232);
and U44465 (N_44465,N_40390,N_42262);
nor U44466 (N_44466,N_40540,N_40561);
nor U44467 (N_44467,N_40490,N_40071);
or U44468 (N_44468,N_40084,N_40556);
or U44469 (N_44469,N_42472,N_40176);
and U44470 (N_44470,N_41981,N_41361);
xnor U44471 (N_44471,N_40870,N_40019);
nor U44472 (N_44472,N_42248,N_41891);
nor U44473 (N_44473,N_42014,N_41653);
nor U44474 (N_44474,N_41391,N_41059);
and U44475 (N_44475,N_41679,N_41340);
xnor U44476 (N_44476,N_42269,N_42119);
xor U44477 (N_44477,N_41624,N_40376);
nand U44478 (N_44478,N_40033,N_42240);
xor U44479 (N_44479,N_40679,N_41161);
or U44480 (N_44480,N_40697,N_42061);
xor U44481 (N_44481,N_40858,N_40329);
nand U44482 (N_44482,N_40142,N_41728);
nor U44483 (N_44483,N_40853,N_40837);
xor U44484 (N_44484,N_41170,N_41003);
nor U44485 (N_44485,N_41982,N_40577);
and U44486 (N_44486,N_41755,N_40560);
nor U44487 (N_44487,N_42359,N_41939);
xnor U44488 (N_44488,N_42244,N_40786);
or U44489 (N_44489,N_42062,N_41766);
xnor U44490 (N_44490,N_42017,N_40330);
and U44491 (N_44491,N_41535,N_40201);
nor U44492 (N_44492,N_40742,N_42302);
xnor U44493 (N_44493,N_42264,N_41298);
or U44494 (N_44494,N_40459,N_41613);
and U44495 (N_44495,N_41347,N_40531);
xnor U44496 (N_44496,N_40071,N_41940);
and U44497 (N_44497,N_40141,N_40537);
or U44498 (N_44498,N_41100,N_41967);
nand U44499 (N_44499,N_40818,N_40088);
and U44500 (N_44500,N_41399,N_42443);
xnor U44501 (N_44501,N_41723,N_40882);
or U44502 (N_44502,N_40048,N_40385);
xnor U44503 (N_44503,N_40384,N_41569);
nor U44504 (N_44504,N_40446,N_40440);
xor U44505 (N_44505,N_41673,N_41363);
and U44506 (N_44506,N_40369,N_41976);
and U44507 (N_44507,N_41884,N_40643);
or U44508 (N_44508,N_42265,N_40625);
and U44509 (N_44509,N_40018,N_41873);
and U44510 (N_44510,N_41061,N_40825);
xor U44511 (N_44511,N_41128,N_40459);
nand U44512 (N_44512,N_41880,N_42047);
nand U44513 (N_44513,N_41924,N_40825);
xnor U44514 (N_44514,N_41938,N_40725);
or U44515 (N_44515,N_41838,N_40302);
or U44516 (N_44516,N_42016,N_41579);
xor U44517 (N_44517,N_41406,N_42480);
and U44518 (N_44518,N_42065,N_41048);
nand U44519 (N_44519,N_41744,N_40528);
or U44520 (N_44520,N_40565,N_40113);
xor U44521 (N_44521,N_40727,N_42006);
xnor U44522 (N_44522,N_40945,N_41469);
and U44523 (N_44523,N_42165,N_40075);
or U44524 (N_44524,N_41682,N_40502);
nand U44525 (N_44525,N_40723,N_42120);
xor U44526 (N_44526,N_42394,N_40807);
and U44527 (N_44527,N_41660,N_40800);
nor U44528 (N_44528,N_40043,N_41919);
or U44529 (N_44529,N_40648,N_40501);
xor U44530 (N_44530,N_41464,N_40437);
nor U44531 (N_44531,N_41053,N_41810);
nand U44532 (N_44532,N_41154,N_42169);
xnor U44533 (N_44533,N_41255,N_40857);
nand U44534 (N_44534,N_41694,N_41943);
or U44535 (N_44535,N_40594,N_41716);
or U44536 (N_44536,N_40614,N_41577);
and U44537 (N_44537,N_41328,N_41824);
nor U44538 (N_44538,N_41886,N_41615);
nor U44539 (N_44539,N_41577,N_42085);
nor U44540 (N_44540,N_42413,N_41343);
and U44541 (N_44541,N_40027,N_40564);
or U44542 (N_44542,N_40364,N_41561);
xnor U44543 (N_44543,N_42278,N_41948);
nor U44544 (N_44544,N_41194,N_41045);
nor U44545 (N_44545,N_40485,N_40787);
nor U44546 (N_44546,N_41131,N_41806);
nor U44547 (N_44547,N_42442,N_40802);
xor U44548 (N_44548,N_41396,N_40836);
xor U44549 (N_44549,N_41346,N_40694);
xnor U44550 (N_44550,N_40622,N_40613);
or U44551 (N_44551,N_42053,N_40033);
or U44552 (N_44552,N_41847,N_41104);
and U44553 (N_44553,N_41061,N_40012);
or U44554 (N_44554,N_40683,N_41024);
nand U44555 (N_44555,N_41823,N_40462);
or U44556 (N_44556,N_41128,N_40254);
or U44557 (N_44557,N_41102,N_41813);
nand U44558 (N_44558,N_41829,N_41014);
xnor U44559 (N_44559,N_42045,N_41662);
or U44560 (N_44560,N_42102,N_41397);
xnor U44561 (N_44561,N_40369,N_42194);
xnor U44562 (N_44562,N_41427,N_41539);
and U44563 (N_44563,N_40046,N_41787);
nor U44564 (N_44564,N_40034,N_41161);
nor U44565 (N_44565,N_40282,N_40011);
xnor U44566 (N_44566,N_41059,N_42046);
or U44567 (N_44567,N_41492,N_40688);
or U44568 (N_44568,N_41997,N_41581);
nor U44569 (N_44569,N_40713,N_41563);
and U44570 (N_44570,N_40847,N_40665);
nor U44571 (N_44571,N_41527,N_40630);
nand U44572 (N_44572,N_40214,N_40193);
nand U44573 (N_44573,N_42145,N_41523);
and U44574 (N_44574,N_42354,N_41842);
nand U44575 (N_44575,N_41365,N_41404);
nor U44576 (N_44576,N_40075,N_40330);
and U44577 (N_44577,N_42091,N_41094);
nor U44578 (N_44578,N_41469,N_41543);
and U44579 (N_44579,N_42358,N_40291);
nand U44580 (N_44580,N_40536,N_40452);
and U44581 (N_44581,N_41780,N_40724);
xnor U44582 (N_44582,N_42392,N_42411);
nand U44583 (N_44583,N_41755,N_40118);
nand U44584 (N_44584,N_42204,N_40764);
nand U44585 (N_44585,N_40781,N_40052);
nor U44586 (N_44586,N_40171,N_42152);
nor U44587 (N_44587,N_40729,N_40896);
or U44588 (N_44588,N_40404,N_40703);
nand U44589 (N_44589,N_41965,N_41785);
xnor U44590 (N_44590,N_42189,N_42006);
nor U44591 (N_44591,N_40239,N_40048);
nor U44592 (N_44592,N_42084,N_40136);
or U44593 (N_44593,N_41190,N_41007);
xnor U44594 (N_44594,N_42423,N_41710);
xor U44595 (N_44595,N_40622,N_41748);
xnor U44596 (N_44596,N_41169,N_40821);
and U44597 (N_44597,N_41266,N_41232);
xor U44598 (N_44598,N_40531,N_41792);
nand U44599 (N_44599,N_42231,N_40903);
nor U44600 (N_44600,N_42167,N_42126);
and U44601 (N_44601,N_41122,N_42479);
nor U44602 (N_44602,N_42421,N_41203);
nor U44603 (N_44603,N_41010,N_40124);
nor U44604 (N_44604,N_40084,N_41195);
and U44605 (N_44605,N_40556,N_41174);
and U44606 (N_44606,N_42350,N_41223);
and U44607 (N_44607,N_40449,N_41439);
and U44608 (N_44608,N_40605,N_41755);
nand U44609 (N_44609,N_40434,N_41391);
or U44610 (N_44610,N_40954,N_40396);
nor U44611 (N_44611,N_40190,N_41916);
xor U44612 (N_44612,N_40986,N_40492);
nand U44613 (N_44613,N_41899,N_40383);
xnor U44614 (N_44614,N_41924,N_40180);
xor U44615 (N_44615,N_40298,N_40960);
or U44616 (N_44616,N_41165,N_41028);
or U44617 (N_44617,N_41900,N_41663);
nand U44618 (N_44618,N_40401,N_41719);
xor U44619 (N_44619,N_40121,N_41072);
or U44620 (N_44620,N_41606,N_41278);
xor U44621 (N_44621,N_40833,N_40794);
or U44622 (N_44622,N_40103,N_41732);
nand U44623 (N_44623,N_41956,N_41757);
and U44624 (N_44624,N_40094,N_40961);
nor U44625 (N_44625,N_42203,N_40263);
nor U44626 (N_44626,N_41033,N_40462);
nand U44627 (N_44627,N_40349,N_40332);
nor U44628 (N_44628,N_41213,N_42248);
and U44629 (N_44629,N_41748,N_41563);
nor U44630 (N_44630,N_40320,N_41382);
xnor U44631 (N_44631,N_41698,N_40677);
nand U44632 (N_44632,N_40142,N_42481);
xor U44633 (N_44633,N_41941,N_41577);
or U44634 (N_44634,N_41542,N_41990);
or U44635 (N_44635,N_40152,N_40737);
nor U44636 (N_44636,N_40446,N_41629);
and U44637 (N_44637,N_42052,N_40885);
nor U44638 (N_44638,N_40724,N_41297);
or U44639 (N_44639,N_40951,N_40835);
or U44640 (N_44640,N_42245,N_42395);
xnor U44641 (N_44641,N_40345,N_41971);
xnor U44642 (N_44642,N_41461,N_41579);
nor U44643 (N_44643,N_40797,N_40773);
or U44644 (N_44644,N_40206,N_42333);
and U44645 (N_44645,N_41296,N_40341);
nor U44646 (N_44646,N_40124,N_40385);
xor U44647 (N_44647,N_40557,N_40617);
nand U44648 (N_44648,N_42216,N_40775);
nand U44649 (N_44649,N_41969,N_41179);
nand U44650 (N_44650,N_41641,N_40269);
or U44651 (N_44651,N_40363,N_41963);
nand U44652 (N_44652,N_40239,N_42300);
or U44653 (N_44653,N_42009,N_40155);
xnor U44654 (N_44654,N_40291,N_41150);
nor U44655 (N_44655,N_41126,N_40800);
xor U44656 (N_44656,N_40693,N_42494);
and U44657 (N_44657,N_41363,N_40618);
xnor U44658 (N_44658,N_41203,N_42346);
or U44659 (N_44659,N_40184,N_41412);
xor U44660 (N_44660,N_41479,N_42443);
nor U44661 (N_44661,N_40395,N_40174);
and U44662 (N_44662,N_40604,N_41916);
or U44663 (N_44663,N_40984,N_40653);
and U44664 (N_44664,N_42397,N_42110);
xor U44665 (N_44665,N_40351,N_40088);
nand U44666 (N_44666,N_42184,N_40046);
or U44667 (N_44667,N_41439,N_41483);
nor U44668 (N_44668,N_41088,N_42178);
xnor U44669 (N_44669,N_41813,N_40859);
and U44670 (N_44670,N_41161,N_41282);
or U44671 (N_44671,N_41182,N_40090);
xnor U44672 (N_44672,N_40161,N_41081);
nor U44673 (N_44673,N_41866,N_40790);
nand U44674 (N_44674,N_41941,N_41882);
and U44675 (N_44675,N_40532,N_41121);
xnor U44676 (N_44676,N_41127,N_40332);
nand U44677 (N_44677,N_40376,N_42408);
and U44678 (N_44678,N_40167,N_41837);
or U44679 (N_44679,N_40232,N_41045);
nor U44680 (N_44680,N_40790,N_41478);
or U44681 (N_44681,N_41392,N_42389);
and U44682 (N_44682,N_41149,N_41558);
and U44683 (N_44683,N_41001,N_41145);
nand U44684 (N_44684,N_41205,N_40651);
or U44685 (N_44685,N_41004,N_40765);
or U44686 (N_44686,N_41831,N_42145);
or U44687 (N_44687,N_41777,N_42280);
xnor U44688 (N_44688,N_41986,N_40368);
xor U44689 (N_44689,N_41950,N_41066);
and U44690 (N_44690,N_41851,N_42046);
or U44691 (N_44691,N_41819,N_42215);
nor U44692 (N_44692,N_40965,N_42001);
nand U44693 (N_44693,N_41381,N_41371);
and U44694 (N_44694,N_41764,N_40448);
and U44695 (N_44695,N_42457,N_40584);
and U44696 (N_44696,N_42190,N_40489);
nor U44697 (N_44697,N_41098,N_42051);
or U44698 (N_44698,N_41184,N_41497);
nand U44699 (N_44699,N_40495,N_40612);
nor U44700 (N_44700,N_41001,N_40552);
nor U44701 (N_44701,N_41206,N_41662);
and U44702 (N_44702,N_41446,N_40201);
nor U44703 (N_44703,N_41915,N_40400);
nor U44704 (N_44704,N_41170,N_42146);
nand U44705 (N_44705,N_40366,N_41282);
or U44706 (N_44706,N_41796,N_41825);
nor U44707 (N_44707,N_41291,N_41756);
or U44708 (N_44708,N_41762,N_41413);
nand U44709 (N_44709,N_42136,N_41329);
and U44710 (N_44710,N_42417,N_40744);
nand U44711 (N_44711,N_41553,N_42011);
xnor U44712 (N_44712,N_40749,N_40213);
and U44713 (N_44713,N_42274,N_41139);
nand U44714 (N_44714,N_41561,N_40279);
or U44715 (N_44715,N_40125,N_42320);
and U44716 (N_44716,N_42132,N_40003);
and U44717 (N_44717,N_41524,N_42168);
and U44718 (N_44718,N_41907,N_41618);
xnor U44719 (N_44719,N_41717,N_40798);
or U44720 (N_44720,N_42179,N_41909);
nand U44721 (N_44721,N_40909,N_41323);
xor U44722 (N_44722,N_40815,N_42476);
or U44723 (N_44723,N_41791,N_40792);
nand U44724 (N_44724,N_41360,N_40385);
and U44725 (N_44725,N_42154,N_41421);
nor U44726 (N_44726,N_42390,N_40665);
nand U44727 (N_44727,N_40823,N_42304);
nor U44728 (N_44728,N_40136,N_41972);
and U44729 (N_44729,N_42112,N_41858);
and U44730 (N_44730,N_41106,N_41746);
nand U44731 (N_44731,N_41952,N_41475);
xor U44732 (N_44732,N_41662,N_40496);
or U44733 (N_44733,N_41209,N_40052);
or U44734 (N_44734,N_40438,N_41409);
or U44735 (N_44735,N_42267,N_41401);
or U44736 (N_44736,N_40000,N_40761);
nor U44737 (N_44737,N_41211,N_42014);
xor U44738 (N_44738,N_42090,N_40276);
nand U44739 (N_44739,N_41307,N_40784);
nand U44740 (N_44740,N_40121,N_41480);
or U44741 (N_44741,N_42399,N_40240);
xnor U44742 (N_44742,N_40559,N_40731);
and U44743 (N_44743,N_40311,N_41928);
or U44744 (N_44744,N_41175,N_41939);
xnor U44745 (N_44745,N_40274,N_40876);
nor U44746 (N_44746,N_40408,N_41255);
nor U44747 (N_44747,N_40022,N_41159);
or U44748 (N_44748,N_41598,N_41438);
xnor U44749 (N_44749,N_42005,N_40933);
and U44750 (N_44750,N_41092,N_40517);
or U44751 (N_44751,N_40799,N_41176);
nand U44752 (N_44752,N_41523,N_42235);
xnor U44753 (N_44753,N_40456,N_41145);
nand U44754 (N_44754,N_40110,N_41482);
or U44755 (N_44755,N_41032,N_41014);
and U44756 (N_44756,N_42396,N_41898);
nor U44757 (N_44757,N_41292,N_41089);
xor U44758 (N_44758,N_41508,N_41160);
or U44759 (N_44759,N_41994,N_42285);
or U44760 (N_44760,N_42488,N_40809);
xor U44761 (N_44761,N_42429,N_42478);
or U44762 (N_44762,N_41822,N_40926);
nor U44763 (N_44763,N_41574,N_41794);
xnor U44764 (N_44764,N_41647,N_40332);
xor U44765 (N_44765,N_41199,N_42165);
or U44766 (N_44766,N_42179,N_40223);
nor U44767 (N_44767,N_41831,N_41905);
or U44768 (N_44768,N_40541,N_41103);
or U44769 (N_44769,N_40462,N_41419);
nand U44770 (N_44770,N_41150,N_40507);
xnor U44771 (N_44771,N_41418,N_40336);
and U44772 (N_44772,N_41500,N_40827);
and U44773 (N_44773,N_41496,N_42154);
nor U44774 (N_44774,N_41603,N_42124);
or U44775 (N_44775,N_42116,N_41751);
or U44776 (N_44776,N_41264,N_40630);
and U44777 (N_44777,N_42044,N_41391);
xor U44778 (N_44778,N_41910,N_41292);
nor U44779 (N_44779,N_40102,N_40208);
xnor U44780 (N_44780,N_42278,N_40674);
xor U44781 (N_44781,N_40534,N_40975);
nor U44782 (N_44782,N_41777,N_41307);
or U44783 (N_44783,N_40685,N_41080);
xnor U44784 (N_44784,N_40974,N_41841);
and U44785 (N_44785,N_42074,N_41515);
and U44786 (N_44786,N_42109,N_40008);
nand U44787 (N_44787,N_40118,N_40109);
xor U44788 (N_44788,N_42183,N_42294);
nand U44789 (N_44789,N_40522,N_40680);
and U44790 (N_44790,N_40046,N_41954);
nor U44791 (N_44791,N_40124,N_40199);
nor U44792 (N_44792,N_40291,N_40701);
or U44793 (N_44793,N_42474,N_40143);
nand U44794 (N_44794,N_42440,N_41684);
and U44795 (N_44795,N_42239,N_40850);
and U44796 (N_44796,N_40172,N_40493);
and U44797 (N_44797,N_40759,N_41908);
nand U44798 (N_44798,N_41000,N_40054);
nor U44799 (N_44799,N_41433,N_41017);
nand U44800 (N_44800,N_41236,N_40154);
and U44801 (N_44801,N_41672,N_40390);
nand U44802 (N_44802,N_40984,N_41469);
nand U44803 (N_44803,N_41565,N_41033);
nand U44804 (N_44804,N_40413,N_41276);
and U44805 (N_44805,N_42035,N_42420);
and U44806 (N_44806,N_40001,N_41987);
nand U44807 (N_44807,N_42249,N_42185);
nor U44808 (N_44808,N_41860,N_42462);
xor U44809 (N_44809,N_41739,N_42276);
xnor U44810 (N_44810,N_40999,N_42399);
nand U44811 (N_44811,N_41241,N_42259);
nor U44812 (N_44812,N_40233,N_42257);
nand U44813 (N_44813,N_42427,N_40869);
nor U44814 (N_44814,N_41581,N_41691);
or U44815 (N_44815,N_40977,N_40666);
xnor U44816 (N_44816,N_40264,N_41630);
or U44817 (N_44817,N_40174,N_42429);
xnor U44818 (N_44818,N_42267,N_41994);
or U44819 (N_44819,N_41316,N_41275);
nand U44820 (N_44820,N_40289,N_42136);
nand U44821 (N_44821,N_42156,N_40521);
nor U44822 (N_44822,N_41881,N_41773);
nand U44823 (N_44823,N_41246,N_40761);
or U44824 (N_44824,N_41301,N_41741);
xnor U44825 (N_44825,N_40544,N_40748);
nand U44826 (N_44826,N_41407,N_41697);
nand U44827 (N_44827,N_42337,N_40955);
and U44828 (N_44828,N_40499,N_40117);
xnor U44829 (N_44829,N_41226,N_40154);
nor U44830 (N_44830,N_41729,N_40398);
xor U44831 (N_44831,N_40079,N_40549);
and U44832 (N_44832,N_40741,N_42412);
or U44833 (N_44833,N_41181,N_41105);
nor U44834 (N_44834,N_40031,N_42326);
xor U44835 (N_44835,N_42202,N_41006);
xor U44836 (N_44836,N_41320,N_41693);
nand U44837 (N_44837,N_42285,N_40340);
nand U44838 (N_44838,N_41289,N_40003);
and U44839 (N_44839,N_41347,N_41101);
or U44840 (N_44840,N_41726,N_40319);
nor U44841 (N_44841,N_41128,N_42381);
xnor U44842 (N_44842,N_41559,N_40470);
and U44843 (N_44843,N_42172,N_40400);
nor U44844 (N_44844,N_40727,N_40406);
nor U44845 (N_44845,N_41386,N_41145);
and U44846 (N_44846,N_40998,N_41208);
nor U44847 (N_44847,N_42404,N_40793);
nand U44848 (N_44848,N_40326,N_41044);
nor U44849 (N_44849,N_40415,N_42257);
xor U44850 (N_44850,N_41722,N_40872);
and U44851 (N_44851,N_41723,N_41286);
nor U44852 (N_44852,N_40485,N_42005);
and U44853 (N_44853,N_41354,N_40590);
xnor U44854 (N_44854,N_41359,N_40640);
nand U44855 (N_44855,N_40869,N_42378);
nand U44856 (N_44856,N_40482,N_40255);
or U44857 (N_44857,N_40684,N_41626);
xnor U44858 (N_44858,N_40758,N_40484);
nand U44859 (N_44859,N_40145,N_40176);
nor U44860 (N_44860,N_42192,N_41711);
and U44861 (N_44861,N_42149,N_41892);
nand U44862 (N_44862,N_42402,N_42333);
nand U44863 (N_44863,N_40220,N_40764);
xor U44864 (N_44864,N_42020,N_42134);
nor U44865 (N_44865,N_41593,N_40412);
nand U44866 (N_44866,N_41976,N_41230);
nand U44867 (N_44867,N_42462,N_41237);
nand U44868 (N_44868,N_42431,N_42011);
and U44869 (N_44869,N_40320,N_42165);
nand U44870 (N_44870,N_41181,N_40191);
nand U44871 (N_44871,N_40291,N_41584);
nand U44872 (N_44872,N_41953,N_41770);
nor U44873 (N_44873,N_40483,N_41408);
and U44874 (N_44874,N_42007,N_42003);
or U44875 (N_44875,N_40122,N_40662);
nand U44876 (N_44876,N_40007,N_40857);
nand U44877 (N_44877,N_41230,N_40893);
nand U44878 (N_44878,N_42068,N_41710);
nor U44879 (N_44879,N_40858,N_40399);
xnor U44880 (N_44880,N_41050,N_40631);
nor U44881 (N_44881,N_40139,N_42231);
nand U44882 (N_44882,N_40670,N_40875);
or U44883 (N_44883,N_40636,N_41537);
or U44884 (N_44884,N_40196,N_41211);
and U44885 (N_44885,N_40788,N_41560);
nand U44886 (N_44886,N_41241,N_40338);
nand U44887 (N_44887,N_41507,N_40054);
and U44888 (N_44888,N_40976,N_41474);
nor U44889 (N_44889,N_41835,N_40644);
and U44890 (N_44890,N_40170,N_41177);
xor U44891 (N_44891,N_41671,N_42043);
and U44892 (N_44892,N_42374,N_41737);
or U44893 (N_44893,N_40827,N_40451);
xor U44894 (N_44894,N_40516,N_41910);
or U44895 (N_44895,N_42230,N_41535);
and U44896 (N_44896,N_40537,N_40128);
nor U44897 (N_44897,N_41115,N_40726);
nand U44898 (N_44898,N_41183,N_41022);
and U44899 (N_44899,N_42461,N_41925);
or U44900 (N_44900,N_42331,N_40045);
nor U44901 (N_44901,N_40379,N_41099);
and U44902 (N_44902,N_41174,N_41433);
nand U44903 (N_44903,N_41008,N_40496);
or U44904 (N_44904,N_40426,N_42447);
nor U44905 (N_44905,N_40194,N_42196);
or U44906 (N_44906,N_41750,N_41990);
xnor U44907 (N_44907,N_41786,N_40536);
nand U44908 (N_44908,N_40915,N_42389);
xor U44909 (N_44909,N_42484,N_40255);
xor U44910 (N_44910,N_40975,N_41000);
nor U44911 (N_44911,N_40063,N_41297);
nand U44912 (N_44912,N_41518,N_40223);
and U44913 (N_44913,N_40854,N_40939);
and U44914 (N_44914,N_41304,N_41736);
nor U44915 (N_44915,N_41281,N_40781);
nor U44916 (N_44916,N_42391,N_42373);
xor U44917 (N_44917,N_41562,N_41414);
and U44918 (N_44918,N_42317,N_42036);
nand U44919 (N_44919,N_41880,N_42079);
nand U44920 (N_44920,N_41586,N_40040);
or U44921 (N_44921,N_40363,N_42072);
nor U44922 (N_44922,N_41704,N_42109);
nand U44923 (N_44923,N_41006,N_41963);
and U44924 (N_44924,N_42104,N_40291);
and U44925 (N_44925,N_41917,N_40763);
or U44926 (N_44926,N_40406,N_40590);
nand U44927 (N_44927,N_40619,N_40478);
or U44928 (N_44928,N_40487,N_41656);
nor U44929 (N_44929,N_41330,N_40284);
or U44930 (N_44930,N_41100,N_41667);
or U44931 (N_44931,N_40155,N_41846);
nand U44932 (N_44932,N_40723,N_41123);
nand U44933 (N_44933,N_40932,N_40849);
and U44934 (N_44934,N_41136,N_40632);
and U44935 (N_44935,N_41551,N_42314);
and U44936 (N_44936,N_40093,N_42169);
xor U44937 (N_44937,N_40989,N_41043);
or U44938 (N_44938,N_41481,N_42117);
nand U44939 (N_44939,N_40585,N_40476);
and U44940 (N_44940,N_40263,N_42473);
xnor U44941 (N_44941,N_40336,N_41332);
and U44942 (N_44942,N_41818,N_41650);
and U44943 (N_44943,N_40057,N_41033);
or U44944 (N_44944,N_42260,N_41905);
or U44945 (N_44945,N_40365,N_41910);
and U44946 (N_44946,N_40024,N_42223);
nor U44947 (N_44947,N_41224,N_40280);
or U44948 (N_44948,N_40644,N_42426);
or U44949 (N_44949,N_42466,N_40325);
nor U44950 (N_44950,N_40256,N_40316);
nand U44951 (N_44951,N_41922,N_40696);
nand U44952 (N_44952,N_42178,N_40015);
xnor U44953 (N_44953,N_40239,N_40570);
xnor U44954 (N_44954,N_40870,N_42176);
nor U44955 (N_44955,N_41834,N_41949);
or U44956 (N_44956,N_40008,N_40038);
nand U44957 (N_44957,N_40362,N_40059);
or U44958 (N_44958,N_41783,N_40931);
nor U44959 (N_44959,N_42384,N_41478);
nor U44960 (N_44960,N_41484,N_40670);
nor U44961 (N_44961,N_41322,N_42423);
nor U44962 (N_44962,N_41744,N_41118);
nor U44963 (N_44963,N_42247,N_42134);
or U44964 (N_44964,N_41523,N_41243);
nor U44965 (N_44965,N_40607,N_41198);
nor U44966 (N_44966,N_40158,N_40511);
nand U44967 (N_44967,N_41375,N_40873);
and U44968 (N_44968,N_40769,N_40846);
nand U44969 (N_44969,N_41922,N_40044);
xnor U44970 (N_44970,N_42342,N_40051);
or U44971 (N_44971,N_40921,N_40301);
and U44972 (N_44972,N_40104,N_42037);
and U44973 (N_44973,N_42305,N_40310);
and U44974 (N_44974,N_42043,N_40905);
nand U44975 (N_44975,N_41443,N_40637);
and U44976 (N_44976,N_41227,N_40847);
nor U44977 (N_44977,N_40536,N_40027);
nand U44978 (N_44978,N_42084,N_41498);
xor U44979 (N_44979,N_41466,N_41637);
and U44980 (N_44980,N_40240,N_40721);
xor U44981 (N_44981,N_40323,N_40341);
and U44982 (N_44982,N_41151,N_41985);
and U44983 (N_44983,N_40722,N_40192);
or U44984 (N_44984,N_41118,N_41212);
or U44985 (N_44985,N_40558,N_41039);
nor U44986 (N_44986,N_40909,N_41787);
or U44987 (N_44987,N_40843,N_40329);
nor U44988 (N_44988,N_42027,N_40958);
and U44989 (N_44989,N_41528,N_40860);
xnor U44990 (N_44990,N_40050,N_41343);
nor U44991 (N_44991,N_40120,N_41810);
xnor U44992 (N_44992,N_41393,N_42163);
xnor U44993 (N_44993,N_40608,N_40433);
and U44994 (N_44994,N_40783,N_42478);
xnor U44995 (N_44995,N_40325,N_40652);
nor U44996 (N_44996,N_40378,N_41142);
nor U44997 (N_44997,N_40390,N_42285);
and U44998 (N_44998,N_42083,N_42154);
nor U44999 (N_44999,N_40634,N_42396);
nand U45000 (N_45000,N_43267,N_44390);
nor U45001 (N_45001,N_44895,N_44146);
or U45002 (N_45002,N_42777,N_42580);
or U45003 (N_45003,N_43220,N_43589);
or U45004 (N_45004,N_43065,N_43173);
nand U45005 (N_45005,N_43757,N_42752);
and U45006 (N_45006,N_42677,N_43855);
nor U45007 (N_45007,N_43043,N_44856);
nor U45008 (N_45008,N_44134,N_44731);
nand U45009 (N_45009,N_44641,N_42874);
nor U45010 (N_45010,N_43133,N_42693);
or U45011 (N_45011,N_43416,N_44019);
xnor U45012 (N_45012,N_44168,N_44876);
and U45013 (N_45013,N_43633,N_44688);
nor U45014 (N_45014,N_42707,N_42720);
xnor U45015 (N_45015,N_44115,N_42996);
nor U45016 (N_45016,N_42814,N_44837);
nor U45017 (N_45017,N_43901,N_42891);
or U45018 (N_45018,N_44334,N_42632);
and U45019 (N_45019,N_43675,N_44872);
nand U45020 (N_45020,N_43816,N_44260);
or U45021 (N_45021,N_42856,N_42786);
nor U45022 (N_45022,N_43139,N_43257);
nor U45023 (N_45023,N_43376,N_42736);
nand U45024 (N_45024,N_44703,N_44306);
nor U45025 (N_45025,N_43134,N_44016);
nand U45026 (N_45026,N_42916,N_43539);
or U45027 (N_45027,N_44196,N_44279);
nand U45028 (N_45028,N_43618,N_44912);
nand U45029 (N_45029,N_44112,N_42972);
or U45030 (N_45030,N_43374,N_42966);
nand U45031 (N_45031,N_42672,N_44948);
xor U45032 (N_45032,N_43559,N_44014);
or U45033 (N_45033,N_44583,N_44282);
or U45034 (N_45034,N_42836,N_43081);
xnor U45035 (N_45035,N_44650,N_42689);
xnor U45036 (N_45036,N_43676,N_43491);
or U45037 (N_45037,N_44612,N_43393);
nor U45038 (N_45038,N_44163,N_44157);
nand U45039 (N_45039,N_44861,N_43206);
xor U45040 (N_45040,N_43907,N_44581);
nor U45041 (N_45041,N_44240,N_44800);
nor U45042 (N_45042,N_44568,N_44771);
or U45043 (N_45043,N_44429,N_44342);
nor U45044 (N_45044,N_44122,N_44313);
xnor U45045 (N_45045,N_43403,N_44721);
xor U45046 (N_45046,N_44285,N_43836);
xnor U45047 (N_45047,N_44497,N_43044);
nor U45048 (N_45048,N_42760,N_42505);
nor U45049 (N_45049,N_44551,N_44414);
and U45050 (N_45050,N_42607,N_42539);
or U45051 (N_45051,N_43874,N_44391);
and U45052 (N_45052,N_43946,N_44759);
or U45053 (N_45053,N_43011,N_42556);
nor U45054 (N_45054,N_44471,N_43256);
nand U45055 (N_45055,N_44576,N_42549);
nand U45056 (N_45056,N_43643,N_42821);
nor U45057 (N_45057,N_44076,N_42599);
and U45058 (N_45058,N_44715,N_43606);
xnor U45059 (N_45059,N_44673,N_42567);
and U45060 (N_45060,N_42535,N_43292);
or U45061 (N_45061,N_42763,N_43725);
nand U45062 (N_45062,N_44248,N_44617);
nor U45063 (N_45063,N_42721,N_42560);
nor U45064 (N_45064,N_44258,N_44781);
nand U45065 (N_45065,N_44807,N_43387);
xor U45066 (N_45066,N_43818,N_44954);
and U45067 (N_45067,N_44220,N_43208);
nor U45068 (N_45068,N_44243,N_43506);
nand U45069 (N_45069,N_43165,N_44758);
and U45070 (N_45070,N_43467,N_44847);
or U45071 (N_45071,N_44147,N_42762);
nor U45072 (N_45072,N_43736,N_44442);
and U45073 (N_45073,N_44035,N_44998);
or U45074 (N_45074,N_44030,N_44364);
xor U45075 (N_45075,N_44064,N_44000);
or U45076 (N_45076,N_43557,N_44791);
xnor U45077 (N_45077,N_43939,N_43678);
and U45078 (N_45078,N_42524,N_44742);
and U45079 (N_45079,N_44644,N_43898);
nand U45080 (N_45080,N_44448,N_43113);
and U45081 (N_45081,N_42719,N_42923);
nand U45082 (N_45082,N_44244,N_42661);
nand U45083 (N_45083,N_44303,N_42589);
nor U45084 (N_45084,N_44133,N_43471);
nor U45085 (N_45085,N_44158,N_44107);
and U45086 (N_45086,N_44149,N_42783);
and U45087 (N_45087,N_44445,N_42812);
nand U45088 (N_45088,N_44614,N_44606);
or U45089 (N_45089,N_44377,N_43435);
xnor U45090 (N_45090,N_43096,N_42603);
xnor U45091 (N_45091,N_44859,N_43789);
nand U45092 (N_45092,N_44275,N_43771);
and U45093 (N_45093,N_44036,N_43249);
xor U45094 (N_45094,N_42994,N_44054);
nor U45095 (N_45095,N_44074,N_44379);
or U45096 (N_45096,N_43042,N_42676);
and U45097 (N_45097,N_43446,N_43852);
and U45098 (N_45098,N_42899,N_43753);
and U45099 (N_45099,N_43677,N_42973);
xor U45100 (N_45100,N_44607,N_44485);
xnor U45101 (N_45101,N_42900,N_44679);
nor U45102 (N_45102,N_44969,N_43494);
or U45103 (N_45103,N_43285,N_43866);
nor U45104 (N_45104,N_43703,N_43190);
nand U45105 (N_45105,N_44575,N_44534);
nor U45106 (N_45106,N_44402,N_42657);
and U45107 (N_45107,N_43910,N_44215);
xor U45108 (N_45108,N_44593,N_44462);
or U45109 (N_45109,N_43649,N_43031);
nand U45110 (N_45110,N_43335,N_43086);
nand U45111 (N_45111,N_42835,N_44329);
and U45112 (N_45112,N_42564,N_44660);
nor U45113 (N_45113,N_42879,N_43068);
or U45114 (N_45114,N_43670,N_43560);
nand U45115 (N_45115,N_42638,N_44709);
and U45116 (N_45116,N_43992,N_43873);
nand U45117 (N_45117,N_44870,N_43452);
or U45118 (N_45118,N_42546,N_43246);
and U45119 (N_45119,N_44068,N_43429);
nand U45120 (N_45120,N_42526,N_44531);
or U45121 (N_45121,N_43895,N_43905);
nor U45122 (N_45122,N_43973,N_43085);
nand U45123 (N_45123,N_42915,N_44691);
nor U45124 (N_45124,N_44528,N_42845);
nand U45125 (N_45125,N_42965,N_44853);
or U45126 (N_45126,N_44444,N_44530);
nand U45127 (N_45127,N_43639,N_44480);
nand U45128 (N_45128,N_42541,N_42969);
xnor U45129 (N_45129,N_43070,N_44836);
or U45130 (N_45130,N_44413,N_44857);
xor U45131 (N_45131,N_43401,N_43218);
and U45132 (N_45132,N_43706,N_43149);
nand U45133 (N_45133,N_44932,N_42788);
nand U45134 (N_45134,N_44230,N_43398);
nor U45135 (N_45135,N_44799,N_44986);
nand U45136 (N_45136,N_44381,N_43822);
or U45137 (N_45137,N_43323,N_42617);
and U45138 (N_45138,N_43769,N_43058);
nor U45139 (N_45139,N_43795,N_44592);
or U45140 (N_45140,N_43720,N_42794);
or U45141 (N_45141,N_44643,N_44401);
xnor U45142 (N_45142,N_44256,N_43164);
xor U45143 (N_45143,N_44967,N_43567);
and U45144 (N_45144,N_44852,N_42608);
and U45145 (N_45145,N_43749,N_43215);
and U45146 (N_45146,N_43313,N_44921);
nor U45147 (N_45147,N_42982,N_42862);
nand U45148 (N_45148,N_44945,N_43899);
xor U45149 (N_45149,N_43603,N_43610);
or U45150 (N_45150,N_43620,N_42967);
xor U45151 (N_45151,N_44189,N_44811);
nand U45152 (N_45152,N_43485,N_44142);
and U45153 (N_45153,N_44524,N_43558);
nand U45154 (N_45154,N_43271,N_42851);
and U45155 (N_45155,N_44116,N_43129);
xnor U45156 (N_45156,N_44446,N_43046);
and U45157 (N_45157,N_44063,N_44411);
xnor U45158 (N_45158,N_44616,N_43005);
nor U45159 (N_45159,N_42907,N_44489);
or U45160 (N_45160,N_42881,N_43858);
or U45161 (N_45161,N_43136,N_44177);
xnor U45162 (N_45162,N_43135,N_44558);
or U45163 (N_45163,N_43177,N_43951);
nand U45164 (N_45164,N_44667,N_44683);
nand U45165 (N_45165,N_43975,N_43646);
nand U45166 (N_45166,N_43409,N_42674);
or U45167 (N_45167,N_43977,N_43423);
nor U45168 (N_45168,N_43351,N_43631);
xor U45169 (N_45169,N_44522,N_43726);
or U45170 (N_45170,N_44152,N_44736);
xnor U45171 (N_45171,N_44977,N_42935);
nand U45172 (N_45172,N_43730,N_43959);
xnor U45173 (N_45173,N_43994,N_43247);
nand U45174 (N_45174,N_44357,N_44712);
xnor U45175 (N_45175,N_42515,N_44510);
xor U45176 (N_45176,N_44713,N_43648);
and U45177 (N_45177,N_43384,N_44624);
and U45178 (N_45178,N_43025,N_44653);
and U45179 (N_45179,N_43377,N_43463);
or U45180 (N_45180,N_44125,N_43709);
nand U45181 (N_45181,N_44761,N_44182);
xnor U45182 (N_45182,N_44015,N_44990);
nand U45183 (N_45183,N_42778,N_42850);
xor U45184 (N_45184,N_43550,N_43608);
xor U45185 (N_45185,N_43735,N_44487);
nand U45186 (N_45186,N_42948,N_44165);
and U45187 (N_45187,N_43521,N_43408);
xor U45188 (N_45188,N_44498,N_43651);
and U45189 (N_45189,N_44809,N_44674);
nor U45190 (N_45190,N_43492,N_43794);
nor U45191 (N_45191,N_43808,N_42548);
and U45192 (N_45192,N_43150,N_42998);
and U45193 (N_45193,N_43502,N_43138);
or U45194 (N_45194,N_44126,N_43094);
or U45195 (N_45195,N_42521,N_43157);
nor U45196 (N_45196,N_44959,N_42991);
or U45197 (N_45197,N_44473,N_42618);
or U45198 (N_45198,N_44976,N_42810);
nor U45199 (N_45199,N_42866,N_43829);
and U45200 (N_45200,N_44003,N_43418);
or U45201 (N_45201,N_43666,N_43536);
or U45202 (N_45202,N_44083,N_44717);
and U45203 (N_45203,N_44491,N_44785);
xnor U45204 (N_45204,N_43207,N_44113);
and U45205 (N_45205,N_43483,N_43211);
nor U45206 (N_45206,N_44832,N_42848);
or U45207 (N_45207,N_44788,N_43441);
nor U45208 (N_45208,N_42807,N_44287);
nand U45209 (N_45209,N_43981,N_43683);
nor U45210 (N_45210,N_44815,N_42680);
nand U45211 (N_45211,N_43188,N_42542);
nand U45212 (N_45212,N_43412,N_42550);
xor U45213 (N_45213,N_43200,N_44826);
nand U45214 (N_45214,N_43312,N_44419);
nor U45215 (N_45215,N_44621,N_43932);
and U45216 (N_45216,N_42612,N_44164);
nand U45217 (N_45217,N_43804,N_43275);
nand U45218 (N_45218,N_43996,N_43270);
and U45219 (N_45219,N_44052,N_42614);
or U45220 (N_45220,N_43698,N_43055);
xor U45221 (N_45221,N_43904,N_43186);
xnor U45222 (N_45222,N_43865,N_42928);
and U45223 (N_45223,N_43014,N_43518);
nor U45224 (N_45224,N_44369,N_42873);
nand U45225 (N_45225,N_43642,N_43078);
xor U45226 (N_45226,N_42748,N_42869);
xor U45227 (N_45227,N_44705,N_44700);
nor U45228 (N_45228,N_44347,N_44002);
nor U45229 (N_45229,N_42849,N_43367);
nor U45230 (N_45230,N_44632,N_43342);
xor U45231 (N_45231,N_43599,N_43655);
nor U45232 (N_45232,N_44151,N_44055);
or U45233 (N_45233,N_43128,N_43628);
and U45234 (N_45234,N_44298,N_44523);
nand U45235 (N_45235,N_44824,N_43303);
nand U45236 (N_45236,N_44246,N_44203);
nand U45237 (N_45237,N_42841,N_44192);
or U45238 (N_45238,N_43854,N_43219);
xnor U45239 (N_45239,N_42668,N_43445);
nor U45240 (N_45240,N_44565,N_43896);
xnor U45241 (N_45241,N_43308,N_44968);
xor U45242 (N_45242,N_43325,N_43686);
xor U45243 (N_45243,N_43847,N_43438);
and U45244 (N_45244,N_44034,N_44823);
nor U45245 (N_45245,N_42839,N_44216);
and U45246 (N_45246,N_43072,N_43688);
nand U45247 (N_45247,N_44596,N_43645);
and U45248 (N_45248,N_44507,N_43381);
and U45249 (N_45249,N_43925,N_43942);
nand U45250 (N_45250,N_42854,N_44816);
and U45251 (N_45251,N_44734,N_44629);
nor U45252 (N_45252,N_43891,N_43505);
nand U45253 (N_45253,N_43486,N_42805);
nand U45254 (N_45254,N_42895,N_43546);
xor U45255 (N_45255,N_43301,N_43613);
or U45256 (N_45256,N_44365,N_43034);
and U45257 (N_45257,N_42844,N_44097);
xnor U45258 (N_45258,N_43669,N_44431);
nand U45259 (N_45259,N_44383,N_43143);
xor U45260 (N_45260,N_43792,N_43080);
nand U45261 (N_45261,N_43974,N_43734);
nor U45262 (N_45262,N_42785,N_42690);
xnor U45263 (N_45263,N_44725,N_44255);
nand U45264 (N_45264,N_43913,N_44975);
nor U45265 (N_45265,N_43402,N_44562);
and U45266 (N_45266,N_44801,N_43033);
nor U45267 (N_45267,N_43050,N_44988);
xor U45268 (N_45268,N_44982,N_44748);
or U45269 (N_45269,N_43109,N_42519);
nor U45270 (N_45270,N_43641,N_42795);
nand U45271 (N_45271,N_43921,N_44337);
or U45272 (N_45272,N_43390,N_43363);
xor U45273 (N_45273,N_43021,N_43315);
and U45274 (N_45274,N_44393,N_43888);
nor U45275 (N_45275,N_42507,N_43812);
nand U45276 (N_45276,N_43878,N_44194);
nand U45277 (N_45277,N_43037,N_44994);
nand U45278 (N_45278,N_43653,N_43747);
or U45279 (N_45279,N_44218,N_42579);
nor U45280 (N_45280,N_43934,N_43316);
nand U45281 (N_45281,N_43075,N_43229);
or U45282 (N_45282,N_43537,N_44655);
or U45283 (N_45283,N_43002,N_42622);
nor U45284 (N_45284,N_44409,N_44407);
nand U45285 (N_45285,N_43579,N_43662);
or U45286 (N_45286,N_44185,N_43105);
nand U45287 (N_45287,N_42951,N_43580);
nand U45288 (N_45288,N_42909,N_44564);
and U45289 (N_45289,N_44041,N_44170);
xor U45290 (N_45290,N_44972,N_43272);
nor U45291 (N_45291,N_43941,N_42553);
and U45292 (N_45292,N_43815,N_44305);
nand U45293 (N_45293,N_44560,N_44187);
and U45294 (N_45294,N_43717,N_42582);
nand U45295 (N_45295,N_44790,N_44099);
or U45296 (N_45296,N_44868,N_44549);
or U45297 (N_45297,N_42766,N_44269);
or U45298 (N_45298,N_44040,N_44955);
nand U45299 (N_45299,N_44946,N_42683);
nand U45300 (N_45300,N_43671,N_44006);
xnor U45301 (N_45301,N_43879,N_44397);
xnor U45302 (N_45302,N_43543,N_44878);
xnor U45303 (N_45303,N_44659,N_42530);
and U45304 (N_45304,N_43029,N_42646);
nand U45305 (N_45305,N_43538,N_44710);
xor U45306 (N_45306,N_44301,N_44698);
nand U45307 (N_45307,N_43405,N_42974);
nand U45308 (N_45308,N_43533,N_44410);
and U45309 (N_45309,N_44367,N_44711);
nand U45310 (N_45310,N_43781,N_42757);
or U45311 (N_45311,N_43222,N_44290);
nor U45312 (N_45312,N_43837,N_42889);
nor U45313 (N_45313,N_44589,N_43496);
or U45314 (N_45314,N_43929,N_44027);
and U45315 (N_45315,N_43885,N_42734);
and U45316 (N_45316,N_42666,N_43772);
nand U45317 (N_45317,N_42738,N_44265);
or U45318 (N_45318,N_43382,N_42883);
nor U45319 (N_45319,N_43235,N_44766);
and U45320 (N_45320,N_44304,N_43245);
nor U45321 (N_45321,N_43013,N_43470);
nor U45322 (N_45322,N_42635,N_42824);
and U45323 (N_45323,N_42703,N_44741);
xor U45324 (N_45324,N_44153,N_44430);
nor U45325 (N_45325,N_43953,N_44834);
or U45326 (N_45326,N_43396,N_44864);
nor U45327 (N_45327,N_43371,N_42648);
xor U45328 (N_45328,N_42691,N_44274);
xor U45329 (N_45329,N_44095,N_42926);
or U45330 (N_45330,N_42919,N_43330);
xor U45331 (N_45331,N_43468,N_44077);
xor U45332 (N_45332,N_44682,N_43764);
nand U45333 (N_45333,N_42700,N_44375);
xnor U45334 (N_45334,N_44727,N_42739);
or U45335 (N_45335,N_44004,N_43227);
nand U45336 (N_45336,N_42876,N_44697);
and U45337 (N_45337,N_43444,N_43790);
xor U45338 (N_45338,N_44828,N_43180);
nand U45339 (N_45339,N_44420,N_44008);
and U45340 (N_45340,N_44166,N_43969);
xor U45341 (N_45341,N_43372,N_42508);
xnor U45342 (N_45342,N_44669,N_44845);
or U45343 (N_45343,N_44378,N_43741);
and U45344 (N_45344,N_43800,N_43447);
nor U45345 (N_45345,N_43540,N_43276);
nor U45346 (N_45346,N_43236,N_44831);
xor U45347 (N_45347,N_43568,N_44642);
nor U45348 (N_45348,N_43439,N_44900);
nor U45349 (N_45349,N_42586,N_44273);
nand U45350 (N_45350,N_44536,N_42569);
nand U45351 (N_45351,N_43225,N_44495);
or U45352 (N_45352,N_44706,N_43392);
nor U45353 (N_45353,N_43967,N_43161);
xnor U45354 (N_45354,N_44930,N_44582);
nor U45355 (N_45355,N_43430,N_43791);
xor U45356 (N_45356,N_43419,N_44208);
nand U45357 (N_45357,N_42981,N_44762);
xnor U45358 (N_45358,N_42660,N_42950);
or U45359 (N_45359,N_44931,N_44663);
and U45360 (N_45360,N_44841,N_43718);
nand U45361 (N_45361,N_42825,N_42831);
xnor U45362 (N_45362,N_44769,N_42826);
or U45363 (N_45363,N_43527,N_43581);
nand U45364 (N_45364,N_44056,N_44059);
and U45365 (N_45365,N_44898,N_44072);
nand U45366 (N_45366,N_43991,N_43489);
or U45367 (N_45367,N_42595,N_44757);
nand U45368 (N_45368,N_44694,N_43886);
nor U45369 (N_45369,N_43184,N_43120);
xor U45370 (N_45370,N_43615,N_43465);
or U45371 (N_45371,N_42894,N_43356);
nand U45372 (N_45372,N_44104,N_44965);
xor U45373 (N_45373,N_44093,N_43838);
nor U45374 (N_45374,N_42536,N_44752);
xnor U45375 (N_45375,N_42575,N_43525);
or U45376 (N_45376,N_44735,N_43743);
nand U45377 (N_45377,N_43722,N_44066);
and U45378 (N_45378,N_43509,N_44111);
and U45379 (N_45379,N_43748,N_42771);
nor U45380 (N_45380,N_44037,N_43048);
and U45381 (N_45381,N_44193,N_43348);
nor U45382 (N_45382,N_42692,N_42852);
nor U45383 (N_45383,N_42816,N_44225);
or U45384 (N_45384,N_43035,N_42888);
xor U45385 (N_45385,N_42540,N_44399);
xor U45386 (N_45386,N_44022,N_44251);
or U45387 (N_45387,N_42934,N_43010);
and U45388 (N_45388,N_44400,N_44594);
and U45389 (N_45389,N_43704,N_43949);
xor U45390 (N_45390,N_44840,N_43336);
nand U45391 (N_45391,N_43205,N_42872);
nor U45392 (N_45392,N_43876,N_44106);
xor U45393 (N_45393,N_43554,N_42609);
nand U45394 (N_45394,N_44120,N_44090);
xnor U45395 (N_45395,N_42598,N_44155);
or U45396 (N_45396,N_43768,N_43632);
or U45397 (N_45397,N_44045,N_43201);
nor U45398 (N_45398,N_44867,N_43425);
and U45399 (N_45399,N_43332,N_44174);
nor U45400 (N_45400,N_42616,N_42561);
and U45401 (N_45401,N_42711,N_43248);
nor U45402 (N_45402,N_43341,N_42625);
nand U45403 (N_45403,N_43146,N_43746);
or U45404 (N_45404,N_42903,N_44792);
and U45405 (N_45405,N_44910,N_42797);
nand U45406 (N_45406,N_42511,N_44050);
nand U45407 (N_45407,N_42741,N_43089);
xor U45408 (N_45408,N_44132,N_44359);
or U45409 (N_45409,N_43846,N_43663);
nor U45410 (N_45410,N_42545,N_43714);
or U45411 (N_45411,N_43260,N_44098);
or U45412 (N_45412,N_42959,N_44708);
nand U45413 (N_45413,N_42910,N_43493);
nor U45414 (N_45414,N_42784,N_42828);
and U45415 (N_45415,N_43118,N_44352);
nand U45416 (N_45416,N_43984,N_44386);
nand U45417 (N_45417,N_44283,N_44468);
and U45418 (N_45418,N_43345,N_42863);
nand U45419 (N_45419,N_42615,N_44728);
nor U45420 (N_45420,N_44351,N_44662);
and U45421 (N_45421,N_43616,N_44753);
and U45422 (N_45422,N_44069,N_42624);
or U45423 (N_45423,N_43880,N_43788);
and U45424 (N_45424,N_44176,N_43331);
nand U45425 (N_45425,N_43321,N_44395);
nor U45426 (N_45426,N_43450,N_43090);
xor U45427 (N_45427,N_44362,N_43240);
or U45428 (N_45428,N_44557,N_44681);
xnor U45429 (N_45429,N_43740,N_43782);
or U45430 (N_45430,N_44206,N_44904);
or U45431 (N_45431,N_44934,N_44724);
nand U45432 (N_45432,N_43024,N_43202);
nor U45433 (N_45433,N_44470,N_42551);
xor U45434 (N_45434,N_44129,N_43250);
nor U45435 (N_45435,N_44631,N_42995);
xnor U45436 (N_45436,N_44684,N_42525);
xnor U45437 (N_45437,N_42843,N_43487);
nor U45438 (N_45438,N_43993,N_42675);
xnor U45439 (N_45439,N_44270,N_43253);
or U45440 (N_45440,N_43867,N_42742);
nor U45441 (N_45441,N_43830,N_43673);
nand U45442 (N_45442,N_44983,N_44819);
xnor U45443 (N_45443,N_44906,N_44880);
nand U45444 (N_45444,N_44775,N_43428);
or U45445 (N_45445,N_43453,N_43827);
nor U45446 (N_45446,N_44490,N_43144);
xor U45447 (N_45447,N_44314,N_42892);
nand U45448 (N_45448,N_44084,N_43166);
nor U45449 (N_45449,N_42880,N_43813);
and U45450 (N_45450,N_42574,N_43665);
nor U45451 (N_45451,N_43712,N_42867);
nor U45452 (N_45452,N_43657,N_44587);
and U45453 (N_45453,N_43826,N_43414);
nor U45454 (N_45454,N_44875,N_42662);
nor U45455 (N_45455,N_44901,N_44324);
and U45456 (N_45456,N_44339,N_42699);
nor U45457 (N_45457,N_44981,N_43406);
xor U45458 (N_45458,N_44743,N_43971);
or U45459 (N_45459,N_42858,N_44529);
nor U45460 (N_45460,N_43775,N_43863);
and U45461 (N_45461,N_43379,N_43385);
nor U45462 (N_45462,N_44685,N_44570);
xnor U45463 (N_45463,N_43727,N_43987);
nand U45464 (N_45464,N_44926,N_44424);
xor U45465 (N_45465,N_42838,N_43158);
nor U45466 (N_45466,N_43283,N_44053);
or U45467 (N_45467,N_43810,N_42510);
and U45468 (N_45468,N_43756,N_42893);
nand U45469 (N_45469,N_42986,N_43451);
or U45470 (N_45470,N_42650,N_44695);
and U45471 (N_45471,N_42887,N_43914);
and U45472 (N_45472,N_44460,N_43373);
nor U45473 (N_45473,N_42952,N_42769);
nor U45474 (N_45474,N_43693,N_44382);
or U45475 (N_45475,N_42740,N_42767);
or U45476 (N_45476,N_44936,N_44545);
or U45477 (N_45477,N_44328,N_44902);
nand U45478 (N_45478,N_44227,N_42754);
nand U45479 (N_45479,N_44309,N_43897);
nor U45480 (N_45480,N_42663,N_43063);
and U45481 (N_45481,N_43306,N_44060);
and U45482 (N_45482,N_43498,N_43304);
or U45483 (N_45483,N_42604,N_43909);
xor U45484 (N_45484,N_43943,N_44426);
xor U45485 (N_45485,N_43586,N_43482);
nor U45486 (N_45486,N_44786,N_44408);
and U45487 (N_45487,N_44162,N_43023);
and U45488 (N_45488,N_44300,N_44319);
xor U45489 (N_45489,N_43347,N_42976);
nand U45490 (N_45490,N_43343,N_43059);
nand U45491 (N_45491,N_43243,N_44584);
nand U45492 (N_45492,N_44295,N_43397);
xnor U45493 (N_45493,N_42573,N_44547);
nand U45494 (N_45494,N_42988,N_44065);
nand U45495 (N_45495,N_43957,N_43716);
xor U45496 (N_45496,N_44101,N_44556);
nand U45497 (N_45497,N_43850,N_44481);
and U45498 (N_45498,N_44299,N_44597);
nor U45499 (N_45499,N_44951,N_43875);
nand U45500 (N_45500,N_43760,N_44810);
and U45501 (N_45501,N_44131,N_42949);
nor U45502 (N_45502,N_43298,N_44465);
and U45503 (N_45503,N_44289,N_44851);
or U45504 (N_45504,N_43983,N_42804);
nand U45505 (N_45505,N_42961,N_43127);
nor U45506 (N_45506,N_44281,N_44894);
or U45507 (N_45507,N_42792,N_43279);
and U45508 (N_45508,N_42694,N_42897);
nand U45509 (N_45509,N_44253,N_43112);
or U45510 (N_45510,N_44276,N_43322);
xor U45511 (N_45511,N_43064,N_44513);
nor U45512 (N_45512,N_44464,N_44200);
and U45513 (N_45513,N_44136,N_43831);
nor U45514 (N_45514,N_44086,N_44169);
or U45515 (N_45515,N_44009,N_43239);
nor U45516 (N_45516,N_44091,N_44353);
or U45517 (N_45517,N_44637,N_43226);
xor U45518 (N_45518,N_43707,N_44428);
or U45519 (N_45519,N_44096,N_42619);
and U45520 (N_45520,N_42842,N_44730);
nor U45521 (N_45521,N_43956,N_43307);
or U45522 (N_45522,N_44915,N_44860);
and U45523 (N_45523,N_43751,N_42640);
or U45524 (N_45524,N_42555,N_42558);
xor U45525 (N_45525,N_44922,N_42855);
nand U45526 (N_45526,N_44608,N_43295);
nor U45527 (N_45527,N_42822,N_44920);
xnor U45528 (N_45528,N_42941,N_43699);
xnor U45529 (N_45529,N_42823,N_44924);
and U45530 (N_45530,N_42906,N_44073);
and U45531 (N_45531,N_43629,N_44751);
or U45532 (N_45532,N_44666,N_43454);
and U45533 (N_45533,N_42702,N_44475);
nand U45534 (N_45534,N_44482,N_44923);
or U45535 (N_45535,N_43199,N_43114);
xor U45536 (N_45536,N_42502,N_44315);
or U45537 (N_45537,N_44574,N_43870);
and U45538 (N_45538,N_43597,N_44241);
nand U45539 (N_45539,N_44588,N_43051);
nor U45540 (N_45540,N_43151,N_44343);
or U45541 (N_45541,N_43488,N_44188);
xor U45542 (N_45542,N_43032,N_42633);
and U45543 (N_45543,N_43619,N_42724);
and U45544 (N_45544,N_42629,N_44813);
and U45545 (N_45545,N_44028,N_44718);
and U45546 (N_45546,N_43106,N_44925);
and U45547 (N_45547,N_43099,N_44331);
or U45548 (N_45548,N_44658,N_43674);
and U45549 (N_45549,N_43333,N_43366);
or U45550 (N_45550,N_44416,N_43012);
xor U45551 (N_45551,N_43765,N_43433);
and U45552 (N_45552,N_44999,N_44318);
and U45553 (N_45553,N_43668,N_44882);
xor U45554 (N_45554,N_42630,N_42588);
nand U45555 (N_45555,N_43162,N_43370);
nand U45556 (N_45556,N_43461,N_42591);
nor U45557 (N_45557,N_44021,N_43759);
xor U45558 (N_45558,N_42983,N_43713);
nor U45559 (N_45559,N_42653,N_44341);
nor U45560 (N_45560,N_44997,N_44294);
or U45561 (N_45561,N_43187,N_43600);
nor U45562 (N_45562,N_44380,N_43224);
or U45563 (N_45563,N_43966,N_43001);
and U45564 (N_45564,N_44388,N_44627);
xnor U45565 (N_45565,N_42912,N_43116);
nor U45566 (N_45566,N_43026,N_42776);
or U45567 (N_45567,N_42658,N_42673);
xor U45568 (N_45568,N_44171,N_43607);
nor U45569 (N_45569,N_43104,N_44159);
and U45570 (N_45570,N_43584,N_43833);
nand U45571 (N_45571,N_43998,N_43097);
xnor U45572 (N_45572,N_44360,N_43737);
nor U45573 (N_45573,N_42583,N_44432);
nand U45574 (N_45574,N_44963,N_44130);
and U45575 (N_45575,N_43448,N_43375);
nand U45576 (N_45576,N_43297,N_44467);
or U45577 (N_45577,N_44927,N_43284);
or U45578 (N_45578,N_43353,N_44443);
or U45579 (N_45579,N_43680,N_44696);
or U45580 (N_45580,N_42898,N_44372);
and U45581 (N_45581,N_44286,N_44437);
nand U45582 (N_45582,N_44061,N_43601);
and U45583 (N_45583,N_43659,N_44726);
or U45584 (N_45584,N_42682,N_44978);
and U45585 (N_45585,N_43352,N_43777);
xor U45586 (N_45586,N_44702,N_44846);
nand U45587 (N_45587,N_42726,N_42980);
and U45588 (N_45588,N_42947,N_44817);
and U45589 (N_45589,N_44238,N_43780);
and U45590 (N_45590,N_44494,N_43900);
nand U45591 (N_45591,N_43935,N_42678);
xnor U45592 (N_45592,N_43803,N_44228);
and U45593 (N_45593,N_43922,N_44292);
or U45594 (N_45594,N_43280,N_42523);
xnor U45595 (N_45595,N_43299,N_44863);
nand U45596 (N_45596,N_44418,N_44526);
nand U45597 (N_45597,N_44942,N_43009);
nand U45598 (N_45598,N_43582,N_44219);
nand U45599 (N_45599,N_43828,N_43516);
or U45600 (N_45600,N_44366,N_42749);
xor U45601 (N_45601,N_43528,N_42924);
and U45602 (N_45602,N_44474,N_44858);
xor U45603 (N_45603,N_43251,N_43621);
nor U45604 (N_45604,N_42764,N_44156);
or U45605 (N_45605,N_43049,N_42857);
xnor U45606 (N_45606,N_43930,N_43823);
or U45607 (N_45607,N_42781,N_43185);
and U45608 (N_45608,N_43413,N_43216);
xor U45609 (N_45609,N_43045,N_44778);
nor U45610 (N_45610,N_44051,N_44833);
nand U45611 (N_45611,N_44542,N_43920);
nand U45612 (N_45612,N_42775,N_42753);
nor U45613 (N_45613,N_43175,N_42637);
and U45614 (N_45614,N_43911,N_44609);
xnor U45615 (N_45615,N_43915,N_44918);
nor U45616 (N_45616,N_44889,N_42568);
and U45617 (N_45617,N_43918,N_44049);
nor U45618 (N_45618,N_44916,N_42819);
xnor U45619 (N_45619,N_44661,N_44719);
xnor U45620 (N_45620,N_42756,N_44770);
or U45621 (N_45621,N_43368,N_42623);
nand U45622 (N_45622,N_43122,N_44320);
nand U45623 (N_45623,N_43431,N_43801);
nor U45624 (N_45624,N_42529,N_44263);
nor U45625 (N_45625,N_44323,N_44532);
nor U45626 (N_45626,N_43857,N_43637);
xnor U45627 (N_45627,N_42606,N_43871);
xor U45628 (N_45628,N_44601,N_44940);
and U45629 (N_45629,N_44332,N_42620);
or U45630 (N_45630,N_43542,N_42723);
xnor U45631 (N_45631,N_43575,N_44223);
or U45632 (N_45632,N_43627,N_43480);
and U45633 (N_45633,N_42670,N_42847);
nand U45634 (N_45634,N_44423,N_44508);
and U45635 (N_45635,N_43176,N_43054);
and U45636 (N_45636,N_43711,N_43587);
xor U45637 (N_45637,N_44628,N_43681);
nor U45638 (N_45638,N_44843,N_43264);
and U45639 (N_45639,N_43721,N_44415);
nand U45640 (N_45640,N_43389,N_43750);
and U45641 (N_45641,N_44245,N_44484);
nor U45642 (N_45642,N_43574,N_44678);
and U45643 (N_45643,N_42868,N_44825);
or U45644 (N_45644,N_43098,N_43708);
nor U45645 (N_45645,N_42761,N_42937);
or U45646 (N_45646,N_42808,N_44615);
xnor U45647 (N_45647,N_43155,N_44505);
or U45648 (N_45648,N_43572,N_43061);
and U45649 (N_45649,N_42944,N_43501);
xnor U45650 (N_45650,N_42509,N_42718);
xor U45651 (N_45651,N_42708,N_43549);
xor U45652 (N_45652,N_43437,N_44939);
or U45653 (N_45653,N_44452,N_44029);
or U45654 (N_45654,N_44755,N_44457);
nor U45655 (N_45655,N_44079,N_43092);
xnor U45656 (N_45656,N_43209,N_43820);
or U45657 (N_45657,N_44236,N_43424);
and U45658 (N_45658,N_44361,N_43019);
nand U45659 (N_45659,N_43577,N_43523);
or U45660 (N_45660,N_42978,N_43917);
xnor U45661 (N_45661,N_42581,N_44435);
nand U45662 (N_45662,N_43872,N_44974);
nand U45663 (N_45663,N_43578,N_42522);
or U45664 (N_45664,N_43853,N_44085);
nor U45665 (N_45665,N_44199,N_43400);
xnor U45666 (N_45666,N_43924,N_44720);
and U45667 (N_45667,N_42576,N_44422);
nor U45668 (N_45668,N_42571,N_44602);
xnor U45669 (N_45669,N_42516,N_43689);
and U45670 (N_45670,N_43329,N_43883);
or U45671 (N_45671,N_43758,N_43961);
and U45672 (N_45672,N_44137,N_42533);
xor U45673 (N_45673,N_44088,N_42806);
nand U45674 (N_45674,N_43635,N_44124);
nor U45675 (N_45675,N_44183,N_43100);
nand U45676 (N_45676,N_44544,N_44865);
xnor U45677 (N_45677,N_44327,N_44818);
and U45678 (N_45678,N_44849,N_43228);
nor U45679 (N_45679,N_43369,N_43626);
nor U45680 (N_45680,N_43544,N_42716);
nand U45681 (N_45681,N_44403,N_43281);
or U45682 (N_45682,N_43310,N_43602);
nand U45683 (N_45683,N_44572,N_44405);
xnor U45684 (N_45684,N_43989,N_42886);
nand U45685 (N_45685,N_44191,N_43142);
xor U45686 (N_45686,N_42600,N_44071);
nand U45687 (N_45687,N_42939,N_44555);
and U45688 (N_45688,N_43232,N_43479);
xnor U45689 (N_45689,N_42593,N_43233);
xnor U45690 (N_45690,N_44321,N_44058);
nor U45691 (N_45691,N_43179,N_43842);
nor U45692 (N_45692,N_44802,N_42728);
xnor U45693 (N_45693,N_43687,N_43466);
xor U45694 (N_45694,N_44783,N_43731);
nor U45695 (N_45695,N_42833,N_44732);
nor U45696 (N_45696,N_43300,N_44550);
nor U45697 (N_45697,N_43576,N_44310);
and U45698 (N_45698,N_44648,N_43504);
xor U45699 (N_45699,N_42904,N_44805);
nor U45700 (N_45700,N_43779,N_43805);
xor U45701 (N_45701,N_44440,N_44119);
and U45702 (N_45702,N_43507,N_43819);
xor U45703 (N_45703,N_44344,N_43126);
and U45704 (N_45704,N_43359,N_43860);
xnor U45705 (N_45705,N_44348,N_42840);
xor U45706 (N_45706,N_44374,N_43745);
nand U45707 (N_45707,N_42861,N_42501);
xor U45708 (N_45708,N_44787,N_44871);
nand U45709 (N_45709,N_44543,N_42931);
xnor U45710 (N_45710,N_42500,N_44259);
nor U45711 (N_45711,N_43115,N_44782);
nor U45712 (N_45712,N_43729,N_43057);
xnor U45713 (N_45713,N_44503,N_43340);
nand U45714 (N_45714,N_43178,N_42747);
nand U45715 (N_45715,N_44385,N_44814);
or U45716 (N_45716,N_43774,N_42911);
and U45717 (N_45717,N_43656,N_43592);
and U45718 (N_45718,N_43360,N_43903);
nor U45719 (N_45719,N_42735,N_43141);
or U45720 (N_45720,N_44447,N_43237);
and U45721 (N_45721,N_42587,N_42544);
and U45722 (N_45722,N_44676,N_42920);
nand U45723 (N_45723,N_42527,N_42554);
nor U45724 (N_45724,N_44161,N_44554);
or U45725 (N_45725,N_43358,N_44249);
and U45726 (N_45726,N_44100,N_44893);
or U45727 (N_45727,N_43378,N_43965);
or U45728 (N_45728,N_42989,N_44675);
nand U45729 (N_45729,N_44668,N_44862);
xnor U45730 (N_45730,N_43947,N_43391);
xnor U45731 (N_45731,N_43529,N_42811);
or U45732 (N_45732,N_44913,N_44567);
xnor U45733 (N_45733,N_44080,N_42954);
and U45734 (N_45734,N_43269,N_43562);
or U45735 (N_45735,N_44605,N_44559);
or U45736 (N_45736,N_44479,N_43334);
nor U45737 (N_45737,N_44025,N_43952);
and U45738 (N_45738,N_44277,N_43497);
xor U45739 (N_45739,N_42979,N_44349);
nand U45740 (N_45740,N_44883,N_44441);
xor U45741 (N_45741,N_44458,N_44140);
nand U45742 (N_45742,N_43317,N_43093);
xnor U45743 (N_45743,N_44167,N_44578);
and U45744 (N_45744,N_43624,N_43147);
nor U45745 (N_45745,N_44143,N_44221);
or U45746 (N_45746,N_43605,N_42987);
nand U45747 (N_45747,N_42933,N_43773);
nor U45748 (N_45748,N_43422,N_42922);
nand U45749 (N_45749,N_42577,N_42532);
nor U45750 (N_45750,N_44154,N_44763);
or U45751 (N_45751,N_42504,N_43761);
and U45752 (N_45752,N_44075,N_43062);
nand U45753 (N_45753,N_43710,N_43311);
nor U45754 (N_45754,N_44611,N_43131);
xor U45755 (N_45755,N_44226,N_44311);
xor U45756 (N_45756,N_44919,N_43754);
or U45757 (N_45757,N_44566,N_42780);
or U45758 (N_45758,N_44671,N_43654);
and U45759 (N_45759,N_44774,N_42557);
and U45760 (N_45760,N_44938,N_42731);
and U45761 (N_45761,N_44291,N_43427);
and U45762 (N_45762,N_43108,N_42789);
nor U45763 (N_45763,N_44242,N_44421);
xor U45764 (N_45764,N_44217,N_44754);
xnor U45765 (N_45765,N_44980,N_43436);
xor U45766 (N_45766,N_44350,N_43950);
and U45767 (N_45767,N_43927,N_43530);
nand U45768 (N_45768,N_44745,N_43887);
nor U45769 (N_45769,N_44042,N_43884);
nor U45770 (N_45770,N_44506,N_43547);
nand U45771 (N_45771,N_43630,N_44387);
xnor U45772 (N_45772,N_43111,N_44995);
and U45773 (N_45773,N_43154,N_43192);
xnor U45774 (N_45774,N_44336,N_44477);
and U45775 (N_45775,N_42528,N_42993);
and U45776 (N_45776,N_44881,N_43552);
and U45777 (N_45777,N_44363,N_44518);
or U45778 (N_45778,N_42611,N_44264);
nand U45779 (N_45779,N_44793,N_44297);
or U45780 (N_45780,N_44639,N_43474);
xor U45781 (N_45781,N_44569,N_44548);
xnor U45782 (N_45782,N_43210,N_43982);
xor U45783 (N_45783,N_43755,N_43835);
xor U45784 (N_45784,N_42665,N_43832);
and U45785 (N_45785,N_43928,N_43526);
or U45786 (N_45786,N_44603,N_44714);
and U45787 (N_45787,N_43354,N_42896);
nor U45788 (N_45788,N_44224,N_44376);
xnor U45789 (N_45789,N_42687,N_42563);
xor U45790 (N_45790,N_43556,N_43500);
nand U45791 (N_45791,N_43604,N_43591);
and U45792 (N_45792,N_44070,N_44960);
xor U45793 (N_45793,N_44947,N_44373);
and U45794 (N_45794,N_43986,N_44384);
nor U45795 (N_45795,N_42940,N_44011);
or U45796 (N_45796,N_42641,N_44123);
nand U45797 (N_45797,N_44231,N_43997);
nand U45798 (N_45798,N_44573,N_42503);
or U45799 (N_45799,N_43916,N_44953);
nand U45800 (N_45800,N_44267,N_43364);
xor U45801 (N_45801,N_43355,N_44501);
xnor U45802 (N_45802,N_43839,N_44322);
nand U45803 (N_45803,N_43339,N_42732);
nor U45804 (N_45804,N_42578,N_44517);
nand U45805 (N_45805,N_43636,N_43084);
and U45806 (N_45806,N_44272,N_43189);
or U45807 (N_45807,N_44184,N_44118);
or U45808 (N_45808,N_44454,N_44312);
nand U45809 (N_45809,N_43732,N_44463);
xnor U45810 (N_45810,N_43573,N_44907);
and U45811 (N_45811,N_42713,N_43357);
or U45812 (N_45812,N_43609,N_44830);
nor U45813 (N_45813,N_43864,N_43395);
and U45814 (N_45814,N_43383,N_44389);
or U45815 (N_45815,N_43785,N_43596);
or U45816 (N_45816,N_43796,N_42914);
nor U45817 (N_45817,N_44135,N_42644);
nand U45818 (N_45818,N_43767,N_44406);
xnor U45819 (N_45819,N_43410,N_42729);
and U45820 (N_45820,N_42943,N_43622);
xor U45821 (N_45821,N_43475,N_42793);
and U45822 (N_45822,N_44527,N_42930);
or U45823 (N_45823,N_43570,N_43697);
xnor U45824 (N_45824,N_43752,N_43933);
nand U45825 (N_45825,N_44110,N_44469);
xnor U45826 (N_45826,N_43148,N_43963);
or U45827 (N_45827,N_44909,N_43893);
nand U45828 (N_45828,N_43945,N_44024);
nand U45829 (N_45829,N_44190,N_42813);
nand U45830 (N_45830,N_44738,N_43263);
and U45831 (N_45831,N_44222,N_44117);
and U45832 (N_45832,N_44618,N_44252);
nor U45833 (N_45833,N_44486,N_44427);
nor U45834 (N_45834,N_42513,N_43856);
and U45835 (N_45835,N_44877,N_42779);
and U45836 (N_45836,N_43107,N_43862);
nand U45837 (N_45837,N_44873,N_44739);
nand U45838 (N_45838,N_42559,N_43784);
nand U45839 (N_45839,N_43503,N_44103);
nand U45840 (N_45840,N_43117,N_42706);
or U45841 (N_45841,N_42877,N_44636);
and U45842 (N_45842,N_43923,N_43380);
nand U45843 (N_45843,N_43937,N_43617);
nor U45844 (N_45844,N_42562,N_42590);
nor U45845 (N_45845,N_43365,N_44496);
nand U45846 (N_45846,N_44317,N_43261);
or U45847 (N_45847,N_43399,N_43744);
and U45848 (N_45848,N_43585,N_44590);
or U45849 (N_45849,N_43970,N_44392);
nor U45850 (N_45850,N_42758,N_44483);
or U45851 (N_45851,N_43223,N_44509);
nand U45852 (N_45852,N_42964,N_43534);
nor U45853 (N_45853,N_44018,N_42697);
or U45854 (N_45854,N_42686,N_44180);
nand U45855 (N_45855,N_44640,N_42927);
and U45856 (N_45856,N_43459,N_42534);
nor U45857 (N_45857,N_42715,N_43724);
nor U45858 (N_45858,N_43309,N_43183);
nand U45859 (N_45859,N_44887,N_44173);
or U45860 (N_45860,N_43481,N_43564);
nand U45861 (N_45861,N_44234,N_44635);
nor U45862 (N_45862,N_42992,N_43571);
nand U45863 (N_45863,N_43244,N_44266);
nor U45864 (N_45864,N_43912,N_44201);
nand U45865 (N_45865,N_42975,N_43770);
nand U45866 (N_45866,N_44519,N_43985);
or U45867 (N_45867,N_44345,N_43834);
nand U45868 (N_45868,N_44330,N_43869);
nor U45869 (N_45869,N_43197,N_43881);
nor U45870 (N_45870,N_44211,N_44520);
nand U45871 (N_45871,N_44057,N_44512);
nand U45872 (N_45872,N_43066,N_44827);
or U45873 (N_45873,N_44233,N_44911);
nor U45874 (N_45874,N_44620,N_43962);
nor U45875 (N_45875,N_44746,N_44005);
or U45876 (N_45876,N_42759,N_44108);
xnor U45877 (N_45877,N_44195,N_43349);
and U45878 (N_45878,N_42832,N_43007);
and U45879 (N_45879,N_44677,N_43036);
or U45880 (N_45880,N_44806,N_42932);
and U45881 (N_45881,N_43404,N_43230);
and U45882 (N_45882,N_44533,N_44472);
and U45883 (N_45883,N_44439,N_43460);
xnor U45884 (N_45884,N_42621,N_44869);
nand U45885 (N_45885,N_44687,N_43259);
nand U45886 (N_45886,N_42518,N_42584);
nand U45887 (N_45887,N_44729,N_44262);
or U45888 (N_45888,N_43289,N_43612);
nand U45889 (N_45889,N_43193,N_44355);
or U45890 (N_45890,N_42696,N_44941);
or U45891 (N_45891,N_43968,N_43783);
nand U45892 (N_45892,N_44598,N_43195);
nand U45893 (N_45893,N_43473,N_42870);
nand U45894 (N_45894,N_43337,N_42860);
or U45895 (N_45895,N_42565,N_42714);
and U45896 (N_45896,N_42865,N_43041);
or U45897 (N_45897,N_44723,N_43194);
nand U45898 (N_45898,N_42538,N_44500);
or U45899 (N_45899,N_44139,N_43456);
xnor U45900 (N_45900,N_44855,N_44914);
and U45901 (N_45901,N_43458,N_44672);
and U45902 (N_45902,N_44899,N_42594);
nor U45903 (N_45903,N_43514,N_44820);
nand U45904 (N_45904,N_42514,N_44772);
xnor U45905 (N_45905,N_43902,N_44121);
nor U45906 (N_45906,N_43477,N_43938);
or U45907 (N_45907,N_44933,N_42963);
xor U45908 (N_45908,N_43182,N_43843);
nand U45909 (N_45909,N_43802,N_42871);
and U45910 (N_45910,N_42750,N_42730);
nor U45911 (N_45911,N_42709,N_42570);
or U45912 (N_45912,N_43825,N_43594);
and U45913 (N_45913,N_44949,N_44094);
nor U45914 (N_45914,N_43238,N_44067);
xnor U45915 (N_45915,N_44571,N_44247);
or U45916 (N_45916,N_43119,N_44504);
or U45917 (N_45917,N_44979,N_43326);
xnor U45918 (N_45918,N_44798,N_42506);
or U45919 (N_45919,N_43255,N_43407);
nor U45920 (N_45920,N_42751,N_44048);
nand U45921 (N_45921,N_43053,N_42566);
nor U45922 (N_45922,N_44645,N_42971);
nor U45923 (N_45923,N_43590,N_42809);
or U45924 (N_45924,N_42787,N_43723);
and U45925 (N_45925,N_44204,N_42875);
and U45926 (N_45926,N_43361,N_44261);
and U45927 (N_45927,N_43478,N_43140);
nand U45928 (N_45928,N_42917,N_43840);
or U45929 (N_45929,N_43644,N_44625);
and U45930 (N_45930,N_43972,N_44577);
and U45931 (N_45931,N_44789,N_42655);
nand U45932 (N_45932,N_44412,N_44210);
and U45933 (N_45933,N_44214,N_44579);
and U45934 (N_45934,N_43082,N_44488);
and U45935 (N_45935,N_43440,N_44396);
or U45936 (N_45936,N_44046,N_43069);
xor U45937 (N_45937,N_44750,N_44693);
xor U45938 (N_45938,N_43027,N_43168);
xnor U45939 (N_45939,N_42743,N_44935);
nand U45940 (N_45940,N_44586,N_44356);
nor U45941 (N_45941,N_44623,N_44760);
or U45942 (N_45942,N_43700,N_43715);
and U45943 (N_45943,N_42746,N_44956);
or U45944 (N_45944,N_43958,N_44768);
nand U45945 (N_45945,N_43017,N_44128);
and U45946 (N_45946,N_43350,N_44613);
xor U45947 (N_45947,N_43787,N_42652);
xor U45948 (N_45948,N_42669,N_43845);
nor U45949 (N_45949,N_44250,N_43565);
nor U45950 (N_45950,N_43520,N_42613);
nor U45951 (N_45951,N_43469,N_44854);
nor U45952 (N_45952,N_43672,N_42936);
nor U45953 (N_45953,N_44561,N_44160);
and U45954 (N_45954,N_44404,N_44952);
or U45955 (N_45955,N_42547,N_43510);
nand U45956 (N_45956,N_42733,N_43277);
xor U45957 (N_45957,N_43944,N_42643);
nor U45958 (N_45958,N_42651,N_42955);
nor U45959 (N_45959,N_42654,N_42717);
nand U45960 (N_45960,N_42945,N_43095);
nor U45961 (N_45961,N_43661,N_43018);
nor U45962 (N_45962,N_44141,N_44716);
xnor U45963 (N_45963,N_43338,N_44459);
nand U45964 (N_45964,N_44943,N_44538);
and U45965 (N_45965,N_43692,N_42790);
xnor U45966 (N_45966,N_44007,N_43074);
xnor U45967 (N_45967,N_44175,N_43524);
xnor U45968 (N_45968,N_42517,N_44371);
xnor U45969 (N_45969,N_44649,N_44476);
or U45970 (N_45970,N_44229,N_42765);
nor U45971 (N_45971,N_44232,N_42782);
nand U45972 (N_45972,N_42925,N_43472);
xnor U45973 (N_45973,N_44634,N_44144);
or U45974 (N_45974,N_43464,N_43006);
nor U45975 (N_45975,N_42631,N_42885);
nand U45976 (N_45976,N_44619,N_42681);
nand U45977 (N_45977,N_43940,N_43015);
nand U45978 (N_45978,N_43978,N_42800);
nand U45979 (N_45979,N_43797,N_44425);
xnor U45980 (N_45980,N_42796,N_42890);
nor U45981 (N_45981,N_42921,N_43305);
nor U45982 (N_45982,N_42942,N_43442);
nor U45983 (N_45983,N_43102,N_44235);
nand U45984 (N_45984,N_44316,N_43926);
xnor U45985 (N_45985,N_42878,N_43052);
and U45986 (N_45986,N_43290,N_44178);
and U45987 (N_45987,N_43719,N_43214);
and U45988 (N_45988,N_43763,N_44047);
and U45989 (N_45989,N_42602,N_43809);
nor U45990 (N_45990,N_44012,N_43125);
xor U45991 (N_45991,N_44511,N_43156);
and U45992 (N_45992,N_42627,N_43696);
nand U45993 (N_45993,N_44089,N_42704);
and U45994 (N_45994,N_44205,N_43844);
nor U45995 (N_45995,N_44885,N_44822);
nand U45996 (N_45996,N_43807,N_43174);
nor U45997 (N_45997,N_44984,N_44656);
nand U45998 (N_45998,N_43705,N_44449);
nor U45999 (N_45999,N_44450,N_43682);
and U46000 (N_46000,N_44664,N_43328);
and U46001 (N_46001,N_42605,N_43088);
xnor U46002 (N_46002,N_44903,N_44127);
xnor U46003 (N_46003,N_44541,N_44202);
or U46004 (N_46004,N_43171,N_42791);
nor U46005 (N_46005,N_42901,N_42829);
nor U46006 (N_46006,N_44087,N_43667);
nand U46007 (N_46007,N_43067,N_43091);
nand U46008 (N_46008,N_44652,N_43955);
nand U46009 (N_46009,N_43541,N_43160);
nand U46010 (N_46010,N_44989,N_43434);
or U46011 (N_46011,N_43060,N_44017);
or U46012 (N_46012,N_43611,N_44552);
and U46013 (N_46013,N_43462,N_43212);
or U46014 (N_46014,N_44928,N_42520);
xor U46015 (N_46015,N_43495,N_43995);
and U46016 (N_46016,N_44929,N_44808);
xor U46017 (N_46017,N_43979,N_42929);
nand U46018 (N_46018,N_43999,N_43004);
nor U46019 (N_46019,N_43694,N_43522);
xnor U46020 (N_46020,N_44749,N_43519);
and U46021 (N_46021,N_42712,N_43124);
or U46022 (N_46022,N_44610,N_44773);
nand U46023 (N_46023,N_42671,N_44784);
xnor U46024 (N_46024,N_43101,N_44370);
nand U46025 (N_46025,N_42985,N_44257);
xor U46026 (N_46026,N_44102,N_43394);
nand U46027 (N_46027,N_43799,N_44804);
nor U46028 (N_46028,N_44780,N_42802);
xor U46029 (N_46029,N_44308,N_44340);
or U46030 (N_46030,N_44866,N_44670);
and U46031 (N_46031,N_44803,N_43455);
xor U46032 (N_46032,N_43548,N_43892);
nand U46033 (N_46033,N_43003,N_43213);
nand U46034 (N_46034,N_43861,N_43684);
xor U46035 (N_46035,N_43623,N_42905);
xnor U46036 (N_46036,N_43685,N_44690);
nor U46037 (N_46037,N_44213,N_44970);
nor U46038 (N_46038,N_42882,N_44993);
or U46039 (N_46039,N_43443,N_43152);
xnor U46040 (N_46040,N_43786,N_42902);
or U46041 (N_46041,N_43679,N_43172);
nor U46042 (N_46042,N_42774,N_43561);
and U46043 (N_46043,N_44971,N_43776);
and U46044 (N_46044,N_42610,N_44455);
nand U46045 (N_46045,N_43288,N_44039);
nand U46046 (N_46046,N_43964,N_42597);
xor U46047 (N_46047,N_44797,N_42938);
nor U46048 (N_46048,N_42628,N_43980);
or U46049 (N_46049,N_43638,N_44835);
nand U46050 (N_46050,N_44138,N_43327);
nand U46051 (N_46051,N_43868,N_44842);
and U46052 (N_46052,N_44850,N_44032);
xor U46053 (N_46053,N_42817,N_44535);
or U46054 (N_46054,N_44657,N_44737);
or U46055 (N_46055,N_42962,N_43889);
xnor U46056 (N_46056,N_44023,N_42837);
or U46057 (N_46057,N_44453,N_44239);
and U46058 (N_46058,N_43695,N_43739);
nor U46059 (N_46059,N_44987,N_43077);
or U46060 (N_46060,N_44964,N_44796);
nand U46061 (N_46061,N_44622,N_43513);
xnor U46062 (N_46062,N_44848,N_44451);
and U46063 (N_46063,N_43566,N_43386);
nand U46064 (N_46064,N_43512,N_44886);
and U46065 (N_46065,N_43103,N_44043);
or U46066 (N_46066,N_43159,N_44812);
and U46067 (N_46067,N_44338,N_44346);
and U46068 (N_46068,N_43508,N_44689);
xor U46069 (N_46069,N_43278,N_42667);
xor U46070 (N_46070,N_44417,N_43204);
nand U46071 (N_46071,N_43079,N_44433);
nand U46072 (N_46072,N_44996,N_44795);
nor U46073 (N_46073,N_43318,N_44209);
or U46074 (N_46074,N_43877,N_43728);
xor U46075 (N_46075,N_43319,N_44268);
and U46076 (N_46076,N_43532,N_43545);
or U46077 (N_46077,N_43563,N_43132);
xnor U46078 (N_46078,N_43936,N_42970);
nand U46079 (N_46079,N_42695,N_44908);
nor U46080 (N_46080,N_44280,N_42827);
nand U46081 (N_46081,N_42956,N_44692);
and U46082 (N_46082,N_44537,N_42685);
nor U46083 (N_46083,N_44747,N_44207);
nor U46084 (N_46084,N_42946,N_44026);
xnor U46085 (N_46085,N_43954,N_42799);
or U46086 (N_46086,N_44961,N_42626);
nor U46087 (N_46087,N_43071,N_44001);
nand U46088 (N_46088,N_43273,N_42585);
xnor U46089 (N_46089,N_42531,N_43421);
nor U46090 (N_46090,N_43762,N_43163);
xor U46091 (N_46091,N_44109,N_44699);
nor U46092 (N_46092,N_44539,N_43793);
or U46093 (N_46093,N_43814,N_43426);
and U46094 (N_46094,N_43988,N_43882);
nor U46095 (N_46095,N_44779,N_42634);
or U46096 (N_46096,N_44966,N_44434);
or U46097 (N_46097,N_43040,N_42818);
xnor U46098 (N_46098,N_44884,N_44992);
and U46099 (N_46099,N_43121,N_43030);
nand U46100 (N_46100,N_44368,N_43287);
nor U46101 (N_46101,N_44105,N_43056);
or U46102 (N_46102,N_42596,N_42884);
nand U46103 (N_46103,N_43008,N_42552);
and U46104 (N_46104,N_43595,N_43598);
nor U46105 (N_46105,N_44905,N_44680);
nand U46106 (N_46106,N_44212,N_44546);
nand U46107 (N_46107,N_43262,N_42913);
xor U46108 (N_46108,N_44563,N_44776);
and U46109 (N_46109,N_42834,N_44580);
or U46110 (N_46110,N_44150,N_44466);
or U46111 (N_46111,N_44540,N_44892);
nor U46112 (N_46112,N_44033,N_44917);
nor U46113 (N_46113,N_43948,N_44358);
nand U46114 (N_46114,N_44897,N_43859);
nor U46115 (N_46115,N_44296,N_42727);
and U46116 (N_46116,N_44765,N_44516);
nor U46117 (N_46117,N_43614,N_43555);
nor U46118 (N_46118,N_43821,N_44354);
or U46119 (N_46119,N_42592,N_43535);
nand U46120 (N_46120,N_44302,N_44092);
xnor U46121 (N_46121,N_42798,N_42957);
and U46122 (N_46122,N_44172,N_42656);
and U46123 (N_46123,N_44525,N_44740);
nand U46124 (N_46124,N_43733,N_44591);
or U46125 (N_46125,N_44879,N_44651);
xnor U46126 (N_46126,N_43742,N_44638);
nand U46127 (N_46127,N_43976,N_43449);
or U46128 (N_46128,N_44686,N_43266);
or U46129 (N_46129,N_42770,N_44515);
or U46130 (N_46130,N_44325,N_44985);
and U46131 (N_46131,N_43234,N_44284);
or U46132 (N_46132,N_43324,N_44962);
nor U46133 (N_46133,N_42647,N_43302);
xor U46134 (N_46134,N_44456,N_42977);
xnor U46135 (N_46135,N_44461,N_43181);
nor U46136 (N_46136,N_43242,N_43314);
nand U46137 (N_46137,N_44839,N_44478);
nor U46138 (N_46138,N_43231,N_42830);
nand U46139 (N_46139,N_42990,N_44794);
nand U46140 (N_46140,N_43960,N_42773);
nor U46141 (N_46141,N_43344,N_43531);
nor U46142 (N_46142,N_43388,N_44333);
and U46143 (N_46143,N_43221,N_42642);
xnor U46144 (N_46144,N_42543,N_43817);
and U46145 (N_46145,N_44733,N_43039);
and U46146 (N_46146,N_43417,N_43087);
nand U46147 (N_46147,N_44890,N_43217);
and U46148 (N_46148,N_43265,N_43241);
nand U46149 (N_46149,N_43990,N_42537);
nor U46150 (N_46150,N_44438,N_42803);
xnor U46151 (N_46151,N_44891,N_43286);
nand U46152 (N_46152,N_44307,N_42737);
nand U46153 (N_46153,N_43282,N_44647);
nand U46154 (N_46154,N_42997,N_42960);
or U46155 (N_46155,N_42801,N_43110);
nand U46156 (N_46156,N_43634,N_44973);
xor U46157 (N_46157,N_42999,N_43553);
nand U46158 (N_46158,N_43919,N_42645);
nand U46159 (N_46159,N_43511,N_44874);
nand U46160 (N_46160,N_44777,N_43268);
xnor U46161 (N_46161,N_43908,N_44896);
xor U46162 (N_46162,N_43457,N_43411);
nand U46163 (N_46163,N_44179,N_43476);
nor U46164 (N_46164,N_44398,N_43890);
xor U46165 (N_46165,N_43028,N_43650);
xor U46166 (N_46166,N_43849,N_43517);
nor U46167 (N_46167,N_44010,N_44704);
and U46168 (N_46168,N_44553,N_44633);
and U46169 (N_46169,N_44958,N_43848);
and U46170 (N_46170,N_44585,N_43691);
and U46171 (N_46171,N_43664,N_43198);
nor U46172 (N_46172,N_42684,N_44821);
nor U46173 (N_46173,N_44626,N_43130);
and U46174 (N_46174,N_44937,N_44020);
xor U46175 (N_46175,N_42722,N_43022);
nand U46176 (N_46176,N_44944,N_44829);
and U46177 (N_46177,N_44271,N_43047);
nand U46178 (N_46178,N_43083,N_43490);
xor U46179 (N_46179,N_43362,N_44148);
xnor U46180 (N_46180,N_43778,N_44888);
and U46181 (N_46181,N_44630,N_43346);
xnor U46182 (N_46182,N_43625,N_44646);
xnor U46183 (N_46183,N_43076,N_42701);
xor U46184 (N_46184,N_42636,N_44278);
or U46185 (N_46185,N_43252,N_44082);
and U46186 (N_46186,N_42725,N_42688);
or U46187 (N_46187,N_42953,N_42908);
nand U46188 (N_46188,N_43320,N_43515);
and U46189 (N_46189,N_44114,N_44838);
and U46190 (N_46190,N_43145,N_44493);
or U46191 (N_46191,N_44186,N_42512);
and U46192 (N_46192,N_44722,N_42710);
nor U46193 (N_46193,N_44767,N_44701);
nand U46194 (N_46194,N_44145,N_42664);
xor U46195 (N_46195,N_44081,N_44198);
and U46196 (N_46196,N_43274,N_42572);
and U46197 (N_46197,N_44031,N_44078);
nor U46198 (N_46198,N_44394,N_43766);
or U46199 (N_46199,N_42820,N_43203);
or U46200 (N_46200,N_42705,N_43073);
and U46201 (N_46201,N_43583,N_43811);
and U46202 (N_46202,N_43123,N_44197);
nand U46203 (N_46203,N_44038,N_43593);
nor U46204 (N_46204,N_43153,N_44600);
nor U46205 (N_46205,N_43551,N_43191);
nand U46206 (N_46206,N_43658,N_44950);
and U46207 (N_46207,N_42864,N_42859);
nor U46208 (N_46208,N_43906,N_43702);
nand U46209 (N_46209,N_42984,N_43931);
nand U46210 (N_46210,N_43020,N_43499);
nand U46211 (N_46211,N_44502,N_44764);
nor U46212 (N_46212,N_43894,N_44521);
xor U46213 (N_46213,N_43016,N_43806);
nand U46214 (N_46214,N_43167,N_42815);
nor U46215 (N_46215,N_42601,N_43170);
nand U46216 (N_46216,N_44599,N_42918);
nand U46217 (N_46217,N_44044,N_43824);
xnor U46218 (N_46218,N_44991,N_42772);
nor U46219 (N_46219,N_44335,N_43569);
and U46220 (N_46220,N_43254,N_42853);
nand U46221 (N_46221,N_43432,N_44744);
nor U46222 (N_46222,N_43038,N_43294);
and U46223 (N_46223,N_43588,N_44436);
and U46224 (N_46224,N_44237,N_43169);
xor U46225 (N_46225,N_44254,N_44665);
or U46226 (N_46226,N_43652,N_44654);
xor U46227 (N_46227,N_44492,N_44844);
nor U46228 (N_46228,N_44181,N_44514);
or U46229 (N_46229,N_42659,N_42968);
nor U46230 (N_46230,N_44604,N_42679);
nand U46231 (N_46231,N_44707,N_42698);
nand U46232 (N_46232,N_43420,N_42745);
nand U46233 (N_46233,N_43701,N_42639);
nor U46234 (N_46234,N_43660,N_42755);
nor U46235 (N_46235,N_44293,N_44326);
xnor U46236 (N_46236,N_43258,N_43640);
nand U46237 (N_46237,N_44288,N_42846);
nor U46238 (N_46238,N_43415,N_42744);
nand U46239 (N_46239,N_42649,N_44062);
or U46240 (N_46240,N_43851,N_43137);
nor U46241 (N_46241,N_43690,N_43484);
nand U46242 (N_46242,N_44499,N_43798);
nand U46243 (N_46243,N_43738,N_42958);
and U46244 (N_46244,N_43647,N_43196);
and U46245 (N_46245,N_44595,N_43291);
or U46246 (N_46246,N_43841,N_44013);
nor U46247 (N_46247,N_43000,N_43293);
xor U46248 (N_46248,N_43296,N_44957);
nor U46249 (N_46249,N_44756,N_42768);
nor U46250 (N_46250,N_44647,N_44856);
and U46251 (N_46251,N_44895,N_43362);
and U46252 (N_46252,N_43659,N_43356);
and U46253 (N_46253,N_44951,N_43231);
nor U46254 (N_46254,N_43348,N_43139);
or U46255 (N_46255,N_42620,N_44032);
nand U46256 (N_46256,N_43665,N_43193);
and U46257 (N_46257,N_42742,N_43523);
and U46258 (N_46258,N_44186,N_42949);
nor U46259 (N_46259,N_43309,N_44937);
or U46260 (N_46260,N_43981,N_43133);
or U46261 (N_46261,N_44424,N_44914);
or U46262 (N_46262,N_42619,N_44774);
nand U46263 (N_46263,N_44320,N_44902);
nand U46264 (N_46264,N_43883,N_43945);
nand U46265 (N_46265,N_43488,N_44443);
xnor U46266 (N_46266,N_44819,N_42939);
nor U46267 (N_46267,N_43334,N_44026);
xnor U46268 (N_46268,N_43353,N_42522);
and U46269 (N_46269,N_43573,N_44526);
xor U46270 (N_46270,N_43508,N_42897);
xor U46271 (N_46271,N_43180,N_43397);
or U46272 (N_46272,N_44211,N_43278);
and U46273 (N_46273,N_44609,N_43110);
and U46274 (N_46274,N_44438,N_42816);
or U46275 (N_46275,N_43197,N_43871);
or U46276 (N_46276,N_43124,N_44651);
xnor U46277 (N_46277,N_44395,N_44552);
nand U46278 (N_46278,N_43358,N_44289);
xor U46279 (N_46279,N_43782,N_44262);
xnor U46280 (N_46280,N_44102,N_44350);
xor U46281 (N_46281,N_44702,N_44323);
nor U46282 (N_46282,N_43961,N_42918);
and U46283 (N_46283,N_42662,N_43900);
nor U46284 (N_46284,N_44011,N_44778);
and U46285 (N_46285,N_43326,N_44521);
xnor U46286 (N_46286,N_42975,N_43394);
or U46287 (N_46287,N_42663,N_43250);
or U46288 (N_46288,N_42550,N_43466);
or U46289 (N_46289,N_44927,N_43331);
nand U46290 (N_46290,N_43610,N_42772);
nand U46291 (N_46291,N_42691,N_44505);
nand U46292 (N_46292,N_44745,N_44933);
and U46293 (N_46293,N_44636,N_44434);
nor U46294 (N_46294,N_43971,N_43858);
or U46295 (N_46295,N_42701,N_43961);
nand U46296 (N_46296,N_44970,N_44880);
nand U46297 (N_46297,N_43082,N_42669);
or U46298 (N_46298,N_43604,N_44797);
xnor U46299 (N_46299,N_43225,N_44783);
or U46300 (N_46300,N_44292,N_44898);
nand U46301 (N_46301,N_42978,N_44332);
xor U46302 (N_46302,N_43137,N_42787);
nor U46303 (N_46303,N_44943,N_43436);
nand U46304 (N_46304,N_44490,N_44592);
and U46305 (N_46305,N_44587,N_43087);
or U46306 (N_46306,N_43395,N_44462);
and U46307 (N_46307,N_43434,N_44361);
or U46308 (N_46308,N_43594,N_42667);
or U46309 (N_46309,N_42826,N_42607);
xnor U46310 (N_46310,N_43469,N_42538);
and U46311 (N_46311,N_43984,N_44628);
nor U46312 (N_46312,N_44672,N_44267);
or U46313 (N_46313,N_44164,N_44264);
nor U46314 (N_46314,N_43526,N_44288);
xnor U46315 (N_46315,N_44932,N_44832);
nor U46316 (N_46316,N_43726,N_44343);
xor U46317 (N_46317,N_44298,N_43607);
or U46318 (N_46318,N_44511,N_42638);
nand U46319 (N_46319,N_44187,N_43899);
or U46320 (N_46320,N_42673,N_43850);
or U46321 (N_46321,N_43255,N_42782);
nor U46322 (N_46322,N_42897,N_43592);
xnor U46323 (N_46323,N_43716,N_44085);
xor U46324 (N_46324,N_43191,N_44104);
and U46325 (N_46325,N_43231,N_43391);
xor U46326 (N_46326,N_43921,N_42590);
nand U46327 (N_46327,N_44601,N_44894);
nand U46328 (N_46328,N_44961,N_44023);
and U46329 (N_46329,N_43841,N_44321);
and U46330 (N_46330,N_44440,N_44786);
and U46331 (N_46331,N_43467,N_44500);
nor U46332 (N_46332,N_42911,N_44476);
nand U46333 (N_46333,N_44648,N_44638);
and U46334 (N_46334,N_42973,N_43803);
xor U46335 (N_46335,N_44507,N_42798);
and U46336 (N_46336,N_44923,N_42631);
nand U46337 (N_46337,N_43301,N_43374);
nor U46338 (N_46338,N_44535,N_44312);
and U46339 (N_46339,N_44513,N_42700);
or U46340 (N_46340,N_42858,N_42668);
nand U46341 (N_46341,N_44125,N_42950);
or U46342 (N_46342,N_43615,N_43910);
or U46343 (N_46343,N_43157,N_44512);
nand U46344 (N_46344,N_44607,N_44597);
nor U46345 (N_46345,N_43566,N_43916);
xor U46346 (N_46346,N_44366,N_43118);
and U46347 (N_46347,N_43528,N_42516);
or U46348 (N_46348,N_44796,N_44698);
xor U46349 (N_46349,N_44007,N_43141);
nor U46350 (N_46350,N_43634,N_44549);
or U46351 (N_46351,N_43566,N_44134);
and U46352 (N_46352,N_44124,N_44388);
and U46353 (N_46353,N_42930,N_43696);
xnor U46354 (N_46354,N_42919,N_44165);
and U46355 (N_46355,N_43159,N_44059);
or U46356 (N_46356,N_42562,N_44781);
nor U46357 (N_46357,N_44947,N_44911);
nand U46358 (N_46358,N_44021,N_43889);
xor U46359 (N_46359,N_44747,N_44273);
nand U46360 (N_46360,N_44980,N_44228);
nor U46361 (N_46361,N_44951,N_44374);
nand U46362 (N_46362,N_44821,N_44075);
and U46363 (N_46363,N_43093,N_44593);
nor U46364 (N_46364,N_42812,N_44254);
nand U46365 (N_46365,N_42820,N_43052);
xnor U46366 (N_46366,N_43027,N_42577);
or U46367 (N_46367,N_43982,N_42942);
and U46368 (N_46368,N_43924,N_43813);
xor U46369 (N_46369,N_43656,N_44121);
nand U46370 (N_46370,N_44501,N_42859);
xor U46371 (N_46371,N_43435,N_42956);
or U46372 (N_46372,N_44416,N_44503);
and U46373 (N_46373,N_44982,N_42813);
xor U46374 (N_46374,N_42687,N_42510);
xnor U46375 (N_46375,N_43007,N_44493);
and U46376 (N_46376,N_42738,N_44674);
nor U46377 (N_46377,N_43825,N_43646);
or U46378 (N_46378,N_43136,N_42772);
xnor U46379 (N_46379,N_43142,N_44546);
xor U46380 (N_46380,N_44966,N_43868);
nor U46381 (N_46381,N_44114,N_42914);
and U46382 (N_46382,N_42734,N_44858);
nor U46383 (N_46383,N_43587,N_44578);
or U46384 (N_46384,N_42615,N_44129);
xnor U46385 (N_46385,N_43511,N_43494);
xor U46386 (N_46386,N_43545,N_42719);
nand U46387 (N_46387,N_44497,N_43247);
nor U46388 (N_46388,N_43900,N_43007);
or U46389 (N_46389,N_44707,N_43886);
and U46390 (N_46390,N_44372,N_42763);
or U46391 (N_46391,N_43847,N_43333);
nor U46392 (N_46392,N_44748,N_44785);
or U46393 (N_46393,N_43111,N_43504);
and U46394 (N_46394,N_44490,N_43888);
or U46395 (N_46395,N_43118,N_43123);
and U46396 (N_46396,N_43717,N_44691);
nor U46397 (N_46397,N_44805,N_44633);
nand U46398 (N_46398,N_44410,N_44389);
nor U46399 (N_46399,N_42803,N_43984);
xor U46400 (N_46400,N_42951,N_44644);
nor U46401 (N_46401,N_44367,N_44873);
xor U46402 (N_46402,N_43785,N_43349);
nand U46403 (N_46403,N_42869,N_44214);
nor U46404 (N_46404,N_42849,N_42547);
xnor U46405 (N_46405,N_43511,N_42847);
xnor U46406 (N_46406,N_44254,N_43031);
nand U46407 (N_46407,N_44651,N_43185);
and U46408 (N_46408,N_42890,N_42778);
and U46409 (N_46409,N_43671,N_43363);
and U46410 (N_46410,N_42907,N_43459);
nand U46411 (N_46411,N_43441,N_43803);
nor U46412 (N_46412,N_44745,N_44673);
and U46413 (N_46413,N_43483,N_44849);
nor U46414 (N_46414,N_43550,N_43038);
nand U46415 (N_46415,N_42951,N_43851);
nor U46416 (N_46416,N_44185,N_44376);
and U46417 (N_46417,N_43183,N_42597);
xnor U46418 (N_46418,N_43473,N_43003);
and U46419 (N_46419,N_43054,N_43675);
and U46420 (N_46420,N_43327,N_44466);
and U46421 (N_46421,N_44909,N_42948);
or U46422 (N_46422,N_43964,N_43373);
nor U46423 (N_46423,N_42578,N_42829);
or U46424 (N_46424,N_43483,N_42898);
and U46425 (N_46425,N_42985,N_44449);
xnor U46426 (N_46426,N_44789,N_42983);
and U46427 (N_46427,N_44046,N_42721);
nand U46428 (N_46428,N_43363,N_43830);
or U46429 (N_46429,N_42774,N_42974);
nand U46430 (N_46430,N_44653,N_44581);
nand U46431 (N_46431,N_43153,N_42638);
and U46432 (N_46432,N_44043,N_44544);
or U46433 (N_46433,N_42559,N_43538);
nand U46434 (N_46434,N_42897,N_42545);
and U46435 (N_46435,N_43200,N_42753);
nor U46436 (N_46436,N_42729,N_43202);
and U46437 (N_46437,N_44208,N_44039);
nand U46438 (N_46438,N_43307,N_42927);
xnor U46439 (N_46439,N_44105,N_43007);
or U46440 (N_46440,N_44472,N_43679);
xor U46441 (N_46441,N_44430,N_42909);
or U46442 (N_46442,N_44706,N_44524);
nand U46443 (N_46443,N_42753,N_42563);
nor U46444 (N_46444,N_44003,N_43203);
nor U46445 (N_46445,N_43346,N_43453);
nor U46446 (N_46446,N_44007,N_44511);
and U46447 (N_46447,N_44008,N_44963);
nand U46448 (N_46448,N_43390,N_44861);
nand U46449 (N_46449,N_43768,N_43955);
xor U46450 (N_46450,N_44255,N_43181);
nor U46451 (N_46451,N_44297,N_44823);
xor U46452 (N_46452,N_44325,N_43910);
or U46453 (N_46453,N_42788,N_44999);
or U46454 (N_46454,N_42659,N_44630);
nor U46455 (N_46455,N_44917,N_43338);
xor U46456 (N_46456,N_44791,N_44827);
xnor U46457 (N_46457,N_43438,N_43918);
nand U46458 (N_46458,N_43672,N_44566);
and U46459 (N_46459,N_44296,N_44657);
nor U46460 (N_46460,N_44354,N_44987);
and U46461 (N_46461,N_43610,N_44273);
nand U46462 (N_46462,N_43081,N_42857);
xor U46463 (N_46463,N_44591,N_44729);
and U46464 (N_46464,N_43424,N_44320);
nand U46465 (N_46465,N_43983,N_43439);
nand U46466 (N_46466,N_42972,N_43636);
or U46467 (N_46467,N_44613,N_44482);
nor U46468 (N_46468,N_43631,N_43873);
or U46469 (N_46469,N_44200,N_42745);
nor U46470 (N_46470,N_43802,N_42834);
or U46471 (N_46471,N_44289,N_44869);
nand U46472 (N_46472,N_43190,N_44740);
or U46473 (N_46473,N_44932,N_42512);
nor U46474 (N_46474,N_42641,N_44304);
and U46475 (N_46475,N_42594,N_43306);
nand U46476 (N_46476,N_43447,N_43653);
nor U46477 (N_46477,N_42814,N_43203);
nor U46478 (N_46478,N_43076,N_43953);
and U46479 (N_46479,N_44580,N_42920);
and U46480 (N_46480,N_42994,N_43211);
or U46481 (N_46481,N_42680,N_43988);
or U46482 (N_46482,N_43046,N_42929);
nand U46483 (N_46483,N_43278,N_43272);
xnor U46484 (N_46484,N_44190,N_42610);
xnor U46485 (N_46485,N_43736,N_44137);
nand U46486 (N_46486,N_42638,N_43927);
and U46487 (N_46487,N_44695,N_44622);
nor U46488 (N_46488,N_42871,N_44606);
xor U46489 (N_46489,N_42832,N_44543);
nand U46490 (N_46490,N_44679,N_44695);
nand U46491 (N_46491,N_42728,N_44045);
and U46492 (N_46492,N_43838,N_43509);
nor U46493 (N_46493,N_44533,N_42654);
nor U46494 (N_46494,N_43470,N_44234);
and U46495 (N_46495,N_44276,N_44461);
xor U46496 (N_46496,N_44930,N_43310);
nand U46497 (N_46497,N_42542,N_43452);
and U46498 (N_46498,N_44611,N_44278);
or U46499 (N_46499,N_44985,N_44263);
or U46500 (N_46500,N_44201,N_43290);
and U46501 (N_46501,N_43378,N_42517);
or U46502 (N_46502,N_43899,N_44086);
nor U46503 (N_46503,N_42895,N_43217);
or U46504 (N_46504,N_43420,N_44493);
or U46505 (N_46505,N_43040,N_43490);
xor U46506 (N_46506,N_43947,N_44347);
or U46507 (N_46507,N_42909,N_43707);
xnor U46508 (N_46508,N_42807,N_43769);
nor U46509 (N_46509,N_42857,N_44246);
nand U46510 (N_46510,N_42659,N_44468);
nand U46511 (N_46511,N_44149,N_43381);
nand U46512 (N_46512,N_43828,N_42949);
nor U46513 (N_46513,N_44551,N_42862);
or U46514 (N_46514,N_44416,N_43472);
or U46515 (N_46515,N_43253,N_42798);
or U46516 (N_46516,N_42598,N_43136);
nand U46517 (N_46517,N_43869,N_42513);
xnor U46518 (N_46518,N_43889,N_44253);
or U46519 (N_46519,N_43694,N_42912);
nand U46520 (N_46520,N_44455,N_44150);
nor U46521 (N_46521,N_43832,N_43207);
nand U46522 (N_46522,N_44895,N_44883);
or U46523 (N_46523,N_43417,N_44388);
nor U46524 (N_46524,N_43637,N_42777);
and U46525 (N_46525,N_43952,N_42667);
xnor U46526 (N_46526,N_43964,N_43358);
xnor U46527 (N_46527,N_42898,N_43399);
nor U46528 (N_46528,N_44496,N_43646);
nand U46529 (N_46529,N_44262,N_43369);
and U46530 (N_46530,N_42573,N_42508);
nand U46531 (N_46531,N_44504,N_43095);
and U46532 (N_46532,N_42795,N_44183);
and U46533 (N_46533,N_42743,N_43427);
and U46534 (N_46534,N_44902,N_42512);
and U46535 (N_46535,N_44347,N_43226);
xor U46536 (N_46536,N_43625,N_42873);
or U46537 (N_46537,N_43380,N_43269);
or U46538 (N_46538,N_43311,N_44882);
nand U46539 (N_46539,N_42759,N_42766);
and U46540 (N_46540,N_42617,N_44313);
nand U46541 (N_46541,N_42906,N_43307);
nor U46542 (N_46542,N_44633,N_42746);
nand U46543 (N_46543,N_43030,N_44425);
nor U46544 (N_46544,N_43871,N_43476);
xor U46545 (N_46545,N_44764,N_43093);
xnor U46546 (N_46546,N_44093,N_42605);
nor U46547 (N_46547,N_44329,N_43946);
nand U46548 (N_46548,N_43781,N_42646);
nand U46549 (N_46549,N_42624,N_42566);
xor U46550 (N_46550,N_43232,N_43220);
xor U46551 (N_46551,N_44438,N_43059);
or U46552 (N_46552,N_44367,N_43435);
nand U46553 (N_46553,N_43045,N_44862);
and U46554 (N_46554,N_43486,N_43936);
nor U46555 (N_46555,N_43396,N_43089);
nor U46556 (N_46556,N_44255,N_43775);
or U46557 (N_46557,N_43103,N_44869);
or U46558 (N_46558,N_42698,N_44546);
and U46559 (N_46559,N_44019,N_43402);
nor U46560 (N_46560,N_42776,N_44640);
or U46561 (N_46561,N_44657,N_43123);
nand U46562 (N_46562,N_44020,N_43864);
nand U46563 (N_46563,N_43172,N_43463);
nand U46564 (N_46564,N_44716,N_44527);
nor U46565 (N_46565,N_43955,N_44900);
nand U46566 (N_46566,N_43695,N_43498);
xor U46567 (N_46567,N_43855,N_44210);
nand U46568 (N_46568,N_43857,N_42830);
and U46569 (N_46569,N_43441,N_43169);
or U46570 (N_46570,N_44932,N_43395);
or U46571 (N_46571,N_43897,N_44183);
nand U46572 (N_46572,N_43788,N_43879);
and U46573 (N_46573,N_44691,N_44041);
nor U46574 (N_46574,N_44584,N_43968);
nand U46575 (N_46575,N_44029,N_42920);
and U46576 (N_46576,N_43702,N_42891);
nor U46577 (N_46577,N_44194,N_42818);
nor U46578 (N_46578,N_42927,N_43514);
xor U46579 (N_46579,N_44900,N_43355);
nand U46580 (N_46580,N_43306,N_44806);
nand U46581 (N_46581,N_44618,N_43383);
and U46582 (N_46582,N_42670,N_43226);
and U46583 (N_46583,N_44474,N_42606);
and U46584 (N_46584,N_44450,N_43808);
nand U46585 (N_46585,N_43887,N_43413);
nand U46586 (N_46586,N_43407,N_44124);
xor U46587 (N_46587,N_43574,N_42914);
nand U46588 (N_46588,N_43786,N_43595);
and U46589 (N_46589,N_43830,N_43348);
and U46590 (N_46590,N_44930,N_42837);
or U46591 (N_46591,N_44635,N_43709);
and U46592 (N_46592,N_44348,N_44733);
xnor U46593 (N_46593,N_43131,N_42970);
nor U46594 (N_46594,N_42698,N_43956);
and U46595 (N_46595,N_43481,N_43883);
nand U46596 (N_46596,N_44920,N_43605);
or U46597 (N_46597,N_43797,N_43152);
xnor U46598 (N_46598,N_43223,N_43462);
xor U46599 (N_46599,N_43593,N_42763);
nor U46600 (N_46600,N_43345,N_43879);
nand U46601 (N_46601,N_44183,N_43419);
xnor U46602 (N_46602,N_42500,N_44539);
nand U46603 (N_46603,N_43804,N_43207);
nor U46604 (N_46604,N_43604,N_43098);
nand U46605 (N_46605,N_43945,N_44966);
nor U46606 (N_46606,N_44507,N_44550);
nand U46607 (N_46607,N_44535,N_44687);
nand U46608 (N_46608,N_44623,N_43798);
xnor U46609 (N_46609,N_43888,N_44827);
nor U46610 (N_46610,N_42581,N_43140);
and U46611 (N_46611,N_43649,N_43343);
nand U46612 (N_46612,N_43927,N_43986);
and U46613 (N_46613,N_43038,N_42569);
nor U46614 (N_46614,N_44816,N_43483);
nor U46615 (N_46615,N_43333,N_43685);
and U46616 (N_46616,N_44847,N_42798);
and U46617 (N_46617,N_43902,N_44970);
and U46618 (N_46618,N_42760,N_43012);
xor U46619 (N_46619,N_44733,N_44493);
and U46620 (N_46620,N_44016,N_43826);
and U46621 (N_46621,N_44031,N_43611);
xnor U46622 (N_46622,N_44516,N_44806);
nand U46623 (N_46623,N_43376,N_43548);
and U46624 (N_46624,N_44334,N_44875);
nor U46625 (N_46625,N_43246,N_43469);
or U46626 (N_46626,N_43171,N_43395);
nand U46627 (N_46627,N_43431,N_44536);
or U46628 (N_46628,N_43970,N_44226);
nand U46629 (N_46629,N_43141,N_44878);
xnor U46630 (N_46630,N_44690,N_44618);
or U46631 (N_46631,N_44156,N_43100);
and U46632 (N_46632,N_42777,N_43943);
or U46633 (N_46633,N_42673,N_43706);
nor U46634 (N_46634,N_43239,N_44649);
and U46635 (N_46635,N_42940,N_44478);
nor U46636 (N_46636,N_44067,N_42563);
and U46637 (N_46637,N_43175,N_44580);
nor U46638 (N_46638,N_43077,N_44335);
or U46639 (N_46639,N_42573,N_43606);
and U46640 (N_46640,N_43348,N_43230);
xnor U46641 (N_46641,N_43285,N_44675);
nor U46642 (N_46642,N_44345,N_43705);
nor U46643 (N_46643,N_43876,N_44549);
or U46644 (N_46644,N_43942,N_43039);
nor U46645 (N_46645,N_44208,N_43977);
nand U46646 (N_46646,N_42668,N_43789);
and U46647 (N_46647,N_43638,N_44060);
nand U46648 (N_46648,N_43274,N_43004);
xnor U46649 (N_46649,N_43010,N_44712);
nor U46650 (N_46650,N_43891,N_44432);
or U46651 (N_46651,N_44969,N_44845);
nand U46652 (N_46652,N_44577,N_43271);
and U46653 (N_46653,N_44524,N_42665);
xor U46654 (N_46654,N_44324,N_43485);
or U46655 (N_46655,N_44106,N_44668);
xnor U46656 (N_46656,N_43497,N_44460);
and U46657 (N_46657,N_43883,N_43889);
or U46658 (N_46658,N_42542,N_43932);
nor U46659 (N_46659,N_43656,N_43538);
and U46660 (N_46660,N_44174,N_44018);
nand U46661 (N_46661,N_43105,N_43060);
nor U46662 (N_46662,N_44492,N_44111);
nor U46663 (N_46663,N_44568,N_42704);
or U46664 (N_46664,N_44247,N_44873);
nand U46665 (N_46665,N_42732,N_43631);
xor U46666 (N_46666,N_43442,N_43607);
or U46667 (N_46667,N_43196,N_42661);
nor U46668 (N_46668,N_44371,N_42633);
nor U46669 (N_46669,N_43231,N_44330);
xor U46670 (N_46670,N_44105,N_44136);
and U46671 (N_46671,N_44343,N_43276);
nand U46672 (N_46672,N_42816,N_43823);
xnor U46673 (N_46673,N_43103,N_42840);
xnor U46674 (N_46674,N_42698,N_43674);
and U46675 (N_46675,N_43689,N_44822);
nand U46676 (N_46676,N_42803,N_44867);
nor U46677 (N_46677,N_43937,N_42519);
nor U46678 (N_46678,N_44622,N_43765);
nor U46679 (N_46679,N_44812,N_44981);
and U46680 (N_46680,N_44463,N_44075);
or U46681 (N_46681,N_44021,N_43368);
nor U46682 (N_46682,N_43429,N_43966);
or U46683 (N_46683,N_44958,N_44885);
or U46684 (N_46684,N_43340,N_43037);
nand U46685 (N_46685,N_43473,N_44172);
or U46686 (N_46686,N_43191,N_43443);
or U46687 (N_46687,N_43366,N_44440);
nand U46688 (N_46688,N_44101,N_43589);
nand U46689 (N_46689,N_42542,N_43989);
nor U46690 (N_46690,N_42590,N_44068);
nor U46691 (N_46691,N_44962,N_44326);
and U46692 (N_46692,N_44137,N_42568);
and U46693 (N_46693,N_43229,N_43820);
nand U46694 (N_46694,N_43826,N_44314);
and U46695 (N_46695,N_44120,N_44726);
or U46696 (N_46696,N_44713,N_43546);
and U46697 (N_46697,N_44890,N_44539);
and U46698 (N_46698,N_42952,N_43958);
nor U46699 (N_46699,N_44890,N_44492);
nor U46700 (N_46700,N_43466,N_44334);
nor U46701 (N_46701,N_42596,N_44195);
xor U46702 (N_46702,N_44285,N_42969);
xor U46703 (N_46703,N_44852,N_43658);
nand U46704 (N_46704,N_42806,N_44186);
nand U46705 (N_46705,N_43097,N_44103);
or U46706 (N_46706,N_44549,N_42910);
nand U46707 (N_46707,N_44621,N_43627);
or U46708 (N_46708,N_44146,N_44943);
xnor U46709 (N_46709,N_44065,N_43826);
nand U46710 (N_46710,N_43387,N_44550);
and U46711 (N_46711,N_43922,N_44525);
nand U46712 (N_46712,N_43165,N_42611);
and U46713 (N_46713,N_42946,N_44104);
xnor U46714 (N_46714,N_44440,N_43057);
nand U46715 (N_46715,N_44381,N_43738);
xor U46716 (N_46716,N_42535,N_44122);
xnor U46717 (N_46717,N_43332,N_42660);
or U46718 (N_46718,N_44050,N_43554);
and U46719 (N_46719,N_43642,N_43800);
and U46720 (N_46720,N_43755,N_43131);
and U46721 (N_46721,N_42523,N_44031);
xor U46722 (N_46722,N_43322,N_43992);
or U46723 (N_46723,N_43994,N_43171);
or U46724 (N_46724,N_43814,N_42846);
nand U46725 (N_46725,N_44452,N_44323);
and U46726 (N_46726,N_43024,N_42803);
xnor U46727 (N_46727,N_43198,N_43646);
and U46728 (N_46728,N_44825,N_44924);
and U46729 (N_46729,N_43273,N_44421);
and U46730 (N_46730,N_44273,N_44742);
and U46731 (N_46731,N_44136,N_44595);
or U46732 (N_46732,N_43556,N_43288);
or U46733 (N_46733,N_43641,N_44078);
nor U46734 (N_46734,N_43547,N_44481);
and U46735 (N_46735,N_44490,N_43702);
xor U46736 (N_46736,N_43426,N_44993);
nand U46737 (N_46737,N_43884,N_43580);
and U46738 (N_46738,N_44668,N_42928);
or U46739 (N_46739,N_44981,N_43253);
or U46740 (N_46740,N_43676,N_43304);
or U46741 (N_46741,N_44771,N_43239);
nor U46742 (N_46742,N_44227,N_43207);
or U46743 (N_46743,N_43989,N_44062);
xnor U46744 (N_46744,N_44572,N_44603);
or U46745 (N_46745,N_43235,N_43429);
and U46746 (N_46746,N_43202,N_43417);
nor U46747 (N_46747,N_42872,N_43471);
nand U46748 (N_46748,N_42973,N_42737);
or U46749 (N_46749,N_43250,N_44740);
nand U46750 (N_46750,N_43221,N_42793);
and U46751 (N_46751,N_44883,N_42585);
nand U46752 (N_46752,N_43381,N_44766);
xnor U46753 (N_46753,N_44007,N_43376);
and U46754 (N_46754,N_44161,N_43012);
or U46755 (N_46755,N_44212,N_44309);
xnor U46756 (N_46756,N_43762,N_44708);
and U46757 (N_46757,N_44036,N_44484);
nand U46758 (N_46758,N_44724,N_43519);
nand U46759 (N_46759,N_42899,N_44890);
xnor U46760 (N_46760,N_43125,N_43560);
and U46761 (N_46761,N_44673,N_42876);
xor U46762 (N_46762,N_43478,N_44735);
nor U46763 (N_46763,N_44837,N_43575);
and U46764 (N_46764,N_43771,N_43633);
and U46765 (N_46765,N_44862,N_43452);
or U46766 (N_46766,N_43342,N_43804);
xnor U46767 (N_46767,N_43316,N_44568);
or U46768 (N_46768,N_43225,N_42830);
nor U46769 (N_46769,N_42578,N_43689);
xnor U46770 (N_46770,N_44572,N_42830);
nand U46771 (N_46771,N_43012,N_43280);
and U46772 (N_46772,N_44866,N_43445);
or U46773 (N_46773,N_44172,N_44739);
nor U46774 (N_46774,N_43703,N_44765);
and U46775 (N_46775,N_42694,N_43319);
xor U46776 (N_46776,N_43682,N_44625);
nand U46777 (N_46777,N_44463,N_42818);
or U46778 (N_46778,N_43785,N_43286);
nand U46779 (N_46779,N_42818,N_44916);
or U46780 (N_46780,N_43529,N_43803);
nand U46781 (N_46781,N_43453,N_44290);
nor U46782 (N_46782,N_43017,N_43319);
or U46783 (N_46783,N_43220,N_44623);
nor U46784 (N_46784,N_43367,N_43106);
and U46785 (N_46785,N_44746,N_42867);
nor U46786 (N_46786,N_44190,N_44963);
or U46787 (N_46787,N_44712,N_43223);
and U46788 (N_46788,N_43169,N_44919);
xor U46789 (N_46789,N_43503,N_42756);
nor U46790 (N_46790,N_43444,N_42697);
and U46791 (N_46791,N_42721,N_43176);
nand U46792 (N_46792,N_44355,N_43713);
or U46793 (N_46793,N_44098,N_44316);
nor U46794 (N_46794,N_43998,N_43937);
nor U46795 (N_46795,N_44491,N_43481);
nor U46796 (N_46796,N_44656,N_43582);
xor U46797 (N_46797,N_44678,N_44286);
xor U46798 (N_46798,N_42523,N_42779);
nor U46799 (N_46799,N_43795,N_44501);
nand U46800 (N_46800,N_43195,N_43130);
and U46801 (N_46801,N_43177,N_43958);
and U46802 (N_46802,N_42812,N_44252);
or U46803 (N_46803,N_43102,N_44739);
nor U46804 (N_46804,N_43923,N_43287);
and U46805 (N_46805,N_43957,N_44077);
nand U46806 (N_46806,N_44068,N_44424);
nor U46807 (N_46807,N_44408,N_43666);
nand U46808 (N_46808,N_43915,N_43209);
nor U46809 (N_46809,N_43547,N_44589);
nor U46810 (N_46810,N_43202,N_44871);
nand U46811 (N_46811,N_42853,N_44886);
and U46812 (N_46812,N_43485,N_42566);
and U46813 (N_46813,N_43351,N_44187);
nor U46814 (N_46814,N_44525,N_43800);
nand U46815 (N_46815,N_43909,N_44973);
nand U46816 (N_46816,N_43221,N_44064);
xnor U46817 (N_46817,N_43990,N_43939);
and U46818 (N_46818,N_44401,N_43467);
nand U46819 (N_46819,N_44474,N_44235);
nor U46820 (N_46820,N_44179,N_42973);
xnor U46821 (N_46821,N_42792,N_43730);
xor U46822 (N_46822,N_43876,N_42802);
nand U46823 (N_46823,N_43629,N_43635);
xnor U46824 (N_46824,N_42544,N_43283);
nand U46825 (N_46825,N_42673,N_42753);
or U46826 (N_46826,N_44243,N_44900);
nand U46827 (N_46827,N_44414,N_42983);
nor U46828 (N_46828,N_43332,N_44088);
or U46829 (N_46829,N_44429,N_43190);
or U46830 (N_46830,N_44197,N_42645);
or U46831 (N_46831,N_44662,N_43720);
nor U46832 (N_46832,N_44053,N_43608);
or U46833 (N_46833,N_43733,N_42671);
or U46834 (N_46834,N_42910,N_44938);
xor U46835 (N_46835,N_43217,N_44482);
or U46836 (N_46836,N_44232,N_43761);
xnor U46837 (N_46837,N_44560,N_43825);
or U46838 (N_46838,N_43207,N_43460);
and U46839 (N_46839,N_44996,N_43614);
or U46840 (N_46840,N_44125,N_42794);
nor U46841 (N_46841,N_44878,N_44781);
nor U46842 (N_46842,N_44563,N_44975);
xor U46843 (N_46843,N_43304,N_43398);
xor U46844 (N_46844,N_43033,N_43337);
xnor U46845 (N_46845,N_44911,N_43461);
or U46846 (N_46846,N_44860,N_43916);
xor U46847 (N_46847,N_44862,N_43856);
nor U46848 (N_46848,N_43033,N_43864);
and U46849 (N_46849,N_44059,N_43155);
and U46850 (N_46850,N_42810,N_44103);
or U46851 (N_46851,N_43897,N_43915);
xnor U46852 (N_46852,N_43160,N_44360);
nand U46853 (N_46853,N_43734,N_44781);
and U46854 (N_46854,N_44782,N_42627);
nor U46855 (N_46855,N_44220,N_43025);
or U46856 (N_46856,N_43929,N_44590);
nor U46857 (N_46857,N_43652,N_42552);
xor U46858 (N_46858,N_43599,N_44944);
nor U46859 (N_46859,N_42877,N_44524);
nor U46860 (N_46860,N_42752,N_44049);
nand U46861 (N_46861,N_44040,N_44437);
and U46862 (N_46862,N_44485,N_42715);
xor U46863 (N_46863,N_43463,N_44803);
nor U46864 (N_46864,N_43306,N_44002);
or U46865 (N_46865,N_43876,N_43947);
nor U46866 (N_46866,N_43252,N_42937);
nor U46867 (N_46867,N_42993,N_43900);
xor U46868 (N_46868,N_44711,N_43585);
nand U46869 (N_46869,N_43409,N_43322);
nand U46870 (N_46870,N_42980,N_44691);
nand U46871 (N_46871,N_42864,N_44618);
xor U46872 (N_46872,N_43430,N_42771);
nand U46873 (N_46873,N_43560,N_44851);
or U46874 (N_46874,N_42946,N_44283);
xor U46875 (N_46875,N_43583,N_44720);
xnor U46876 (N_46876,N_42824,N_43358);
nor U46877 (N_46877,N_43183,N_42716);
and U46878 (N_46878,N_43780,N_42841);
nand U46879 (N_46879,N_43866,N_44683);
xnor U46880 (N_46880,N_43982,N_43144);
nand U46881 (N_46881,N_42734,N_44256);
nor U46882 (N_46882,N_44111,N_44799);
or U46883 (N_46883,N_43841,N_43571);
nand U46884 (N_46884,N_43809,N_44930);
or U46885 (N_46885,N_44627,N_43340);
or U46886 (N_46886,N_42786,N_43234);
nand U46887 (N_46887,N_42919,N_44435);
nor U46888 (N_46888,N_44755,N_43762);
and U46889 (N_46889,N_43064,N_44585);
nor U46890 (N_46890,N_44605,N_42959);
and U46891 (N_46891,N_42804,N_44745);
nand U46892 (N_46892,N_44152,N_43781);
nand U46893 (N_46893,N_43871,N_43908);
and U46894 (N_46894,N_43734,N_42729);
or U46895 (N_46895,N_44093,N_44479);
nand U46896 (N_46896,N_44687,N_43983);
nor U46897 (N_46897,N_44067,N_42744);
or U46898 (N_46898,N_44898,N_43517);
xnor U46899 (N_46899,N_43908,N_43827);
xnor U46900 (N_46900,N_42744,N_42869);
nand U46901 (N_46901,N_44209,N_42916);
nand U46902 (N_46902,N_44408,N_43434);
nor U46903 (N_46903,N_44641,N_42991);
nor U46904 (N_46904,N_43014,N_42566);
and U46905 (N_46905,N_43259,N_43329);
xor U46906 (N_46906,N_44647,N_44066);
or U46907 (N_46907,N_42722,N_44465);
and U46908 (N_46908,N_43115,N_42960);
xor U46909 (N_46909,N_44693,N_44323);
nor U46910 (N_46910,N_44869,N_43327);
nor U46911 (N_46911,N_43254,N_43282);
and U46912 (N_46912,N_43107,N_44282);
xnor U46913 (N_46913,N_43348,N_43468);
nor U46914 (N_46914,N_44758,N_43684);
or U46915 (N_46915,N_44470,N_44338);
or U46916 (N_46916,N_42887,N_43344);
xor U46917 (N_46917,N_43470,N_44688);
or U46918 (N_46918,N_42930,N_44308);
nand U46919 (N_46919,N_43439,N_44278);
or U46920 (N_46920,N_44963,N_42559);
and U46921 (N_46921,N_42683,N_42950);
and U46922 (N_46922,N_42896,N_43537);
and U46923 (N_46923,N_42789,N_42530);
nor U46924 (N_46924,N_42916,N_44282);
or U46925 (N_46925,N_43500,N_43690);
xnor U46926 (N_46926,N_43611,N_43237);
xnor U46927 (N_46927,N_44992,N_43504);
or U46928 (N_46928,N_44520,N_42969);
or U46929 (N_46929,N_44722,N_43462);
nand U46930 (N_46930,N_44827,N_42801);
xor U46931 (N_46931,N_43538,N_42746);
nor U46932 (N_46932,N_44196,N_44787);
nand U46933 (N_46933,N_43055,N_42712);
or U46934 (N_46934,N_44427,N_43715);
xnor U46935 (N_46935,N_44530,N_44752);
xor U46936 (N_46936,N_43033,N_43569);
nor U46937 (N_46937,N_42740,N_42624);
xnor U46938 (N_46938,N_43387,N_44144);
nand U46939 (N_46939,N_42864,N_43144);
nand U46940 (N_46940,N_44661,N_42917);
nand U46941 (N_46941,N_43397,N_43189);
nand U46942 (N_46942,N_44525,N_44347);
xor U46943 (N_46943,N_43597,N_44359);
and U46944 (N_46944,N_42935,N_43306);
or U46945 (N_46945,N_44059,N_43791);
xor U46946 (N_46946,N_44963,N_42896);
nand U46947 (N_46947,N_44117,N_42746);
xnor U46948 (N_46948,N_42545,N_44732);
or U46949 (N_46949,N_43462,N_42701);
xnor U46950 (N_46950,N_43567,N_43148);
xor U46951 (N_46951,N_44936,N_44253);
nor U46952 (N_46952,N_43368,N_43519);
xnor U46953 (N_46953,N_43890,N_43567);
and U46954 (N_46954,N_43907,N_42788);
xnor U46955 (N_46955,N_43005,N_44040);
and U46956 (N_46956,N_43866,N_42797);
nor U46957 (N_46957,N_43178,N_44349);
nor U46958 (N_46958,N_43283,N_44687);
nand U46959 (N_46959,N_44212,N_43405);
and U46960 (N_46960,N_44041,N_44704);
xnor U46961 (N_46961,N_42707,N_44085);
or U46962 (N_46962,N_43110,N_44257);
xor U46963 (N_46963,N_44075,N_43025);
xor U46964 (N_46964,N_43595,N_44644);
nand U46965 (N_46965,N_43618,N_44549);
nand U46966 (N_46966,N_43775,N_42845);
and U46967 (N_46967,N_43925,N_44199);
xnor U46968 (N_46968,N_44437,N_44680);
nand U46969 (N_46969,N_43479,N_44634);
nand U46970 (N_46970,N_44900,N_42549);
nand U46971 (N_46971,N_43456,N_43308);
xor U46972 (N_46972,N_44902,N_44077);
xor U46973 (N_46973,N_44379,N_43932);
xnor U46974 (N_46974,N_43422,N_43070);
and U46975 (N_46975,N_42737,N_43777);
xnor U46976 (N_46976,N_44125,N_42863);
nand U46977 (N_46977,N_42507,N_42780);
and U46978 (N_46978,N_43887,N_42747);
or U46979 (N_46979,N_44022,N_44588);
or U46980 (N_46980,N_44465,N_42774);
xnor U46981 (N_46981,N_43247,N_43938);
xnor U46982 (N_46982,N_43497,N_43864);
nor U46983 (N_46983,N_44919,N_44058);
xnor U46984 (N_46984,N_42836,N_42675);
nor U46985 (N_46985,N_42690,N_44061);
and U46986 (N_46986,N_43222,N_42654);
xnor U46987 (N_46987,N_42735,N_44837);
xnor U46988 (N_46988,N_43834,N_42570);
or U46989 (N_46989,N_43878,N_44950);
and U46990 (N_46990,N_43844,N_44082);
and U46991 (N_46991,N_43287,N_44863);
xnor U46992 (N_46992,N_44863,N_44997);
nand U46993 (N_46993,N_44110,N_43445);
nor U46994 (N_46994,N_44712,N_43916);
xnor U46995 (N_46995,N_44709,N_44872);
nand U46996 (N_46996,N_43244,N_44622);
or U46997 (N_46997,N_44758,N_43418);
nor U46998 (N_46998,N_43597,N_42789);
and U46999 (N_46999,N_43881,N_44247);
and U47000 (N_47000,N_44991,N_44194);
xor U47001 (N_47001,N_43974,N_44286);
xor U47002 (N_47002,N_42886,N_44553);
nor U47003 (N_47003,N_42617,N_42775);
nand U47004 (N_47004,N_44695,N_43542);
xnor U47005 (N_47005,N_43200,N_43111);
xnor U47006 (N_47006,N_43062,N_43749);
or U47007 (N_47007,N_43438,N_44972);
nand U47008 (N_47008,N_43446,N_42977);
or U47009 (N_47009,N_44306,N_43310);
xnor U47010 (N_47010,N_43985,N_43584);
and U47011 (N_47011,N_42685,N_43207);
nand U47012 (N_47012,N_43179,N_44878);
and U47013 (N_47013,N_43279,N_44382);
nor U47014 (N_47014,N_43332,N_42646);
nand U47015 (N_47015,N_42598,N_43066);
xnor U47016 (N_47016,N_44240,N_42524);
nand U47017 (N_47017,N_44726,N_42934);
and U47018 (N_47018,N_43035,N_44319);
and U47019 (N_47019,N_43382,N_43063);
or U47020 (N_47020,N_44305,N_43890);
xor U47021 (N_47021,N_44610,N_44450);
and U47022 (N_47022,N_42688,N_42981);
or U47023 (N_47023,N_44288,N_42608);
xor U47024 (N_47024,N_44260,N_43598);
xnor U47025 (N_47025,N_42858,N_42813);
nand U47026 (N_47026,N_42890,N_43599);
or U47027 (N_47027,N_44786,N_44587);
nor U47028 (N_47028,N_44862,N_44220);
nand U47029 (N_47029,N_43722,N_43239);
xnor U47030 (N_47030,N_42631,N_42804);
and U47031 (N_47031,N_43805,N_43789);
and U47032 (N_47032,N_44841,N_43304);
or U47033 (N_47033,N_43401,N_43807);
nor U47034 (N_47034,N_43629,N_43784);
or U47035 (N_47035,N_42851,N_43075);
and U47036 (N_47036,N_44811,N_44680);
and U47037 (N_47037,N_43185,N_44088);
nor U47038 (N_47038,N_43766,N_44657);
nand U47039 (N_47039,N_43548,N_42872);
nand U47040 (N_47040,N_43511,N_44769);
xnor U47041 (N_47041,N_43087,N_43795);
and U47042 (N_47042,N_44083,N_44412);
xnor U47043 (N_47043,N_44941,N_43476);
and U47044 (N_47044,N_44425,N_43987);
xor U47045 (N_47045,N_44682,N_42863);
nor U47046 (N_47046,N_43028,N_43668);
or U47047 (N_47047,N_44742,N_44843);
nand U47048 (N_47048,N_44543,N_42702);
nand U47049 (N_47049,N_44680,N_44386);
or U47050 (N_47050,N_43179,N_44066);
xor U47051 (N_47051,N_44858,N_44641);
nand U47052 (N_47052,N_43277,N_42603);
and U47053 (N_47053,N_43644,N_43139);
nand U47054 (N_47054,N_44981,N_42890);
and U47055 (N_47055,N_44691,N_43213);
nand U47056 (N_47056,N_43419,N_44995);
or U47057 (N_47057,N_43035,N_43065);
and U47058 (N_47058,N_43066,N_44356);
xor U47059 (N_47059,N_43290,N_43379);
nand U47060 (N_47060,N_43629,N_44825);
and U47061 (N_47061,N_43212,N_44920);
nor U47062 (N_47062,N_43694,N_44431);
xnor U47063 (N_47063,N_43554,N_42885);
nand U47064 (N_47064,N_43114,N_43998);
and U47065 (N_47065,N_43500,N_44906);
xor U47066 (N_47066,N_44188,N_43332);
nand U47067 (N_47067,N_42832,N_43863);
nand U47068 (N_47068,N_44792,N_43257);
nor U47069 (N_47069,N_43560,N_42998);
nor U47070 (N_47070,N_43345,N_42603);
and U47071 (N_47071,N_42919,N_43152);
nor U47072 (N_47072,N_43826,N_43243);
nand U47073 (N_47073,N_43373,N_44183);
nor U47074 (N_47074,N_42711,N_43561);
or U47075 (N_47075,N_43981,N_44079);
and U47076 (N_47076,N_44934,N_42567);
xor U47077 (N_47077,N_42597,N_43198);
nand U47078 (N_47078,N_44967,N_44248);
or U47079 (N_47079,N_43105,N_43816);
xor U47080 (N_47080,N_44534,N_44834);
or U47081 (N_47081,N_43661,N_44332);
nand U47082 (N_47082,N_44541,N_44212);
or U47083 (N_47083,N_43135,N_42596);
and U47084 (N_47084,N_43894,N_44463);
nor U47085 (N_47085,N_43576,N_43640);
nand U47086 (N_47086,N_43316,N_44008);
and U47087 (N_47087,N_43389,N_43121);
nor U47088 (N_47088,N_44487,N_42884);
xor U47089 (N_47089,N_44283,N_42841);
nor U47090 (N_47090,N_43868,N_42729);
or U47091 (N_47091,N_43601,N_43812);
or U47092 (N_47092,N_42689,N_43756);
and U47093 (N_47093,N_43153,N_43735);
and U47094 (N_47094,N_43999,N_42808);
and U47095 (N_47095,N_44255,N_42884);
nor U47096 (N_47096,N_44492,N_44984);
nand U47097 (N_47097,N_42529,N_44445);
or U47098 (N_47098,N_44034,N_42849);
nor U47099 (N_47099,N_43430,N_42875);
nand U47100 (N_47100,N_43429,N_44681);
and U47101 (N_47101,N_44524,N_42714);
xor U47102 (N_47102,N_43571,N_42786);
nand U47103 (N_47103,N_44791,N_43788);
xnor U47104 (N_47104,N_42556,N_43032);
nor U47105 (N_47105,N_44446,N_43414);
xnor U47106 (N_47106,N_43841,N_44176);
xnor U47107 (N_47107,N_43165,N_43951);
nand U47108 (N_47108,N_42578,N_43452);
nor U47109 (N_47109,N_44921,N_42914);
xor U47110 (N_47110,N_43282,N_44862);
xnor U47111 (N_47111,N_42868,N_44690);
or U47112 (N_47112,N_42797,N_43349);
nor U47113 (N_47113,N_44605,N_43053);
and U47114 (N_47114,N_44818,N_42726);
or U47115 (N_47115,N_44314,N_42945);
or U47116 (N_47116,N_44743,N_44429);
nor U47117 (N_47117,N_43601,N_43487);
or U47118 (N_47118,N_42619,N_43980);
nand U47119 (N_47119,N_43821,N_43588);
or U47120 (N_47120,N_43389,N_43114);
nand U47121 (N_47121,N_42586,N_43380);
nand U47122 (N_47122,N_43874,N_43744);
xor U47123 (N_47123,N_44500,N_44071);
and U47124 (N_47124,N_44685,N_42787);
and U47125 (N_47125,N_43139,N_43610);
and U47126 (N_47126,N_42518,N_44234);
xnor U47127 (N_47127,N_44194,N_42884);
nand U47128 (N_47128,N_44243,N_43742);
nor U47129 (N_47129,N_42700,N_43077);
nor U47130 (N_47130,N_44347,N_43706);
xnor U47131 (N_47131,N_42909,N_42523);
or U47132 (N_47132,N_43951,N_43538);
or U47133 (N_47133,N_44723,N_43925);
nor U47134 (N_47134,N_44685,N_44139);
xnor U47135 (N_47135,N_44991,N_44081);
or U47136 (N_47136,N_43335,N_43935);
nor U47137 (N_47137,N_43032,N_42956);
or U47138 (N_47138,N_44416,N_42931);
nand U47139 (N_47139,N_43097,N_44714);
nor U47140 (N_47140,N_43409,N_44190);
nand U47141 (N_47141,N_43989,N_44450);
and U47142 (N_47142,N_42994,N_44616);
xor U47143 (N_47143,N_44476,N_44903);
and U47144 (N_47144,N_43206,N_43231);
nor U47145 (N_47145,N_44325,N_44560);
nor U47146 (N_47146,N_42920,N_43823);
nor U47147 (N_47147,N_43456,N_44364);
nand U47148 (N_47148,N_43088,N_43049);
nor U47149 (N_47149,N_44399,N_44657);
xor U47150 (N_47150,N_44444,N_44769);
xnor U47151 (N_47151,N_42916,N_43777);
and U47152 (N_47152,N_44373,N_43315);
or U47153 (N_47153,N_43831,N_43839);
or U47154 (N_47154,N_43417,N_44045);
nand U47155 (N_47155,N_44915,N_43311);
nand U47156 (N_47156,N_44409,N_44938);
and U47157 (N_47157,N_43812,N_43123);
and U47158 (N_47158,N_42735,N_44779);
or U47159 (N_47159,N_43268,N_43388);
and U47160 (N_47160,N_44882,N_43820);
nand U47161 (N_47161,N_44548,N_43692);
xor U47162 (N_47162,N_43086,N_43911);
nand U47163 (N_47163,N_44419,N_44197);
or U47164 (N_47164,N_42906,N_43539);
and U47165 (N_47165,N_42582,N_44614);
or U47166 (N_47166,N_44769,N_44258);
nand U47167 (N_47167,N_43804,N_44171);
xnor U47168 (N_47168,N_44915,N_44525);
or U47169 (N_47169,N_44020,N_43835);
or U47170 (N_47170,N_42707,N_43404);
nor U47171 (N_47171,N_44236,N_44991);
nand U47172 (N_47172,N_44364,N_43503);
or U47173 (N_47173,N_43864,N_44990);
or U47174 (N_47174,N_43842,N_43336);
xnor U47175 (N_47175,N_42756,N_42550);
xnor U47176 (N_47176,N_43744,N_44153);
and U47177 (N_47177,N_42637,N_43603);
and U47178 (N_47178,N_42989,N_43497);
nor U47179 (N_47179,N_42951,N_42994);
or U47180 (N_47180,N_43168,N_43668);
nor U47181 (N_47181,N_42652,N_43713);
nor U47182 (N_47182,N_44360,N_43888);
xnor U47183 (N_47183,N_42877,N_42514);
nor U47184 (N_47184,N_43524,N_44059);
nand U47185 (N_47185,N_43588,N_44035);
nand U47186 (N_47186,N_43403,N_43556);
xnor U47187 (N_47187,N_42532,N_44380);
or U47188 (N_47188,N_43456,N_44854);
xnor U47189 (N_47189,N_44142,N_44500);
or U47190 (N_47190,N_44069,N_44155);
and U47191 (N_47191,N_42526,N_43452);
or U47192 (N_47192,N_44880,N_43168);
xnor U47193 (N_47193,N_44951,N_43152);
nand U47194 (N_47194,N_44632,N_44730);
nor U47195 (N_47195,N_43564,N_44634);
and U47196 (N_47196,N_43605,N_42988);
and U47197 (N_47197,N_44956,N_42840);
nor U47198 (N_47198,N_44977,N_42649);
or U47199 (N_47199,N_43028,N_44899);
or U47200 (N_47200,N_44012,N_44465);
nor U47201 (N_47201,N_43925,N_43192);
nor U47202 (N_47202,N_43358,N_44625);
and U47203 (N_47203,N_43440,N_44482);
nand U47204 (N_47204,N_43038,N_44831);
and U47205 (N_47205,N_44253,N_42764);
xor U47206 (N_47206,N_44894,N_44367);
and U47207 (N_47207,N_43538,N_44381);
or U47208 (N_47208,N_43094,N_44760);
xnor U47209 (N_47209,N_44002,N_42787);
nor U47210 (N_47210,N_44508,N_42961);
nor U47211 (N_47211,N_43227,N_43109);
nor U47212 (N_47212,N_44365,N_42914);
xor U47213 (N_47213,N_44339,N_43230);
or U47214 (N_47214,N_43367,N_44994);
xnor U47215 (N_47215,N_43468,N_43131);
or U47216 (N_47216,N_44693,N_43846);
and U47217 (N_47217,N_42600,N_43711);
and U47218 (N_47218,N_43882,N_43518);
or U47219 (N_47219,N_44575,N_43588);
nand U47220 (N_47220,N_43078,N_44149);
nor U47221 (N_47221,N_44020,N_43679);
or U47222 (N_47222,N_44082,N_42966);
or U47223 (N_47223,N_42853,N_42863);
nand U47224 (N_47224,N_43251,N_44554);
xnor U47225 (N_47225,N_44056,N_44980);
or U47226 (N_47226,N_44753,N_43523);
nor U47227 (N_47227,N_44863,N_43458);
and U47228 (N_47228,N_44415,N_44961);
or U47229 (N_47229,N_42712,N_42873);
nand U47230 (N_47230,N_43029,N_44343);
nand U47231 (N_47231,N_44041,N_44924);
xnor U47232 (N_47232,N_42696,N_42743);
nor U47233 (N_47233,N_44484,N_43715);
and U47234 (N_47234,N_42642,N_44342);
and U47235 (N_47235,N_44342,N_42846);
xor U47236 (N_47236,N_43080,N_44094);
or U47237 (N_47237,N_44888,N_43574);
nor U47238 (N_47238,N_44136,N_44718);
nand U47239 (N_47239,N_43918,N_43039);
or U47240 (N_47240,N_44097,N_43233);
nand U47241 (N_47241,N_42568,N_44927);
nor U47242 (N_47242,N_44013,N_44643);
xor U47243 (N_47243,N_44594,N_43233);
nor U47244 (N_47244,N_42530,N_43453);
or U47245 (N_47245,N_44418,N_42693);
or U47246 (N_47246,N_44297,N_44620);
or U47247 (N_47247,N_43851,N_43590);
nor U47248 (N_47248,N_44301,N_43795);
and U47249 (N_47249,N_44463,N_44930);
nand U47250 (N_47250,N_44557,N_44134);
nand U47251 (N_47251,N_44832,N_44374);
and U47252 (N_47252,N_44995,N_43742);
nor U47253 (N_47253,N_44969,N_44423);
nor U47254 (N_47254,N_43363,N_44421);
nor U47255 (N_47255,N_44482,N_44434);
nand U47256 (N_47256,N_43458,N_42758);
nand U47257 (N_47257,N_44260,N_44945);
nor U47258 (N_47258,N_44227,N_42545);
and U47259 (N_47259,N_44809,N_43563);
and U47260 (N_47260,N_43267,N_43595);
or U47261 (N_47261,N_44888,N_42534);
nor U47262 (N_47262,N_43253,N_43486);
or U47263 (N_47263,N_43641,N_43221);
nand U47264 (N_47264,N_44160,N_43637);
or U47265 (N_47265,N_43304,N_44800);
and U47266 (N_47266,N_44046,N_44680);
or U47267 (N_47267,N_44213,N_43217);
nand U47268 (N_47268,N_42877,N_42665);
nand U47269 (N_47269,N_43537,N_44266);
or U47270 (N_47270,N_43716,N_44922);
nor U47271 (N_47271,N_44401,N_44325);
and U47272 (N_47272,N_42800,N_43539);
or U47273 (N_47273,N_44741,N_44429);
nand U47274 (N_47274,N_43082,N_43003);
nor U47275 (N_47275,N_42962,N_42813);
or U47276 (N_47276,N_43519,N_44229);
nor U47277 (N_47277,N_44951,N_43372);
or U47278 (N_47278,N_44206,N_43192);
nor U47279 (N_47279,N_43276,N_44063);
or U47280 (N_47280,N_42892,N_43494);
or U47281 (N_47281,N_43897,N_42508);
or U47282 (N_47282,N_42812,N_43575);
or U47283 (N_47283,N_43249,N_43799);
nor U47284 (N_47284,N_42892,N_43587);
nand U47285 (N_47285,N_44210,N_43773);
or U47286 (N_47286,N_43447,N_43871);
nor U47287 (N_47287,N_43962,N_42583);
and U47288 (N_47288,N_44142,N_44438);
xor U47289 (N_47289,N_42565,N_44647);
nand U47290 (N_47290,N_44710,N_44761);
and U47291 (N_47291,N_42835,N_44009);
xnor U47292 (N_47292,N_43767,N_43742);
xor U47293 (N_47293,N_44143,N_44042);
xnor U47294 (N_47294,N_44176,N_42607);
xnor U47295 (N_47295,N_43783,N_42892);
nand U47296 (N_47296,N_44752,N_42635);
or U47297 (N_47297,N_43556,N_43619);
nand U47298 (N_47298,N_43015,N_44688);
nand U47299 (N_47299,N_43862,N_44738);
xor U47300 (N_47300,N_44623,N_43625);
or U47301 (N_47301,N_44858,N_44210);
nand U47302 (N_47302,N_44347,N_44420);
nor U47303 (N_47303,N_43889,N_44381);
nor U47304 (N_47304,N_44242,N_43978);
or U47305 (N_47305,N_44028,N_43825);
nor U47306 (N_47306,N_44405,N_44755);
nor U47307 (N_47307,N_43215,N_44069);
and U47308 (N_47308,N_42667,N_44369);
or U47309 (N_47309,N_44770,N_44081);
and U47310 (N_47310,N_44559,N_43422);
and U47311 (N_47311,N_43522,N_44977);
nand U47312 (N_47312,N_43558,N_42639);
nand U47313 (N_47313,N_42671,N_42652);
xor U47314 (N_47314,N_44331,N_44668);
and U47315 (N_47315,N_44936,N_44129);
or U47316 (N_47316,N_42549,N_43946);
nor U47317 (N_47317,N_43892,N_44028);
or U47318 (N_47318,N_43866,N_44951);
xor U47319 (N_47319,N_44653,N_43705);
and U47320 (N_47320,N_43537,N_43249);
xor U47321 (N_47321,N_43319,N_44318);
and U47322 (N_47322,N_44964,N_42984);
or U47323 (N_47323,N_42848,N_44364);
or U47324 (N_47324,N_44770,N_44556);
nand U47325 (N_47325,N_44893,N_43167);
xnor U47326 (N_47326,N_43550,N_42681);
xnor U47327 (N_47327,N_43878,N_43135);
and U47328 (N_47328,N_44662,N_43888);
and U47329 (N_47329,N_42826,N_44219);
or U47330 (N_47330,N_42832,N_43398);
xor U47331 (N_47331,N_43464,N_44546);
or U47332 (N_47332,N_44760,N_42978);
and U47333 (N_47333,N_43439,N_43991);
and U47334 (N_47334,N_43624,N_43124);
nand U47335 (N_47335,N_43855,N_44997);
or U47336 (N_47336,N_44724,N_44905);
nor U47337 (N_47337,N_43301,N_44330);
and U47338 (N_47338,N_42939,N_43976);
nand U47339 (N_47339,N_42624,N_44481);
xnor U47340 (N_47340,N_42995,N_42635);
or U47341 (N_47341,N_42833,N_44141);
or U47342 (N_47342,N_43938,N_42621);
or U47343 (N_47343,N_44850,N_44294);
and U47344 (N_47344,N_44799,N_44035);
xnor U47345 (N_47345,N_44580,N_44739);
nor U47346 (N_47346,N_44310,N_44393);
nor U47347 (N_47347,N_42932,N_44797);
nor U47348 (N_47348,N_43112,N_43550);
or U47349 (N_47349,N_44011,N_44134);
or U47350 (N_47350,N_44210,N_44117);
or U47351 (N_47351,N_42693,N_43373);
and U47352 (N_47352,N_43932,N_44412);
or U47353 (N_47353,N_43033,N_43945);
xnor U47354 (N_47354,N_44219,N_42925);
xor U47355 (N_47355,N_42940,N_43284);
or U47356 (N_47356,N_43530,N_43824);
and U47357 (N_47357,N_42708,N_43128);
nand U47358 (N_47358,N_44321,N_43396);
and U47359 (N_47359,N_42736,N_43236);
and U47360 (N_47360,N_44199,N_43630);
and U47361 (N_47361,N_44023,N_44370);
and U47362 (N_47362,N_43061,N_42888);
nand U47363 (N_47363,N_43571,N_43401);
nor U47364 (N_47364,N_43219,N_44837);
or U47365 (N_47365,N_44771,N_43398);
and U47366 (N_47366,N_42875,N_43094);
nor U47367 (N_47367,N_43915,N_42706);
and U47368 (N_47368,N_43739,N_43530);
and U47369 (N_47369,N_44558,N_43223);
nor U47370 (N_47370,N_43441,N_44067);
xor U47371 (N_47371,N_42898,N_42560);
nor U47372 (N_47372,N_44438,N_44843);
nand U47373 (N_47373,N_42637,N_42714);
and U47374 (N_47374,N_44078,N_42537);
xnor U47375 (N_47375,N_42830,N_43552);
nand U47376 (N_47376,N_44334,N_44358);
nor U47377 (N_47377,N_44886,N_44441);
or U47378 (N_47378,N_43750,N_44093);
xnor U47379 (N_47379,N_44177,N_43748);
nor U47380 (N_47380,N_43694,N_44086);
xnor U47381 (N_47381,N_42846,N_44534);
or U47382 (N_47382,N_43143,N_43634);
nor U47383 (N_47383,N_44161,N_44571);
or U47384 (N_47384,N_43035,N_43708);
xor U47385 (N_47385,N_43318,N_43986);
or U47386 (N_47386,N_44379,N_44461);
and U47387 (N_47387,N_43971,N_43066);
nor U47388 (N_47388,N_44202,N_43776);
xnor U47389 (N_47389,N_43845,N_43005);
and U47390 (N_47390,N_44606,N_44920);
or U47391 (N_47391,N_43796,N_42797);
and U47392 (N_47392,N_43210,N_44964);
xor U47393 (N_47393,N_44092,N_44291);
nand U47394 (N_47394,N_44809,N_42988);
xnor U47395 (N_47395,N_43856,N_42985);
and U47396 (N_47396,N_43764,N_43312);
nand U47397 (N_47397,N_42986,N_44272);
xnor U47398 (N_47398,N_44028,N_43210);
nand U47399 (N_47399,N_44273,N_42512);
nand U47400 (N_47400,N_44516,N_43129);
nand U47401 (N_47401,N_44565,N_44216);
nand U47402 (N_47402,N_43157,N_43874);
or U47403 (N_47403,N_44875,N_44201);
and U47404 (N_47404,N_43832,N_44450);
nor U47405 (N_47405,N_44018,N_44123);
and U47406 (N_47406,N_44079,N_44711);
nand U47407 (N_47407,N_43309,N_43343);
nand U47408 (N_47408,N_44268,N_43008);
nor U47409 (N_47409,N_43545,N_44694);
xor U47410 (N_47410,N_43357,N_44435);
and U47411 (N_47411,N_44570,N_42918);
xor U47412 (N_47412,N_42706,N_43765);
nor U47413 (N_47413,N_42887,N_43438);
or U47414 (N_47414,N_43500,N_42697);
or U47415 (N_47415,N_43458,N_44608);
nand U47416 (N_47416,N_43067,N_43092);
nand U47417 (N_47417,N_44714,N_42935);
nand U47418 (N_47418,N_43539,N_43228);
and U47419 (N_47419,N_44553,N_44409);
xnor U47420 (N_47420,N_42982,N_44670);
and U47421 (N_47421,N_44540,N_43571);
and U47422 (N_47422,N_43264,N_44090);
and U47423 (N_47423,N_43839,N_43457);
nand U47424 (N_47424,N_44365,N_43950);
or U47425 (N_47425,N_43643,N_44588);
and U47426 (N_47426,N_42876,N_44946);
or U47427 (N_47427,N_44776,N_44191);
and U47428 (N_47428,N_43387,N_42877);
nor U47429 (N_47429,N_43353,N_44247);
and U47430 (N_47430,N_43977,N_44997);
and U47431 (N_47431,N_43647,N_44663);
and U47432 (N_47432,N_43506,N_43476);
and U47433 (N_47433,N_43914,N_42679);
or U47434 (N_47434,N_43202,N_42522);
xor U47435 (N_47435,N_44144,N_44789);
nand U47436 (N_47436,N_43014,N_43657);
and U47437 (N_47437,N_43627,N_43634);
nand U47438 (N_47438,N_43001,N_43928);
nand U47439 (N_47439,N_43379,N_44899);
nor U47440 (N_47440,N_44320,N_44002);
or U47441 (N_47441,N_43491,N_42634);
nor U47442 (N_47442,N_42557,N_42843);
or U47443 (N_47443,N_43542,N_44720);
and U47444 (N_47444,N_42795,N_44480);
or U47445 (N_47445,N_43069,N_44609);
and U47446 (N_47446,N_44296,N_43418);
nand U47447 (N_47447,N_43620,N_44581);
or U47448 (N_47448,N_43111,N_44589);
nor U47449 (N_47449,N_42844,N_43627);
nor U47450 (N_47450,N_43494,N_44825);
nor U47451 (N_47451,N_44204,N_42786);
nor U47452 (N_47452,N_42570,N_42904);
and U47453 (N_47453,N_44355,N_42693);
or U47454 (N_47454,N_44104,N_43332);
xnor U47455 (N_47455,N_42865,N_44447);
xnor U47456 (N_47456,N_42569,N_44325);
and U47457 (N_47457,N_43133,N_42516);
nor U47458 (N_47458,N_43827,N_44747);
nand U47459 (N_47459,N_43773,N_43375);
and U47460 (N_47460,N_43877,N_44718);
nor U47461 (N_47461,N_43058,N_44835);
nand U47462 (N_47462,N_43642,N_43662);
nand U47463 (N_47463,N_43511,N_44450);
nand U47464 (N_47464,N_43057,N_42843);
nand U47465 (N_47465,N_43615,N_44464);
or U47466 (N_47466,N_43648,N_43198);
nand U47467 (N_47467,N_44300,N_43602);
or U47468 (N_47468,N_43438,N_44878);
xnor U47469 (N_47469,N_44048,N_43576);
and U47470 (N_47470,N_43481,N_44904);
nand U47471 (N_47471,N_43820,N_43956);
nand U47472 (N_47472,N_44525,N_42744);
nor U47473 (N_47473,N_43940,N_44747);
nor U47474 (N_47474,N_44038,N_43742);
and U47475 (N_47475,N_42976,N_43713);
nor U47476 (N_47476,N_42778,N_42721);
xor U47477 (N_47477,N_42981,N_44173);
xnor U47478 (N_47478,N_44864,N_43996);
xor U47479 (N_47479,N_42986,N_44228);
xnor U47480 (N_47480,N_42770,N_44815);
nor U47481 (N_47481,N_42539,N_44918);
or U47482 (N_47482,N_42612,N_44126);
or U47483 (N_47483,N_44934,N_43288);
nor U47484 (N_47484,N_43170,N_42963);
xnor U47485 (N_47485,N_44455,N_43646);
xor U47486 (N_47486,N_42701,N_42607);
xor U47487 (N_47487,N_44920,N_42644);
xnor U47488 (N_47488,N_43717,N_44493);
or U47489 (N_47489,N_43601,N_44998);
and U47490 (N_47490,N_43973,N_42800);
and U47491 (N_47491,N_43479,N_43953);
or U47492 (N_47492,N_43010,N_44547);
nand U47493 (N_47493,N_44630,N_44963);
and U47494 (N_47494,N_44475,N_43581);
xnor U47495 (N_47495,N_42617,N_43354);
and U47496 (N_47496,N_42662,N_43445);
and U47497 (N_47497,N_44719,N_44781);
nand U47498 (N_47498,N_44910,N_43531);
nor U47499 (N_47499,N_44969,N_42856);
nor U47500 (N_47500,N_45548,N_46478);
xor U47501 (N_47501,N_45091,N_46960);
nor U47502 (N_47502,N_46619,N_46859);
and U47503 (N_47503,N_47446,N_45365);
and U47504 (N_47504,N_47338,N_46028);
nor U47505 (N_47505,N_45845,N_47314);
xnor U47506 (N_47506,N_45562,N_45471);
and U47507 (N_47507,N_47247,N_47017);
nor U47508 (N_47508,N_45516,N_45639);
nand U47509 (N_47509,N_47142,N_46537);
and U47510 (N_47510,N_45820,N_45283);
xnor U47511 (N_47511,N_45224,N_46474);
xor U47512 (N_47512,N_45268,N_45398);
and U47513 (N_47513,N_45729,N_45782);
xnor U47514 (N_47514,N_45744,N_45607);
or U47515 (N_47515,N_46422,N_45446);
nand U47516 (N_47516,N_45602,N_45727);
nand U47517 (N_47517,N_47367,N_46126);
nand U47518 (N_47518,N_45111,N_47465);
and U47519 (N_47519,N_45512,N_45768);
and U47520 (N_47520,N_46773,N_45640);
xor U47521 (N_47521,N_45530,N_45250);
nor U47522 (N_47522,N_47140,N_46276);
nor U47523 (N_47523,N_45711,N_46535);
nand U47524 (N_47524,N_47114,N_47412);
nor U47525 (N_47525,N_46930,N_45348);
and U47526 (N_47526,N_47374,N_46265);
nor U47527 (N_47527,N_45498,N_45067);
and U47528 (N_47528,N_45472,N_46409);
and U47529 (N_47529,N_46944,N_46086);
xor U47530 (N_47530,N_46001,N_45673);
and U47531 (N_47531,N_46708,N_46900);
or U47532 (N_47532,N_47405,N_45217);
or U47533 (N_47533,N_45948,N_46845);
nand U47534 (N_47534,N_46852,N_46136);
or U47535 (N_47535,N_45157,N_46951);
xnor U47536 (N_47536,N_47003,N_47193);
xnor U47537 (N_47537,N_47148,N_46521);
and U47538 (N_47538,N_46074,N_46371);
and U47539 (N_47539,N_47448,N_45231);
nor U47540 (N_47540,N_46687,N_46048);
nor U47541 (N_47541,N_45451,N_45691);
or U47542 (N_47542,N_46005,N_46091);
and U47543 (N_47543,N_47282,N_46143);
xor U47544 (N_47544,N_45865,N_46228);
or U47545 (N_47545,N_45872,N_46090);
nor U47546 (N_47546,N_47369,N_45620);
xor U47547 (N_47547,N_45608,N_45414);
or U47548 (N_47548,N_46479,N_45591);
nor U47549 (N_47549,N_46551,N_46405);
xor U47550 (N_47550,N_47452,N_46331);
and U47551 (N_47551,N_45552,N_47327);
nor U47552 (N_47552,N_46853,N_45368);
or U47553 (N_47553,N_46599,N_46706);
xnor U47554 (N_47554,N_46467,N_46718);
nand U47555 (N_47555,N_46985,N_45925);
nand U47556 (N_47556,N_47104,N_46035);
nand U47557 (N_47557,N_45226,N_45528);
nand U47558 (N_47558,N_45359,N_45965);
xnor U47559 (N_47559,N_47416,N_46233);
nand U47560 (N_47560,N_46080,N_45357);
nand U47561 (N_47561,N_45045,N_46281);
nand U47562 (N_47562,N_45001,N_47007);
nand U47563 (N_47563,N_46895,N_46770);
nand U47564 (N_47564,N_46396,N_46545);
nand U47565 (N_47565,N_47407,N_45382);
xnor U47566 (N_47566,N_45324,N_47313);
or U47567 (N_47567,N_47368,N_46697);
or U47568 (N_47568,N_45893,N_45523);
nor U47569 (N_47569,N_45143,N_47495);
and U47570 (N_47570,N_47281,N_45779);
or U47571 (N_47571,N_46221,N_45606);
nand U47572 (N_47572,N_45173,N_46620);
or U47573 (N_47573,N_46270,N_45052);
nor U47574 (N_47574,N_45982,N_46591);
and U47575 (N_47575,N_45294,N_47294);
and U47576 (N_47576,N_45080,N_45106);
or U47577 (N_47577,N_46686,N_47037);
or U47578 (N_47578,N_45875,N_45669);
or U47579 (N_47579,N_47413,N_46257);
nand U47580 (N_47580,N_45330,N_45578);
nand U47581 (N_47581,N_47402,N_46804);
xor U47582 (N_47582,N_45486,N_45722);
nor U47583 (N_47583,N_45582,N_45439);
xor U47584 (N_47584,N_46273,N_46349);
or U47585 (N_47585,N_46471,N_47418);
xnor U47586 (N_47586,N_45209,N_47083);
nor U47587 (N_47587,N_47320,N_46542);
xnor U47588 (N_47588,N_45637,N_46514);
or U47589 (N_47589,N_46294,N_46056);
and U47590 (N_47590,N_45990,N_46735);
or U47591 (N_47591,N_46592,N_46940);
and U47592 (N_47592,N_45979,N_46446);
and U47593 (N_47593,N_45254,N_45029);
and U47594 (N_47594,N_47190,N_46942);
nand U47595 (N_47595,N_45087,N_46589);
or U47596 (N_47596,N_47437,N_47039);
xor U47597 (N_47597,N_45536,N_47065);
and U47598 (N_47598,N_45424,N_45407);
nand U47599 (N_47599,N_46099,N_45580);
xor U47600 (N_47600,N_46814,N_46500);
nand U47601 (N_47601,N_46746,N_45053);
or U47602 (N_47602,N_45549,N_45302);
nand U47603 (N_47603,N_46555,N_45935);
nand U47604 (N_47604,N_45553,N_47173);
xnor U47605 (N_47605,N_45886,N_46047);
or U47606 (N_47606,N_46936,N_45487);
and U47607 (N_47607,N_47122,N_45346);
or U47608 (N_47608,N_45454,N_45649);
or U47609 (N_47609,N_45186,N_46284);
or U47610 (N_47610,N_45320,N_45629);
xor U47611 (N_47611,N_46308,N_46565);
xnor U47612 (N_47612,N_46106,N_46890);
nor U47613 (N_47613,N_46886,N_46849);
xnor U47614 (N_47614,N_46206,N_46782);
nand U47615 (N_47615,N_45885,N_46881);
or U47616 (N_47616,N_47260,N_47225);
nor U47617 (N_47617,N_45958,N_46470);
or U47618 (N_47618,N_45137,N_45650);
nand U47619 (N_47619,N_46524,N_46484);
xor U47620 (N_47620,N_46832,N_46953);
nor U47621 (N_47621,N_46963,N_45815);
nor U47622 (N_47622,N_45912,N_46650);
nand U47623 (N_47623,N_46200,N_47154);
nand U47624 (N_47624,N_46375,N_45785);
nand U47625 (N_47625,N_45969,N_46462);
and U47626 (N_47626,N_46546,N_47274);
xor U47627 (N_47627,N_45437,N_45689);
nor U47628 (N_47628,N_45311,N_46637);
and U47629 (N_47629,N_47363,N_46178);
and U47630 (N_47630,N_45394,N_45643);
or U47631 (N_47631,N_45120,N_46626);
xor U47632 (N_47632,N_45298,N_47490);
nand U47633 (N_47633,N_45460,N_46410);
or U47634 (N_47634,N_47047,N_47441);
or U47635 (N_47635,N_46863,N_47426);
xor U47636 (N_47636,N_46938,N_47400);
or U47637 (N_47637,N_46865,N_45638);
xor U47638 (N_47638,N_45550,N_45896);
xnor U47639 (N_47639,N_46914,N_46887);
and U47640 (N_47640,N_45203,N_46125);
or U47641 (N_47641,N_46685,N_46185);
and U47642 (N_47642,N_46986,N_46646);
xnor U47643 (N_47643,N_47155,N_45763);
and U47644 (N_47644,N_47172,N_45725);
or U47645 (N_47645,N_45301,N_45757);
nand U47646 (N_47646,N_46093,N_45849);
and U47647 (N_47647,N_45628,N_45293);
xor U47648 (N_47648,N_47290,N_47415);
nand U47649 (N_47649,N_45573,N_45568);
nor U47650 (N_47650,N_45028,N_45430);
xor U47651 (N_47651,N_46290,N_45064);
nand U47652 (N_47652,N_45975,N_46385);
xnor U47653 (N_47653,N_46825,N_46039);
or U47654 (N_47654,N_45808,N_45743);
or U47655 (N_47655,N_47326,N_46651);
nand U47656 (N_47656,N_45450,N_45477);
nor U47657 (N_47657,N_46867,N_47456);
or U47658 (N_47658,N_45289,N_46073);
or U47659 (N_47659,N_46869,N_47386);
nor U47660 (N_47660,N_47224,N_45739);
and U47661 (N_47661,N_46128,N_47271);
nand U47662 (N_47662,N_46821,N_45118);
nand U47663 (N_47663,N_46883,N_46991);
nor U47664 (N_47664,N_47138,N_47470);
nand U47665 (N_47665,N_46884,N_46016);
and U47666 (N_47666,N_47477,N_46495);
xor U47667 (N_47667,N_45144,N_45513);
and U47668 (N_47668,N_45208,N_46598);
or U47669 (N_47669,N_46754,N_46292);
nor U47670 (N_47670,N_46282,N_45465);
nand U47671 (N_47671,N_46823,N_46417);
or U47672 (N_47672,N_46232,N_46088);
nand U47673 (N_47673,N_47417,N_46952);
and U47674 (N_47674,N_47375,N_46252);
nand U47675 (N_47675,N_47161,N_46267);
nand U47676 (N_47676,N_46360,N_46915);
nor U47677 (N_47677,N_45705,N_47000);
nor U47678 (N_47678,N_47088,N_45981);
or U47679 (N_47679,N_47031,N_47250);
and U47680 (N_47680,N_46269,N_47236);
and U47681 (N_47681,N_45720,N_45488);
and U47682 (N_47682,N_45404,N_45280);
nand U47683 (N_47683,N_46400,N_46922);
and U47684 (N_47684,N_46286,N_47279);
and U47685 (N_47685,N_45184,N_45692);
nor U47686 (N_47686,N_46486,N_47177);
and U47687 (N_47687,N_45766,N_46969);
and U47688 (N_47688,N_45764,N_46764);
nand U47689 (N_47689,N_45244,N_45018);
nor U47690 (N_47690,N_47466,N_46085);
nand U47691 (N_47691,N_47382,N_46731);
or U47692 (N_47692,N_47340,N_47066);
and U47693 (N_47693,N_45006,N_46289);
xnor U47694 (N_47694,N_46601,N_45119);
xor U47695 (N_47695,N_46447,N_47032);
or U47696 (N_47696,N_46435,N_45895);
nand U47697 (N_47697,N_45961,N_46775);
nand U47698 (N_47698,N_46729,N_45457);
xor U47699 (N_47699,N_45461,N_46391);
and U47700 (N_47700,N_45211,N_46006);
nor U47701 (N_47701,N_45690,N_46095);
or U47702 (N_47702,N_47178,N_46215);
xnor U47703 (N_47703,N_45155,N_45570);
xnor U47704 (N_47704,N_45599,N_45964);
nor U47705 (N_47705,N_47199,N_45574);
or U47706 (N_47706,N_46184,N_45632);
nand U47707 (N_47707,N_46612,N_47233);
and U47708 (N_47708,N_45993,N_46777);
and U47709 (N_47709,N_45219,N_46054);
or U47710 (N_47710,N_47409,N_46694);
nor U47711 (N_47711,N_46235,N_47043);
nand U47712 (N_47712,N_46947,N_45834);
nor U47713 (N_47713,N_46576,N_45288);
xor U47714 (N_47714,N_47480,N_45222);
nor U47715 (N_47715,N_47054,N_47112);
nor U47716 (N_47716,N_46330,N_46012);
xor U47717 (N_47717,N_46161,N_47115);
and U47718 (N_47718,N_45112,N_46424);
nand U47719 (N_47719,N_46496,N_47468);
nand U47720 (N_47720,N_45332,N_45651);
nand U47721 (N_47721,N_45532,N_45827);
xor U47722 (N_47722,N_45862,N_46581);
and U47723 (N_47723,N_45544,N_45127);
nand U47724 (N_47724,N_46656,N_47401);
nand U47725 (N_47725,N_45376,N_45065);
nor U47726 (N_47726,N_46271,N_45710);
xor U47727 (N_47727,N_45468,N_46137);
nor U47728 (N_47728,N_45076,N_46045);
and U47729 (N_47729,N_45585,N_46982);
nor U47730 (N_47730,N_45493,N_46748);
nand U47731 (N_47731,N_45277,N_45115);
and U47732 (N_47732,N_45889,N_45243);
nor U47733 (N_47733,N_46266,N_46856);
nand U47734 (N_47734,N_46665,N_47451);
or U47735 (N_47735,N_46031,N_45605);
nand U47736 (N_47736,N_46188,N_45342);
and U47737 (N_47737,N_45917,N_45178);
and U47738 (N_47738,N_46209,N_45387);
nand U47739 (N_47739,N_47280,N_45462);
xnor U47740 (N_47740,N_45588,N_47149);
nor U47741 (N_47741,N_47385,N_46477);
xor U47742 (N_47742,N_46783,N_45802);
xor U47743 (N_47743,N_46212,N_45467);
nor U47744 (N_47744,N_47309,N_46318);
or U47745 (N_47745,N_45929,N_45617);
or U47746 (N_47746,N_45646,N_46354);
nand U47747 (N_47747,N_45829,N_47158);
and U47748 (N_47748,N_45547,N_47038);
and U47749 (N_47749,N_47316,N_47258);
nor U47750 (N_47750,N_46350,N_45379);
nor U47751 (N_47751,N_45242,N_45494);
xnor U47752 (N_47752,N_45049,N_46324);
xor U47753 (N_47753,N_45923,N_45936);
xnor U47754 (N_47754,N_46536,N_45726);
nand U47755 (N_47755,N_45305,N_46101);
xor U47756 (N_47756,N_45631,N_45022);
nor U47757 (N_47757,N_47317,N_45758);
xor U47758 (N_47758,N_47208,N_47132);
xor U47759 (N_47759,N_47145,N_45682);
xnor U47760 (N_47760,N_47336,N_46568);
nor U47761 (N_47761,N_47330,N_45125);
nand U47762 (N_47762,N_46459,N_45527);
and U47763 (N_47763,N_46710,N_45977);
xor U47764 (N_47764,N_46245,N_46672);
and U47765 (N_47765,N_46113,N_46690);
nor U47766 (N_47766,N_45662,N_47455);
or U47767 (N_47767,N_45113,N_46872);
or U47768 (N_47768,N_46961,N_45777);
or U47769 (N_47769,N_47086,N_45275);
and U47770 (N_47770,N_45361,N_46629);
xnor U47771 (N_47771,N_46109,N_47435);
nor U47772 (N_47772,N_47135,N_46339);
nor U47773 (N_47773,N_45432,N_45499);
xnor U47774 (N_47774,N_47453,N_46874);
nand U47775 (N_47775,N_46122,N_46653);
nand U47776 (N_47776,N_45678,N_47079);
xor U47777 (N_47777,N_45040,N_47443);
nor U47778 (N_47778,N_46489,N_46140);
xnor U47779 (N_47779,N_46858,N_45563);
xor U47780 (N_47780,N_46671,N_45199);
nor U47781 (N_47781,N_45378,N_45851);
nand U47782 (N_47782,N_46485,N_46190);
nand U47783 (N_47783,N_45321,N_45482);
xor U47784 (N_47784,N_45952,N_46624);
and U47785 (N_47785,N_45017,N_45656);
nand U47786 (N_47786,N_46450,N_45273);
or U47787 (N_47787,N_47075,N_45401);
or U47788 (N_47788,N_47109,N_47085);
xnor U47789 (N_47789,N_45101,N_46377);
nand U47790 (N_47790,N_45783,N_46306);
nand U47791 (N_47791,N_46901,N_45962);
nor U47792 (N_47792,N_47182,N_47144);
nor U47793 (N_47793,N_45138,N_45162);
nor U47794 (N_47794,N_46844,N_46413);
xor U47795 (N_47795,N_46104,N_47380);
xnor U47796 (N_47796,N_45240,N_45919);
nand U47797 (N_47797,N_47276,N_45481);
and U47798 (N_47798,N_47439,N_46483);
nor U47799 (N_47799,N_47323,N_47168);
xnor U47800 (N_47800,N_46896,N_47100);
or U47801 (N_47801,N_46837,N_46611);
nand U47802 (N_47802,N_46750,N_45931);
nand U47803 (N_47803,N_47218,N_46558);
nand U47804 (N_47804,N_46813,N_46995);
and U47805 (N_47805,N_46970,N_45519);
xor U47806 (N_47806,N_47183,N_46302);
nor U47807 (N_47807,N_45391,N_46443);
xor U47808 (N_47808,N_46441,N_45041);
nand U47809 (N_47809,N_45025,N_45676);
or U47810 (N_47810,N_45652,N_46795);
nand U47811 (N_47811,N_46150,N_46716);
and U47812 (N_47812,N_45237,N_46526);
or U47813 (N_47813,N_45295,N_45927);
or U47814 (N_47814,N_47248,N_47061);
or U47815 (N_47815,N_46255,N_45042);
xnor U47816 (N_47816,N_45433,N_47227);
and U47817 (N_47817,N_47176,N_45255);
nor U47818 (N_47818,N_45071,N_46147);
or U47819 (N_47819,N_47034,N_46034);
xor U47820 (N_47820,N_45205,N_45134);
nor U47821 (N_47821,N_47259,N_47345);
nand U47822 (N_47822,N_45469,N_45507);
or U47823 (N_47823,N_46374,N_45223);
nor U47824 (N_47824,N_45371,N_45664);
and U47825 (N_47825,N_46341,N_47378);
or U47826 (N_47826,N_45846,N_46657);
or U47827 (N_47827,N_47499,N_45239);
xnor U47828 (N_47828,N_45510,N_46550);
or U47829 (N_47829,N_45296,N_47201);
or U47830 (N_47830,N_47342,N_47344);
nor U47831 (N_47831,N_45759,N_46022);
or U47832 (N_47832,N_45716,N_45836);
nor U47833 (N_47833,N_46638,N_47261);
xnor U47834 (N_47834,N_45201,N_45306);
and U47835 (N_47835,N_47243,N_47487);
nand U47836 (N_47836,N_45683,N_46246);
or U47837 (N_47837,N_47133,N_47389);
nand U47838 (N_47838,N_47460,N_46802);
nand U47839 (N_47839,N_46340,N_45164);
nor U47840 (N_47840,N_45667,N_46510);
or U47841 (N_47841,N_46593,N_47373);
or U47842 (N_47842,N_45480,N_47063);
or U47843 (N_47843,N_46162,N_45350);
xor U47844 (N_47844,N_47381,N_45934);
nand U47845 (N_47845,N_45983,N_46300);
xor U47846 (N_47846,N_45470,N_47228);
nor U47847 (N_47847,N_45136,N_45695);
nor U47848 (N_47848,N_46287,N_47312);
xnor U47849 (N_47849,N_46024,N_46158);
and U47850 (N_47850,N_45366,N_46427);
nand U47851 (N_47851,N_46328,N_46538);
xor U47852 (N_47852,N_46418,N_47223);
nand U47853 (N_47853,N_46401,N_45791);
xnor U47854 (N_47854,N_46351,N_45781);
xor U47855 (N_47855,N_45741,N_46717);
or U47856 (N_47856,N_46641,N_46316);
xnor U47857 (N_47857,N_46967,N_46168);
nand U47858 (N_47858,N_46700,N_46303);
nand U47859 (N_47859,N_45644,N_47289);
xnor U47860 (N_47860,N_45438,N_45908);
and U47861 (N_47861,N_46705,N_45543);
nor U47862 (N_47862,N_46841,N_45245);
xnor U47863 (N_47863,N_46812,N_45175);
nor U47864 (N_47864,N_46571,N_45755);
xor U47865 (N_47865,N_46298,N_45973);
nand U47866 (N_47866,N_45621,N_46149);
xor U47867 (N_47867,N_46127,N_45060);
xnor U47868 (N_47868,N_45150,N_46138);
or U47869 (N_47869,N_45110,N_46518);
or U47870 (N_47870,N_45329,N_46414);
nand U47871 (N_47871,N_45787,N_45614);
or U47872 (N_47872,N_46684,N_45776);
and U47873 (N_47873,N_46451,N_45007);
nor U47874 (N_47874,N_47220,N_45009);
or U47875 (N_47875,N_46166,N_45166);
xnor U47876 (N_47876,N_45884,N_45408);
or U47877 (N_47877,N_45730,N_45707);
and U47878 (N_47878,N_45215,N_45954);
nand U47879 (N_47879,N_47348,N_45084);
or U47880 (N_47880,N_46893,N_45020);
or U47881 (N_47881,N_45805,N_46440);
and U47882 (N_47882,N_45586,N_47226);
xnor U47883 (N_47883,N_47077,N_46752);
nand U47884 (N_47884,N_45323,N_45309);
and U47885 (N_47885,N_47048,N_46507);
nor U47886 (N_47886,N_46636,N_46481);
nand U47887 (N_47887,N_46909,N_46789);
or U47888 (N_47888,N_45626,N_46709);
and U47889 (N_47889,N_46030,N_46491);
and U47890 (N_47890,N_45272,N_46038);
nand U47891 (N_47891,N_46046,N_46213);
nand U47892 (N_47892,N_47153,N_46996);
nor U47893 (N_47893,N_46283,N_46457);
nor U47894 (N_47894,N_45904,N_45714);
xnor U47895 (N_47895,N_46562,N_45967);
nor U47896 (N_47896,N_46381,N_45444);
or U47897 (N_47897,N_46019,N_47440);
or U47898 (N_47898,N_45390,N_45657);
nor U47899 (N_47899,N_47050,N_45515);
xnor U47900 (N_47900,N_45225,N_47310);
or U47901 (N_47901,N_45595,N_45955);
nand U47902 (N_47902,N_45600,N_45396);
xor U47903 (N_47903,N_45126,N_46627);
and U47904 (N_47904,N_47181,N_46042);
and U47905 (N_47905,N_46192,N_45476);
nand U47906 (N_47906,N_47496,N_46923);
or U47907 (N_47907,N_46337,N_46103);
xor U47908 (N_47908,N_46299,N_46556);
nor U47909 (N_47909,N_47377,N_46756);
and U47910 (N_47910,N_45998,N_46726);
nand U47911 (N_47911,N_47163,N_46439);
nand U47912 (N_47912,N_46766,N_45419);
xnor U47913 (N_47913,N_45442,N_45859);
nor U47914 (N_47914,N_46943,N_47303);
nand U47915 (N_47915,N_45381,N_45284);
and U47916 (N_47916,N_45459,N_45016);
xnor U47917 (N_47917,N_45317,N_47307);
and U47918 (N_47918,N_45957,N_45310);
xor U47919 (N_47919,N_46956,N_46021);
and U47920 (N_47920,N_46359,N_47484);
or U47921 (N_47921,N_47053,N_45956);
or U47922 (N_47922,N_45502,N_46583);
xnor U47923 (N_47923,N_46892,N_45098);
or U47924 (N_47924,N_45590,N_45351);
and U47925 (N_47925,N_45539,N_47391);
xor U47926 (N_47926,N_46421,N_46226);
xor U47927 (N_47927,N_45655,N_45848);
or U47928 (N_47928,N_47205,N_46513);
nand U47929 (N_47929,N_46151,N_45878);
nand U47930 (N_47930,N_47390,N_47301);
and U47931 (N_47931,N_45423,N_46553);
nand U47932 (N_47932,N_45061,N_46714);
nand U47933 (N_47933,N_46987,N_45044);
and U47934 (N_47934,N_45107,N_45630);
and U47935 (N_47935,N_46724,N_46179);
nand U47936 (N_47936,N_46933,N_47213);
nor U47937 (N_47937,N_45821,N_47014);
nor U47938 (N_47938,N_46262,N_45503);
nor U47939 (N_47939,N_45531,N_46403);
nor U47940 (N_47940,N_46688,N_46208);
and U47941 (N_47941,N_45760,N_47489);
or U47942 (N_47942,N_46368,N_45596);
nand U47943 (N_47943,N_45731,N_45256);
xor U47944 (N_47944,N_45870,N_46240);
nand U47945 (N_47945,N_45267,N_45835);
or U47946 (N_47946,N_45723,N_46975);
xor U47947 (N_47947,N_47025,N_45194);
nand U47948 (N_47948,N_46668,N_45496);
and U47949 (N_47949,N_46224,N_47318);
and U47950 (N_47950,N_46805,N_46345);
nand U47951 (N_47951,N_46383,N_45943);
nand U47952 (N_47952,N_47497,N_45997);
nor U47953 (N_47953,N_45816,N_47333);
nor U47954 (N_47954,N_45218,N_46954);
nor U47955 (N_47955,N_46683,N_45202);
xnor U47956 (N_47956,N_45790,N_46058);
or U47957 (N_47957,N_45609,N_46305);
nor U47958 (N_47958,N_47068,N_46721);
xnor U47959 (N_47959,N_47240,N_46380);
and U47960 (N_47960,N_45828,N_45319);
nand U47961 (N_47961,N_45322,N_46701);
or U47962 (N_47962,N_45123,N_45039);
nor U47963 (N_47963,N_47089,N_45855);
xor U47964 (N_47964,N_47215,N_46755);
or U47965 (N_47965,N_46788,N_46780);
xnor U47966 (N_47966,N_46608,N_47387);
and U47967 (N_47967,N_47353,N_45535);
nand U47968 (N_47968,N_46156,N_46616);
and U47969 (N_47969,N_45135,N_46473);
nor U47970 (N_47970,N_47354,N_46769);
xnor U47971 (N_47971,N_45734,N_45994);
nand U47972 (N_47972,N_46402,N_46512);
xnor U47973 (N_47973,N_45565,N_46904);
or U47974 (N_47974,N_47410,N_46965);
nor U47975 (N_47975,N_45385,N_45556);
xor U47976 (N_47976,N_45648,N_45132);
and U47977 (N_47977,N_46250,N_45452);
nand U47978 (N_47978,N_46355,N_46171);
nor U47979 (N_47979,N_47001,N_47212);
nand U47980 (N_47980,N_45762,N_45765);
nor U47981 (N_47981,N_47403,N_47167);
nor U47982 (N_47982,N_45699,N_46927);
xor U47983 (N_47983,N_45625,N_47267);
and U47984 (N_47984,N_45684,N_46395);
xnor U47985 (N_47985,N_45511,N_45894);
nand U47986 (N_47986,N_47319,N_46920);
nand U47987 (N_47987,N_46154,N_47095);
nand U47988 (N_47988,N_45117,N_45745);
or U47989 (N_47989,N_46310,N_45265);
nor U47990 (N_47990,N_45004,N_47408);
or U47991 (N_47991,N_47450,N_45304);
xnor U47992 (N_47992,N_46864,N_45197);
or U47993 (N_47993,N_46875,N_45924);
or U47994 (N_47994,N_47244,N_45313);
nor U47995 (N_47995,N_45524,N_45794);
nand U47996 (N_47996,N_46198,N_45561);
nand U47997 (N_47997,N_47036,N_46811);
or U47998 (N_47998,N_47196,N_46807);
nor U47999 (N_47999,N_46816,N_46993);
and U48000 (N_48000,N_46772,N_46519);
xor U48001 (N_48001,N_45073,N_47099);
xnor U48002 (N_48002,N_47019,N_46587);
nor U48003 (N_48003,N_45772,N_45140);
nand U48004 (N_48004,N_45784,N_45393);
nand U48005 (N_48005,N_45478,N_45636);
nor U48006 (N_48006,N_45702,N_47081);
xnor U48007 (N_48007,N_45907,N_45221);
and U48008 (N_48008,N_47297,N_47346);
or U48009 (N_48009,N_46361,N_46574);
nor U48010 (N_48010,N_46382,N_46707);
nand U48011 (N_48011,N_46373,N_47306);
nand U48012 (N_48012,N_45857,N_46370);
xor U48013 (N_48013,N_46399,N_45789);
and U48014 (N_48014,N_45069,N_47252);
nor U48015 (N_48015,N_45837,N_45403);
nand U48016 (N_48016,N_46389,N_46720);
xor U48017 (N_48017,N_45397,N_45594);
nor U48018 (N_48018,N_45405,N_47355);
xnor U48019 (N_48019,N_46606,N_45798);
or U48020 (N_48020,N_45058,N_46843);
and U48021 (N_48021,N_45021,N_46984);
or U48022 (N_48022,N_45034,N_47082);
nand U48023 (N_48023,N_45160,N_46977);
nand U48024 (N_48024,N_47268,N_46958);
xnor U48025 (N_48025,N_46488,N_46704);
xor U48026 (N_48026,N_45083,N_46681);
xor U48027 (N_48027,N_45700,N_46817);
nand U48028 (N_48028,N_46026,N_45863);
nor U48029 (N_48029,N_45756,N_47479);
or U48030 (N_48030,N_46411,N_46695);
xor U48031 (N_48031,N_46741,N_45966);
nand U48032 (N_48032,N_47438,N_46135);
and U48033 (N_48033,N_45501,N_46068);
xor U48034 (N_48034,N_47383,N_45560);
nand U48035 (N_48035,N_45603,N_45104);
and U48036 (N_48036,N_47308,N_45139);
nand U48037 (N_48037,N_46165,N_45773);
and U48038 (N_48038,N_45661,N_46830);
nor U48039 (N_48039,N_45939,N_45786);
nor U48040 (N_48040,N_46288,N_46220);
nand U48041 (N_48041,N_46888,N_46326);
xor U48042 (N_48042,N_45068,N_45168);
nand U48043 (N_48043,N_46464,N_46738);
nor U48044 (N_48044,N_45417,N_45897);
and U48045 (N_48045,N_46529,N_46312);
nor U48046 (N_48046,N_47008,N_45075);
nor U48047 (N_48047,N_45372,N_45338);
or U48048 (N_48048,N_45458,N_47364);
nor U48049 (N_48049,N_46734,N_46761);
and U48050 (N_48050,N_46971,N_46670);
and U48051 (N_48051,N_45362,N_47207);
xor U48052 (N_48052,N_45900,N_46736);
nand U48053 (N_48053,N_46279,N_47291);
nand U48054 (N_48054,N_45873,N_46949);
nor U48055 (N_48055,N_46669,N_45987);
or U48056 (N_48056,N_46549,N_46673);
xor U48057 (N_48057,N_46013,N_47206);
xnor U48058 (N_48058,N_45384,N_45995);
and U48059 (N_48059,N_45169,N_47349);
xnor U48060 (N_48060,N_47249,N_45592);
nand U48061 (N_48061,N_46876,N_46263);
or U48062 (N_48062,N_45945,N_45860);
xor U48063 (N_48063,N_45627,N_46586);
and U48064 (N_48064,N_46087,N_46515);
nor U48065 (N_48065,N_46251,N_46494);
nor U48066 (N_48066,N_45569,N_46384);
nand U48067 (N_48067,N_45063,N_46108);
and U48068 (N_48068,N_46652,N_46862);
nor U48069 (N_48069,N_46141,N_46067);
nor U48070 (N_48070,N_46527,N_47137);
or U48071 (N_48071,N_45999,N_47266);
and U48072 (N_48072,N_45497,N_47094);
and U48073 (N_48073,N_45694,N_45074);
or U48074 (N_48074,N_47339,N_46778);
nor U48075 (N_48075,N_45316,N_47445);
xnor U48076 (N_48076,N_45559,N_47431);
and U48077 (N_48077,N_46541,N_46723);
nor U48078 (N_48078,N_45048,N_46544);
and U48079 (N_48079,N_46454,N_45748);
xnor U48080 (N_48080,N_47035,N_46719);
nor U48081 (N_48081,N_46195,N_47130);
or U48082 (N_48082,N_47126,N_47098);
or U48083 (N_48083,N_46857,N_47253);
nand U48084 (N_48084,N_46990,N_45434);
nand U48085 (N_48085,N_45866,N_45318);
xor U48086 (N_48086,N_45858,N_46819);
xnor U48087 (N_48087,N_46703,N_47092);
and U48088 (N_48088,N_46966,N_46057);
or U48089 (N_48089,N_45207,N_45619);
nor U48090 (N_48090,N_46835,N_47395);
or U48091 (N_48091,N_45426,N_45261);
xor U48092 (N_48092,N_46560,N_47096);
nand U48093 (N_48093,N_45431,N_46666);
nand U48094 (N_48094,N_47419,N_45367);
nor U48095 (N_48095,N_45830,N_45095);
or U48096 (N_48096,N_45133,N_47476);
nand U48097 (N_48097,N_47049,N_47129);
nand U48098 (N_48098,N_46912,N_46983);
or U48099 (N_48099,N_45797,N_47072);
nand U48100 (N_48100,N_45970,N_46428);
xor U48101 (N_48101,N_45266,N_47146);
nor U48102 (N_48102,N_46277,N_45879);
and U48103 (N_48103,N_45057,N_45986);
nor U48104 (N_48104,N_46745,N_45803);
nand U48105 (N_48105,N_45300,N_46335);
nand U48106 (N_48106,N_45555,N_45747);
or U48107 (N_48107,N_45011,N_45066);
nor U48108 (N_48108,N_47420,N_47481);
and U48109 (N_48109,N_45809,N_46398);
nand U48110 (N_48110,N_47045,N_46051);
xor U48111 (N_48111,N_46522,N_45712);
xor U48112 (N_48112,N_46787,N_45200);
nor U48113 (N_48113,N_46498,N_47069);
xor U48114 (N_48114,N_45492,N_46531);
and U48115 (N_48115,N_46050,N_46274);
xnor U48116 (N_48116,N_46010,N_46580);
or U48117 (N_48117,N_45767,N_45593);
nand U48118 (N_48118,N_45930,N_46548);
and U48119 (N_48119,N_45370,N_45788);
xor U48120 (N_48120,N_45171,N_45415);
nand U48121 (N_48121,N_46800,N_45941);
nand U48122 (N_48122,N_45703,N_46032);
nand U48123 (N_48123,N_45037,N_45308);
nand U48124 (N_48124,N_45754,N_45704);
nor U48125 (N_48125,N_46183,N_45911);
nor U48126 (N_48126,N_45416,N_46501);
xnor U48127 (N_48127,N_46357,N_46182);
and U48128 (N_48128,N_47027,N_46419);
nand U48129 (N_48129,N_47493,N_45564);
nand U48130 (N_48130,N_47234,N_46979);
nor U48131 (N_48131,N_45109,N_45545);
nor U48132 (N_48132,N_46831,N_46810);
or U48133 (N_48133,N_45072,N_47337);
nor U48134 (N_48134,N_47051,N_46196);
nand U48135 (N_48135,N_47262,N_46539);
or U48136 (N_48136,N_45914,N_46663);
xor U48137 (N_48137,N_45024,N_46177);
nor U48138 (N_48138,N_46121,N_45634);
or U48139 (N_48139,N_45947,N_45474);
nand U48140 (N_48140,N_47322,N_47341);
nand U48141 (N_48141,N_47189,N_45642);
nand U48142 (N_48142,N_46790,N_46758);
nand U48143 (N_48143,N_45811,N_45336);
and U48144 (N_48144,N_45279,N_46442);
nand U48145 (N_48145,N_45801,N_46379);
nor U48146 (N_48146,N_45435,N_45206);
and U48147 (N_48147,N_45780,N_46071);
nor U48148 (N_48148,N_45891,N_47270);
or U48149 (N_48149,N_46497,N_46827);
and U48150 (N_48150,N_45228,N_45709);
nand U48151 (N_48151,N_46160,N_46855);
nand U48152 (N_48152,N_45005,N_45428);
xnor U48153 (N_48153,N_46452,N_47231);
nand U48154 (N_48154,N_46793,N_45395);
xnor U48155 (N_48155,N_45951,N_46517);
nand U48156 (N_48156,N_45546,N_47239);
xnor U48157 (N_48157,N_46002,N_45932);
or U48158 (N_48158,N_46083,N_46230);
xnor U48159 (N_48159,N_45092,N_46333);
or U48160 (N_48160,N_45877,N_45571);
or U48161 (N_48161,N_46948,N_46076);
and U48162 (N_48162,N_47120,N_46490);
or U48163 (N_48163,N_45033,N_46625);
or U48164 (N_48164,N_46540,N_46897);
and U48165 (N_48165,N_45185,N_45421);
xnor U48166 (N_48166,N_46674,N_47087);
nor U48167 (N_48167,N_45070,N_45946);
nor U48168 (N_48168,N_47216,N_47472);
nor U48169 (N_48169,N_47255,N_46765);
xnor U48170 (N_48170,N_46244,N_45713);
xnor U48171 (N_48171,N_46343,N_46794);
nand U48172 (N_48172,N_47214,N_46332);
or U48173 (N_48173,N_46989,N_46603);
nand U48174 (N_48174,N_45575,N_45752);
xor U48175 (N_48175,N_45436,N_45286);
and U48176 (N_48176,N_47191,N_45291);
xnor U48177 (N_48177,N_46623,N_46590);
nor U48178 (N_48178,N_47041,N_45750);
and U48179 (N_48179,N_46009,N_46771);
or U48180 (N_48180,N_45094,N_46430);
or U48181 (N_48181,N_46415,N_45213);
nor U48182 (N_48182,N_46585,N_47422);
xor U48183 (N_48183,N_45441,N_45715);
and U48184 (N_48184,N_46348,N_45842);
nor U48185 (N_48185,N_45096,N_46436);
and U48186 (N_48186,N_45799,N_47024);
and U48187 (N_48187,N_46268,N_45824);
xnor U48188 (N_48188,N_45718,N_46469);
nand U48189 (N_48189,N_45950,N_45910);
xnor U48190 (N_48190,N_45191,N_45409);
nand U48191 (N_48191,N_46509,N_46199);
nand U48192 (N_48192,N_45996,N_45013);
and U48193 (N_48193,N_47232,N_46614);
or U48194 (N_48194,N_46078,N_45183);
or U48195 (N_48195,N_45447,N_45121);
nor U48196 (N_48196,N_47067,N_47180);
nand U48197 (N_48197,N_47358,N_47021);
nor U48198 (N_48198,N_45737,N_45898);
nor U48199 (N_48199,N_47474,N_47221);
and U48200 (N_48200,N_45116,N_46014);
nor U48201 (N_48201,N_46525,N_46163);
nor U48202 (N_48202,N_46607,N_47332);
and U48203 (N_48203,N_47052,N_45509);
nand U48204 (N_48204,N_47288,N_46313);
or U48205 (N_48205,N_45838,N_46846);
and U48206 (N_48206,N_46564,N_46075);
nand U48207 (N_48207,N_46004,N_45972);
or U48208 (N_48208,N_45679,N_45082);
nor U48209 (N_48209,N_46202,N_46826);
nor U48210 (N_48210,N_45274,N_46878);
xor U48211 (N_48211,N_46640,N_45775);
and U48212 (N_48212,N_45012,N_46219);
xor U48213 (N_48213,N_46552,N_46079);
xor U48214 (N_48214,N_45352,N_45774);
nand U48215 (N_48215,N_46997,N_46908);
or U48216 (N_48216,N_45864,N_47179);
or U48217 (N_48217,N_45355,N_47238);
nand U48218 (N_48218,N_45665,N_45325);
xor U48219 (N_48219,N_46820,N_46115);
or U48220 (N_48220,N_46066,N_47195);
or U48221 (N_48221,N_47028,N_46466);
nand U48222 (N_48222,N_46836,N_45055);
or U48223 (N_48223,N_45852,N_45448);
nand U48224 (N_48224,N_46234,N_46781);
or U48225 (N_48225,N_45373,N_45483);
nor U48226 (N_48226,N_47469,N_45235);
xnor U48227 (N_48227,N_46456,N_47242);
xor U48228 (N_48228,N_45192,N_46907);
nor U48229 (N_48229,N_45062,N_46691);
xor U48230 (N_48230,N_46847,N_46605);
xor U48231 (N_48231,N_46642,N_46029);
nor U48232 (N_48232,N_46879,N_45102);
xnor U48233 (N_48233,N_45960,N_46434);
nor U48234 (N_48234,N_45701,N_45010);
and U48235 (N_48235,N_45195,N_45968);
and U48236 (N_48236,N_46596,N_46148);
xor U48237 (N_48237,N_46502,N_45813);
nand U48238 (N_48238,N_45331,N_45047);
xnor U48239 (N_48239,N_45888,N_46533);
nor U48240 (N_48240,N_45400,N_46662);
nand U48241 (N_48241,N_45181,N_45922);
or U48242 (N_48242,N_46449,N_47429);
nor U48243 (N_48243,N_45988,N_46577);
and U48244 (N_48244,N_46314,N_46675);
or U48245 (N_48245,N_47204,N_45167);
and U48246 (N_48246,N_45262,N_47160);
nand U48247 (N_48247,N_46579,N_45795);
nor U48248 (N_48248,N_45647,N_45161);
nor U48249 (N_48249,N_46667,N_46145);
nor U48250 (N_48250,N_46100,N_47388);
or U48251 (N_48251,N_46660,N_46499);
nor U48252 (N_48252,N_47269,N_46352);
xor U48253 (N_48253,N_45363,N_45380);
nor U48254 (N_48254,N_45152,N_46633);
nand U48255 (N_48255,N_46898,N_46146);
xnor U48256 (N_48256,N_46053,N_46264);
and U48257 (N_48257,N_47277,N_46570);
nand U48258 (N_48258,N_46362,N_47362);
nand U48259 (N_48259,N_45270,N_45833);
nand U48260 (N_48260,N_45508,N_46261);
xor U48261 (N_48261,N_46785,N_46647);
xnor U48262 (N_48262,N_47324,N_47005);
xnor U48263 (N_48263,N_46204,N_45533);
and U48264 (N_48264,N_45899,N_46397);
nor U48265 (N_48265,N_45976,N_46630);
nand U48266 (N_48266,N_46319,N_46017);
and U48267 (N_48267,N_46120,N_46444);
nor U48268 (N_48268,N_46272,N_47074);
xor U48269 (N_48269,N_45992,N_46461);
nor U48270 (N_48270,N_46939,N_46732);
nor U48271 (N_48271,N_47475,N_46278);
and U48272 (N_48272,N_46950,N_46798);
nand U48273 (N_48273,N_45333,N_45740);
or U48274 (N_48274,N_45892,N_46463);
nor U48275 (N_48275,N_46223,N_47198);
or U48276 (N_48276,N_46801,N_46645);
and U48277 (N_48277,N_45902,N_46678);
nor U48278 (N_48278,N_45771,N_46404);
and U48279 (N_48279,N_46760,N_46394);
or U48280 (N_48280,N_47241,N_45869);
or U48281 (N_48281,N_46242,N_45840);
nor U48282 (N_48282,N_46926,N_45587);
and U48283 (N_48283,N_46241,N_45314);
xor U48284 (N_48284,N_47127,N_45281);
and U48285 (N_48285,N_45660,N_47424);
xnor U48286 (N_48286,N_46155,N_46973);
or U48287 (N_48287,N_45108,N_46425);
nand U48288 (N_48288,N_46885,N_47057);
nor U48289 (N_48289,N_47064,N_46600);
nand U48290 (N_48290,N_45554,N_45360);
or U48291 (N_48291,N_45149,N_46776);
nand U48292 (N_48292,N_45659,N_45114);
nor U48293 (N_48293,N_45823,N_47404);
or U48294 (N_48294,N_47272,N_45529);
or U48295 (N_48295,N_47406,N_47350);
nand U48296 (N_48296,N_46604,N_45292);
and U48297 (N_48297,N_47293,N_45234);
and U48298 (N_48298,N_46860,N_46217);
xor U48299 (N_48299,N_46191,N_47396);
xnor U48300 (N_48300,N_47105,N_45282);
and U48301 (N_48301,N_45880,N_45854);
or U48302 (N_48302,N_45290,N_45340);
and U48303 (N_48303,N_45410,N_47329);
nand U48304 (N_48304,N_45085,N_46713);
and U48305 (N_48305,N_45027,N_47370);
and U48306 (N_48306,N_45356,N_46725);
nand U48307 (N_48307,N_45375,N_46052);
nand U48308 (N_48308,N_46311,N_47136);
nand U48309 (N_48309,N_46036,N_46877);
xnor U48310 (N_48310,N_45504,N_47491);
and U48311 (N_48311,N_45187,N_46482);
xor U48312 (N_48312,N_46167,N_45440);
nand U48313 (N_48313,N_47188,N_46285);
and U48314 (N_48314,N_46569,N_46347);
nor U48315 (N_48315,N_45056,N_45697);
and U48316 (N_48316,N_45540,N_46868);
nand U48317 (N_48317,N_45358,N_45227);
xor U48318 (N_48318,N_46677,N_45841);
and U48319 (N_48319,N_46315,N_47097);
nor U48320 (N_48320,N_46992,N_46153);
nand U48321 (N_48321,N_47073,N_46743);
xor U48322 (N_48322,N_46530,N_47128);
xor U48323 (N_48323,N_45618,N_47311);
xnor U48324 (N_48324,N_45672,N_45505);
nor U48325 (N_48325,N_46894,N_47296);
and U48326 (N_48326,N_46711,N_47011);
or U48327 (N_48327,N_45724,N_46172);
and U48328 (N_48328,N_47352,N_45598);
and U48329 (N_48329,N_46107,N_46910);
nor U48330 (N_48330,N_46406,N_45537);
xnor U48331 (N_48331,N_45165,N_47209);
xor U48332 (N_48332,N_45422,N_45696);
nor U48333 (N_48333,N_47125,N_47151);
xnor U48334 (N_48334,N_47357,N_47090);
or U48335 (N_48335,N_45031,N_46139);
nand U48336 (N_48336,N_45130,N_47471);
nand U48337 (N_48337,N_45220,N_46475);
nor U48338 (N_48338,N_46918,N_46578);
nand U48339 (N_48339,N_46472,N_47194);
nor U48340 (N_48340,N_46774,N_45814);
or U48341 (N_48341,N_45369,N_46152);
or U48342 (N_48342,N_45008,N_46649);
xnor U48343 (N_48343,N_46203,N_47287);
nand U48344 (N_48344,N_45804,N_46176);
nand U48345 (N_48345,N_47411,N_46157);
or U48346 (N_48346,N_45466,N_46258);
nand U48347 (N_48347,N_46988,N_46275);
or U48348 (N_48348,N_46505,N_45258);
or U48349 (N_48349,N_46218,N_47492);
xor U48350 (N_48350,N_45686,N_45026);
nand U48351 (N_48351,N_47284,N_46069);
or U48352 (N_48352,N_45832,N_46468);
xor U48353 (N_48353,N_46429,N_45377);
nand U48354 (N_48354,N_46309,N_47245);
nor U48355 (N_48355,N_46321,N_46205);
and U48356 (N_48356,N_46407,N_45861);
nor U48357 (N_48357,N_46737,N_45844);
or U48358 (N_48358,N_46655,N_45198);
nand U48359 (N_48359,N_46870,N_47157);
xor U48360 (N_48360,N_47488,N_45736);
xor U48361 (N_48361,N_47152,N_45182);
and U48362 (N_48362,N_45717,N_46130);
nand U48363 (N_48363,N_45163,N_46664);
xnor U48364 (N_48364,N_46296,N_46532);
nor U48365 (N_48365,N_46248,N_45920);
xnor U48366 (N_48366,N_47399,N_46077);
or U48367 (N_48367,N_47343,N_46211);
or U48368 (N_48368,N_45589,N_45312);
nand U48369 (N_48369,N_45542,N_47325);
nor U48370 (N_48370,N_46999,N_46534);
and U48371 (N_48371,N_46327,N_45937);
nand U48372 (N_48372,N_46247,N_47170);
xnor U48373 (N_48373,N_47080,N_46609);
nor U48374 (N_48374,N_46508,N_45349);
xnor U48375 (N_48375,N_46210,N_45671);
and U48376 (N_48376,N_46613,N_46236);
or U48377 (N_48377,N_47016,N_47174);
or U48378 (N_48378,N_46061,N_46027);
nand U48379 (N_48379,N_46320,N_45260);
or U48380 (N_48380,N_45733,N_46448);
nor U48381 (N_48381,N_46903,N_46225);
or U48382 (N_48382,N_46480,N_46547);
or U48383 (N_48383,N_45938,N_47263);
xnor U48384 (N_48384,N_47393,N_45328);
and U48385 (N_48385,N_45374,N_47444);
nand U48386 (N_48386,N_46423,N_46941);
or U48387 (N_48387,N_46572,N_45915);
nor U48388 (N_48388,N_46516,N_47304);
and U48389 (N_48389,N_46976,N_45204);
or U48390 (N_48390,N_47091,N_45190);
and U48391 (N_48391,N_45077,N_46453);
nor U48392 (N_48392,N_47464,N_46431);
or U48393 (N_48393,N_45153,N_47018);
xnor U48394 (N_48394,N_47107,N_45604);
nand U48395 (N_48395,N_45903,N_46123);
or U48396 (N_48396,N_46420,N_46338);
nor U48397 (N_48397,N_47116,N_46757);
or U48398 (N_48398,N_45247,N_46173);
and U48399 (N_48399,N_46945,N_46994);
or U48400 (N_48400,N_46037,N_47186);
nor U48401 (N_48401,N_45819,N_46597);
and U48402 (N_48402,N_46260,N_46751);
nand U48403 (N_48403,N_47070,N_46323);
and U48404 (N_48404,N_45525,N_45749);
or U48405 (N_48405,N_46861,N_46925);
nand U48406 (N_48406,N_45521,N_45287);
and U48407 (N_48407,N_46358,N_45216);
and U48408 (N_48408,N_46455,N_47071);
or U48409 (N_48409,N_47478,N_47013);
nor U48410 (N_48410,N_45719,N_46055);
and U48411 (N_48411,N_46216,N_47458);
nor U48412 (N_48412,N_46806,N_47078);
and U48413 (N_48413,N_45241,N_45663);
or U48414 (N_48414,N_46566,N_46712);
and U48415 (N_48415,N_47482,N_45796);
xor U48416 (N_48416,N_46784,N_45383);
and U48417 (N_48417,N_46180,N_46119);
nand U48418 (N_48418,N_47421,N_47111);
nor U48419 (N_48419,N_45670,N_46561);
nand U48420 (N_48420,N_45728,N_46229);
nor U48421 (N_48421,N_45792,N_47278);
nor U48422 (N_48422,N_47101,N_45971);
nor U48423 (N_48423,N_45263,N_47108);
nor U48424 (N_48424,N_46390,N_45271);
or U48425 (N_48425,N_45761,N_46882);
xor U48426 (N_48426,N_47432,N_46946);
nand U48427 (N_48427,N_47365,N_47347);
and U48428 (N_48428,N_45577,N_46679);
or U48429 (N_48429,N_46291,N_45229);
xnor U48430 (N_48430,N_45567,N_47210);
and U48431 (N_48431,N_46175,N_46563);
nor U48432 (N_48432,N_45156,N_46972);
nor U48433 (N_48433,N_45978,N_46833);
nor U48434 (N_48434,N_45354,N_45520);
nor U48435 (N_48435,N_45386,N_45399);
and U48436 (N_48436,N_45097,N_46043);
or U48437 (N_48437,N_45335,N_46008);
xnor U48438 (N_48438,N_46065,N_47434);
or U48439 (N_48439,N_45825,N_47187);
nor U48440 (N_48440,N_45706,N_45874);
nand U48441 (N_48441,N_45449,N_46070);
nand U48442 (N_48442,N_45822,N_45036);
or U48443 (N_48443,N_45753,N_47459);
or U48444 (N_48444,N_46935,N_47302);
xnor U48445 (N_48445,N_47428,N_46631);
xor U48446 (N_48446,N_47498,N_47219);
xor U48447 (N_48447,N_46998,N_45913);
xor U48448 (N_48448,N_46854,N_46214);
and U48449 (N_48449,N_45597,N_47305);
xor U48450 (N_48450,N_47059,N_47159);
xor U48451 (N_48451,N_45959,N_46227);
and U48452 (N_48452,N_46387,N_45581);
nand U48453 (N_48453,N_45246,N_47467);
or U48454 (N_48454,N_45032,N_46346);
xnor U48455 (N_48455,N_46818,N_46072);
nor U48456 (N_48456,N_45249,N_47351);
xor U48457 (N_48457,N_45014,N_47361);
and U48458 (N_48458,N_46293,N_46964);
nor U48459 (N_48459,N_45489,N_45193);
and U48460 (N_48460,N_46129,N_47033);
or U48461 (N_48461,N_46408,N_46044);
nand U48462 (N_48462,N_47165,N_45867);
nor U48463 (N_48463,N_45850,N_47237);
and U48464 (N_48464,N_45624,N_45522);
or U48465 (N_48465,N_47076,N_45212);
nor U48466 (N_48466,N_45800,N_45343);
xor U48467 (N_48467,N_46588,N_45974);
nor U48468 (N_48468,N_46369,N_45666);
nor U48469 (N_48469,N_46367,N_45526);
and U48470 (N_48470,N_47162,N_46392);
xnor U48471 (N_48471,N_45500,N_46181);
or U48472 (N_48472,N_45019,N_47192);
nand U48473 (N_48473,N_45353,N_45392);
nor U48474 (N_48474,N_47171,N_46796);
nor U48475 (N_48475,N_45576,N_46959);
nand U48476 (N_48476,N_47298,N_45681);
and U48477 (N_48477,N_45675,N_45248);
or U48478 (N_48478,N_46492,N_46520);
nand U48479 (N_48479,N_46644,N_46253);
or U48480 (N_48480,N_45023,N_46715);
or U48481 (N_48481,N_46438,N_45674);
nor U48482 (N_48482,N_45236,N_46201);
and U48483 (N_48483,N_45677,N_45572);
nand U48484 (N_48484,N_45050,N_46891);
nand U48485 (N_48485,N_45214,N_47427);
and U48486 (N_48486,N_45297,N_47398);
nand U48487 (N_48487,N_45413,N_46025);
xnor U48488 (N_48488,N_46365,N_47392);
nor U48489 (N_48489,N_45145,N_47359);
nor U48490 (N_48490,N_46840,N_45517);
and U48491 (N_48491,N_46353,N_46799);
and U48492 (N_48492,N_45746,N_47372);
nor U48493 (N_48493,N_47222,N_47376);
nand U48494 (N_48494,N_46767,N_45326);
or U48495 (N_48495,N_46931,N_46133);
and U48496 (N_48496,N_46911,N_45615);
xnor U48497 (N_48497,N_46322,N_47335);
nor U48498 (N_48498,N_46256,N_45693);
xor U48499 (N_48499,N_46363,N_46194);
or U48500 (N_48500,N_47292,N_45412);
nor U48501 (N_48501,N_47217,N_45616);
nand U48502 (N_48502,N_47121,N_45443);
nand U48503 (N_48503,N_45653,N_47143);
nand U48504 (N_48504,N_46779,N_46699);
xor U48505 (N_48505,N_45141,N_47030);
or U48506 (N_48506,N_46692,N_46000);
and U48507 (N_48507,N_46124,N_47113);
nor U48508 (N_48508,N_45843,N_45538);
xor U48509 (N_48509,N_46924,N_47457);
nor U48510 (N_48510,N_47315,N_47295);
nand U48511 (N_48511,N_45817,N_47486);
nor U48512 (N_48512,N_46759,N_46503);
or U48513 (N_48513,N_46112,N_46238);
xnor U48514 (N_48514,N_46062,N_47134);
nand U48515 (N_48515,N_45514,N_46231);
or U48516 (N_48516,N_47384,N_46899);
or U48517 (N_48517,N_46378,N_46064);
xor U48518 (N_48518,N_46602,N_46364);
nor U48519 (N_48519,N_45583,N_46848);
or U48520 (N_48520,N_46676,N_46617);
and U48521 (N_48521,N_45551,N_46880);
nor U48522 (N_48522,N_46237,N_47461);
nor U48523 (N_48523,N_46615,N_45847);
and U48524 (N_48524,N_46243,N_45105);
and U48525 (N_48525,N_47485,N_45940);
xor U48526 (N_48526,N_45687,N_45051);
and U48527 (N_48527,N_46639,N_45035);
xnor U48528 (N_48528,N_47366,N_45475);
or U48529 (N_48529,N_46786,N_45484);
nor U48530 (N_48530,N_47397,N_47110);
xnor U48531 (N_48531,N_46554,N_45890);
xor U48532 (N_48532,N_46301,N_45030);
and U48533 (N_48533,N_46511,N_46957);
or U48534 (N_48534,N_45868,N_45278);
nor U48535 (N_48535,N_46344,N_46432);
xor U48536 (N_48536,N_46791,N_45751);
nand U48537 (N_48537,N_46388,N_45856);
xor U48538 (N_48538,N_47414,N_47042);
and U48539 (N_48539,N_45807,N_46280);
nor U48540 (N_48540,N_45876,N_45129);
nand U48541 (N_48541,N_47026,N_46458);
and U48542 (N_48542,N_47156,N_46334);
nor U48543 (N_48543,N_46197,N_45926);
and U48544 (N_48544,N_46749,N_47235);
nor U48545 (N_48545,N_46727,N_45142);
xor U48546 (N_48546,N_47002,N_45633);
xnor U48547 (N_48547,N_45853,N_46023);
nor U48548 (N_48548,N_46366,N_45455);
or U48549 (N_48549,N_47425,N_46905);
or U48550 (N_48550,N_46174,N_47184);
and U48551 (N_48551,N_45613,N_47055);
xnor U48552 (N_48552,N_46768,N_47494);
nor U48553 (N_48553,N_46295,N_46934);
nor U48554 (N_48554,N_45871,N_47246);
or U48555 (N_48555,N_47283,N_46851);
xor U48556 (N_48556,N_45645,N_46543);
and U48557 (N_48557,N_46020,N_45818);
and U48558 (N_48558,N_45347,N_45654);
xnor U48559 (N_48559,N_47169,N_46763);
and U48560 (N_48560,N_45464,N_46722);
xnor U48561 (N_48561,N_45337,N_46557);
xor U48562 (N_48562,N_46033,N_45658);
xor U48563 (N_48563,N_46003,N_45420);
nand U48564 (N_48564,N_46063,N_46682);
xor U48565 (N_48565,N_47185,N_46105);
nor U48566 (N_48566,N_46372,N_45601);
and U48567 (N_48567,N_46259,N_47058);
or U48568 (N_48568,N_45698,N_47462);
nand U48569 (N_48569,N_47200,N_45089);
or U48570 (N_48570,N_46634,N_46974);
nand U48571 (N_48571,N_47139,N_45933);
nor U48572 (N_48572,N_46386,N_46834);
nor U48573 (N_48573,N_47454,N_46747);
nor U48574 (N_48574,N_45307,N_46919);
nand U48575 (N_48575,N_46528,N_47040);
nor U48576 (N_48576,N_46193,N_45490);
and U48577 (N_48577,N_45131,N_47117);
nor U48578 (N_48578,N_46376,N_46102);
nand U48579 (N_48579,N_47275,N_46207);
nor U48580 (N_48580,N_47394,N_47062);
nor U48581 (N_48581,N_47423,N_46249);
nor U48582 (N_48582,N_46504,N_45485);
nor U48583 (N_48583,N_45406,N_45081);
and U48584 (N_48584,N_45269,N_46635);
xor U48585 (N_48585,N_45339,N_45610);
xnor U48586 (N_48586,N_46117,N_45463);
and U48587 (N_48587,N_46873,N_47166);
and U48588 (N_48588,N_45991,N_46164);
or U48589 (N_48589,N_46110,N_45176);
nor U48590 (N_48590,N_45928,N_46828);
nand U48591 (N_48591,N_47447,N_46018);
nor U48592 (N_48592,N_46628,N_45151);
or U48593 (N_48593,N_46092,N_45388);
nor U48594 (N_48594,N_45189,N_46015);
nor U48595 (N_48595,N_46239,N_45344);
nand U48596 (N_48596,N_45078,N_45953);
xor U48597 (N_48597,N_45918,N_47056);
and U48598 (N_48598,N_45146,N_45148);
nand U48599 (N_48599,N_46222,N_45491);
xnor U48600 (N_48600,N_47093,N_45251);
and U48601 (N_48601,N_46643,N_47230);
nand U48602 (N_48602,N_46082,N_46968);
or U48603 (N_48603,N_46134,N_45088);
xnor U48604 (N_48604,N_45909,N_45159);
xor U48605 (N_48605,N_45147,N_47360);
nor U48606 (N_48606,N_45812,N_46733);
xor U48607 (N_48607,N_46089,N_46906);
or U48608 (N_48608,N_46084,N_46189);
nand U48609 (N_48609,N_45883,N_45093);
nor U48610 (N_48610,N_46170,N_45557);
xnor U48611 (N_48611,N_47442,N_46622);
or U48612 (N_48612,N_45881,N_46007);
and U48613 (N_48613,N_47118,N_47009);
or U48614 (N_48614,N_45230,N_47175);
xnor U48615 (N_48615,N_45738,N_45103);
and U48616 (N_48616,N_45232,N_45299);
xor U48617 (N_48617,N_45154,N_45541);
or U48618 (N_48618,N_46928,N_46060);
and U48619 (N_48619,N_46559,N_46573);
xor U48620 (N_48620,N_45364,N_46329);
or U48621 (N_48621,N_45315,N_47103);
or U48622 (N_48622,N_45128,N_47264);
and U48623 (N_48623,N_45887,N_45622);
and U48624 (N_48624,N_46803,N_45425);
nand U48625 (N_48625,N_47211,N_46680);
xnor U48626 (N_48626,N_45685,N_45418);
nand U48627 (N_48627,N_45905,N_46594);
nor U48628 (N_48628,N_45980,N_45172);
nand U48629 (N_48629,N_47285,N_46902);
xor U48630 (N_48630,N_45334,N_45303);
and U48631 (N_48631,N_46917,N_46582);
xnor U48632 (N_48632,N_45196,N_45506);
xor U48633 (N_48633,N_45534,N_46304);
nor U48634 (N_48634,N_45090,N_45611);
nand U48635 (N_48635,N_45456,N_47123);
or U48636 (N_48636,N_45099,N_46476);
nor U48637 (N_48637,N_47473,N_45793);
nand U48638 (N_48638,N_46696,N_46980);
or U48639 (N_48639,N_45276,N_46698);
xor U48640 (N_48640,N_45810,N_46412);
nand U48641 (N_48641,N_46913,N_46661);
xnor U48642 (N_48642,N_46187,N_45327);
nor U48643 (N_48643,N_46822,N_47202);
and U48644 (N_48644,N_45921,N_45170);
xor U48645 (N_48645,N_45949,N_45059);
or U48646 (N_48646,N_45916,N_47257);
and U48647 (N_48647,N_46728,N_46808);
nor U48648 (N_48648,N_45769,N_46433);
or U48649 (N_48649,N_46839,N_45839);
xor U48650 (N_48650,N_45038,N_46838);
nor U48651 (N_48651,N_46094,N_46114);
nand U48652 (N_48652,N_45054,N_46297);
nor U48653 (N_48653,N_47449,N_46739);
or U48654 (N_48654,N_46648,N_45233);
and U48655 (N_48655,N_46815,N_47022);
and U48656 (N_48656,N_46740,N_47299);
and U48657 (N_48657,N_45708,N_45453);
nand U48658 (N_48658,N_47106,N_46702);
or U48659 (N_48659,N_46792,N_45188);
xor U48660 (N_48660,N_45259,N_45179);
nand U48661 (N_48661,N_46744,N_47331);
xor U48662 (N_48662,N_47102,N_46981);
xor U48663 (N_48663,N_46144,N_45264);
and U48664 (N_48664,N_46040,N_45257);
and U48665 (N_48665,N_46797,N_46753);
nand U48666 (N_48666,N_46116,N_45015);
xor U48667 (N_48667,N_46098,N_45688);
nand U48668 (N_48668,N_47044,N_47150);
xor U48669 (N_48669,N_46575,N_46487);
or U48670 (N_48670,N_47119,N_47147);
xnor U48671 (N_48671,N_45210,N_46932);
xor U48672 (N_48672,N_46689,N_46506);
and U48673 (N_48673,N_45046,N_45389);
or U48674 (N_48674,N_47379,N_47321);
and U48675 (N_48675,N_47029,N_45253);
or U48676 (N_48676,N_46131,N_45732);
xor U48677 (N_48677,N_46325,N_45963);
nand U48678 (N_48678,N_47265,N_45473);
xor U48679 (N_48679,N_47012,N_47273);
and U48680 (N_48680,N_45806,N_46659);
nor U48681 (N_48681,N_45252,N_46842);
nor U48682 (N_48682,N_46610,N_47010);
and U48683 (N_48683,N_45079,N_46621);
nand U48684 (N_48684,N_45003,N_46693);
nor U48685 (N_48685,N_46866,N_46809);
or U48686 (N_48686,N_46445,N_47124);
xor U48687 (N_48687,N_46342,N_45680);
nand U48688 (N_48688,N_46186,N_45518);
or U48689 (N_48689,N_45495,N_47371);
or U48690 (N_48690,N_46097,N_46730);
xor U48691 (N_48691,N_46829,N_47300);
nor U48692 (N_48692,N_47141,N_47254);
and U48693 (N_48693,N_46871,N_47356);
and U48694 (N_48694,N_45180,N_45445);
nand U48695 (N_48695,N_46307,N_47006);
xor U48696 (N_48696,N_45944,N_46493);
xor U48697 (N_48697,N_45742,N_45984);
and U48698 (N_48698,N_46132,N_45002);
or U48699 (N_48699,N_46584,N_45341);
and U48700 (N_48700,N_45906,N_47164);
xor U48701 (N_48701,N_46523,N_46142);
and U48702 (N_48702,N_47197,N_46393);
or U48703 (N_48703,N_47436,N_45826);
nor U48704 (N_48704,N_45989,N_46658);
nand U48705 (N_48705,N_47328,N_46929);
and U48706 (N_48706,N_46465,N_46978);
nor U48707 (N_48707,N_47483,N_46254);
nor U48708 (N_48708,N_47286,N_45942);
xor U48709 (N_48709,N_46850,N_45635);
and U48710 (N_48710,N_46916,N_45122);
or U48711 (N_48711,N_47131,N_46437);
xor U48712 (N_48712,N_45623,N_45566);
nand U48713 (N_48713,N_45479,N_46955);
nand U48714 (N_48714,N_46618,N_46632);
or U48715 (N_48715,N_46742,N_46336);
xor U48716 (N_48716,N_45831,N_45285);
xor U48717 (N_48717,N_45177,N_47463);
and U48718 (N_48718,N_46356,N_45427);
nand U48719 (N_48719,N_46317,N_45882);
nand U48720 (N_48720,N_45000,N_47251);
nor U48721 (N_48721,N_45778,N_45770);
nor U48722 (N_48722,N_46118,N_47256);
nand U48723 (N_48723,N_46426,N_47046);
and U48724 (N_48724,N_46937,N_46962);
nor U48725 (N_48725,N_46081,N_45901);
nor U48726 (N_48726,N_45238,N_45641);
xnor U48727 (N_48727,N_46567,N_45558);
nor U48728 (N_48728,N_47084,N_46824);
nor U48729 (N_48729,N_45429,N_46889);
or U48730 (N_48730,N_47060,N_45086);
nor U48731 (N_48731,N_45124,N_45174);
nor U48732 (N_48732,N_47229,N_47203);
xnor U48733 (N_48733,N_47430,N_46169);
and U48734 (N_48734,N_45345,N_47023);
and U48735 (N_48735,N_46096,N_47433);
nand U48736 (N_48736,N_47020,N_46921);
nor U48737 (N_48737,N_45402,N_46011);
and U48738 (N_48738,N_47015,N_46159);
xor U48739 (N_48739,N_46460,N_46111);
or U48740 (N_48740,N_45043,N_45612);
nand U48741 (N_48741,N_46762,N_46654);
or U48742 (N_48742,N_45985,N_47004);
and U48743 (N_48743,N_45584,N_47334);
nand U48744 (N_48744,N_45579,N_46059);
and U48745 (N_48745,N_45100,N_45735);
nor U48746 (N_48746,N_45411,N_46041);
xnor U48747 (N_48747,N_46416,N_46049);
and U48748 (N_48748,N_45668,N_45721);
nand U48749 (N_48749,N_46595,N_45158);
or U48750 (N_48750,N_46731,N_45316);
nor U48751 (N_48751,N_47432,N_46754);
nand U48752 (N_48752,N_46789,N_45994);
nor U48753 (N_48753,N_46118,N_45367);
xnor U48754 (N_48754,N_45959,N_46660);
and U48755 (N_48755,N_46561,N_46588);
nand U48756 (N_48756,N_45631,N_47169);
xor U48757 (N_48757,N_47451,N_45351);
and U48758 (N_48758,N_46823,N_47349);
nor U48759 (N_48759,N_46943,N_46099);
xor U48760 (N_48760,N_46457,N_45777);
xor U48761 (N_48761,N_46347,N_46736);
xnor U48762 (N_48762,N_47187,N_45206);
nor U48763 (N_48763,N_45029,N_46367);
nand U48764 (N_48764,N_45272,N_46059);
and U48765 (N_48765,N_47142,N_45043);
nand U48766 (N_48766,N_46172,N_45136);
and U48767 (N_48767,N_45906,N_45887);
or U48768 (N_48768,N_45706,N_45363);
nor U48769 (N_48769,N_45467,N_45942);
xnor U48770 (N_48770,N_46577,N_46158);
nor U48771 (N_48771,N_46545,N_47388);
nor U48772 (N_48772,N_45169,N_45572);
nor U48773 (N_48773,N_46741,N_45269);
nand U48774 (N_48774,N_46911,N_47259);
xor U48775 (N_48775,N_46091,N_46908);
nor U48776 (N_48776,N_45797,N_46814);
or U48777 (N_48777,N_46887,N_47005);
nand U48778 (N_48778,N_45834,N_47070);
nor U48779 (N_48779,N_46864,N_46473);
nand U48780 (N_48780,N_47095,N_45708);
xnor U48781 (N_48781,N_46468,N_46136);
xor U48782 (N_48782,N_45489,N_46903);
nor U48783 (N_48783,N_46504,N_45285);
xnor U48784 (N_48784,N_45141,N_47399);
nand U48785 (N_48785,N_47397,N_45916);
nand U48786 (N_48786,N_46632,N_45403);
nor U48787 (N_48787,N_46516,N_47368);
or U48788 (N_48788,N_45189,N_45251);
xnor U48789 (N_48789,N_46052,N_45084);
and U48790 (N_48790,N_46515,N_46445);
nand U48791 (N_48791,N_46280,N_46264);
nor U48792 (N_48792,N_45471,N_46884);
and U48793 (N_48793,N_46571,N_46384);
nand U48794 (N_48794,N_46194,N_45117);
xnor U48795 (N_48795,N_46079,N_46345);
or U48796 (N_48796,N_45304,N_46997);
or U48797 (N_48797,N_45820,N_45132);
nand U48798 (N_48798,N_46857,N_47234);
nand U48799 (N_48799,N_47085,N_45376);
or U48800 (N_48800,N_47432,N_46195);
or U48801 (N_48801,N_46578,N_45172);
and U48802 (N_48802,N_46693,N_46302);
xor U48803 (N_48803,N_45397,N_45792);
xor U48804 (N_48804,N_46158,N_45028);
and U48805 (N_48805,N_46577,N_45186);
or U48806 (N_48806,N_46313,N_45337);
or U48807 (N_48807,N_45302,N_45602);
and U48808 (N_48808,N_45420,N_46582);
xnor U48809 (N_48809,N_46119,N_45484);
xor U48810 (N_48810,N_46574,N_45797);
nand U48811 (N_48811,N_46134,N_46494);
and U48812 (N_48812,N_47030,N_47466);
or U48813 (N_48813,N_46443,N_47323);
and U48814 (N_48814,N_46309,N_47384);
xor U48815 (N_48815,N_46335,N_46525);
nand U48816 (N_48816,N_47135,N_46786);
nand U48817 (N_48817,N_46602,N_46892);
or U48818 (N_48818,N_45151,N_46809);
nor U48819 (N_48819,N_45624,N_45236);
or U48820 (N_48820,N_46366,N_46891);
or U48821 (N_48821,N_46347,N_46948);
nor U48822 (N_48822,N_45659,N_45716);
nand U48823 (N_48823,N_47155,N_45417);
or U48824 (N_48824,N_45320,N_46576);
nor U48825 (N_48825,N_46627,N_45054);
xor U48826 (N_48826,N_46180,N_45407);
nor U48827 (N_48827,N_46547,N_46751);
nand U48828 (N_48828,N_46067,N_45490);
and U48829 (N_48829,N_45713,N_45069);
and U48830 (N_48830,N_46781,N_47410);
and U48831 (N_48831,N_47051,N_45776);
nor U48832 (N_48832,N_46963,N_47138);
nor U48833 (N_48833,N_46666,N_47000);
or U48834 (N_48834,N_46390,N_45825);
nand U48835 (N_48835,N_45878,N_46227);
and U48836 (N_48836,N_47036,N_46697);
xnor U48837 (N_48837,N_46694,N_47108);
nor U48838 (N_48838,N_45748,N_47188);
and U48839 (N_48839,N_46241,N_45149);
xnor U48840 (N_48840,N_46042,N_46741);
nor U48841 (N_48841,N_46549,N_47117);
nor U48842 (N_48842,N_45437,N_47020);
or U48843 (N_48843,N_46077,N_46657);
and U48844 (N_48844,N_47024,N_46819);
or U48845 (N_48845,N_47410,N_47194);
nor U48846 (N_48846,N_45838,N_45304);
and U48847 (N_48847,N_47435,N_47259);
and U48848 (N_48848,N_47217,N_46515);
nor U48849 (N_48849,N_45833,N_45047);
nand U48850 (N_48850,N_45788,N_45668);
and U48851 (N_48851,N_46086,N_45148);
and U48852 (N_48852,N_45869,N_46373);
or U48853 (N_48853,N_46047,N_45238);
nor U48854 (N_48854,N_45491,N_45208);
and U48855 (N_48855,N_45419,N_45731);
or U48856 (N_48856,N_46242,N_46491);
or U48857 (N_48857,N_47393,N_45281);
or U48858 (N_48858,N_45976,N_46858);
or U48859 (N_48859,N_46290,N_45946);
nand U48860 (N_48860,N_47255,N_45522);
nand U48861 (N_48861,N_47448,N_46396);
or U48862 (N_48862,N_45606,N_45896);
nand U48863 (N_48863,N_46106,N_46423);
nor U48864 (N_48864,N_46532,N_47055);
and U48865 (N_48865,N_46287,N_45479);
or U48866 (N_48866,N_45695,N_47089);
and U48867 (N_48867,N_46675,N_46695);
nor U48868 (N_48868,N_46271,N_46077);
nand U48869 (N_48869,N_47351,N_46621);
and U48870 (N_48870,N_45517,N_47216);
nor U48871 (N_48871,N_46506,N_46538);
xor U48872 (N_48872,N_47265,N_45355);
nor U48873 (N_48873,N_46770,N_46359);
xor U48874 (N_48874,N_46445,N_46149);
or U48875 (N_48875,N_45404,N_45851);
nor U48876 (N_48876,N_46167,N_47190);
xnor U48877 (N_48877,N_46370,N_46904);
xor U48878 (N_48878,N_47033,N_46013);
and U48879 (N_48879,N_46952,N_45106);
xnor U48880 (N_48880,N_45511,N_46125);
nand U48881 (N_48881,N_45025,N_45488);
xor U48882 (N_48882,N_45685,N_45573);
nor U48883 (N_48883,N_47214,N_45575);
nand U48884 (N_48884,N_46086,N_46789);
nor U48885 (N_48885,N_46847,N_46777);
nand U48886 (N_48886,N_45073,N_46272);
nor U48887 (N_48887,N_46265,N_47411);
nor U48888 (N_48888,N_46470,N_46411);
or U48889 (N_48889,N_45679,N_45196);
xor U48890 (N_48890,N_45985,N_45937);
nor U48891 (N_48891,N_45635,N_46611);
nand U48892 (N_48892,N_45784,N_46737);
and U48893 (N_48893,N_45289,N_46717);
nor U48894 (N_48894,N_45154,N_46115);
and U48895 (N_48895,N_45030,N_46437);
xor U48896 (N_48896,N_46317,N_46041);
xnor U48897 (N_48897,N_47442,N_46395);
xor U48898 (N_48898,N_46841,N_45412);
nand U48899 (N_48899,N_45552,N_46284);
and U48900 (N_48900,N_45050,N_46858);
nor U48901 (N_48901,N_46435,N_46565);
nand U48902 (N_48902,N_46900,N_46703);
nor U48903 (N_48903,N_47438,N_47237);
xor U48904 (N_48904,N_46778,N_45238);
and U48905 (N_48905,N_46828,N_46096);
nand U48906 (N_48906,N_45362,N_46570);
nor U48907 (N_48907,N_47079,N_45598);
or U48908 (N_48908,N_45686,N_46176);
and U48909 (N_48909,N_47435,N_46352);
nor U48910 (N_48910,N_46234,N_45929);
xor U48911 (N_48911,N_47129,N_45198);
nor U48912 (N_48912,N_46175,N_46968);
and U48913 (N_48913,N_46033,N_46332);
nor U48914 (N_48914,N_46782,N_46871);
and U48915 (N_48915,N_46005,N_47299);
or U48916 (N_48916,N_45622,N_45545);
and U48917 (N_48917,N_45899,N_46738);
or U48918 (N_48918,N_46849,N_46842);
or U48919 (N_48919,N_45569,N_46950);
or U48920 (N_48920,N_45998,N_46109);
nor U48921 (N_48921,N_45889,N_47152);
or U48922 (N_48922,N_46194,N_45049);
nor U48923 (N_48923,N_45652,N_45655);
and U48924 (N_48924,N_46130,N_45715);
or U48925 (N_48925,N_46859,N_46449);
nor U48926 (N_48926,N_46241,N_47247);
nor U48927 (N_48927,N_46330,N_45945);
nand U48928 (N_48928,N_46800,N_46638);
and U48929 (N_48929,N_46804,N_45470);
nand U48930 (N_48930,N_46296,N_45258);
nand U48931 (N_48931,N_46633,N_46429);
or U48932 (N_48932,N_46966,N_46232);
nand U48933 (N_48933,N_45673,N_45607);
nor U48934 (N_48934,N_45653,N_47081);
nor U48935 (N_48935,N_46276,N_46579);
nor U48936 (N_48936,N_46186,N_45898);
nor U48937 (N_48937,N_46341,N_46735);
nand U48938 (N_48938,N_46757,N_46772);
xnor U48939 (N_48939,N_46815,N_46030);
nor U48940 (N_48940,N_46695,N_45612);
nand U48941 (N_48941,N_46377,N_45663);
nor U48942 (N_48942,N_45452,N_46926);
and U48943 (N_48943,N_46676,N_46105);
xor U48944 (N_48944,N_45867,N_45564);
or U48945 (N_48945,N_46531,N_47218);
nor U48946 (N_48946,N_45458,N_47131);
nand U48947 (N_48947,N_46153,N_47049);
nor U48948 (N_48948,N_45069,N_46290);
xor U48949 (N_48949,N_47039,N_47074);
and U48950 (N_48950,N_46144,N_46914);
or U48951 (N_48951,N_45332,N_45563);
and U48952 (N_48952,N_47317,N_46268);
nor U48953 (N_48953,N_46669,N_46691);
xnor U48954 (N_48954,N_46041,N_45317);
nand U48955 (N_48955,N_47186,N_45940);
or U48956 (N_48956,N_46770,N_45346);
nand U48957 (N_48957,N_46249,N_46887);
xnor U48958 (N_48958,N_45902,N_45408);
nor U48959 (N_48959,N_45328,N_46911);
and U48960 (N_48960,N_45245,N_45821);
nor U48961 (N_48961,N_45558,N_46431);
nor U48962 (N_48962,N_45922,N_46138);
nor U48963 (N_48963,N_46431,N_45138);
or U48964 (N_48964,N_45537,N_45908);
and U48965 (N_48965,N_47267,N_46091);
and U48966 (N_48966,N_45664,N_46523);
and U48967 (N_48967,N_47376,N_47469);
xor U48968 (N_48968,N_45394,N_45230);
xor U48969 (N_48969,N_46042,N_45400);
nor U48970 (N_48970,N_46593,N_47134);
or U48971 (N_48971,N_45397,N_45515);
nor U48972 (N_48972,N_45103,N_46384);
nand U48973 (N_48973,N_45904,N_46129);
xnor U48974 (N_48974,N_46258,N_45498);
nor U48975 (N_48975,N_46586,N_45954);
xor U48976 (N_48976,N_45289,N_47006);
nor U48977 (N_48977,N_45191,N_45742);
nor U48978 (N_48978,N_45608,N_45199);
nor U48979 (N_48979,N_45011,N_46999);
nand U48980 (N_48980,N_46698,N_47493);
nand U48981 (N_48981,N_46218,N_46718);
xor U48982 (N_48982,N_45769,N_46087);
nand U48983 (N_48983,N_46080,N_47402);
nor U48984 (N_48984,N_45254,N_45968);
or U48985 (N_48985,N_45377,N_45391);
or U48986 (N_48986,N_46563,N_47480);
xnor U48987 (N_48987,N_45292,N_45300);
or U48988 (N_48988,N_46814,N_45474);
xnor U48989 (N_48989,N_46242,N_46116);
nor U48990 (N_48990,N_45647,N_45385);
nor U48991 (N_48991,N_46511,N_45471);
and U48992 (N_48992,N_46087,N_45056);
nand U48993 (N_48993,N_47484,N_46710);
and U48994 (N_48994,N_45210,N_45373);
xnor U48995 (N_48995,N_46567,N_46926);
xnor U48996 (N_48996,N_46227,N_45931);
or U48997 (N_48997,N_46307,N_45522);
nor U48998 (N_48998,N_45053,N_47249);
xor U48999 (N_48999,N_46439,N_46691);
or U49000 (N_49000,N_47313,N_46486);
and U49001 (N_49001,N_47232,N_47409);
nor U49002 (N_49002,N_45052,N_46298);
nand U49003 (N_49003,N_46059,N_46395);
nor U49004 (N_49004,N_46200,N_45872);
xnor U49005 (N_49005,N_45720,N_46767);
nor U49006 (N_49006,N_45850,N_46226);
and U49007 (N_49007,N_47307,N_47106);
or U49008 (N_49008,N_47365,N_46324);
or U49009 (N_49009,N_45173,N_46381);
and U49010 (N_49010,N_46038,N_46210);
nor U49011 (N_49011,N_46695,N_45586);
nor U49012 (N_49012,N_46784,N_45869);
nor U49013 (N_49013,N_45263,N_46007);
xnor U49014 (N_49014,N_46844,N_45698);
or U49015 (N_49015,N_46431,N_46425);
nand U49016 (N_49016,N_45958,N_47273);
nor U49017 (N_49017,N_46358,N_45301);
nor U49018 (N_49018,N_46143,N_46179);
and U49019 (N_49019,N_46681,N_47110);
or U49020 (N_49020,N_46590,N_46629);
and U49021 (N_49021,N_45125,N_45635);
xor U49022 (N_49022,N_46880,N_45625);
and U49023 (N_49023,N_47079,N_46465);
nand U49024 (N_49024,N_46137,N_45067);
or U49025 (N_49025,N_46722,N_46199);
nor U49026 (N_49026,N_46618,N_47171);
xor U49027 (N_49027,N_46113,N_46282);
nor U49028 (N_49028,N_46407,N_45575);
nand U49029 (N_49029,N_46885,N_45384);
and U49030 (N_49030,N_47215,N_47224);
or U49031 (N_49031,N_45048,N_46825);
xor U49032 (N_49032,N_45192,N_45880);
nand U49033 (N_49033,N_45039,N_45089);
or U49034 (N_49034,N_46869,N_46625);
and U49035 (N_49035,N_47039,N_45235);
nor U49036 (N_49036,N_45208,N_45599);
xor U49037 (N_49037,N_45574,N_47486);
and U49038 (N_49038,N_45767,N_46936);
nand U49039 (N_49039,N_47272,N_45255);
xor U49040 (N_49040,N_46496,N_45608);
xnor U49041 (N_49041,N_47304,N_46405);
or U49042 (N_49042,N_46589,N_46095);
nand U49043 (N_49043,N_46231,N_47008);
nor U49044 (N_49044,N_47220,N_47438);
nand U49045 (N_49045,N_46658,N_47265);
xor U49046 (N_49046,N_46218,N_45807);
or U49047 (N_49047,N_46458,N_47273);
or U49048 (N_49048,N_47466,N_47160);
xor U49049 (N_49049,N_45632,N_46317);
nand U49050 (N_49050,N_45894,N_46143);
nand U49051 (N_49051,N_46718,N_47035);
nor U49052 (N_49052,N_47070,N_45446);
nand U49053 (N_49053,N_45658,N_47259);
xnor U49054 (N_49054,N_46773,N_46501);
nand U49055 (N_49055,N_46447,N_45801);
nand U49056 (N_49056,N_45618,N_46206);
nor U49057 (N_49057,N_45133,N_46385);
nand U49058 (N_49058,N_45531,N_46236);
xnor U49059 (N_49059,N_46917,N_46757);
and U49060 (N_49060,N_45753,N_45467);
or U49061 (N_49061,N_45335,N_46117);
and U49062 (N_49062,N_46338,N_45916);
nor U49063 (N_49063,N_46895,N_46168);
nand U49064 (N_49064,N_45461,N_45478);
and U49065 (N_49065,N_46070,N_46787);
or U49066 (N_49066,N_45336,N_45598);
and U49067 (N_49067,N_45443,N_45326);
nand U49068 (N_49068,N_47235,N_45058);
and U49069 (N_49069,N_47316,N_45688);
nor U49070 (N_49070,N_46143,N_47363);
nand U49071 (N_49071,N_47442,N_46484);
xnor U49072 (N_49072,N_45702,N_46650);
nand U49073 (N_49073,N_45890,N_45114);
or U49074 (N_49074,N_45033,N_47280);
and U49075 (N_49075,N_45763,N_46391);
nand U49076 (N_49076,N_46593,N_45726);
nor U49077 (N_49077,N_45361,N_45537);
nand U49078 (N_49078,N_46628,N_46991);
or U49079 (N_49079,N_45684,N_46798);
nand U49080 (N_49080,N_46238,N_46770);
nor U49081 (N_49081,N_45834,N_45359);
nand U49082 (N_49082,N_45332,N_46342);
or U49083 (N_49083,N_45349,N_46868);
or U49084 (N_49084,N_46765,N_45957);
or U49085 (N_49085,N_47133,N_45801);
nor U49086 (N_49086,N_46094,N_45592);
xor U49087 (N_49087,N_47402,N_45350);
nor U49088 (N_49088,N_45575,N_47272);
or U49089 (N_49089,N_47034,N_47318);
xor U49090 (N_49090,N_45226,N_46156);
and U49091 (N_49091,N_45630,N_47182);
nand U49092 (N_49092,N_45707,N_47174);
xor U49093 (N_49093,N_45379,N_45449);
xor U49094 (N_49094,N_47386,N_47015);
and U49095 (N_49095,N_47499,N_45606);
nor U49096 (N_49096,N_46785,N_47160);
and U49097 (N_49097,N_46060,N_45437);
or U49098 (N_49098,N_45792,N_47163);
and U49099 (N_49099,N_45339,N_47337);
xor U49100 (N_49100,N_46253,N_46705);
nand U49101 (N_49101,N_46179,N_45847);
and U49102 (N_49102,N_45409,N_45938);
and U49103 (N_49103,N_45374,N_46518);
or U49104 (N_49104,N_45687,N_47307);
or U49105 (N_49105,N_45719,N_47221);
and U49106 (N_49106,N_46931,N_46677);
nand U49107 (N_49107,N_46863,N_45884);
and U49108 (N_49108,N_47200,N_46702);
nor U49109 (N_49109,N_47004,N_47198);
or U49110 (N_49110,N_45519,N_45630);
xor U49111 (N_49111,N_46822,N_47253);
or U49112 (N_49112,N_45026,N_46042);
and U49113 (N_49113,N_47102,N_46377);
nor U49114 (N_49114,N_46229,N_46762);
and U49115 (N_49115,N_45649,N_45979);
nand U49116 (N_49116,N_45246,N_46632);
nor U49117 (N_49117,N_47279,N_45577);
nand U49118 (N_49118,N_46406,N_46164);
or U49119 (N_49119,N_46360,N_46017);
nand U49120 (N_49120,N_45769,N_47446);
xnor U49121 (N_49121,N_45276,N_46625);
and U49122 (N_49122,N_45568,N_45706);
or U49123 (N_49123,N_46428,N_47004);
or U49124 (N_49124,N_45392,N_46854);
and U49125 (N_49125,N_46786,N_45456);
and U49126 (N_49126,N_47290,N_46032);
or U49127 (N_49127,N_45633,N_45762);
and U49128 (N_49128,N_45089,N_45133);
nand U49129 (N_49129,N_46347,N_45598);
xnor U49130 (N_49130,N_47357,N_46157);
or U49131 (N_49131,N_46608,N_46076);
nor U49132 (N_49132,N_47009,N_45728);
or U49133 (N_49133,N_46276,N_46673);
nor U49134 (N_49134,N_47289,N_45406);
nand U49135 (N_49135,N_45348,N_46722);
nor U49136 (N_49136,N_46199,N_45586);
nand U49137 (N_49137,N_45835,N_47255);
or U49138 (N_49138,N_46335,N_47408);
and U49139 (N_49139,N_46867,N_46746);
nand U49140 (N_49140,N_46974,N_46862);
and U49141 (N_49141,N_46802,N_47115);
nor U49142 (N_49142,N_45040,N_47268);
nor U49143 (N_49143,N_47102,N_47281);
xnor U49144 (N_49144,N_46587,N_47248);
nor U49145 (N_49145,N_45562,N_46017);
nand U49146 (N_49146,N_46293,N_45287);
and U49147 (N_49147,N_45499,N_45626);
or U49148 (N_49148,N_46525,N_47384);
and U49149 (N_49149,N_45568,N_47154);
nand U49150 (N_49150,N_47390,N_47311);
xor U49151 (N_49151,N_47131,N_46654);
nand U49152 (N_49152,N_46925,N_45798);
nand U49153 (N_49153,N_46972,N_46131);
xnor U49154 (N_49154,N_46607,N_46622);
nand U49155 (N_49155,N_45789,N_46434);
nand U49156 (N_49156,N_45308,N_45178);
or U49157 (N_49157,N_45635,N_47097);
and U49158 (N_49158,N_45707,N_45679);
and U49159 (N_49159,N_47341,N_47206);
xor U49160 (N_49160,N_45892,N_46287);
or U49161 (N_49161,N_46864,N_46988);
and U49162 (N_49162,N_47456,N_46118);
or U49163 (N_49163,N_45123,N_46144);
and U49164 (N_49164,N_46627,N_47243);
nor U49165 (N_49165,N_47379,N_47006);
nand U49166 (N_49166,N_47073,N_45479);
or U49167 (N_49167,N_47421,N_47023);
or U49168 (N_49168,N_47156,N_45038);
and U49169 (N_49169,N_45410,N_45124);
and U49170 (N_49170,N_47211,N_46937);
xor U49171 (N_49171,N_46156,N_46681);
and U49172 (N_49172,N_47079,N_47394);
nand U49173 (N_49173,N_46153,N_45168);
nor U49174 (N_49174,N_46283,N_45891);
or U49175 (N_49175,N_47168,N_47020);
nor U49176 (N_49176,N_45622,N_45665);
nand U49177 (N_49177,N_46648,N_45071);
nor U49178 (N_49178,N_46085,N_45241);
or U49179 (N_49179,N_46437,N_46317);
and U49180 (N_49180,N_46709,N_47027);
and U49181 (N_49181,N_46139,N_46235);
or U49182 (N_49182,N_45526,N_46282);
or U49183 (N_49183,N_46726,N_45675);
nor U49184 (N_49184,N_45753,N_46802);
or U49185 (N_49185,N_45050,N_47023);
or U49186 (N_49186,N_46817,N_47084);
xnor U49187 (N_49187,N_47002,N_46847);
and U49188 (N_49188,N_46576,N_45845);
xor U49189 (N_49189,N_46177,N_45922);
xnor U49190 (N_49190,N_45031,N_45130);
nor U49191 (N_49191,N_47342,N_46218);
xor U49192 (N_49192,N_46680,N_45422);
nor U49193 (N_49193,N_47099,N_47055);
xor U49194 (N_49194,N_46148,N_47093);
nand U49195 (N_49195,N_45325,N_45723);
nor U49196 (N_49196,N_45866,N_46066);
and U49197 (N_49197,N_45393,N_45508);
and U49198 (N_49198,N_46854,N_47224);
nand U49199 (N_49199,N_46037,N_46491);
nand U49200 (N_49200,N_45716,N_47445);
or U49201 (N_49201,N_46513,N_47137);
xor U49202 (N_49202,N_45468,N_46837);
nand U49203 (N_49203,N_45099,N_46840);
and U49204 (N_49204,N_46035,N_45930);
nand U49205 (N_49205,N_46588,N_47351);
nor U49206 (N_49206,N_47398,N_46890);
xor U49207 (N_49207,N_47115,N_45984);
and U49208 (N_49208,N_46649,N_47242);
and U49209 (N_49209,N_46342,N_46360);
xor U49210 (N_49210,N_47262,N_45247);
and U49211 (N_49211,N_45865,N_46774);
or U49212 (N_49212,N_46303,N_46204);
or U49213 (N_49213,N_45313,N_45292);
nand U49214 (N_49214,N_46410,N_46952);
xor U49215 (N_49215,N_46577,N_46752);
and U49216 (N_49216,N_45106,N_46325);
and U49217 (N_49217,N_45170,N_46971);
xnor U49218 (N_49218,N_45403,N_45207);
xor U49219 (N_49219,N_45866,N_45954);
or U49220 (N_49220,N_47373,N_46484);
or U49221 (N_49221,N_45232,N_45991);
and U49222 (N_49222,N_46247,N_45155);
nand U49223 (N_49223,N_46235,N_45522);
nor U49224 (N_49224,N_46990,N_47492);
and U49225 (N_49225,N_45711,N_47158);
and U49226 (N_49226,N_46767,N_46453);
nor U49227 (N_49227,N_45927,N_45584);
or U49228 (N_49228,N_45900,N_46936);
nor U49229 (N_49229,N_47370,N_46746);
xor U49230 (N_49230,N_47221,N_47004);
xnor U49231 (N_49231,N_46992,N_47276);
and U49232 (N_49232,N_46550,N_45711);
nor U49233 (N_49233,N_45218,N_45664);
or U49234 (N_49234,N_46070,N_46334);
and U49235 (N_49235,N_47022,N_46921);
or U49236 (N_49236,N_46073,N_45349);
nor U49237 (N_49237,N_46547,N_46464);
or U49238 (N_49238,N_46072,N_45465);
nor U49239 (N_49239,N_46268,N_47325);
nand U49240 (N_49240,N_46388,N_47287);
nor U49241 (N_49241,N_45934,N_45421);
nand U49242 (N_49242,N_46159,N_45695);
nor U49243 (N_49243,N_46369,N_46826);
nand U49244 (N_49244,N_45130,N_47300);
or U49245 (N_49245,N_45772,N_46130);
and U49246 (N_49246,N_47340,N_45709);
xnor U49247 (N_49247,N_45187,N_45086);
xnor U49248 (N_49248,N_45900,N_45618);
nand U49249 (N_49249,N_45410,N_47437);
and U49250 (N_49250,N_45237,N_47103);
nor U49251 (N_49251,N_46884,N_45858);
or U49252 (N_49252,N_47274,N_46140);
xor U49253 (N_49253,N_45296,N_46261);
nor U49254 (N_49254,N_45424,N_45104);
xnor U49255 (N_49255,N_45504,N_47439);
nand U49256 (N_49256,N_45112,N_46146);
nor U49257 (N_49257,N_46707,N_46470);
and U49258 (N_49258,N_45424,N_47321);
nor U49259 (N_49259,N_46102,N_47421);
or U49260 (N_49260,N_47117,N_46495);
or U49261 (N_49261,N_47025,N_45859);
nor U49262 (N_49262,N_45842,N_46651);
or U49263 (N_49263,N_45509,N_46838);
nand U49264 (N_49264,N_46432,N_46254);
nor U49265 (N_49265,N_46127,N_45578);
or U49266 (N_49266,N_45054,N_46249);
xor U49267 (N_49267,N_46049,N_46007);
nor U49268 (N_49268,N_45665,N_47376);
xnor U49269 (N_49269,N_45794,N_46825);
and U49270 (N_49270,N_47154,N_45476);
xor U49271 (N_49271,N_46349,N_45803);
or U49272 (N_49272,N_45700,N_46772);
nand U49273 (N_49273,N_45218,N_46999);
or U49274 (N_49274,N_45586,N_46468);
or U49275 (N_49275,N_47173,N_45090);
xnor U49276 (N_49276,N_45980,N_45483);
xnor U49277 (N_49277,N_47481,N_45836);
and U49278 (N_49278,N_46123,N_45335);
and U49279 (N_49279,N_46693,N_45232);
and U49280 (N_49280,N_45562,N_46438);
xnor U49281 (N_49281,N_45844,N_47152);
nand U49282 (N_49282,N_45643,N_46717);
and U49283 (N_49283,N_45213,N_47360);
nand U49284 (N_49284,N_47178,N_45027);
nor U49285 (N_49285,N_45875,N_46091);
nor U49286 (N_49286,N_47275,N_45872);
nand U49287 (N_49287,N_47160,N_45976);
and U49288 (N_49288,N_45468,N_46974);
xnor U49289 (N_49289,N_45655,N_47121);
xor U49290 (N_49290,N_46429,N_46350);
or U49291 (N_49291,N_45227,N_47078);
nand U49292 (N_49292,N_45581,N_46274);
nand U49293 (N_49293,N_45795,N_46736);
and U49294 (N_49294,N_46283,N_47084);
nor U49295 (N_49295,N_45134,N_45038);
or U49296 (N_49296,N_46694,N_46056);
nand U49297 (N_49297,N_45866,N_45718);
and U49298 (N_49298,N_46383,N_46125);
nor U49299 (N_49299,N_45845,N_46568);
nor U49300 (N_49300,N_45180,N_46724);
xnor U49301 (N_49301,N_46833,N_45773);
nand U49302 (N_49302,N_46112,N_45326);
xor U49303 (N_49303,N_47097,N_45934);
nor U49304 (N_49304,N_45074,N_45872);
xnor U49305 (N_49305,N_47294,N_46617);
xnor U49306 (N_49306,N_47498,N_47098);
xnor U49307 (N_49307,N_45553,N_47281);
or U49308 (N_49308,N_45736,N_46630);
or U49309 (N_49309,N_45887,N_46061);
nand U49310 (N_49310,N_45766,N_45641);
and U49311 (N_49311,N_45525,N_46629);
and U49312 (N_49312,N_45419,N_47081);
or U49313 (N_49313,N_45754,N_46426);
or U49314 (N_49314,N_45450,N_45944);
xnor U49315 (N_49315,N_47181,N_45098);
nor U49316 (N_49316,N_46057,N_45432);
nor U49317 (N_49317,N_45392,N_46768);
xnor U49318 (N_49318,N_45449,N_45589);
nor U49319 (N_49319,N_46336,N_46193);
xnor U49320 (N_49320,N_46394,N_47102);
nand U49321 (N_49321,N_45411,N_47170);
or U49322 (N_49322,N_45632,N_46658);
nand U49323 (N_49323,N_45502,N_47112);
nor U49324 (N_49324,N_45141,N_47469);
nor U49325 (N_49325,N_45688,N_45178);
nand U49326 (N_49326,N_46365,N_47448);
nor U49327 (N_49327,N_45424,N_47136);
nand U49328 (N_49328,N_47489,N_45741);
or U49329 (N_49329,N_46450,N_46082);
xnor U49330 (N_49330,N_47444,N_47151);
and U49331 (N_49331,N_45870,N_47248);
xnor U49332 (N_49332,N_45702,N_47096);
xor U49333 (N_49333,N_46843,N_47186);
nand U49334 (N_49334,N_46845,N_46837);
or U49335 (N_49335,N_46398,N_47045);
nand U49336 (N_49336,N_45864,N_46666);
nand U49337 (N_49337,N_47005,N_46946);
xor U49338 (N_49338,N_45430,N_45032);
nor U49339 (N_49339,N_47132,N_45597);
nand U49340 (N_49340,N_47080,N_47153);
xor U49341 (N_49341,N_45541,N_46527);
nand U49342 (N_49342,N_45905,N_45314);
nand U49343 (N_49343,N_45397,N_47038);
xor U49344 (N_49344,N_45344,N_45396);
or U49345 (N_49345,N_46360,N_46402);
and U49346 (N_49346,N_46160,N_47170);
nor U49347 (N_49347,N_45921,N_46918);
nor U49348 (N_49348,N_46487,N_47052);
and U49349 (N_49349,N_46826,N_45939);
and U49350 (N_49350,N_45684,N_45473);
xnor U49351 (N_49351,N_45541,N_45247);
and U49352 (N_49352,N_45958,N_46245);
xnor U49353 (N_49353,N_45196,N_46088);
and U49354 (N_49354,N_45612,N_47044);
xnor U49355 (N_49355,N_47262,N_47415);
and U49356 (N_49356,N_47292,N_46797);
and U49357 (N_49357,N_45339,N_45790);
and U49358 (N_49358,N_45314,N_45613);
nand U49359 (N_49359,N_46167,N_45459);
nor U49360 (N_49360,N_45861,N_46257);
and U49361 (N_49361,N_45799,N_47092);
or U49362 (N_49362,N_45629,N_46085);
nand U49363 (N_49363,N_47262,N_46803);
and U49364 (N_49364,N_47035,N_46547);
nor U49365 (N_49365,N_47449,N_45264);
and U49366 (N_49366,N_46678,N_47357);
xnor U49367 (N_49367,N_45338,N_46978);
nor U49368 (N_49368,N_46679,N_45338);
or U49369 (N_49369,N_46270,N_47439);
nor U49370 (N_49370,N_45606,N_45995);
xor U49371 (N_49371,N_45687,N_46198);
or U49372 (N_49372,N_46358,N_45012);
or U49373 (N_49373,N_45053,N_45130);
and U49374 (N_49374,N_47464,N_46719);
or U49375 (N_49375,N_47213,N_47362);
nor U49376 (N_49376,N_47362,N_46139);
or U49377 (N_49377,N_45450,N_46616);
nor U49378 (N_49378,N_46094,N_45378);
and U49379 (N_49379,N_47067,N_47353);
and U49380 (N_49380,N_45880,N_45580);
xnor U49381 (N_49381,N_46781,N_46555);
nand U49382 (N_49382,N_46488,N_47066);
nand U49383 (N_49383,N_47356,N_45295);
xnor U49384 (N_49384,N_47053,N_46238);
nand U49385 (N_49385,N_46995,N_45610);
xnor U49386 (N_49386,N_45221,N_45695);
or U49387 (N_49387,N_46261,N_46264);
xor U49388 (N_49388,N_45012,N_45575);
and U49389 (N_49389,N_46378,N_45987);
or U49390 (N_49390,N_46815,N_46289);
xor U49391 (N_49391,N_47462,N_47092);
or U49392 (N_49392,N_46310,N_47107);
and U49393 (N_49393,N_46073,N_46750);
nand U49394 (N_49394,N_47388,N_45856);
xnor U49395 (N_49395,N_47040,N_46856);
and U49396 (N_49396,N_46816,N_45675);
or U49397 (N_49397,N_45913,N_45791);
nand U49398 (N_49398,N_45048,N_47333);
nand U49399 (N_49399,N_45557,N_45140);
or U49400 (N_49400,N_45427,N_46852);
nand U49401 (N_49401,N_45616,N_46997);
xor U49402 (N_49402,N_45144,N_45023);
and U49403 (N_49403,N_45791,N_45671);
xnor U49404 (N_49404,N_46892,N_46494);
xor U49405 (N_49405,N_45735,N_45517);
or U49406 (N_49406,N_46787,N_45168);
nor U49407 (N_49407,N_46897,N_45555);
or U49408 (N_49408,N_45002,N_45948);
nor U49409 (N_49409,N_46472,N_47098);
xor U49410 (N_49410,N_47221,N_46710);
xnor U49411 (N_49411,N_45395,N_46090);
and U49412 (N_49412,N_45973,N_46909);
nand U49413 (N_49413,N_45254,N_46146);
nor U49414 (N_49414,N_46225,N_45159);
nand U49415 (N_49415,N_46772,N_45098);
or U49416 (N_49416,N_45706,N_46557);
xor U49417 (N_49417,N_46574,N_46129);
nand U49418 (N_49418,N_46711,N_45245);
nor U49419 (N_49419,N_46362,N_47396);
nor U49420 (N_49420,N_46153,N_46315);
xor U49421 (N_49421,N_46096,N_46848);
or U49422 (N_49422,N_47305,N_46860);
and U49423 (N_49423,N_45626,N_46083);
xor U49424 (N_49424,N_45170,N_47124);
or U49425 (N_49425,N_45912,N_45479);
and U49426 (N_49426,N_47248,N_45545);
xnor U49427 (N_49427,N_46247,N_47363);
or U49428 (N_49428,N_46632,N_45118);
and U49429 (N_49429,N_45327,N_47188);
or U49430 (N_49430,N_46864,N_45830);
nor U49431 (N_49431,N_45574,N_45061);
nor U49432 (N_49432,N_46831,N_46992);
xnor U49433 (N_49433,N_45056,N_47163);
and U49434 (N_49434,N_45274,N_45988);
nand U49435 (N_49435,N_46057,N_47300);
nor U49436 (N_49436,N_47489,N_46306);
or U49437 (N_49437,N_46442,N_45517);
xor U49438 (N_49438,N_45879,N_47380);
xor U49439 (N_49439,N_46991,N_45347);
nor U49440 (N_49440,N_46262,N_45638);
or U49441 (N_49441,N_45187,N_46785);
nor U49442 (N_49442,N_45895,N_47150);
or U49443 (N_49443,N_46634,N_47244);
and U49444 (N_49444,N_46599,N_45624);
or U49445 (N_49445,N_45151,N_45429);
xnor U49446 (N_49446,N_46335,N_45980);
or U49447 (N_49447,N_45233,N_46879);
and U49448 (N_49448,N_45596,N_47050);
and U49449 (N_49449,N_45162,N_45486);
xnor U49450 (N_49450,N_46507,N_45805);
nor U49451 (N_49451,N_45367,N_46016);
and U49452 (N_49452,N_46439,N_46276);
nor U49453 (N_49453,N_46295,N_47195);
xor U49454 (N_49454,N_45780,N_47177);
and U49455 (N_49455,N_46594,N_46891);
xnor U49456 (N_49456,N_45853,N_47226);
or U49457 (N_49457,N_45126,N_46329);
and U49458 (N_49458,N_47382,N_46050);
xor U49459 (N_49459,N_46226,N_46614);
or U49460 (N_49460,N_46584,N_46641);
nand U49461 (N_49461,N_45597,N_46217);
nand U49462 (N_49462,N_47231,N_47464);
xnor U49463 (N_49463,N_45362,N_45212);
or U49464 (N_49464,N_46240,N_47029);
nor U49465 (N_49465,N_47063,N_47139);
nand U49466 (N_49466,N_45750,N_47224);
and U49467 (N_49467,N_46864,N_46440);
and U49468 (N_49468,N_46228,N_46089);
or U49469 (N_49469,N_46848,N_46966);
and U49470 (N_49470,N_45720,N_46568);
xor U49471 (N_49471,N_46049,N_46533);
and U49472 (N_49472,N_45960,N_45170);
nor U49473 (N_49473,N_47054,N_46933);
nand U49474 (N_49474,N_45441,N_45145);
or U49475 (N_49475,N_46811,N_46167);
and U49476 (N_49476,N_47195,N_46457);
nand U49477 (N_49477,N_46179,N_47144);
or U49478 (N_49478,N_45723,N_47333);
nand U49479 (N_49479,N_45095,N_46055);
and U49480 (N_49480,N_46505,N_45879);
nor U49481 (N_49481,N_47334,N_46844);
nand U49482 (N_49482,N_46634,N_46334);
or U49483 (N_49483,N_46726,N_46063);
xor U49484 (N_49484,N_46956,N_46598);
nor U49485 (N_49485,N_47122,N_45786);
and U49486 (N_49486,N_45492,N_46764);
or U49487 (N_49487,N_47061,N_45231);
xor U49488 (N_49488,N_46074,N_45967);
nor U49489 (N_49489,N_46565,N_46392);
or U49490 (N_49490,N_45953,N_46212);
xnor U49491 (N_49491,N_46073,N_46162);
nor U49492 (N_49492,N_45427,N_45733);
and U49493 (N_49493,N_45140,N_45821);
and U49494 (N_49494,N_47357,N_46740);
nor U49495 (N_49495,N_45646,N_46047);
and U49496 (N_49496,N_46701,N_46026);
nand U49497 (N_49497,N_47084,N_46607);
xor U49498 (N_49498,N_46258,N_45859);
nor U49499 (N_49499,N_46070,N_46884);
nor U49500 (N_49500,N_45866,N_47434);
and U49501 (N_49501,N_46780,N_45267);
and U49502 (N_49502,N_46689,N_45180);
nand U49503 (N_49503,N_47298,N_45194);
xnor U49504 (N_49504,N_45339,N_45499);
and U49505 (N_49505,N_47145,N_46496);
nor U49506 (N_49506,N_46691,N_45201);
nor U49507 (N_49507,N_46619,N_47403);
and U49508 (N_49508,N_46188,N_47338);
xor U49509 (N_49509,N_45279,N_45899);
xor U49510 (N_49510,N_45082,N_46876);
xor U49511 (N_49511,N_46715,N_45693);
xnor U49512 (N_49512,N_45154,N_46943);
or U49513 (N_49513,N_45926,N_45339);
nor U49514 (N_49514,N_45798,N_47006);
or U49515 (N_49515,N_45307,N_46993);
or U49516 (N_49516,N_45540,N_45720);
and U49517 (N_49517,N_45039,N_45372);
and U49518 (N_49518,N_45369,N_45115);
or U49519 (N_49519,N_45613,N_47101);
and U49520 (N_49520,N_45771,N_45316);
nor U49521 (N_49521,N_47120,N_45921);
nor U49522 (N_49522,N_45814,N_46998);
and U49523 (N_49523,N_47414,N_46547);
or U49524 (N_49524,N_45600,N_46023);
xor U49525 (N_49525,N_46915,N_46955);
nor U49526 (N_49526,N_46280,N_45827);
or U49527 (N_49527,N_45249,N_46841);
nor U49528 (N_49528,N_46460,N_47023);
and U49529 (N_49529,N_45489,N_45299);
and U49530 (N_49530,N_45546,N_45067);
and U49531 (N_49531,N_45069,N_45714);
nand U49532 (N_49532,N_46236,N_45643);
nand U49533 (N_49533,N_45439,N_45210);
xnor U49534 (N_49534,N_47476,N_47233);
or U49535 (N_49535,N_47329,N_46395);
or U49536 (N_49536,N_45385,N_46608);
nand U49537 (N_49537,N_47377,N_47452);
or U49538 (N_49538,N_45279,N_45982);
nand U49539 (N_49539,N_46303,N_45219);
nor U49540 (N_49540,N_46594,N_47272);
xnor U49541 (N_49541,N_46393,N_45456);
or U49542 (N_49542,N_45704,N_45238);
or U49543 (N_49543,N_47012,N_45668);
nand U49544 (N_49544,N_45349,N_46966);
xnor U49545 (N_49545,N_46077,N_45189);
and U49546 (N_49546,N_46398,N_46457);
or U49547 (N_49547,N_45092,N_45743);
or U49548 (N_49548,N_45456,N_46860);
or U49549 (N_49549,N_45107,N_47359);
xor U49550 (N_49550,N_46763,N_46525);
and U49551 (N_49551,N_45129,N_45283);
and U49552 (N_49552,N_45134,N_47468);
and U49553 (N_49553,N_45126,N_46130);
and U49554 (N_49554,N_46654,N_46411);
nand U49555 (N_49555,N_46497,N_45347);
xnor U49556 (N_49556,N_46608,N_46225);
xnor U49557 (N_49557,N_45896,N_46162);
xnor U49558 (N_49558,N_46527,N_45521);
or U49559 (N_49559,N_45300,N_46131);
and U49560 (N_49560,N_45749,N_47256);
xor U49561 (N_49561,N_45625,N_45062);
and U49562 (N_49562,N_46080,N_45351);
nand U49563 (N_49563,N_46069,N_45087);
nand U49564 (N_49564,N_47322,N_47023);
nor U49565 (N_49565,N_46865,N_45545);
nand U49566 (N_49566,N_45978,N_45299);
nor U49567 (N_49567,N_46705,N_45115);
nand U49568 (N_49568,N_46669,N_45007);
nand U49569 (N_49569,N_46873,N_46573);
or U49570 (N_49570,N_46554,N_46836);
and U49571 (N_49571,N_46507,N_45732);
nand U49572 (N_49572,N_45455,N_46303);
and U49573 (N_49573,N_45165,N_46071);
xor U49574 (N_49574,N_46427,N_45304);
nor U49575 (N_49575,N_45369,N_45187);
or U49576 (N_49576,N_45637,N_45531);
nand U49577 (N_49577,N_45753,N_45832);
nor U49578 (N_49578,N_45898,N_46016);
xor U49579 (N_49579,N_45135,N_46639);
nand U49580 (N_49580,N_46897,N_46722);
nand U49581 (N_49581,N_46524,N_45287);
xnor U49582 (N_49582,N_46144,N_46975);
or U49583 (N_49583,N_47301,N_46368);
or U49584 (N_49584,N_45760,N_46989);
nor U49585 (N_49585,N_46095,N_45203);
and U49586 (N_49586,N_47089,N_45055);
nor U49587 (N_49587,N_46813,N_46008);
or U49588 (N_49588,N_46067,N_45601);
xor U49589 (N_49589,N_45380,N_46283);
nor U49590 (N_49590,N_47316,N_47018);
nand U49591 (N_49591,N_47460,N_46779);
nor U49592 (N_49592,N_47107,N_46172);
and U49593 (N_49593,N_46845,N_45143);
nor U49594 (N_49594,N_46488,N_45996);
nand U49595 (N_49595,N_46698,N_46945);
or U49596 (N_49596,N_46448,N_45643);
and U49597 (N_49597,N_46034,N_46165);
nand U49598 (N_49598,N_47265,N_47204);
or U49599 (N_49599,N_46261,N_47305);
xor U49600 (N_49600,N_46866,N_46028);
nor U49601 (N_49601,N_47480,N_45303);
nor U49602 (N_49602,N_47321,N_46952);
nand U49603 (N_49603,N_45806,N_46387);
nand U49604 (N_49604,N_47461,N_45474);
nand U49605 (N_49605,N_45897,N_46641);
nand U49606 (N_49606,N_46726,N_46482);
nand U49607 (N_49607,N_45899,N_45506);
or U49608 (N_49608,N_45740,N_46810);
and U49609 (N_49609,N_46884,N_45195);
nor U49610 (N_49610,N_47233,N_45510);
nand U49611 (N_49611,N_47489,N_46184);
xnor U49612 (N_49612,N_45672,N_46617);
nand U49613 (N_49613,N_45742,N_45604);
nand U49614 (N_49614,N_47017,N_46994);
or U49615 (N_49615,N_46095,N_45102);
and U49616 (N_49616,N_45315,N_45481);
xor U49617 (N_49617,N_47251,N_47060);
nor U49618 (N_49618,N_47318,N_45205);
or U49619 (N_49619,N_45258,N_45615);
nor U49620 (N_49620,N_46368,N_46422);
xnor U49621 (N_49621,N_46373,N_47249);
and U49622 (N_49622,N_47076,N_46858);
or U49623 (N_49623,N_46117,N_46362);
and U49624 (N_49624,N_45025,N_45353);
and U49625 (N_49625,N_46565,N_45967);
xor U49626 (N_49626,N_47420,N_45439);
nand U49627 (N_49627,N_46015,N_46423);
nand U49628 (N_49628,N_46181,N_46075);
and U49629 (N_49629,N_47134,N_45365);
xnor U49630 (N_49630,N_46578,N_45669);
nand U49631 (N_49631,N_47489,N_46647);
xnor U49632 (N_49632,N_46001,N_46893);
or U49633 (N_49633,N_45873,N_46749);
nand U49634 (N_49634,N_45056,N_47221);
xnor U49635 (N_49635,N_46577,N_46366);
xor U49636 (N_49636,N_46330,N_47194);
nor U49637 (N_49637,N_45772,N_45666);
nand U49638 (N_49638,N_45322,N_45066);
nand U49639 (N_49639,N_46715,N_46530);
nand U49640 (N_49640,N_45133,N_45408);
or U49641 (N_49641,N_45124,N_47287);
nor U49642 (N_49642,N_45975,N_45971);
or U49643 (N_49643,N_46183,N_45997);
nor U49644 (N_49644,N_45368,N_46004);
or U49645 (N_49645,N_45069,N_47180);
nand U49646 (N_49646,N_46566,N_46339);
or U49647 (N_49647,N_47133,N_46108);
nor U49648 (N_49648,N_46074,N_47495);
nand U49649 (N_49649,N_46298,N_46990);
nand U49650 (N_49650,N_45664,N_45662);
or U49651 (N_49651,N_46118,N_47339);
or U49652 (N_49652,N_46806,N_46152);
xor U49653 (N_49653,N_45836,N_46950);
and U49654 (N_49654,N_45985,N_47109);
and U49655 (N_49655,N_46205,N_47191);
nand U49656 (N_49656,N_45028,N_45898);
nor U49657 (N_49657,N_45235,N_46007);
nor U49658 (N_49658,N_45706,N_46789);
nor U49659 (N_49659,N_45160,N_45745);
nor U49660 (N_49660,N_47179,N_45314);
and U49661 (N_49661,N_46676,N_47460);
nor U49662 (N_49662,N_46878,N_46721);
and U49663 (N_49663,N_46334,N_47194);
or U49664 (N_49664,N_47393,N_45473);
xnor U49665 (N_49665,N_45053,N_45554);
nor U49666 (N_49666,N_46102,N_46724);
or U49667 (N_49667,N_45443,N_45624);
xnor U49668 (N_49668,N_45729,N_46183);
nor U49669 (N_49669,N_47178,N_45686);
xor U49670 (N_49670,N_45207,N_45935);
nand U49671 (N_49671,N_46601,N_45978);
nand U49672 (N_49672,N_47275,N_46846);
nor U49673 (N_49673,N_46641,N_45400);
nand U49674 (N_49674,N_46926,N_46911);
xnor U49675 (N_49675,N_47392,N_46803);
xor U49676 (N_49676,N_45764,N_46413);
and U49677 (N_49677,N_45976,N_46366);
nand U49678 (N_49678,N_45354,N_45167);
or U49679 (N_49679,N_45154,N_47314);
nand U49680 (N_49680,N_45745,N_45607);
or U49681 (N_49681,N_46851,N_46792);
nor U49682 (N_49682,N_45372,N_45925);
xor U49683 (N_49683,N_46184,N_45121);
nor U49684 (N_49684,N_46547,N_45672);
or U49685 (N_49685,N_46589,N_45539);
or U49686 (N_49686,N_47326,N_45062);
nand U49687 (N_49687,N_46918,N_46530);
nand U49688 (N_49688,N_46660,N_46511);
nor U49689 (N_49689,N_46448,N_46387);
nor U49690 (N_49690,N_47384,N_45137);
or U49691 (N_49691,N_47295,N_46792);
or U49692 (N_49692,N_46699,N_45521);
nand U49693 (N_49693,N_46599,N_45510);
nand U49694 (N_49694,N_46418,N_46054);
or U49695 (N_49695,N_45688,N_47075);
and U49696 (N_49696,N_46129,N_46572);
xnor U49697 (N_49697,N_46199,N_45093);
and U49698 (N_49698,N_47216,N_46829);
and U49699 (N_49699,N_46010,N_45513);
or U49700 (N_49700,N_47425,N_47479);
or U49701 (N_49701,N_46855,N_46964);
and U49702 (N_49702,N_45050,N_46620);
or U49703 (N_49703,N_45315,N_47314);
and U49704 (N_49704,N_45755,N_45110);
nand U49705 (N_49705,N_45375,N_45678);
nor U49706 (N_49706,N_46234,N_45653);
nand U49707 (N_49707,N_45452,N_47018);
xor U49708 (N_49708,N_47181,N_45634);
nor U49709 (N_49709,N_45797,N_46037);
and U49710 (N_49710,N_46118,N_46428);
or U49711 (N_49711,N_46990,N_45816);
nor U49712 (N_49712,N_45108,N_46044);
nor U49713 (N_49713,N_45484,N_46090);
or U49714 (N_49714,N_46624,N_46929);
and U49715 (N_49715,N_46759,N_46910);
or U49716 (N_49716,N_46713,N_45441);
or U49717 (N_49717,N_45127,N_45453);
nor U49718 (N_49718,N_46577,N_47186);
nor U49719 (N_49719,N_46190,N_45062);
nor U49720 (N_49720,N_46888,N_46531);
and U49721 (N_49721,N_46677,N_45198);
nor U49722 (N_49722,N_47195,N_47428);
nand U49723 (N_49723,N_46483,N_47417);
xnor U49724 (N_49724,N_45016,N_46742);
or U49725 (N_49725,N_45573,N_45244);
xnor U49726 (N_49726,N_45337,N_46362);
xnor U49727 (N_49727,N_46010,N_47166);
nand U49728 (N_49728,N_46651,N_47407);
xor U49729 (N_49729,N_46723,N_46273);
nor U49730 (N_49730,N_45474,N_46124);
nor U49731 (N_49731,N_45470,N_46217);
nor U49732 (N_49732,N_45769,N_46587);
nor U49733 (N_49733,N_47075,N_47366);
xor U49734 (N_49734,N_45840,N_46660);
xnor U49735 (N_49735,N_46693,N_45436);
nor U49736 (N_49736,N_46139,N_46712);
nor U49737 (N_49737,N_45457,N_46547);
nor U49738 (N_49738,N_46481,N_46579);
nor U49739 (N_49739,N_45017,N_45934);
nand U49740 (N_49740,N_47066,N_46379);
or U49741 (N_49741,N_46354,N_47275);
or U49742 (N_49742,N_45885,N_46742);
xor U49743 (N_49743,N_45661,N_45981);
or U49744 (N_49744,N_46404,N_45769);
xor U49745 (N_49745,N_45469,N_45084);
nor U49746 (N_49746,N_47372,N_46479);
and U49747 (N_49747,N_46120,N_46777);
or U49748 (N_49748,N_45181,N_46779);
and U49749 (N_49749,N_46215,N_45635);
or U49750 (N_49750,N_45877,N_45265);
nand U49751 (N_49751,N_47496,N_45979);
and U49752 (N_49752,N_45842,N_45304);
xor U49753 (N_49753,N_46804,N_45305);
or U49754 (N_49754,N_46153,N_45052);
nand U49755 (N_49755,N_46824,N_47285);
and U49756 (N_49756,N_45069,N_45007);
nand U49757 (N_49757,N_45989,N_46277);
or U49758 (N_49758,N_47448,N_46505);
and U49759 (N_49759,N_46244,N_46670);
and U49760 (N_49760,N_46037,N_45486);
nor U49761 (N_49761,N_45680,N_45386);
or U49762 (N_49762,N_47422,N_45292);
nand U49763 (N_49763,N_46541,N_46263);
nand U49764 (N_49764,N_46018,N_46687);
and U49765 (N_49765,N_46305,N_46093);
xnor U49766 (N_49766,N_46842,N_46360);
or U49767 (N_49767,N_46775,N_46308);
xnor U49768 (N_49768,N_47395,N_47149);
and U49769 (N_49769,N_46344,N_47302);
and U49770 (N_49770,N_46748,N_45687);
nand U49771 (N_49771,N_46966,N_46442);
nor U49772 (N_49772,N_45823,N_47016);
xor U49773 (N_49773,N_46773,N_46889);
or U49774 (N_49774,N_46810,N_45507);
nand U49775 (N_49775,N_47398,N_47016);
and U49776 (N_49776,N_45457,N_46362);
and U49777 (N_49777,N_46303,N_45023);
and U49778 (N_49778,N_46991,N_46224);
nand U49779 (N_49779,N_46556,N_45540);
and U49780 (N_49780,N_46257,N_45130);
xor U49781 (N_49781,N_47202,N_45963);
and U49782 (N_49782,N_47349,N_45014);
nand U49783 (N_49783,N_47079,N_45264);
nor U49784 (N_49784,N_46659,N_46266);
or U49785 (N_49785,N_46561,N_46691);
nor U49786 (N_49786,N_46878,N_45022);
or U49787 (N_49787,N_45351,N_45475);
or U49788 (N_49788,N_46405,N_45655);
nor U49789 (N_49789,N_47104,N_47386);
xnor U49790 (N_49790,N_45541,N_47002);
nand U49791 (N_49791,N_45590,N_45403);
and U49792 (N_49792,N_47429,N_46638);
nand U49793 (N_49793,N_45430,N_46641);
and U49794 (N_49794,N_46617,N_45848);
nor U49795 (N_49795,N_45336,N_45979);
nor U49796 (N_49796,N_47291,N_46897);
and U49797 (N_49797,N_46545,N_46962);
and U49798 (N_49798,N_46953,N_45006);
nand U49799 (N_49799,N_46364,N_45844);
and U49800 (N_49800,N_46274,N_46059);
or U49801 (N_49801,N_45000,N_46734);
nor U49802 (N_49802,N_45065,N_47232);
nand U49803 (N_49803,N_46712,N_46676);
xor U49804 (N_49804,N_47416,N_46743);
or U49805 (N_49805,N_47132,N_47138);
nand U49806 (N_49806,N_46922,N_45185);
nor U49807 (N_49807,N_46491,N_45285);
and U49808 (N_49808,N_47315,N_46590);
and U49809 (N_49809,N_45783,N_46903);
xnor U49810 (N_49810,N_47441,N_45254);
and U49811 (N_49811,N_46470,N_47475);
and U49812 (N_49812,N_45700,N_45549);
nand U49813 (N_49813,N_47467,N_45227);
nor U49814 (N_49814,N_46661,N_46108);
or U49815 (N_49815,N_46002,N_46929);
and U49816 (N_49816,N_47339,N_45868);
and U49817 (N_49817,N_46058,N_45545);
xor U49818 (N_49818,N_46667,N_45061);
or U49819 (N_49819,N_45520,N_46939);
or U49820 (N_49820,N_45063,N_46265);
or U49821 (N_49821,N_45296,N_46937);
nor U49822 (N_49822,N_47305,N_45530);
nand U49823 (N_49823,N_45450,N_47064);
and U49824 (N_49824,N_47465,N_46606);
xor U49825 (N_49825,N_45485,N_46967);
and U49826 (N_49826,N_46339,N_46326);
xor U49827 (N_49827,N_45717,N_46675);
nand U49828 (N_49828,N_46938,N_45124);
or U49829 (N_49829,N_46294,N_47124);
nor U49830 (N_49830,N_45718,N_46246);
xnor U49831 (N_49831,N_45951,N_45984);
xnor U49832 (N_49832,N_46867,N_45822);
or U49833 (N_49833,N_46726,N_45407);
and U49834 (N_49834,N_46258,N_45753);
or U49835 (N_49835,N_45077,N_45030);
or U49836 (N_49836,N_45647,N_45072);
xnor U49837 (N_49837,N_46383,N_45052);
nand U49838 (N_49838,N_46198,N_45744);
xor U49839 (N_49839,N_45609,N_47062);
or U49840 (N_49840,N_46393,N_45723);
and U49841 (N_49841,N_46772,N_46962);
nand U49842 (N_49842,N_46376,N_45106);
xor U49843 (N_49843,N_45750,N_46763);
nand U49844 (N_49844,N_47389,N_47390);
and U49845 (N_49845,N_45825,N_47373);
nand U49846 (N_49846,N_46677,N_45645);
nor U49847 (N_49847,N_46434,N_47158);
and U49848 (N_49848,N_46501,N_46779);
and U49849 (N_49849,N_45419,N_46600);
nand U49850 (N_49850,N_46325,N_47249);
nor U49851 (N_49851,N_46535,N_45887);
xnor U49852 (N_49852,N_45152,N_45726);
and U49853 (N_49853,N_46279,N_46665);
xnor U49854 (N_49854,N_46412,N_46133);
xor U49855 (N_49855,N_46583,N_47252);
and U49856 (N_49856,N_47049,N_47435);
or U49857 (N_49857,N_46265,N_45698);
or U49858 (N_49858,N_45815,N_46703);
nor U49859 (N_49859,N_46267,N_47339);
and U49860 (N_49860,N_46094,N_47056);
and U49861 (N_49861,N_47242,N_45959);
or U49862 (N_49862,N_45802,N_46480);
and U49863 (N_49863,N_46048,N_45006);
nor U49864 (N_49864,N_45563,N_46981);
nand U49865 (N_49865,N_46728,N_47132);
or U49866 (N_49866,N_46274,N_46535);
or U49867 (N_49867,N_46724,N_45384);
xnor U49868 (N_49868,N_46537,N_45803);
nor U49869 (N_49869,N_45593,N_45225);
or U49870 (N_49870,N_45393,N_45700);
xor U49871 (N_49871,N_46968,N_46566);
nand U49872 (N_49872,N_45612,N_47018);
nor U49873 (N_49873,N_47080,N_46942);
nor U49874 (N_49874,N_45192,N_47212);
nand U49875 (N_49875,N_47455,N_47375);
nor U49876 (N_49876,N_47209,N_45451);
xor U49877 (N_49877,N_45894,N_47365);
xor U49878 (N_49878,N_46778,N_45439);
nor U49879 (N_49879,N_47001,N_46800);
and U49880 (N_49880,N_47324,N_46998);
nor U49881 (N_49881,N_47372,N_46737);
nor U49882 (N_49882,N_45281,N_47364);
xnor U49883 (N_49883,N_45379,N_46797);
nor U49884 (N_49884,N_46770,N_47269);
nand U49885 (N_49885,N_45539,N_47385);
nand U49886 (N_49886,N_47431,N_46002);
nor U49887 (N_49887,N_45151,N_47096);
and U49888 (N_49888,N_47299,N_47363);
xnor U49889 (N_49889,N_46632,N_45946);
nand U49890 (N_49890,N_46374,N_45318);
and U49891 (N_49891,N_45823,N_47119);
xor U49892 (N_49892,N_45337,N_47340);
and U49893 (N_49893,N_46064,N_46276);
xor U49894 (N_49894,N_47239,N_45758);
or U49895 (N_49895,N_46513,N_45739);
xnor U49896 (N_49896,N_46121,N_45530);
nor U49897 (N_49897,N_46102,N_47153);
nor U49898 (N_49898,N_47380,N_47029);
or U49899 (N_49899,N_46567,N_46911);
or U49900 (N_49900,N_45743,N_46163);
nand U49901 (N_49901,N_46199,N_46936);
xor U49902 (N_49902,N_46576,N_45916);
and U49903 (N_49903,N_45595,N_45283);
nor U49904 (N_49904,N_45578,N_46527);
or U49905 (N_49905,N_45327,N_47078);
xnor U49906 (N_49906,N_45661,N_47082);
xnor U49907 (N_49907,N_45122,N_46145);
nand U49908 (N_49908,N_46354,N_45531);
xnor U49909 (N_49909,N_46188,N_46140);
nand U49910 (N_49910,N_47207,N_45937);
or U49911 (N_49911,N_45884,N_46777);
nand U49912 (N_49912,N_46548,N_46103);
or U49913 (N_49913,N_46500,N_47184);
nand U49914 (N_49914,N_45874,N_46768);
nor U49915 (N_49915,N_47058,N_46554);
or U49916 (N_49916,N_46630,N_45328);
or U49917 (N_49917,N_46911,N_46862);
nand U49918 (N_49918,N_46683,N_45376);
and U49919 (N_49919,N_46801,N_45035);
or U49920 (N_49920,N_46459,N_46564);
and U49921 (N_49921,N_46173,N_47209);
xor U49922 (N_49922,N_46037,N_45684);
nand U49923 (N_49923,N_47409,N_45227);
xnor U49924 (N_49924,N_45043,N_46263);
or U49925 (N_49925,N_46655,N_45416);
or U49926 (N_49926,N_46279,N_45852);
nand U49927 (N_49927,N_47019,N_47388);
nor U49928 (N_49928,N_45764,N_47221);
and U49929 (N_49929,N_47477,N_45459);
xnor U49930 (N_49930,N_46660,N_46117);
xor U49931 (N_49931,N_45209,N_45615);
or U49932 (N_49932,N_45383,N_45074);
nor U49933 (N_49933,N_45656,N_46756);
xor U49934 (N_49934,N_46734,N_45646);
or U49935 (N_49935,N_45345,N_45821);
nand U49936 (N_49936,N_47473,N_45565);
xor U49937 (N_49937,N_46816,N_45427);
and U49938 (N_49938,N_45771,N_45085);
xor U49939 (N_49939,N_46647,N_45973);
and U49940 (N_49940,N_46537,N_47280);
or U49941 (N_49941,N_46580,N_47240);
nor U49942 (N_49942,N_46920,N_45603);
and U49943 (N_49943,N_45986,N_46493);
and U49944 (N_49944,N_45235,N_45179);
nand U49945 (N_49945,N_46461,N_47205);
nor U49946 (N_49946,N_45330,N_46190);
and U49947 (N_49947,N_46408,N_45540);
nand U49948 (N_49948,N_47449,N_47026);
and U49949 (N_49949,N_45678,N_45029);
nand U49950 (N_49950,N_45753,N_45461);
or U49951 (N_49951,N_45920,N_45779);
or U49952 (N_49952,N_46870,N_47307);
nor U49953 (N_49953,N_45772,N_46868);
and U49954 (N_49954,N_45869,N_46223);
or U49955 (N_49955,N_46707,N_46687);
xnor U49956 (N_49956,N_46224,N_46739);
or U49957 (N_49957,N_47269,N_46839);
xor U49958 (N_49958,N_46132,N_46343);
nor U49959 (N_49959,N_46616,N_45110);
nor U49960 (N_49960,N_45507,N_45459);
and U49961 (N_49961,N_46888,N_45040);
or U49962 (N_49962,N_46625,N_45793);
nor U49963 (N_49963,N_46921,N_46968);
nand U49964 (N_49964,N_46805,N_46403);
xor U49965 (N_49965,N_45414,N_47438);
nand U49966 (N_49966,N_47015,N_45154);
nand U49967 (N_49967,N_45126,N_47437);
xnor U49968 (N_49968,N_45084,N_46414);
xnor U49969 (N_49969,N_45211,N_47233);
nand U49970 (N_49970,N_45794,N_46174);
nand U49971 (N_49971,N_45039,N_45952);
and U49972 (N_49972,N_46537,N_45736);
nand U49973 (N_49973,N_46283,N_46597);
xnor U49974 (N_49974,N_47039,N_45644);
or U49975 (N_49975,N_47429,N_45176);
and U49976 (N_49976,N_46821,N_46536);
nand U49977 (N_49977,N_46425,N_45898);
nor U49978 (N_49978,N_45475,N_45069);
and U49979 (N_49979,N_47386,N_46431);
nand U49980 (N_49980,N_47144,N_45297);
nor U49981 (N_49981,N_45147,N_46161);
nand U49982 (N_49982,N_47190,N_46487);
or U49983 (N_49983,N_45085,N_46773);
and U49984 (N_49984,N_45989,N_45303);
nor U49985 (N_49985,N_45362,N_47193);
and U49986 (N_49986,N_47352,N_46190);
or U49987 (N_49987,N_46496,N_46656);
xnor U49988 (N_49988,N_47309,N_45582);
or U49989 (N_49989,N_46375,N_46060);
and U49990 (N_49990,N_47293,N_46798);
and U49991 (N_49991,N_45138,N_47411);
xnor U49992 (N_49992,N_45267,N_46413);
and U49993 (N_49993,N_45099,N_46315);
xnor U49994 (N_49994,N_45878,N_45448);
nand U49995 (N_49995,N_45769,N_47364);
xor U49996 (N_49996,N_46161,N_46517);
or U49997 (N_49997,N_45915,N_45979);
xnor U49998 (N_49998,N_46071,N_46450);
nor U49999 (N_49999,N_46351,N_47174);
or UO_0 (O_0,N_49634,N_49669);
and UO_1 (O_1,N_49788,N_48331);
and UO_2 (O_2,N_49495,N_47835);
xor UO_3 (O_3,N_49789,N_47674);
nor UO_4 (O_4,N_48425,N_48947);
nand UO_5 (O_5,N_49313,N_47891);
and UO_6 (O_6,N_49794,N_47780);
xor UO_7 (O_7,N_49717,N_49890);
or UO_8 (O_8,N_48574,N_49768);
nand UO_9 (O_9,N_48495,N_47613);
xor UO_10 (O_10,N_48522,N_47616);
xor UO_11 (O_11,N_48848,N_47562);
nand UO_12 (O_12,N_48176,N_48036);
xnor UO_13 (O_13,N_48248,N_47718);
xnor UO_14 (O_14,N_48695,N_47893);
and UO_15 (O_15,N_48724,N_48198);
or UO_16 (O_16,N_48426,N_47501);
and UO_17 (O_17,N_48090,N_49830);
nand UO_18 (O_18,N_49976,N_47820);
nand UO_19 (O_19,N_48776,N_47691);
nor UO_20 (O_20,N_47945,N_48725);
or UO_21 (O_21,N_49998,N_49568);
xor UO_22 (O_22,N_49737,N_49918);
xor UO_23 (O_23,N_49856,N_48917);
xnor UO_24 (O_24,N_47715,N_49384);
and UO_25 (O_25,N_47664,N_49652);
and UO_26 (O_26,N_49999,N_49357);
or UO_27 (O_27,N_49572,N_48301);
nor UO_28 (O_28,N_47872,N_47581);
nor UO_29 (O_29,N_48847,N_49702);
and UO_30 (O_30,N_49287,N_49651);
or UO_31 (O_31,N_47941,N_49847);
or UO_32 (O_32,N_48812,N_49969);
or UO_33 (O_33,N_48702,N_49275);
xnor UO_34 (O_34,N_47589,N_49136);
nand UO_35 (O_35,N_49104,N_49885);
nor UO_36 (O_36,N_47964,N_49808);
and UO_37 (O_37,N_48743,N_48335);
and UO_38 (O_38,N_49750,N_49538);
xnor UO_39 (O_39,N_49775,N_49234);
nor UO_40 (O_40,N_48348,N_48011);
nor UO_41 (O_41,N_49195,N_48570);
or UO_42 (O_42,N_48329,N_49564);
and UO_43 (O_43,N_48544,N_48951);
xnor UO_44 (O_44,N_49601,N_49403);
and UO_45 (O_45,N_49837,N_47905);
xor UO_46 (O_46,N_47706,N_48799);
nor UO_47 (O_47,N_48444,N_49467);
and UO_48 (O_48,N_49628,N_47742);
nand UO_49 (O_49,N_48611,N_49552);
nor UO_50 (O_50,N_47770,N_48406);
and UO_51 (O_51,N_48673,N_47607);
and UO_52 (O_52,N_48212,N_49703);
nor UO_53 (O_53,N_49610,N_49282);
and UO_54 (O_54,N_49945,N_47600);
and UO_55 (O_55,N_48370,N_48551);
or UO_56 (O_56,N_48225,N_47594);
nand UO_57 (O_57,N_49807,N_49631);
nor UO_58 (O_58,N_49835,N_48085);
nand UO_59 (O_59,N_48565,N_48018);
nor UO_60 (O_60,N_49772,N_47752);
or UO_61 (O_61,N_49370,N_47663);
nand UO_62 (O_62,N_49782,N_49562);
xor UO_63 (O_63,N_49710,N_49230);
or UO_64 (O_64,N_48784,N_49249);
xor UO_65 (O_65,N_48572,N_47885);
xor UO_66 (O_66,N_48906,N_49067);
xor UO_67 (O_67,N_47727,N_47703);
and UO_68 (O_68,N_47816,N_48648);
nand UO_69 (O_69,N_49225,N_48150);
and UO_70 (O_70,N_49490,N_48671);
xnor UO_71 (O_71,N_48427,N_48942);
nand UO_72 (O_72,N_47667,N_48638);
or UO_73 (O_73,N_49845,N_49368);
nand UO_74 (O_74,N_49228,N_48059);
nand UO_75 (O_75,N_49217,N_49585);
and UO_76 (O_76,N_49209,N_49690);
xor UO_77 (O_77,N_48435,N_48775);
xor UO_78 (O_78,N_49781,N_48726);
and UO_79 (O_79,N_49280,N_48626);
or UO_80 (O_80,N_48106,N_48378);
or UO_81 (O_81,N_48629,N_49365);
nor UO_82 (O_82,N_49901,N_48490);
nor UO_83 (O_83,N_48834,N_49107);
nor UO_84 (O_84,N_47712,N_48468);
nor UO_85 (O_85,N_48622,N_47505);
or UO_86 (O_86,N_49747,N_47684);
or UO_87 (O_87,N_47856,N_49689);
xor UO_88 (O_88,N_48679,N_48575);
and UO_89 (O_89,N_49617,N_48911);
xnor UO_90 (O_90,N_48828,N_48524);
and UO_91 (O_91,N_48571,N_47847);
and UO_92 (O_92,N_49298,N_49135);
or UO_93 (O_93,N_49472,N_48956);
nand UO_94 (O_94,N_47629,N_49052);
or UO_95 (O_95,N_49510,N_47588);
nand UO_96 (O_96,N_48503,N_47568);
and UO_97 (O_97,N_49650,N_47697);
and UO_98 (O_98,N_49148,N_48669);
nand UO_99 (O_99,N_48430,N_47688);
xor UO_100 (O_100,N_47982,N_48485);
or UO_101 (O_101,N_47827,N_48417);
nand UO_102 (O_102,N_47965,N_49066);
nand UO_103 (O_103,N_48636,N_48904);
or UO_104 (O_104,N_49749,N_47782);
nand UO_105 (O_105,N_47639,N_48149);
nor UO_106 (O_106,N_48082,N_49959);
and UO_107 (O_107,N_49192,N_47832);
or UO_108 (O_108,N_48664,N_47519);
xnor UO_109 (O_109,N_49680,N_48445);
xnor UO_110 (O_110,N_49663,N_47615);
nand UO_111 (O_111,N_49711,N_47755);
and UO_112 (O_112,N_48609,N_47644);
nand UO_113 (O_113,N_48122,N_49700);
xor UO_114 (O_114,N_48344,N_49972);
nor UO_115 (O_115,N_49765,N_49397);
nand UO_116 (O_116,N_49262,N_49461);
xor UO_117 (O_117,N_49960,N_48305);
and UO_118 (O_118,N_48761,N_48438);
nand UO_119 (O_119,N_47554,N_48965);
or UO_120 (O_120,N_47537,N_49968);
xor UO_121 (O_121,N_47636,N_49730);
xnor UO_122 (O_122,N_49787,N_48578);
or UO_123 (O_123,N_49991,N_48778);
or UO_124 (O_124,N_49425,N_48589);
or UO_125 (O_125,N_47928,N_47936);
nand UO_126 (O_126,N_49762,N_48733);
nor UO_127 (O_127,N_49222,N_49798);
xor UO_128 (O_128,N_48088,N_47753);
or UO_129 (O_129,N_48857,N_48160);
and UO_130 (O_130,N_48974,N_47888);
or UO_131 (O_131,N_48976,N_49994);
xor UO_132 (O_132,N_48772,N_47987);
nand UO_133 (O_133,N_49134,N_48236);
xor UO_134 (O_134,N_48294,N_48549);
nor UO_135 (O_135,N_49892,N_49076);
or UO_136 (O_136,N_49696,N_47592);
nand UO_137 (O_137,N_48306,N_48615);
nand UO_138 (O_138,N_48759,N_49598);
nand UO_139 (O_139,N_47808,N_49444);
or UO_140 (O_140,N_48890,N_49074);
and UO_141 (O_141,N_48881,N_49944);
or UO_142 (O_142,N_48252,N_48810);
nand UO_143 (O_143,N_48140,N_49408);
nor UO_144 (O_144,N_49919,N_49253);
or UO_145 (O_145,N_48498,N_48732);
nor UO_146 (O_146,N_47678,N_49031);
or UO_147 (O_147,N_49186,N_49530);
or UO_148 (O_148,N_47989,N_48270);
or UO_149 (O_149,N_48255,N_48020);
or UO_150 (O_150,N_47659,N_48148);
and UO_151 (O_151,N_49009,N_49388);
and UO_152 (O_152,N_48802,N_47759);
and UO_153 (O_153,N_48910,N_48533);
xnor UO_154 (O_154,N_48844,N_48142);
or UO_155 (O_155,N_49058,N_49443);
nor UO_156 (O_156,N_47870,N_48944);
xnor UO_157 (O_157,N_48060,N_49200);
or UO_158 (O_158,N_49528,N_49333);
xor UO_159 (O_159,N_47698,N_47617);
nor UO_160 (O_160,N_48573,N_49926);
xor UO_161 (O_161,N_49630,N_49435);
xnor UO_162 (O_162,N_49242,N_48756);
nand UO_163 (O_163,N_48357,N_49424);
nor UO_164 (O_164,N_47791,N_48870);
and UO_165 (O_165,N_47851,N_49288);
or UO_166 (O_166,N_48397,N_48663);
nor UO_167 (O_167,N_49477,N_49439);
and UO_168 (O_168,N_48318,N_47907);
or UO_169 (O_169,N_49805,N_49817);
nor UO_170 (O_170,N_49797,N_47542);
or UO_171 (O_171,N_49422,N_49672);
xor UO_172 (O_172,N_49579,N_49004);
and UO_173 (O_173,N_48026,N_48337);
xor UO_174 (O_174,N_49353,N_48442);
xor UO_175 (O_175,N_49119,N_48658);
and UO_176 (O_176,N_49406,N_48126);
nand UO_177 (O_177,N_48966,N_49311);
or UO_178 (O_178,N_49813,N_49214);
or UO_179 (O_179,N_49592,N_48882);
and UO_180 (O_180,N_49533,N_49973);
nor UO_181 (O_181,N_49014,N_47774);
xnor UO_182 (O_182,N_48083,N_49522);
and UO_183 (O_183,N_49942,N_49984);
xnor UO_184 (O_184,N_47574,N_48672);
or UO_185 (O_185,N_48089,N_48066);
or UO_186 (O_186,N_47878,N_49350);
xnor UO_187 (O_187,N_48271,N_49773);
and UO_188 (O_188,N_48184,N_49733);
or UO_189 (O_189,N_49843,N_48385);
and UO_190 (O_190,N_47834,N_48460);
nand UO_191 (O_191,N_48511,N_49812);
and UO_192 (O_192,N_49433,N_48913);
and UO_193 (O_193,N_48576,N_48437);
nor UO_194 (O_194,N_49643,N_49882);
and UO_195 (O_195,N_49393,N_48798);
nor UO_196 (O_196,N_49305,N_47836);
and UO_197 (O_197,N_49654,N_49922);
xor UO_198 (O_198,N_49716,N_48719);
and UO_199 (O_199,N_49671,N_47601);
nand UO_200 (O_200,N_47572,N_48705);
or UO_201 (O_201,N_49336,N_47794);
xnor UO_202 (O_202,N_49325,N_48390);
nand UO_203 (O_203,N_47829,N_49400);
nand UO_204 (O_204,N_48204,N_49487);
or UO_205 (O_205,N_47988,N_49824);
and UO_206 (O_206,N_47952,N_49500);
nor UO_207 (O_207,N_49011,N_49352);
or UO_208 (O_208,N_47523,N_48620);
or UO_209 (O_209,N_47547,N_48903);
and UO_210 (O_210,N_47733,N_48601);
nand UO_211 (O_211,N_47821,N_48901);
and UO_212 (O_212,N_49641,N_48139);
nor UO_213 (O_213,N_47510,N_49731);
xor UO_214 (O_214,N_48800,N_48037);
or UO_215 (O_215,N_49827,N_47802);
nand UO_216 (O_216,N_48209,N_49905);
nor UO_217 (O_217,N_48831,N_49299);
or UO_218 (O_218,N_49906,N_48053);
nand UO_219 (O_219,N_47894,N_48431);
and UO_220 (O_220,N_48072,N_49168);
nand UO_221 (O_221,N_49895,N_48721);
or UO_222 (O_222,N_49719,N_49339);
or UO_223 (O_223,N_48462,N_47911);
or UO_224 (O_224,N_48228,N_48013);
nor UO_225 (O_225,N_48519,N_48119);
xnor UO_226 (O_226,N_48528,N_47558);
and UO_227 (O_227,N_49129,N_48559);
or UO_228 (O_228,N_47557,N_47853);
and UO_229 (O_229,N_49925,N_47545);
xor UO_230 (O_230,N_49608,N_47979);
xnor UO_231 (O_231,N_47561,N_49402);
or UO_232 (O_232,N_49741,N_49810);
or UO_233 (O_233,N_48830,N_48937);
or UO_234 (O_234,N_48630,N_48550);
xnor UO_235 (O_235,N_49158,N_49875);
nand UO_236 (O_236,N_49611,N_48424);
nand UO_237 (O_237,N_49904,N_48746);
or UO_238 (O_238,N_48720,N_48793);
and UO_239 (O_239,N_48189,N_49923);
xor UO_240 (O_240,N_48593,N_49289);
nand UO_241 (O_241,N_48411,N_49176);
nand UO_242 (O_242,N_48699,N_47506);
or UO_243 (O_243,N_49848,N_48009);
nand UO_244 (O_244,N_47694,N_47998);
xnor UO_245 (O_245,N_47876,N_49975);
nor UO_246 (O_246,N_49887,N_48501);
nand UO_247 (O_247,N_48736,N_48398);
nor UO_248 (O_248,N_49100,N_48824);
nand UO_249 (O_249,N_47981,N_48814);
xnor UO_250 (O_250,N_47809,N_47514);
nor UO_251 (O_251,N_47551,N_47543);
nand UO_252 (O_252,N_47756,N_49092);
and UO_253 (O_253,N_48635,N_49556);
or UO_254 (O_254,N_48166,N_49117);
and UO_255 (O_255,N_48708,N_49012);
nor UO_256 (O_256,N_48553,N_47923);
nor UO_257 (O_257,N_48476,N_49019);
nor UO_258 (O_258,N_48716,N_48299);
or UO_259 (O_259,N_49385,N_49734);
and UO_260 (O_260,N_49331,N_48044);
nand UO_261 (O_261,N_48960,N_49502);
or UO_262 (O_262,N_48447,N_48543);
or UO_263 (O_263,N_49779,N_49484);
or UO_264 (O_264,N_48757,N_48436);
nor UO_265 (O_265,N_48194,N_49769);
nand UO_266 (O_266,N_49886,N_48597);
xnor UO_267 (O_267,N_48779,N_49596);
xor UO_268 (O_268,N_49417,N_48742);
xnor UO_269 (O_269,N_47909,N_48339);
and UO_270 (O_270,N_49532,N_47735);
nor UO_271 (O_271,N_48224,N_48482);
and UO_272 (O_272,N_49981,N_48652);
or UO_273 (O_273,N_49525,N_48540);
xor UO_274 (O_274,N_47977,N_48035);
and UO_275 (O_275,N_47552,N_48675);
xor UO_276 (O_276,N_47749,N_49979);
and UO_277 (O_277,N_48807,N_47502);
xnor UO_278 (O_278,N_49213,N_47689);
and UO_279 (O_279,N_47884,N_48461);
nor UO_280 (O_280,N_48769,N_48165);
and UO_281 (O_281,N_49018,N_49594);
or UO_282 (O_282,N_49446,N_49632);
nor UO_283 (O_283,N_49040,N_47769);
nor UO_284 (O_284,N_47729,N_49237);
or UO_285 (O_285,N_48115,N_47926);
and UO_286 (O_286,N_48826,N_48833);
nor UO_287 (O_287,N_49872,N_49953);
nand UO_288 (O_288,N_49088,N_48939);
xor UO_289 (O_289,N_48446,N_47704);
or UO_290 (O_290,N_49492,N_49606);
nor UO_291 (O_291,N_49952,N_49142);
xnor UO_292 (O_292,N_48595,N_49478);
and UO_293 (O_293,N_49898,N_49414);
nor UO_294 (O_294,N_48213,N_48114);
nor UO_295 (O_295,N_49185,N_47709);
and UO_296 (O_296,N_49266,N_48883);
xor UO_297 (O_297,N_48879,N_48829);
and UO_298 (O_298,N_49553,N_48481);
or UO_299 (O_299,N_49614,N_49770);
nor UO_300 (O_300,N_48324,N_47883);
xor UO_301 (O_301,N_47553,N_49183);
nor UO_302 (O_302,N_47651,N_48354);
nand UO_303 (O_303,N_48872,N_49983);
xor UO_304 (O_304,N_47570,N_49995);
nor UO_305 (O_305,N_49304,N_47806);
nor UO_306 (O_306,N_49364,N_47932);
and UO_307 (O_307,N_47719,N_47968);
xnor UO_308 (O_308,N_48092,N_49448);
and UO_309 (O_309,N_49246,N_48924);
nor UO_310 (O_310,N_48214,N_49701);
and UO_311 (O_311,N_49527,N_48545);
nor UO_312 (O_312,N_49619,N_49196);
xnor UO_313 (O_313,N_49445,N_49583);
nor UO_314 (O_314,N_48471,N_47761);
nand UO_315 (O_315,N_47737,N_49748);
or UO_316 (O_316,N_47889,N_48432);
nor UO_317 (O_317,N_49721,N_47705);
xnor UO_318 (O_318,N_49025,N_49296);
nand UO_319 (O_319,N_47521,N_48369);
xor UO_320 (O_320,N_49429,N_49163);
and UO_321 (O_321,N_47931,N_49753);
and UO_322 (O_322,N_49871,N_48560);
xor UO_323 (O_323,N_48862,N_49174);
nor UO_324 (O_324,N_48986,N_48838);
or UO_325 (O_325,N_49398,N_48731);
nand UO_326 (O_326,N_49034,N_47728);
or UO_327 (O_327,N_49114,N_49269);
or UO_328 (O_328,N_47608,N_48920);
nor UO_329 (O_329,N_49394,N_48584);
xnor UO_330 (O_330,N_49259,N_49274);
xor UO_331 (O_331,N_49561,N_48623);
or UO_332 (O_332,N_48983,N_49577);
xnor UO_333 (O_333,N_47943,N_48741);
nand UO_334 (O_334,N_49109,N_48178);
nor UO_335 (O_335,N_47959,N_48242);
or UO_336 (O_336,N_48005,N_49054);
or UO_337 (O_337,N_49464,N_49850);
or UO_338 (O_338,N_49535,N_47963);
and UO_339 (O_339,N_48347,N_49539);
nand UO_340 (O_340,N_49774,N_49743);
and UO_341 (O_341,N_48617,N_48130);
nor UO_342 (O_342,N_48030,N_48941);
xor UO_343 (O_343,N_49358,N_49233);
and UO_344 (O_344,N_48727,N_48223);
nand UO_345 (O_345,N_47699,N_49876);
or UO_346 (O_346,N_48842,N_49838);
xor UO_347 (O_347,N_47621,N_49308);
and UO_348 (O_348,N_48373,N_49471);
nor UO_349 (O_349,N_47942,N_49566);
and UO_350 (O_350,N_48328,N_49363);
nor UO_351 (O_351,N_48266,N_49440);
nand UO_352 (O_352,N_47530,N_48161);
nor UO_353 (O_353,N_49961,N_48541);
and UO_354 (O_354,N_47680,N_48052);
xor UO_355 (O_355,N_48441,N_49361);
nor UO_356 (O_356,N_48863,N_48116);
xnor UO_357 (O_357,N_48624,N_48867);
or UO_358 (O_358,N_48645,N_47717);
nand UO_359 (O_359,N_48400,N_48456);
nor UO_360 (O_360,N_48309,N_48021);
nand UO_361 (O_361,N_49625,N_48728);
or UO_362 (O_362,N_49957,N_47969);
xor UO_363 (O_363,N_49780,N_48422);
nor UO_364 (O_364,N_48317,N_49754);
nand UO_365 (O_365,N_47813,N_48368);
and UO_366 (O_366,N_47500,N_49373);
and UO_367 (O_367,N_49996,N_48203);
nor UO_368 (O_368,N_47803,N_48386);
or UO_369 (O_369,N_47692,N_48978);
xnor UO_370 (O_370,N_49869,N_48790);
or UO_371 (O_371,N_49581,N_47929);
xor UO_372 (O_372,N_48237,N_48217);
and UO_373 (O_373,N_49714,N_47582);
nand UO_374 (O_374,N_49218,N_49613);
nand UO_375 (O_375,N_49125,N_48680);
nand UO_376 (O_376,N_48892,N_47564);
nand UO_377 (O_377,N_49989,N_49801);
nand UO_378 (O_378,N_48136,N_49574);
nand UO_379 (O_379,N_47677,N_49198);
xor UO_380 (O_380,N_48327,N_49724);
or UO_381 (O_381,N_48621,N_47976);
nand UO_382 (O_382,N_48693,N_47593);
nand UO_383 (O_383,N_49436,N_49524);
or UO_384 (O_384,N_49752,N_49624);
xor UO_385 (O_385,N_48210,N_49191);
or UO_386 (O_386,N_47881,N_47599);
or UO_387 (O_387,N_49226,N_48310);
xor UO_388 (O_388,N_47960,N_48585);
or UO_389 (O_389,N_49518,N_47840);
nand UO_390 (O_390,N_49565,N_49818);
xor UO_391 (O_391,N_48943,N_47586);
xnor UO_392 (O_392,N_48889,N_49924);
xnor UO_393 (O_393,N_47575,N_47711);
or UO_394 (O_394,N_49599,N_48508);
and UO_395 (O_395,N_48326,N_47933);
nand UO_396 (O_396,N_49124,N_47950);
nand UO_397 (O_397,N_49479,N_49793);
xnor UO_398 (O_398,N_49544,N_47906);
xor UO_399 (O_399,N_49958,N_47902);
or UO_400 (O_400,N_48192,N_48396);
nor UO_401 (O_401,N_49369,N_49506);
xor UO_402 (O_402,N_49437,N_49884);
xor UO_403 (O_403,N_49633,N_49459);
nor UO_404 (O_404,N_49697,N_48958);
nor UO_405 (O_405,N_48654,N_47669);
xnor UO_406 (O_406,N_49110,N_49639);
xor UO_407 (O_407,N_49560,N_49591);
and UO_408 (O_408,N_47916,N_48909);
nor UO_409 (O_409,N_49164,N_49016);
xnor UO_410 (O_410,N_48579,N_48646);
and UO_411 (O_411,N_48952,N_49132);
or UO_412 (O_412,N_49851,N_48455);
or UO_413 (O_413,N_48591,N_48234);
nand UO_414 (O_414,N_48325,N_48269);
or UO_415 (O_415,N_48185,N_49783);
nand UO_416 (O_416,N_49473,N_47700);
nor UO_417 (O_417,N_47555,N_48065);
or UO_418 (O_418,N_48345,N_49790);
and UO_419 (O_419,N_47993,N_48016);
xor UO_420 (O_420,N_49795,N_49170);
nand UO_421 (O_421,N_48656,N_48668);
nand UO_422 (O_422,N_48632,N_48649);
or UO_423 (O_423,N_49197,N_48245);
or UO_424 (O_424,N_47672,N_49260);
or UO_425 (O_425,N_49220,N_48866);
nand UO_426 (O_426,N_49194,N_49912);
nand UO_427 (O_427,N_49708,N_49179);
nor UO_428 (O_428,N_49858,N_47640);
xor UO_429 (O_429,N_48667,N_48902);
and UO_430 (O_430,N_49207,N_48938);
or UO_431 (O_431,N_47512,N_48962);
nor UO_432 (O_432,N_48614,N_48118);
nand UO_433 (O_433,N_49413,N_48566);
nor UO_434 (O_434,N_48979,N_47956);
xor UO_435 (O_435,N_48227,N_48916);
or UO_436 (O_436,N_47804,N_47649);
nor UO_437 (O_437,N_48141,N_48758);
and UO_438 (O_438,N_48767,N_48061);
xor UO_439 (O_439,N_48180,N_47790);
or UO_440 (O_440,N_48749,N_49864);
nor UO_441 (O_441,N_47676,N_47620);
nor UO_442 (O_442,N_49030,N_48808);
and UO_443 (O_443,N_49570,N_48860);
nor UO_444 (O_444,N_48312,N_49006);
xor UO_445 (O_445,N_49345,N_49038);
nand UO_446 (O_446,N_48568,N_48521);
and UO_447 (O_447,N_47797,N_47671);
xor UO_448 (O_448,N_48283,N_49636);
xor UO_449 (O_449,N_48280,N_48463);
nand UO_450 (O_450,N_48235,N_49640);
xor UO_451 (O_451,N_48405,N_47522);
xor UO_452 (O_452,N_48489,N_47868);
xnor UO_453 (O_453,N_49949,N_48459);
nor UO_454 (O_454,N_49064,N_48590);
and UO_455 (O_455,N_47722,N_48101);
xor UO_456 (O_456,N_49929,N_47800);
and UO_457 (O_457,N_48592,N_49137);
and UO_458 (O_458,N_48249,N_49022);
nand UO_459 (O_459,N_49354,N_49677);
xor UO_460 (O_460,N_49964,N_48998);
xnor UO_461 (O_461,N_48171,N_48637);
nand UO_462 (O_462,N_48665,N_47540);
nor UO_463 (O_463,N_49381,N_47788);
and UO_464 (O_464,N_48858,N_49335);
nand UO_465 (O_465,N_48969,N_48581);
nand UO_466 (O_466,N_48275,N_49130);
nor UO_467 (O_467,N_48478,N_48949);
and UO_468 (O_468,N_48536,N_49021);
nor UO_469 (O_469,N_47842,N_47643);
xor UO_470 (O_470,N_48651,N_49003);
or UO_471 (O_471,N_47972,N_48316);
nor UO_472 (O_472,N_48027,N_47799);
nor UO_473 (O_473,N_47745,N_48647);
nand UO_474 (O_474,N_47648,N_49239);
xor UO_475 (O_475,N_48413,N_49070);
xor UO_476 (O_476,N_49279,N_48558);
and UO_477 (O_477,N_48694,N_47900);
xnor UO_478 (O_478,N_47548,N_49300);
or UO_479 (O_479,N_49557,N_49656);
xnor UO_480 (O_480,N_49102,N_47930);
or UO_481 (O_481,N_47739,N_48111);
and UO_482 (O_482,N_49878,N_49988);
nor UO_483 (O_483,N_47973,N_48697);
and UO_484 (O_484,N_49224,N_49540);
nor UO_485 (O_485,N_47587,N_48019);
nor UO_486 (O_486,N_49238,N_47645);
nand UO_487 (O_487,N_47508,N_48314);
nand UO_488 (O_488,N_49720,N_48084);
nand UO_489 (O_489,N_48894,N_48097);
xor UO_490 (O_490,N_49943,N_48682);
and UO_491 (O_491,N_49216,N_49569);
xnor UO_492 (O_492,N_49491,N_48100);
and UO_493 (O_493,N_49166,N_49044);
or UO_494 (O_494,N_48710,N_48279);
xor UO_495 (O_495,N_49673,N_49831);
xor UO_496 (O_496,N_49267,N_47638);
xnor UO_497 (O_497,N_48977,N_49615);
nor UO_498 (O_498,N_49203,N_49589);
and UO_499 (O_499,N_49799,N_48359);
or UO_500 (O_500,N_49684,N_49676);
nor UO_501 (O_501,N_49231,N_47897);
and UO_502 (O_502,N_48602,N_49526);
nor UO_503 (O_503,N_48957,N_47880);
nor UO_504 (O_504,N_48268,N_49551);
or UO_505 (O_505,N_47518,N_48113);
xnor UO_506 (O_506,N_49455,N_48067);
nand UO_507 (O_507,N_49938,N_48530);
nor UO_508 (O_508,N_49415,N_49534);
and UO_509 (O_509,N_49160,N_48404);
nand UO_510 (O_510,N_49879,N_47525);
or UO_511 (O_511,N_48674,N_49341);
nand UO_512 (O_512,N_49050,N_48750);
nor UO_513 (O_513,N_47863,N_49096);
or UO_514 (O_514,N_48534,N_48355);
xnor UO_515 (O_515,N_48908,N_48764);
nand UO_516 (O_516,N_49802,N_48263);
or UO_517 (O_517,N_48929,N_47634);
nand UO_518 (O_518,N_49286,N_48817);
and UO_519 (O_519,N_48276,N_48449);
xnor UO_520 (O_520,N_48515,N_47614);
nor UO_521 (O_521,N_49832,N_48313);
nor UO_522 (O_522,N_49877,N_47690);
and UO_523 (O_523,N_49784,N_49997);
nor UO_524 (O_524,N_48439,N_47970);
nor UO_525 (O_525,N_47862,N_48017);
nor UO_526 (O_526,N_48512,N_47624);
nand UO_527 (O_527,N_48897,N_48156);
and UO_528 (O_528,N_48876,N_48465);
and UO_529 (O_529,N_48105,N_49008);
xnor UO_530 (O_530,N_48412,N_48989);
nand UO_531 (O_531,N_47708,N_48231);
nor UO_532 (O_532,N_48492,N_48163);
nand UO_533 (O_533,N_49431,N_47631);
xnor UO_534 (O_534,N_49140,N_48032);
or UO_535 (O_535,N_49057,N_49726);
xor UO_536 (O_536,N_48531,N_47910);
nor UO_537 (O_537,N_48243,N_48290);
or UO_538 (O_538,N_47838,N_48744);
nor UO_539 (O_539,N_47686,N_49699);
and UO_540 (O_540,N_47796,N_48634);
nand UO_541 (O_541,N_48821,N_48984);
nand UO_542 (O_542,N_48968,N_48552);
or UO_543 (O_543,N_47618,N_47875);
nand UO_544 (O_544,N_47927,N_48771);
nor UO_545 (O_545,N_48625,N_48657);
or UO_546 (O_546,N_49974,N_48878);
nor UO_547 (O_547,N_48040,N_47819);
nor UO_548 (O_548,N_49855,N_49985);
xnor UO_549 (O_549,N_48698,N_48109);
or UO_550 (O_550,N_47990,N_47815);
nand UO_551 (O_551,N_49681,N_47653);
xnor UO_552 (O_552,N_48745,N_49815);
nand UO_553 (O_553,N_48296,N_49405);
or UO_554 (O_554,N_49542,N_48048);
xnor UO_555 (O_555,N_48098,N_49758);
nor UO_556 (O_556,N_48755,N_49232);
or UO_557 (O_557,N_48010,N_47939);
and UO_558 (O_558,N_49811,N_47795);
xor UO_559 (O_559,N_49276,N_48349);
nand UO_560 (O_560,N_47556,N_48265);
nor UO_561 (O_561,N_49543,N_49764);
nor UO_562 (O_562,N_49411,N_48803);
xor UO_563 (O_563,N_47903,N_48954);
and UO_564 (O_564,N_47997,N_49272);
nand UO_565 (O_565,N_49638,N_47611);
xor UO_566 (O_566,N_48377,N_49839);
nor UO_567 (O_567,N_49537,N_47504);
xor UO_568 (O_568,N_49891,N_49965);
nand UO_569 (O_569,N_49982,N_49587);
nand UO_570 (O_570,N_49881,N_47527);
and UO_571 (O_571,N_48278,N_47713);
nor UO_572 (O_572,N_48360,N_49616);
xor UO_573 (O_573,N_49120,N_48475);
and UO_574 (O_574,N_48070,N_48479);
nand UO_575 (O_575,N_48055,N_47605);
nand UO_576 (O_576,N_48707,N_49508);
or UO_577 (O_577,N_47983,N_49162);
or UO_578 (O_578,N_48025,N_48391);
or UO_579 (O_579,N_48365,N_49908);
and UO_580 (O_580,N_48786,N_49061);
and UO_581 (O_581,N_48477,N_47954);
nor UO_582 (O_582,N_47660,N_48284);
nor UO_583 (O_583,N_48056,N_48599);
xor UO_584 (O_584,N_49268,N_49893);
xnor UO_585 (O_585,N_49270,N_47904);
and UO_586 (O_586,N_49597,N_49065);
or UO_587 (O_587,N_49558,N_49707);
xor UO_588 (O_588,N_48416,N_47751);
nor UO_589 (O_589,N_49909,N_48421);
or UO_590 (O_590,N_49829,N_48197);
and UO_591 (O_591,N_49840,N_48752);
or UO_592 (O_592,N_49027,N_47913);
nand UO_593 (O_593,N_48953,N_48190);
nor UO_594 (O_594,N_49321,N_49432);
xor UO_595 (O_595,N_49029,N_47563);
nor UO_596 (O_596,N_47971,N_47890);
nor UO_597 (O_597,N_49644,N_49428);
nor UO_598 (O_598,N_49059,N_49612);
nand UO_599 (O_599,N_48473,N_47901);
or UO_600 (O_600,N_49513,N_48520);
or UO_601 (O_601,N_47787,N_49967);
or UO_602 (O_602,N_48509,N_49005);
xnor UO_603 (O_603,N_48900,N_48007);
and UO_604 (O_604,N_47824,N_48959);
nor UO_605 (O_605,N_49852,N_48014);
xor UO_606 (O_606,N_47810,N_49159);
nand UO_607 (O_607,N_48094,N_47886);
xnor UO_608 (O_608,N_47567,N_49853);
and UO_609 (O_609,N_47994,N_48940);
or UO_610 (O_610,N_48073,N_47789);
nor UO_611 (O_611,N_47583,N_49883);
xor UO_612 (O_612,N_48739,N_49048);
nor UO_613 (O_613,N_48823,N_49935);
xnor UO_614 (O_614,N_47873,N_49169);
nor UO_615 (O_615,N_49138,N_49247);
nand UO_616 (O_616,N_47961,N_48076);
nand UO_617 (O_617,N_48666,N_49121);
xor UO_618 (O_618,N_48244,N_49705);
nor UO_619 (O_619,N_49920,N_49629);
xnor UO_620 (O_620,N_49483,N_49201);
nor UO_621 (O_621,N_48760,N_47647);
xnor UO_622 (O_622,N_48627,N_48295);
nor UO_623 (O_623,N_48548,N_48605);
or UO_624 (O_624,N_49037,N_48740);
xor UO_625 (O_625,N_48864,N_48186);
xnor UO_626 (O_626,N_49911,N_47685);
nand UO_627 (O_627,N_48737,N_49682);
xnor UO_628 (O_628,N_48419,N_48921);
xor UO_629 (O_629,N_47566,N_48852);
or UO_630 (O_630,N_48174,N_49778);
and UO_631 (O_631,N_48353,N_48898);
or UO_632 (O_632,N_49692,N_49379);
and UO_633 (O_633,N_49190,N_49177);
or UO_634 (O_634,N_49150,N_49206);
nor UO_635 (O_635,N_49010,N_49695);
nor UO_636 (O_636,N_49356,N_47823);
xor UO_637 (O_637,N_49963,N_48091);
and UO_638 (O_638,N_49307,N_47822);
nor UO_639 (O_639,N_48992,N_49273);
or UO_640 (O_640,N_47786,N_47559);
xnor UO_641 (O_641,N_48062,N_47598);
nor UO_642 (O_642,N_49874,N_48361);
nor UO_643 (O_643,N_48458,N_48333);
xnor UO_644 (O_644,N_47534,N_48818);
and UO_645 (O_645,N_47917,N_48851);
xor UO_646 (O_646,N_47702,N_47517);
nor UO_647 (O_647,N_48029,N_48321);
xnor UO_648 (O_648,N_49603,N_49880);
or UO_649 (O_649,N_49834,N_48117);
nor UO_650 (O_650,N_49127,N_49442);
xnor UO_651 (O_651,N_49825,N_48873);
nand UO_652 (O_652,N_49235,N_48643);
or UO_653 (O_653,N_48660,N_48713);
and UO_654 (O_654,N_49727,N_48922);
or UO_655 (O_655,N_48493,N_49115);
nor UO_656 (O_656,N_49343,N_48208);
or UO_657 (O_657,N_49804,N_48051);
nor UO_658 (O_658,N_48711,N_47953);
xnor UO_659 (O_659,N_47777,N_48781);
and UO_660 (O_660,N_47576,N_49987);
or UO_661 (O_661,N_47738,N_47668);
nand UO_662 (O_662,N_49956,N_48600);
nor UO_663 (O_663,N_48613,N_47516);
xnor UO_664 (O_664,N_48905,N_47841);
or UO_665 (O_665,N_49660,N_48683);
nor UO_666 (O_666,N_48557,N_49468);
nor UO_667 (O_667,N_48024,N_47693);
nor UO_668 (O_668,N_48687,N_48392);
nor UO_669 (O_669,N_48927,N_47665);
xnor UO_670 (O_670,N_48414,N_49015);
nor UO_671 (O_671,N_47736,N_49649);
and UO_672 (O_672,N_49056,N_48454);
and UO_673 (O_673,N_48811,N_47743);
nand UO_674 (O_674,N_49101,N_47503);
nand UO_675 (O_675,N_48580,N_48125);
xnor UO_676 (O_676,N_49978,N_48990);
and UO_677 (O_677,N_48893,N_47716);
nor UO_678 (O_678,N_49863,N_49072);
and UO_679 (O_679,N_48099,N_48789);
or UO_680 (O_680,N_49401,N_48855);
xor UO_681 (O_681,N_48429,N_49451);
nor UO_682 (O_682,N_49359,N_48448);
or UO_683 (O_683,N_47513,N_49248);
or UO_684 (O_684,N_48895,N_49188);
nor UO_685 (O_685,N_48322,N_47744);
nor UO_686 (O_686,N_49496,N_48045);
or UO_687 (O_687,N_48928,N_47871);
xnor UO_688 (O_688,N_48738,N_49453);
or UO_689 (O_689,N_49531,N_48081);
nand UO_690 (O_690,N_47603,N_48257);
xnor UO_691 (O_691,N_47626,N_48219);
xnor UO_692 (O_692,N_49563,N_48352);
nor UO_693 (O_693,N_47746,N_48407);
and UO_694 (O_694,N_49763,N_48616);
nor UO_695 (O_695,N_48253,N_48583);
nand UO_696 (O_696,N_47654,N_49128);
xor UO_697 (O_697,N_49051,N_47683);
or UO_698 (O_698,N_49873,N_48782);
or UO_699 (O_699,N_49899,N_49658);
nand UO_700 (O_700,N_48987,N_49318);
xnor UO_701 (O_701,N_48050,N_48964);
or UO_702 (O_702,N_49111,N_49693);
or UO_703 (O_703,N_49055,N_48610);
xnor UO_704 (O_704,N_49328,N_49079);
xor UO_705 (O_705,N_48506,N_47679);
and UO_706 (O_706,N_49725,N_49167);
nand UO_707 (O_707,N_49093,N_49258);
nand UO_708 (O_708,N_49306,N_48988);
and UO_709 (O_709,N_49536,N_49947);
or UO_710 (O_710,N_48804,N_49303);
nand UO_711 (O_711,N_48604,N_47539);
nand UO_712 (O_712,N_49053,N_47784);
and UO_713 (O_713,N_49946,N_49241);
or UO_714 (O_714,N_48715,N_48388);
and UO_715 (O_715,N_47763,N_49154);
nor UO_716 (O_716,N_47732,N_47807);
nand UO_717 (O_717,N_47934,N_48640);
or UO_718 (O_718,N_48806,N_49301);
xor UO_719 (O_719,N_49028,N_48075);
nand UO_720 (O_720,N_47805,N_48538);
and UO_721 (O_721,N_49903,N_47839);
or UO_722 (O_722,N_48525,N_48012);
nor UO_723 (O_723,N_47656,N_48896);
xnor UO_724 (O_724,N_49295,N_48837);
nand UO_725 (O_725,N_48158,N_49122);
and UO_726 (O_726,N_48961,N_49450);
nor UO_727 (O_727,N_48232,N_49655);
xnor UO_728 (O_728,N_47661,N_49867);
nand UO_729 (O_729,N_47785,N_49816);
xor UO_730 (O_730,N_49380,N_47549);
and UO_731 (O_731,N_48193,N_49073);
or UO_732 (O_732,N_49080,N_47940);
nand UO_733 (O_733,N_48780,N_48079);
or UO_734 (O_734,N_48343,N_49208);
nand UO_735 (O_735,N_47999,N_49746);
nand UO_736 (O_736,N_49980,N_49766);
xnor UO_737 (O_737,N_48285,N_48086);
xor UO_738 (O_738,N_48856,N_47757);
nor UO_739 (O_739,N_47892,N_48262);
xor UO_740 (O_740,N_49131,N_48043);
and UO_741 (O_741,N_49933,N_49509);
xnor UO_742 (O_742,N_48588,N_49555);
xor UO_743 (O_743,N_49745,N_49627);
or UO_744 (O_744,N_49047,N_49108);
or UO_745 (O_745,N_48472,N_49896);
xnor UO_746 (O_746,N_48201,N_48188);
nand UO_747 (O_747,N_48303,N_48108);
and UO_748 (O_748,N_49171,N_49857);
or UO_749 (O_749,N_48514,N_48700);
xnor UO_750 (O_750,N_49657,N_47515);
or UO_751 (O_751,N_48334,N_49516);
and UO_752 (O_752,N_49327,N_48004);
nor UO_753 (O_753,N_49454,N_49465);
nand UO_754 (O_754,N_48907,N_49205);
and UO_755 (O_755,N_49776,N_49550);
or UO_756 (O_756,N_48692,N_48137);
nor UO_757 (O_757,N_48287,N_47628);
xor UO_758 (O_758,N_49285,N_47610);
and UO_759 (O_759,N_48875,N_48777);
or UO_760 (O_760,N_48152,N_48678);
or UO_761 (O_761,N_49767,N_48751);
nor UO_762 (O_762,N_49347,N_48871);
nor UO_763 (O_763,N_48001,N_48450);
and UO_764 (O_764,N_49297,N_49082);
or UO_765 (O_765,N_49387,N_49712);
nor UO_766 (O_766,N_49921,N_48612);
nor UO_767 (O_767,N_48644,N_49375);
nor UO_768 (O_768,N_48499,N_47627);
nand UO_769 (O_769,N_47673,N_48470);
and UO_770 (O_770,N_48845,N_47675);
nand UO_771 (O_771,N_49497,N_48696);
xor UO_772 (O_772,N_49330,N_47741);
nor UO_773 (O_773,N_47825,N_48526);
and UO_774 (O_774,N_49736,N_48577);
nand UO_775 (O_775,N_49256,N_49548);
nand UO_776 (O_776,N_48315,N_48110);
and UO_777 (O_777,N_48206,N_49661);
nor UO_778 (O_778,N_49744,N_49458);
and UO_779 (O_779,N_48135,N_48443);
nor UO_780 (O_780,N_47793,N_48500);
and UO_781 (O_781,N_49118,N_48104);
and UO_782 (O_782,N_49165,N_48918);
nor UO_783 (O_783,N_48561,N_49902);
nand UO_784 (O_784,N_48691,N_49932);
nand UO_785 (O_785,N_48350,N_48815);
and UO_786 (O_786,N_47578,N_48132);
nand UO_787 (O_787,N_49936,N_48794);
xnor UO_788 (O_788,N_48735,N_49441);
nor UO_789 (O_789,N_47710,N_48134);
or UO_790 (O_790,N_48991,N_47612);
or UO_791 (O_791,N_47866,N_47507);
and UO_792 (O_792,N_47948,N_47573);
or UO_793 (O_793,N_48537,N_49155);
and UO_794 (O_794,N_48399,N_48123);
xnor UO_795 (O_795,N_48281,N_49694);
nand UO_796 (O_796,N_48797,N_49323);
nand UO_797 (O_797,N_47846,N_49930);
nand UO_798 (O_798,N_48078,N_49738);
xor UO_799 (O_799,N_48195,N_48556);
nor UO_800 (O_800,N_48323,N_49043);
nor UO_801 (O_801,N_49860,N_48701);
and UO_802 (O_802,N_47655,N_47833);
nand UO_803 (O_803,N_49265,N_49407);
or UO_804 (O_804,N_49144,N_47852);
and UO_805 (O_805,N_48730,N_48096);
xor UO_806 (O_806,N_48997,N_48211);
or UO_807 (O_807,N_49340,N_49755);
nand UO_808 (O_808,N_47765,N_49410);
xnor UO_809 (O_809,N_48849,N_49593);
nor UO_810 (O_810,N_47925,N_49934);
and UO_811 (O_811,N_47859,N_49713);
or UO_812 (O_812,N_49404,N_49284);
xor UO_813 (O_813,N_48063,N_48143);
nand UO_814 (O_814,N_48183,N_49002);
nor UO_815 (O_815,N_49007,N_49683);
nand UO_816 (O_816,N_47858,N_48395);
xor UO_817 (O_817,N_48259,N_47622);
xnor UO_818 (O_818,N_49621,N_47721);
or UO_819 (O_819,N_49777,N_49147);
or UO_820 (O_820,N_49046,N_49828);
or UO_821 (O_821,N_49547,N_48809);
or UO_822 (O_822,N_47978,N_49489);
nand UO_823 (O_823,N_49020,N_47869);
and UO_824 (O_824,N_48690,N_49157);
and UO_825 (O_825,N_49281,N_48594);
nand UO_826 (O_826,N_48338,N_48077);
nand UO_827 (O_827,N_49722,N_49223);
nor UO_828 (O_828,N_49941,N_47682);
xor UO_829 (O_829,N_49126,N_48586);
nor UO_830 (O_830,N_47848,N_49937);
or UO_831 (O_831,N_49447,N_48546);
xor UO_832 (O_832,N_48467,N_47571);
or UO_833 (O_833,N_48362,N_49184);
nor UO_834 (O_834,N_48022,N_48420);
or UO_835 (O_835,N_48884,N_48058);
and UO_836 (O_836,N_49571,N_47924);
or UO_837 (O_837,N_49685,N_49302);
and UO_838 (O_838,N_49152,N_48162);
nand UO_839 (O_839,N_48356,N_48220);
xnor UO_840 (O_840,N_49106,N_48451);
nor UO_841 (O_841,N_48371,N_48222);
and UO_842 (O_842,N_49145,N_48563);
nor UO_843 (O_843,N_48491,N_48216);
or UO_844 (O_844,N_48440,N_49310);
or UO_845 (O_845,N_49665,N_48805);
nand UO_846 (O_846,N_48003,N_49001);
xnor UO_847 (O_847,N_49870,N_48054);
nor UO_848 (O_848,N_48181,N_48517);
xnor UO_849 (O_849,N_49822,N_49187);
nand UO_850 (O_850,N_47544,N_48791);
and UO_851 (O_851,N_49939,N_47625);
nand UO_852 (O_852,N_47766,N_49814);
and UO_853 (O_853,N_49086,N_49245);
and UO_854 (O_854,N_47767,N_49662);
and UO_855 (O_855,N_48480,N_49607);
xor UO_856 (O_856,N_49348,N_47580);
or UO_857 (O_857,N_49481,N_49252);
xnor UO_858 (O_858,N_48469,N_49362);
nand UO_859 (O_859,N_48205,N_48304);
and UO_860 (O_860,N_49739,N_47760);
and UO_861 (O_861,N_48933,N_49156);
nand UO_862 (O_862,N_49376,N_49240);
nand UO_863 (O_863,N_49732,N_49360);
and UO_864 (O_864,N_49081,N_49604);
xnor UO_865 (O_865,N_48401,N_49452);
xor UO_866 (O_866,N_48418,N_48564);
and UO_867 (O_867,N_49293,N_48008);
or UO_868 (O_868,N_48128,N_47874);
and UO_869 (O_869,N_47962,N_49674);
xnor UO_870 (O_870,N_49861,N_49740);
nand UO_871 (O_871,N_48292,N_47855);
nor UO_872 (O_872,N_48880,N_48466);
nand UO_873 (O_873,N_48704,N_49412);
nand UO_874 (O_874,N_47877,N_49578);
xor UO_875 (O_875,N_47864,N_48642);
or UO_876 (O_876,N_49244,N_49421);
nor UO_877 (O_877,N_49180,N_48963);
xnor UO_878 (O_878,N_48330,N_47635);
nand UO_879 (O_879,N_48182,N_48187);
nor UO_880 (O_880,N_49161,N_49688);
nand UO_881 (O_881,N_47779,N_48835);
nor UO_882 (O_882,N_49499,N_49063);
nor UO_883 (O_883,N_49512,N_48207);
and UO_884 (O_884,N_49049,N_49507);
nor UO_885 (O_885,N_47771,N_48948);
xor UO_886 (O_886,N_48433,N_48785);
and UO_887 (O_887,N_47696,N_48753);
nand UO_888 (O_888,N_49642,N_49024);
nor UO_889 (O_889,N_48754,N_47946);
nand UO_890 (O_890,N_47811,N_47529);
nand UO_891 (O_891,N_48955,N_49312);
nor UO_892 (O_892,N_48332,N_49666);
nor UO_893 (O_893,N_48367,N_48930);
xor UO_894 (O_894,N_49520,N_49515);
nor UO_895 (O_895,N_49646,N_49503);
and UO_896 (O_896,N_48714,N_47778);
nand UO_897 (O_897,N_48765,N_47687);
nand UO_898 (O_898,N_47662,N_48218);
nor UO_899 (O_899,N_48685,N_48677);
nor UO_900 (O_900,N_47526,N_48147);
and UO_901 (O_901,N_49757,N_49045);
nor UO_902 (O_902,N_48410,N_49419);
nand UO_903 (O_903,N_48971,N_48298);
or UO_904 (O_904,N_48241,N_47831);
nor UO_905 (O_905,N_47641,N_48972);
xor UO_906 (O_906,N_49493,N_49586);
xor UO_907 (O_907,N_49559,N_48023);
nand UO_908 (O_908,N_48483,N_49862);
xnor UO_909 (O_909,N_47650,N_48861);
nor UO_910 (O_910,N_49277,N_49718);
nor UO_911 (O_911,N_49914,N_49664);
nor UO_912 (O_912,N_49098,N_49210);
nand UO_913 (O_913,N_49456,N_48071);
nor UO_914 (O_914,N_49263,N_48729);
xor UO_915 (O_915,N_49849,N_48822);
nand UO_916 (O_916,N_48628,N_49836);
and UO_917 (O_917,N_48154,N_49133);
or UO_918 (O_918,N_48859,N_49486);
nand UO_919 (O_919,N_48006,N_49760);
and UO_920 (O_920,N_48215,N_48919);
nor UO_921 (O_921,N_48311,N_49355);
or UO_922 (O_922,N_47898,N_48832);
and UO_923 (O_923,N_48783,N_49833);
nand UO_924 (O_924,N_49342,N_49800);
nor UO_925 (O_925,N_48996,N_49605);
xor UO_926 (O_926,N_47896,N_48042);
and UO_927 (O_927,N_49041,N_49123);
nor UO_928 (O_928,N_49069,N_47918);
and UO_929 (O_929,N_48164,N_49383);
nor UO_930 (O_930,N_48510,N_49377);
nand UO_931 (O_931,N_48151,N_49488);
or UO_932 (O_932,N_47541,N_49236);
xor UO_933 (O_933,N_48120,N_48995);
xor UO_934 (O_934,N_48226,N_47758);
xor UO_935 (O_935,N_48670,N_47520);
or UO_936 (O_936,N_48256,N_47536);
xor UO_937 (O_937,N_48934,N_47569);
xor UO_938 (O_938,N_48926,N_47602);
nand UO_939 (O_939,N_49077,N_49309);
and UO_940 (O_940,N_49821,N_48080);
xor UO_941 (O_941,N_49409,N_48346);
nand UO_942 (O_942,N_48403,N_48596);
or UO_943 (O_943,N_47637,N_48912);
or UO_944 (O_944,N_47590,N_47681);
or UO_945 (O_945,N_49291,N_48379);
nand UO_946 (O_946,N_47623,N_49584);
xnor UO_947 (O_947,N_47772,N_49243);
nand UO_948 (O_948,N_49426,N_48925);
xnor UO_949 (O_949,N_48827,N_47707);
and UO_950 (O_950,N_49389,N_48773);
nor UO_951 (O_951,N_49951,N_49868);
nor UO_952 (O_952,N_49590,N_47750);
nand UO_953 (O_953,N_49761,N_48931);
nor UO_954 (O_954,N_47633,N_48034);
nor UO_955 (O_955,N_49278,N_48840);
nor UO_956 (O_956,N_49475,N_49576);
nand UO_957 (O_957,N_48428,N_48282);
or UO_958 (O_958,N_49173,N_47922);
xnor UO_959 (O_959,N_47801,N_48196);
nor UO_960 (O_960,N_48289,N_48307);
and UO_961 (O_961,N_49514,N_49523);
and UO_962 (O_962,N_48650,N_49466);
xor UO_963 (O_963,N_48843,N_47734);
nand UO_964 (O_964,N_49283,N_49457);
and UO_965 (O_965,N_49470,N_47882);
nor UO_966 (O_966,N_49742,N_48747);
nor UO_967 (O_967,N_48277,N_47857);
and UO_968 (O_968,N_47937,N_48788);
nor UO_969 (O_969,N_49622,N_49966);
nand UO_970 (O_970,N_49250,N_49314);
or UO_971 (O_971,N_49992,N_48046);
nor UO_972 (O_972,N_47991,N_47879);
or UO_973 (O_973,N_47604,N_48074);
and UO_974 (O_974,N_49322,N_48681);
and UO_975 (O_975,N_49382,N_49193);
or UO_976 (O_976,N_47701,N_48069);
or UO_977 (O_977,N_48607,N_49151);
nand UO_978 (O_978,N_49670,N_48274);
or UO_979 (O_979,N_47865,N_49146);
nand UO_980 (O_980,N_49255,N_48661);
and UO_981 (O_981,N_48529,N_49900);
xnor UO_982 (O_982,N_49678,N_47666);
or UO_983 (O_983,N_48841,N_49970);
nand UO_984 (O_984,N_48047,N_48676);
nor UO_985 (O_985,N_49954,N_49251);
or UO_986 (O_986,N_49476,N_48202);
and UO_987 (O_987,N_47935,N_48452);
and UO_988 (O_988,N_49910,N_48703);
xor UO_989 (O_989,N_47914,N_47915);
nand UO_990 (O_990,N_48107,N_48655);
xnor UO_991 (O_991,N_48363,N_49917);
nand UO_992 (O_992,N_48229,N_49659);
nor UO_993 (O_993,N_48319,N_48393);
xnor UO_994 (O_994,N_49647,N_49986);
xor UO_995 (O_995,N_49257,N_48886);
nand UO_996 (O_996,N_49416,N_49032);
and UO_997 (O_997,N_48587,N_47596);
nand UO_998 (O_998,N_49955,N_48532);
nand UO_999 (O_999,N_49993,N_49141);
or UO_1000 (O_1000,N_49723,N_47714);
nand UO_1001 (O_1001,N_47642,N_49316);
or UO_1002 (O_1002,N_49469,N_48434);
nor UO_1003 (O_1003,N_48762,N_49090);
or UO_1004 (O_1004,N_49889,N_49686);
nand UO_1005 (O_1005,N_48868,N_49915);
nand UO_1006 (O_1006,N_48877,N_49013);
nor UO_1007 (O_1007,N_48103,N_47723);
and UO_1008 (O_1008,N_48121,N_49498);
nor UO_1009 (O_1009,N_47826,N_48064);
or UO_1010 (O_1010,N_48133,N_49715);
xnor UO_1011 (O_1011,N_47951,N_49463);
nand UO_1012 (O_1012,N_48238,N_49083);
nand UO_1013 (O_1013,N_48712,N_48504);
nor UO_1014 (O_1014,N_47509,N_48748);
nand UO_1015 (O_1015,N_49819,N_48031);
nand UO_1016 (O_1016,N_47609,N_49378);
or UO_1017 (O_1017,N_49791,N_48813);
nor UO_1018 (O_1018,N_47984,N_48260);
or UO_1019 (O_1019,N_48175,N_48891);
xnor UO_1020 (O_1020,N_47591,N_49521);
nor UO_1021 (O_1021,N_48796,N_47646);
xor UO_1022 (O_1022,N_49315,N_47966);
xor UO_1023 (O_1023,N_48766,N_48041);
xnor UO_1024 (O_1024,N_47670,N_48127);
nor UO_1025 (O_1025,N_48763,N_49317);
and UO_1026 (O_1026,N_49977,N_49679);
nand UO_1027 (O_1027,N_48129,N_48273);
nor UO_1028 (O_1028,N_47754,N_49948);
nor UO_1029 (O_1029,N_48639,N_47531);
and UO_1030 (O_1030,N_49573,N_48177);
nand UO_1031 (O_1031,N_47818,N_49371);
or UO_1032 (O_1032,N_48686,N_48179);
and UO_1033 (O_1033,N_48342,N_48825);
or UO_1034 (O_1034,N_47938,N_48946);
or UO_1035 (O_1035,N_48505,N_49337);
nor UO_1036 (O_1036,N_48464,N_49913);
nor UO_1037 (O_1037,N_47773,N_49888);
nand UO_1038 (O_1038,N_47985,N_49212);
nor UO_1039 (O_1039,N_47949,N_48375);
xnor UO_1040 (O_1040,N_48569,N_49653);
or UO_1041 (O_1041,N_47546,N_49324);
nor UO_1042 (O_1042,N_48516,N_48869);
or UO_1043 (O_1043,N_47814,N_48351);
nor UO_1044 (O_1044,N_47783,N_48366);
nor UO_1045 (O_1045,N_48145,N_47792);
nand UO_1046 (O_1046,N_47528,N_47958);
or UO_1047 (O_1047,N_48684,N_48146);
nand UO_1048 (O_1048,N_48820,N_48709);
nor UO_1049 (O_1049,N_49927,N_49820);
and UO_1050 (O_1050,N_48474,N_48722);
nand UO_1051 (O_1051,N_48049,N_48853);
nor UO_1052 (O_1052,N_48792,N_49189);
xnor UO_1053 (O_1053,N_48539,N_48251);
or UO_1054 (O_1054,N_47921,N_49149);
and UO_1055 (O_1055,N_49806,N_48970);
and UO_1056 (O_1056,N_49785,N_49026);
or UO_1057 (O_1057,N_48409,N_48484);
xor UO_1058 (O_1058,N_48172,N_49071);
nor UO_1059 (O_1059,N_47812,N_48994);
nand UO_1060 (O_1060,N_49675,N_49254);
xnor UO_1061 (O_1061,N_49423,N_49319);
xor UO_1062 (O_1062,N_49462,N_49931);
or UO_1063 (O_1063,N_48167,N_47695);
or UO_1064 (O_1064,N_49854,N_49372);
nand UO_1065 (O_1065,N_48888,N_49215);
or UO_1066 (O_1066,N_49396,N_48087);
and UO_1067 (O_1067,N_47630,N_48153);
or UO_1068 (O_1068,N_48402,N_49035);
xor UO_1069 (O_1069,N_49418,N_49460);
nand UO_1070 (O_1070,N_47908,N_48555);
nand UO_1071 (O_1071,N_48608,N_48717);
and UO_1072 (O_1072,N_49623,N_48199);
nand UO_1073 (O_1073,N_49928,N_49786);
and UO_1074 (O_1074,N_49438,N_49329);
nor UO_1075 (O_1075,N_48932,N_47538);
xor UO_1076 (O_1076,N_48002,N_47830);
or UO_1077 (O_1077,N_48381,N_48358);
and UO_1078 (O_1078,N_48308,N_49706);
xor UO_1079 (O_1079,N_48923,N_47619);
nor UO_1080 (O_1080,N_49338,N_48408);
nand UO_1081 (O_1081,N_49178,N_48618);
xor UO_1082 (O_1082,N_48102,N_49430);
nor UO_1083 (O_1083,N_47895,N_47843);
xor UO_1084 (O_1084,N_49826,N_48453);
or UO_1085 (O_1085,N_49667,N_49139);
xor UO_1086 (O_1086,N_48157,N_47798);
nor UO_1087 (O_1087,N_48423,N_48973);
nor UO_1088 (O_1088,N_47657,N_49894);
and UO_1089 (O_1089,N_49000,N_49227);
xnor UO_1090 (O_1090,N_48068,N_48770);
nor UO_1091 (O_1091,N_49427,N_48297);
and UO_1092 (O_1092,N_49264,N_48899);
and UO_1093 (O_1093,N_48554,N_48945);
nand UO_1094 (O_1094,N_48567,N_49709);
and UO_1095 (O_1095,N_49175,N_48967);
nor UO_1096 (O_1096,N_49729,N_49897);
and UO_1097 (O_1097,N_49068,N_47850);
xnor UO_1098 (O_1098,N_49392,N_49844);
nor UO_1099 (O_1099,N_47724,N_49841);
xnor UO_1100 (O_1100,N_48497,N_49735);
nor UO_1101 (O_1101,N_48015,N_47726);
xor UO_1102 (O_1102,N_49085,N_48885);
xor UO_1103 (O_1103,N_49103,N_47944);
or UO_1104 (O_1104,N_49698,N_48836);
or UO_1105 (O_1105,N_48718,N_49084);
or UO_1106 (O_1106,N_49501,N_48494);
nor UO_1107 (O_1107,N_48787,N_49349);
xor UO_1108 (O_1108,N_48341,N_48170);
nor UO_1109 (O_1109,N_47781,N_49386);
nand UO_1110 (O_1110,N_49219,N_48457);
nand UO_1111 (O_1111,N_49618,N_47585);
nor UO_1112 (O_1112,N_47867,N_48302);
xnor UO_1113 (O_1113,N_49172,N_47947);
xnor UO_1114 (O_1114,N_47861,N_48384);
nand UO_1115 (O_1115,N_49796,N_48057);
or UO_1116 (O_1116,N_48999,N_48246);
nand UO_1117 (O_1117,N_49609,N_49691);
xor UO_1118 (O_1118,N_49023,N_49859);
and UO_1119 (O_1119,N_49199,N_47775);
or UO_1120 (O_1120,N_49271,N_49771);
and UO_1121 (O_1121,N_48138,N_47817);
xnor UO_1122 (O_1122,N_49866,N_49204);
nand UO_1123 (O_1123,N_49907,N_49575);
nand UO_1124 (O_1124,N_49990,N_47764);
nor UO_1125 (O_1125,N_49221,N_49211);
and UO_1126 (O_1126,N_49648,N_49112);
xor UO_1127 (O_1127,N_49113,N_48688);
xor UO_1128 (O_1128,N_48502,N_49060);
nand UO_1129 (O_1129,N_49519,N_47511);
or UO_1130 (O_1130,N_48364,N_49390);
nor UO_1131 (O_1131,N_48112,N_48496);
nand UO_1132 (O_1132,N_48850,N_47632);
or UO_1133 (O_1133,N_49326,N_49505);
or UO_1134 (O_1134,N_49803,N_49334);
and UO_1135 (O_1135,N_47560,N_47837);
and UO_1136 (O_1136,N_49704,N_48689);
xor UO_1137 (O_1137,N_49950,N_47606);
nor UO_1138 (O_1138,N_49261,N_48993);
nor UO_1139 (O_1139,N_48233,N_49099);
and UO_1140 (O_1140,N_49626,N_47579);
nor UO_1141 (O_1141,N_47860,N_49062);
nor UO_1142 (O_1142,N_47849,N_48272);
or UO_1143 (O_1143,N_48200,N_49105);
nor UO_1144 (O_1144,N_48168,N_47658);
xnor UO_1145 (O_1145,N_49399,N_48606);
or UO_1146 (O_1146,N_49042,N_48633);
nand UO_1147 (O_1147,N_49620,N_48169);
nand UO_1148 (O_1148,N_48774,N_48267);
nand UO_1149 (O_1149,N_47957,N_49637);
xnor UO_1150 (O_1150,N_49545,N_48394);
nor UO_1151 (O_1151,N_48985,N_48523);
xor UO_1152 (O_1152,N_48582,N_47996);
and UO_1153 (O_1153,N_48734,N_49374);
nor UO_1154 (O_1154,N_48488,N_47955);
xnor UO_1155 (O_1155,N_47652,N_48653);
xnor UO_1156 (O_1156,N_48095,N_49792);
xor UO_1157 (O_1157,N_48159,N_49367);
or UO_1158 (O_1158,N_49097,N_49504);
nor UO_1159 (O_1159,N_49116,N_48093);
xor UO_1160 (O_1160,N_49420,N_48603);
nand UO_1161 (O_1161,N_49078,N_47597);
nand UO_1162 (O_1162,N_49482,N_48340);
or UO_1163 (O_1163,N_48854,N_49434);
xnor UO_1164 (O_1164,N_49351,N_48336);
or UO_1165 (O_1165,N_48518,N_49751);
nor UO_1166 (O_1166,N_48247,N_48000);
or UO_1167 (O_1167,N_49366,N_48507);
xnor UO_1168 (O_1168,N_47731,N_49668);
nor UO_1169 (O_1169,N_49332,N_47887);
and UO_1170 (O_1170,N_49320,N_48250);
or UO_1171 (O_1171,N_47844,N_49182);
and UO_1172 (O_1172,N_49017,N_48935);
nand UO_1173 (O_1173,N_49480,N_49292);
xor UO_1174 (O_1174,N_48487,N_48535);
nand UO_1175 (O_1175,N_47828,N_49567);
nand UO_1176 (O_1176,N_49588,N_48619);
or UO_1177 (O_1177,N_49595,N_49962);
nor UO_1178 (O_1178,N_47748,N_48874);
nor UO_1179 (O_1179,N_47725,N_49294);
xor UO_1180 (O_1180,N_49580,N_49075);
xnor UO_1181 (O_1181,N_47532,N_48547);
nand UO_1182 (O_1182,N_49687,N_48486);
nand UO_1183 (O_1183,N_48801,N_48293);
or UO_1184 (O_1184,N_49842,N_47577);
and UO_1185 (O_1185,N_48383,N_49602);
nand UO_1186 (O_1186,N_48239,N_48038);
nand UO_1187 (O_1187,N_48981,N_49474);
nand UO_1188 (O_1188,N_49202,N_47912);
xor UO_1189 (O_1189,N_47762,N_48387);
xor UO_1190 (O_1190,N_49823,N_49846);
nand UO_1191 (O_1191,N_48950,N_48846);
xnor UO_1192 (O_1192,N_49549,N_49346);
nand UO_1193 (O_1193,N_49095,N_48258);
or UO_1194 (O_1194,N_48795,N_47919);
or UO_1195 (O_1195,N_49759,N_47747);
and UO_1196 (O_1196,N_48144,N_49485);
and UO_1197 (O_1197,N_47975,N_48374);
nor UO_1198 (O_1198,N_48221,N_47776);
nand UO_1199 (O_1199,N_48527,N_49091);
or UO_1200 (O_1200,N_47740,N_49344);
and UO_1201 (O_1201,N_48631,N_47967);
xor UO_1202 (O_1202,N_48415,N_47524);
or UO_1203 (O_1203,N_48288,N_49541);
or UO_1204 (O_1204,N_49728,N_49290);
nor UO_1205 (O_1205,N_48865,N_48376);
xor UO_1206 (O_1206,N_48155,N_49143);
nand UO_1207 (O_1207,N_47974,N_48039);
xnor UO_1208 (O_1208,N_47595,N_48264);
nor UO_1209 (O_1209,N_48768,N_48286);
nor UO_1210 (O_1210,N_49517,N_48598);
or UO_1211 (O_1211,N_48980,N_48173);
xor UO_1212 (O_1212,N_49600,N_47550);
or UO_1213 (O_1213,N_47995,N_48291);
or UO_1214 (O_1214,N_48562,N_49494);
nand UO_1215 (O_1215,N_47986,N_49087);
xnor UO_1216 (O_1216,N_49089,N_48839);
xor UO_1217 (O_1217,N_47980,N_48819);
nor UO_1218 (O_1218,N_48706,N_49554);
and UO_1219 (O_1219,N_49635,N_48380);
and UO_1220 (O_1220,N_48662,N_47768);
nor UO_1221 (O_1221,N_49645,N_48914);
or UO_1222 (O_1222,N_48382,N_49449);
xor UO_1223 (O_1223,N_47533,N_48131);
xnor UO_1224 (O_1224,N_49229,N_48254);
xor UO_1225 (O_1225,N_49529,N_47992);
or UO_1226 (O_1226,N_49033,N_49039);
and UO_1227 (O_1227,N_48124,N_48300);
xnor UO_1228 (O_1228,N_47535,N_48887);
nor UO_1229 (O_1229,N_48372,N_49809);
and UO_1230 (O_1230,N_48191,N_47899);
nor UO_1231 (O_1231,N_47845,N_48033);
or UO_1232 (O_1232,N_48641,N_49181);
nor UO_1233 (O_1233,N_49546,N_49153);
and UO_1234 (O_1234,N_49971,N_49036);
xor UO_1235 (O_1235,N_49582,N_47584);
xor UO_1236 (O_1236,N_48936,N_48723);
and UO_1237 (O_1237,N_48975,N_47565);
and UO_1238 (O_1238,N_49916,N_48230);
or UO_1239 (O_1239,N_48320,N_48659);
nand UO_1240 (O_1240,N_48513,N_47920);
xor UO_1241 (O_1241,N_49391,N_48028);
xnor UO_1242 (O_1242,N_49940,N_48816);
xnor UO_1243 (O_1243,N_48240,N_48542);
xnor UO_1244 (O_1244,N_48389,N_49395);
nand UO_1245 (O_1245,N_48982,N_49094);
or UO_1246 (O_1246,N_48261,N_47720);
nor UO_1247 (O_1247,N_47854,N_49756);
and UO_1248 (O_1248,N_48915,N_49865);
and UO_1249 (O_1249,N_49511,N_47730);
or UO_1250 (O_1250,N_48191,N_49996);
or UO_1251 (O_1251,N_47546,N_48109);
xnor UO_1252 (O_1252,N_48338,N_48622);
nor UO_1253 (O_1253,N_48573,N_48973);
or UO_1254 (O_1254,N_48007,N_49486);
nor UO_1255 (O_1255,N_48324,N_47605);
or UO_1256 (O_1256,N_48432,N_48267);
xnor UO_1257 (O_1257,N_48915,N_48405);
and UO_1258 (O_1258,N_49096,N_47686);
nand UO_1259 (O_1259,N_49495,N_48886);
nor UO_1260 (O_1260,N_48352,N_49558);
and UO_1261 (O_1261,N_48650,N_49667);
nor UO_1262 (O_1262,N_49620,N_48234);
xnor UO_1263 (O_1263,N_49683,N_49345);
and UO_1264 (O_1264,N_47637,N_48183);
nor UO_1265 (O_1265,N_48125,N_49791);
nand UO_1266 (O_1266,N_48733,N_48045);
and UO_1267 (O_1267,N_47822,N_49751);
nor UO_1268 (O_1268,N_47880,N_48927);
nor UO_1269 (O_1269,N_48242,N_49448);
nor UO_1270 (O_1270,N_49916,N_49374);
or UO_1271 (O_1271,N_48321,N_49170);
xnor UO_1272 (O_1272,N_47973,N_49599);
and UO_1273 (O_1273,N_48628,N_48581);
nand UO_1274 (O_1274,N_48846,N_47816);
xor UO_1275 (O_1275,N_49990,N_49078);
nor UO_1276 (O_1276,N_48297,N_49417);
nor UO_1277 (O_1277,N_48029,N_48244);
or UO_1278 (O_1278,N_47632,N_48570);
nor UO_1279 (O_1279,N_49629,N_48594);
or UO_1280 (O_1280,N_48296,N_49982);
nor UO_1281 (O_1281,N_49834,N_47863);
and UO_1282 (O_1282,N_48578,N_49203);
and UO_1283 (O_1283,N_49342,N_47641);
xor UO_1284 (O_1284,N_48461,N_48895);
xnor UO_1285 (O_1285,N_49211,N_49419);
or UO_1286 (O_1286,N_49158,N_49884);
nand UO_1287 (O_1287,N_48238,N_48472);
and UO_1288 (O_1288,N_48752,N_48916);
xor UO_1289 (O_1289,N_48872,N_48236);
nor UO_1290 (O_1290,N_49328,N_47548);
nor UO_1291 (O_1291,N_48865,N_49492);
nand UO_1292 (O_1292,N_47501,N_47840);
xnor UO_1293 (O_1293,N_48677,N_48360);
and UO_1294 (O_1294,N_48665,N_49446);
or UO_1295 (O_1295,N_48751,N_47912);
or UO_1296 (O_1296,N_48568,N_48538);
or UO_1297 (O_1297,N_48949,N_49346);
xor UO_1298 (O_1298,N_49505,N_49354);
and UO_1299 (O_1299,N_49486,N_49918);
nor UO_1300 (O_1300,N_49698,N_48150);
nand UO_1301 (O_1301,N_47761,N_48814);
and UO_1302 (O_1302,N_49930,N_48953);
or UO_1303 (O_1303,N_49272,N_48601);
nand UO_1304 (O_1304,N_47769,N_47656);
and UO_1305 (O_1305,N_48892,N_49363);
nand UO_1306 (O_1306,N_49170,N_48861);
or UO_1307 (O_1307,N_49826,N_48313);
xnor UO_1308 (O_1308,N_48913,N_49797);
or UO_1309 (O_1309,N_48835,N_48364);
nor UO_1310 (O_1310,N_48241,N_48426);
or UO_1311 (O_1311,N_47586,N_47571);
nand UO_1312 (O_1312,N_47530,N_49867);
or UO_1313 (O_1313,N_47690,N_48307);
and UO_1314 (O_1314,N_49558,N_48365);
and UO_1315 (O_1315,N_47605,N_47592);
and UO_1316 (O_1316,N_48908,N_48415);
nor UO_1317 (O_1317,N_47943,N_48987);
nand UO_1318 (O_1318,N_48016,N_48420);
or UO_1319 (O_1319,N_49089,N_47712);
and UO_1320 (O_1320,N_49043,N_48663);
nor UO_1321 (O_1321,N_47726,N_49491);
and UO_1322 (O_1322,N_49333,N_49313);
or UO_1323 (O_1323,N_49390,N_48560);
or UO_1324 (O_1324,N_48935,N_47936);
nor UO_1325 (O_1325,N_47951,N_48794);
nor UO_1326 (O_1326,N_47853,N_48928);
or UO_1327 (O_1327,N_49235,N_47955);
nor UO_1328 (O_1328,N_49861,N_48195);
nor UO_1329 (O_1329,N_48408,N_48756);
xor UO_1330 (O_1330,N_47885,N_49029);
xnor UO_1331 (O_1331,N_49590,N_48452);
or UO_1332 (O_1332,N_48415,N_49738);
nand UO_1333 (O_1333,N_47582,N_49290);
and UO_1334 (O_1334,N_49664,N_48447);
or UO_1335 (O_1335,N_48322,N_48282);
and UO_1336 (O_1336,N_48044,N_49375);
nor UO_1337 (O_1337,N_48834,N_48294);
and UO_1338 (O_1338,N_47814,N_48827);
and UO_1339 (O_1339,N_49237,N_48569);
and UO_1340 (O_1340,N_48635,N_47645);
nand UO_1341 (O_1341,N_48221,N_48825);
or UO_1342 (O_1342,N_48424,N_48561);
and UO_1343 (O_1343,N_48907,N_48879);
xnor UO_1344 (O_1344,N_48455,N_49066);
nand UO_1345 (O_1345,N_47667,N_48069);
nand UO_1346 (O_1346,N_47799,N_49669);
nand UO_1347 (O_1347,N_48851,N_48779);
nor UO_1348 (O_1348,N_48466,N_48915);
nor UO_1349 (O_1349,N_49389,N_48023);
or UO_1350 (O_1350,N_48484,N_49527);
nor UO_1351 (O_1351,N_48311,N_47503);
nor UO_1352 (O_1352,N_48800,N_47980);
and UO_1353 (O_1353,N_49934,N_47713);
and UO_1354 (O_1354,N_49962,N_49978);
nand UO_1355 (O_1355,N_49823,N_48078);
nand UO_1356 (O_1356,N_48406,N_48151);
nand UO_1357 (O_1357,N_48819,N_48781);
and UO_1358 (O_1358,N_47922,N_49726);
and UO_1359 (O_1359,N_49561,N_48919);
or UO_1360 (O_1360,N_49958,N_49679);
or UO_1361 (O_1361,N_47770,N_49060);
xnor UO_1362 (O_1362,N_47800,N_49498);
and UO_1363 (O_1363,N_48316,N_47592);
nor UO_1364 (O_1364,N_49608,N_48013);
and UO_1365 (O_1365,N_49636,N_47815);
and UO_1366 (O_1366,N_47966,N_49435);
or UO_1367 (O_1367,N_48243,N_49749);
and UO_1368 (O_1368,N_48096,N_48590);
nand UO_1369 (O_1369,N_47523,N_49288);
nand UO_1370 (O_1370,N_47766,N_49327);
and UO_1371 (O_1371,N_47892,N_48849);
nand UO_1372 (O_1372,N_48978,N_48626);
or UO_1373 (O_1373,N_48828,N_49095);
xor UO_1374 (O_1374,N_49769,N_49427);
or UO_1375 (O_1375,N_48747,N_47919);
or UO_1376 (O_1376,N_49360,N_49112);
xnor UO_1377 (O_1377,N_47955,N_48001);
nor UO_1378 (O_1378,N_48866,N_49298);
nand UO_1379 (O_1379,N_49214,N_48608);
nand UO_1380 (O_1380,N_48540,N_48462);
nand UO_1381 (O_1381,N_49405,N_48637);
xnor UO_1382 (O_1382,N_48631,N_49269);
xor UO_1383 (O_1383,N_48157,N_48501);
nor UO_1384 (O_1384,N_48665,N_49856);
and UO_1385 (O_1385,N_48403,N_49659);
and UO_1386 (O_1386,N_49418,N_49889);
or UO_1387 (O_1387,N_48363,N_48005);
nand UO_1388 (O_1388,N_48832,N_49543);
nor UO_1389 (O_1389,N_47996,N_48795);
nand UO_1390 (O_1390,N_49726,N_49904);
nand UO_1391 (O_1391,N_48292,N_49756);
nand UO_1392 (O_1392,N_48009,N_47968);
or UO_1393 (O_1393,N_48387,N_49184);
nor UO_1394 (O_1394,N_48327,N_49052);
xnor UO_1395 (O_1395,N_48141,N_49680);
and UO_1396 (O_1396,N_48698,N_49914);
xnor UO_1397 (O_1397,N_49652,N_49234);
or UO_1398 (O_1398,N_49091,N_49167);
nand UO_1399 (O_1399,N_48640,N_49907);
nand UO_1400 (O_1400,N_48856,N_48652);
xor UO_1401 (O_1401,N_49172,N_47734);
and UO_1402 (O_1402,N_47780,N_49819);
or UO_1403 (O_1403,N_49849,N_47656);
xor UO_1404 (O_1404,N_48306,N_48830);
nand UO_1405 (O_1405,N_49116,N_49018);
nor UO_1406 (O_1406,N_48580,N_48794);
and UO_1407 (O_1407,N_47567,N_49053);
nor UO_1408 (O_1408,N_48084,N_48871);
and UO_1409 (O_1409,N_48912,N_49567);
and UO_1410 (O_1410,N_48981,N_49458);
xor UO_1411 (O_1411,N_49946,N_49981);
or UO_1412 (O_1412,N_48720,N_48143);
or UO_1413 (O_1413,N_49208,N_48668);
xnor UO_1414 (O_1414,N_49404,N_48074);
and UO_1415 (O_1415,N_49223,N_49167);
or UO_1416 (O_1416,N_47576,N_49441);
xnor UO_1417 (O_1417,N_48662,N_47651);
xor UO_1418 (O_1418,N_47509,N_49270);
nor UO_1419 (O_1419,N_48263,N_47547);
xnor UO_1420 (O_1420,N_49843,N_48049);
and UO_1421 (O_1421,N_48058,N_49642);
or UO_1422 (O_1422,N_49949,N_47889);
xor UO_1423 (O_1423,N_48758,N_48972);
nand UO_1424 (O_1424,N_48648,N_47870);
and UO_1425 (O_1425,N_49391,N_49069);
or UO_1426 (O_1426,N_48246,N_48770);
nor UO_1427 (O_1427,N_47503,N_49340);
nor UO_1428 (O_1428,N_49313,N_47652);
xor UO_1429 (O_1429,N_49034,N_47827);
or UO_1430 (O_1430,N_47901,N_48924);
xor UO_1431 (O_1431,N_48392,N_48044);
and UO_1432 (O_1432,N_48801,N_49346);
or UO_1433 (O_1433,N_49611,N_48816);
and UO_1434 (O_1434,N_49491,N_49995);
or UO_1435 (O_1435,N_48714,N_49813);
xnor UO_1436 (O_1436,N_49573,N_49518);
nor UO_1437 (O_1437,N_47930,N_49160);
nor UO_1438 (O_1438,N_49105,N_47905);
xor UO_1439 (O_1439,N_48467,N_47631);
xor UO_1440 (O_1440,N_47527,N_48058);
xor UO_1441 (O_1441,N_47531,N_48392);
or UO_1442 (O_1442,N_49154,N_49139);
nor UO_1443 (O_1443,N_47894,N_47893);
nor UO_1444 (O_1444,N_48165,N_49953);
nand UO_1445 (O_1445,N_49689,N_48930);
xnor UO_1446 (O_1446,N_49956,N_49864);
nand UO_1447 (O_1447,N_49785,N_49207);
xnor UO_1448 (O_1448,N_49137,N_47878);
xnor UO_1449 (O_1449,N_48158,N_48803);
nor UO_1450 (O_1450,N_47520,N_48295);
nand UO_1451 (O_1451,N_49175,N_49309);
nand UO_1452 (O_1452,N_48655,N_47704);
xnor UO_1453 (O_1453,N_48558,N_47898);
or UO_1454 (O_1454,N_49838,N_47695);
nor UO_1455 (O_1455,N_48684,N_49741);
or UO_1456 (O_1456,N_48601,N_48078);
and UO_1457 (O_1457,N_49908,N_48939);
nor UO_1458 (O_1458,N_47908,N_48316);
nand UO_1459 (O_1459,N_49674,N_47563);
nor UO_1460 (O_1460,N_49294,N_49328);
nand UO_1461 (O_1461,N_49480,N_47996);
nor UO_1462 (O_1462,N_49261,N_48717);
nor UO_1463 (O_1463,N_49074,N_49082);
xor UO_1464 (O_1464,N_48145,N_49903);
xor UO_1465 (O_1465,N_47501,N_47782);
nor UO_1466 (O_1466,N_48912,N_49235);
nor UO_1467 (O_1467,N_49671,N_48450);
xnor UO_1468 (O_1468,N_47654,N_49299);
nor UO_1469 (O_1469,N_48570,N_49670);
and UO_1470 (O_1470,N_47981,N_49718);
nand UO_1471 (O_1471,N_48130,N_48410);
xor UO_1472 (O_1472,N_49168,N_49606);
xnor UO_1473 (O_1473,N_48293,N_48976);
or UO_1474 (O_1474,N_49125,N_48601);
or UO_1475 (O_1475,N_49868,N_49100);
nand UO_1476 (O_1476,N_48087,N_49637);
nand UO_1477 (O_1477,N_48016,N_47904);
and UO_1478 (O_1478,N_49600,N_47700);
and UO_1479 (O_1479,N_49062,N_47794);
and UO_1480 (O_1480,N_48258,N_48911);
nand UO_1481 (O_1481,N_47865,N_47958);
and UO_1482 (O_1482,N_48163,N_47609);
or UO_1483 (O_1483,N_47934,N_48545);
nor UO_1484 (O_1484,N_47613,N_49546);
nor UO_1485 (O_1485,N_48743,N_48036);
nand UO_1486 (O_1486,N_49393,N_49507);
xnor UO_1487 (O_1487,N_49727,N_48392);
or UO_1488 (O_1488,N_48716,N_49989);
xor UO_1489 (O_1489,N_49053,N_49802);
and UO_1490 (O_1490,N_48720,N_49130);
or UO_1491 (O_1491,N_47918,N_49028);
nand UO_1492 (O_1492,N_47994,N_48733);
or UO_1493 (O_1493,N_49388,N_49329);
nor UO_1494 (O_1494,N_49365,N_48037);
nand UO_1495 (O_1495,N_48553,N_49775);
nand UO_1496 (O_1496,N_48281,N_48569);
nand UO_1497 (O_1497,N_48068,N_49715);
or UO_1498 (O_1498,N_48621,N_49189);
and UO_1499 (O_1499,N_49108,N_48813);
xor UO_1500 (O_1500,N_48253,N_47907);
and UO_1501 (O_1501,N_49546,N_48629);
and UO_1502 (O_1502,N_49087,N_47924);
nor UO_1503 (O_1503,N_49324,N_48870);
nor UO_1504 (O_1504,N_47635,N_48392);
nand UO_1505 (O_1505,N_48969,N_47934);
nor UO_1506 (O_1506,N_48398,N_48227);
xnor UO_1507 (O_1507,N_47657,N_49989);
xor UO_1508 (O_1508,N_48829,N_49761);
or UO_1509 (O_1509,N_49043,N_49317);
or UO_1510 (O_1510,N_49543,N_48624);
or UO_1511 (O_1511,N_48720,N_48986);
nor UO_1512 (O_1512,N_48196,N_48621);
and UO_1513 (O_1513,N_48456,N_48539);
and UO_1514 (O_1514,N_47724,N_47521);
nand UO_1515 (O_1515,N_49376,N_48968);
xor UO_1516 (O_1516,N_48759,N_48981);
nand UO_1517 (O_1517,N_48177,N_49818);
and UO_1518 (O_1518,N_47831,N_47546);
and UO_1519 (O_1519,N_49255,N_49503);
nand UO_1520 (O_1520,N_49883,N_47644);
and UO_1521 (O_1521,N_49713,N_48467);
or UO_1522 (O_1522,N_49536,N_47761);
and UO_1523 (O_1523,N_49420,N_49772);
nor UO_1524 (O_1524,N_49101,N_49872);
and UO_1525 (O_1525,N_48068,N_48665);
or UO_1526 (O_1526,N_48885,N_48512);
and UO_1527 (O_1527,N_47811,N_49042);
nand UO_1528 (O_1528,N_48188,N_48265);
xor UO_1529 (O_1529,N_49147,N_48808);
nand UO_1530 (O_1530,N_48331,N_49309);
nor UO_1531 (O_1531,N_48546,N_49191);
xnor UO_1532 (O_1532,N_49973,N_47607);
xor UO_1533 (O_1533,N_49968,N_47653);
xnor UO_1534 (O_1534,N_47855,N_48695);
and UO_1535 (O_1535,N_47629,N_49953);
and UO_1536 (O_1536,N_49127,N_49655);
nor UO_1537 (O_1537,N_49405,N_48608);
or UO_1538 (O_1538,N_49392,N_49370);
nor UO_1539 (O_1539,N_49970,N_47877);
nand UO_1540 (O_1540,N_48807,N_48686);
or UO_1541 (O_1541,N_47598,N_48701);
or UO_1542 (O_1542,N_47944,N_49394);
or UO_1543 (O_1543,N_48304,N_48215);
xnor UO_1544 (O_1544,N_49769,N_48704);
and UO_1545 (O_1545,N_47791,N_49193);
nor UO_1546 (O_1546,N_48119,N_47573);
or UO_1547 (O_1547,N_48648,N_48933);
nand UO_1548 (O_1548,N_49491,N_48631);
or UO_1549 (O_1549,N_48841,N_49881);
nor UO_1550 (O_1550,N_47635,N_48017);
and UO_1551 (O_1551,N_48171,N_49696);
or UO_1552 (O_1552,N_48516,N_48925);
and UO_1553 (O_1553,N_49358,N_49697);
nand UO_1554 (O_1554,N_49875,N_49300);
nor UO_1555 (O_1555,N_47641,N_47808);
nor UO_1556 (O_1556,N_49512,N_48747);
and UO_1557 (O_1557,N_49169,N_49717);
or UO_1558 (O_1558,N_47820,N_48000);
xnor UO_1559 (O_1559,N_48675,N_47893);
and UO_1560 (O_1560,N_47939,N_48093);
or UO_1561 (O_1561,N_48028,N_48054);
or UO_1562 (O_1562,N_49490,N_47624);
and UO_1563 (O_1563,N_47936,N_47891);
xnor UO_1564 (O_1564,N_48388,N_49510);
or UO_1565 (O_1565,N_48276,N_48964);
xor UO_1566 (O_1566,N_49578,N_48539);
xor UO_1567 (O_1567,N_48176,N_49303);
or UO_1568 (O_1568,N_49359,N_48416);
and UO_1569 (O_1569,N_49175,N_49374);
or UO_1570 (O_1570,N_49901,N_48371);
nand UO_1571 (O_1571,N_48360,N_48532);
nor UO_1572 (O_1572,N_49655,N_49171);
nor UO_1573 (O_1573,N_48990,N_49049);
and UO_1574 (O_1574,N_48503,N_48112);
nand UO_1575 (O_1575,N_49980,N_48215);
xnor UO_1576 (O_1576,N_48615,N_47710);
xnor UO_1577 (O_1577,N_49226,N_49447);
or UO_1578 (O_1578,N_48323,N_49151);
and UO_1579 (O_1579,N_48196,N_48793);
or UO_1580 (O_1580,N_48716,N_48261);
and UO_1581 (O_1581,N_48800,N_48577);
or UO_1582 (O_1582,N_48491,N_47838);
nor UO_1583 (O_1583,N_49480,N_49067);
nand UO_1584 (O_1584,N_47534,N_47618);
nand UO_1585 (O_1585,N_48644,N_48429);
or UO_1586 (O_1586,N_49947,N_49822);
and UO_1587 (O_1587,N_47593,N_49176);
xnor UO_1588 (O_1588,N_49685,N_48396);
nor UO_1589 (O_1589,N_49579,N_47811);
nand UO_1590 (O_1590,N_47624,N_48858);
nand UO_1591 (O_1591,N_49217,N_49509);
and UO_1592 (O_1592,N_48348,N_48492);
nor UO_1593 (O_1593,N_49587,N_47776);
xnor UO_1594 (O_1594,N_47916,N_49565);
and UO_1595 (O_1595,N_48460,N_48505);
or UO_1596 (O_1596,N_48533,N_48767);
or UO_1597 (O_1597,N_49827,N_48357);
nand UO_1598 (O_1598,N_49297,N_49516);
and UO_1599 (O_1599,N_49710,N_49013);
xnor UO_1600 (O_1600,N_48942,N_48917);
and UO_1601 (O_1601,N_49432,N_48667);
or UO_1602 (O_1602,N_48463,N_47636);
xnor UO_1603 (O_1603,N_49224,N_47595);
xor UO_1604 (O_1604,N_49486,N_47970);
or UO_1605 (O_1605,N_49622,N_49423);
nor UO_1606 (O_1606,N_49972,N_49450);
xnor UO_1607 (O_1607,N_48792,N_47888);
nand UO_1608 (O_1608,N_47976,N_49481);
nand UO_1609 (O_1609,N_49414,N_49569);
nand UO_1610 (O_1610,N_48163,N_48251);
nand UO_1611 (O_1611,N_48141,N_48399);
nor UO_1612 (O_1612,N_48401,N_48841);
and UO_1613 (O_1613,N_48296,N_47595);
and UO_1614 (O_1614,N_49331,N_47543);
nand UO_1615 (O_1615,N_47694,N_48329);
nand UO_1616 (O_1616,N_48282,N_49688);
xor UO_1617 (O_1617,N_47506,N_49772);
xor UO_1618 (O_1618,N_48954,N_49012);
nand UO_1619 (O_1619,N_48343,N_48320);
and UO_1620 (O_1620,N_48170,N_48614);
and UO_1621 (O_1621,N_48159,N_49885);
xor UO_1622 (O_1622,N_48403,N_48994);
xor UO_1623 (O_1623,N_49635,N_48911);
and UO_1624 (O_1624,N_48351,N_47843);
or UO_1625 (O_1625,N_47769,N_49070);
or UO_1626 (O_1626,N_48225,N_49215);
and UO_1627 (O_1627,N_49223,N_47826);
xnor UO_1628 (O_1628,N_48832,N_48657);
nor UO_1629 (O_1629,N_48174,N_48205);
and UO_1630 (O_1630,N_49100,N_49555);
or UO_1631 (O_1631,N_48586,N_48092);
nand UO_1632 (O_1632,N_48851,N_49241);
xor UO_1633 (O_1633,N_49303,N_49871);
xnor UO_1634 (O_1634,N_49180,N_48983);
xor UO_1635 (O_1635,N_49105,N_48348);
and UO_1636 (O_1636,N_48477,N_49716);
nand UO_1637 (O_1637,N_48120,N_47582);
nor UO_1638 (O_1638,N_47807,N_49718);
xnor UO_1639 (O_1639,N_47696,N_47503);
nor UO_1640 (O_1640,N_49027,N_49340);
nor UO_1641 (O_1641,N_48552,N_49390);
nor UO_1642 (O_1642,N_47886,N_49711);
nor UO_1643 (O_1643,N_47904,N_49471);
xor UO_1644 (O_1644,N_48873,N_48834);
nor UO_1645 (O_1645,N_47741,N_48982);
xnor UO_1646 (O_1646,N_48427,N_47788);
xor UO_1647 (O_1647,N_49539,N_47991);
xnor UO_1648 (O_1648,N_48165,N_47590);
nand UO_1649 (O_1649,N_49847,N_48780);
nand UO_1650 (O_1650,N_49892,N_48184);
or UO_1651 (O_1651,N_49930,N_48891);
and UO_1652 (O_1652,N_49595,N_49186);
and UO_1653 (O_1653,N_48985,N_47996);
nor UO_1654 (O_1654,N_48628,N_48632);
nor UO_1655 (O_1655,N_48588,N_49796);
or UO_1656 (O_1656,N_49716,N_48155);
and UO_1657 (O_1657,N_48193,N_47748);
xor UO_1658 (O_1658,N_47832,N_47697);
xor UO_1659 (O_1659,N_48807,N_47715);
and UO_1660 (O_1660,N_47731,N_48764);
nor UO_1661 (O_1661,N_49735,N_47546);
or UO_1662 (O_1662,N_49680,N_49464);
and UO_1663 (O_1663,N_47571,N_47627);
nand UO_1664 (O_1664,N_48020,N_48660);
xnor UO_1665 (O_1665,N_49771,N_48362);
xor UO_1666 (O_1666,N_48042,N_48547);
or UO_1667 (O_1667,N_48361,N_49313);
and UO_1668 (O_1668,N_49826,N_48919);
xor UO_1669 (O_1669,N_47652,N_49132);
or UO_1670 (O_1670,N_48711,N_48510);
nor UO_1671 (O_1671,N_49685,N_49493);
nand UO_1672 (O_1672,N_49351,N_49280);
nor UO_1673 (O_1673,N_49401,N_48773);
or UO_1674 (O_1674,N_49456,N_47604);
nor UO_1675 (O_1675,N_47675,N_47505);
or UO_1676 (O_1676,N_49428,N_49870);
or UO_1677 (O_1677,N_47504,N_47638);
or UO_1678 (O_1678,N_49146,N_49125);
nor UO_1679 (O_1679,N_48224,N_47506);
xor UO_1680 (O_1680,N_48331,N_49597);
nor UO_1681 (O_1681,N_48932,N_49504);
nor UO_1682 (O_1682,N_49693,N_48445);
or UO_1683 (O_1683,N_47578,N_47554);
nor UO_1684 (O_1684,N_49826,N_48115);
and UO_1685 (O_1685,N_48004,N_48962);
or UO_1686 (O_1686,N_48483,N_48705);
and UO_1687 (O_1687,N_49172,N_47591);
and UO_1688 (O_1688,N_49786,N_49340);
xor UO_1689 (O_1689,N_48856,N_49233);
nand UO_1690 (O_1690,N_49152,N_48670);
or UO_1691 (O_1691,N_48531,N_49497);
and UO_1692 (O_1692,N_49170,N_47839);
nor UO_1693 (O_1693,N_49793,N_47945);
nand UO_1694 (O_1694,N_49131,N_47762);
nor UO_1695 (O_1695,N_48971,N_48150);
nand UO_1696 (O_1696,N_49721,N_48177);
or UO_1697 (O_1697,N_49032,N_48945);
xor UO_1698 (O_1698,N_49739,N_49848);
nand UO_1699 (O_1699,N_49828,N_47782);
nor UO_1700 (O_1700,N_48636,N_48673);
or UO_1701 (O_1701,N_48383,N_48836);
or UO_1702 (O_1702,N_47521,N_48093);
nand UO_1703 (O_1703,N_49600,N_48204);
nor UO_1704 (O_1704,N_49212,N_49343);
xnor UO_1705 (O_1705,N_49704,N_47720);
and UO_1706 (O_1706,N_48973,N_49153);
or UO_1707 (O_1707,N_48085,N_49366);
and UO_1708 (O_1708,N_47573,N_47967);
xor UO_1709 (O_1709,N_48229,N_48231);
nand UO_1710 (O_1710,N_49784,N_48787);
nor UO_1711 (O_1711,N_49876,N_49814);
nand UO_1712 (O_1712,N_49229,N_48033);
nand UO_1713 (O_1713,N_48861,N_48801);
xor UO_1714 (O_1714,N_49556,N_48431);
and UO_1715 (O_1715,N_47841,N_47815);
and UO_1716 (O_1716,N_48317,N_49005);
and UO_1717 (O_1717,N_49792,N_47654);
nand UO_1718 (O_1718,N_48108,N_48793);
or UO_1719 (O_1719,N_47783,N_48132);
nand UO_1720 (O_1720,N_49698,N_48261);
nor UO_1721 (O_1721,N_49278,N_49821);
nand UO_1722 (O_1722,N_48334,N_49656);
nor UO_1723 (O_1723,N_49988,N_47805);
xnor UO_1724 (O_1724,N_47519,N_49285);
or UO_1725 (O_1725,N_48697,N_48544);
or UO_1726 (O_1726,N_49622,N_48101);
or UO_1727 (O_1727,N_47899,N_47798);
nand UO_1728 (O_1728,N_47905,N_48542);
and UO_1729 (O_1729,N_48174,N_48720);
and UO_1730 (O_1730,N_49852,N_47693);
or UO_1731 (O_1731,N_49263,N_49861);
nand UO_1732 (O_1732,N_49153,N_47564);
nand UO_1733 (O_1733,N_49864,N_49210);
or UO_1734 (O_1734,N_49256,N_47935);
nor UO_1735 (O_1735,N_47873,N_49993);
xor UO_1736 (O_1736,N_49628,N_49846);
nor UO_1737 (O_1737,N_48909,N_47969);
xor UO_1738 (O_1738,N_47902,N_49859);
nor UO_1739 (O_1739,N_48386,N_48794);
or UO_1740 (O_1740,N_49291,N_47526);
nor UO_1741 (O_1741,N_49924,N_49095);
xnor UO_1742 (O_1742,N_48879,N_48945);
or UO_1743 (O_1743,N_48039,N_49282);
or UO_1744 (O_1744,N_47531,N_49665);
nor UO_1745 (O_1745,N_49977,N_49082);
xor UO_1746 (O_1746,N_48817,N_49469);
or UO_1747 (O_1747,N_49351,N_49020);
or UO_1748 (O_1748,N_48160,N_47626);
xnor UO_1749 (O_1749,N_49123,N_49130);
and UO_1750 (O_1750,N_47546,N_48597);
or UO_1751 (O_1751,N_48720,N_47900);
and UO_1752 (O_1752,N_49815,N_49554);
nor UO_1753 (O_1753,N_48088,N_48906);
nand UO_1754 (O_1754,N_49615,N_48351);
xor UO_1755 (O_1755,N_48066,N_49348);
nor UO_1756 (O_1756,N_49566,N_48962);
nor UO_1757 (O_1757,N_48117,N_49066);
xor UO_1758 (O_1758,N_49442,N_47976);
nor UO_1759 (O_1759,N_47809,N_48219);
xnor UO_1760 (O_1760,N_48024,N_47514);
and UO_1761 (O_1761,N_49279,N_49433);
nor UO_1762 (O_1762,N_48387,N_47827);
or UO_1763 (O_1763,N_48061,N_48775);
nor UO_1764 (O_1764,N_49940,N_48463);
nand UO_1765 (O_1765,N_49333,N_49990);
and UO_1766 (O_1766,N_49650,N_48252);
nor UO_1767 (O_1767,N_47848,N_48237);
nor UO_1768 (O_1768,N_49619,N_47909);
and UO_1769 (O_1769,N_49466,N_49206);
nor UO_1770 (O_1770,N_47542,N_47996);
nor UO_1771 (O_1771,N_49326,N_48731);
xnor UO_1772 (O_1772,N_48832,N_49110);
and UO_1773 (O_1773,N_47744,N_49630);
or UO_1774 (O_1774,N_49456,N_48513);
or UO_1775 (O_1775,N_49294,N_47857);
nand UO_1776 (O_1776,N_49990,N_48439);
or UO_1777 (O_1777,N_49128,N_48081);
nor UO_1778 (O_1778,N_48184,N_48620);
or UO_1779 (O_1779,N_49107,N_49388);
nor UO_1780 (O_1780,N_49379,N_48626);
nor UO_1781 (O_1781,N_47921,N_48146);
and UO_1782 (O_1782,N_48515,N_48404);
nand UO_1783 (O_1783,N_49752,N_48736);
nor UO_1784 (O_1784,N_49455,N_48544);
or UO_1785 (O_1785,N_48664,N_48737);
and UO_1786 (O_1786,N_49123,N_49182);
nand UO_1787 (O_1787,N_47835,N_49209);
or UO_1788 (O_1788,N_47852,N_49390);
nand UO_1789 (O_1789,N_49889,N_49103);
nand UO_1790 (O_1790,N_47993,N_48690);
nor UO_1791 (O_1791,N_49103,N_49102);
nor UO_1792 (O_1792,N_49605,N_47712);
xor UO_1793 (O_1793,N_48451,N_49671);
nand UO_1794 (O_1794,N_48157,N_49041);
or UO_1795 (O_1795,N_47577,N_48238);
nand UO_1796 (O_1796,N_47578,N_47926);
and UO_1797 (O_1797,N_47506,N_48692);
and UO_1798 (O_1798,N_49129,N_49530);
nor UO_1799 (O_1799,N_48548,N_49323);
nand UO_1800 (O_1800,N_48378,N_48892);
nand UO_1801 (O_1801,N_48103,N_47555);
xor UO_1802 (O_1802,N_49489,N_49144);
nor UO_1803 (O_1803,N_48376,N_48464);
xor UO_1804 (O_1804,N_47889,N_49071);
nor UO_1805 (O_1805,N_48948,N_48978);
and UO_1806 (O_1806,N_48974,N_47913);
nor UO_1807 (O_1807,N_49518,N_49351);
or UO_1808 (O_1808,N_47615,N_47913);
xor UO_1809 (O_1809,N_47648,N_48166);
and UO_1810 (O_1810,N_48507,N_48771);
or UO_1811 (O_1811,N_47533,N_49067);
nand UO_1812 (O_1812,N_47637,N_48437);
and UO_1813 (O_1813,N_47993,N_48575);
or UO_1814 (O_1814,N_48458,N_47508);
nor UO_1815 (O_1815,N_49576,N_47770);
and UO_1816 (O_1816,N_48697,N_48442);
and UO_1817 (O_1817,N_49968,N_48195);
xnor UO_1818 (O_1818,N_49639,N_48496);
xnor UO_1819 (O_1819,N_48264,N_49472);
nor UO_1820 (O_1820,N_48547,N_49783);
xnor UO_1821 (O_1821,N_47727,N_49758);
nor UO_1822 (O_1822,N_47520,N_48032);
nor UO_1823 (O_1823,N_49305,N_49315);
nor UO_1824 (O_1824,N_47893,N_49330);
xor UO_1825 (O_1825,N_49636,N_49484);
xnor UO_1826 (O_1826,N_49788,N_49064);
and UO_1827 (O_1827,N_48782,N_48678);
nand UO_1828 (O_1828,N_48801,N_49787);
nand UO_1829 (O_1829,N_48516,N_48857);
or UO_1830 (O_1830,N_48497,N_48043);
nand UO_1831 (O_1831,N_49429,N_47663);
nor UO_1832 (O_1832,N_47795,N_49965);
nand UO_1833 (O_1833,N_48245,N_48395);
and UO_1834 (O_1834,N_49232,N_48426);
nand UO_1835 (O_1835,N_49818,N_48643);
nand UO_1836 (O_1836,N_49637,N_48747);
nand UO_1837 (O_1837,N_49732,N_49435);
and UO_1838 (O_1838,N_48623,N_47833);
xor UO_1839 (O_1839,N_47624,N_47555);
nor UO_1840 (O_1840,N_49039,N_49462);
or UO_1841 (O_1841,N_47924,N_48547);
xor UO_1842 (O_1842,N_48082,N_49616);
or UO_1843 (O_1843,N_49828,N_48016);
or UO_1844 (O_1844,N_48079,N_48515);
nand UO_1845 (O_1845,N_48700,N_49419);
or UO_1846 (O_1846,N_48047,N_48356);
and UO_1847 (O_1847,N_48166,N_47910);
or UO_1848 (O_1848,N_49825,N_49277);
xor UO_1849 (O_1849,N_48603,N_49616);
xnor UO_1850 (O_1850,N_47606,N_48152);
or UO_1851 (O_1851,N_49269,N_48605);
nor UO_1852 (O_1852,N_48470,N_49475);
nor UO_1853 (O_1853,N_48420,N_47563);
nor UO_1854 (O_1854,N_48593,N_48561);
xor UO_1855 (O_1855,N_47845,N_49872);
nor UO_1856 (O_1856,N_47959,N_47538);
and UO_1857 (O_1857,N_48049,N_48354);
or UO_1858 (O_1858,N_48080,N_49769);
or UO_1859 (O_1859,N_49074,N_49811);
nor UO_1860 (O_1860,N_47796,N_48665);
nor UO_1861 (O_1861,N_49298,N_47894);
xor UO_1862 (O_1862,N_48105,N_49871);
xnor UO_1863 (O_1863,N_49566,N_47575);
and UO_1864 (O_1864,N_48595,N_49639);
nor UO_1865 (O_1865,N_49124,N_48994);
nor UO_1866 (O_1866,N_49695,N_49941);
xor UO_1867 (O_1867,N_47868,N_49023);
nor UO_1868 (O_1868,N_47843,N_48724);
nor UO_1869 (O_1869,N_49976,N_48509);
nor UO_1870 (O_1870,N_48247,N_47656);
xor UO_1871 (O_1871,N_49893,N_47560);
and UO_1872 (O_1872,N_47935,N_47579);
or UO_1873 (O_1873,N_48339,N_49630);
or UO_1874 (O_1874,N_47811,N_48467);
and UO_1875 (O_1875,N_49398,N_49283);
or UO_1876 (O_1876,N_48827,N_49022);
or UO_1877 (O_1877,N_49675,N_48572);
nor UO_1878 (O_1878,N_48470,N_48425);
and UO_1879 (O_1879,N_47697,N_47742);
or UO_1880 (O_1880,N_49929,N_49316);
or UO_1881 (O_1881,N_49771,N_49783);
or UO_1882 (O_1882,N_49477,N_49638);
and UO_1883 (O_1883,N_49205,N_48672);
xor UO_1884 (O_1884,N_48338,N_48997);
and UO_1885 (O_1885,N_49969,N_49486);
nor UO_1886 (O_1886,N_49417,N_48267);
and UO_1887 (O_1887,N_48784,N_48530);
xor UO_1888 (O_1888,N_48006,N_47889);
and UO_1889 (O_1889,N_47781,N_48037);
and UO_1890 (O_1890,N_47690,N_49168);
nand UO_1891 (O_1891,N_48287,N_49244);
and UO_1892 (O_1892,N_49311,N_47905);
or UO_1893 (O_1893,N_48303,N_48051);
and UO_1894 (O_1894,N_49622,N_48768);
or UO_1895 (O_1895,N_49277,N_48397);
and UO_1896 (O_1896,N_48030,N_47708);
and UO_1897 (O_1897,N_48684,N_47525);
or UO_1898 (O_1898,N_48898,N_48146);
nand UO_1899 (O_1899,N_47658,N_49053);
nor UO_1900 (O_1900,N_48703,N_49467);
nand UO_1901 (O_1901,N_47737,N_49854);
and UO_1902 (O_1902,N_48064,N_48700);
xor UO_1903 (O_1903,N_48568,N_48372);
nand UO_1904 (O_1904,N_49320,N_47667);
or UO_1905 (O_1905,N_49884,N_49501);
xnor UO_1906 (O_1906,N_47897,N_48255);
nand UO_1907 (O_1907,N_49584,N_49596);
and UO_1908 (O_1908,N_49909,N_48385);
and UO_1909 (O_1909,N_49669,N_49376);
xnor UO_1910 (O_1910,N_48546,N_47701);
and UO_1911 (O_1911,N_47827,N_48676);
nor UO_1912 (O_1912,N_49081,N_49243);
nand UO_1913 (O_1913,N_47998,N_47625);
nand UO_1914 (O_1914,N_47590,N_47857);
nor UO_1915 (O_1915,N_48746,N_48210);
nand UO_1916 (O_1916,N_49056,N_49777);
and UO_1917 (O_1917,N_49219,N_49141);
and UO_1918 (O_1918,N_49075,N_48782);
nor UO_1919 (O_1919,N_47543,N_49127);
nor UO_1920 (O_1920,N_47722,N_49213);
nor UO_1921 (O_1921,N_49629,N_49049);
and UO_1922 (O_1922,N_48670,N_49591);
xnor UO_1923 (O_1923,N_49145,N_48183);
nor UO_1924 (O_1924,N_48829,N_47647);
xor UO_1925 (O_1925,N_48140,N_49048);
and UO_1926 (O_1926,N_49341,N_48715);
nand UO_1927 (O_1927,N_49795,N_48508);
xor UO_1928 (O_1928,N_47755,N_49758);
xnor UO_1929 (O_1929,N_49509,N_48674);
nand UO_1930 (O_1930,N_48112,N_47630);
xnor UO_1931 (O_1931,N_49675,N_47734);
nand UO_1932 (O_1932,N_49910,N_48152);
nor UO_1933 (O_1933,N_49334,N_49940);
xor UO_1934 (O_1934,N_49719,N_48464);
nand UO_1935 (O_1935,N_48626,N_49068);
or UO_1936 (O_1936,N_48021,N_47976);
or UO_1937 (O_1937,N_49607,N_48388);
nand UO_1938 (O_1938,N_48093,N_48207);
or UO_1939 (O_1939,N_48274,N_47783);
xor UO_1940 (O_1940,N_48618,N_48873);
or UO_1941 (O_1941,N_48689,N_47725);
nor UO_1942 (O_1942,N_49293,N_49432);
nand UO_1943 (O_1943,N_48434,N_47528);
or UO_1944 (O_1944,N_47866,N_49178);
and UO_1945 (O_1945,N_47999,N_47901);
nand UO_1946 (O_1946,N_49436,N_49190);
or UO_1947 (O_1947,N_48079,N_47529);
nand UO_1948 (O_1948,N_49594,N_48336);
and UO_1949 (O_1949,N_49555,N_49184);
xor UO_1950 (O_1950,N_49383,N_48800);
nor UO_1951 (O_1951,N_47915,N_48945);
xor UO_1952 (O_1952,N_49124,N_49772);
nand UO_1953 (O_1953,N_49526,N_49730);
nor UO_1954 (O_1954,N_47822,N_49285);
xnor UO_1955 (O_1955,N_49306,N_48921);
and UO_1956 (O_1956,N_49568,N_48587);
or UO_1957 (O_1957,N_48090,N_48120);
and UO_1958 (O_1958,N_48622,N_49931);
xnor UO_1959 (O_1959,N_48620,N_49716);
xnor UO_1960 (O_1960,N_48408,N_49874);
and UO_1961 (O_1961,N_49792,N_49315);
nand UO_1962 (O_1962,N_49747,N_47812);
and UO_1963 (O_1963,N_47549,N_49509);
xor UO_1964 (O_1964,N_49801,N_48399);
xnor UO_1965 (O_1965,N_49797,N_49013);
xor UO_1966 (O_1966,N_47713,N_47550);
and UO_1967 (O_1967,N_49308,N_48463);
nor UO_1968 (O_1968,N_49507,N_48079);
nand UO_1969 (O_1969,N_47518,N_48659);
xor UO_1970 (O_1970,N_48479,N_49049);
xnor UO_1971 (O_1971,N_49119,N_47622);
or UO_1972 (O_1972,N_48993,N_49074);
and UO_1973 (O_1973,N_48012,N_48226);
and UO_1974 (O_1974,N_47625,N_48845);
xor UO_1975 (O_1975,N_48390,N_47718);
and UO_1976 (O_1976,N_49655,N_48061);
nand UO_1977 (O_1977,N_48400,N_47746);
nand UO_1978 (O_1978,N_49789,N_47913);
or UO_1979 (O_1979,N_49852,N_49944);
nand UO_1980 (O_1980,N_49834,N_49425);
and UO_1981 (O_1981,N_48336,N_48948);
nor UO_1982 (O_1982,N_49415,N_48667);
and UO_1983 (O_1983,N_49087,N_47901);
xor UO_1984 (O_1984,N_48775,N_49338);
or UO_1985 (O_1985,N_49383,N_47598);
xor UO_1986 (O_1986,N_48380,N_49964);
nand UO_1987 (O_1987,N_48113,N_49574);
and UO_1988 (O_1988,N_49562,N_48217);
xor UO_1989 (O_1989,N_47662,N_48663);
xor UO_1990 (O_1990,N_49395,N_48279);
or UO_1991 (O_1991,N_47711,N_47877);
nand UO_1992 (O_1992,N_49703,N_48806);
nor UO_1993 (O_1993,N_49385,N_49612);
nor UO_1994 (O_1994,N_48157,N_47556);
nor UO_1995 (O_1995,N_49048,N_49239);
nand UO_1996 (O_1996,N_49348,N_49059);
and UO_1997 (O_1997,N_49224,N_48549);
nand UO_1998 (O_1998,N_48867,N_48262);
xnor UO_1999 (O_1999,N_48297,N_48407);
xor UO_2000 (O_2000,N_49429,N_47963);
nand UO_2001 (O_2001,N_49137,N_47982);
nor UO_2002 (O_2002,N_49981,N_49979);
nor UO_2003 (O_2003,N_48083,N_48879);
and UO_2004 (O_2004,N_48962,N_49504);
nor UO_2005 (O_2005,N_48026,N_48221);
nand UO_2006 (O_2006,N_49098,N_48151);
or UO_2007 (O_2007,N_48075,N_47644);
nand UO_2008 (O_2008,N_47942,N_49644);
xnor UO_2009 (O_2009,N_49621,N_48984);
nor UO_2010 (O_2010,N_49916,N_49171);
nand UO_2011 (O_2011,N_48381,N_47527);
nor UO_2012 (O_2012,N_48862,N_49270);
xor UO_2013 (O_2013,N_48277,N_48291);
nand UO_2014 (O_2014,N_48075,N_49244);
and UO_2015 (O_2015,N_49745,N_48643);
or UO_2016 (O_2016,N_49198,N_48823);
nor UO_2017 (O_2017,N_47956,N_49363);
xnor UO_2018 (O_2018,N_47582,N_49145);
or UO_2019 (O_2019,N_48837,N_48127);
or UO_2020 (O_2020,N_48038,N_49491);
or UO_2021 (O_2021,N_49431,N_48665);
nand UO_2022 (O_2022,N_49014,N_47863);
and UO_2023 (O_2023,N_49433,N_48836);
or UO_2024 (O_2024,N_48296,N_49490);
nor UO_2025 (O_2025,N_47821,N_48062);
xor UO_2026 (O_2026,N_48936,N_48222);
xnor UO_2027 (O_2027,N_49060,N_48704);
nand UO_2028 (O_2028,N_49023,N_49905);
or UO_2029 (O_2029,N_47808,N_49646);
nand UO_2030 (O_2030,N_49106,N_48692);
nor UO_2031 (O_2031,N_49678,N_47858);
nand UO_2032 (O_2032,N_49391,N_48270);
xnor UO_2033 (O_2033,N_48150,N_49513);
nor UO_2034 (O_2034,N_47558,N_49228);
and UO_2035 (O_2035,N_48643,N_48633);
xnor UO_2036 (O_2036,N_48590,N_47929);
xor UO_2037 (O_2037,N_49094,N_49725);
nor UO_2038 (O_2038,N_47583,N_49496);
or UO_2039 (O_2039,N_48312,N_47970);
xnor UO_2040 (O_2040,N_48455,N_49057);
xnor UO_2041 (O_2041,N_48947,N_48649);
nand UO_2042 (O_2042,N_47846,N_48978);
and UO_2043 (O_2043,N_48354,N_49816);
and UO_2044 (O_2044,N_48166,N_47894);
nand UO_2045 (O_2045,N_49093,N_49656);
or UO_2046 (O_2046,N_48202,N_47749);
xnor UO_2047 (O_2047,N_47647,N_49964);
xor UO_2048 (O_2048,N_47889,N_48956);
xor UO_2049 (O_2049,N_48953,N_48779);
nor UO_2050 (O_2050,N_49480,N_49485);
xor UO_2051 (O_2051,N_48688,N_49930);
or UO_2052 (O_2052,N_49224,N_49142);
or UO_2053 (O_2053,N_48803,N_48870);
or UO_2054 (O_2054,N_48953,N_48597);
and UO_2055 (O_2055,N_49827,N_49485);
nor UO_2056 (O_2056,N_48229,N_48836);
nand UO_2057 (O_2057,N_49521,N_49105);
xnor UO_2058 (O_2058,N_49426,N_47911);
and UO_2059 (O_2059,N_47581,N_48086);
or UO_2060 (O_2060,N_48334,N_49021);
or UO_2061 (O_2061,N_49075,N_48636);
xnor UO_2062 (O_2062,N_49375,N_49181);
xnor UO_2063 (O_2063,N_48316,N_49293);
or UO_2064 (O_2064,N_48171,N_48639);
nand UO_2065 (O_2065,N_48565,N_48741);
or UO_2066 (O_2066,N_47785,N_49704);
or UO_2067 (O_2067,N_47911,N_47663);
and UO_2068 (O_2068,N_47593,N_49847);
nand UO_2069 (O_2069,N_48344,N_47840);
xnor UO_2070 (O_2070,N_49085,N_47974);
xnor UO_2071 (O_2071,N_49192,N_48105);
nand UO_2072 (O_2072,N_48264,N_47950);
xnor UO_2073 (O_2073,N_47843,N_49560);
xor UO_2074 (O_2074,N_48627,N_48465);
xnor UO_2075 (O_2075,N_48995,N_48747);
nand UO_2076 (O_2076,N_48387,N_48582);
and UO_2077 (O_2077,N_48274,N_47902);
and UO_2078 (O_2078,N_48801,N_48723);
nand UO_2079 (O_2079,N_48475,N_47712);
xor UO_2080 (O_2080,N_48805,N_49010);
nand UO_2081 (O_2081,N_49907,N_49100);
xnor UO_2082 (O_2082,N_49461,N_47538);
nor UO_2083 (O_2083,N_48150,N_49322);
and UO_2084 (O_2084,N_48679,N_48310);
xor UO_2085 (O_2085,N_47919,N_47917);
nand UO_2086 (O_2086,N_48466,N_47894);
nor UO_2087 (O_2087,N_49292,N_48962);
or UO_2088 (O_2088,N_48429,N_48486);
and UO_2089 (O_2089,N_48330,N_47860);
nand UO_2090 (O_2090,N_49536,N_49065);
xnor UO_2091 (O_2091,N_49203,N_48747);
and UO_2092 (O_2092,N_49218,N_49244);
nor UO_2093 (O_2093,N_49004,N_48187);
or UO_2094 (O_2094,N_49227,N_48696);
nor UO_2095 (O_2095,N_48131,N_49411);
or UO_2096 (O_2096,N_48929,N_49662);
nand UO_2097 (O_2097,N_48722,N_47562);
and UO_2098 (O_2098,N_48244,N_48986);
xor UO_2099 (O_2099,N_49484,N_49490);
or UO_2100 (O_2100,N_48854,N_48480);
and UO_2101 (O_2101,N_48247,N_49727);
and UO_2102 (O_2102,N_48117,N_49886);
nand UO_2103 (O_2103,N_47595,N_49486);
xor UO_2104 (O_2104,N_47792,N_47780);
xor UO_2105 (O_2105,N_49314,N_48383);
and UO_2106 (O_2106,N_49814,N_47855);
and UO_2107 (O_2107,N_47614,N_48727);
or UO_2108 (O_2108,N_48542,N_47543);
nor UO_2109 (O_2109,N_49330,N_47557);
nor UO_2110 (O_2110,N_49400,N_48880);
nor UO_2111 (O_2111,N_47944,N_48667);
xnor UO_2112 (O_2112,N_47818,N_48702);
nor UO_2113 (O_2113,N_49725,N_48755);
or UO_2114 (O_2114,N_47685,N_48647);
xnor UO_2115 (O_2115,N_47746,N_47992);
nand UO_2116 (O_2116,N_49472,N_49947);
or UO_2117 (O_2117,N_47535,N_49184);
and UO_2118 (O_2118,N_47926,N_49565);
nand UO_2119 (O_2119,N_48522,N_48433);
and UO_2120 (O_2120,N_48307,N_49608);
nor UO_2121 (O_2121,N_49143,N_48732);
nand UO_2122 (O_2122,N_49078,N_48439);
nand UO_2123 (O_2123,N_48583,N_47753);
nand UO_2124 (O_2124,N_49344,N_48190);
and UO_2125 (O_2125,N_48025,N_49271);
xor UO_2126 (O_2126,N_48115,N_47605);
or UO_2127 (O_2127,N_48727,N_48919);
or UO_2128 (O_2128,N_49597,N_48624);
and UO_2129 (O_2129,N_47602,N_49618);
nor UO_2130 (O_2130,N_48814,N_49910);
and UO_2131 (O_2131,N_47927,N_48155);
xor UO_2132 (O_2132,N_49247,N_48703);
or UO_2133 (O_2133,N_47990,N_47572);
xnor UO_2134 (O_2134,N_49974,N_49108);
nor UO_2135 (O_2135,N_49180,N_49534);
xnor UO_2136 (O_2136,N_48130,N_49487);
nor UO_2137 (O_2137,N_49183,N_48938);
nor UO_2138 (O_2138,N_48305,N_48762);
nor UO_2139 (O_2139,N_47745,N_49743);
and UO_2140 (O_2140,N_48791,N_48316);
and UO_2141 (O_2141,N_49897,N_49119);
nor UO_2142 (O_2142,N_48256,N_48493);
nor UO_2143 (O_2143,N_47791,N_47841);
xor UO_2144 (O_2144,N_49852,N_48752);
or UO_2145 (O_2145,N_49624,N_47771);
or UO_2146 (O_2146,N_47839,N_48816);
nand UO_2147 (O_2147,N_48258,N_49398);
or UO_2148 (O_2148,N_49714,N_49115);
nor UO_2149 (O_2149,N_49750,N_48591);
nor UO_2150 (O_2150,N_49771,N_48144);
nand UO_2151 (O_2151,N_48558,N_49340);
nor UO_2152 (O_2152,N_49938,N_48274);
nor UO_2153 (O_2153,N_48652,N_48903);
xor UO_2154 (O_2154,N_48985,N_49789);
nor UO_2155 (O_2155,N_48289,N_48185);
or UO_2156 (O_2156,N_49379,N_48503);
nand UO_2157 (O_2157,N_48553,N_48094);
nor UO_2158 (O_2158,N_48617,N_49239);
and UO_2159 (O_2159,N_47519,N_48579);
and UO_2160 (O_2160,N_48311,N_48100);
nor UO_2161 (O_2161,N_48407,N_49898);
and UO_2162 (O_2162,N_49697,N_49097);
xnor UO_2163 (O_2163,N_47508,N_49029);
xor UO_2164 (O_2164,N_49353,N_48198);
xor UO_2165 (O_2165,N_48812,N_47785);
and UO_2166 (O_2166,N_49843,N_47594);
nor UO_2167 (O_2167,N_49728,N_48473);
nand UO_2168 (O_2168,N_49381,N_49849);
nor UO_2169 (O_2169,N_49491,N_48851);
or UO_2170 (O_2170,N_49209,N_48177);
nor UO_2171 (O_2171,N_49037,N_49702);
and UO_2172 (O_2172,N_49784,N_48189);
and UO_2173 (O_2173,N_49959,N_47516);
or UO_2174 (O_2174,N_48852,N_47685);
and UO_2175 (O_2175,N_49624,N_47956);
and UO_2176 (O_2176,N_49807,N_49062);
and UO_2177 (O_2177,N_47726,N_49164);
and UO_2178 (O_2178,N_48461,N_48842);
and UO_2179 (O_2179,N_49751,N_47539);
or UO_2180 (O_2180,N_48096,N_49029);
nor UO_2181 (O_2181,N_48937,N_47754);
nor UO_2182 (O_2182,N_49739,N_47787);
or UO_2183 (O_2183,N_49348,N_48109);
nor UO_2184 (O_2184,N_49533,N_49839);
xor UO_2185 (O_2185,N_49411,N_48226);
nor UO_2186 (O_2186,N_49487,N_49577);
nand UO_2187 (O_2187,N_48090,N_47842);
nand UO_2188 (O_2188,N_48748,N_48590);
nand UO_2189 (O_2189,N_49541,N_48002);
nor UO_2190 (O_2190,N_49853,N_49135);
nand UO_2191 (O_2191,N_48518,N_48953);
xnor UO_2192 (O_2192,N_48654,N_49716);
nor UO_2193 (O_2193,N_49918,N_47810);
nand UO_2194 (O_2194,N_49020,N_47968);
nand UO_2195 (O_2195,N_47975,N_48083);
xor UO_2196 (O_2196,N_49421,N_48736);
or UO_2197 (O_2197,N_49069,N_49830);
nor UO_2198 (O_2198,N_49745,N_48168);
or UO_2199 (O_2199,N_49522,N_48693);
and UO_2200 (O_2200,N_49130,N_47815);
nand UO_2201 (O_2201,N_49613,N_49147);
or UO_2202 (O_2202,N_47765,N_48328);
nor UO_2203 (O_2203,N_49810,N_47759);
nor UO_2204 (O_2204,N_47780,N_48607);
nand UO_2205 (O_2205,N_49579,N_48873);
xnor UO_2206 (O_2206,N_48624,N_48684);
and UO_2207 (O_2207,N_48032,N_48501);
or UO_2208 (O_2208,N_48650,N_48209);
and UO_2209 (O_2209,N_49968,N_49030);
nor UO_2210 (O_2210,N_49989,N_49313);
nand UO_2211 (O_2211,N_48918,N_48284);
or UO_2212 (O_2212,N_49772,N_49418);
or UO_2213 (O_2213,N_48436,N_49712);
nor UO_2214 (O_2214,N_48966,N_48820);
nand UO_2215 (O_2215,N_47828,N_49341);
or UO_2216 (O_2216,N_49885,N_49083);
and UO_2217 (O_2217,N_49523,N_49586);
nor UO_2218 (O_2218,N_49757,N_48181);
nand UO_2219 (O_2219,N_48055,N_49858);
nor UO_2220 (O_2220,N_49596,N_48679);
nor UO_2221 (O_2221,N_49599,N_48547);
and UO_2222 (O_2222,N_47800,N_47688);
or UO_2223 (O_2223,N_48613,N_48985);
xnor UO_2224 (O_2224,N_47757,N_49249);
xnor UO_2225 (O_2225,N_49836,N_47819);
xnor UO_2226 (O_2226,N_47847,N_47531);
nor UO_2227 (O_2227,N_47729,N_47749);
or UO_2228 (O_2228,N_48518,N_49979);
and UO_2229 (O_2229,N_49707,N_47606);
and UO_2230 (O_2230,N_48358,N_48610);
nand UO_2231 (O_2231,N_49768,N_49174);
nand UO_2232 (O_2232,N_48434,N_48127);
nor UO_2233 (O_2233,N_48119,N_48300);
nor UO_2234 (O_2234,N_48396,N_48991);
xnor UO_2235 (O_2235,N_49629,N_49869);
nor UO_2236 (O_2236,N_49710,N_49678);
nand UO_2237 (O_2237,N_49514,N_49527);
xor UO_2238 (O_2238,N_49532,N_49182);
and UO_2239 (O_2239,N_49873,N_49476);
nand UO_2240 (O_2240,N_49954,N_48416);
nand UO_2241 (O_2241,N_47790,N_48908);
nor UO_2242 (O_2242,N_48625,N_49246);
nor UO_2243 (O_2243,N_48400,N_48032);
or UO_2244 (O_2244,N_48186,N_48924);
nand UO_2245 (O_2245,N_47901,N_47791);
xnor UO_2246 (O_2246,N_49903,N_49054);
nand UO_2247 (O_2247,N_48647,N_49858);
nand UO_2248 (O_2248,N_49484,N_48565);
xnor UO_2249 (O_2249,N_47735,N_48447);
or UO_2250 (O_2250,N_48092,N_49963);
nand UO_2251 (O_2251,N_48422,N_48603);
nand UO_2252 (O_2252,N_47563,N_48440);
nor UO_2253 (O_2253,N_49423,N_49839);
nand UO_2254 (O_2254,N_47679,N_49470);
or UO_2255 (O_2255,N_49037,N_49513);
and UO_2256 (O_2256,N_49710,N_49582);
and UO_2257 (O_2257,N_48691,N_49317);
or UO_2258 (O_2258,N_48555,N_49873);
nor UO_2259 (O_2259,N_49650,N_49258);
nand UO_2260 (O_2260,N_48633,N_49909);
nor UO_2261 (O_2261,N_49868,N_48673);
nor UO_2262 (O_2262,N_47633,N_48763);
and UO_2263 (O_2263,N_49018,N_48525);
or UO_2264 (O_2264,N_48919,N_49221);
nor UO_2265 (O_2265,N_49777,N_49520);
or UO_2266 (O_2266,N_49633,N_49011);
or UO_2267 (O_2267,N_47861,N_48645);
or UO_2268 (O_2268,N_49865,N_48191);
or UO_2269 (O_2269,N_47738,N_48836);
nor UO_2270 (O_2270,N_47855,N_48461);
xor UO_2271 (O_2271,N_48921,N_49287);
nand UO_2272 (O_2272,N_47738,N_49083);
nor UO_2273 (O_2273,N_48746,N_49513);
and UO_2274 (O_2274,N_48314,N_49301);
and UO_2275 (O_2275,N_49943,N_48758);
nand UO_2276 (O_2276,N_49911,N_49006);
xnor UO_2277 (O_2277,N_48643,N_48447);
nor UO_2278 (O_2278,N_48094,N_48481);
nor UO_2279 (O_2279,N_47879,N_49726);
nand UO_2280 (O_2280,N_47522,N_49856);
or UO_2281 (O_2281,N_49644,N_48373);
or UO_2282 (O_2282,N_47543,N_48723);
or UO_2283 (O_2283,N_49342,N_49078);
and UO_2284 (O_2284,N_48932,N_47733);
and UO_2285 (O_2285,N_49511,N_48061);
nand UO_2286 (O_2286,N_49296,N_49110);
nor UO_2287 (O_2287,N_49845,N_47989);
or UO_2288 (O_2288,N_47735,N_48107);
xor UO_2289 (O_2289,N_48800,N_47806);
nor UO_2290 (O_2290,N_48851,N_47801);
nor UO_2291 (O_2291,N_48929,N_48868);
xor UO_2292 (O_2292,N_49248,N_48462);
and UO_2293 (O_2293,N_49417,N_48775);
xor UO_2294 (O_2294,N_47601,N_48648);
nand UO_2295 (O_2295,N_49549,N_49666);
and UO_2296 (O_2296,N_48879,N_48713);
nand UO_2297 (O_2297,N_47876,N_48558);
or UO_2298 (O_2298,N_49664,N_48282);
nor UO_2299 (O_2299,N_49242,N_48387);
xnor UO_2300 (O_2300,N_47962,N_49248);
or UO_2301 (O_2301,N_48215,N_48191);
or UO_2302 (O_2302,N_48520,N_48604);
xor UO_2303 (O_2303,N_48672,N_49231);
xor UO_2304 (O_2304,N_49562,N_49076);
and UO_2305 (O_2305,N_49501,N_48490);
nor UO_2306 (O_2306,N_47953,N_48553);
nand UO_2307 (O_2307,N_47812,N_48356);
xnor UO_2308 (O_2308,N_49032,N_49351);
and UO_2309 (O_2309,N_49446,N_48379);
nor UO_2310 (O_2310,N_48688,N_48954);
nor UO_2311 (O_2311,N_49889,N_49187);
and UO_2312 (O_2312,N_48599,N_49085);
nand UO_2313 (O_2313,N_47511,N_49512);
xor UO_2314 (O_2314,N_49030,N_49435);
or UO_2315 (O_2315,N_48407,N_48041);
xor UO_2316 (O_2316,N_48541,N_49769);
or UO_2317 (O_2317,N_48471,N_49761);
or UO_2318 (O_2318,N_49296,N_49718);
nor UO_2319 (O_2319,N_48582,N_48029);
nor UO_2320 (O_2320,N_48877,N_47531);
or UO_2321 (O_2321,N_48234,N_49750);
and UO_2322 (O_2322,N_49855,N_47680);
xor UO_2323 (O_2323,N_49457,N_48401);
xor UO_2324 (O_2324,N_49921,N_49376);
xor UO_2325 (O_2325,N_47931,N_49743);
and UO_2326 (O_2326,N_48549,N_47590);
xnor UO_2327 (O_2327,N_49399,N_48938);
nor UO_2328 (O_2328,N_49978,N_47562);
xnor UO_2329 (O_2329,N_48209,N_48713);
nand UO_2330 (O_2330,N_48689,N_48619);
or UO_2331 (O_2331,N_49692,N_49500);
and UO_2332 (O_2332,N_47603,N_48475);
xor UO_2333 (O_2333,N_48539,N_49961);
xor UO_2334 (O_2334,N_49580,N_48946);
or UO_2335 (O_2335,N_48364,N_49900);
or UO_2336 (O_2336,N_48623,N_49130);
or UO_2337 (O_2337,N_48877,N_48204);
nor UO_2338 (O_2338,N_47575,N_48773);
xor UO_2339 (O_2339,N_48630,N_48611);
nor UO_2340 (O_2340,N_48151,N_49258);
nand UO_2341 (O_2341,N_48657,N_48760);
nor UO_2342 (O_2342,N_48769,N_49761);
or UO_2343 (O_2343,N_47511,N_49711);
or UO_2344 (O_2344,N_49219,N_49458);
xor UO_2345 (O_2345,N_47531,N_49765);
or UO_2346 (O_2346,N_48347,N_47923);
and UO_2347 (O_2347,N_49980,N_49624);
xnor UO_2348 (O_2348,N_49767,N_47784);
and UO_2349 (O_2349,N_48342,N_48360);
nand UO_2350 (O_2350,N_47840,N_48865);
xor UO_2351 (O_2351,N_49106,N_47674);
nor UO_2352 (O_2352,N_48866,N_49165);
nor UO_2353 (O_2353,N_48031,N_47768);
and UO_2354 (O_2354,N_47974,N_49027);
and UO_2355 (O_2355,N_49728,N_47979);
xor UO_2356 (O_2356,N_49434,N_47777);
xnor UO_2357 (O_2357,N_49632,N_48521);
nor UO_2358 (O_2358,N_47534,N_48307);
and UO_2359 (O_2359,N_49427,N_49328);
and UO_2360 (O_2360,N_48183,N_48266);
xor UO_2361 (O_2361,N_48267,N_48568);
nand UO_2362 (O_2362,N_47918,N_48017);
and UO_2363 (O_2363,N_48164,N_49922);
and UO_2364 (O_2364,N_49178,N_49568);
and UO_2365 (O_2365,N_47843,N_47901);
nor UO_2366 (O_2366,N_48221,N_49688);
xor UO_2367 (O_2367,N_47605,N_48807);
nand UO_2368 (O_2368,N_48649,N_48057);
xor UO_2369 (O_2369,N_48604,N_48974);
or UO_2370 (O_2370,N_47986,N_49441);
nor UO_2371 (O_2371,N_48749,N_47929);
xor UO_2372 (O_2372,N_47695,N_49455);
nand UO_2373 (O_2373,N_49804,N_49458);
nor UO_2374 (O_2374,N_47773,N_49104);
or UO_2375 (O_2375,N_48804,N_49527);
xor UO_2376 (O_2376,N_47767,N_47739);
nor UO_2377 (O_2377,N_47586,N_49666);
nor UO_2378 (O_2378,N_47710,N_48860);
or UO_2379 (O_2379,N_47610,N_49920);
nor UO_2380 (O_2380,N_49115,N_49162);
nand UO_2381 (O_2381,N_48122,N_48107);
or UO_2382 (O_2382,N_48796,N_49660);
xor UO_2383 (O_2383,N_48238,N_48334);
and UO_2384 (O_2384,N_48552,N_47839);
and UO_2385 (O_2385,N_48098,N_48287);
nand UO_2386 (O_2386,N_49080,N_48514);
xnor UO_2387 (O_2387,N_48443,N_49806);
or UO_2388 (O_2388,N_47990,N_49268);
nand UO_2389 (O_2389,N_49466,N_48516);
and UO_2390 (O_2390,N_48328,N_49569);
nor UO_2391 (O_2391,N_48037,N_48146);
nand UO_2392 (O_2392,N_49973,N_49654);
xor UO_2393 (O_2393,N_49625,N_48514);
or UO_2394 (O_2394,N_47980,N_48240);
xnor UO_2395 (O_2395,N_47925,N_47589);
nand UO_2396 (O_2396,N_49217,N_49027);
or UO_2397 (O_2397,N_48225,N_49483);
and UO_2398 (O_2398,N_49086,N_48537);
or UO_2399 (O_2399,N_48425,N_48482);
nor UO_2400 (O_2400,N_48820,N_48968);
nor UO_2401 (O_2401,N_49458,N_49931);
nor UO_2402 (O_2402,N_49629,N_49443);
and UO_2403 (O_2403,N_48434,N_49628);
xor UO_2404 (O_2404,N_48053,N_48568);
nand UO_2405 (O_2405,N_49237,N_49912);
or UO_2406 (O_2406,N_49763,N_49771);
and UO_2407 (O_2407,N_47758,N_47531);
nor UO_2408 (O_2408,N_48742,N_47622);
nor UO_2409 (O_2409,N_48856,N_49303);
xnor UO_2410 (O_2410,N_49744,N_48369);
and UO_2411 (O_2411,N_48245,N_48460);
and UO_2412 (O_2412,N_49865,N_47601);
xor UO_2413 (O_2413,N_47821,N_48486);
xor UO_2414 (O_2414,N_48433,N_49963);
xor UO_2415 (O_2415,N_48748,N_47572);
nand UO_2416 (O_2416,N_48361,N_49244);
xor UO_2417 (O_2417,N_47672,N_49331);
nor UO_2418 (O_2418,N_47924,N_47878);
or UO_2419 (O_2419,N_47922,N_48111);
xor UO_2420 (O_2420,N_47694,N_48541);
nand UO_2421 (O_2421,N_47906,N_48438);
xor UO_2422 (O_2422,N_47846,N_48301);
nor UO_2423 (O_2423,N_49017,N_49864);
or UO_2424 (O_2424,N_49318,N_48611);
and UO_2425 (O_2425,N_49412,N_48062);
and UO_2426 (O_2426,N_48160,N_49882);
nor UO_2427 (O_2427,N_48647,N_48991);
or UO_2428 (O_2428,N_49504,N_48703);
nand UO_2429 (O_2429,N_49407,N_48319);
nor UO_2430 (O_2430,N_47904,N_49769);
nor UO_2431 (O_2431,N_48929,N_48686);
and UO_2432 (O_2432,N_48206,N_47668);
nor UO_2433 (O_2433,N_48546,N_49097);
nor UO_2434 (O_2434,N_48850,N_47742);
nor UO_2435 (O_2435,N_48787,N_49581);
nand UO_2436 (O_2436,N_49759,N_49511);
xor UO_2437 (O_2437,N_48277,N_47710);
xnor UO_2438 (O_2438,N_48901,N_48819);
and UO_2439 (O_2439,N_47538,N_48943);
nand UO_2440 (O_2440,N_47504,N_49094);
or UO_2441 (O_2441,N_49972,N_49681);
or UO_2442 (O_2442,N_48670,N_48062);
nand UO_2443 (O_2443,N_47598,N_48194);
nor UO_2444 (O_2444,N_48050,N_48889);
nor UO_2445 (O_2445,N_49216,N_48352);
and UO_2446 (O_2446,N_48667,N_48806);
or UO_2447 (O_2447,N_48300,N_49068);
xor UO_2448 (O_2448,N_49187,N_47909);
and UO_2449 (O_2449,N_49938,N_48322);
xnor UO_2450 (O_2450,N_48408,N_47710);
or UO_2451 (O_2451,N_47992,N_47938);
nor UO_2452 (O_2452,N_48420,N_49025);
xnor UO_2453 (O_2453,N_49363,N_48040);
xor UO_2454 (O_2454,N_47988,N_47522);
and UO_2455 (O_2455,N_48643,N_49086);
or UO_2456 (O_2456,N_47902,N_47811);
and UO_2457 (O_2457,N_48109,N_49451);
and UO_2458 (O_2458,N_49130,N_47769);
and UO_2459 (O_2459,N_49776,N_47532);
xnor UO_2460 (O_2460,N_48227,N_49395);
and UO_2461 (O_2461,N_48069,N_49676);
and UO_2462 (O_2462,N_47773,N_48728);
xor UO_2463 (O_2463,N_49879,N_48805);
and UO_2464 (O_2464,N_49085,N_49499);
nand UO_2465 (O_2465,N_49960,N_49001);
or UO_2466 (O_2466,N_47875,N_49389);
nand UO_2467 (O_2467,N_49993,N_49243);
or UO_2468 (O_2468,N_48232,N_48479);
xnor UO_2469 (O_2469,N_49950,N_48816);
or UO_2470 (O_2470,N_48003,N_47807);
nor UO_2471 (O_2471,N_48015,N_49153);
and UO_2472 (O_2472,N_48551,N_47572);
or UO_2473 (O_2473,N_47604,N_48276);
or UO_2474 (O_2474,N_48810,N_48041);
or UO_2475 (O_2475,N_48005,N_49992);
or UO_2476 (O_2476,N_48400,N_48931);
and UO_2477 (O_2477,N_49610,N_49798);
or UO_2478 (O_2478,N_49156,N_49622);
and UO_2479 (O_2479,N_49895,N_49693);
or UO_2480 (O_2480,N_47720,N_48813);
and UO_2481 (O_2481,N_49174,N_48045);
or UO_2482 (O_2482,N_49008,N_47747);
xnor UO_2483 (O_2483,N_47793,N_49943);
xor UO_2484 (O_2484,N_49081,N_49559);
xor UO_2485 (O_2485,N_49136,N_49132);
nor UO_2486 (O_2486,N_48133,N_48994);
or UO_2487 (O_2487,N_49081,N_47641);
and UO_2488 (O_2488,N_47503,N_47839);
or UO_2489 (O_2489,N_48914,N_48255);
and UO_2490 (O_2490,N_49143,N_48995);
nand UO_2491 (O_2491,N_47845,N_47660);
nand UO_2492 (O_2492,N_49040,N_48457);
nor UO_2493 (O_2493,N_47876,N_49724);
nand UO_2494 (O_2494,N_48205,N_49156);
nand UO_2495 (O_2495,N_47749,N_48849);
and UO_2496 (O_2496,N_48778,N_48023);
nor UO_2497 (O_2497,N_48053,N_47963);
xor UO_2498 (O_2498,N_47981,N_48140);
or UO_2499 (O_2499,N_49034,N_48585);
or UO_2500 (O_2500,N_48304,N_48060);
nor UO_2501 (O_2501,N_48642,N_49457);
xor UO_2502 (O_2502,N_47703,N_49195);
or UO_2503 (O_2503,N_48569,N_47894);
xnor UO_2504 (O_2504,N_48576,N_49745);
and UO_2505 (O_2505,N_49006,N_48059);
nor UO_2506 (O_2506,N_49603,N_49780);
nor UO_2507 (O_2507,N_47993,N_49041);
and UO_2508 (O_2508,N_48235,N_49688);
nor UO_2509 (O_2509,N_48589,N_48083);
nand UO_2510 (O_2510,N_49669,N_48256);
or UO_2511 (O_2511,N_48955,N_49464);
nand UO_2512 (O_2512,N_47619,N_49004);
nor UO_2513 (O_2513,N_47507,N_49983);
and UO_2514 (O_2514,N_47796,N_48109);
xnor UO_2515 (O_2515,N_48788,N_49582);
and UO_2516 (O_2516,N_48912,N_48948);
or UO_2517 (O_2517,N_47807,N_49486);
nor UO_2518 (O_2518,N_49525,N_48440);
or UO_2519 (O_2519,N_47708,N_49438);
or UO_2520 (O_2520,N_48708,N_47606);
nand UO_2521 (O_2521,N_48818,N_49743);
nand UO_2522 (O_2522,N_48004,N_48055);
nand UO_2523 (O_2523,N_49432,N_49690);
xnor UO_2524 (O_2524,N_47988,N_47818);
nor UO_2525 (O_2525,N_49362,N_48491);
xnor UO_2526 (O_2526,N_47955,N_48011);
xnor UO_2527 (O_2527,N_48716,N_48325);
xor UO_2528 (O_2528,N_47536,N_49115);
or UO_2529 (O_2529,N_48239,N_48822);
xor UO_2530 (O_2530,N_49021,N_48754);
xor UO_2531 (O_2531,N_47912,N_47520);
or UO_2532 (O_2532,N_47719,N_49120);
xor UO_2533 (O_2533,N_49932,N_48038);
and UO_2534 (O_2534,N_48412,N_47819);
nor UO_2535 (O_2535,N_49469,N_49916);
nor UO_2536 (O_2536,N_47902,N_48263);
xnor UO_2537 (O_2537,N_47585,N_49915);
nand UO_2538 (O_2538,N_47844,N_49332);
nand UO_2539 (O_2539,N_47851,N_49342);
nand UO_2540 (O_2540,N_49998,N_47693);
or UO_2541 (O_2541,N_49650,N_47701);
nand UO_2542 (O_2542,N_48058,N_47763);
xor UO_2543 (O_2543,N_49895,N_49640);
or UO_2544 (O_2544,N_48435,N_47892);
nand UO_2545 (O_2545,N_49901,N_49423);
or UO_2546 (O_2546,N_49849,N_48757);
or UO_2547 (O_2547,N_47821,N_47887);
and UO_2548 (O_2548,N_48185,N_48054);
xnor UO_2549 (O_2549,N_47634,N_48651);
nor UO_2550 (O_2550,N_49830,N_49858);
xnor UO_2551 (O_2551,N_49939,N_48209);
or UO_2552 (O_2552,N_49094,N_49194);
nor UO_2553 (O_2553,N_49751,N_49599);
and UO_2554 (O_2554,N_48750,N_49906);
nand UO_2555 (O_2555,N_49215,N_48584);
or UO_2556 (O_2556,N_48474,N_48986);
xnor UO_2557 (O_2557,N_48074,N_47799);
or UO_2558 (O_2558,N_48697,N_48471);
and UO_2559 (O_2559,N_48627,N_48998);
nand UO_2560 (O_2560,N_48594,N_48506);
or UO_2561 (O_2561,N_48181,N_48163);
and UO_2562 (O_2562,N_47577,N_48256);
and UO_2563 (O_2563,N_48866,N_49241);
nand UO_2564 (O_2564,N_48605,N_48325);
or UO_2565 (O_2565,N_49319,N_49799);
and UO_2566 (O_2566,N_48147,N_49367);
nand UO_2567 (O_2567,N_49340,N_49398);
xnor UO_2568 (O_2568,N_47634,N_49122);
xor UO_2569 (O_2569,N_49670,N_49516);
nand UO_2570 (O_2570,N_48395,N_48607);
or UO_2571 (O_2571,N_48808,N_49208);
xnor UO_2572 (O_2572,N_49133,N_49495);
xor UO_2573 (O_2573,N_49922,N_48228);
xor UO_2574 (O_2574,N_49971,N_47552);
and UO_2575 (O_2575,N_49674,N_47671);
and UO_2576 (O_2576,N_49223,N_49987);
xor UO_2577 (O_2577,N_48020,N_49845);
and UO_2578 (O_2578,N_48567,N_47553);
or UO_2579 (O_2579,N_48972,N_49368);
nor UO_2580 (O_2580,N_49067,N_49852);
nor UO_2581 (O_2581,N_47582,N_48547);
nor UO_2582 (O_2582,N_47803,N_47569);
nand UO_2583 (O_2583,N_47521,N_49922);
nand UO_2584 (O_2584,N_48332,N_49475);
xor UO_2585 (O_2585,N_48690,N_48124);
and UO_2586 (O_2586,N_47622,N_48499);
and UO_2587 (O_2587,N_48833,N_49378);
or UO_2588 (O_2588,N_49537,N_48438);
or UO_2589 (O_2589,N_49170,N_49011);
and UO_2590 (O_2590,N_49048,N_48085);
or UO_2591 (O_2591,N_48496,N_47956);
nand UO_2592 (O_2592,N_48424,N_49133);
or UO_2593 (O_2593,N_49833,N_49134);
xor UO_2594 (O_2594,N_48598,N_48364);
nor UO_2595 (O_2595,N_48626,N_48603);
xor UO_2596 (O_2596,N_48309,N_47771);
or UO_2597 (O_2597,N_47582,N_48721);
nor UO_2598 (O_2598,N_48820,N_49184);
and UO_2599 (O_2599,N_49987,N_49485);
nor UO_2600 (O_2600,N_49912,N_47692);
nand UO_2601 (O_2601,N_49235,N_49202);
or UO_2602 (O_2602,N_49320,N_49662);
nand UO_2603 (O_2603,N_49809,N_49039);
nor UO_2604 (O_2604,N_47904,N_49945);
nor UO_2605 (O_2605,N_49986,N_49080);
nand UO_2606 (O_2606,N_49667,N_48499);
or UO_2607 (O_2607,N_49019,N_47583);
nor UO_2608 (O_2608,N_49530,N_49935);
or UO_2609 (O_2609,N_47770,N_47550);
xor UO_2610 (O_2610,N_48804,N_49503);
xor UO_2611 (O_2611,N_47573,N_49663);
and UO_2612 (O_2612,N_48463,N_48606);
and UO_2613 (O_2613,N_49629,N_48282);
xnor UO_2614 (O_2614,N_48152,N_49902);
xor UO_2615 (O_2615,N_49541,N_49397);
xor UO_2616 (O_2616,N_48708,N_49566);
xnor UO_2617 (O_2617,N_49993,N_49819);
nand UO_2618 (O_2618,N_48609,N_48626);
xor UO_2619 (O_2619,N_47705,N_49548);
nor UO_2620 (O_2620,N_49257,N_48531);
xor UO_2621 (O_2621,N_48147,N_49278);
xor UO_2622 (O_2622,N_48125,N_48380);
nor UO_2623 (O_2623,N_49197,N_48001);
or UO_2624 (O_2624,N_48733,N_47792);
and UO_2625 (O_2625,N_48098,N_48442);
nor UO_2626 (O_2626,N_49948,N_49341);
xor UO_2627 (O_2627,N_49402,N_47986);
and UO_2628 (O_2628,N_47869,N_49368);
xor UO_2629 (O_2629,N_48209,N_47923);
and UO_2630 (O_2630,N_49953,N_49135);
and UO_2631 (O_2631,N_48227,N_47588);
xnor UO_2632 (O_2632,N_48842,N_49834);
or UO_2633 (O_2633,N_49655,N_48139);
or UO_2634 (O_2634,N_48794,N_48591);
or UO_2635 (O_2635,N_48934,N_49736);
and UO_2636 (O_2636,N_48303,N_49760);
or UO_2637 (O_2637,N_48863,N_49387);
xnor UO_2638 (O_2638,N_47805,N_48415);
nor UO_2639 (O_2639,N_47811,N_47631);
and UO_2640 (O_2640,N_47909,N_48945);
nor UO_2641 (O_2641,N_47983,N_48474);
nand UO_2642 (O_2642,N_48628,N_48431);
or UO_2643 (O_2643,N_47619,N_49347);
or UO_2644 (O_2644,N_48192,N_49565);
nand UO_2645 (O_2645,N_49809,N_49995);
or UO_2646 (O_2646,N_49853,N_47886);
nor UO_2647 (O_2647,N_49157,N_49465);
nor UO_2648 (O_2648,N_49162,N_47524);
nor UO_2649 (O_2649,N_48206,N_49410);
or UO_2650 (O_2650,N_49722,N_48252);
nor UO_2651 (O_2651,N_49672,N_49538);
or UO_2652 (O_2652,N_49336,N_48527);
nand UO_2653 (O_2653,N_49142,N_49416);
xor UO_2654 (O_2654,N_48042,N_48298);
xor UO_2655 (O_2655,N_49535,N_48708);
or UO_2656 (O_2656,N_48038,N_48182);
and UO_2657 (O_2657,N_47902,N_47960);
or UO_2658 (O_2658,N_49933,N_49237);
and UO_2659 (O_2659,N_48739,N_49397);
xnor UO_2660 (O_2660,N_48827,N_49596);
nor UO_2661 (O_2661,N_48032,N_48865);
and UO_2662 (O_2662,N_49970,N_49070);
xor UO_2663 (O_2663,N_47569,N_49357);
and UO_2664 (O_2664,N_48572,N_47961);
nor UO_2665 (O_2665,N_49570,N_49630);
nand UO_2666 (O_2666,N_47719,N_47980);
and UO_2667 (O_2667,N_48806,N_49163);
and UO_2668 (O_2668,N_49003,N_49602);
nand UO_2669 (O_2669,N_48609,N_47923);
and UO_2670 (O_2670,N_49821,N_48938);
and UO_2671 (O_2671,N_49001,N_47637);
xor UO_2672 (O_2672,N_48652,N_47856);
nand UO_2673 (O_2673,N_48795,N_48664);
nand UO_2674 (O_2674,N_49085,N_48117);
nand UO_2675 (O_2675,N_48956,N_48598);
nor UO_2676 (O_2676,N_48703,N_47957);
and UO_2677 (O_2677,N_49483,N_49894);
and UO_2678 (O_2678,N_49998,N_48494);
and UO_2679 (O_2679,N_49320,N_48302);
nor UO_2680 (O_2680,N_48695,N_49208);
nand UO_2681 (O_2681,N_47792,N_48008);
nor UO_2682 (O_2682,N_49317,N_49453);
xor UO_2683 (O_2683,N_47782,N_49144);
nor UO_2684 (O_2684,N_48161,N_49063);
and UO_2685 (O_2685,N_48150,N_49580);
xnor UO_2686 (O_2686,N_47904,N_47754);
or UO_2687 (O_2687,N_49128,N_47942);
or UO_2688 (O_2688,N_48495,N_48120);
or UO_2689 (O_2689,N_49984,N_49980);
and UO_2690 (O_2690,N_47605,N_48233);
nand UO_2691 (O_2691,N_47876,N_48544);
or UO_2692 (O_2692,N_47768,N_48724);
or UO_2693 (O_2693,N_49090,N_49973);
or UO_2694 (O_2694,N_48373,N_47864);
nor UO_2695 (O_2695,N_47611,N_49826);
or UO_2696 (O_2696,N_48666,N_49266);
xnor UO_2697 (O_2697,N_49473,N_49624);
nand UO_2698 (O_2698,N_47667,N_49033);
nand UO_2699 (O_2699,N_49968,N_49764);
or UO_2700 (O_2700,N_48488,N_49037);
or UO_2701 (O_2701,N_48730,N_49219);
and UO_2702 (O_2702,N_49831,N_49981);
nand UO_2703 (O_2703,N_48627,N_49979);
xor UO_2704 (O_2704,N_49815,N_47575);
and UO_2705 (O_2705,N_48981,N_48715);
xnor UO_2706 (O_2706,N_47904,N_48670);
and UO_2707 (O_2707,N_48106,N_48343);
nand UO_2708 (O_2708,N_49875,N_48971);
xor UO_2709 (O_2709,N_48095,N_48113);
nor UO_2710 (O_2710,N_49630,N_47516);
or UO_2711 (O_2711,N_48482,N_49089);
and UO_2712 (O_2712,N_48484,N_49316);
and UO_2713 (O_2713,N_49263,N_48335);
nand UO_2714 (O_2714,N_49121,N_48295);
or UO_2715 (O_2715,N_48754,N_48975);
nand UO_2716 (O_2716,N_49360,N_48441);
nor UO_2717 (O_2717,N_49007,N_48669);
nor UO_2718 (O_2718,N_49677,N_49024);
nor UO_2719 (O_2719,N_47566,N_48072);
nor UO_2720 (O_2720,N_47855,N_48123);
xnor UO_2721 (O_2721,N_48001,N_49715);
nor UO_2722 (O_2722,N_48527,N_49407);
xor UO_2723 (O_2723,N_48430,N_48377);
or UO_2724 (O_2724,N_49161,N_47740);
nand UO_2725 (O_2725,N_48618,N_48177);
xnor UO_2726 (O_2726,N_47888,N_49977);
nand UO_2727 (O_2727,N_48599,N_47751);
or UO_2728 (O_2728,N_49678,N_49265);
or UO_2729 (O_2729,N_49909,N_48924);
or UO_2730 (O_2730,N_48144,N_49007);
nor UO_2731 (O_2731,N_48336,N_47606);
xnor UO_2732 (O_2732,N_48972,N_48566);
and UO_2733 (O_2733,N_49830,N_48652);
and UO_2734 (O_2734,N_48546,N_49498);
nand UO_2735 (O_2735,N_48356,N_49400);
and UO_2736 (O_2736,N_49494,N_49889);
nand UO_2737 (O_2737,N_49007,N_48026);
or UO_2738 (O_2738,N_48683,N_49037);
or UO_2739 (O_2739,N_49082,N_49439);
and UO_2740 (O_2740,N_49587,N_49039);
xor UO_2741 (O_2741,N_47724,N_48701);
nand UO_2742 (O_2742,N_48374,N_48338);
and UO_2743 (O_2743,N_48025,N_48933);
nor UO_2744 (O_2744,N_49391,N_47876);
nor UO_2745 (O_2745,N_49050,N_48412);
or UO_2746 (O_2746,N_49649,N_48951);
and UO_2747 (O_2747,N_47557,N_48721);
or UO_2748 (O_2748,N_47515,N_48033);
nand UO_2749 (O_2749,N_48989,N_48804);
xor UO_2750 (O_2750,N_49402,N_48452);
nor UO_2751 (O_2751,N_48938,N_48078);
or UO_2752 (O_2752,N_49412,N_48562);
nor UO_2753 (O_2753,N_49903,N_48564);
or UO_2754 (O_2754,N_48595,N_49310);
nor UO_2755 (O_2755,N_47737,N_49485);
nand UO_2756 (O_2756,N_49845,N_49661);
nand UO_2757 (O_2757,N_48549,N_48297);
nand UO_2758 (O_2758,N_49565,N_48270);
and UO_2759 (O_2759,N_49676,N_49852);
nand UO_2760 (O_2760,N_49446,N_47765);
nand UO_2761 (O_2761,N_47703,N_49185);
nor UO_2762 (O_2762,N_49651,N_49220);
and UO_2763 (O_2763,N_49198,N_47554);
nand UO_2764 (O_2764,N_47987,N_49711);
nor UO_2765 (O_2765,N_48512,N_49466);
and UO_2766 (O_2766,N_47782,N_47901);
and UO_2767 (O_2767,N_49859,N_48314);
or UO_2768 (O_2768,N_48705,N_48105);
nor UO_2769 (O_2769,N_47847,N_48777);
or UO_2770 (O_2770,N_48543,N_49155);
and UO_2771 (O_2771,N_47709,N_47859);
and UO_2772 (O_2772,N_48728,N_49343);
or UO_2773 (O_2773,N_48060,N_47922);
nand UO_2774 (O_2774,N_47615,N_49781);
nor UO_2775 (O_2775,N_48960,N_48470);
and UO_2776 (O_2776,N_49827,N_49880);
nor UO_2777 (O_2777,N_48718,N_49214);
nor UO_2778 (O_2778,N_48312,N_48131);
xnor UO_2779 (O_2779,N_47591,N_49896);
or UO_2780 (O_2780,N_47769,N_48389);
nand UO_2781 (O_2781,N_48058,N_48958);
nor UO_2782 (O_2782,N_49083,N_48020);
or UO_2783 (O_2783,N_48004,N_47998);
nand UO_2784 (O_2784,N_49429,N_48693);
nand UO_2785 (O_2785,N_49119,N_47867);
and UO_2786 (O_2786,N_48133,N_48499);
xor UO_2787 (O_2787,N_48852,N_47700);
or UO_2788 (O_2788,N_47561,N_47615);
or UO_2789 (O_2789,N_47629,N_49312);
nor UO_2790 (O_2790,N_48821,N_47505);
xnor UO_2791 (O_2791,N_49090,N_49369);
and UO_2792 (O_2792,N_47507,N_49986);
or UO_2793 (O_2793,N_48830,N_48249);
nor UO_2794 (O_2794,N_48945,N_47951);
and UO_2795 (O_2795,N_49864,N_49326);
nor UO_2796 (O_2796,N_48927,N_49550);
nor UO_2797 (O_2797,N_48417,N_47896);
xnor UO_2798 (O_2798,N_47658,N_48591);
nand UO_2799 (O_2799,N_48162,N_48648);
or UO_2800 (O_2800,N_48700,N_49084);
or UO_2801 (O_2801,N_49554,N_48270);
xnor UO_2802 (O_2802,N_48252,N_47813);
nand UO_2803 (O_2803,N_49155,N_49630);
or UO_2804 (O_2804,N_48380,N_48679);
xor UO_2805 (O_2805,N_49795,N_47954);
nor UO_2806 (O_2806,N_49733,N_48576);
nor UO_2807 (O_2807,N_49389,N_49436);
nor UO_2808 (O_2808,N_49302,N_48498);
and UO_2809 (O_2809,N_47877,N_47810);
and UO_2810 (O_2810,N_48812,N_49579);
nand UO_2811 (O_2811,N_48191,N_49501);
or UO_2812 (O_2812,N_49174,N_47541);
and UO_2813 (O_2813,N_48965,N_49438);
nand UO_2814 (O_2814,N_47997,N_47872);
xnor UO_2815 (O_2815,N_49212,N_48684);
and UO_2816 (O_2816,N_48796,N_48869);
nor UO_2817 (O_2817,N_48759,N_48908);
and UO_2818 (O_2818,N_48685,N_49853);
nand UO_2819 (O_2819,N_47941,N_47760);
xnor UO_2820 (O_2820,N_47797,N_47718);
nand UO_2821 (O_2821,N_48434,N_47600);
and UO_2822 (O_2822,N_48216,N_49700);
nand UO_2823 (O_2823,N_49478,N_49045);
and UO_2824 (O_2824,N_48835,N_49228);
or UO_2825 (O_2825,N_48599,N_48156);
nor UO_2826 (O_2826,N_49664,N_48360);
nor UO_2827 (O_2827,N_49712,N_48058);
or UO_2828 (O_2828,N_49487,N_48085);
and UO_2829 (O_2829,N_49505,N_49591);
or UO_2830 (O_2830,N_49977,N_49120);
xor UO_2831 (O_2831,N_47518,N_47976);
nor UO_2832 (O_2832,N_48143,N_49539);
or UO_2833 (O_2833,N_49465,N_49722);
or UO_2834 (O_2834,N_47658,N_49140);
nand UO_2835 (O_2835,N_48578,N_48516);
xor UO_2836 (O_2836,N_47997,N_48956);
nor UO_2837 (O_2837,N_48001,N_49935);
xnor UO_2838 (O_2838,N_48307,N_48395);
xnor UO_2839 (O_2839,N_48117,N_49427);
nor UO_2840 (O_2840,N_48109,N_49182);
nand UO_2841 (O_2841,N_48317,N_48115);
nand UO_2842 (O_2842,N_49548,N_47886);
xor UO_2843 (O_2843,N_47929,N_49967);
xnor UO_2844 (O_2844,N_47901,N_49638);
xnor UO_2845 (O_2845,N_49255,N_49485);
nand UO_2846 (O_2846,N_47874,N_49538);
or UO_2847 (O_2847,N_48967,N_48990);
nor UO_2848 (O_2848,N_49373,N_48849);
and UO_2849 (O_2849,N_47748,N_48211);
nand UO_2850 (O_2850,N_48828,N_47650);
or UO_2851 (O_2851,N_47718,N_48555);
nand UO_2852 (O_2852,N_49083,N_47538);
or UO_2853 (O_2853,N_48980,N_47655);
xor UO_2854 (O_2854,N_48327,N_47803);
xnor UO_2855 (O_2855,N_49554,N_47843);
xor UO_2856 (O_2856,N_47940,N_48912);
nand UO_2857 (O_2857,N_48014,N_49413);
or UO_2858 (O_2858,N_47925,N_48436);
or UO_2859 (O_2859,N_49807,N_48354);
nor UO_2860 (O_2860,N_49695,N_47991);
nand UO_2861 (O_2861,N_48139,N_47706);
and UO_2862 (O_2862,N_47772,N_48906);
nand UO_2863 (O_2863,N_47611,N_47906);
xor UO_2864 (O_2864,N_49308,N_49129);
nand UO_2865 (O_2865,N_49812,N_49336);
and UO_2866 (O_2866,N_48328,N_49108);
or UO_2867 (O_2867,N_49968,N_49826);
and UO_2868 (O_2868,N_49435,N_49237);
or UO_2869 (O_2869,N_49054,N_47725);
nand UO_2870 (O_2870,N_49914,N_49495);
xnor UO_2871 (O_2871,N_49956,N_48132);
or UO_2872 (O_2872,N_48219,N_49342);
or UO_2873 (O_2873,N_49020,N_48945);
nand UO_2874 (O_2874,N_47721,N_49168);
nor UO_2875 (O_2875,N_47630,N_48186);
or UO_2876 (O_2876,N_48907,N_49792);
nor UO_2877 (O_2877,N_47550,N_48102);
or UO_2878 (O_2878,N_47917,N_48428);
or UO_2879 (O_2879,N_49440,N_49098);
or UO_2880 (O_2880,N_49247,N_48317);
nor UO_2881 (O_2881,N_47915,N_48121);
or UO_2882 (O_2882,N_48219,N_49318);
and UO_2883 (O_2883,N_49210,N_47762);
nand UO_2884 (O_2884,N_48721,N_47975);
and UO_2885 (O_2885,N_49373,N_48138);
or UO_2886 (O_2886,N_49740,N_48521);
nor UO_2887 (O_2887,N_48271,N_47992);
xnor UO_2888 (O_2888,N_49039,N_48250);
nand UO_2889 (O_2889,N_48619,N_48999);
nor UO_2890 (O_2890,N_49082,N_48487);
or UO_2891 (O_2891,N_47550,N_47839);
nor UO_2892 (O_2892,N_48317,N_48728);
xnor UO_2893 (O_2893,N_49755,N_48126);
xor UO_2894 (O_2894,N_48341,N_49222);
and UO_2895 (O_2895,N_47637,N_47630);
xnor UO_2896 (O_2896,N_48891,N_49487);
and UO_2897 (O_2897,N_49854,N_49316);
or UO_2898 (O_2898,N_47771,N_49779);
and UO_2899 (O_2899,N_49358,N_47503);
xnor UO_2900 (O_2900,N_49153,N_48433);
and UO_2901 (O_2901,N_48987,N_48596);
and UO_2902 (O_2902,N_49924,N_48305);
xnor UO_2903 (O_2903,N_48148,N_48788);
and UO_2904 (O_2904,N_47763,N_48290);
nand UO_2905 (O_2905,N_48243,N_49988);
xor UO_2906 (O_2906,N_49468,N_48215);
nand UO_2907 (O_2907,N_49807,N_48306);
or UO_2908 (O_2908,N_49789,N_49833);
or UO_2909 (O_2909,N_47629,N_48297);
nor UO_2910 (O_2910,N_47506,N_48320);
or UO_2911 (O_2911,N_47809,N_49636);
nor UO_2912 (O_2912,N_49033,N_48724);
and UO_2913 (O_2913,N_48826,N_49918);
nor UO_2914 (O_2914,N_49116,N_47663);
or UO_2915 (O_2915,N_48002,N_49003);
or UO_2916 (O_2916,N_49864,N_49157);
or UO_2917 (O_2917,N_47910,N_48849);
nor UO_2918 (O_2918,N_49761,N_49362);
nand UO_2919 (O_2919,N_49727,N_47751);
and UO_2920 (O_2920,N_49919,N_48046);
or UO_2921 (O_2921,N_47757,N_49903);
nor UO_2922 (O_2922,N_48620,N_49228);
nor UO_2923 (O_2923,N_48476,N_48165);
nor UO_2924 (O_2924,N_49382,N_49402);
or UO_2925 (O_2925,N_47652,N_48406);
and UO_2926 (O_2926,N_49582,N_47912);
or UO_2927 (O_2927,N_49520,N_49543);
xnor UO_2928 (O_2928,N_47874,N_47611);
xor UO_2929 (O_2929,N_49297,N_49793);
or UO_2930 (O_2930,N_48254,N_48153);
nor UO_2931 (O_2931,N_49418,N_48589);
xnor UO_2932 (O_2932,N_48531,N_49932);
and UO_2933 (O_2933,N_48814,N_48927);
nor UO_2934 (O_2934,N_49781,N_48327);
and UO_2935 (O_2935,N_49093,N_49835);
and UO_2936 (O_2936,N_49706,N_48575);
nand UO_2937 (O_2937,N_49707,N_47992);
nor UO_2938 (O_2938,N_49447,N_49705);
nand UO_2939 (O_2939,N_47806,N_48366);
and UO_2940 (O_2940,N_49198,N_47775);
or UO_2941 (O_2941,N_47549,N_48370);
and UO_2942 (O_2942,N_48500,N_48270);
nand UO_2943 (O_2943,N_48583,N_48902);
and UO_2944 (O_2944,N_49189,N_48068);
and UO_2945 (O_2945,N_49594,N_48457);
or UO_2946 (O_2946,N_48294,N_49759);
or UO_2947 (O_2947,N_49758,N_49286);
or UO_2948 (O_2948,N_49398,N_48617);
xnor UO_2949 (O_2949,N_48963,N_48896);
xor UO_2950 (O_2950,N_49163,N_49638);
or UO_2951 (O_2951,N_48669,N_48530);
xor UO_2952 (O_2952,N_48450,N_49815);
nand UO_2953 (O_2953,N_48966,N_47970);
and UO_2954 (O_2954,N_49765,N_47618);
nand UO_2955 (O_2955,N_49753,N_49938);
nand UO_2956 (O_2956,N_47825,N_47535);
nor UO_2957 (O_2957,N_47741,N_49732);
or UO_2958 (O_2958,N_48284,N_49104);
and UO_2959 (O_2959,N_48007,N_49145);
nor UO_2960 (O_2960,N_48267,N_47898);
nor UO_2961 (O_2961,N_48600,N_47924);
nor UO_2962 (O_2962,N_49826,N_49755);
or UO_2963 (O_2963,N_48913,N_47791);
and UO_2964 (O_2964,N_48396,N_47986);
nor UO_2965 (O_2965,N_47916,N_48758);
nor UO_2966 (O_2966,N_49027,N_47996);
nand UO_2967 (O_2967,N_49492,N_49519);
xnor UO_2968 (O_2968,N_49626,N_49184);
nand UO_2969 (O_2969,N_49174,N_47603);
xor UO_2970 (O_2970,N_49308,N_49577);
or UO_2971 (O_2971,N_49402,N_48709);
or UO_2972 (O_2972,N_47723,N_48687);
or UO_2973 (O_2973,N_47808,N_49155);
and UO_2974 (O_2974,N_47686,N_49260);
nand UO_2975 (O_2975,N_48669,N_47640);
and UO_2976 (O_2976,N_48686,N_49409);
and UO_2977 (O_2977,N_48032,N_47971);
and UO_2978 (O_2978,N_49103,N_48715);
nand UO_2979 (O_2979,N_48649,N_48931);
xor UO_2980 (O_2980,N_48645,N_48794);
nand UO_2981 (O_2981,N_47925,N_49664);
nor UO_2982 (O_2982,N_49608,N_48476);
nor UO_2983 (O_2983,N_47770,N_49177);
nor UO_2984 (O_2984,N_48338,N_47909);
and UO_2985 (O_2985,N_47687,N_49340);
and UO_2986 (O_2986,N_49897,N_48403);
nor UO_2987 (O_2987,N_49084,N_49827);
nor UO_2988 (O_2988,N_48020,N_49964);
or UO_2989 (O_2989,N_49076,N_48283);
xor UO_2990 (O_2990,N_48171,N_48662);
nand UO_2991 (O_2991,N_49941,N_48221);
or UO_2992 (O_2992,N_48880,N_49275);
nor UO_2993 (O_2993,N_49176,N_48962);
and UO_2994 (O_2994,N_48879,N_48708);
and UO_2995 (O_2995,N_48655,N_48868);
and UO_2996 (O_2996,N_49396,N_47880);
nor UO_2997 (O_2997,N_49518,N_48520);
and UO_2998 (O_2998,N_49549,N_47819);
xor UO_2999 (O_2999,N_47865,N_47650);
and UO_3000 (O_3000,N_48002,N_48776);
nor UO_3001 (O_3001,N_49879,N_48852);
or UO_3002 (O_3002,N_49829,N_49071);
nand UO_3003 (O_3003,N_49862,N_49295);
nand UO_3004 (O_3004,N_47684,N_49290);
and UO_3005 (O_3005,N_49882,N_47935);
nor UO_3006 (O_3006,N_48426,N_48783);
or UO_3007 (O_3007,N_48896,N_47633);
nor UO_3008 (O_3008,N_49170,N_48673);
nor UO_3009 (O_3009,N_49222,N_47539);
nand UO_3010 (O_3010,N_49075,N_49303);
and UO_3011 (O_3011,N_49811,N_47525);
or UO_3012 (O_3012,N_47625,N_49402);
and UO_3013 (O_3013,N_47701,N_49724);
and UO_3014 (O_3014,N_48474,N_49287);
or UO_3015 (O_3015,N_48547,N_49851);
nor UO_3016 (O_3016,N_49189,N_49112);
nor UO_3017 (O_3017,N_47520,N_49213);
xnor UO_3018 (O_3018,N_49010,N_47924);
nand UO_3019 (O_3019,N_48203,N_48749);
nor UO_3020 (O_3020,N_48889,N_47555);
or UO_3021 (O_3021,N_49773,N_49764);
nor UO_3022 (O_3022,N_48810,N_48248);
nor UO_3023 (O_3023,N_47900,N_48725);
nand UO_3024 (O_3024,N_47557,N_48802);
and UO_3025 (O_3025,N_48061,N_49866);
xor UO_3026 (O_3026,N_47821,N_47844);
xnor UO_3027 (O_3027,N_49901,N_48449);
and UO_3028 (O_3028,N_49482,N_47737);
nor UO_3029 (O_3029,N_49758,N_49228);
xnor UO_3030 (O_3030,N_49325,N_49428);
or UO_3031 (O_3031,N_49557,N_49167);
nand UO_3032 (O_3032,N_49951,N_49677);
nand UO_3033 (O_3033,N_47612,N_48696);
xnor UO_3034 (O_3034,N_48252,N_48470);
xnor UO_3035 (O_3035,N_49124,N_47998);
nor UO_3036 (O_3036,N_49445,N_48079);
xnor UO_3037 (O_3037,N_49553,N_49984);
or UO_3038 (O_3038,N_48570,N_48059);
and UO_3039 (O_3039,N_48180,N_48309);
nor UO_3040 (O_3040,N_48032,N_48319);
xnor UO_3041 (O_3041,N_49239,N_48201);
nand UO_3042 (O_3042,N_48599,N_48619);
or UO_3043 (O_3043,N_48802,N_47798);
nor UO_3044 (O_3044,N_48430,N_48684);
nor UO_3045 (O_3045,N_49292,N_48950);
or UO_3046 (O_3046,N_47797,N_49406);
nand UO_3047 (O_3047,N_49159,N_48277);
nand UO_3048 (O_3048,N_49569,N_48673);
xnor UO_3049 (O_3049,N_48478,N_48889);
xor UO_3050 (O_3050,N_49604,N_48016);
xor UO_3051 (O_3051,N_49285,N_48056);
and UO_3052 (O_3052,N_48834,N_48674);
nand UO_3053 (O_3053,N_47799,N_48439);
nand UO_3054 (O_3054,N_47942,N_48750);
nor UO_3055 (O_3055,N_47932,N_49069);
or UO_3056 (O_3056,N_49383,N_48246);
and UO_3057 (O_3057,N_48328,N_48198);
and UO_3058 (O_3058,N_49119,N_49937);
or UO_3059 (O_3059,N_48609,N_48618);
nor UO_3060 (O_3060,N_47511,N_49494);
or UO_3061 (O_3061,N_48536,N_49674);
nor UO_3062 (O_3062,N_47964,N_49863);
nor UO_3063 (O_3063,N_49969,N_49264);
and UO_3064 (O_3064,N_49928,N_49288);
nor UO_3065 (O_3065,N_49672,N_48157);
nand UO_3066 (O_3066,N_47605,N_49392);
nand UO_3067 (O_3067,N_49471,N_49103);
xor UO_3068 (O_3068,N_48655,N_49367);
nand UO_3069 (O_3069,N_49261,N_48653);
nand UO_3070 (O_3070,N_49791,N_47985);
nor UO_3071 (O_3071,N_47507,N_47597);
and UO_3072 (O_3072,N_49495,N_49150);
nor UO_3073 (O_3073,N_48283,N_49275);
or UO_3074 (O_3074,N_47684,N_49172);
or UO_3075 (O_3075,N_48150,N_49113);
xor UO_3076 (O_3076,N_48232,N_48213);
or UO_3077 (O_3077,N_49799,N_48462);
nor UO_3078 (O_3078,N_48473,N_47643);
or UO_3079 (O_3079,N_49535,N_48484);
xnor UO_3080 (O_3080,N_48229,N_47522);
and UO_3081 (O_3081,N_49706,N_47536);
xnor UO_3082 (O_3082,N_47553,N_48379);
xor UO_3083 (O_3083,N_48245,N_47752);
nor UO_3084 (O_3084,N_47879,N_49931);
xor UO_3085 (O_3085,N_48632,N_48895);
and UO_3086 (O_3086,N_49473,N_48248);
nand UO_3087 (O_3087,N_48600,N_47749);
nor UO_3088 (O_3088,N_49303,N_47643);
xnor UO_3089 (O_3089,N_47580,N_48045);
and UO_3090 (O_3090,N_47652,N_48111);
nand UO_3091 (O_3091,N_49807,N_48856);
nor UO_3092 (O_3092,N_47548,N_48181);
and UO_3093 (O_3093,N_49211,N_47738);
nor UO_3094 (O_3094,N_47889,N_48465);
nor UO_3095 (O_3095,N_49558,N_48545);
nand UO_3096 (O_3096,N_48323,N_49033);
or UO_3097 (O_3097,N_47961,N_48321);
xnor UO_3098 (O_3098,N_49306,N_47504);
or UO_3099 (O_3099,N_49079,N_48243);
nand UO_3100 (O_3100,N_48822,N_49985);
xnor UO_3101 (O_3101,N_48752,N_48121);
and UO_3102 (O_3102,N_49407,N_47705);
and UO_3103 (O_3103,N_47653,N_49777);
nor UO_3104 (O_3104,N_49127,N_49871);
or UO_3105 (O_3105,N_49238,N_49534);
nor UO_3106 (O_3106,N_49923,N_48518);
or UO_3107 (O_3107,N_47905,N_49847);
xnor UO_3108 (O_3108,N_48404,N_48384);
nor UO_3109 (O_3109,N_48955,N_48268);
nor UO_3110 (O_3110,N_48709,N_48328);
or UO_3111 (O_3111,N_49589,N_48545);
nor UO_3112 (O_3112,N_48240,N_48980);
or UO_3113 (O_3113,N_48464,N_47609);
nand UO_3114 (O_3114,N_49454,N_48552);
nor UO_3115 (O_3115,N_49073,N_49346);
nor UO_3116 (O_3116,N_48665,N_47974);
and UO_3117 (O_3117,N_49600,N_48797);
nor UO_3118 (O_3118,N_49756,N_49509);
and UO_3119 (O_3119,N_47752,N_49782);
nor UO_3120 (O_3120,N_48481,N_49240);
nor UO_3121 (O_3121,N_48372,N_47598);
xor UO_3122 (O_3122,N_48015,N_48274);
or UO_3123 (O_3123,N_49189,N_49604);
xnor UO_3124 (O_3124,N_48806,N_47591);
xor UO_3125 (O_3125,N_49810,N_49029);
and UO_3126 (O_3126,N_48974,N_48942);
and UO_3127 (O_3127,N_48888,N_48833);
and UO_3128 (O_3128,N_48324,N_48364);
nor UO_3129 (O_3129,N_49882,N_47883);
nor UO_3130 (O_3130,N_48837,N_47795);
xor UO_3131 (O_3131,N_48486,N_48010);
xnor UO_3132 (O_3132,N_49697,N_47831);
nand UO_3133 (O_3133,N_48389,N_49192);
xnor UO_3134 (O_3134,N_48351,N_49727);
xor UO_3135 (O_3135,N_49536,N_49904);
and UO_3136 (O_3136,N_49754,N_48688);
and UO_3137 (O_3137,N_48638,N_47525);
nor UO_3138 (O_3138,N_49210,N_48038);
nand UO_3139 (O_3139,N_49849,N_49384);
xor UO_3140 (O_3140,N_48003,N_47947);
nor UO_3141 (O_3141,N_48114,N_49255);
nand UO_3142 (O_3142,N_49763,N_47950);
nand UO_3143 (O_3143,N_48941,N_49172);
or UO_3144 (O_3144,N_48843,N_49576);
or UO_3145 (O_3145,N_47581,N_49570);
xnor UO_3146 (O_3146,N_49384,N_49098);
or UO_3147 (O_3147,N_49522,N_48406);
nor UO_3148 (O_3148,N_49238,N_49903);
or UO_3149 (O_3149,N_49380,N_48667);
and UO_3150 (O_3150,N_47737,N_49363);
and UO_3151 (O_3151,N_49728,N_49046);
or UO_3152 (O_3152,N_49541,N_48899);
and UO_3153 (O_3153,N_48677,N_48786);
nand UO_3154 (O_3154,N_47828,N_48723);
nand UO_3155 (O_3155,N_49979,N_49186);
nor UO_3156 (O_3156,N_48937,N_49880);
and UO_3157 (O_3157,N_48048,N_48908);
nand UO_3158 (O_3158,N_48378,N_48932);
or UO_3159 (O_3159,N_47804,N_48275);
xor UO_3160 (O_3160,N_49114,N_49568);
and UO_3161 (O_3161,N_48722,N_49930);
and UO_3162 (O_3162,N_49381,N_48521);
and UO_3163 (O_3163,N_49039,N_47517);
nor UO_3164 (O_3164,N_49489,N_49335);
nand UO_3165 (O_3165,N_47998,N_47689);
nor UO_3166 (O_3166,N_48636,N_48163);
and UO_3167 (O_3167,N_49494,N_49759);
nand UO_3168 (O_3168,N_49258,N_49611);
xnor UO_3169 (O_3169,N_47836,N_48508);
or UO_3170 (O_3170,N_49372,N_47734);
and UO_3171 (O_3171,N_48321,N_49739);
nand UO_3172 (O_3172,N_47547,N_47807);
or UO_3173 (O_3173,N_49506,N_47944);
nand UO_3174 (O_3174,N_48390,N_47717);
xnor UO_3175 (O_3175,N_49292,N_49581);
nor UO_3176 (O_3176,N_48273,N_48780);
xnor UO_3177 (O_3177,N_49781,N_49772);
nor UO_3178 (O_3178,N_47679,N_47916);
nand UO_3179 (O_3179,N_47732,N_49341);
nor UO_3180 (O_3180,N_48589,N_48875);
nand UO_3181 (O_3181,N_48437,N_49269);
nand UO_3182 (O_3182,N_47873,N_48972);
and UO_3183 (O_3183,N_48148,N_48155);
nor UO_3184 (O_3184,N_49071,N_48685);
or UO_3185 (O_3185,N_48648,N_49929);
or UO_3186 (O_3186,N_47734,N_49304);
nand UO_3187 (O_3187,N_49588,N_48137);
nor UO_3188 (O_3188,N_48430,N_48286);
or UO_3189 (O_3189,N_47582,N_47939);
xnor UO_3190 (O_3190,N_47544,N_48215);
xnor UO_3191 (O_3191,N_49716,N_48617);
nor UO_3192 (O_3192,N_48717,N_49809);
and UO_3193 (O_3193,N_48097,N_49272);
xor UO_3194 (O_3194,N_47947,N_47566);
xor UO_3195 (O_3195,N_49090,N_47576);
xor UO_3196 (O_3196,N_49110,N_47615);
and UO_3197 (O_3197,N_48054,N_47706);
or UO_3198 (O_3198,N_48936,N_48815);
and UO_3199 (O_3199,N_49361,N_47894);
nor UO_3200 (O_3200,N_48756,N_49359);
and UO_3201 (O_3201,N_47736,N_48847);
nor UO_3202 (O_3202,N_48686,N_49293);
nand UO_3203 (O_3203,N_47989,N_49100);
nor UO_3204 (O_3204,N_48707,N_48027);
or UO_3205 (O_3205,N_49513,N_49304);
xnor UO_3206 (O_3206,N_47743,N_48552);
or UO_3207 (O_3207,N_49932,N_48334);
or UO_3208 (O_3208,N_49379,N_49812);
or UO_3209 (O_3209,N_48492,N_49677);
nor UO_3210 (O_3210,N_48421,N_48616);
or UO_3211 (O_3211,N_49189,N_49206);
xnor UO_3212 (O_3212,N_48302,N_49886);
nor UO_3213 (O_3213,N_48013,N_49605);
xnor UO_3214 (O_3214,N_48860,N_48308);
nand UO_3215 (O_3215,N_47714,N_48171);
nand UO_3216 (O_3216,N_48810,N_48211);
and UO_3217 (O_3217,N_48020,N_47839);
or UO_3218 (O_3218,N_47960,N_47898);
and UO_3219 (O_3219,N_49069,N_49633);
or UO_3220 (O_3220,N_49932,N_48540);
nand UO_3221 (O_3221,N_48233,N_49436);
and UO_3222 (O_3222,N_48239,N_49166);
nor UO_3223 (O_3223,N_47570,N_48761);
and UO_3224 (O_3224,N_49254,N_48583);
or UO_3225 (O_3225,N_48120,N_48723);
nor UO_3226 (O_3226,N_48687,N_48425);
nand UO_3227 (O_3227,N_49741,N_48938);
xnor UO_3228 (O_3228,N_49588,N_48259);
nor UO_3229 (O_3229,N_48775,N_49511);
and UO_3230 (O_3230,N_48486,N_48445);
xnor UO_3231 (O_3231,N_47922,N_49794);
and UO_3232 (O_3232,N_48935,N_49568);
nor UO_3233 (O_3233,N_49463,N_48112);
or UO_3234 (O_3234,N_47915,N_49264);
or UO_3235 (O_3235,N_48138,N_49197);
and UO_3236 (O_3236,N_48901,N_49301);
nand UO_3237 (O_3237,N_47972,N_49517);
nor UO_3238 (O_3238,N_49522,N_49438);
and UO_3239 (O_3239,N_49871,N_49902);
nand UO_3240 (O_3240,N_48530,N_48462);
nor UO_3241 (O_3241,N_47575,N_49884);
xnor UO_3242 (O_3242,N_48886,N_47967);
or UO_3243 (O_3243,N_47813,N_48582);
xnor UO_3244 (O_3244,N_48052,N_47581);
nand UO_3245 (O_3245,N_47967,N_49838);
or UO_3246 (O_3246,N_48556,N_48525);
and UO_3247 (O_3247,N_49884,N_49490);
xor UO_3248 (O_3248,N_47592,N_47554);
nor UO_3249 (O_3249,N_49282,N_49283);
nand UO_3250 (O_3250,N_48136,N_49759);
xnor UO_3251 (O_3251,N_48021,N_49143);
nor UO_3252 (O_3252,N_49328,N_49179);
xnor UO_3253 (O_3253,N_48103,N_49658);
or UO_3254 (O_3254,N_47562,N_49094);
nor UO_3255 (O_3255,N_47723,N_49256);
or UO_3256 (O_3256,N_48984,N_48936);
nand UO_3257 (O_3257,N_49487,N_47994);
xor UO_3258 (O_3258,N_49399,N_49254);
and UO_3259 (O_3259,N_49733,N_48307);
or UO_3260 (O_3260,N_49024,N_48429);
and UO_3261 (O_3261,N_48492,N_48144);
xor UO_3262 (O_3262,N_48396,N_49966);
nor UO_3263 (O_3263,N_47588,N_48582);
nand UO_3264 (O_3264,N_47590,N_48532);
nor UO_3265 (O_3265,N_47996,N_47905);
or UO_3266 (O_3266,N_49400,N_49084);
nand UO_3267 (O_3267,N_48041,N_48919);
nand UO_3268 (O_3268,N_49733,N_48757);
xnor UO_3269 (O_3269,N_48911,N_47957);
or UO_3270 (O_3270,N_48839,N_49602);
nand UO_3271 (O_3271,N_47962,N_48499);
and UO_3272 (O_3272,N_49510,N_48534);
nand UO_3273 (O_3273,N_48777,N_49836);
nand UO_3274 (O_3274,N_48724,N_49621);
and UO_3275 (O_3275,N_48029,N_48773);
xor UO_3276 (O_3276,N_49910,N_47918);
xor UO_3277 (O_3277,N_49091,N_49018);
or UO_3278 (O_3278,N_47923,N_48663);
nor UO_3279 (O_3279,N_49720,N_49650);
and UO_3280 (O_3280,N_48310,N_49278);
and UO_3281 (O_3281,N_48210,N_47506);
nor UO_3282 (O_3282,N_48106,N_47982);
xnor UO_3283 (O_3283,N_48316,N_49450);
nor UO_3284 (O_3284,N_49253,N_48109);
xnor UO_3285 (O_3285,N_48852,N_49918);
nor UO_3286 (O_3286,N_48303,N_49280);
or UO_3287 (O_3287,N_49374,N_49293);
nand UO_3288 (O_3288,N_49991,N_49481);
or UO_3289 (O_3289,N_49919,N_49546);
or UO_3290 (O_3290,N_48088,N_49536);
and UO_3291 (O_3291,N_48115,N_49923);
or UO_3292 (O_3292,N_49316,N_47835);
or UO_3293 (O_3293,N_48178,N_49784);
xor UO_3294 (O_3294,N_49626,N_48773);
xnor UO_3295 (O_3295,N_48355,N_48022);
and UO_3296 (O_3296,N_48496,N_47979);
and UO_3297 (O_3297,N_48346,N_49349);
nand UO_3298 (O_3298,N_47769,N_49778);
xnor UO_3299 (O_3299,N_49058,N_49683);
and UO_3300 (O_3300,N_48674,N_48631);
and UO_3301 (O_3301,N_47966,N_47745);
nand UO_3302 (O_3302,N_47628,N_48455);
nor UO_3303 (O_3303,N_48935,N_48552);
or UO_3304 (O_3304,N_47725,N_48009);
xor UO_3305 (O_3305,N_47968,N_49898);
nand UO_3306 (O_3306,N_49160,N_49061);
xnor UO_3307 (O_3307,N_48413,N_48127);
nor UO_3308 (O_3308,N_49764,N_48543);
and UO_3309 (O_3309,N_49641,N_49218);
and UO_3310 (O_3310,N_48114,N_49688);
nor UO_3311 (O_3311,N_48404,N_49688);
nor UO_3312 (O_3312,N_48002,N_48869);
nor UO_3313 (O_3313,N_48912,N_49878);
nor UO_3314 (O_3314,N_49255,N_47976);
nand UO_3315 (O_3315,N_47693,N_48095);
or UO_3316 (O_3316,N_48060,N_47577);
nand UO_3317 (O_3317,N_48486,N_48659);
or UO_3318 (O_3318,N_48296,N_48456);
or UO_3319 (O_3319,N_48369,N_49957);
and UO_3320 (O_3320,N_49531,N_49217);
nand UO_3321 (O_3321,N_49282,N_49753);
or UO_3322 (O_3322,N_49146,N_47841);
nor UO_3323 (O_3323,N_47673,N_49747);
nand UO_3324 (O_3324,N_48120,N_48354);
and UO_3325 (O_3325,N_49896,N_49979);
nand UO_3326 (O_3326,N_47593,N_48427);
nand UO_3327 (O_3327,N_47808,N_49835);
nor UO_3328 (O_3328,N_49711,N_48366);
nor UO_3329 (O_3329,N_48707,N_49168);
nand UO_3330 (O_3330,N_48072,N_49419);
nand UO_3331 (O_3331,N_48420,N_47515);
and UO_3332 (O_3332,N_47900,N_48261);
and UO_3333 (O_3333,N_48587,N_47506);
nand UO_3334 (O_3334,N_48680,N_47675);
or UO_3335 (O_3335,N_49047,N_49243);
nor UO_3336 (O_3336,N_47741,N_49039);
xnor UO_3337 (O_3337,N_49172,N_48364);
and UO_3338 (O_3338,N_49652,N_47984);
or UO_3339 (O_3339,N_48138,N_48120);
nor UO_3340 (O_3340,N_48840,N_48862);
nor UO_3341 (O_3341,N_47659,N_49643);
nand UO_3342 (O_3342,N_49414,N_49577);
xor UO_3343 (O_3343,N_48969,N_48314);
nand UO_3344 (O_3344,N_49780,N_48462);
xnor UO_3345 (O_3345,N_48368,N_48040);
and UO_3346 (O_3346,N_48956,N_47760);
or UO_3347 (O_3347,N_48623,N_48506);
xor UO_3348 (O_3348,N_47946,N_49254);
and UO_3349 (O_3349,N_49278,N_48137);
nand UO_3350 (O_3350,N_47665,N_47624);
and UO_3351 (O_3351,N_48310,N_47571);
nand UO_3352 (O_3352,N_47896,N_48788);
xnor UO_3353 (O_3353,N_47768,N_48940);
xor UO_3354 (O_3354,N_48087,N_49493);
nor UO_3355 (O_3355,N_49634,N_48880);
nand UO_3356 (O_3356,N_47555,N_48739);
xor UO_3357 (O_3357,N_49303,N_47538);
xnor UO_3358 (O_3358,N_48014,N_49923);
nor UO_3359 (O_3359,N_49230,N_48218);
nor UO_3360 (O_3360,N_49934,N_49444);
or UO_3361 (O_3361,N_48534,N_48724);
and UO_3362 (O_3362,N_49079,N_47641);
nand UO_3363 (O_3363,N_49060,N_49262);
nor UO_3364 (O_3364,N_47714,N_48553);
nor UO_3365 (O_3365,N_48141,N_48449);
or UO_3366 (O_3366,N_49421,N_47712);
nand UO_3367 (O_3367,N_48427,N_47932);
or UO_3368 (O_3368,N_49659,N_47658);
and UO_3369 (O_3369,N_49078,N_49232);
or UO_3370 (O_3370,N_47983,N_49221);
nand UO_3371 (O_3371,N_48642,N_47883);
and UO_3372 (O_3372,N_48864,N_49587);
xnor UO_3373 (O_3373,N_49898,N_49372);
nor UO_3374 (O_3374,N_49809,N_48750);
xnor UO_3375 (O_3375,N_47817,N_49789);
and UO_3376 (O_3376,N_47717,N_48477);
or UO_3377 (O_3377,N_49505,N_49382);
nand UO_3378 (O_3378,N_48530,N_48328);
xnor UO_3379 (O_3379,N_49220,N_47934);
or UO_3380 (O_3380,N_47648,N_49540);
or UO_3381 (O_3381,N_48552,N_49069);
nor UO_3382 (O_3382,N_48487,N_48861);
nor UO_3383 (O_3383,N_47859,N_49627);
or UO_3384 (O_3384,N_47716,N_49300);
nand UO_3385 (O_3385,N_47764,N_49035);
xor UO_3386 (O_3386,N_48859,N_47507);
xor UO_3387 (O_3387,N_48502,N_49041);
nor UO_3388 (O_3388,N_47601,N_48679);
or UO_3389 (O_3389,N_48778,N_47753);
nand UO_3390 (O_3390,N_47594,N_49803);
nor UO_3391 (O_3391,N_49233,N_49277);
nor UO_3392 (O_3392,N_48504,N_49297);
and UO_3393 (O_3393,N_49516,N_48899);
or UO_3394 (O_3394,N_48454,N_47698);
nand UO_3395 (O_3395,N_49320,N_49606);
nor UO_3396 (O_3396,N_48492,N_49112);
and UO_3397 (O_3397,N_48518,N_48351);
or UO_3398 (O_3398,N_49612,N_47908);
or UO_3399 (O_3399,N_48807,N_49976);
nor UO_3400 (O_3400,N_49199,N_49302);
nand UO_3401 (O_3401,N_49913,N_49238);
nor UO_3402 (O_3402,N_49652,N_48721);
and UO_3403 (O_3403,N_49297,N_47639);
and UO_3404 (O_3404,N_49113,N_48593);
nand UO_3405 (O_3405,N_47522,N_48005);
or UO_3406 (O_3406,N_49975,N_48476);
and UO_3407 (O_3407,N_48738,N_47848);
nor UO_3408 (O_3408,N_48472,N_49005);
nand UO_3409 (O_3409,N_48860,N_49245);
or UO_3410 (O_3410,N_49896,N_49702);
nor UO_3411 (O_3411,N_49594,N_47794);
or UO_3412 (O_3412,N_47906,N_47722);
or UO_3413 (O_3413,N_49951,N_49735);
and UO_3414 (O_3414,N_49411,N_48660);
and UO_3415 (O_3415,N_49949,N_48847);
nand UO_3416 (O_3416,N_48923,N_47607);
xnor UO_3417 (O_3417,N_47753,N_48284);
xor UO_3418 (O_3418,N_48618,N_48853);
xnor UO_3419 (O_3419,N_47538,N_48211);
xor UO_3420 (O_3420,N_47565,N_48807);
or UO_3421 (O_3421,N_48068,N_48420);
or UO_3422 (O_3422,N_49805,N_49896);
or UO_3423 (O_3423,N_48142,N_47741);
or UO_3424 (O_3424,N_48382,N_49832);
xor UO_3425 (O_3425,N_48730,N_48820);
nand UO_3426 (O_3426,N_49399,N_49291);
nor UO_3427 (O_3427,N_49904,N_48135);
or UO_3428 (O_3428,N_48825,N_49386);
xor UO_3429 (O_3429,N_48535,N_48151);
xor UO_3430 (O_3430,N_49111,N_48793);
and UO_3431 (O_3431,N_49188,N_49434);
nand UO_3432 (O_3432,N_49944,N_49777);
or UO_3433 (O_3433,N_47894,N_47899);
nand UO_3434 (O_3434,N_47705,N_49905);
nor UO_3435 (O_3435,N_48143,N_49458);
xor UO_3436 (O_3436,N_49200,N_49145);
or UO_3437 (O_3437,N_49894,N_48762);
and UO_3438 (O_3438,N_48542,N_49659);
and UO_3439 (O_3439,N_48054,N_48248);
xor UO_3440 (O_3440,N_47929,N_48914);
nand UO_3441 (O_3441,N_48227,N_49988);
or UO_3442 (O_3442,N_49267,N_49242);
or UO_3443 (O_3443,N_49128,N_48017);
nand UO_3444 (O_3444,N_49548,N_49281);
nor UO_3445 (O_3445,N_49834,N_48134);
or UO_3446 (O_3446,N_47550,N_48326);
nor UO_3447 (O_3447,N_48063,N_47550);
or UO_3448 (O_3448,N_48681,N_49159);
nor UO_3449 (O_3449,N_48536,N_48533);
nand UO_3450 (O_3450,N_49502,N_47533);
nand UO_3451 (O_3451,N_48326,N_48824);
nand UO_3452 (O_3452,N_49624,N_47869);
nand UO_3453 (O_3453,N_48136,N_48592);
nor UO_3454 (O_3454,N_48615,N_49481);
xnor UO_3455 (O_3455,N_48291,N_48993);
nand UO_3456 (O_3456,N_48378,N_49226);
xnor UO_3457 (O_3457,N_49704,N_47790);
xor UO_3458 (O_3458,N_49190,N_48658);
or UO_3459 (O_3459,N_48604,N_48990);
nand UO_3460 (O_3460,N_48555,N_47899);
xnor UO_3461 (O_3461,N_48759,N_48000);
nor UO_3462 (O_3462,N_49318,N_48733);
nor UO_3463 (O_3463,N_49988,N_48591);
nor UO_3464 (O_3464,N_49116,N_48353);
xor UO_3465 (O_3465,N_48102,N_48311);
nand UO_3466 (O_3466,N_48321,N_49232);
or UO_3467 (O_3467,N_48285,N_49395);
xor UO_3468 (O_3468,N_49063,N_49308);
nor UO_3469 (O_3469,N_49837,N_49490);
xnor UO_3470 (O_3470,N_48505,N_48045);
and UO_3471 (O_3471,N_48380,N_47711);
and UO_3472 (O_3472,N_47597,N_49981);
nand UO_3473 (O_3473,N_47859,N_47570);
or UO_3474 (O_3474,N_49708,N_48128);
nor UO_3475 (O_3475,N_48726,N_49909);
and UO_3476 (O_3476,N_48961,N_49348);
and UO_3477 (O_3477,N_49800,N_48815);
nor UO_3478 (O_3478,N_47523,N_48074);
xor UO_3479 (O_3479,N_48165,N_49947);
xor UO_3480 (O_3480,N_49314,N_49557);
and UO_3481 (O_3481,N_48640,N_49865);
and UO_3482 (O_3482,N_48813,N_47627);
nand UO_3483 (O_3483,N_48650,N_49268);
xor UO_3484 (O_3484,N_49677,N_49855);
xnor UO_3485 (O_3485,N_48633,N_47629);
or UO_3486 (O_3486,N_48788,N_49850);
nand UO_3487 (O_3487,N_47534,N_49998);
nand UO_3488 (O_3488,N_48370,N_47564);
nand UO_3489 (O_3489,N_48395,N_47597);
nand UO_3490 (O_3490,N_49243,N_47744);
and UO_3491 (O_3491,N_48967,N_49508);
nor UO_3492 (O_3492,N_48674,N_49604);
nand UO_3493 (O_3493,N_47507,N_47658);
xnor UO_3494 (O_3494,N_49105,N_48648);
nand UO_3495 (O_3495,N_48114,N_49240);
or UO_3496 (O_3496,N_49930,N_49299);
or UO_3497 (O_3497,N_49534,N_48685);
nand UO_3498 (O_3498,N_48458,N_48877);
xnor UO_3499 (O_3499,N_48202,N_49688);
xnor UO_3500 (O_3500,N_48925,N_47720);
xnor UO_3501 (O_3501,N_49514,N_47629);
nand UO_3502 (O_3502,N_48495,N_49946);
or UO_3503 (O_3503,N_48427,N_49704);
and UO_3504 (O_3504,N_49171,N_48459);
and UO_3505 (O_3505,N_48641,N_48851);
xnor UO_3506 (O_3506,N_49850,N_49877);
and UO_3507 (O_3507,N_48382,N_47917);
xnor UO_3508 (O_3508,N_47782,N_48324);
nor UO_3509 (O_3509,N_48479,N_49458);
nor UO_3510 (O_3510,N_48966,N_48325);
or UO_3511 (O_3511,N_48958,N_48029);
nand UO_3512 (O_3512,N_47758,N_48553);
nor UO_3513 (O_3513,N_48915,N_48794);
and UO_3514 (O_3514,N_48067,N_48431);
nor UO_3515 (O_3515,N_47509,N_49010);
nand UO_3516 (O_3516,N_49212,N_48264);
and UO_3517 (O_3517,N_47879,N_48560);
nand UO_3518 (O_3518,N_48302,N_48751);
and UO_3519 (O_3519,N_48564,N_47790);
nand UO_3520 (O_3520,N_49157,N_49066);
xnor UO_3521 (O_3521,N_48190,N_49633);
and UO_3522 (O_3522,N_49391,N_48108);
xor UO_3523 (O_3523,N_49074,N_48283);
xor UO_3524 (O_3524,N_48617,N_47924);
and UO_3525 (O_3525,N_48203,N_48552);
nor UO_3526 (O_3526,N_48903,N_47612);
nand UO_3527 (O_3527,N_48425,N_47821);
nand UO_3528 (O_3528,N_47873,N_49233);
nand UO_3529 (O_3529,N_48774,N_48133);
and UO_3530 (O_3530,N_48503,N_49423);
xnor UO_3531 (O_3531,N_49790,N_49265);
and UO_3532 (O_3532,N_49931,N_47799);
or UO_3533 (O_3533,N_48260,N_49003);
and UO_3534 (O_3534,N_49595,N_49637);
xor UO_3535 (O_3535,N_49308,N_48623);
nand UO_3536 (O_3536,N_47540,N_47538);
xnor UO_3537 (O_3537,N_49624,N_48063);
nor UO_3538 (O_3538,N_48808,N_47727);
and UO_3539 (O_3539,N_48670,N_49791);
or UO_3540 (O_3540,N_49234,N_48045);
xnor UO_3541 (O_3541,N_47582,N_47589);
nand UO_3542 (O_3542,N_49433,N_49500);
xor UO_3543 (O_3543,N_47595,N_49113);
and UO_3544 (O_3544,N_48050,N_49567);
nand UO_3545 (O_3545,N_47981,N_49988);
xnor UO_3546 (O_3546,N_49940,N_47729);
xor UO_3547 (O_3547,N_48678,N_49797);
or UO_3548 (O_3548,N_47890,N_48182);
xnor UO_3549 (O_3549,N_48235,N_48230);
xor UO_3550 (O_3550,N_48534,N_49104);
or UO_3551 (O_3551,N_47650,N_49868);
nor UO_3552 (O_3552,N_49279,N_48862);
nand UO_3553 (O_3553,N_47874,N_47510);
nand UO_3554 (O_3554,N_48464,N_48653);
or UO_3555 (O_3555,N_48281,N_48384);
nor UO_3556 (O_3556,N_49274,N_49102);
nand UO_3557 (O_3557,N_48246,N_48427);
nand UO_3558 (O_3558,N_49745,N_47657);
nand UO_3559 (O_3559,N_49691,N_47602);
or UO_3560 (O_3560,N_49122,N_49812);
or UO_3561 (O_3561,N_49582,N_48243);
and UO_3562 (O_3562,N_49879,N_48096);
or UO_3563 (O_3563,N_49916,N_47781);
nor UO_3564 (O_3564,N_49720,N_48361);
or UO_3565 (O_3565,N_47558,N_49878);
nor UO_3566 (O_3566,N_49154,N_48209);
xor UO_3567 (O_3567,N_47823,N_49363);
nor UO_3568 (O_3568,N_48597,N_48521);
xor UO_3569 (O_3569,N_48988,N_47758);
xor UO_3570 (O_3570,N_48139,N_48458);
and UO_3571 (O_3571,N_48598,N_48003);
xnor UO_3572 (O_3572,N_47773,N_47841);
or UO_3573 (O_3573,N_49263,N_47815);
or UO_3574 (O_3574,N_47866,N_48137);
and UO_3575 (O_3575,N_48532,N_49797);
xnor UO_3576 (O_3576,N_49690,N_48793);
nand UO_3577 (O_3577,N_48239,N_48248);
nand UO_3578 (O_3578,N_49985,N_47679);
nand UO_3579 (O_3579,N_48072,N_49407);
and UO_3580 (O_3580,N_49396,N_47588);
or UO_3581 (O_3581,N_49777,N_49829);
or UO_3582 (O_3582,N_49787,N_48012);
nor UO_3583 (O_3583,N_49842,N_47744);
nand UO_3584 (O_3584,N_48023,N_47848);
nand UO_3585 (O_3585,N_49005,N_49724);
xnor UO_3586 (O_3586,N_49611,N_48180);
xnor UO_3587 (O_3587,N_47535,N_47648);
xor UO_3588 (O_3588,N_48927,N_49925);
nand UO_3589 (O_3589,N_47500,N_47910);
xnor UO_3590 (O_3590,N_49524,N_49685);
or UO_3591 (O_3591,N_48858,N_48228);
nand UO_3592 (O_3592,N_48892,N_48032);
or UO_3593 (O_3593,N_48441,N_49452);
nand UO_3594 (O_3594,N_49517,N_48878);
or UO_3595 (O_3595,N_48686,N_48039);
nand UO_3596 (O_3596,N_48688,N_47655);
and UO_3597 (O_3597,N_48962,N_48344);
and UO_3598 (O_3598,N_48505,N_49940);
and UO_3599 (O_3599,N_49653,N_47646);
or UO_3600 (O_3600,N_49010,N_48644);
or UO_3601 (O_3601,N_48191,N_49105);
nand UO_3602 (O_3602,N_49975,N_49135);
and UO_3603 (O_3603,N_48392,N_47917);
xor UO_3604 (O_3604,N_49225,N_48374);
xnor UO_3605 (O_3605,N_49954,N_49135);
xnor UO_3606 (O_3606,N_49791,N_48395);
nor UO_3607 (O_3607,N_49949,N_48657);
or UO_3608 (O_3608,N_47876,N_49351);
nand UO_3609 (O_3609,N_49923,N_48274);
or UO_3610 (O_3610,N_49513,N_48353);
nor UO_3611 (O_3611,N_49622,N_48830);
xnor UO_3612 (O_3612,N_47834,N_48638);
nor UO_3613 (O_3613,N_48699,N_48909);
xnor UO_3614 (O_3614,N_49685,N_49902);
and UO_3615 (O_3615,N_48608,N_48034);
xor UO_3616 (O_3616,N_49508,N_48485);
xnor UO_3617 (O_3617,N_47519,N_48331);
and UO_3618 (O_3618,N_47901,N_48314);
nor UO_3619 (O_3619,N_48784,N_48045);
nand UO_3620 (O_3620,N_49344,N_48709);
nor UO_3621 (O_3621,N_48658,N_48477);
or UO_3622 (O_3622,N_48019,N_47713);
xnor UO_3623 (O_3623,N_49944,N_48587);
nor UO_3624 (O_3624,N_47678,N_48070);
nor UO_3625 (O_3625,N_47621,N_49914);
nand UO_3626 (O_3626,N_47713,N_49744);
or UO_3627 (O_3627,N_49591,N_48276);
nor UO_3628 (O_3628,N_48234,N_48317);
nor UO_3629 (O_3629,N_48411,N_49303);
and UO_3630 (O_3630,N_48245,N_48096);
or UO_3631 (O_3631,N_48638,N_49267);
or UO_3632 (O_3632,N_48165,N_47720);
or UO_3633 (O_3633,N_49109,N_49692);
nand UO_3634 (O_3634,N_47526,N_47825);
and UO_3635 (O_3635,N_48816,N_49302);
nor UO_3636 (O_3636,N_48973,N_47702);
nor UO_3637 (O_3637,N_47788,N_48142);
and UO_3638 (O_3638,N_49355,N_49356);
and UO_3639 (O_3639,N_49598,N_48259);
xor UO_3640 (O_3640,N_49996,N_48056);
and UO_3641 (O_3641,N_47884,N_48751);
and UO_3642 (O_3642,N_48151,N_49519);
nand UO_3643 (O_3643,N_47583,N_48767);
and UO_3644 (O_3644,N_49009,N_49763);
or UO_3645 (O_3645,N_47631,N_49432);
xor UO_3646 (O_3646,N_48942,N_47929);
and UO_3647 (O_3647,N_47855,N_47826);
xor UO_3648 (O_3648,N_47620,N_48042);
and UO_3649 (O_3649,N_47832,N_47690);
nand UO_3650 (O_3650,N_49180,N_49558);
and UO_3651 (O_3651,N_48460,N_47791);
xnor UO_3652 (O_3652,N_48605,N_49040);
nor UO_3653 (O_3653,N_49808,N_48515);
xor UO_3654 (O_3654,N_49675,N_48953);
nand UO_3655 (O_3655,N_49083,N_48816);
nor UO_3656 (O_3656,N_49959,N_49353);
and UO_3657 (O_3657,N_49989,N_48547);
nor UO_3658 (O_3658,N_48152,N_47792);
nand UO_3659 (O_3659,N_48591,N_49343);
nor UO_3660 (O_3660,N_47927,N_49405);
or UO_3661 (O_3661,N_49374,N_48633);
and UO_3662 (O_3662,N_49382,N_48462);
nand UO_3663 (O_3663,N_48106,N_48945);
xor UO_3664 (O_3664,N_48126,N_48021);
or UO_3665 (O_3665,N_47923,N_47911);
nand UO_3666 (O_3666,N_49582,N_49420);
nand UO_3667 (O_3667,N_48047,N_48197);
or UO_3668 (O_3668,N_47598,N_47693);
and UO_3669 (O_3669,N_49523,N_48598);
and UO_3670 (O_3670,N_49513,N_47587);
xnor UO_3671 (O_3671,N_47650,N_48168);
or UO_3672 (O_3672,N_49647,N_47718);
xor UO_3673 (O_3673,N_49744,N_47564);
xor UO_3674 (O_3674,N_48387,N_49634);
and UO_3675 (O_3675,N_48782,N_48131);
or UO_3676 (O_3676,N_49492,N_48503);
nor UO_3677 (O_3677,N_49436,N_48507);
and UO_3678 (O_3678,N_48730,N_48983);
nand UO_3679 (O_3679,N_48522,N_48228);
xnor UO_3680 (O_3680,N_47760,N_49187);
or UO_3681 (O_3681,N_49657,N_48561);
nand UO_3682 (O_3682,N_49455,N_49501);
xnor UO_3683 (O_3683,N_48586,N_48852);
nor UO_3684 (O_3684,N_48922,N_48251);
xnor UO_3685 (O_3685,N_49588,N_47511);
nand UO_3686 (O_3686,N_48337,N_49347);
or UO_3687 (O_3687,N_48202,N_48422);
or UO_3688 (O_3688,N_49617,N_48576);
or UO_3689 (O_3689,N_48267,N_48978);
and UO_3690 (O_3690,N_49454,N_48389);
xor UO_3691 (O_3691,N_49129,N_49564);
xnor UO_3692 (O_3692,N_47834,N_48640);
and UO_3693 (O_3693,N_47721,N_48856);
and UO_3694 (O_3694,N_47751,N_49848);
or UO_3695 (O_3695,N_47529,N_49978);
nor UO_3696 (O_3696,N_49941,N_48739);
or UO_3697 (O_3697,N_47613,N_48128);
xnor UO_3698 (O_3698,N_48444,N_49768);
xor UO_3699 (O_3699,N_48492,N_48374);
or UO_3700 (O_3700,N_49174,N_49701);
xor UO_3701 (O_3701,N_47619,N_48143);
and UO_3702 (O_3702,N_49962,N_49508);
or UO_3703 (O_3703,N_49964,N_49591);
and UO_3704 (O_3704,N_48324,N_48813);
or UO_3705 (O_3705,N_47504,N_47676);
xor UO_3706 (O_3706,N_47935,N_49638);
and UO_3707 (O_3707,N_49428,N_49840);
nor UO_3708 (O_3708,N_48311,N_48332);
and UO_3709 (O_3709,N_49587,N_47929);
xor UO_3710 (O_3710,N_47668,N_48086);
and UO_3711 (O_3711,N_49401,N_47958);
nor UO_3712 (O_3712,N_47821,N_48756);
xor UO_3713 (O_3713,N_47545,N_48150);
nor UO_3714 (O_3714,N_48868,N_47752);
and UO_3715 (O_3715,N_48283,N_49502);
or UO_3716 (O_3716,N_48941,N_49853);
and UO_3717 (O_3717,N_49768,N_47696);
and UO_3718 (O_3718,N_48521,N_49806);
nand UO_3719 (O_3719,N_48830,N_48514);
and UO_3720 (O_3720,N_47979,N_49091);
nor UO_3721 (O_3721,N_48380,N_49467);
and UO_3722 (O_3722,N_49764,N_49110);
xnor UO_3723 (O_3723,N_49087,N_49682);
and UO_3724 (O_3724,N_48589,N_49504);
and UO_3725 (O_3725,N_48861,N_49176);
and UO_3726 (O_3726,N_49629,N_49190);
nand UO_3727 (O_3727,N_49420,N_47784);
and UO_3728 (O_3728,N_48463,N_49116);
xor UO_3729 (O_3729,N_49274,N_48887);
xnor UO_3730 (O_3730,N_48470,N_48043);
nand UO_3731 (O_3731,N_49489,N_48024);
nand UO_3732 (O_3732,N_48203,N_48862);
xor UO_3733 (O_3733,N_48274,N_49246);
and UO_3734 (O_3734,N_48900,N_49021);
nand UO_3735 (O_3735,N_48272,N_49836);
and UO_3736 (O_3736,N_48458,N_47535);
or UO_3737 (O_3737,N_47590,N_47599);
or UO_3738 (O_3738,N_48374,N_47573);
nor UO_3739 (O_3739,N_48598,N_49336);
nand UO_3740 (O_3740,N_48161,N_48833);
nand UO_3741 (O_3741,N_48095,N_48493);
xor UO_3742 (O_3742,N_47928,N_47877);
nand UO_3743 (O_3743,N_48349,N_48292);
and UO_3744 (O_3744,N_49648,N_49195);
and UO_3745 (O_3745,N_48889,N_49743);
and UO_3746 (O_3746,N_49127,N_49140);
and UO_3747 (O_3747,N_47502,N_49617);
or UO_3748 (O_3748,N_49794,N_49126);
or UO_3749 (O_3749,N_49520,N_49432);
nand UO_3750 (O_3750,N_49754,N_48504);
and UO_3751 (O_3751,N_47658,N_47601);
or UO_3752 (O_3752,N_49421,N_48745);
and UO_3753 (O_3753,N_49736,N_48335);
nand UO_3754 (O_3754,N_48426,N_49252);
nor UO_3755 (O_3755,N_47607,N_47896);
or UO_3756 (O_3756,N_48237,N_48464);
xor UO_3757 (O_3757,N_48905,N_48348);
or UO_3758 (O_3758,N_49049,N_48546);
and UO_3759 (O_3759,N_49948,N_48071);
nand UO_3760 (O_3760,N_48085,N_49712);
xnor UO_3761 (O_3761,N_47840,N_48662);
nand UO_3762 (O_3762,N_49688,N_47774);
nor UO_3763 (O_3763,N_48005,N_49200);
xor UO_3764 (O_3764,N_48827,N_48124);
and UO_3765 (O_3765,N_49224,N_49569);
xnor UO_3766 (O_3766,N_48601,N_47979);
or UO_3767 (O_3767,N_48090,N_49942);
nor UO_3768 (O_3768,N_49179,N_49798);
nor UO_3769 (O_3769,N_49442,N_48228);
and UO_3770 (O_3770,N_49934,N_47760);
xnor UO_3771 (O_3771,N_49775,N_48187);
and UO_3772 (O_3772,N_49797,N_48381);
and UO_3773 (O_3773,N_47781,N_48023);
nand UO_3774 (O_3774,N_49092,N_49435);
xnor UO_3775 (O_3775,N_48174,N_49521);
nand UO_3776 (O_3776,N_49678,N_47638);
and UO_3777 (O_3777,N_48335,N_48963);
or UO_3778 (O_3778,N_47778,N_47803);
xor UO_3779 (O_3779,N_48351,N_48345);
xor UO_3780 (O_3780,N_49722,N_47828);
nand UO_3781 (O_3781,N_48035,N_49786);
nor UO_3782 (O_3782,N_47840,N_48335);
or UO_3783 (O_3783,N_48143,N_48215);
and UO_3784 (O_3784,N_48942,N_47761);
nor UO_3785 (O_3785,N_49551,N_47675);
or UO_3786 (O_3786,N_49193,N_48298);
nor UO_3787 (O_3787,N_48985,N_48707);
xor UO_3788 (O_3788,N_49892,N_49444);
or UO_3789 (O_3789,N_48141,N_48925);
nor UO_3790 (O_3790,N_48426,N_48613);
or UO_3791 (O_3791,N_48614,N_49630);
nor UO_3792 (O_3792,N_49257,N_48586);
and UO_3793 (O_3793,N_47740,N_47844);
nor UO_3794 (O_3794,N_49427,N_47882);
or UO_3795 (O_3795,N_47825,N_47785);
nor UO_3796 (O_3796,N_49845,N_48723);
or UO_3797 (O_3797,N_47804,N_48400);
nand UO_3798 (O_3798,N_48916,N_47784);
and UO_3799 (O_3799,N_47770,N_47564);
xor UO_3800 (O_3800,N_47961,N_48111);
nor UO_3801 (O_3801,N_48977,N_47741);
nand UO_3802 (O_3802,N_47770,N_48540);
and UO_3803 (O_3803,N_47722,N_48858);
and UO_3804 (O_3804,N_47550,N_47726);
nor UO_3805 (O_3805,N_49678,N_49563);
and UO_3806 (O_3806,N_49714,N_47987);
xor UO_3807 (O_3807,N_48284,N_47987);
or UO_3808 (O_3808,N_49868,N_48488);
or UO_3809 (O_3809,N_49113,N_48260);
or UO_3810 (O_3810,N_47976,N_47741);
xnor UO_3811 (O_3811,N_49225,N_49584);
xor UO_3812 (O_3812,N_49079,N_49950);
or UO_3813 (O_3813,N_48014,N_49202);
xnor UO_3814 (O_3814,N_49809,N_48253);
nand UO_3815 (O_3815,N_47981,N_48507);
nand UO_3816 (O_3816,N_48736,N_49923);
xnor UO_3817 (O_3817,N_49134,N_49669);
xnor UO_3818 (O_3818,N_47619,N_48557);
xnor UO_3819 (O_3819,N_48883,N_49398);
xor UO_3820 (O_3820,N_48767,N_48695);
or UO_3821 (O_3821,N_48583,N_47856);
nor UO_3822 (O_3822,N_48439,N_48918);
xor UO_3823 (O_3823,N_48378,N_47637);
and UO_3824 (O_3824,N_49095,N_47589);
xor UO_3825 (O_3825,N_48079,N_49492);
nor UO_3826 (O_3826,N_49703,N_49680);
nor UO_3827 (O_3827,N_48758,N_49655);
nand UO_3828 (O_3828,N_48930,N_48616);
nand UO_3829 (O_3829,N_48364,N_49331);
nand UO_3830 (O_3830,N_49415,N_48274);
nor UO_3831 (O_3831,N_48609,N_48777);
nand UO_3832 (O_3832,N_48277,N_47763);
or UO_3833 (O_3833,N_48100,N_49389);
nand UO_3834 (O_3834,N_49945,N_49852);
xor UO_3835 (O_3835,N_47944,N_49979);
and UO_3836 (O_3836,N_49850,N_47656);
or UO_3837 (O_3837,N_49608,N_48815);
xor UO_3838 (O_3838,N_47932,N_49003);
xor UO_3839 (O_3839,N_48284,N_48077);
or UO_3840 (O_3840,N_49256,N_47844);
nand UO_3841 (O_3841,N_48009,N_48580);
or UO_3842 (O_3842,N_48117,N_48599);
and UO_3843 (O_3843,N_49013,N_47561);
nor UO_3844 (O_3844,N_49817,N_49775);
and UO_3845 (O_3845,N_48513,N_47837);
nor UO_3846 (O_3846,N_48128,N_49644);
nand UO_3847 (O_3847,N_48068,N_48804);
nor UO_3848 (O_3848,N_47630,N_49391);
or UO_3849 (O_3849,N_49114,N_48069);
or UO_3850 (O_3850,N_47689,N_49606);
or UO_3851 (O_3851,N_49270,N_48611);
and UO_3852 (O_3852,N_49309,N_47870);
and UO_3853 (O_3853,N_48677,N_48942);
and UO_3854 (O_3854,N_48973,N_49835);
and UO_3855 (O_3855,N_47948,N_49652);
and UO_3856 (O_3856,N_48555,N_49152);
nor UO_3857 (O_3857,N_49326,N_48575);
nor UO_3858 (O_3858,N_49246,N_49765);
xnor UO_3859 (O_3859,N_47602,N_48033);
nand UO_3860 (O_3860,N_49755,N_49232);
nor UO_3861 (O_3861,N_48108,N_47842);
and UO_3862 (O_3862,N_49302,N_48745);
or UO_3863 (O_3863,N_48033,N_49840);
and UO_3864 (O_3864,N_49595,N_49891);
xnor UO_3865 (O_3865,N_48210,N_49840);
or UO_3866 (O_3866,N_49216,N_47804);
and UO_3867 (O_3867,N_48798,N_47527);
xnor UO_3868 (O_3868,N_48383,N_49818);
or UO_3869 (O_3869,N_48837,N_47996);
nor UO_3870 (O_3870,N_49282,N_49622);
and UO_3871 (O_3871,N_49367,N_48369);
nor UO_3872 (O_3872,N_49678,N_48523);
and UO_3873 (O_3873,N_49822,N_47644);
and UO_3874 (O_3874,N_49362,N_47701);
nand UO_3875 (O_3875,N_47822,N_48238);
nor UO_3876 (O_3876,N_48568,N_48314);
nand UO_3877 (O_3877,N_48215,N_49590);
nor UO_3878 (O_3878,N_47764,N_47849);
nor UO_3879 (O_3879,N_48766,N_49283);
or UO_3880 (O_3880,N_47809,N_49835);
xnor UO_3881 (O_3881,N_49323,N_49998);
nor UO_3882 (O_3882,N_48116,N_48767);
nor UO_3883 (O_3883,N_48517,N_47996);
or UO_3884 (O_3884,N_47684,N_48601);
nand UO_3885 (O_3885,N_49338,N_49381);
nand UO_3886 (O_3886,N_48862,N_49660);
or UO_3887 (O_3887,N_48865,N_49904);
nand UO_3888 (O_3888,N_49717,N_49611);
xor UO_3889 (O_3889,N_48822,N_48332);
and UO_3890 (O_3890,N_49672,N_49516);
and UO_3891 (O_3891,N_49426,N_49059);
or UO_3892 (O_3892,N_48812,N_47765);
and UO_3893 (O_3893,N_49020,N_48040);
and UO_3894 (O_3894,N_47706,N_48076);
or UO_3895 (O_3895,N_48155,N_49003);
or UO_3896 (O_3896,N_49882,N_47867);
nor UO_3897 (O_3897,N_47918,N_49174);
xnor UO_3898 (O_3898,N_48184,N_47757);
and UO_3899 (O_3899,N_47642,N_48684);
or UO_3900 (O_3900,N_48091,N_48506);
and UO_3901 (O_3901,N_49503,N_49450);
xnor UO_3902 (O_3902,N_49579,N_49326);
and UO_3903 (O_3903,N_49955,N_47923);
nand UO_3904 (O_3904,N_49843,N_49480);
xor UO_3905 (O_3905,N_48698,N_47904);
or UO_3906 (O_3906,N_49342,N_48116);
or UO_3907 (O_3907,N_48494,N_47610);
nor UO_3908 (O_3908,N_47666,N_49281);
and UO_3909 (O_3909,N_49884,N_49351);
nor UO_3910 (O_3910,N_48191,N_49629);
nand UO_3911 (O_3911,N_48292,N_49992);
and UO_3912 (O_3912,N_48381,N_49595);
and UO_3913 (O_3913,N_48564,N_47988);
xnor UO_3914 (O_3914,N_47590,N_47894);
and UO_3915 (O_3915,N_48605,N_47881);
nor UO_3916 (O_3916,N_49882,N_48834);
xor UO_3917 (O_3917,N_48820,N_49516);
or UO_3918 (O_3918,N_48726,N_48724);
and UO_3919 (O_3919,N_49728,N_47731);
or UO_3920 (O_3920,N_48699,N_48728);
and UO_3921 (O_3921,N_49026,N_48593);
nor UO_3922 (O_3922,N_47897,N_49397);
xnor UO_3923 (O_3923,N_49626,N_48226);
or UO_3924 (O_3924,N_47963,N_48009);
nand UO_3925 (O_3925,N_49640,N_49790);
or UO_3926 (O_3926,N_49547,N_48460);
nor UO_3927 (O_3927,N_47849,N_49350);
or UO_3928 (O_3928,N_49759,N_49302);
or UO_3929 (O_3929,N_49929,N_48813);
or UO_3930 (O_3930,N_48139,N_49249);
nand UO_3931 (O_3931,N_49731,N_48048);
nand UO_3932 (O_3932,N_49830,N_49692);
nor UO_3933 (O_3933,N_48438,N_49465);
nor UO_3934 (O_3934,N_48648,N_49425);
xnor UO_3935 (O_3935,N_48966,N_48781);
or UO_3936 (O_3936,N_47527,N_47565);
nand UO_3937 (O_3937,N_49574,N_48283);
nor UO_3938 (O_3938,N_48365,N_47760);
nor UO_3939 (O_3939,N_49100,N_49582);
nand UO_3940 (O_3940,N_48033,N_47987);
xnor UO_3941 (O_3941,N_47810,N_48218);
nand UO_3942 (O_3942,N_48254,N_48211);
and UO_3943 (O_3943,N_49296,N_48648);
xnor UO_3944 (O_3944,N_49418,N_47841);
nor UO_3945 (O_3945,N_48336,N_49973);
nand UO_3946 (O_3946,N_49086,N_48700);
or UO_3947 (O_3947,N_48718,N_49860);
and UO_3948 (O_3948,N_48258,N_48438);
or UO_3949 (O_3949,N_49874,N_48673);
nor UO_3950 (O_3950,N_49755,N_48826);
nand UO_3951 (O_3951,N_48442,N_48356);
and UO_3952 (O_3952,N_49885,N_48630);
nand UO_3953 (O_3953,N_47629,N_49209);
or UO_3954 (O_3954,N_49751,N_48787);
nor UO_3955 (O_3955,N_47718,N_49882);
nor UO_3956 (O_3956,N_48959,N_48197);
xor UO_3957 (O_3957,N_49590,N_49399);
or UO_3958 (O_3958,N_49126,N_49805);
or UO_3959 (O_3959,N_48378,N_49334);
or UO_3960 (O_3960,N_48511,N_48739);
xnor UO_3961 (O_3961,N_48349,N_48975);
xnor UO_3962 (O_3962,N_47505,N_48017);
xor UO_3963 (O_3963,N_47888,N_47908);
or UO_3964 (O_3964,N_47594,N_49953);
nand UO_3965 (O_3965,N_48956,N_47897);
or UO_3966 (O_3966,N_48567,N_49211);
and UO_3967 (O_3967,N_48126,N_49142);
and UO_3968 (O_3968,N_49290,N_48533);
nand UO_3969 (O_3969,N_48564,N_47682);
or UO_3970 (O_3970,N_48271,N_48885);
and UO_3971 (O_3971,N_49348,N_47630);
and UO_3972 (O_3972,N_48054,N_49051);
and UO_3973 (O_3973,N_48028,N_49470);
xor UO_3974 (O_3974,N_48470,N_48779);
nand UO_3975 (O_3975,N_47955,N_48782);
or UO_3976 (O_3976,N_49105,N_47827);
or UO_3977 (O_3977,N_47756,N_48105);
xor UO_3978 (O_3978,N_48993,N_48819);
or UO_3979 (O_3979,N_47992,N_48495);
xor UO_3980 (O_3980,N_49390,N_48986);
xor UO_3981 (O_3981,N_47963,N_49711);
or UO_3982 (O_3982,N_47648,N_47723);
xnor UO_3983 (O_3983,N_48926,N_48533);
or UO_3984 (O_3984,N_49649,N_48636);
or UO_3985 (O_3985,N_48638,N_49237);
xnor UO_3986 (O_3986,N_48128,N_49491);
nor UO_3987 (O_3987,N_49256,N_48975);
or UO_3988 (O_3988,N_48416,N_49040);
or UO_3989 (O_3989,N_49511,N_49108);
and UO_3990 (O_3990,N_49541,N_48038);
nor UO_3991 (O_3991,N_49498,N_49939);
and UO_3992 (O_3992,N_48081,N_47920);
nor UO_3993 (O_3993,N_47557,N_49780);
or UO_3994 (O_3994,N_48823,N_47753);
nor UO_3995 (O_3995,N_49739,N_49615);
or UO_3996 (O_3996,N_49768,N_49639);
nand UO_3997 (O_3997,N_47655,N_48710);
and UO_3998 (O_3998,N_49681,N_49945);
and UO_3999 (O_3999,N_47635,N_47778);
nand UO_4000 (O_4000,N_47806,N_49436);
or UO_4001 (O_4001,N_48183,N_49048);
and UO_4002 (O_4002,N_49508,N_47996);
nor UO_4003 (O_4003,N_48494,N_49752);
xor UO_4004 (O_4004,N_49564,N_49507);
and UO_4005 (O_4005,N_48590,N_48136);
xor UO_4006 (O_4006,N_48218,N_49326);
nand UO_4007 (O_4007,N_49512,N_48661);
nand UO_4008 (O_4008,N_49642,N_49273);
xor UO_4009 (O_4009,N_48695,N_47921);
nand UO_4010 (O_4010,N_49794,N_48522);
or UO_4011 (O_4011,N_48547,N_49086);
and UO_4012 (O_4012,N_49788,N_47849);
nand UO_4013 (O_4013,N_47751,N_49201);
nor UO_4014 (O_4014,N_47693,N_49355);
nor UO_4015 (O_4015,N_49084,N_48505);
and UO_4016 (O_4016,N_49589,N_48653);
nand UO_4017 (O_4017,N_49093,N_47961);
nor UO_4018 (O_4018,N_48314,N_47671);
nor UO_4019 (O_4019,N_48266,N_48515);
or UO_4020 (O_4020,N_49745,N_48851);
xor UO_4021 (O_4021,N_49266,N_48358);
nor UO_4022 (O_4022,N_48174,N_47546);
nand UO_4023 (O_4023,N_49529,N_49741);
or UO_4024 (O_4024,N_48765,N_47873);
and UO_4025 (O_4025,N_49481,N_49288);
or UO_4026 (O_4026,N_48334,N_48903);
nor UO_4027 (O_4027,N_49623,N_47999);
or UO_4028 (O_4028,N_47765,N_47761);
xor UO_4029 (O_4029,N_49338,N_49685);
nor UO_4030 (O_4030,N_48643,N_48432);
and UO_4031 (O_4031,N_48579,N_49393);
nor UO_4032 (O_4032,N_48366,N_48632);
or UO_4033 (O_4033,N_48496,N_47510);
or UO_4034 (O_4034,N_48640,N_48568);
nor UO_4035 (O_4035,N_47525,N_49822);
or UO_4036 (O_4036,N_49285,N_49542);
nand UO_4037 (O_4037,N_49685,N_48754);
and UO_4038 (O_4038,N_49735,N_48401);
nor UO_4039 (O_4039,N_49553,N_47887);
or UO_4040 (O_4040,N_47926,N_49140);
nand UO_4041 (O_4041,N_47678,N_48355);
nor UO_4042 (O_4042,N_49698,N_49817);
and UO_4043 (O_4043,N_49083,N_48450);
nor UO_4044 (O_4044,N_49069,N_49730);
or UO_4045 (O_4045,N_49537,N_48723);
nor UO_4046 (O_4046,N_48232,N_47799);
nand UO_4047 (O_4047,N_48716,N_47631);
nand UO_4048 (O_4048,N_47993,N_48624);
xnor UO_4049 (O_4049,N_48353,N_48428);
xor UO_4050 (O_4050,N_48333,N_49400);
or UO_4051 (O_4051,N_48728,N_47706);
nand UO_4052 (O_4052,N_47736,N_49479);
or UO_4053 (O_4053,N_48078,N_48209);
nand UO_4054 (O_4054,N_47864,N_49568);
and UO_4055 (O_4055,N_48397,N_49348);
nor UO_4056 (O_4056,N_48482,N_49198);
xor UO_4057 (O_4057,N_47570,N_48988);
nand UO_4058 (O_4058,N_48738,N_49501);
xor UO_4059 (O_4059,N_49386,N_48693);
xnor UO_4060 (O_4060,N_47515,N_49627);
nand UO_4061 (O_4061,N_48135,N_49302);
nor UO_4062 (O_4062,N_49017,N_49454);
nand UO_4063 (O_4063,N_48462,N_48380);
nand UO_4064 (O_4064,N_49081,N_47598);
nor UO_4065 (O_4065,N_48592,N_48272);
xor UO_4066 (O_4066,N_48854,N_48210);
or UO_4067 (O_4067,N_49140,N_47837);
and UO_4068 (O_4068,N_48376,N_48035);
and UO_4069 (O_4069,N_47862,N_48421);
nand UO_4070 (O_4070,N_48079,N_47852);
nand UO_4071 (O_4071,N_49752,N_49707);
or UO_4072 (O_4072,N_48853,N_49582);
nor UO_4073 (O_4073,N_49664,N_48890);
xor UO_4074 (O_4074,N_48375,N_48551);
and UO_4075 (O_4075,N_47813,N_48051);
or UO_4076 (O_4076,N_48894,N_48088);
or UO_4077 (O_4077,N_48146,N_49924);
nor UO_4078 (O_4078,N_47996,N_48671);
xnor UO_4079 (O_4079,N_48989,N_47944);
nor UO_4080 (O_4080,N_49608,N_48151);
nor UO_4081 (O_4081,N_48550,N_48245);
or UO_4082 (O_4082,N_49517,N_49377);
or UO_4083 (O_4083,N_49040,N_47965);
or UO_4084 (O_4084,N_47883,N_48577);
xor UO_4085 (O_4085,N_49285,N_49136);
nand UO_4086 (O_4086,N_47905,N_49885);
or UO_4087 (O_4087,N_47515,N_48355);
nor UO_4088 (O_4088,N_48765,N_49444);
and UO_4089 (O_4089,N_48061,N_49562);
xnor UO_4090 (O_4090,N_48466,N_49439);
xnor UO_4091 (O_4091,N_49707,N_48410);
and UO_4092 (O_4092,N_49691,N_47693);
or UO_4093 (O_4093,N_48115,N_48066);
nor UO_4094 (O_4094,N_49116,N_49645);
xnor UO_4095 (O_4095,N_49725,N_49644);
xnor UO_4096 (O_4096,N_49145,N_47591);
xor UO_4097 (O_4097,N_49083,N_48595);
xnor UO_4098 (O_4098,N_49660,N_49449);
nand UO_4099 (O_4099,N_49168,N_49721);
xor UO_4100 (O_4100,N_48222,N_49854);
or UO_4101 (O_4101,N_49937,N_48017);
xor UO_4102 (O_4102,N_48676,N_49354);
nand UO_4103 (O_4103,N_47746,N_47618);
nor UO_4104 (O_4104,N_47565,N_48701);
or UO_4105 (O_4105,N_49766,N_49818);
nor UO_4106 (O_4106,N_49212,N_48165);
or UO_4107 (O_4107,N_48990,N_48095);
and UO_4108 (O_4108,N_49083,N_47945);
nor UO_4109 (O_4109,N_49688,N_48977);
and UO_4110 (O_4110,N_49576,N_48748);
xnor UO_4111 (O_4111,N_49281,N_47642);
and UO_4112 (O_4112,N_48052,N_48609);
nor UO_4113 (O_4113,N_48673,N_47978);
nor UO_4114 (O_4114,N_49508,N_47647);
xor UO_4115 (O_4115,N_49801,N_49320);
xor UO_4116 (O_4116,N_49345,N_48216);
xor UO_4117 (O_4117,N_47504,N_48218);
nor UO_4118 (O_4118,N_48037,N_49565);
nand UO_4119 (O_4119,N_47966,N_49546);
xor UO_4120 (O_4120,N_49340,N_49030);
or UO_4121 (O_4121,N_47571,N_48000);
nor UO_4122 (O_4122,N_49853,N_49295);
and UO_4123 (O_4123,N_49133,N_49361);
or UO_4124 (O_4124,N_47559,N_49650);
nor UO_4125 (O_4125,N_48409,N_49277);
and UO_4126 (O_4126,N_49798,N_48222);
nor UO_4127 (O_4127,N_49645,N_48708);
and UO_4128 (O_4128,N_47774,N_49701);
nand UO_4129 (O_4129,N_48403,N_49605);
and UO_4130 (O_4130,N_49847,N_48234);
xnor UO_4131 (O_4131,N_49145,N_49173);
nand UO_4132 (O_4132,N_47513,N_49593);
nor UO_4133 (O_4133,N_48576,N_47757);
or UO_4134 (O_4134,N_48517,N_47968);
and UO_4135 (O_4135,N_49045,N_48357);
xor UO_4136 (O_4136,N_49178,N_49274);
and UO_4137 (O_4137,N_49417,N_48767);
nor UO_4138 (O_4138,N_49489,N_49730);
nand UO_4139 (O_4139,N_49170,N_48310);
nand UO_4140 (O_4140,N_47817,N_48077);
nor UO_4141 (O_4141,N_49415,N_49697);
or UO_4142 (O_4142,N_49177,N_48397);
xor UO_4143 (O_4143,N_49490,N_48466);
xor UO_4144 (O_4144,N_48957,N_47694);
and UO_4145 (O_4145,N_49980,N_48798);
or UO_4146 (O_4146,N_49777,N_49026);
nor UO_4147 (O_4147,N_48212,N_49228);
and UO_4148 (O_4148,N_49469,N_47935);
or UO_4149 (O_4149,N_48944,N_48746);
xnor UO_4150 (O_4150,N_48828,N_48472);
nand UO_4151 (O_4151,N_48505,N_49272);
nand UO_4152 (O_4152,N_48123,N_47526);
nor UO_4153 (O_4153,N_47857,N_47568);
nor UO_4154 (O_4154,N_49778,N_47745);
nand UO_4155 (O_4155,N_48030,N_49262);
nand UO_4156 (O_4156,N_49912,N_48247);
or UO_4157 (O_4157,N_47989,N_47629);
nor UO_4158 (O_4158,N_47875,N_47683);
or UO_4159 (O_4159,N_48687,N_47720);
xor UO_4160 (O_4160,N_49964,N_48949);
nor UO_4161 (O_4161,N_48921,N_49926);
xnor UO_4162 (O_4162,N_49738,N_47900);
xor UO_4163 (O_4163,N_49267,N_49874);
and UO_4164 (O_4164,N_48314,N_47730);
and UO_4165 (O_4165,N_49984,N_49309);
nand UO_4166 (O_4166,N_48089,N_47805);
nand UO_4167 (O_4167,N_47945,N_49327);
and UO_4168 (O_4168,N_48888,N_49754);
nand UO_4169 (O_4169,N_48818,N_49206);
nor UO_4170 (O_4170,N_49750,N_48248);
nand UO_4171 (O_4171,N_49818,N_48070);
or UO_4172 (O_4172,N_48092,N_48479);
xor UO_4173 (O_4173,N_49019,N_48804);
xnor UO_4174 (O_4174,N_48046,N_48422);
nor UO_4175 (O_4175,N_49432,N_49565);
nor UO_4176 (O_4176,N_48097,N_49146);
and UO_4177 (O_4177,N_47601,N_47738);
and UO_4178 (O_4178,N_47966,N_49326);
xnor UO_4179 (O_4179,N_49250,N_49483);
nor UO_4180 (O_4180,N_48945,N_48189);
nor UO_4181 (O_4181,N_49191,N_49448);
xnor UO_4182 (O_4182,N_47683,N_47500);
xnor UO_4183 (O_4183,N_48935,N_48891);
nor UO_4184 (O_4184,N_47655,N_48449);
nand UO_4185 (O_4185,N_48991,N_47996);
xor UO_4186 (O_4186,N_47903,N_49922);
nor UO_4187 (O_4187,N_49886,N_47809);
or UO_4188 (O_4188,N_48956,N_48264);
and UO_4189 (O_4189,N_48471,N_48305);
and UO_4190 (O_4190,N_48044,N_47984);
or UO_4191 (O_4191,N_48632,N_49063);
and UO_4192 (O_4192,N_48443,N_49439);
and UO_4193 (O_4193,N_47723,N_49755);
nor UO_4194 (O_4194,N_49076,N_48152);
nand UO_4195 (O_4195,N_48227,N_49257);
or UO_4196 (O_4196,N_48925,N_49314);
or UO_4197 (O_4197,N_49756,N_49765);
nor UO_4198 (O_4198,N_47754,N_49470);
nand UO_4199 (O_4199,N_47899,N_49225);
xnor UO_4200 (O_4200,N_49443,N_49072);
xor UO_4201 (O_4201,N_47626,N_49189);
nor UO_4202 (O_4202,N_47984,N_48060);
xnor UO_4203 (O_4203,N_48348,N_49818);
or UO_4204 (O_4204,N_48682,N_49771);
nand UO_4205 (O_4205,N_49747,N_49701);
and UO_4206 (O_4206,N_47506,N_48192);
xnor UO_4207 (O_4207,N_48730,N_48274);
and UO_4208 (O_4208,N_48372,N_49588);
nor UO_4209 (O_4209,N_48559,N_48472);
or UO_4210 (O_4210,N_47674,N_49695);
xor UO_4211 (O_4211,N_48419,N_48555);
and UO_4212 (O_4212,N_48200,N_49805);
and UO_4213 (O_4213,N_49528,N_48517);
and UO_4214 (O_4214,N_49040,N_48594);
xnor UO_4215 (O_4215,N_47597,N_47842);
and UO_4216 (O_4216,N_48871,N_49107);
nor UO_4217 (O_4217,N_47633,N_49685);
xor UO_4218 (O_4218,N_49128,N_48478);
nor UO_4219 (O_4219,N_49043,N_48760);
nand UO_4220 (O_4220,N_47542,N_49984);
or UO_4221 (O_4221,N_48950,N_49416);
nand UO_4222 (O_4222,N_48075,N_48741);
nor UO_4223 (O_4223,N_49537,N_47919);
nor UO_4224 (O_4224,N_49926,N_48756);
xor UO_4225 (O_4225,N_49092,N_49849);
nand UO_4226 (O_4226,N_49664,N_49221);
nor UO_4227 (O_4227,N_48640,N_49843);
nor UO_4228 (O_4228,N_48865,N_49006);
nor UO_4229 (O_4229,N_48647,N_49729);
or UO_4230 (O_4230,N_49629,N_49938);
and UO_4231 (O_4231,N_49324,N_49312);
xor UO_4232 (O_4232,N_47714,N_48430);
or UO_4233 (O_4233,N_47785,N_49507);
xnor UO_4234 (O_4234,N_47724,N_48507);
nor UO_4235 (O_4235,N_48766,N_48606);
nor UO_4236 (O_4236,N_49899,N_49218);
and UO_4237 (O_4237,N_49644,N_49949);
or UO_4238 (O_4238,N_47559,N_48005);
nor UO_4239 (O_4239,N_49349,N_49520);
or UO_4240 (O_4240,N_49357,N_48679);
xor UO_4241 (O_4241,N_48953,N_47668);
nor UO_4242 (O_4242,N_47864,N_48113);
xor UO_4243 (O_4243,N_48755,N_49637);
or UO_4244 (O_4244,N_48364,N_48405);
nor UO_4245 (O_4245,N_49303,N_49462);
or UO_4246 (O_4246,N_49794,N_49691);
and UO_4247 (O_4247,N_47831,N_49930);
or UO_4248 (O_4248,N_48665,N_47966);
xnor UO_4249 (O_4249,N_48246,N_49074);
and UO_4250 (O_4250,N_48655,N_47620);
xor UO_4251 (O_4251,N_48028,N_49146);
nand UO_4252 (O_4252,N_48848,N_47763);
and UO_4253 (O_4253,N_48239,N_49923);
nor UO_4254 (O_4254,N_48358,N_49772);
xor UO_4255 (O_4255,N_48848,N_48538);
xor UO_4256 (O_4256,N_47566,N_47957);
or UO_4257 (O_4257,N_49960,N_47794);
xnor UO_4258 (O_4258,N_48446,N_48645);
and UO_4259 (O_4259,N_49400,N_48878);
and UO_4260 (O_4260,N_48391,N_48500);
nand UO_4261 (O_4261,N_47545,N_49203);
nand UO_4262 (O_4262,N_49085,N_48390);
or UO_4263 (O_4263,N_49522,N_48413);
nor UO_4264 (O_4264,N_48433,N_49411);
xnor UO_4265 (O_4265,N_48370,N_49860);
and UO_4266 (O_4266,N_48181,N_48502);
and UO_4267 (O_4267,N_47770,N_49598);
nand UO_4268 (O_4268,N_49071,N_49040);
nor UO_4269 (O_4269,N_47844,N_49080);
nor UO_4270 (O_4270,N_48086,N_48302);
nand UO_4271 (O_4271,N_49915,N_49275);
nor UO_4272 (O_4272,N_48174,N_48485);
and UO_4273 (O_4273,N_49246,N_48181);
and UO_4274 (O_4274,N_48858,N_47603);
nand UO_4275 (O_4275,N_48012,N_47699);
nor UO_4276 (O_4276,N_49874,N_47700);
nor UO_4277 (O_4277,N_49237,N_47617);
or UO_4278 (O_4278,N_47827,N_48840);
and UO_4279 (O_4279,N_48140,N_49335);
xnor UO_4280 (O_4280,N_48868,N_48954);
and UO_4281 (O_4281,N_49236,N_49426);
and UO_4282 (O_4282,N_48383,N_49456);
nor UO_4283 (O_4283,N_47889,N_48393);
xnor UO_4284 (O_4284,N_48187,N_49263);
nand UO_4285 (O_4285,N_48302,N_47916);
or UO_4286 (O_4286,N_48078,N_48182);
or UO_4287 (O_4287,N_48209,N_49972);
nor UO_4288 (O_4288,N_48317,N_48955);
xor UO_4289 (O_4289,N_48932,N_49676);
xnor UO_4290 (O_4290,N_48942,N_48499);
nand UO_4291 (O_4291,N_49862,N_49219);
or UO_4292 (O_4292,N_49415,N_48409);
xnor UO_4293 (O_4293,N_49079,N_48153);
and UO_4294 (O_4294,N_49888,N_48357);
or UO_4295 (O_4295,N_47859,N_48994);
xnor UO_4296 (O_4296,N_49154,N_48965);
nor UO_4297 (O_4297,N_48767,N_49223);
nand UO_4298 (O_4298,N_49221,N_48011);
nand UO_4299 (O_4299,N_47539,N_49646);
xnor UO_4300 (O_4300,N_49566,N_49379);
or UO_4301 (O_4301,N_47958,N_48474);
nand UO_4302 (O_4302,N_48836,N_48732);
and UO_4303 (O_4303,N_48302,N_48363);
nand UO_4304 (O_4304,N_49808,N_47686);
nand UO_4305 (O_4305,N_48543,N_48667);
xor UO_4306 (O_4306,N_47726,N_48124);
and UO_4307 (O_4307,N_49832,N_49114);
nor UO_4308 (O_4308,N_49868,N_49547);
and UO_4309 (O_4309,N_49741,N_49493);
or UO_4310 (O_4310,N_49425,N_49530);
and UO_4311 (O_4311,N_48962,N_48379);
nand UO_4312 (O_4312,N_49939,N_48359);
xor UO_4313 (O_4313,N_49904,N_48222);
or UO_4314 (O_4314,N_49771,N_49124);
xor UO_4315 (O_4315,N_49131,N_49908);
or UO_4316 (O_4316,N_49323,N_48430);
xnor UO_4317 (O_4317,N_49435,N_49542);
nor UO_4318 (O_4318,N_49473,N_49970);
xor UO_4319 (O_4319,N_48426,N_49700);
and UO_4320 (O_4320,N_48026,N_48806);
nor UO_4321 (O_4321,N_49346,N_48876);
or UO_4322 (O_4322,N_47557,N_47642);
xnor UO_4323 (O_4323,N_47985,N_49960);
or UO_4324 (O_4324,N_47542,N_48349);
nand UO_4325 (O_4325,N_48488,N_48604);
or UO_4326 (O_4326,N_48629,N_48081);
or UO_4327 (O_4327,N_48596,N_47738);
nand UO_4328 (O_4328,N_49182,N_47576);
nor UO_4329 (O_4329,N_48171,N_48126);
and UO_4330 (O_4330,N_47616,N_47792);
nor UO_4331 (O_4331,N_47735,N_49854);
or UO_4332 (O_4332,N_49715,N_49425);
nand UO_4333 (O_4333,N_49224,N_48124);
nor UO_4334 (O_4334,N_49801,N_48212);
nand UO_4335 (O_4335,N_48007,N_49424);
or UO_4336 (O_4336,N_49073,N_48723);
and UO_4337 (O_4337,N_48841,N_47611);
xnor UO_4338 (O_4338,N_48936,N_47759);
and UO_4339 (O_4339,N_48492,N_49553);
nor UO_4340 (O_4340,N_49469,N_48646);
xnor UO_4341 (O_4341,N_47535,N_48197);
and UO_4342 (O_4342,N_47719,N_49020);
xnor UO_4343 (O_4343,N_47778,N_49276);
and UO_4344 (O_4344,N_48066,N_48621);
nor UO_4345 (O_4345,N_48672,N_47937);
nand UO_4346 (O_4346,N_48233,N_48118);
xor UO_4347 (O_4347,N_49970,N_48528);
nand UO_4348 (O_4348,N_48379,N_48573);
and UO_4349 (O_4349,N_48544,N_47522);
or UO_4350 (O_4350,N_49346,N_49330);
or UO_4351 (O_4351,N_49442,N_49099);
nand UO_4352 (O_4352,N_48212,N_47753);
nor UO_4353 (O_4353,N_48641,N_49988);
xor UO_4354 (O_4354,N_48925,N_48669);
xnor UO_4355 (O_4355,N_49567,N_48388);
nor UO_4356 (O_4356,N_48861,N_48075);
nor UO_4357 (O_4357,N_48983,N_47713);
nand UO_4358 (O_4358,N_48586,N_47663);
nand UO_4359 (O_4359,N_48880,N_48109);
xor UO_4360 (O_4360,N_48651,N_48266);
nor UO_4361 (O_4361,N_48565,N_49473);
nor UO_4362 (O_4362,N_48956,N_49854);
or UO_4363 (O_4363,N_49342,N_47685);
and UO_4364 (O_4364,N_49786,N_48728);
xor UO_4365 (O_4365,N_48407,N_48763);
nand UO_4366 (O_4366,N_48890,N_47970);
or UO_4367 (O_4367,N_49178,N_47752);
and UO_4368 (O_4368,N_49202,N_49752);
or UO_4369 (O_4369,N_47634,N_48763);
xnor UO_4370 (O_4370,N_48479,N_48761);
and UO_4371 (O_4371,N_47592,N_49429);
or UO_4372 (O_4372,N_49715,N_49770);
xnor UO_4373 (O_4373,N_48015,N_49105);
nand UO_4374 (O_4374,N_48523,N_47501);
nand UO_4375 (O_4375,N_48539,N_49100);
and UO_4376 (O_4376,N_48782,N_49122);
xor UO_4377 (O_4377,N_49354,N_48383);
or UO_4378 (O_4378,N_47644,N_48610);
nand UO_4379 (O_4379,N_47584,N_49341);
nor UO_4380 (O_4380,N_48782,N_49298);
nand UO_4381 (O_4381,N_49078,N_49085);
nor UO_4382 (O_4382,N_48785,N_49518);
and UO_4383 (O_4383,N_49481,N_47643);
nand UO_4384 (O_4384,N_48924,N_48447);
nand UO_4385 (O_4385,N_47827,N_48545);
nand UO_4386 (O_4386,N_49440,N_48136);
xnor UO_4387 (O_4387,N_49158,N_49303);
or UO_4388 (O_4388,N_49211,N_47754);
xnor UO_4389 (O_4389,N_48753,N_48825);
and UO_4390 (O_4390,N_47777,N_48868);
nand UO_4391 (O_4391,N_49653,N_49056);
nor UO_4392 (O_4392,N_48484,N_49806);
xor UO_4393 (O_4393,N_48418,N_47899);
xor UO_4394 (O_4394,N_49127,N_47661);
xor UO_4395 (O_4395,N_48527,N_47940);
nand UO_4396 (O_4396,N_49177,N_47703);
nor UO_4397 (O_4397,N_48862,N_48099);
nand UO_4398 (O_4398,N_49287,N_49139);
nand UO_4399 (O_4399,N_49870,N_48184);
nor UO_4400 (O_4400,N_48341,N_47703);
nand UO_4401 (O_4401,N_47556,N_49142);
and UO_4402 (O_4402,N_48257,N_48511);
xor UO_4403 (O_4403,N_49519,N_48838);
xor UO_4404 (O_4404,N_49053,N_49103);
nor UO_4405 (O_4405,N_49572,N_48838);
xor UO_4406 (O_4406,N_49854,N_48350);
nor UO_4407 (O_4407,N_47780,N_48722);
nand UO_4408 (O_4408,N_48267,N_49719);
nand UO_4409 (O_4409,N_48127,N_49489);
nor UO_4410 (O_4410,N_48206,N_47635);
nand UO_4411 (O_4411,N_48851,N_49526);
and UO_4412 (O_4412,N_49252,N_49348);
and UO_4413 (O_4413,N_49510,N_48017);
nand UO_4414 (O_4414,N_48566,N_48827);
and UO_4415 (O_4415,N_47737,N_47556);
or UO_4416 (O_4416,N_48883,N_49992);
or UO_4417 (O_4417,N_49965,N_47811);
or UO_4418 (O_4418,N_49377,N_49047);
nand UO_4419 (O_4419,N_49447,N_49831);
xnor UO_4420 (O_4420,N_48125,N_48653);
xor UO_4421 (O_4421,N_48541,N_48216);
xnor UO_4422 (O_4422,N_49060,N_49113);
nor UO_4423 (O_4423,N_49366,N_48075);
xnor UO_4424 (O_4424,N_48143,N_47680);
nor UO_4425 (O_4425,N_47808,N_48626);
nand UO_4426 (O_4426,N_47858,N_49597);
nand UO_4427 (O_4427,N_49736,N_49592);
xnor UO_4428 (O_4428,N_49264,N_47842);
xnor UO_4429 (O_4429,N_48483,N_49806);
nand UO_4430 (O_4430,N_49952,N_49345);
or UO_4431 (O_4431,N_49657,N_48021);
or UO_4432 (O_4432,N_48693,N_48301);
xnor UO_4433 (O_4433,N_48967,N_47828);
or UO_4434 (O_4434,N_47715,N_48645);
nand UO_4435 (O_4435,N_48917,N_49734);
nor UO_4436 (O_4436,N_48647,N_48227);
nand UO_4437 (O_4437,N_49209,N_49222);
nor UO_4438 (O_4438,N_47941,N_49629);
nor UO_4439 (O_4439,N_48836,N_49243);
nand UO_4440 (O_4440,N_49541,N_49733);
xor UO_4441 (O_4441,N_49378,N_47535);
nand UO_4442 (O_4442,N_48899,N_48014);
xnor UO_4443 (O_4443,N_47811,N_49184);
nand UO_4444 (O_4444,N_48815,N_48573);
xor UO_4445 (O_4445,N_48928,N_48751);
nor UO_4446 (O_4446,N_47507,N_49352);
nand UO_4447 (O_4447,N_48347,N_49828);
or UO_4448 (O_4448,N_49131,N_49266);
or UO_4449 (O_4449,N_49730,N_48455);
or UO_4450 (O_4450,N_47789,N_48605);
or UO_4451 (O_4451,N_49504,N_48104);
xor UO_4452 (O_4452,N_48194,N_49025);
xor UO_4453 (O_4453,N_48123,N_47616);
or UO_4454 (O_4454,N_49719,N_47781);
and UO_4455 (O_4455,N_47680,N_48503);
nand UO_4456 (O_4456,N_49222,N_49367);
and UO_4457 (O_4457,N_47534,N_48347);
nand UO_4458 (O_4458,N_49445,N_49355);
nand UO_4459 (O_4459,N_48759,N_47511);
nor UO_4460 (O_4460,N_47938,N_49811);
nand UO_4461 (O_4461,N_48829,N_49330);
nand UO_4462 (O_4462,N_48038,N_48793);
nor UO_4463 (O_4463,N_48608,N_47578);
xnor UO_4464 (O_4464,N_49302,N_49431);
nand UO_4465 (O_4465,N_49004,N_47784);
nand UO_4466 (O_4466,N_47706,N_48597);
nor UO_4467 (O_4467,N_49614,N_47827);
or UO_4468 (O_4468,N_48407,N_49774);
xor UO_4469 (O_4469,N_48922,N_48694);
xnor UO_4470 (O_4470,N_49404,N_48621);
and UO_4471 (O_4471,N_49924,N_47847);
nand UO_4472 (O_4472,N_48065,N_49865);
and UO_4473 (O_4473,N_48661,N_49996);
nor UO_4474 (O_4474,N_48278,N_48283);
or UO_4475 (O_4475,N_48648,N_49740);
or UO_4476 (O_4476,N_49633,N_48794);
xor UO_4477 (O_4477,N_49672,N_49000);
xor UO_4478 (O_4478,N_48351,N_47609);
xnor UO_4479 (O_4479,N_48558,N_49183);
or UO_4480 (O_4480,N_49570,N_48754);
nand UO_4481 (O_4481,N_48622,N_49454);
or UO_4482 (O_4482,N_49563,N_49872);
or UO_4483 (O_4483,N_48880,N_48928);
or UO_4484 (O_4484,N_49483,N_49765);
and UO_4485 (O_4485,N_47831,N_49824);
and UO_4486 (O_4486,N_48207,N_49924);
xor UO_4487 (O_4487,N_47775,N_47941);
nor UO_4488 (O_4488,N_49164,N_48399);
and UO_4489 (O_4489,N_49124,N_49828);
and UO_4490 (O_4490,N_49349,N_47765);
nor UO_4491 (O_4491,N_48248,N_49418);
or UO_4492 (O_4492,N_49326,N_48135);
and UO_4493 (O_4493,N_49589,N_49742);
nand UO_4494 (O_4494,N_49584,N_49720);
and UO_4495 (O_4495,N_49605,N_49832);
nand UO_4496 (O_4496,N_48200,N_48466);
nand UO_4497 (O_4497,N_49945,N_49423);
and UO_4498 (O_4498,N_49685,N_49281);
xnor UO_4499 (O_4499,N_48967,N_49790);
nand UO_4500 (O_4500,N_48783,N_49756);
xor UO_4501 (O_4501,N_49269,N_48720);
and UO_4502 (O_4502,N_49320,N_48013);
xnor UO_4503 (O_4503,N_47893,N_49925);
or UO_4504 (O_4504,N_49382,N_49788);
xor UO_4505 (O_4505,N_48595,N_49237);
and UO_4506 (O_4506,N_49881,N_48594);
nor UO_4507 (O_4507,N_48311,N_48528);
or UO_4508 (O_4508,N_47906,N_49275);
or UO_4509 (O_4509,N_49039,N_47681);
xnor UO_4510 (O_4510,N_49033,N_47788);
or UO_4511 (O_4511,N_49939,N_49550);
nand UO_4512 (O_4512,N_49865,N_49475);
nand UO_4513 (O_4513,N_49767,N_49400);
or UO_4514 (O_4514,N_49183,N_48419);
nor UO_4515 (O_4515,N_48312,N_49779);
or UO_4516 (O_4516,N_49852,N_49976);
or UO_4517 (O_4517,N_48992,N_48901);
or UO_4518 (O_4518,N_49180,N_48701);
or UO_4519 (O_4519,N_49369,N_47739);
or UO_4520 (O_4520,N_49652,N_48133);
and UO_4521 (O_4521,N_49816,N_48704);
and UO_4522 (O_4522,N_48280,N_48582);
and UO_4523 (O_4523,N_49718,N_47716);
xor UO_4524 (O_4524,N_47597,N_49024);
nand UO_4525 (O_4525,N_47758,N_48440);
and UO_4526 (O_4526,N_47576,N_49712);
nand UO_4527 (O_4527,N_49830,N_49896);
nand UO_4528 (O_4528,N_49011,N_48459);
or UO_4529 (O_4529,N_48072,N_48893);
nand UO_4530 (O_4530,N_47613,N_49972);
nand UO_4531 (O_4531,N_49853,N_47926);
nand UO_4532 (O_4532,N_48196,N_49742);
and UO_4533 (O_4533,N_49629,N_49050);
nor UO_4534 (O_4534,N_47581,N_49938);
nor UO_4535 (O_4535,N_48167,N_47562);
nor UO_4536 (O_4536,N_47928,N_48138);
and UO_4537 (O_4537,N_49698,N_49240);
and UO_4538 (O_4538,N_49475,N_49531);
or UO_4539 (O_4539,N_47789,N_49435);
or UO_4540 (O_4540,N_48279,N_47865);
xnor UO_4541 (O_4541,N_49507,N_49994);
nand UO_4542 (O_4542,N_48520,N_47541);
nor UO_4543 (O_4543,N_49930,N_48114);
nand UO_4544 (O_4544,N_47596,N_48733);
and UO_4545 (O_4545,N_47820,N_48313);
and UO_4546 (O_4546,N_48512,N_49847);
nor UO_4547 (O_4547,N_49588,N_49339);
or UO_4548 (O_4548,N_47791,N_48462);
nand UO_4549 (O_4549,N_48637,N_47873);
and UO_4550 (O_4550,N_49432,N_49981);
or UO_4551 (O_4551,N_48415,N_47995);
xor UO_4552 (O_4552,N_49126,N_47612);
xor UO_4553 (O_4553,N_48463,N_48581);
nand UO_4554 (O_4554,N_48110,N_49141);
and UO_4555 (O_4555,N_49442,N_49574);
xor UO_4556 (O_4556,N_49255,N_48982);
xor UO_4557 (O_4557,N_47555,N_47888);
xnor UO_4558 (O_4558,N_49933,N_49596);
xor UO_4559 (O_4559,N_48666,N_49751);
nor UO_4560 (O_4560,N_49751,N_48214);
and UO_4561 (O_4561,N_49676,N_48576);
xor UO_4562 (O_4562,N_48785,N_49457);
or UO_4563 (O_4563,N_49090,N_48210);
or UO_4564 (O_4564,N_47525,N_48948);
xor UO_4565 (O_4565,N_48459,N_49601);
or UO_4566 (O_4566,N_47828,N_49055);
nor UO_4567 (O_4567,N_48890,N_48431);
nand UO_4568 (O_4568,N_48227,N_49334);
xnor UO_4569 (O_4569,N_47536,N_47874);
or UO_4570 (O_4570,N_49808,N_49564);
xnor UO_4571 (O_4571,N_48884,N_49395);
xor UO_4572 (O_4572,N_49309,N_49658);
xor UO_4573 (O_4573,N_48829,N_49401);
nand UO_4574 (O_4574,N_48102,N_48048);
nor UO_4575 (O_4575,N_49502,N_48956);
and UO_4576 (O_4576,N_47618,N_49417);
nand UO_4577 (O_4577,N_48732,N_49823);
nand UO_4578 (O_4578,N_48064,N_49328);
and UO_4579 (O_4579,N_48846,N_48763);
nor UO_4580 (O_4580,N_47992,N_48704);
and UO_4581 (O_4581,N_49615,N_48462);
or UO_4582 (O_4582,N_48909,N_49616);
and UO_4583 (O_4583,N_49555,N_47597);
or UO_4584 (O_4584,N_47739,N_48879);
and UO_4585 (O_4585,N_48481,N_48414);
xnor UO_4586 (O_4586,N_47813,N_48672);
xor UO_4587 (O_4587,N_48358,N_49396);
xor UO_4588 (O_4588,N_49566,N_49261);
xor UO_4589 (O_4589,N_49338,N_47949);
and UO_4590 (O_4590,N_47801,N_48164);
and UO_4591 (O_4591,N_49109,N_47979);
xor UO_4592 (O_4592,N_49743,N_49681);
and UO_4593 (O_4593,N_49623,N_48024);
and UO_4594 (O_4594,N_48911,N_47725);
xnor UO_4595 (O_4595,N_49245,N_47623);
and UO_4596 (O_4596,N_48100,N_47957);
nand UO_4597 (O_4597,N_49485,N_49148);
and UO_4598 (O_4598,N_48263,N_48744);
xnor UO_4599 (O_4599,N_47860,N_49190);
nor UO_4600 (O_4600,N_47548,N_49062);
nand UO_4601 (O_4601,N_48335,N_49364);
nand UO_4602 (O_4602,N_49675,N_48637);
and UO_4603 (O_4603,N_49988,N_48838);
nand UO_4604 (O_4604,N_49470,N_48247);
or UO_4605 (O_4605,N_47910,N_48881);
xnor UO_4606 (O_4606,N_49150,N_47504);
and UO_4607 (O_4607,N_49740,N_49132);
nor UO_4608 (O_4608,N_49463,N_48731);
xor UO_4609 (O_4609,N_48530,N_48472);
nor UO_4610 (O_4610,N_47746,N_48070);
and UO_4611 (O_4611,N_48402,N_47624);
xor UO_4612 (O_4612,N_48349,N_49096);
nand UO_4613 (O_4613,N_48699,N_48091);
xor UO_4614 (O_4614,N_49717,N_49014);
nand UO_4615 (O_4615,N_48068,N_48583);
or UO_4616 (O_4616,N_48747,N_47791);
xnor UO_4617 (O_4617,N_48065,N_47578);
nor UO_4618 (O_4618,N_49240,N_49800);
or UO_4619 (O_4619,N_49887,N_48392);
or UO_4620 (O_4620,N_49579,N_48583);
and UO_4621 (O_4621,N_47925,N_47686);
nor UO_4622 (O_4622,N_49040,N_49466);
nand UO_4623 (O_4623,N_47856,N_49288);
xnor UO_4624 (O_4624,N_49785,N_48518);
nand UO_4625 (O_4625,N_47770,N_49985);
xnor UO_4626 (O_4626,N_49473,N_48174);
xnor UO_4627 (O_4627,N_49510,N_49954);
nand UO_4628 (O_4628,N_49454,N_49779);
and UO_4629 (O_4629,N_49483,N_49602);
nor UO_4630 (O_4630,N_48413,N_49013);
nand UO_4631 (O_4631,N_47577,N_48396);
or UO_4632 (O_4632,N_47964,N_48878);
nand UO_4633 (O_4633,N_49699,N_49978);
and UO_4634 (O_4634,N_49480,N_49901);
or UO_4635 (O_4635,N_49183,N_47959);
nand UO_4636 (O_4636,N_47929,N_47720);
or UO_4637 (O_4637,N_49840,N_47930);
or UO_4638 (O_4638,N_49492,N_47598);
xor UO_4639 (O_4639,N_48919,N_49139);
nand UO_4640 (O_4640,N_48487,N_48747);
xor UO_4641 (O_4641,N_47861,N_48371);
xor UO_4642 (O_4642,N_49967,N_49542);
and UO_4643 (O_4643,N_47778,N_49676);
or UO_4644 (O_4644,N_49641,N_48476);
or UO_4645 (O_4645,N_47550,N_49528);
xor UO_4646 (O_4646,N_49406,N_48300);
nor UO_4647 (O_4647,N_49238,N_49968);
nand UO_4648 (O_4648,N_49374,N_48645);
nand UO_4649 (O_4649,N_49886,N_49716);
xnor UO_4650 (O_4650,N_49300,N_49321);
nor UO_4651 (O_4651,N_49471,N_48374);
nand UO_4652 (O_4652,N_49356,N_49275);
or UO_4653 (O_4653,N_48316,N_49649);
nand UO_4654 (O_4654,N_48526,N_48025);
nor UO_4655 (O_4655,N_47767,N_48192);
nor UO_4656 (O_4656,N_47737,N_49427);
nor UO_4657 (O_4657,N_48601,N_49400);
xnor UO_4658 (O_4658,N_49797,N_48395);
nand UO_4659 (O_4659,N_48692,N_47850);
nor UO_4660 (O_4660,N_49448,N_48433);
xor UO_4661 (O_4661,N_49374,N_49354);
nor UO_4662 (O_4662,N_47797,N_47678);
and UO_4663 (O_4663,N_49629,N_49518);
nor UO_4664 (O_4664,N_48797,N_48086);
nand UO_4665 (O_4665,N_47843,N_48938);
or UO_4666 (O_4666,N_49791,N_49403);
nor UO_4667 (O_4667,N_48099,N_47855);
nor UO_4668 (O_4668,N_48583,N_49181);
and UO_4669 (O_4669,N_49343,N_49827);
xor UO_4670 (O_4670,N_49092,N_48715);
nor UO_4671 (O_4671,N_48339,N_49686);
or UO_4672 (O_4672,N_47808,N_47577);
nand UO_4673 (O_4673,N_47518,N_48338);
nand UO_4674 (O_4674,N_48462,N_49421);
or UO_4675 (O_4675,N_47636,N_49202);
xor UO_4676 (O_4676,N_49953,N_47631);
nand UO_4677 (O_4677,N_49616,N_48980);
or UO_4678 (O_4678,N_48285,N_48863);
xor UO_4679 (O_4679,N_49260,N_48528);
nand UO_4680 (O_4680,N_48065,N_49706);
and UO_4681 (O_4681,N_49392,N_49507);
nor UO_4682 (O_4682,N_48327,N_49142);
nand UO_4683 (O_4683,N_48063,N_49879);
xnor UO_4684 (O_4684,N_49275,N_47748);
and UO_4685 (O_4685,N_47863,N_48618);
nand UO_4686 (O_4686,N_47834,N_48634);
xor UO_4687 (O_4687,N_48685,N_48096);
nor UO_4688 (O_4688,N_49931,N_49859);
and UO_4689 (O_4689,N_49911,N_49346);
xnor UO_4690 (O_4690,N_48827,N_48425);
or UO_4691 (O_4691,N_47662,N_49204);
and UO_4692 (O_4692,N_49875,N_48072);
nand UO_4693 (O_4693,N_48280,N_49987);
xnor UO_4694 (O_4694,N_48700,N_49874);
nand UO_4695 (O_4695,N_48370,N_49561);
nor UO_4696 (O_4696,N_48200,N_49288);
nand UO_4697 (O_4697,N_49055,N_49361);
and UO_4698 (O_4698,N_47651,N_49048);
nor UO_4699 (O_4699,N_49198,N_48976);
xor UO_4700 (O_4700,N_47876,N_48392);
nand UO_4701 (O_4701,N_49520,N_49127);
nand UO_4702 (O_4702,N_48064,N_49656);
nand UO_4703 (O_4703,N_49005,N_48323);
nor UO_4704 (O_4704,N_48398,N_47529);
or UO_4705 (O_4705,N_47604,N_49050);
or UO_4706 (O_4706,N_47853,N_48270);
and UO_4707 (O_4707,N_48798,N_49477);
or UO_4708 (O_4708,N_48252,N_49836);
and UO_4709 (O_4709,N_49179,N_48979);
xor UO_4710 (O_4710,N_47713,N_49782);
or UO_4711 (O_4711,N_47800,N_47997);
or UO_4712 (O_4712,N_48088,N_48240);
nand UO_4713 (O_4713,N_48434,N_48882);
or UO_4714 (O_4714,N_47970,N_49981);
or UO_4715 (O_4715,N_49420,N_49329);
nand UO_4716 (O_4716,N_49031,N_48098);
nor UO_4717 (O_4717,N_48938,N_49598);
and UO_4718 (O_4718,N_49222,N_47773);
nand UO_4719 (O_4719,N_48315,N_49509);
nand UO_4720 (O_4720,N_49851,N_49494);
nand UO_4721 (O_4721,N_47776,N_49148);
or UO_4722 (O_4722,N_48156,N_47864);
or UO_4723 (O_4723,N_48995,N_47578);
nor UO_4724 (O_4724,N_48175,N_48420);
xor UO_4725 (O_4725,N_48199,N_47588);
nand UO_4726 (O_4726,N_48863,N_48372);
nand UO_4727 (O_4727,N_49701,N_48780);
nand UO_4728 (O_4728,N_49020,N_47737);
and UO_4729 (O_4729,N_49709,N_48306);
and UO_4730 (O_4730,N_48886,N_48486);
nor UO_4731 (O_4731,N_47936,N_49164);
nand UO_4732 (O_4732,N_47608,N_48746);
nor UO_4733 (O_4733,N_47739,N_48954);
nand UO_4734 (O_4734,N_48670,N_48726);
or UO_4735 (O_4735,N_48364,N_49580);
or UO_4736 (O_4736,N_48895,N_48291);
nand UO_4737 (O_4737,N_49396,N_48870);
nor UO_4738 (O_4738,N_47509,N_47515);
nand UO_4739 (O_4739,N_49553,N_47596);
and UO_4740 (O_4740,N_47821,N_48060);
or UO_4741 (O_4741,N_49605,N_48511);
and UO_4742 (O_4742,N_48914,N_49719);
nor UO_4743 (O_4743,N_48410,N_49163);
or UO_4744 (O_4744,N_48286,N_47961);
xor UO_4745 (O_4745,N_48145,N_47701);
and UO_4746 (O_4746,N_48137,N_47625);
xnor UO_4747 (O_4747,N_48026,N_47621);
nand UO_4748 (O_4748,N_48266,N_49029);
xor UO_4749 (O_4749,N_47888,N_48690);
and UO_4750 (O_4750,N_49168,N_48494);
nand UO_4751 (O_4751,N_48317,N_48191);
xor UO_4752 (O_4752,N_47842,N_47894);
or UO_4753 (O_4753,N_48455,N_48774);
nor UO_4754 (O_4754,N_49960,N_49938);
and UO_4755 (O_4755,N_49162,N_49895);
and UO_4756 (O_4756,N_49585,N_49299);
nor UO_4757 (O_4757,N_49990,N_47876);
xor UO_4758 (O_4758,N_48347,N_47922);
xnor UO_4759 (O_4759,N_48339,N_47745);
xnor UO_4760 (O_4760,N_49547,N_48429);
xor UO_4761 (O_4761,N_48415,N_48039);
nor UO_4762 (O_4762,N_49805,N_47696);
nand UO_4763 (O_4763,N_47881,N_47742);
nand UO_4764 (O_4764,N_48500,N_48068);
and UO_4765 (O_4765,N_48173,N_47749);
and UO_4766 (O_4766,N_49508,N_48284);
and UO_4767 (O_4767,N_49031,N_47917);
and UO_4768 (O_4768,N_49028,N_49996);
nor UO_4769 (O_4769,N_47834,N_49067);
nor UO_4770 (O_4770,N_49795,N_47609);
nor UO_4771 (O_4771,N_48695,N_48999);
nand UO_4772 (O_4772,N_49599,N_48868);
or UO_4773 (O_4773,N_49053,N_48873);
and UO_4774 (O_4774,N_48054,N_48356);
and UO_4775 (O_4775,N_48804,N_49346);
and UO_4776 (O_4776,N_48827,N_47918);
nand UO_4777 (O_4777,N_49300,N_49794);
and UO_4778 (O_4778,N_47881,N_48029);
nand UO_4779 (O_4779,N_47598,N_49545);
xor UO_4780 (O_4780,N_48166,N_49568);
or UO_4781 (O_4781,N_48490,N_49458);
nand UO_4782 (O_4782,N_49643,N_49914);
nor UO_4783 (O_4783,N_47607,N_49390);
nand UO_4784 (O_4784,N_47535,N_47987);
nand UO_4785 (O_4785,N_48262,N_49040);
and UO_4786 (O_4786,N_48965,N_49678);
nand UO_4787 (O_4787,N_47885,N_47565);
and UO_4788 (O_4788,N_49160,N_49957);
and UO_4789 (O_4789,N_49277,N_47845);
and UO_4790 (O_4790,N_49692,N_47939);
xnor UO_4791 (O_4791,N_47670,N_48318);
nor UO_4792 (O_4792,N_48008,N_47850);
xnor UO_4793 (O_4793,N_49330,N_48640);
xor UO_4794 (O_4794,N_49330,N_48729);
and UO_4795 (O_4795,N_49618,N_47794);
nand UO_4796 (O_4796,N_49616,N_48844);
or UO_4797 (O_4797,N_47841,N_49327);
nor UO_4798 (O_4798,N_49345,N_49698);
nor UO_4799 (O_4799,N_49226,N_47966);
nand UO_4800 (O_4800,N_48225,N_49853);
nand UO_4801 (O_4801,N_48788,N_48075);
and UO_4802 (O_4802,N_49060,N_47815);
nor UO_4803 (O_4803,N_48651,N_49659);
nor UO_4804 (O_4804,N_47519,N_47745);
xnor UO_4805 (O_4805,N_47584,N_47589);
or UO_4806 (O_4806,N_47776,N_48298);
nor UO_4807 (O_4807,N_49691,N_49612);
or UO_4808 (O_4808,N_49253,N_48340);
and UO_4809 (O_4809,N_47799,N_48748);
nand UO_4810 (O_4810,N_49943,N_48974);
nor UO_4811 (O_4811,N_49735,N_48723);
or UO_4812 (O_4812,N_49899,N_49747);
and UO_4813 (O_4813,N_48449,N_49340);
nor UO_4814 (O_4814,N_49596,N_48095);
and UO_4815 (O_4815,N_47734,N_49431);
xor UO_4816 (O_4816,N_47907,N_47904);
and UO_4817 (O_4817,N_48321,N_48596);
nand UO_4818 (O_4818,N_48458,N_49197);
xnor UO_4819 (O_4819,N_49578,N_48210);
xnor UO_4820 (O_4820,N_48531,N_48621);
and UO_4821 (O_4821,N_48615,N_49921);
nor UO_4822 (O_4822,N_48855,N_49763);
xnor UO_4823 (O_4823,N_49025,N_47697);
xnor UO_4824 (O_4824,N_48115,N_48567);
and UO_4825 (O_4825,N_49572,N_49412);
nor UO_4826 (O_4826,N_48976,N_49439);
or UO_4827 (O_4827,N_49238,N_49842);
nand UO_4828 (O_4828,N_48947,N_49549);
nand UO_4829 (O_4829,N_47696,N_47568);
nand UO_4830 (O_4830,N_49062,N_48890);
nor UO_4831 (O_4831,N_48538,N_49154);
nand UO_4832 (O_4832,N_48019,N_49245);
xnor UO_4833 (O_4833,N_49258,N_48410);
and UO_4834 (O_4834,N_48007,N_47567);
nand UO_4835 (O_4835,N_49453,N_49143);
nand UO_4836 (O_4836,N_49983,N_48539);
and UO_4837 (O_4837,N_49019,N_49599);
and UO_4838 (O_4838,N_49275,N_48312);
xor UO_4839 (O_4839,N_49183,N_49054);
and UO_4840 (O_4840,N_49037,N_48154);
or UO_4841 (O_4841,N_49142,N_48340);
or UO_4842 (O_4842,N_48305,N_48089);
or UO_4843 (O_4843,N_48575,N_47563);
xor UO_4844 (O_4844,N_48675,N_48789);
nor UO_4845 (O_4845,N_47934,N_47887);
or UO_4846 (O_4846,N_48797,N_49280);
xor UO_4847 (O_4847,N_49376,N_47670);
and UO_4848 (O_4848,N_47998,N_48143);
or UO_4849 (O_4849,N_48129,N_49975);
and UO_4850 (O_4850,N_47965,N_49521);
nand UO_4851 (O_4851,N_48148,N_48624);
or UO_4852 (O_4852,N_48374,N_49170);
xor UO_4853 (O_4853,N_48536,N_48858);
nand UO_4854 (O_4854,N_48935,N_47974);
nor UO_4855 (O_4855,N_48726,N_48627);
and UO_4856 (O_4856,N_48671,N_47882);
nand UO_4857 (O_4857,N_48581,N_47772);
and UO_4858 (O_4858,N_48709,N_49466);
nand UO_4859 (O_4859,N_49732,N_48997);
or UO_4860 (O_4860,N_49023,N_49193);
xnor UO_4861 (O_4861,N_49756,N_48881);
and UO_4862 (O_4862,N_49118,N_49335);
or UO_4863 (O_4863,N_49939,N_48548);
or UO_4864 (O_4864,N_48976,N_48916);
xor UO_4865 (O_4865,N_48739,N_47825);
and UO_4866 (O_4866,N_49042,N_49325);
and UO_4867 (O_4867,N_48674,N_47852);
nor UO_4868 (O_4868,N_49835,N_48127);
nand UO_4869 (O_4869,N_49493,N_49989);
nor UO_4870 (O_4870,N_49510,N_49665);
nand UO_4871 (O_4871,N_48187,N_48865);
or UO_4872 (O_4872,N_49286,N_48074);
and UO_4873 (O_4873,N_47681,N_48265);
or UO_4874 (O_4874,N_48912,N_49804);
xnor UO_4875 (O_4875,N_48397,N_49379);
and UO_4876 (O_4876,N_49482,N_49273);
xnor UO_4877 (O_4877,N_49742,N_48397);
and UO_4878 (O_4878,N_49202,N_48551);
or UO_4879 (O_4879,N_48899,N_47606);
nor UO_4880 (O_4880,N_49672,N_48347);
nand UO_4881 (O_4881,N_49053,N_47510);
nand UO_4882 (O_4882,N_49638,N_49331);
nor UO_4883 (O_4883,N_48705,N_49953);
xnor UO_4884 (O_4884,N_47567,N_48392);
xnor UO_4885 (O_4885,N_48592,N_48514);
nand UO_4886 (O_4886,N_48704,N_48059);
and UO_4887 (O_4887,N_48575,N_49671);
xnor UO_4888 (O_4888,N_49921,N_48279);
and UO_4889 (O_4889,N_47547,N_48121);
xor UO_4890 (O_4890,N_47816,N_47644);
xnor UO_4891 (O_4891,N_47648,N_49361);
xor UO_4892 (O_4892,N_49903,N_48328);
xnor UO_4893 (O_4893,N_47941,N_48749);
nor UO_4894 (O_4894,N_49694,N_48889);
xor UO_4895 (O_4895,N_49381,N_47977);
or UO_4896 (O_4896,N_49899,N_49339);
or UO_4897 (O_4897,N_49986,N_48438);
and UO_4898 (O_4898,N_48756,N_48200);
xor UO_4899 (O_4899,N_48733,N_48291);
and UO_4900 (O_4900,N_48958,N_49637);
nand UO_4901 (O_4901,N_49579,N_47709);
and UO_4902 (O_4902,N_49048,N_47697);
nand UO_4903 (O_4903,N_48699,N_49859);
nand UO_4904 (O_4904,N_47899,N_48734);
nand UO_4905 (O_4905,N_49942,N_47564);
nor UO_4906 (O_4906,N_49897,N_49828);
xnor UO_4907 (O_4907,N_47938,N_49533);
nor UO_4908 (O_4908,N_48429,N_47910);
xor UO_4909 (O_4909,N_49052,N_49406);
nand UO_4910 (O_4910,N_48157,N_49596);
and UO_4911 (O_4911,N_48982,N_47938);
xor UO_4912 (O_4912,N_49654,N_47916);
xnor UO_4913 (O_4913,N_49097,N_48568);
xnor UO_4914 (O_4914,N_48194,N_48960);
or UO_4915 (O_4915,N_49371,N_49128);
nor UO_4916 (O_4916,N_49081,N_48283);
and UO_4917 (O_4917,N_48056,N_48602);
nand UO_4918 (O_4918,N_47606,N_49150);
nor UO_4919 (O_4919,N_49620,N_49819);
xnor UO_4920 (O_4920,N_49540,N_48373);
and UO_4921 (O_4921,N_49117,N_47943);
and UO_4922 (O_4922,N_48150,N_49254);
xnor UO_4923 (O_4923,N_47630,N_48731);
and UO_4924 (O_4924,N_49378,N_48154);
or UO_4925 (O_4925,N_48797,N_49923);
or UO_4926 (O_4926,N_48438,N_49098);
or UO_4927 (O_4927,N_49060,N_47648);
nand UO_4928 (O_4928,N_47828,N_47931);
nor UO_4929 (O_4929,N_49247,N_49995);
xor UO_4930 (O_4930,N_48899,N_48046);
xnor UO_4931 (O_4931,N_48177,N_47938);
xor UO_4932 (O_4932,N_48730,N_47826);
nand UO_4933 (O_4933,N_49695,N_48457);
and UO_4934 (O_4934,N_48173,N_49192);
nor UO_4935 (O_4935,N_48026,N_49946);
xor UO_4936 (O_4936,N_49936,N_48899);
and UO_4937 (O_4937,N_49562,N_49910);
xnor UO_4938 (O_4938,N_48836,N_47840);
or UO_4939 (O_4939,N_47636,N_48689);
nor UO_4940 (O_4940,N_47668,N_48852);
nand UO_4941 (O_4941,N_48535,N_48168);
xnor UO_4942 (O_4942,N_47508,N_49210);
nor UO_4943 (O_4943,N_49851,N_47562);
nand UO_4944 (O_4944,N_48959,N_48495);
nor UO_4945 (O_4945,N_49603,N_49259);
nor UO_4946 (O_4946,N_48790,N_47971);
xor UO_4947 (O_4947,N_49724,N_49004);
nand UO_4948 (O_4948,N_47771,N_49413);
nand UO_4949 (O_4949,N_48998,N_49303);
and UO_4950 (O_4950,N_48834,N_48554);
or UO_4951 (O_4951,N_47702,N_47670);
xor UO_4952 (O_4952,N_48449,N_48068);
nand UO_4953 (O_4953,N_49928,N_48903);
nor UO_4954 (O_4954,N_48884,N_48578);
or UO_4955 (O_4955,N_49396,N_48460);
and UO_4956 (O_4956,N_48457,N_49844);
or UO_4957 (O_4957,N_48747,N_47628);
nand UO_4958 (O_4958,N_49399,N_49246);
and UO_4959 (O_4959,N_48851,N_49901);
or UO_4960 (O_4960,N_48617,N_48266);
or UO_4961 (O_4961,N_49727,N_49470);
or UO_4962 (O_4962,N_49319,N_48737);
nand UO_4963 (O_4963,N_47648,N_47518);
and UO_4964 (O_4964,N_49136,N_49602);
xor UO_4965 (O_4965,N_49130,N_48574);
xnor UO_4966 (O_4966,N_49138,N_48308);
or UO_4967 (O_4967,N_47579,N_49994);
nand UO_4968 (O_4968,N_48543,N_49582);
and UO_4969 (O_4969,N_49889,N_49101);
nor UO_4970 (O_4970,N_49494,N_47922);
and UO_4971 (O_4971,N_49920,N_48416);
xor UO_4972 (O_4972,N_49466,N_47587);
or UO_4973 (O_4973,N_48444,N_49963);
xor UO_4974 (O_4974,N_48615,N_47942);
nand UO_4975 (O_4975,N_49176,N_48979);
nor UO_4976 (O_4976,N_48837,N_48263);
or UO_4977 (O_4977,N_48842,N_49021);
nor UO_4978 (O_4978,N_48311,N_47520);
and UO_4979 (O_4979,N_47577,N_47692);
xor UO_4980 (O_4980,N_48194,N_48539);
or UO_4981 (O_4981,N_47763,N_49746);
and UO_4982 (O_4982,N_49084,N_48871);
and UO_4983 (O_4983,N_49859,N_47698);
xor UO_4984 (O_4984,N_49155,N_49355);
xor UO_4985 (O_4985,N_48817,N_49119);
xnor UO_4986 (O_4986,N_48928,N_49896);
nand UO_4987 (O_4987,N_47930,N_48240);
xnor UO_4988 (O_4988,N_48263,N_47526);
and UO_4989 (O_4989,N_47555,N_49918);
nand UO_4990 (O_4990,N_49263,N_48284);
nand UO_4991 (O_4991,N_48758,N_49462);
nand UO_4992 (O_4992,N_49175,N_47633);
nor UO_4993 (O_4993,N_49289,N_49265);
and UO_4994 (O_4994,N_48920,N_48677);
and UO_4995 (O_4995,N_48482,N_47699);
or UO_4996 (O_4996,N_48139,N_49753);
xnor UO_4997 (O_4997,N_47549,N_49844);
nand UO_4998 (O_4998,N_49622,N_48532);
or UO_4999 (O_4999,N_49863,N_47823);
endmodule