module basic_1000_10000_1500_4_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nand U0 (N_0,In_580,In_51);
or U1 (N_1,In_944,In_832);
and U2 (N_2,In_567,In_57);
nor U3 (N_3,In_984,In_824);
xnor U4 (N_4,In_309,In_971);
nand U5 (N_5,In_574,In_578);
nor U6 (N_6,In_925,In_412);
xnor U7 (N_7,In_263,In_127);
nor U8 (N_8,In_349,In_674);
and U9 (N_9,In_593,In_600);
xnor U10 (N_10,In_129,In_555);
or U11 (N_11,In_371,In_59);
nand U12 (N_12,In_415,In_22);
or U13 (N_13,In_115,In_377);
nor U14 (N_14,In_262,In_691);
nor U15 (N_15,In_446,In_778);
and U16 (N_16,In_547,In_135);
or U17 (N_17,In_788,In_267);
xnor U18 (N_18,In_724,In_861);
nand U19 (N_19,In_546,In_467);
nor U20 (N_20,In_151,In_763);
or U21 (N_21,In_562,In_896);
nor U22 (N_22,In_474,In_764);
and U23 (N_23,In_903,In_254);
xnor U24 (N_24,In_950,In_240);
nor U25 (N_25,In_176,In_797);
nand U26 (N_26,In_17,In_959);
or U27 (N_27,In_384,In_95);
or U28 (N_28,In_440,In_613);
xnor U29 (N_29,In_529,In_952);
nand U30 (N_30,In_475,In_623);
xor U31 (N_31,In_740,In_496);
xor U32 (N_32,In_414,In_809);
or U33 (N_33,In_927,In_65);
or U34 (N_34,In_715,In_926);
and U35 (N_35,In_268,In_31);
and U36 (N_36,In_448,In_160);
nor U37 (N_37,In_921,In_808);
nor U38 (N_38,In_500,In_589);
xor U39 (N_39,In_329,In_11);
and U40 (N_40,In_295,In_779);
xor U41 (N_41,In_66,In_429);
xor U42 (N_42,In_15,In_835);
and U43 (N_43,In_131,In_834);
nor U44 (N_44,In_596,In_234);
xor U45 (N_45,In_445,In_469);
nor U46 (N_46,In_464,In_677);
nand U47 (N_47,In_848,In_482);
or U48 (N_48,In_790,In_292);
xnor U49 (N_49,In_58,In_557);
nand U50 (N_50,In_199,In_0);
and U51 (N_51,In_172,In_275);
nor U52 (N_52,In_558,In_897);
nand U53 (N_53,In_726,In_618);
or U54 (N_54,In_791,In_599);
or U55 (N_55,In_661,In_439);
and U56 (N_56,In_857,In_82);
and U57 (N_57,In_785,In_717);
nand U58 (N_58,In_539,In_990);
or U59 (N_59,In_572,In_901);
or U60 (N_60,In_163,In_957);
and U61 (N_61,In_992,In_205);
or U62 (N_62,In_209,In_516);
or U63 (N_63,In_276,In_781);
or U64 (N_64,In_895,In_284);
nand U65 (N_65,In_468,In_281);
nand U66 (N_66,In_583,In_391);
or U67 (N_67,In_755,In_657);
xor U68 (N_68,In_62,In_366);
or U69 (N_69,In_194,In_739);
xnor U70 (N_70,In_41,In_345);
and U71 (N_71,In_481,In_751);
nand U72 (N_72,In_916,In_149);
xnor U73 (N_73,In_928,In_289);
and U74 (N_74,In_322,In_710);
nor U75 (N_75,In_706,In_455);
nor U76 (N_76,In_633,In_113);
nor U77 (N_77,In_940,In_510);
nand U78 (N_78,In_884,In_659);
nor U79 (N_79,In_90,In_307);
or U80 (N_80,In_830,In_25);
or U81 (N_81,In_478,In_827);
and U82 (N_82,In_712,In_491);
nor U83 (N_83,In_817,In_932);
and U84 (N_84,In_609,In_994);
nand U85 (N_85,In_296,In_372);
xnor U86 (N_86,In_69,In_261);
nor U87 (N_87,In_577,In_531);
or U88 (N_88,In_140,In_612);
xor U89 (N_89,In_356,In_308);
nor U90 (N_90,In_846,In_663);
nor U91 (N_91,In_383,In_148);
nand U92 (N_92,In_625,In_795);
nand U93 (N_93,In_631,In_907);
and U94 (N_94,In_53,In_452);
or U95 (N_95,In_286,In_882);
xnor U96 (N_96,In_967,In_693);
and U97 (N_97,In_590,In_762);
or U98 (N_98,In_550,In_158);
and U99 (N_99,In_894,In_509);
or U100 (N_100,In_368,In_310);
xnor U101 (N_101,In_568,In_634);
nor U102 (N_102,In_997,In_863);
or U103 (N_103,In_416,In_694);
nor U104 (N_104,In_771,In_876);
nand U105 (N_105,In_576,In_406);
nor U106 (N_106,In_201,In_251);
or U107 (N_107,In_141,In_999);
nand U108 (N_108,In_887,In_192);
and U109 (N_109,In_662,In_867);
xor U110 (N_110,In_741,In_956);
nand U111 (N_111,In_421,In_21);
and U112 (N_112,In_128,In_881);
or U113 (N_113,In_112,In_167);
nor U114 (N_114,In_981,In_313);
xnor U115 (N_115,In_472,In_266);
nor U116 (N_116,In_891,In_423);
nand U117 (N_117,In_551,In_389);
nand U118 (N_118,In_731,In_92);
nand U119 (N_119,In_6,In_498);
and U120 (N_120,In_507,In_290);
and U121 (N_121,In_875,In_961);
nand U122 (N_122,In_330,In_264);
and U123 (N_123,In_379,In_864);
nand U124 (N_124,In_769,In_231);
nor U125 (N_125,In_923,In_180);
nor U126 (N_126,In_906,In_913);
nor U127 (N_127,In_336,In_637);
nor U128 (N_128,In_941,In_660);
xnor U129 (N_129,In_460,In_648);
xor U130 (N_130,In_407,In_513);
and U131 (N_131,In_506,In_859);
nor U132 (N_132,In_304,In_963);
nand U133 (N_133,In_86,In_658);
xnor U134 (N_134,In_239,In_342);
xor U135 (N_135,In_444,In_252);
nor U136 (N_136,In_611,In_890);
or U137 (N_137,In_560,In_838);
and U138 (N_138,In_530,In_986);
nand U139 (N_139,In_137,In_341);
and U140 (N_140,In_222,In_899);
nand U141 (N_141,In_493,In_87);
nor U142 (N_142,In_584,In_632);
or U143 (N_143,In_398,In_705);
or U144 (N_144,In_975,In_753);
nand U145 (N_145,In_43,In_607);
nand U146 (N_146,In_48,In_74);
and U147 (N_147,In_118,In_619);
and U148 (N_148,In_968,In_9);
and U149 (N_149,In_579,In_554);
nand U150 (N_150,In_422,In_425);
or U151 (N_151,In_219,In_652);
and U152 (N_152,In_316,In_453);
nand U153 (N_153,In_136,In_980);
and U154 (N_154,In_616,In_919);
nor U155 (N_155,In_459,In_285);
xor U156 (N_156,In_72,In_883);
and U157 (N_157,In_256,In_768);
xnor U158 (N_158,In_435,In_484);
or U159 (N_159,In_936,In_299);
or U160 (N_160,In_47,In_335);
or U161 (N_161,In_247,In_365);
nor U162 (N_162,In_678,In_643);
xor U163 (N_163,In_945,In_536);
or U164 (N_164,In_738,In_178);
or U165 (N_165,In_543,In_338);
and U166 (N_166,In_965,In_248);
or U167 (N_167,In_253,In_426);
or U168 (N_168,In_725,In_357);
and U169 (N_169,In_886,In_54);
xor U170 (N_170,In_328,In_799);
nand U171 (N_171,In_775,In_120);
and U172 (N_172,In_359,In_332);
and U173 (N_173,In_979,In_76);
nor U174 (N_174,In_541,In_465);
nor U175 (N_175,In_798,In_733);
nand U176 (N_176,In_278,In_38);
and U177 (N_177,In_471,In_436);
and U178 (N_178,In_215,In_32);
or U179 (N_179,In_796,In_703);
nand U180 (N_180,In_5,In_851);
nand U181 (N_181,In_63,In_535);
or U182 (N_182,In_918,In_696);
nor U183 (N_183,In_517,In_184);
or U184 (N_184,In_362,In_348);
or U185 (N_185,In_855,In_563);
xor U186 (N_186,In_317,In_300);
or U187 (N_187,In_282,In_973);
nor U188 (N_188,In_628,In_917);
nand U189 (N_189,In_872,In_494);
or U190 (N_190,In_404,In_102);
and U191 (N_191,In_807,In_719);
nor U192 (N_192,In_879,In_972);
nand U193 (N_193,In_364,In_243);
and U194 (N_194,In_470,In_321);
nand U195 (N_195,In_238,In_327);
and U196 (N_196,In_559,In_649);
nor U197 (N_197,In_224,In_323);
or U198 (N_198,In_697,In_138);
and U199 (N_199,In_164,In_44);
or U200 (N_200,In_33,In_642);
nor U201 (N_201,In_360,In_608);
or U202 (N_202,In_193,In_314);
nand U203 (N_203,In_487,In_523);
xor U204 (N_204,In_951,In_743);
nand U205 (N_205,In_433,In_647);
xnor U206 (N_206,In_594,In_269);
nor U207 (N_207,In_280,In_37);
nand U208 (N_208,In_67,In_331);
and U209 (N_209,In_626,In_56);
nor U210 (N_210,In_214,In_991);
and U211 (N_211,In_424,In_68);
or U212 (N_212,In_392,In_671);
or U213 (N_213,In_303,In_221);
nor U214 (N_214,In_822,In_676);
xor U215 (N_215,In_888,In_746);
or U216 (N_216,In_34,In_1);
nor U217 (N_217,In_169,In_728);
nand U218 (N_218,In_977,In_93);
nand U219 (N_219,In_443,In_854);
nor U220 (N_220,In_143,In_675);
and U221 (N_221,In_191,In_98);
nand U222 (N_222,In_985,In_512);
xnor U223 (N_223,In_124,In_587);
xnor U224 (N_224,In_575,In_302);
nor U225 (N_225,In_157,In_792);
or U226 (N_226,In_198,In_130);
and U227 (N_227,In_108,In_374);
or U228 (N_228,In_187,In_966);
nor U229 (N_229,In_103,In_672);
nand U230 (N_230,In_821,In_730);
or U231 (N_231,In_905,In_858);
xor U232 (N_232,In_721,In_376);
or U233 (N_233,In_434,In_85);
nand U234 (N_234,In_339,In_598);
nor U235 (N_235,In_355,In_704);
and U236 (N_236,In_334,In_777);
xor U237 (N_237,In_104,In_670);
or U238 (N_238,In_499,In_639);
xnor U239 (N_239,In_350,In_183);
and U240 (N_240,In_2,In_767);
and U241 (N_241,In_566,In_549);
xor U242 (N_242,In_766,In_418);
and U243 (N_243,In_570,In_789);
xor U244 (N_244,In_97,In_734);
nor U245 (N_245,In_301,In_116);
and U246 (N_246,In_892,In_390);
or U247 (N_247,In_89,In_351);
or U248 (N_248,In_942,In_868);
or U249 (N_249,In_159,In_630);
nand U250 (N_250,In_606,In_912);
or U251 (N_251,In_837,In_24);
or U252 (N_252,In_408,In_603);
nor U253 (N_253,In_688,In_409);
nand U254 (N_254,In_381,In_430);
nor U255 (N_255,In_370,In_569);
or U256 (N_256,In_841,In_154);
and U257 (N_257,In_196,In_353);
nand U258 (N_258,In_524,In_451);
and U259 (N_259,In_490,In_644);
and U260 (N_260,In_902,In_689);
and U261 (N_261,In_312,In_477);
nor U262 (N_262,In_935,In_400);
xor U263 (N_263,In_571,In_417);
nor U264 (N_264,In_748,In_287);
or U265 (N_265,In_197,In_23);
and U266 (N_266,In_449,In_126);
and U267 (N_267,In_319,In_969);
nand U268 (N_268,In_700,In_88);
nor U269 (N_269,In_654,In_121);
or U270 (N_270,In_403,In_656);
nand U271 (N_271,In_166,In_757);
or U272 (N_272,In_582,In_621);
nor U273 (N_273,In_650,In_745);
or U274 (N_274,In_702,In_119);
nand U275 (N_275,In_801,In_52);
or U276 (N_276,In_291,In_7);
nor U277 (N_277,In_683,In_288);
and U278 (N_278,In_16,In_604);
xor U279 (N_279,In_463,In_19);
and U280 (N_280,In_271,In_347);
and U281 (N_281,In_836,In_784);
or U282 (N_282,In_709,In_640);
and U283 (N_283,In_908,In_525);
xnor U284 (N_284,In_318,In_20);
and U285 (N_285,In_889,In_948);
nand U286 (N_286,In_714,In_871);
xnor U287 (N_287,In_727,In_615);
xor U288 (N_288,In_367,In_235);
nand U289 (N_289,In_344,In_823);
xor U290 (N_290,In_458,In_614);
xor U291 (N_291,In_283,In_489);
xnor U292 (N_292,In_50,In_847);
and U293 (N_293,In_190,In_242);
or U294 (N_294,In_962,In_937);
nor U295 (N_295,In_776,In_189);
nand U296 (N_296,In_849,In_686);
xor U297 (N_297,In_664,In_825);
and U298 (N_298,In_79,In_810);
nand U299 (N_299,In_915,In_910);
xnor U300 (N_300,In_358,In_842);
or U301 (N_301,In_49,In_736);
or U302 (N_302,In_690,In_761);
xor U303 (N_303,In_179,In_211);
or U304 (N_304,In_732,In_18);
nor U305 (N_305,In_207,In_538);
xor U306 (N_306,In_259,In_852);
or U307 (N_307,In_635,In_305);
nor U308 (N_308,In_363,In_99);
nand U309 (N_309,In_955,In_396);
or U310 (N_310,In_713,In_518);
xnor U311 (N_311,In_64,In_28);
nor U312 (N_312,In_954,In_636);
nor U313 (N_313,In_929,In_241);
or U314 (N_314,In_174,In_641);
nand U315 (N_315,In_816,In_900);
nor U316 (N_316,In_337,In_12);
and U317 (N_317,In_306,In_814);
and U318 (N_318,In_134,In_315);
nor U319 (N_319,In_682,In_142);
and U320 (N_320,In_354,In_601);
xor U321 (N_321,In_39,In_185);
and U322 (N_322,In_186,In_441);
or U323 (N_323,In_820,In_976);
and U324 (N_324,In_236,In_934);
and U325 (N_325,In_399,In_35);
nand U326 (N_326,In_805,In_462);
nor U327 (N_327,In_447,In_685);
nand U328 (N_328,In_831,In_3);
nand U329 (N_329,In_534,In_324);
and U330 (N_330,In_216,In_898);
xor U331 (N_331,In_46,In_856);
or U332 (N_332,In_100,In_553);
nand U333 (N_333,In_77,In_387);
and U334 (N_334,In_556,In_749);
or U335 (N_335,In_701,In_161);
and U336 (N_336,In_212,In_495);
nand U337 (N_337,In_655,In_297);
xor U338 (N_338,In_385,In_438);
nor U339 (N_339,In_270,In_27);
or U340 (N_340,In_233,In_497);
and U341 (N_341,In_146,In_819);
nor U342 (N_342,In_218,In_565);
or U343 (N_343,In_226,In_537);
or U344 (N_344,In_772,In_953);
xnor U345 (N_345,In_720,In_737);
and U346 (N_346,In_504,In_723);
xnor U347 (N_347,In_274,In_73);
xnor U348 (N_348,In_812,In_585);
or U349 (N_349,In_393,In_346);
or U350 (N_350,In_420,In_800);
nand U351 (N_351,In_803,In_227);
nor U352 (N_352,In_277,In_26);
xnor U353 (N_353,In_419,In_844);
xor U354 (N_354,In_681,In_60);
nor U355 (N_355,In_114,In_101);
and U356 (N_356,In_181,In_454);
nand U357 (N_357,In_480,In_561);
nor U358 (N_358,In_109,In_150);
and U359 (N_359,In_911,In_665);
nand U360 (N_360,In_786,In_747);
and U361 (N_361,In_29,In_182);
or U362 (N_362,In_492,In_30);
or U363 (N_363,In_502,In_545);
and U364 (N_364,In_442,In_145);
nor U365 (N_365,In_208,In_228);
or U366 (N_366,In_437,In_380);
xnor U367 (N_367,In_605,In_760);
xnor U368 (N_368,In_8,In_202);
nor U369 (N_369,In_361,In_397);
nor U370 (N_370,In_729,In_210);
nand U371 (N_371,In_853,In_645);
nor U372 (N_372,In_744,In_943);
nor U373 (N_373,In_684,In_326);
nand U374 (N_374,In_987,In_461);
or U375 (N_375,In_177,In_405);
xor U376 (N_376,In_257,In_806);
and U377 (N_377,In_175,In_410);
nor U378 (N_378,In_610,In_272);
nor U379 (N_379,In_964,In_107);
xnor U380 (N_380,In_666,In_42);
nand U381 (N_381,In_217,In_783);
nand U382 (N_382,In_687,In_970);
nand U383 (N_383,In_933,In_14);
nand U384 (N_384,In_246,In_520);
and U385 (N_385,In_388,In_223);
xnor U386 (N_386,In_958,In_938);
and U387 (N_387,In_488,In_787);
xnor U388 (N_388,In_55,In_105);
nand U389 (N_389,In_110,In_793);
xor U390 (N_390,In_770,In_515);
or U391 (N_391,In_220,In_230);
nand U392 (N_392,In_111,In_695);
and U393 (N_393,In_865,In_765);
and U394 (N_394,In_548,In_949);
nand U395 (N_395,In_860,In_503);
xnor U396 (N_396,In_298,In_818);
xor U397 (N_397,In_843,In_45);
or U398 (N_398,In_117,In_586);
or U399 (N_399,In_265,In_123);
nand U400 (N_400,In_617,In_828);
nand U401 (N_401,In_249,In_139);
or U402 (N_402,In_974,In_813);
and U403 (N_403,In_947,In_996);
and U404 (N_404,In_431,In_144);
or U405 (N_405,In_156,In_840);
or U406 (N_406,In_718,In_564);
and U407 (N_407,In_369,In_382);
and U408 (N_408,In_526,In_622);
nand U409 (N_409,In_125,In_244);
or U410 (N_410,In_815,In_946);
nor U411 (N_411,In_83,In_833);
and U412 (N_412,In_213,In_106);
xor U413 (N_413,In_669,In_204);
nor U414 (N_414,In_78,In_75);
nand U415 (N_415,In_773,In_542);
and U416 (N_416,In_91,In_165);
nor U417 (N_417,In_255,In_511);
xnor U418 (N_418,In_80,In_699);
and U419 (N_419,In_680,In_153);
and U420 (N_420,In_528,In_132);
nor U421 (N_421,In_411,In_707);
or U422 (N_422,In_450,In_758);
and U423 (N_423,In_620,In_544);
or U424 (N_424,In_311,In_826);
nor U425 (N_425,In_237,In_839);
nand U426 (N_426,In_624,In_36);
nand U427 (N_427,In_522,In_229);
nand U428 (N_428,In_802,In_780);
and U429 (N_429,In_508,In_862);
nor U430 (N_430,In_206,In_155);
nor U431 (N_431,In_457,In_988);
and U432 (N_432,In_920,In_147);
nor U433 (N_433,In_716,In_260);
nor U434 (N_434,In_646,In_386);
nor U435 (N_435,In_325,In_850);
or U436 (N_436,In_873,In_651);
nand U437 (N_437,In_479,In_294);
and U438 (N_438,In_162,In_878);
xor U439 (N_439,In_394,In_375);
nand U440 (N_440,In_486,In_874);
and U441 (N_441,In_668,In_340);
xor U442 (N_442,In_70,In_152);
nand U443 (N_443,In_61,In_232);
or U444 (N_444,In_845,In_759);
nand U445 (N_445,In_171,In_735);
nand U446 (N_446,In_993,In_84);
nand U447 (N_447,In_595,In_627);
xor U448 (N_448,In_428,In_893);
xnor U449 (N_449,In_811,In_983);
and U450 (N_450,In_667,In_320);
or U451 (N_451,In_245,In_982);
nand U452 (N_452,In_195,In_914);
and U453 (N_453,In_752,In_989);
nor U454 (N_454,In_456,In_673);
or U455 (N_455,In_200,In_505);
nor U456 (N_456,In_514,In_692);
and U457 (N_457,In_880,In_592);
and U458 (N_458,In_13,In_343);
or U459 (N_459,In_395,In_333);
nand U460 (N_460,In_432,In_533);
nor U461 (N_461,In_476,In_960);
xor U462 (N_462,In_413,In_597);
nor U463 (N_463,In_273,In_532);
nand U464 (N_464,In_591,In_552);
and U465 (N_465,In_225,In_250);
and U466 (N_466,In_527,In_373);
or U467 (N_467,In_402,In_638);
or U468 (N_468,In_679,In_94);
xor U469 (N_469,In_10,In_466);
nand U470 (N_470,In_922,In_754);
nand U471 (N_471,In_203,In_698);
or U472 (N_472,In_750,In_653);
and U473 (N_473,In_540,In_40);
xnor U474 (N_474,In_427,In_170);
nand U475 (N_475,In_774,In_978);
or U476 (N_476,In_794,In_473);
or U477 (N_477,In_869,In_279);
or U478 (N_478,In_877,In_71);
nor U479 (N_479,In_588,In_939);
and U480 (N_480,In_519,In_168);
nor U481 (N_481,In_782,In_96);
xnor U482 (N_482,In_188,In_4);
nor U483 (N_483,In_122,In_581);
xor U484 (N_484,In_352,In_501);
nor U485 (N_485,In_378,In_173);
and U486 (N_486,In_870,In_885);
and U487 (N_487,In_930,In_904);
nor U488 (N_488,In_924,In_258);
nor U489 (N_489,In_931,In_133);
or U490 (N_490,In_866,In_804);
nor U491 (N_491,In_602,In_742);
and U492 (N_492,In_711,In_81);
and U493 (N_493,In_708,In_756);
and U494 (N_494,In_521,In_485);
and U495 (N_495,In_909,In_573);
and U496 (N_496,In_722,In_995);
xor U497 (N_497,In_629,In_829);
nor U498 (N_498,In_293,In_483);
and U499 (N_499,In_998,In_401);
and U500 (N_500,In_269,In_560);
nor U501 (N_501,In_160,In_413);
or U502 (N_502,In_48,In_284);
xnor U503 (N_503,In_941,In_291);
nand U504 (N_504,In_730,In_900);
or U505 (N_505,In_186,In_164);
and U506 (N_506,In_590,In_63);
nand U507 (N_507,In_9,In_426);
nand U508 (N_508,In_221,In_963);
xnor U509 (N_509,In_796,In_49);
nor U510 (N_510,In_425,In_531);
or U511 (N_511,In_81,In_458);
or U512 (N_512,In_906,In_817);
nor U513 (N_513,In_482,In_616);
nand U514 (N_514,In_650,In_997);
or U515 (N_515,In_861,In_382);
xnor U516 (N_516,In_976,In_300);
or U517 (N_517,In_612,In_891);
and U518 (N_518,In_165,In_445);
nand U519 (N_519,In_959,In_199);
nor U520 (N_520,In_712,In_90);
or U521 (N_521,In_594,In_567);
xor U522 (N_522,In_202,In_644);
nand U523 (N_523,In_102,In_581);
xor U524 (N_524,In_121,In_849);
nor U525 (N_525,In_555,In_773);
xnor U526 (N_526,In_548,In_295);
xnor U527 (N_527,In_928,In_320);
nor U528 (N_528,In_997,In_430);
nand U529 (N_529,In_151,In_866);
or U530 (N_530,In_2,In_566);
nor U531 (N_531,In_618,In_83);
nor U532 (N_532,In_109,In_909);
nor U533 (N_533,In_327,In_351);
or U534 (N_534,In_67,In_825);
or U535 (N_535,In_579,In_591);
nor U536 (N_536,In_95,In_544);
or U537 (N_537,In_632,In_695);
nor U538 (N_538,In_239,In_334);
nand U539 (N_539,In_92,In_708);
or U540 (N_540,In_922,In_716);
nand U541 (N_541,In_281,In_752);
nand U542 (N_542,In_241,In_562);
and U543 (N_543,In_345,In_436);
nand U544 (N_544,In_472,In_638);
xnor U545 (N_545,In_769,In_608);
xor U546 (N_546,In_139,In_752);
and U547 (N_547,In_530,In_858);
xor U548 (N_548,In_579,In_578);
or U549 (N_549,In_74,In_809);
xnor U550 (N_550,In_59,In_82);
nand U551 (N_551,In_240,In_41);
nand U552 (N_552,In_466,In_212);
or U553 (N_553,In_623,In_358);
nor U554 (N_554,In_35,In_165);
or U555 (N_555,In_975,In_517);
nor U556 (N_556,In_226,In_815);
nand U557 (N_557,In_703,In_423);
nor U558 (N_558,In_79,In_99);
nor U559 (N_559,In_250,In_578);
and U560 (N_560,In_543,In_594);
or U561 (N_561,In_772,In_582);
nor U562 (N_562,In_577,In_760);
nor U563 (N_563,In_389,In_716);
nand U564 (N_564,In_816,In_536);
and U565 (N_565,In_18,In_896);
nor U566 (N_566,In_692,In_393);
and U567 (N_567,In_717,In_484);
and U568 (N_568,In_303,In_429);
nand U569 (N_569,In_541,In_942);
xnor U570 (N_570,In_956,In_914);
or U571 (N_571,In_395,In_621);
nor U572 (N_572,In_842,In_221);
nand U573 (N_573,In_532,In_628);
nand U574 (N_574,In_51,In_172);
and U575 (N_575,In_378,In_282);
or U576 (N_576,In_810,In_749);
xor U577 (N_577,In_905,In_529);
and U578 (N_578,In_55,In_799);
or U579 (N_579,In_831,In_944);
or U580 (N_580,In_914,In_708);
or U581 (N_581,In_7,In_916);
or U582 (N_582,In_283,In_227);
and U583 (N_583,In_55,In_18);
and U584 (N_584,In_892,In_361);
nand U585 (N_585,In_858,In_701);
or U586 (N_586,In_281,In_915);
xor U587 (N_587,In_919,In_813);
nand U588 (N_588,In_858,In_550);
or U589 (N_589,In_585,In_836);
or U590 (N_590,In_586,In_615);
or U591 (N_591,In_407,In_162);
or U592 (N_592,In_82,In_259);
nor U593 (N_593,In_84,In_665);
nand U594 (N_594,In_612,In_488);
nand U595 (N_595,In_201,In_493);
xor U596 (N_596,In_352,In_823);
nand U597 (N_597,In_105,In_651);
xnor U598 (N_598,In_6,In_586);
xor U599 (N_599,In_854,In_595);
or U600 (N_600,In_380,In_929);
nand U601 (N_601,In_338,In_354);
and U602 (N_602,In_738,In_639);
xnor U603 (N_603,In_251,In_300);
nand U604 (N_604,In_328,In_653);
nor U605 (N_605,In_86,In_295);
nor U606 (N_606,In_491,In_974);
nand U607 (N_607,In_550,In_868);
xnor U608 (N_608,In_259,In_806);
nor U609 (N_609,In_406,In_276);
xnor U610 (N_610,In_7,In_141);
or U611 (N_611,In_48,In_218);
nor U612 (N_612,In_307,In_124);
nor U613 (N_613,In_388,In_475);
and U614 (N_614,In_187,In_175);
or U615 (N_615,In_644,In_307);
or U616 (N_616,In_265,In_473);
and U617 (N_617,In_335,In_979);
and U618 (N_618,In_695,In_840);
nor U619 (N_619,In_990,In_101);
nor U620 (N_620,In_196,In_699);
nand U621 (N_621,In_387,In_274);
and U622 (N_622,In_522,In_976);
or U623 (N_623,In_95,In_174);
nor U624 (N_624,In_55,In_874);
or U625 (N_625,In_717,In_463);
or U626 (N_626,In_198,In_14);
nand U627 (N_627,In_954,In_23);
and U628 (N_628,In_383,In_998);
nand U629 (N_629,In_673,In_877);
or U630 (N_630,In_889,In_485);
nor U631 (N_631,In_915,In_257);
nor U632 (N_632,In_355,In_991);
nor U633 (N_633,In_22,In_655);
and U634 (N_634,In_517,In_175);
or U635 (N_635,In_514,In_348);
and U636 (N_636,In_825,In_565);
nor U637 (N_637,In_266,In_707);
and U638 (N_638,In_179,In_355);
nand U639 (N_639,In_209,In_908);
and U640 (N_640,In_953,In_274);
nor U641 (N_641,In_858,In_56);
nor U642 (N_642,In_908,In_314);
and U643 (N_643,In_527,In_589);
nor U644 (N_644,In_929,In_618);
nor U645 (N_645,In_964,In_469);
nand U646 (N_646,In_449,In_283);
nand U647 (N_647,In_631,In_687);
nor U648 (N_648,In_836,In_942);
or U649 (N_649,In_153,In_196);
xnor U650 (N_650,In_140,In_495);
or U651 (N_651,In_535,In_244);
and U652 (N_652,In_652,In_637);
and U653 (N_653,In_982,In_161);
xnor U654 (N_654,In_778,In_101);
nor U655 (N_655,In_531,In_495);
nand U656 (N_656,In_812,In_946);
nand U657 (N_657,In_359,In_629);
xnor U658 (N_658,In_381,In_914);
or U659 (N_659,In_244,In_614);
or U660 (N_660,In_38,In_754);
nand U661 (N_661,In_510,In_305);
or U662 (N_662,In_204,In_135);
nand U663 (N_663,In_915,In_814);
nor U664 (N_664,In_804,In_661);
and U665 (N_665,In_114,In_964);
nor U666 (N_666,In_538,In_143);
nand U667 (N_667,In_378,In_369);
nor U668 (N_668,In_565,In_976);
nand U669 (N_669,In_772,In_272);
nor U670 (N_670,In_993,In_139);
nor U671 (N_671,In_176,In_279);
xnor U672 (N_672,In_777,In_149);
or U673 (N_673,In_208,In_536);
nor U674 (N_674,In_226,In_472);
or U675 (N_675,In_352,In_378);
nand U676 (N_676,In_255,In_505);
nand U677 (N_677,In_334,In_237);
nor U678 (N_678,In_906,In_437);
xnor U679 (N_679,In_484,In_40);
nand U680 (N_680,In_773,In_406);
or U681 (N_681,In_851,In_369);
or U682 (N_682,In_840,In_87);
nor U683 (N_683,In_899,In_303);
nor U684 (N_684,In_54,In_561);
nand U685 (N_685,In_723,In_802);
or U686 (N_686,In_589,In_677);
nor U687 (N_687,In_144,In_735);
xor U688 (N_688,In_185,In_232);
xnor U689 (N_689,In_161,In_206);
nor U690 (N_690,In_460,In_683);
xnor U691 (N_691,In_939,In_910);
nand U692 (N_692,In_613,In_864);
nor U693 (N_693,In_967,In_741);
or U694 (N_694,In_995,In_720);
nand U695 (N_695,In_398,In_599);
nor U696 (N_696,In_391,In_569);
or U697 (N_697,In_462,In_725);
and U698 (N_698,In_815,In_8);
or U699 (N_699,In_389,In_122);
nor U700 (N_700,In_3,In_402);
and U701 (N_701,In_442,In_74);
or U702 (N_702,In_817,In_752);
nor U703 (N_703,In_499,In_916);
nor U704 (N_704,In_189,In_790);
or U705 (N_705,In_503,In_881);
nor U706 (N_706,In_748,In_772);
or U707 (N_707,In_636,In_716);
nand U708 (N_708,In_848,In_132);
or U709 (N_709,In_104,In_218);
and U710 (N_710,In_712,In_262);
and U711 (N_711,In_101,In_927);
and U712 (N_712,In_474,In_311);
nand U713 (N_713,In_530,In_344);
nand U714 (N_714,In_305,In_677);
xor U715 (N_715,In_314,In_395);
nor U716 (N_716,In_358,In_863);
xnor U717 (N_717,In_687,In_907);
nor U718 (N_718,In_162,In_206);
and U719 (N_719,In_197,In_666);
and U720 (N_720,In_720,In_569);
nand U721 (N_721,In_928,In_562);
nor U722 (N_722,In_419,In_318);
xnor U723 (N_723,In_259,In_466);
xnor U724 (N_724,In_945,In_433);
and U725 (N_725,In_259,In_464);
or U726 (N_726,In_704,In_926);
xor U727 (N_727,In_151,In_709);
or U728 (N_728,In_812,In_589);
and U729 (N_729,In_639,In_663);
xnor U730 (N_730,In_994,In_514);
and U731 (N_731,In_914,In_857);
or U732 (N_732,In_908,In_536);
or U733 (N_733,In_754,In_212);
or U734 (N_734,In_205,In_847);
and U735 (N_735,In_976,In_891);
nand U736 (N_736,In_884,In_13);
xor U737 (N_737,In_945,In_776);
or U738 (N_738,In_348,In_127);
nor U739 (N_739,In_772,In_353);
and U740 (N_740,In_986,In_751);
or U741 (N_741,In_469,In_23);
nor U742 (N_742,In_489,In_718);
nor U743 (N_743,In_436,In_693);
or U744 (N_744,In_775,In_126);
nand U745 (N_745,In_40,In_432);
nand U746 (N_746,In_92,In_69);
or U747 (N_747,In_458,In_926);
nand U748 (N_748,In_778,In_675);
and U749 (N_749,In_435,In_344);
and U750 (N_750,In_333,In_185);
xnor U751 (N_751,In_538,In_216);
nor U752 (N_752,In_589,In_772);
and U753 (N_753,In_435,In_746);
or U754 (N_754,In_692,In_783);
or U755 (N_755,In_940,In_902);
nor U756 (N_756,In_309,In_986);
xnor U757 (N_757,In_59,In_47);
or U758 (N_758,In_586,In_317);
nand U759 (N_759,In_350,In_252);
xor U760 (N_760,In_121,In_921);
or U761 (N_761,In_597,In_667);
nor U762 (N_762,In_962,In_530);
and U763 (N_763,In_649,In_8);
xor U764 (N_764,In_371,In_158);
and U765 (N_765,In_686,In_159);
nand U766 (N_766,In_148,In_744);
or U767 (N_767,In_228,In_877);
nand U768 (N_768,In_664,In_252);
nor U769 (N_769,In_112,In_474);
and U770 (N_770,In_27,In_159);
nand U771 (N_771,In_921,In_12);
nand U772 (N_772,In_591,In_301);
nand U773 (N_773,In_285,In_427);
or U774 (N_774,In_249,In_686);
or U775 (N_775,In_340,In_732);
nand U776 (N_776,In_355,In_405);
and U777 (N_777,In_552,In_43);
xnor U778 (N_778,In_98,In_872);
and U779 (N_779,In_201,In_613);
or U780 (N_780,In_614,In_77);
xnor U781 (N_781,In_325,In_833);
and U782 (N_782,In_515,In_180);
xnor U783 (N_783,In_58,In_307);
and U784 (N_784,In_909,In_117);
xor U785 (N_785,In_936,In_573);
xnor U786 (N_786,In_59,In_254);
and U787 (N_787,In_985,In_203);
xor U788 (N_788,In_726,In_783);
nand U789 (N_789,In_432,In_337);
and U790 (N_790,In_387,In_691);
xor U791 (N_791,In_429,In_243);
or U792 (N_792,In_69,In_283);
or U793 (N_793,In_993,In_677);
or U794 (N_794,In_891,In_654);
and U795 (N_795,In_527,In_501);
xor U796 (N_796,In_898,In_501);
xor U797 (N_797,In_158,In_944);
and U798 (N_798,In_670,In_219);
xnor U799 (N_799,In_717,In_41);
xnor U800 (N_800,In_353,In_771);
nand U801 (N_801,In_676,In_428);
and U802 (N_802,In_160,In_40);
nor U803 (N_803,In_396,In_405);
or U804 (N_804,In_516,In_884);
and U805 (N_805,In_914,In_784);
or U806 (N_806,In_503,In_83);
nor U807 (N_807,In_880,In_850);
and U808 (N_808,In_750,In_858);
or U809 (N_809,In_905,In_857);
or U810 (N_810,In_178,In_10);
xnor U811 (N_811,In_499,In_244);
xor U812 (N_812,In_576,In_747);
xnor U813 (N_813,In_777,In_702);
nor U814 (N_814,In_827,In_383);
xnor U815 (N_815,In_46,In_249);
xnor U816 (N_816,In_667,In_770);
and U817 (N_817,In_75,In_434);
nand U818 (N_818,In_885,In_522);
nand U819 (N_819,In_936,In_252);
and U820 (N_820,In_805,In_745);
or U821 (N_821,In_723,In_149);
or U822 (N_822,In_367,In_473);
or U823 (N_823,In_404,In_383);
nor U824 (N_824,In_829,In_875);
and U825 (N_825,In_420,In_94);
nor U826 (N_826,In_382,In_43);
nor U827 (N_827,In_183,In_823);
and U828 (N_828,In_357,In_359);
xor U829 (N_829,In_904,In_831);
nor U830 (N_830,In_216,In_582);
or U831 (N_831,In_762,In_183);
and U832 (N_832,In_129,In_800);
and U833 (N_833,In_15,In_96);
nor U834 (N_834,In_251,In_774);
nor U835 (N_835,In_957,In_352);
xnor U836 (N_836,In_341,In_955);
nor U837 (N_837,In_44,In_453);
or U838 (N_838,In_135,In_39);
or U839 (N_839,In_991,In_771);
or U840 (N_840,In_380,In_595);
and U841 (N_841,In_737,In_593);
xnor U842 (N_842,In_782,In_601);
nor U843 (N_843,In_905,In_988);
xnor U844 (N_844,In_271,In_448);
nand U845 (N_845,In_852,In_72);
or U846 (N_846,In_575,In_867);
and U847 (N_847,In_914,In_910);
nand U848 (N_848,In_605,In_984);
and U849 (N_849,In_655,In_626);
and U850 (N_850,In_297,In_112);
and U851 (N_851,In_47,In_209);
nor U852 (N_852,In_647,In_653);
or U853 (N_853,In_613,In_0);
nand U854 (N_854,In_989,In_784);
and U855 (N_855,In_524,In_782);
xnor U856 (N_856,In_663,In_736);
and U857 (N_857,In_419,In_380);
nand U858 (N_858,In_197,In_251);
or U859 (N_859,In_14,In_824);
nor U860 (N_860,In_805,In_581);
nand U861 (N_861,In_421,In_654);
xnor U862 (N_862,In_588,In_148);
xnor U863 (N_863,In_362,In_296);
nand U864 (N_864,In_641,In_915);
nand U865 (N_865,In_95,In_482);
and U866 (N_866,In_176,In_641);
or U867 (N_867,In_667,In_634);
nand U868 (N_868,In_140,In_589);
nor U869 (N_869,In_522,In_397);
and U870 (N_870,In_480,In_503);
xnor U871 (N_871,In_460,In_23);
or U872 (N_872,In_506,In_303);
or U873 (N_873,In_236,In_182);
nor U874 (N_874,In_352,In_89);
xor U875 (N_875,In_829,In_624);
or U876 (N_876,In_780,In_713);
nor U877 (N_877,In_315,In_200);
and U878 (N_878,In_9,In_990);
nor U879 (N_879,In_222,In_549);
nor U880 (N_880,In_47,In_281);
nand U881 (N_881,In_244,In_188);
xor U882 (N_882,In_59,In_488);
or U883 (N_883,In_887,In_252);
or U884 (N_884,In_536,In_405);
xnor U885 (N_885,In_335,In_791);
or U886 (N_886,In_482,In_489);
nor U887 (N_887,In_877,In_560);
nand U888 (N_888,In_74,In_249);
xor U889 (N_889,In_450,In_109);
xor U890 (N_890,In_939,In_535);
or U891 (N_891,In_891,In_58);
or U892 (N_892,In_650,In_946);
and U893 (N_893,In_452,In_933);
and U894 (N_894,In_912,In_161);
or U895 (N_895,In_7,In_980);
or U896 (N_896,In_52,In_788);
xor U897 (N_897,In_335,In_948);
nor U898 (N_898,In_756,In_420);
nor U899 (N_899,In_35,In_445);
nor U900 (N_900,In_721,In_100);
nand U901 (N_901,In_534,In_767);
and U902 (N_902,In_994,In_473);
nor U903 (N_903,In_337,In_540);
nor U904 (N_904,In_310,In_743);
or U905 (N_905,In_751,In_434);
nand U906 (N_906,In_109,In_732);
or U907 (N_907,In_422,In_932);
xor U908 (N_908,In_104,In_8);
and U909 (N_909,In_461,In_135);
or U910 (N_910,In_557,In_366);
xnor U911 (N_911,In_191,In_643);
or U912 (N_912,In_10,In_111);
nor U913 (N_913,In_506,In_243);
nand U914 (N_914,In_474,In_667);
xnor U915 (N_915,In_409,In_838);
and U916 (N_916,In_834,In_892);
or U917 (N_917,In_379,In_555);
nand U918 (N_918,In_483,In_809);
nor U919 (N_919,In_279,In_77);
nor U920 (N_920,In_791,In_103);
and U921 (N_921,In_42,In_402);
xnor U922 (N_922,In_133,In_614);
nand U923 (N_923,In_522,In_655);
and U924 (N_924,In_493,In_618);
or U925 (N_925,In_461,In_296);
xnor U926 (N_926,In_918,In_93);
xnor U927 (N_927,In_47,In_900);
nand U928 (N_928,In_652,In_773);
nor U929 (N_929,In_731,In_374);
nor U930 (N_930,In_83,In_653);
nor U931 (N_931,In_258,In_842);
or U932 (N_932,In_766,In_351);
nand U933 (N_933,In_584,In_772);
xnor U934 (N_934,In_162,In_872);
nor U935 (N_935,In_210,In_764);
xnor U936 (N_936,In_882,In_704);
xnor U937 (N_937,In_624,In_590);
nor U938 (N_938,In_708,In_477);
and U939 (N_939,In_80,In_163);
or U940 (N_940,In_194,In_933);
xnor U941 (N_941,In_798,In_204);
and U942 (N_942,In_640,In_860);
xnor U943 (N_943,In_152,In_900);
nor U944 (N_944,In_165,In_659);
or U945 (N_945,In_574,In_918);
nand U946 (N_946,In_7,In_22);
and U947 (N_947,In_982,In_87);
or U948 (N_948,In_963,In_582);
nor U949 (N_949,In_287,In_796);
or U950 (N_950,In_750,In_949);
nor U951 (N_951,In_329,In_470);
xor U952 (N_952,In_167,In_658);
or U953 (N_953,In_839,In_888);
and U954 (N_954,In_2,In_466);
and U955 (N_955,In_352,In_413);
nand U956 (N_956,In_368,In_80);
nor U957 (N_957,In_387,In_266);
nand U958 (N_958,In_2,In_667);
nor U959 (N_959,In_643,In_575);
nor U960 (N_960,In_762,In_363);
xor U961 (N_961,In_208,In_32);
nor U962 (N_962,In_482,In_220);
nor U963 (N_963,In_457,In_950);
nand U964 (N_964,In_608,In_425);
and U965 (N_965,In_417,In_214);
or U966 (N_966,In_450,In_479);
xor U967 (N_967,In_978,In_474);
or U968 (N_968,In_941,In_925);
and U969 (N_969,In_402,In_543);
or U970 (N_970,In_746,In_206);
or U971 (N_971,In_403,In_742);
xor U972 (N_972,In_148,In_703);
and U973 (N_973,In_210,In_292);
xor U974 (N_974,In_420,In_634);
xor U975 (N_975,In_939,In_242);
nand U976 (N_976,In_80,In_831);
or U977 (N_977,In_383,In_78);
nor U978 (N_978,In_833,In_706);
and U979 (N_979,In_758,In_40);
nand U980 (N_980,In_891,In_576);
xnor U981 (N_981,In_367,In_848);
or U982 (N_982,In_279,In_718);
nor U983 (N_983,In_825,In_403);
and U984 (N_984,In_82,In_175);
or U985 (N_985,In_228,In_137);
nor U986 (N_986,In_351,In_9);
nand U987 (N_987,In_563,In_414);
nand U988 (N_988,In_520,In_344);
nand U989 (N_989,In_13,In_782);
nand U990 (N_990,In_250,In_25);
nand U991 (N_991,In_403,In_293);
nor U992 (N_992,In_536,In_476);
or U993 (N_993,In_617,In_78);
or U994 (N_994,In_986,In_792);
xor U995 (N_995,In_335,In_190);
xor U996 (N_996,In_540,In_759);
nor U997 (N_997,In_946,In_559);
nand U998 (N_998,In_318,In_632);
or U999 (N_999,In_154,In_801);
nor U1000 (N_1000,In_838,In_902);
nor U1001 (N_1001,In_876,In_370);
and U1002 (N_1002,In_624,In_791);
xor U1003 (N_1003,In_73,In_252);
nor U1004 (N_1004,In_534,In_552);
nor U1005 (N_1005,In_183,In_794);
and U1006 (N_1006,In_629,In_706);
and U1007 (N_1007,In_698,In_562);
and U1008 (N_1008,In_822,In_462);
and U1009 (N_1009,In_963,In_544);
nand U1010 (N_1010,In_57,In_968);
and U1011 (N_1011,In_904,In_606);
or U1012 (N_1012,In_342,In_173);
xnor U1013 (N_1013,In_101,In_807);
or U1014 (N_1014,In_955,In_645);
nand U1015 (N_1015,In_815,In_267);
and U1016 (N_1016,In_647,In_472);
nor U1017 (N_1017,In_200,In_876);
nor U1018 (N_1018,In_649,In_462);
nor U1019 (N_1019,In_257,In_32);
nor U1020 (N_1020,In_328,In_171);
or U1021 (N_1021,In_81,In_21);
or U1022 (N_1022,In_65,In_304);
or U1023 (N_1023,In_785,In_650);
nand U1024 (N_1024,In_986,In_777);
and U1025 (N_1025,In_303,In_662);
nand U1026 (N_1026,In_389,In_762);
and U1027 (N_1027,In_731,In_139);
or U1028 (N_1028,In_47,In_989);
nor U1029 (N_1029,In_142,In_712);
nand U1030 (N_1030,In_114,In_547);
nand U1031 (N_1031,In_631,In_831);
nor U1032 (N_1032,In_313,In_67);
nor U1033 (N_1033,In_878,In_747);
nand U1034 (N_1034,In_914,In_999);
or U1035 (N_1035,In_193,In_964);
xor U1036 (N_1036,In_74,In_398);
or U1037 (N_1037,In_29,In_706);
nor U1038 (N_1038,In_61,In_655);
or U1039 (N_1039,In_815,In_487);
nor U1040 (N_1040,In_677,In_905);
nor U1041 (N_1041,In_540,In_279);
nor U1042 (N_1042,In_423,In_979);
xnor U1043 (N_1043,In_586,In_291);
or U1044 (N_1044,In_167,In_223);
or U1045 (N_1045,In_812,In_713);
and U1046 (N_1046,In_913,In_674);
xnor U1047 (N_1047,In_138,In_256);
and U1048 (N_1048,In_315,In_233);
and U1049 (N_1049,In_201,In_944);
nor U1050 (N_1050,In_569,In_971);
nand U1051 (N_1051,In_967,In_366);
nor U1052 (N_1052,In_879,In_220);
nor U1053 (N_1053,In_204,In_159);
nand U1054 (N_1054,In_162,In_738);
or U1055 (N_1055,In_392,In_408);
and U1056 (N_1056,In_206,In_69);
xnor U1057 (N_1057,In_190,In_235);
nor U1058 (N_1058,In_854,In_630);
nand U1059 (N_1059,In_925,In_999);
nor U1060 (N_1060,In_526,In_120);
or U1061 (N_1061,In_517,In_192);
nor U1062 (N_1062,In_897,In_354);
nor U1063 (N_1063,In_18,In_124);
or U1064 (N_1064,In_159,In_120);
or U1065 (N_1065,In_310,In_252);
nor U1066 (N_1066,In_832,In_322);
or U1067 (N_1067,In_941,In_721);
nand U1068 (N_1068,In_391,In_351);
nor U1069 (N_1069,In_912,In_867);
nand U1070 (N_1070,In_914,In_580);
or U1071 (N_1071,In_406,In_497);
or U1072 (N_1072,In_988,In_296);
xnor U1073 (N_1073,In_163,In_842);
nand U1074 (N_1074,In_828,In_971);
nand U1075 (N_1075,In_61,In_528);
xor U1076 (N_1076,In_711,In_488);
nor U1077 (N_1077,In_703,In_953);
nand U1078 (N_1078,In_310,In_42);
nand U1079 (N_1079,In_522,In_247);
nand U1080 (N_1080,In_152,In_219);
nand U1081 (N_1081,In_405,In_673);
nor U1082 (N_1082,In_549,In_59);
or U1083 (N_1083,In_505,In_214);
nand U1084 (N_1084,In_841,In_401);
nor U1085 (N_1085,In_397,In_528);
or U1086 (N_1086,In_280,In_589);
or U1087 (N_1087,In_438,In_443);
and U1088 (N_1088,In_907,In_37);
or U1089 (N_1089,In_129,In_782);
or U1090 (N_1090,In_144,In_335);
nor U1091 (N_1091,In_416,In_664);
nor U1092 (N_1092,In_616,In_575);
xor U1093 (N_1093,In_338,In_138);
or U1094 (N_1094,In_301,In_603);
or U1095 (N_1095,In_216,In_847);
nor U1096 (N_1096,In_517,In_234);
or U1097 (N_1097,In_618,In_478);
nor U1098 (N_1098,In_120,In_121);
or U1099 (N_1099,In_843,In_528);
or U1100 (N_1100,In_527,In_547);
nand U1101 (N_1101,In_505,In_37);
xnor U1102 (N_1102,In_87,In_147);
nor U1103 (N_1103,In_841,In_663);
and U1104 (N_1104,In_932,In_943);
and U1105 (N_1105,In_949,In_628);
xor U1106 (N_1106,In_779,In_164);
or U1107 (N_1107,In_374,In_507);
nor U1108 (N_1108,In_139,In_596);
nand U1109 (N_1109,In_620,In_626);
or U1110 (N_1110,In_23,In_961);
xnor U1111 (N_1111,In_128,In_721);
nand U1112 (N_1112,In_245,In_492);
xnor U1113 (N_1113,In_208,In_250);
nand U1114 (N_1114,In_861,In_843);
or U1115 (N_1115,In_887,In_149);
nand U1116 (N_1116,In_953,In_114);
xnor U1117 (N_1117,In_646,In_141);
nand U1118 (N_1118,In_435,In_768);
or U1119 (N_1119,In_915,In_709);
xor U1120 (N_1120,In_436,In_40);
nand U1121 (N_1121,In_522,In_234);
nor U1122 (N_1122,In_529,In_254);
xnor U1123 (N_1123,In_266,In_742);
nor U1124 (N_1124,In_573,In_51);
nand U1125 (N_1125,In_503,In_662);
nor U1126 (N_1126,In_598,In_10);
xnor U1127 (N_1127,In_658,In_57);
xnor U1128 (N_1128,In_401,In_622);
nor U1129 (N_1129,In_905,In_560);
nor U1130 (N_1130,In_560,In_824);
xnor U1131 (N_1131,In_517,In_28);
or U1132 (N_1132,In_345,In_648);
xnor U1133 (N_1133,In_422,In_678);
or U1134 (N_1134,In_519,In_882);
xnor U1135 (N_1135,In_630,In_206);
nor U1136 (N_1136,In_102,In_822);
or U1137 (N_1137,In_49,In_159);
and U1138 (N_1138,In_427,In_317);
or U1139 (N_1139,In_431,In_401);
xor U1140 (N_1140,In_41,In_763);
nand U1141 (N_1141,In_361,In_473);
or U1142 (N_1142,In_345,In_221);
and U1143 (N_1143,In_240,In_325);
xor U1144 (N_1144,In_186,In_415);
or U1145 (N_1145,In_431,In_967);
nand U1146 (N_1146,In_344,In_901);
nor U1147 (N_1147,In_920,In_118);
nor U1148 (N_1148,In_320,In_509);
nor U1149 (N_1149,In_465,In_412);
nor U1150 (N_1150,In_438,In_843);
nand U1151 (N_1151,In_198,In_233);
nor U1152 (N_1152,In_982,In_428);
nand U1153 (N_1153,In_616,In_314);
xnor U1154 (N_1154,In_565,In_188);
nand U1155 (N_1155,In_610,In_151);
or U1156 (N_1156,In_297,In_111);
nand U1157 (N_1157,In_985,In_767);
nand U1158 (N_1158,In_837,In_761);
or U1159 (N_1159,In_403,In_964);
and U1160 (N_1160,In_971,In_575);
or U1161 (N_1161,In_429,In_716);
or U1162 (N_1162,In_829,In_676);
or U1163 (N_1163,In_768,In_407);
nor U1164 (N_1164,In_226,In_640);
xnor U1165 (N_1165,In_514,In_946);
nand U1166 (N_1166,In_296,In_403);
or U1167 (N_1167,In_876,In_67);
and U1168 (N_1168,In_789,In_687);
nor U1169 (N_1169,In_951,In_532);
nor U1170 (N_1170,In_883,In_225);
or U1171 (N_1171,In_936,In_335);
and U1172 (N_1172,In_973,In_134);
and U1173 (N_1173,In_9,In_360);
and U1174 (N_1174,In_35,In_543);
and U1175 (N_1175,In_431,In_631);
and U1176 (N_1176,In_472,In_440);
and U1177 (N_1177,In_415,In_626);
nor U1178 (N_1178,In_791,In_797);
xnor U1179 (N_1179,In_678,In_378);
and U1180 (N_1180,In_406,In_807);
nor U1181 (N_1181,In_668,In_222);
and U1182 (N_1182,In_712,In_580);
and U1183 (N_1183,In_719,In_581);
xor U1184 (N_1184,In_560,In_551);
and U1185 (N_1185,In_58,In_858);
nor U1186 (N_1186,In_605,In_583);
and U1187 (N_1187,In_689,In_826);
nand U1188 (N_1188,In_220,In_136);
nor U1189 (N_1189,In_971,In_811);
and U1190 (N_1190,In_347,In_633);
nor U1191 (N_1191,In_930,In_685);
and U1192 (N_1192,In_629,In_500);
xnor U1193 (N_1193,In_86,In_834);
or U1194 (N_1194,In_713,In_813);
xor U1195 (N_1195,In_876,In_130);
and U1196 (N_1196,In_645,In_595);
nand U1197 (N_1197,In_687,In_778);
nand U1198 (N_1198,In_314,In_336);
nand U1199 (N_1199,In_640,In_775);
and U1200 (N_1200,In_415,In_525);
or U1201 (N_1201,In_211,In_1);
nand U1202 (N_1202,In_879,In_288);
and U1203 (N_1203,In_349,In_431);
and U1204 (N_1204,In_830,In_738);
xor U1205 (N_1205,In_446,In_430);
and U1206 (N_1206,In_853,In_114);
nor U1207 (N_1207,In_612,In_866);
nor U1208 (N_1208,In_605,In_219);
xor U1209 (N_1209,In_182,In_242);
nand U1210 (N_1210,In_228,In_170);
nand U1211 (N_1211,In_732,In_1);
or U1212 (N_1212,In_882,In_672);
nor U1213 (N_1213,In_779,In_385);
nor U1214 (N_1214,In_865,In_753);
or U1215 (N_1215,In_73,In_958);
nand U1216 (N_1216,In_105,In_284);
or U1217 (N_1217,In_179,In_875);
or U1218 (N_1218,In_893,In_978);
xor U1219 (N_1219,In_186,In_566);
and U1220 (N_1220,In_21,In_400);
or U1221 (N_1221,In_880,In_261);
xor U1222 (N_1222,In_183,In_855);
or U1223 (N_1223,In_936,In_742);
or U1224 (N_1224,In_478,In_415);
and U1225 (N_1225,In_589,In_430);
or U1226 (N_1226,In_821,In_713);
nand U1227 (N_1227,In_158,In_147);
nor U1228 (N_1228,In_484,In_69);
nand U1229 (N_1229,In_88,In_728);
nand U1230 (N_1230,In_227,In_7);
xor U1231 (N_1231,In_492,In_638);
or U1232 (N_1232,In_164,In_742);
or U1233 (N_1233,In_430,In_50);
nor U1234 (N_1234,In_231,In_452);
nand U1235 (N_1235,In_7,In_415);
nor U1236 (N_1236,In_506,In_886);
or U1237 (N_1237,In_443,In_554);
xnor U1238 (N_1238,In_487,In_491);
and U1239 (N_1239,In_655,In_705);
or U1240 (N_1240,In_6,In_925);
nand U1241 (N_1241,In_580,In_14);
and U1242 (N_1242,In_512,In_442);
nand U1243 (N_1243,In_854,In_817);
nand U1244 (N_1244,In_95,In_369);
or U1245 (N_1245,In_589,In_552);
or U1246 (N_1246,In_710,In_780);
nand U1247 (N_1247,In_796,In_953);
nor U1248 (N_1248,In_185,In_997);
xor U1249 (N_1249,In_448,In_845);
xor U1250 (N_1250,In_606,In_511);
xor U1251 (N_1251,In_127,In_208);
nor U1252 (N_1252,In_255,In_256);
or U1253 (N_1253,In_414,In_825);
xor U1254 (N_1254,In_443,In_159);
and U1255 (N_1255,In_172,In_809);
or U1256 (N_1256,In_450,In_206);
and U1257 (N_1257,In_719,In_867);
and U1258 (N_1258,In_139,In_694);
nor U1259 (N_1259,In_2,In_383);
or U1260 (N_1260,In_317,In_349);
xor U1261 (N_1261,In_979,In_918);
xnor U1262 (N_1262,In_944,In_907);
nor U1263 (N_1263,In_206,In_252);
xnor U1264 (N_1264,In_993,In_445);
xnor U1265 (N_1265,In_499,In_670);
nand U1266 (N_1266,In_811,In_200);
nand U1267 (N_1267,In_774,In_929);
and U1268 (N_1268,In_99,In_882);
and U1269 (N_1269,In_592,In_663);
and U1270 (N_1270,In_336,In_538);
xnor U1271 (N_1271,In_875,In_936);
and U1272 (N_1272,In_686,In_919);
nor U1273 (N_1273,In_661,In_680);
nor U1274 (N_1274,In_93,In_998);
nor U1275 (N_1275,In_135,In_877);
and U1276 (N_1276,In_101,In_276);
and U1277 (N_1277,In_317,In_251);
nand U1278 (N_1278,In_61,In_842);
and U1279 (N_1279,In_350,In_953);
or U1280 (N_1280,In_281,In_901);
or U1281 (N_1281,In_189,In_981);
xnor U1282 (N_1282,In_593,In_915);
nor U1283 (N_1283,In_572,In_760);
nor U1284 (N_1284,In_622,In_233);
xnor U1285 (N_1285,In_964,In_600);
and U1286 (N_1286,In_215,In_114);
and U1287 (N_1287,In_226,In_814);
and U1288 (N_1288,In_698,In_658);
nor U1289 (N_1289,In_294,In_203);
and U1290 (N_1290,In_576,In_18);
nand U1291 (N_1291,In_120,In_50);
xor U1292 (N_1292,In_999,In_184);
or U1293 (N_1293,In_965,In_411);
nand U1294 (N_1294,In_866,In_155);
xor U1295 (N_1295,In_645,In_708);
xor U1296 (N_1296,In_358,In_428);
nand U1297 (N_1297,In_291,In_795);
or U1298 (N_1298,In_681,In_428);
nand U1299 (N_1299,In_393,In_429);
xnor U1300 (N_1300,In_315,In_774);
xor U1301 (N_1301,In_659,In_830);
xor U1302 (N_1302,In_964,In_289);
xnor U1303 (N_1303,In_715,In_845);
xor U1304 (N_1304,In_9,In_378);
nand U1305 (N_1305,In_624,In_271);
nor U1306 (N_1306,In_557,In_797);
nand U1307 (N_1307,In_305,In_408);
and U1308 (N_1308,In_457,In_50);
nand U1309 (N_1309,In_450,In_935);
or U1310 (N_1310,In_144,In_58);
xnor U1311 (N_1311,In_364,In_633);
nor U1312 (N_1312,In_332,In_803);
xor U1313 (N_1313,In_995,In_981);
and U1314 (N_1314,In_644,In_326);
and U1315 (N_1315,In_66,In_489);
nand U1316 (N_1316,In_116,In_291);
nand U1317 (N_1317,In_636,In_129);
and U1318 (N_1318,In_270,In_970);
or U1319 (N_1319,In_965,In_63);
or U1320 (N_1320,In_723,In_846);
or U1321 (N_1321,In_935,In_770);
nand U1322 (N_1322,In_405,In_335);
nand U1323 (N_1323,In_892,In_408);
xnor U1324 (N_1324,In_847,In_128);
xnor U1325 (N_1325,In_592,In_530);
nand U1326 (N_1326,In_567,In_852);
nor U1327 (N_1327,In_759,In_409);
and U1328 (N_1328,In_785,In_656);
or U1329 (N_1329,In_373,In_54);
nand U1330 (N_1330,In_199,In_61);
nand U1331 (N_1331,In_141,In_403);
xnor U1332 (N_1332,In_853,In_461);
or U1333 (N_1333,In_670,In_899);
xnor U1334 (N_1334,In_998,In_841);
nor U1335 (N_1335,In_304,In_531);
xor U1336 (N_1336,In_703,In_100);
and U1337 (N_1337,In_118,In_460);
xor U1338 (N_1338,In_872,In_780);
and U1339 (N_1339,In_983,In_918);
and U1340 (N_1340,In_938,In_685);
and U1341 (N_1341,In_47,In_808);
nor U1342 (N_1342,In_623,In_677);
xnor U1343 (N_1343,In_610,In_15);
xor U1344 (N_1344,In_617,In_562);
nor U1345 (N_1345,In_558,In_223);
and U1346 (N_1346,In_116,In_743);
xor U1347 (N_1347,In_971,In_712);
or U1348 (N_1348,In_786,In_677);
or U1349 (N_1349,In_590,In_230);
nor U1350 (N_1350,In_264,In_474);
nor U1351 (N_1351,In_119,In_186);
or U1352 (N_1352,In_716,In_226);
or U1353 (N_1353,In_328,In_966);
nand U1354 (N_1354,In_489,In_492);
xnor U1355 (N_1355,In_932,In_424);
or U1356 (N_1356,In_932,In_761);
nor U1357 (N_1357,In_785,In_378);
xnor U1358 (N_1358,In_436,In_216);
nor U1359 (N_1359,In_92,In_453);
and U1360 (N_1360,In_231,In_577);
or U1361 (N_1361,In_627,In_817);
or U1362 (N_1362,In_149,In_844);
nand U1363 (N_1363,In_634,In_244);
nand U1364 (N_1364,In_258,In_291);
xnor U1365 (N_1365,In_768,In_51);
or U1366 (N_1366,In_843,In_746);
or U1367 (N_1367,In_364,In_844);
xor U1368 (N_1368,In_46,In_366);
nand U1369 (N_1369,In_603,In_969);
xnor U1370 (N_1370,In_948,In_857);
nand U1371 (N_1371,In_309,In_236);
and U1372 (N_1372,In_650,In_99);
or U1373 (N_1373,In_788,In_928);
nand U1374 (N_1374,In_372,In_654);
xor U1375 (N_1375,In_732,In_752);
or U1376 (N_1376,In_355,In_988);
nor U1377 (N_1377,In_257,In_142);
xor U1378 (N_1378,In_278,In_749);
or U1379 (N_1379,In_496,In_481);
nand U1380 (N_1380,In_420,In_833);
xor U1381 (N_1381,In_898,In_369);
nor U1382 (N_1382,In_489,In_491);
nor U1383 (N_1383,In_90,In_880);
nand U1384 (N_1384,In_422,In_960);
and U1385 (N_1385,In_903,In_69);
nand U1386 (N_1386,In_372,In_605);
nor U1387 (N_1387,In_880,In_692);
or U1388 (N_1388,In_391,In_284);
nor U1389 (N_1389,In_92,In_697);
and U1390 (N_1390,In_154,In_343);
and U1391 (N_1391,In_745,In_939);
and U1392 (N_1392,In_188,In_362);
and U1393 (N_1393,In_430,In_631);
nand U1394 (N_1394,In_905,In_137);
or U1395 (N_1395,In_534,In_944);
nor U1396 (N_1396,In_321,In_747);
and U1397 (N_1397,In_169,In_751);
xnor U1398 (N_1398,In_305,In_501);
or U1399 (N_1399,In_986,In_628);
nor U1400 (N_1400,In_506,In_902);
or U1401 (N_1401,In_282,In_415);
nand U1402 (N_1402,In_66,In_944);
nor U1403 (N_1403,In_401,In_131);
nand U1404 (N_1404,In_337,In_381);
nand U1405 (N_1405,In_913,In_500);
nand U1406 (N_1406,In_435,In_25);
and U1407 (N_1407,In_857,In_656);
nand U1408 (N_1408,In_513,In_569);
and U1409 (N_1409,In_340,In_10);
or U1410 (N_1410,In_824,In_458);
nand U1411 (N_1411,In_916,In_305);
and U1412 (N_1412,In_90,In_152);
nand U1413 (N_1413,In_324,In_653);
nor U1414 (N_1414,In_480,In_469);
or U1415 (N_1415,In_601,In_504);
xnor U1416 (N_1416,In_276,In_899);
or U1417 (N_1417,In_474,In_320);
or U1418 (N_1418,In_348,In_42);
or U1419 (N_1419,In_36,In_625);
nand U1420 (N_1420,In_378,In_19);
nor U1421 (N_1421,In_976,In_250);
xnor U1422 (N_1422,In_342,In_911);
nand U1423 (N_1423,In_876,In_113);
and U1424 (N_1424,In_398,In_581);
xnor U1425 (N_1425,In_335,In_963);
or U1426 (N_1426,In_69,In_953);
nand U1427 (N_1427,In_769,In_198);
or U1428 (N_1428,In_139,In_0);
nor U1429 (N_1429,In_452,In_696);
nand U1430 (N_1430,In_980,In_392);
nor U1431 (N_1431,In_485,In_947);
xor U1432 (N_1432,In_84,In_510);
and U1433 (N_1433,In_508,In_316);
xnor U1434 (N_1434,In_80,In_318);
and U1435 (N_1435,In_10,In_582);
nand U1436 (N_1436,In_641,In_971);
and U1437 (N_1437,In_203,In_261);
xnor U1438 (N_1438,In_804,In_988);
and U1439 (N_1439,In_855,In_354);
nor U1440 (N_1440,In_896,In_869);
nand U1441 (N_1441,In_9,In_147);
nor U1442 (N_1442,In_272,In_91);
xor U1443 (N_1443,In_449,In_908);
xnor U1444 (N_1444,In_205,In_778);
nor U1445 (N_1445,In_947,In_689);
and U1446 (N_1446,In_803,In_782);
nor U1447 (N_1447,In_872,In_993);
nor U1448 (N_1448,In_998,In_680);
xor U1449 (N_1449,In_518,In_630);
xor U1450 (N_1450,In_621,In_251);
and U1451 (N_1451,In_301,In_209);
and U1452 (N_1452,In_190,In_315);
xor U1453 (N_1453,In_815,In_24);
nand U1454 (N_1454,In_4,In_456);
nor U1455 (N_1455,In_94,In_854);
and U1456 (N_1456,In_465,In_366);
xor U1457 (N_1457,In_20,In_846);
and U1458 (N_1458,In_458,In_138);
nand U1459 (N_1459,In_631,In_256);
nor U1460 (N_1460,In_714,In_529);
nand U1461 (N_1461,In_6,In_469);
or U1462 (N_1462,In_514,In_762);
nor U1463 (N_1463,In_651,In_168);
xor U1464 (N_1464,In_216,In_975);
nor U1465 (N_1465,In_92,In_87);
and U1466 (N_1466,In_922,In_994);
nand U1467 (N_1467,In_278,In_190);
nand U1468 (N_1468,In_82,In_107);
and U1469 (N_1469,In_956,In_994);
or U1470 (N_1470,In_404,In_26);
nor U1471 (N_1471,In_500,In_384);
nor U1472 (N_1472,In_207,In_862);
nand U1473 (N_1473,In_507,In_950);
nor U1474 (N_1474,In_621,In_11);
or U1475 (N_1475,In_9,In_507);
and U1476 (N_1476,In_913,In_343);
nand U1477 (N_1477,In_605,In_474);
and U1478 (N_1478,In_195,In_729);
nand U1479 (N_1479,In_41,In_623);
xor U1480 (N_1480,In_708,In_431);
nand U1481 (N_1481,In_635,In_76);
or U1482 (N_1482,In_983,In_363);
and U1483 (N_1483,In_195,In_345);
xor U1484 (N_1484,In_802,In_712);
nor U1485 (N_1485,In_583,In_44);
nand U1486 (N_1486,In_854,In_179);
and U1487 (N_1487,In_697,In_483);
nand U1488 (N_1488,In_612,In_453);
and U1489 (N_1489,In_444,In_410);
nand U1490 (N_1490,In_113,In_798);
nand U1491 (N_1491,In_341,In_3);
xor U1492 (N_1492,In_915,In_219);
nor U1493 (N_1493,In_626,In_779);
nor U1494 (N_1494,In_786,In_876);
nand U1495 (N_1495,In_649,In_83);
or U1496 (N_1496,In_613,In_527);
or U1497 (N_1497,In_997,In_885);
or U1498 (N_1498,In_44,In_515);
nor U1499 (N_1499,In_985,In_42);
or U1500 (N_1500,In_796,In_339);
or U1501 (N_1501,In_496,In_686);
nand U1502 (N_1502,In_559,In_966);
or U1503 (N_1503,In_212,In_583);
or U1504 (N_1504,In_600,In_94);
nor U1505 (N_1505,In_28,In_877);
or U1506 (N_1506,In_181,In_74);
and U1507 (N_1507,In_665,In_469);
nand U1508 (N_1508,In_26,In_859);
or U1509 (N_1509,In_997,In_26);
or U1510 (N_1510,In_502,In_805);
xnor U1511 (N_1511,In_184,In_709);
and U1512 (N_1512,In_152,In_572);
xnor U1513 (N_1513,In_441,In_183);
or U1514 (N_1514,In_936,In_172);
nand U1515 (N_1515,In_886,In_317);
nor U1516 (N_1516,In_65,In_446);
or U1517 (N_1517,In_750,In_94);
nand U1518 (N_1518,In_69,In_442);
nand U1519 (N_1519,In_3,In_104);
or U1520 (N_1520,In_788,In_305);
xnor U1521 (N_1521,In_716,In_409);
nand U1522 (N_1522,In_780,In_26);
xnor U1523 (N_1523,In_622,In_798);
nor U1524 (N_1524,In_667,In_510);
nand U1525 (N_1525,In_803,In_699);
nand U1526 (N_1526,In_981,In_146);
nand U1527 (N_1527,In_807,In_455);
nand U1528 (N_1528,In_814,In_81);
and U1529 (N_1529,In_331,In_616);
xnor U1530 (N_1530,In_954,In_48);
and U1531 (N_1531,In_580,In_697);
or U1532 (N_1532,In_446,In_235);
xnor U1533 (N_1533,In_237,In_320);
xnor U1534 (N_1534,In_562,In_913);
and U1535 (N_1535,In_651,In_392);
nand U1536 (N_1536,In_741,In_799);
xnor U1537 (N_1537,In_681,In_278);
or U1538 (N_1538,In_306,In_823);
and U1539 (N_1539,In_321,In_648);
xnor U1540 (N_1540,In_61,In_305);
or U1541 (N_1541,In_883,In_956);
nor U1542 (N_1542,In_450,In_926);
nand U1543 (N_1543,In_35,In_714);
or U1544 (N_1544,In_258,In_502);
nand U1545 (N_1545,In_802,In_375);
nand U1546 (N_1546,In_790,In_549);
nand U1547 (N_1547,In_56,In_947);
nand U1548 (N_1548,In_660,In_578);
nor U1549 (N_1549,In_775,In_295);
and U1550 (N_1550,In_630,In_626);
or U1551 (N_1551,In_166,In_326);
or U1552 (N_1552,In_176,In_611);
nand U1553 (N_1553,In_650,In_950);
nor U1554 (N_1554,In_95,In_258);
nand U1555 (N_1555,In_764,In_562);
or U1556 (N_1556,In_606,In_22);
nor U1557 (N_1557,In_303,In_959);
xor U1558 (N_1558,In_264,In_800);
or U1559 (N_1559,In_100,In_930);
or U1560 (N_1560,In_66,In_528);
nor U1561 (N_1561,In_363,In_958);
nor U1562 (N_1562,In_200,In_606);
nor U1563 (N_1563,In_382,In_792);
xor U1564 (N_1564,In_852,In_397);
nor U1565 (N_1565,In_234,In_367);
nor U1566 (N_1566,In_796,In_827);
nand U1567 (N_1567,In_229,In_889);
xor U1568 (N_1568,In_171,In_476);
and U1569 (N_1569,In_733,In_750);
xor U1570 (N_1570,In_850,In_953);
or U1571 (N_1571,In_807,In_125);
and U1572 (N_1572,In_454,In_438);
and U1573 (N_1573,In_412,In_69);
and U1574 (N_1574,In_869,In_304);
xor U1575 (N_1575,In_636,In_386);
nand U1576 (N_1576,In_893,In_834);
nand U1577 (N_1577,In_323,In_591);
or U1578 (N_1578,In_12,In_555);
and U1579 (N_1579,In_132,In_282);
nor U1580 (N_1580,In_973,In_714);
or U1581 (N_1581,In_264,In_705);
or U1582 (N_1582,In_353,In_395);
and U1583 (N_1583,In_577,In_252);
xnor U1584 (N_1584,In_7,In_113);
xnor U1585 (N_1585,In_837,In_425);
or U1586 (N_1586,In_686,In_881);
nand U1587 (N_1587,In_193,In_892);
nor U1588 (N_1588,In_180,In_329);
and U1589 (N_1589,In_171,In_737);
or U1590 (N_1590,In_57,In_249);
nor U1591 (N_1591,In_344,In_535);
or U1592 (N_1592,In_365,In_166);
and U1593 (N_1593,In_548,In_727);
nor U1594 (N_1594,In_75,In_109);
or U1595 (N_1595,In_848,In_312);
and U1596 (N_1596,In_876,In_359);
xnor U1597 (N_1597,In_200,In_211);
xnor U1598 (N_1598,In_338,In_983);
xnor U1599 (N_1599,In_713,In_599);
and U1600 (N_1600,In_572,In_704);
xnor U1601 (N_1601,In_697,In_669);
nor U1602 (N_1602,In_96,In_568);
nor U1603 (N_1603,In_51,In_927);
or U1604 (N_1604,In_454,In_419);
or U1605 (N_1605,In_767,In_559);
and U1606 (N_1606,In_244,In_226);
xnor U1607 (N_1607,In_164,In_65);
or U1608 (N_1608,In_554,In_96);
nand U1609 (N_1609,In_150,In_981);
and U1610 (N_1610,In_746,In_127);
or U1611 (N_1611,In_918,In_911);
nand U1612 (N_1612,In_181,In_484);
or U1613 (N_1613,In_774,In_749);
or U1614 (N_1614,In_87,In_349);
xnor U1615 (N_1615,In_279,In_74);
or U1616 (N_1616,In_386,In_582);
nor U1617 (N_1617,In_801,In_483);
nand U1618 (N_1618,In_134,In_282);
or U1619 (N_1619,In_699,In_376);
nand U1620 (N_1620,In_43,In_149);
nand U1621 (N_1621,In_299,In_53);
and U1622 (N_1622,In_421,In_766);
xnor U1623 (N_1623,In_784,In_64);
or U1624 (N_1624,In_736,In_197);
nand U1625 (N_1625,In_418,In_868);
nor U1626 (N_1626,In_834,In_481);
nand U1627 (N_1627,In_689,In_5);
or U1628 (N_1628,In_971,In_775);
and U1629 (N_1629,In_549,In_693);
xnor U1630 (N_1630,In_450,In_133);
or U1631 (N_1631,In_131,In_952);
nand U1632 (N_1632,In_326,In_849);
xor U1633 (N_1633,In_305,In_656);
nor U1634 (N_1634,In_537,In_267);
xor U1635 (N_1635,In_845,In_495);
and U1636 (N_1636,In_359,In_889);
xor U1637 (N_1637,In_37,In_365);
or U1638 (N_1638,In_192,In_821);
xnor U1639 (N_1639,In_320,In_450);
xnor U1640 (N_1640,In_692,In_430);
xor U1641 (N_1641,In_118,In_209);
xnor U1642 (N_1642,In_471,In_845);
xor U1643 (N_1643,In_143,In_4);
or U1644 (N_1644,In_833,In_61);
xnor U1645 (N_1645,In_123,In_572);
and U1646 (N_1646,In_371,In_351);
or U1647 (N_1647,In_193,In_403);
or U1648 (N_1648,In_734,In_375);
nor U1649 (N_1649,In_272,In_257);
and U1650 (N_1650,In_142,In_447);
xnor U1651 (N_1651,In_760,In_122);
or U1652 (N_1652,In_862,In_987);
nand U1653 (N_1653,In_865,In_609);
nor U1654 (N_1654,In_651,In_998);
and U1655 (N_1655,In_802,In_68);
xor U1656 (N_1656,In_424,In_255);
xor U1657 (N_1657,In_73,In_68);
xor U1658 (N_1658,In_71,In_425);
xor U1659 (N_1659,In_849,In_310);
xnor U1660 (N_1660,In_955,In_262);
xor U1661 (N_1661,In_476,In_886);
nand U1662 (N_1662,In_420,In_636);
xor U1663 (N_1663,In_835,In_539);
or U1664 (N_1664,In_325,In_478);
xnor U1665 (N_1665,In_925,In_973);
and U1666 (N_1666,In_494,In_605);
xnor U1667 (N_1667,In_477,In_671);
nand U1668 (N_1668,In_63,In_817);
and U1669 (N_1669,In_935,In_700);
or U1670 (N_1670,In_623,In_508);
and U1671 (N_1671,In_341,In_838);
or U1672 (N_1672,In_44,In_780);
nor U1673 (N_1673,In_366,In_244);
and U1674 (N_1674,In_824,In_441);
nand U1675 (N_1675,In_35,In_342);
nor U1676 (N_1676,In_329,In_804);
nor U1677 (N_1677,In_813,In_97);
and U1678 (N_1678,In_877,In_747);
or U1679 (N_1679,In_600,In_331);
and U1680 (N_1680,In_799,In_320);
or U1681 (N_1681,In_920,In_728);
and U1682 (N_1682,In_430,In_985);
nor U1683 (N_1683,In_233,In_846);
xnor U1684 (N_1684,In_916,In_723);
nand U1685 (N_1685,In_601,In_958);
xnor U1686 (N_1686,In_102,In_199);
nand U1687 (N_1687,In_788,In_218);
and U1688 (N_1688,In_204,In_904);
and U1689 (N_1689,In_178,In_674);
or U1690 (N_1690,In_98,In_558);
nand U1691 (N_1691,In_72,In_328);
nor U1692 (N_1692,In_442,In_110);
xor U1693 (N_1693,In_845,In_959);
and U1694 (N_1694,In_854,In_485);
xnor U1695 (N_1695,In_983,In_797);
xor U1696 (N_1696,In_424,In_675);
or U1697 (N_1697,In_473,In_174);
nor U1698 (N_1698,In_29,In_175);
or U1699 (N_1699,In_23,In_816);
xor U1700 (N_1700,In_263,In_795);
and U1701 (N_1701,In_881,In_123);
and U1702 (N_1702,In_839,In_545);
nor U1703 (N_1703,In_431,In_862);
nor U1704 (N_1704,In_845,In_393);
xnor U1705 (N_1705,In_653,In_443);
xnor U1706 (N_1706,In_427,In_999);
nor U1707 (N_1707,In_568,In_938);
nor U1708 (N_1708,In_514,In_209);
nor U1709 (N_1709,In_221,In_494);
xnor U1710 (N_1710,In_884,In_499);
xor U1711 (N_1711,In_490,In_293);
and U1712 (N_1712,In_25,In_593);
or U1713 (N_1713,In_270,In_547);
nor U1714 (N_1714,In_546,In_584);
or U1715 (N_1715,In_239,In_221);
and U1716 (N_1716,In_64,In_32);
xnor U1717 (N_1717,In_389,In_463);
and U1718 (N_1718,In_838,In_512);
xnor U1719 (N_1719,In_261,In_702);
or U1720 (N_1720,In_855,In_783);
nor U1721 (N_1721,In_581,In_35);
nor U1722 (N_1722,In_242,In_687);
or U1723 (N_1723,In_268,In_773);
xor U1724 (N_1724,In_963,In_951);
xnor U1725 (N_1725,In_46,In_713);
xnor U1726 (N_1726,In_309,In_311);
or U1727 (N_1727,In_166,In_193);
or U1728 (N_1728,In_640,In_100);
and U1729 (N_1729,In_661,In_892);
nor U1730 (N_1730,In_541,In_430);
nor U1731 (N_1731,In_489,In_696);
xor U1732 (N_1732,In_783,In_944);
and U1733 (N_1733,In_54,In_322);
nor U1734 (N_1734,In_399,In_978);
nand U1735 (N_1735,In_111,In_153);
xor U1736 (N_1736,In_108,In_102);
nand U1737 (N_1737,In_779,In_19);
xor U1738 (N_1738,In_697,In_670);
xor U1739 (N_1739,In_12,In_696);
xnor U1740 (N_1740,In_404,In_778);
nor U1741 (N_1741,In_277,In_383);
nand U1742 (N_1742,In_656,In_468);
and U1743 (N_1743,In_947,In_644);
nand U1744 (N_1744,In_623,In_436);
nor U1745 (N_1745,In_841,In_945);
or U1746 (N_1746,In_684,In_662);
or U1747 (N_1747,In_797,In_724);
and U1748 (N_1748,In_829,In_907);
nor U1749 (N_1749,In_169,In_587);
or U1750 (N_1750,In_363,In_393);
nand U1751 (N_1751,In_202,In_614);
nand U1752 (N_1752,In_657,In_561);
xor U1753 (N_1753,In_68,In_107);
nand U1754 (N_1754,In_202,In_950);
nand U1755 (N_1755,In_351,In_626);
and U1756 (N_1756,In_621,In_222);
and U1757 (N_1757,In_648,In_758);
nor U1758 (N_1758,In_191,In_436);
and U1759 (N_1759,In_326,In_433);
nor U1760 (N_1760,In_752,In_489);
nor U1761 (N_1761,In_119,In_919);
and U1762 (N_1762,In_174,In_432);
xnor U1763 (N_1763,In_622,In_366);
nand U1764 (N_1764,In_772,In_655);
and U1765 (N_1765,In_475,In_778);
and U1766 (N_1766,In_528,In_233);
nand U1767 (N_1767,In_360,In_609);
nand U1768 (N_1768,In_969,In_564);
or U1769 (N_1769,In_621,In_527);
nand U1770 (N_1770,In_158,In_75);
xnor U1771 (N_1771,In_512,In_533);
nor U1772 (N_1772,In_179,In_346);
or U1773 (N_1773,In_794,In_379);
nor U1774 (N_1774,In_116,In_687);
nor U1775 (N_1775,In_154,In_526);
nand U1776 (N_1776,In_29,In_177);
nor U1777 (N_1777,In_360,In_512);
nand U1778 (N_1778,In_701,In_806);
xor U1779 (N_1779,In_283,In_309);
or U1780 (N_1780,In_703,In_277);
nor U1781 (N_1781,In_68,In_859);
nor U1782 (N_1782,In_265,In_861);
xnor U1783 (N_1783,In_366,In_159);
and U1784 (N_1784,In_332,In_340);
xor U1785 (N_1785,In_431,In_655);
nand U1786 (N_1786,In_234,In_192);
nand U1787 (N_1787,In_461,In_90);
nor U1788 (N_1788,In_579,In_133);
or U1789 (N_1789,In_910,In_778);
nand U1790 (N_1790,In_586,In_680);
nor U1791 (N_1791,In_127,In_506);
and U1792 (N_1792,In_882,In_741);
and U1793 (N_1793,In_797,In_195);
or U1794 (N_1794,In_598,In_545);
and U1795 (N_1795,In_89,In_182);
nand U1796 (N_1796,In_834,In_297);
or U1797 (N_1797,In_666,In_488);
or U1798 (N_1798,In_956,In_696);
nand U1799 (N_1799,In_810,In_23);
and U1800 (N_1800,In_434,In_606);
xnor U1801 (N_1801,In_286,In_438);
and U1802 (N_1802,In_614,In_771);
and U1803 (N_1803,In_532,In_851);
or U1804 (N_1804,In_781,In_961);
or U1805 (N_1805,In_680,In_865);
nand U1806 (N_1806,In_194,In_903);
or U1807 (N_1807,In_409,In_7);
nor U1808 (N_1808,In_95,In_429);
and U1809 (N_1809,In_360,In_778);
or U1810 (N_1810,In_414,In_779);
nand U1811 (N_1811,In_484,In_186);
nor U1812 (N_1812,In_588,In_5);
xor U1813 (N_1813,In_579,In_258);
xor U1814 (N_1814,In_919,In_903);
or U1815 (N_1815,In_966,In_541);
nor U1816 (N_1816,In_243,In_777);
nand U1817 (N_1817,In_499,In_716);
or U1818 (N_1818,In_329,In_290);
xnor U1819 (N_1819,In_754,In_859);
xnor U1820 (N_1820,In_453,In_139);
xnor U1821 (N_1821,In_270,In_385);
or U1822 (N_1822,In_470,In_196);
xnor U1823 (N_1823,In_63,In_841);
and U1824 (N_1824,In_345,In_713);
and U1825 (N_1825,In_665,In_718);
and U1826 (N_1826,In_94,In_589);
nand U1827 (N_1827,In_673,In_469);
nor U1828 (N_1828,In_422,In_336);
nand U1829 (N_1829,In_695,In_748);
nor U1830 (N_1830,In_193,In_386);
nor U1831 (N_1831,In_656,In_808);
or U1832 (N_1832,In_836,In_387);
and U1833 (N_1833,In_546,In_749);
or U1834 (N_1834,In_648,In_828);
nand U1835 (N_1835,In_48,In_475);
or U1836 (N_1836,In_946,In_523);
nand U1837 (N_1837,In_620,In_498);
nor U1838 (N_1838,In_232,In_770);
xor U1839 (N_1839,In_29,In_669);
xnor U1840 (N_1840,In_509,In_619);
nor U1841 (N_1841,In_648,In_777);
or U1842 (N_1842,In_238,In_431);
or U1843 (N_1843,In_584,In_400);
or U1844 (N_1844,In_178,In_423);
xor U1845 (N_1845,In_815,In_830);
xnor U1846 (N_1846,In_563,In_753);
and U1847 (N_1847,In_908,In_621);
or U1848 (N_1848,In_867,In_285);
nand U1849 (N_1849,In_822,In_795);
xor U1850 (N_1850,In_875,In_561);
or U1851 (N_1851,In_229,In_583);
and U1852 (N_1852,In_732,In_329);
or U1853 (N_1853,In_617,In_642);
nor U1854 (N_1854,In_918,In_602);
xnor U1855 (N_1855,In_37,In_76);
nor U1856 (N_1856,In_239,In_271);
nand U1857 (N_1857,In_31,In_275);
xnor U1858 (N_1858,In_21,In_445);
nand U1859 (N_1859,In_804,In_983);
xnor U1860 (N_1860,In_904,In_282);
or U1861 (N_1861,In_895,In_249);
and U1862 (N_1862,In_544,In_674);
nand U1863 (N_1863,In_854,In_943);
xnor U1864 (N_1864,In_477,In_919);
or U1865 (N_1865,In_567,In_274);
nand U1866 (N_1866,In_839,In_98);
nor U1867 (N_1867,In_352,In_241);
xor U1868 (N_1868,In_946,In_867);
and U1869 (N_1869,In_237,In_59);
xnor U1870 (N_1870,In_825,In_695);
nand U1871 (N_1871,In_960,In_43);
xor U1872 (N_1872,In_303,In_82);
or U1873 (N_1873,In_305,In_831);
nand U1874 (N_1874,In_418,In_441);
or U1875 (N_1875,In_10,In_716);
xor U1876 (N_1876,In_68,In_850);
nand U1877 (N_1877,In_140,In_53);
and U1878 (N_1878,In_967,In_597);
xor U1879 (N_1879,In_645,In_823);
nor U1880 (N_1880,In_680,In_499);
and U1881 (N_1881,In_598,In_671);
or U1882 (N_1882,In_338,In_187);
nor U1883 (N_1883,In_603,In_222);
nand U1884 (N_1884,In_643,In_853);
nor U1885 (N_1885,In_251,In_771);
nand U1886 (N_1886,In_824,In_291);
or U1887 (N_1887,In_628,In_698);
nand U1888 (N_1888,In_749,In_508);
nand U1889 (N_1889,In_12,In_303);
or U1890 (N_1890,In_577,In_163);
and U1891 (N_1891,In_159,In_731);
nand U1892 (N_1892,In_154,In_660);
nor U1893 (N_1893,In_721,In_53);
nor U1894 (N_1894,In_55,In_909);
xor U1895 (N_1895,In_138,In_981);
xnor U1896 (N_1896,In_272,In_755);
xnor U1897 (N_1897,In_121,In_476);
xor U1898 (N_1898,In_839,In_768);
nor U1899 (N_1899,In_555,In_394);
nor U1900 (N_1900,In_327,In_494);
nand U1901 (N_1901,In_953,In_685);
and U1902 (N_1902,In_455,In_911);
xor U1903 (N_1903,In_867,In_550);
nor U1904 (N_1904,In_872,In_995);
nor U1905 (N_1905,In_943,In_254);
and U1906 (N_1906,In_899,In_271);
nand U1907 (N_1907,In_578,In_291);
xor U1908 (N_1908,In_398,In_320);
and U1909 (N_1909,In_176,In_670);
and U1910 (N_1910,In_193,In_529);
nor U1911 (N_1911,In_777,In_250);
nand U1912 (N_1912,In_116,In_42);
nand U1913 (N_1913,In_850,In_678);
or U1914 (N_1914,In_299,In_141);
nand U1915 (N_1915,In_280,In_73);
nand U1916 (N_1916,In_802,In_701);
and U1917 (N_1917,In_292,In_696);
or U1918 (N_1918,In_1,In_16);
nor U1919 (N_1919,In_234,In_923);
and U1920 (N_1920,In_872,In_703);
xnor U1921 (N_1921,In_997,In_334);
nor U1922 (N_1922,In_472,In_846);
nor U1923 (N_1923,In_834,In_5);
or U1924 (N_1924,In_670,In_339);
xor U1925 (N_1925,In_136,In_898);
xor U1926 (N_1926,In_811,In_141);
nand U1927 (N_1927,In_200,In_225);
nor U1928 (N_1928,In_65,In_240);
nor U1929 (N_1929,In_924,In_524);
xor U1930 (N_1930,In_631,In_328);
or U1931 (N_1931,In_831,In_42);
nand U1932 (N_1932,In_450,In_116);
nor U1933 (N_1933,In_12,In_604);
nor U1934 (N_1934,In_513,In_312);
nor U1935 (N_1935,In_294,In_236);
xnor U1936 (N_1936,In_937,In_459);
or U1937 (N_1937,In_789,In_751);
nand U1938 (N_1938,In_448,In_469);
or U1939 (N_1939,In_82,In_963);
and U1940 (N_1940,In_558,In_323);
or U1941 (N_1941,In_70,In_731);
xor U1942 (N_1942,In_66,In_543);
or U1943 (N_1943,In_258,In_369);
or U1944 (N_1944,In_683,In_73);
or U1945 (N_1945,In_906,In_138);
or U1946 (N_1946,In_498,In_321);
nand U1947 (N_1947,In_940,In_409);
and U1948 (N_1948,In_147,In_838);
xor U1949 (N_1949,In_258,In_474);
nor U1950 (N_1950,In_327,In_309);
or U1951 (N_1951,In_104,In_726);
nor U1952 (N_1952,In_574,In_860);
xnor U1953 (N_1953,In_893,In_892);
nand U1954 (N_1954,In_846,In_826);
xor U1955 (N_1955,In_383,In_535);
or U1956 (N_1956,In_7,In_371);
nor U1957 (N_1957,In_77,In_636);
or U1958 (N_1958,In_921,In_748);
or U1959 (N_1959,In_690,In_362);
or U1960 (N_1960,In_482,In_869);
nor U1961 (N_1961,In_79,In_595);
or U1962 (N_1962,In_332,In_377);
or U1963 (N_1963,In_110,In_106);
and U1964 (N_1964,In_698,In_586);
nor U1965 (N_1965,In_197,In_610);
nor U1966 (N_1966,In_605,In_722);
nor U1967 (N_1967,In_87,In_695);
and U1968 (N_1968,In_660,In_571);
nor U1969 (N_1969,In_585,In_965);
xor U1970 (N_1970,In_469,In_240);
nor U1971 (N_1971,In_490,In_301);
nand U1972 (N_1972,In_145,In_100);
xnor U1973 (N_1973,In_21,In_125);
and U1974 (N_1974,In_793,In_38);
xor U1975 (N_1975,In_981,In_431);
and U1976 (N_1976,In_243,In_979);
nor U1977 (N_1977,In_231,In_224);
and U1978 (N_1978,In_221,In_515);
nor U1979 (N_1979,In_561,In_878);
nand U1980 (N_1980,In_820,In_829);
nor U1981 (N_1981,In_496,In_279);
nor U1982 (N_1982,In_649,In_307);
nor U1983 (N_1983,In_417,In_466);
and U1984 (N_1984,In_319,In_254);
xnor U1985 (N_1985,In_879,In_45);
xor U1986 (N_1986,In_68,In_234);
and U1987 (N_1987,In_35,In_351);
nor U1988 (N_1988,In_121,In_7);
and U1989 (N_1989,In_751,In_889);
xnor U1990 (N_1990,In_738,In_59);
and U1991 (N_1991,In_572,In_978);
and U1992 (N_1992,In_572,In_348);
nor U1993 (N_1993,In_441,In_166);
nand U1994 (N_1994,In_303,In_696);
xor U1995 (N_1995,In_756,In_680);
nand U1996 (N_1996,In_643,In_871);
or U1997 (N_1997,In_577,In_514);
nor U1998 (N_1998,In_864,In_699);
or U1999 (N_1999,In_671,In_192);
xnor U2000 (N_2000,In_71,In_35);
nor U2001 (N_2001,In_226,In_252);
nor U2002 (N_2002,In_522,In_313);
nor U2003 (N_2003,In_179,In_548);
and U2004 (N_2004,In_88,In_192);
and U2005 (N_2005,In_478,In_990);
or U2006 (N_2006,In_351,In_969);
and U2007 (N_2007,In_594,In_375);
and U2008 (N_2008,In_848,In_978);
or U2009 (N_2009,In_733,In_825);
and U2010 (N_2010,In_472,In_942);
and U2011 (N_2011,In_227,In_568);
and U2012 (N_2012,In_566,In_355);
nor U2013 (N_2013,In_418,In_451);
xor U2014 (N_2014,In_835,In_319);
xor U2015 (N_2015,In_960,In_316);
xor U2016 (N_2016,In_667,In_917);
nor U2017 (N_2017,In_655,In_771);
or U2018 (N_2018,In_616,In_196);
nor U2019 (N_2019,In_346,In_703);
xnor U2020 (N_2020,In_265,In_622);
nand U2021 (N_2021,In_430,In_816);
and U2022 (N_2022,In_386,In_990);
or U2023 (N_2023,In_248,In_823);
or U2024 (N_2024,In_927,In_221);
nor U2025 (N_2025,In_905,In_261);
nor U2026 (N_2026,In_248,In_133);
nand U2027 (N_2027,In_586,In_415);
xnor U2028 (N_2028,In_38,In_157);
nand U2029 (N_2029,In_792,In_136);
nor U2030 (N_2030,In_231,In_571);
xor U2031 (N_2031,In_227,In_942);
and U2032 (N_2032,In_357,In_898);
nand U2033 (N_2033,In_576,In_204);
and U2034 (N_2034,In_362,In_317);
and U2035 (N_2035,In_698,In_311);
xor U2036 (N_2036,In_600,In_307);
nand U2037 (N_2037,In_130,In_933);
nor U2038 (N_2038,In_876,In_928);
nand U2039 (N_2039,In_903,In_729);
nor U2040 (N_2040,In_360,In_880);
nand U2041 (N_2041,In_816,In_48);
xnor U2042 (N_2042,In_29,In_258);
and U2043 (N_2043,In_487,In_371);
nand U2044 (N_2044,In_789,In_461);
xnor U2045 (N_2045,In_335,In_582);
nand U2046 (N_2046,In_619,In_418);
and U2047 (N_2047,In_760,In_693);
nor U2048 (N_2048,In_421,In_454);
or U2049 (N_2049,In_562,In_137);
nor U2050 (N_2050,In_4,In_941);
nand U2051 (N_2051,In_534,In_399);
xor U2052 (N_2052,In_120,In_325);
and U2053 (N_2053,In_797,In_613);
and U2054 (N_2054,In_270,In_796);
and U2055 (N_2055,In_967,In_453);
and U2056 (N_2056,In_236,In_881);
or U2057 (N_2057,In_101,In_129);
nand U2058 (N_2058,In_341,In_397);
xor U2059 (N_2059,In_304,In_54);
and U2060 (N_2060,In_24,In_55);
xnor U2061 (N_2061,In_161,In_622);
or U2062 (N_2062,In_431,In_292);
nand U2063 (N_2063,In_356,In_103);
or U2064 (N_2064,In_470,In_113);
or U2065 (N_2065,In_831,In_280);
xor U2066 (N_2066,In_337,In_120);
and U2067 (N_2067,In_746,In_488);
and U2068 (N_2068,In_637,In_956);
and U2069 (N_2069,In_945,In_886);
and U2070 (N_2070,In_5,In_24);
xnor U2071 (N_2071,In_376,In_327);
nor U2072 (N_2072,In_105,In_931);
nor U2073 (N_2073,In_859,In_367);
and U2074 (N_2074,In_276,In_274);
or U2075 (N_2075,In_902,In_99);
and U2076 (N_2076,In_651,In_675);
xor U2077 (N_2077,In_720,In_945);
or U2078 (N_2078,In_782,In_289);
nor U2079 (N_2079,In_552,In_716);
or U2080 (N_2080,In_479,In_425);
or U2081 (N_2081,In_298,In_415);
and U2082 (N_2082,In_381,In_203);
xnor U2083 (N_2083,In_885,In_450);
xnor U2084 (N_2084,In_965,In_985);
and U2085 (N_2085,In_280,In_872);
or U2086 (N_2086,In_800,In_100);
xor U2087 (N_2087,In_865,In_497);
nor U2088 (N_2088,In_28,In_992);
and U2089 (N_2089,In_378,In_824);
or U2090 (N_2090,In_876,In_851);
nor U2091 (N_2091,In_977,In_542);
or U2092 (N_2092,In_383,In_262);
and U2093 (N_2093,In_21,In_955);
nor U2094 (N_2094,In_390,In_342);
and U2095 (N_2095,In_558,In_5);
or U2096 (N_2096,In_212,In_275);
and U2097 (N_2097,In_521,In_115);
nand U2098 (N_2098,In_224,In_133);
xnor U2099 (N_2099,In_756,In_87);
or U2100 (N_2100,In_479,In_10);
or U2101 (N_2101,In_640,In_287);
or U2102 (N_2102,In_389,In_730);
nand U2103 (N_2103,In_428,In_542);
nand U2104 (N_2104,In_794,In_954);
nand U2105 (N_2105,In_579,In_678);
nand U2106 (N_2106,In_27,In_724);
or U2107 (N_2107,In_961,In_173);
or U2108 (N_2108,In_817,In_314);
xor U2109 (N_2109,In_22,In_778);
nand U2110 (N_2110,In_761,In_602);
or U2111 (N_2111,In_242,In_743);
xnor U2112 (N_2112,In_126,In_221);
nand U2113 (N_2113,In_53,In_421);
and U2114 (N_2114,In_16,In_919);
xnor U2115 (N_2115,In_909,In_214);
xnor U2116 (N_2116,In_732,In_979);
or U2117 (N_2117,In_726,In_647);
nand U2118 (N_2118,In_811,In_838);
nand U2119 (N_2119,In_743,In_374);
nand U2120 (N_2120,In_856,In_864);
or U2121 (N_2121,In_58,In_192);
nor U2122 (N_2122,In_938,In_715);
xor U2123 (N_2123,In_640,In_815);
xor U2124 (N_2124,In_343,In_174);
and U2125 (N_2125,In_749,In_41);
xnor U2126 (N_2126,In_461,In_878);
and U2127 (N_2127,In_897,In_733);
nor U2128 (N_2128,In_774,In_633);
nand U2129 (N_2129,In_545,In_257);
or U2130 (N_2130,In_662,In_989);
or U2131 (N_2131,In_696,In_229);
or U2132 (N_2132,In_880,In_690);
xnor U2133 (N_2133,In_47,In_147);
nor U2134 (N_2134,In_516,In_38);
nor U2135 (N_2135,In_840,In_627);
nand U2136 (N_2136,In_220,In_29);
xnor U2137 (N_2137,In_860,In_26);
nand U2138 (N_2138,In_314,In_49);
nor U2139 (N_2139,In_496,In_400);
nor U2140 (N_2140,In_811,In_106);
or U2141 (N_2141,In_602,In_361);
nor U2142 (N_2142,In_238,In_280);
and U2143 (N_2143,In_702,In_255);
or U2144 (N_2144,In_18,In_773);
xnor U2145 (N_2145,In_180,In_859);
xor U2146 (N_2146,In_335,In_507);
or U2147 (N_2147,In_99,In_613);
xnor U2148 (N_2148,In_740,In_720);
nand U2149 (N_2149,In_566,In_54);
nand U2150 (N_2150,In_379,In_819);
xor U2151 (N_2151,In_320,In_591);
nor U2152 (N_2152,In_115,In_551);
nor U2153 (N_2153,In_666,In_643);
nor U2154 (N_2154,In_433,In_89);
xor U2155 (N_2155,In_309,In_176);
or U2156 (N_2156,In_488,In_335);
or U2157 (N_2157,In_482,In_885);
or U2158 (N_2158,In_544,In_685);
nor U2159 (N_2159,In_947,In_204);
nor U2160 (N_2160,In_892,In_476);
xor U2161 (N_2161,In_924,In_201);
xnor U2162 (N_2162,In_338,In_97);
nor U2163 (N_2163,In_683,In_695);
nor U2164 (N_2164,In_30,In_700);
nand U2165 (N_2165,In_246,In_594);
and U2166 (N_2166,In_312,In_924);
or U2167 (N_2167,In_130,In_209);
xnor U2168 (N_2168,In_214,In_948);
nor U2169 (N_2169,In_71,In_904);
or U2170 (N_2170,In_572,In_964);
xor U2171 (N_2171,In_878,In_718);
xnor U2172 (N_2172,In_189,In_191);
and U2173 (N_2173,In_871,In_149);
and U2174 (N_2174,In_850,In_51);
xor U2175 (N_2175,In_897,In_953);
or U2176 (N_2176,In_844,In_411);
xnor U2177 (N_2177,In_965,In_16);
xor U2178 (N_2178,In_43,In_921);
nor U2179 (N_2179,In_217,In_815);
nand U2180 (N_2180,In_575,In_898);
nor U2181 (N_2181,In_790,In_750);
nor U2182 (N_2182,In_493,In_652);
nor U2183 (N_2183,In_602,In_907);
xnor U2184 (N_2184,In_239,In_351);
nor U2185 (N_2185,In_942,In_903);
or U2186 (N_2186,In_978,In_342);
or U2187 (N_2187,In_176,In_298);
and U2188 (N_2188,In_386,In_679);
nand U2189 (N_2189,In_528,In_274);
xor U2190 (N_2190,In_303,In_545);
nor U2191 (N_2191,In_749,In_686);
nor U2192 (N_2192,In_605,In_574);
nor U2193 (N_2193,In_115,In_168);
nor U2194 (N_2194,In_219,In_265);
nor U2195 (N_2195,In_613,In_665);
and U2196 (N_2196,In_547,In_331);
nand U2197 (N_2197,In_918,In_358);
and U2198 (N_2198,In_913,In_305);
nor U2199 (N_2199,In_542,In_9);
and U2200 (N_2200,In_28,In_264);
nor U2201 (N_2201,In_97,In_363);
nor U2202 (N_2202,In_634,In_315);
xnor U2203 (N_2203,In_856,In_549);
nand U2204 (N_2204,In_923,In_269);
nand U2205 (N_2205,In_246,In_920);
and U2206 (N_2206,In_422,In_30);
nor U2207 (N_2207,In_571,In_347);
nand U2208 (N_2208,In_774,In_378);
and U2209 (N_2209,In_872,In_682);
xor U2210 (N_2210,In_995,In_133);
nand U2211 (N_2211,In_379,In_471);
nor U2212 (N_2212,In_71,In_830);
or U2213 (N_2213,In_917,In_859);
and U2214 (N_2214,In_251,In_227);
xor U2215 (N_2215,In_804,In_682);
nor U2216 (N_2216,In_722,In_179);
and U2217 (N_2217,In_33,In_925);
or U2218 (N_2218,In_303,In_463);
nor U2219 (N_2219,In_593,In_750);
and U2220 (N_2220,In_596,In_520);
nand U2221 (N_2221,In_790,In_373);
or U2222 (N_2222,In_41,In_352);
and U2223 (N_2223,In_562,In_345);
xnor U2224 (N_2224,In_732,In_812);
and U2225 (N_2225,In_166,In_60);
xor U2226 (N_2226,In_483,In_399);
and U2227 (N_2227,In_290,In_458);
nand U2228 (N_2228,In_269,In_931);
and U2229 (N_2229,In_40,In_210);
and U2230 (N_2230,In_812,In_923);
nor U2231 (N_2231,In_975,In_676);
nand U2232 (N_2232,In_775,In_424);
nand U2233 (N_2233,In_680,In_801);
or U2234 (N_2234,In_920,In_994);
xor U2235 (N_2235,In_856,In_728);
or U2236 (N_2236,In_631,In_43);
xnor U2237 (N_2237,In_814,In_842);
nor U2238 (N_2238,In_857,In_159);
nor U2239 (N_2239,In_269,In_300);
or U2240 (N_2240,In_616,In_808);
and U2241 (N_2241,In_711,In_941);
nand U2242 (N_2242,In_240,In_212);
and U2243 (N_2243,In_954,In_554);
xor U2244 (N_2244,In_55,In_449);
nor U2245 (N_2245,In_735,In_826);
xor U2246 (N_2246,In_991,In_101);
nor U2247 (N_2247,In_846,In_578);
nor U2248 (N_2248,In_557,In_961);
and U2249 (N_2249,In_686,In_180);
xnor U2250 (N_2250,In_307,In_339);
and U2251 (N_2251,In_684,In_304);
and U2252 (N_2252,In_629,In_83);
or U2253 (N_2253,In_776,In_396);
or U2254 (N_2254,In_956,In_447);
or U2255 (N_2255,In_62,In_676);
xnor U2256 (N_2256,In_783,In_793);
and U2257 (N_2257,In_744,In_587);
or U2258 (N_2258,In_821,In_218);
nand U2259 (N_2259,In_503,In_220);
or U2260 (N_2260,In_654,In_191);
nor U2261 (N_2261,In_609,In_598);
or U2262 (N_2262,In_648,In_162);
nor U2263 (N_2263,In_634,In_377);
or U2264 (N_2264,In_214,In_282);
and U2265 (N_2265,In_238,In_306);
and U2266 (N_2266,In_885,In_136);
nor U2267 (N_2267,In_891,In_544);
or U2268 (N_2268,In_432,In_58);
or U2269 (N_2269,In_191,In_837);
or U2270 (N_2270,In_355,In_419);
or U2271 (N_2271,In_124,In_413);
or U2272 (N_2272,In_932,In_135);
xnor U2273 (N_2273,In_875,In_774);
xnor U2274 (N_2274,In_339,In_422);
nor U2275 (N_2275,In_691,In_788);
and U2276 (N_2276,In_142,In_903);
xnor U2277 (N_2277,In_764,In_803);
xor U2278 (N_2278,In_206,In_782);
nand U2279 (N_2279,In_340,In_361);
or U2280 (N_2280,In_472,In_608);
nor U2281 (N_2281,In_872,In_462);
xnor U2282 (N_2282,In_432,In_927);
xor U2283 (N_2283,In_157,In_354);
or U2284 (N_2284,In_190,In_802);
xor U2285 (N_2285,In_896,In_3);
or U2286 (N_2286,In_253,In_954);
xnor U2287 (N_2287,In_822,In_156);
xor U2288 (N_2288,In_79,In_150);
xnor U2289 (N_2289,In_417,In_976);
nor U2290 (N_2290,In_860,In_488);
nand U2291 (N_2291,In_663,In_97);
nand U2292 (N_2292,In_443,In_407);
nor U2293 (N_2293,In_887,In_964);
nor U2294 (N_2294,In_764,In_409);
or U2295 (N_2295,In_915,In_742);
xnor U2296 (N_2296,In_398,In_242);
and U2297 (N_2297,In_19,In_369);
nor U2298 (N_2298,In_885,In_98);
xnor U2299 (N_2299,In_772,In_386);
xor U2300 (N_2300,In_504,In_443);
and U2301 (N_2301,In_688,In_228);
nand U2302 (N_2302,In_903,In_275);
and U2303 (N_2303,In_573,In_961);
nand U2304 (N_2304,In_832,In_646);
nor U2305 (N_2305,In_749,In_623);
or U2306 (N_2306,In_200,In_437);
nand U2307 (N_2307,In_750,In_268);
xnor U2308 (N_2308,In_428,In_806);
nor U2309 (N_2309,In_365,In_991);
or U2310 (N_2310,In_979,In_928);
or U2311 (N_2311,In_138,In_632);
xor U2312 (N_2312,In_927,In_441);
xnor U2313 (N_2313,In_240,In_314);
nor U2314 (N_2314,In_537,In_218);
xor U2315 (N_2315,In_711,In_16);
or U2316 (N_2316,In_61,In_393);
nor U2317 (N_2317,In_898,In_757);
xnor U2318 (N_2318,In_764,In_788);
nor U2319 (N_2319,In_316,In_793);
or U2320 (N_2320,In_81,In_356);
nand U2321 (N_2321,In_681,In_493);
nor U2322 (N_2322,In_644,In_500);
nand U2323 (N_2323,In_941,In_787);
nor U2324 (N_2324,In_877,In_763);
nand U2325 (N_2325,In_622,In_891);
and U2326 (N_2326,In_585,In_429);
xnor U2327 (N_2327,In_220,In_635);
and U2328 (N_2328,In_735,In_271);
or U2329 (N_2329,In_593,In_192);
or U2330 (N_2330,In_585,In_979);
nor U2331 (N_2331,In_744,In_407);
nor U2332 (N_2332,In_790,In_99);
nand U2333 (N_2333,In_597,In_522);
nand U2334 (N_2334,In_743,In_827);
or U2335 (N_2335,In_462,In_85);
or U2336 (N_2336,In_457,In_6);
nor U2337 (N_2337,In_67,In_354);
and U2338 (N_2338,In_954,In_285);
and U2339 (N_2339,In_780,In_472);
and U2340 (N_2340,In_534,In_731);
nor U2341 (N_2341,In_627,In_550);
xor U2342 (N_2342,In_59,In_176);
nor U2343 (N_2343,In_484,In_189);
xnor U2344 (N_2344,In_121,In_996);
nor U2345 (N_2345,In_730,In_161);
nor U2346 (N_2346,In_615,In_57);
and U2347 (N_2347,In_307,In_48);
and U2348 (N_2348,In_825,In_339);
and U2349 (N_2349,In_806,In_897);
or U2350 (N_2350,In_693,In_702);
nand U2351 (N_2351,In_103,In_184);
nor U2352 (N_2352,In_60,In_119);
nand U2353 (N_2353,In_865,In_404);
nor U2354 (N_2354,In_738,In_231);
and U2355 (N_2355,In_94,In_647);
or U2356 (N_2356,In_704,In_797);
xnor U2357 (N_2357,In_343,In_191);
nor U2358 (N_2358,In_991,In_418);
and U2359 (N_2359,In_597,In_592);
or U2360 (N_2360,In_334,In_847);
or U2361 (N_2361,In_174,In_134);
or U2362 (N_2362,In_450,In_12);
and U2363 (N_2363,In_86,In_479);
and U2364 (N_2364,In_248,In_884);
nand U2365 (N_2365,In_590,In_689);
xor U2366 (N_2366,In_254,In_180);
nor U2367 (N_2367,In_486,In_303);
nor U2368 (N_2368,In_201,In_464);
xnor U2369 (N_2369,In_319,In_439);
and U2370 (N_2370,In_33,In_244);
nor U2371 (N_2371,In_710,In_714);
nor U2372 (N_2372,In_778,In_415);
nand U2373 (N_2373,In_708,In_812);
nand U2374 (N_2374,In_318,In_422);
and U2375 (N_2375,In_947,In_671);
or U2376 (N_2376,In_572,In_794);
xnor U2377 (N_2377,In_676,In_55);
nand U2378 (N_2378,In_794,In_770);
and U2379 (N_2379,In_355,In_310);
or U2380 (N_2380,In_152,In_227);
nor U2381 (N_2381,In_905,In_933);
and U2382 (N_2382,In_270,In_114);
nor U2383 (N_2383,In_854,In_699);
and U2384 (N_2384,In_486,In_555);
or U2385 (N_2385,In_757,In_377);
and U2386 (N_2386,In_718,In_899);
xnor U2387 (N_2387,In_710,In_12);
or U2388 (N_2388,In_681,In_144);
nand U2389 (N_2389,In_644,In_641);
xnor U2390 (N_2390,In_192,In_755);
nor U2391 (N_2391,In_350,In_488);
nand U2392 (N_2392,In_196,In_615);
and U2393 (N_2393,In_119,In_211);
and U2394 (N_2394,In_322,In_906);
nor U2395 (N_2395,In_102,In_599);
nand U2396 (N_2396,In_494,In_987);
nand U2397 (N_2397,In_492,In_501);
xnor U2398 (N_2398,In_221,In_831);
nor U2399 (N_2399,In_101,In_764);
or U2400 (N_2400,In_148,In_624);
nand U2401 (N_2401,In_70,In_330);
nor U2402 (N_2402,In_677,In_233);
and U2403 (N_2403,In_913,In_536);
xnor U2404 (N_2404,In_310,In_443);
xor U2405 (N_2405,In_90,In_24);
or U2406 (N_2406,In_345,In_193);
or U2407 (N_2407,In_823,In_120);
or U2408 (N_2408,In_67,In_736);
nand U2409 (N_2409,In_799,In_446);
xor U2410 (N_2410,In_878,In_96);
or U2411 (N_2411,In_149,In_457);
nand U2412 (N_2412,In_7,In_129);
nand U2413 (N_2413,In_564,In_525);
or U2414 (N_2414,In_716,In_679);
and U2415 (N_2415,In_692,In_238);
or U2416 (N_2416,In_384,In_973);
nand U2417 (N_2417,In_331,In_115);
nor U2418 (N_2418,In_53,In_990);
xnor U2419 (N_2419,In_347,In_379);
or U2420 (N_2420,In_495,In_537);
and U2421 (N_2421,In_921,In_370);
xnor U2422 (N_2422,In_633,In_839);
or U2423 (N_2423,In_436,In_87);
xor U2424 (N_2424,In_999,In_637);
or U2425 (N_2425,In_945,In_101);
nand U2426 (N_2426,In_234,In_131);
nand U2427 (N_2427,In_30,In_949);
or U2428 (N_2428,In_210,In_281);
nor U2429 (N_2429,In_145,In_541);
nor U2430 (N_2430,In_561,In_126);
and U2431 (N_2431,In_852,In_278);
nor U2432 (N_2432,In_255,In_182);
xnor U2433 (N_2433,In_825,In_93);
nand U2434 (N_2434,In_632,In_912);
or U2435 (N_2435,In_818,In_1);
nor U2436 (N_2436,In_502,In_445);
or U2437 (N_2437,In_929,In_31);
xnor U2438 (N_2438,In_400,In_224);
and U2439 (N_2439,In_351,In_929);
or U2440 (N_2440,In_875,In_833);
or U2441 (N_2441,In_35,In_953);
nor U2442 (N_2442,In_832,In_45);
or U2443 (N_2443,In_78,In_105);
nor U2444 (N_2444,In_635,In_64);
xnor U2445 (N_2445,In_581,In_265);
nor U2446 (N_2446,In_396,In_823);
xor U2447 (N_2447,In_216,In_846);
xor U2448 (N_2448,In_888,In_116);
xnor U2449 (N_2449,In_462,In_26);
nor U2450 (N_2450,In_479,In_881);
xor U2451 (N_2451,In_929,In_654);
xnor U2452 (N_2452,In_874,In_229);
and U2453 (N_2453,In_948,In_468);
nand U2454 (N_2454,In_532,In_719);
nor U2455 (N_2455,In_550,In_631);
xor U2456 (N_2456,In_633,In_883);
nor U2457 (N_2457,In_995,In_717);
and U2458 (N_2458,In_798,In_838);
or U2459 (N_2459,In_727,In_679);
nor U2460 (N_2460,In_894,In_405);
nand U2461 (N_2461,In_326,In_695);
xor U2462 (N_2462,In_557,In_746);
and U2463 (N_2463,In_870,In_552);
or U2464 (N_2464,In_514,In_991);
and U2465 (N_2465,In_232,In_903);
xnor U2466 (N_2466,In_928,In_833);
nor U2467 (N_2467,In_198,In_540);
and U2468 (N_2468,In_165,In_742);
xor U2469 (N_2469,In_521,In_7);
nor U2470 (N_2470,In_745,In_334);
or U2471 (N_2471,In_537,In_33);
xor U2472 (N_2472,In_406,In_451);
or U2473 (N_2473,In_25,In_791);
and U2474 (N_2474,In_313,In_493);
nor U2475 (N_2475,In_400,In_276);
xnor U2476 (N_2476,In_159,In_227);
or U2477 (N_2477,In_905,In_325);
xnor U2478 (N_2478,In_380,In_560);
and U2479 (N_2479,In_981,In_465);
or U2480 (N_2480,In_558,In_561);
nor U2481 (N_2481,In_991,In_496);
nand U2482 (N_2482,In_60,In_16);
nand U2483 (N_2483,In_98,In_933);
and U2484 (N_2484,In_193,In_977);
xnor U2485 (N_2485,In_78,In_740);
xor U2486 (N_2486,In_194,In_375);
or U2487 (N_2487,In_428,In_102);
nand U2488 (N_2488,In_97,In_820);
nor U2489 (N_2489,In_473,In_949);
nand U2490 (N_2490,In_847,In_29);
nand U2491 (N_2491,In_835,In_263);
nor U2492 (N_2492,In_223,In_580);
and U2493 (N_2493,In_112,In_687);
nand U2494 (N_2494,In_71,In_289);
or U2495 (N_2495,In_154,In_897);
xor U2496 (N_2496,In_153,In_48);
xor U2497 (N_2497,In_895,In_751);
nand U2498 (N_2498,In_398,In_288);
or U2499 (N_2499,In_258,In_701);
xnor U2500 (N_2500,N_991,N_366);
and U2501 (N_2501,N_279,N_126);
or U2502 (N_2502,N_1443,N_1897);
or U2503 (N_2503,N_2399,N_904);
or U2504 (N_2504,N_1522,N_2008);
and U2505 (N_2505,N_200,N_321);
and U2506 (N_2506,N_8,N_1416);
nor U2507 (N_2507,N_2291,N_1590);
nand U2508 (N_2508,N_125,N_620);
xnor U2509 (N_2509,N_2035,N_331);
nor U2510 (N_2510,N_1637,N_1566);
and U2511 (N_2511,N_1963,N_1164);
nand U2512 (N_2512,N_1193,N_1041);
nor U2513 (N_2513,N_1926,N_654);
xor U2514 (N_2514,N_116,N_1050);
and U2515 (N_2515,N_839,N_2211);
xor U2516 (N_2516,N_1757,N_712);
or U2517 (N_2517,N_2121,N_1170);
nor U2518 (N_2518,N_2122,N_6);
nand U2519 (N_2519,N_2204,N_906);
nor U2520 (N_2520,N_2178,N_1955);
nor U2521 (N_2521,N_1207,N_2208);
and U2522 (N_2522,N_1005,N_2369);
xnor U2523 (N_2523,N_1221,N_1343);
nand U2524 (N_2524,N_2056,N_2415);
or U2525 (N_2525,N_1849,N_1957);
nor U2526 (N_2526,N_2433,N_1237);
nor U2527 (N_2527,N_575,N_1327);
and U2528 (N_2528,N_1846,N_1727);
or U2529 (N_2529,N_2314,N_296);
nor U2530 (N_2530,N_1117,N_2240);
or U2531 (N_2531,N_510,N_1304);
nand U2532 (N_2532,N_104,N_840);
nand U2533 (N_2533,N_1949,N_2315);
and U2534 (N_2534,N_710,N_1806);
nand U2535 (N_2535,N_878,N_1791);
and U2536 (N_2536,N_2265,N_693);
nor U2537 (N_2537,N_1652,N_1712);
xnor U2538 (N_2538,N_2063,N_2264);
and U2539 (N_2539,N_1553,N_2141);
or U2540 (N_2540,N_1022,N_2320);
and U2541 (N_2541,N_1625,N_1179);
or U2542 (N_2542,N_1009,N_618);
xnor U2543 (N_2543,N_1430,N_72);
nand U2544 (N_2544,N_1558,N_178);
nand U2545 (N_2545,N_64,N_1576);
nand U2546 (N_2546,N_1456,N_272);
nor U2547 (N_2547,N_1749,N_302);
nor U2548 (N_2548,N_2263,N_56);
or U2549 (N_2549,N_1115,N_534);
xnor U2550 (N_2550,N_1363,N_2042);
xnor U2551 (N_2551,N_1153,N_648);
nor U2552 (N_2552,N_1671,N_2000);
nand U2553 (N_2553,N_2431,N_1200);
and U2554 (N_2554,N_1542,N_2031);
or U2555 (N_2555,N_1580,N_1105);
nand U2556 (N_2556,N_294,N_1503);
nor U2557 (N_2557,N_2229,N_2447);
or U2558 (N_2558,N_303,N_2199);
xnor U2559 (N_2559,N_512,N_60);
and U2560 (N_2560,N_1433,N_1912);
xnor U2561 (N_2561,N_633,N_1687);
or U2562 (N_2562,N_305,N_2302);
nand U2563 (N_2563,N_1025,N_684);
xor U2564 (N_2564,N_2391,N_1265);
or U2565 (N_2565,N_925,N_1701);
nor U2566 (N_2566,N_516,N_386);
nor U2567 (N_2567,N_1906,N_795);
nand U2568 (N_2568,N_7,N_1403);
and U2569 (N_2569,N_66,N_809);
or U2570 (N_2570,N_554,N_1006);
nor U2571 (N_2571,N_424,N_2059);
nand U2572 (N_2572,N_1861,N_664);
or U2573 (N_2573,N_1458,N_727);
xnor U2574 (N_2574,N_1719,N_1695);
xnor U2575 (N_2575,N_1877,N_429);
or U2576 (N_2576,N_781,N_341);
nand U2577 (N_2577,N_49,N_770);
nor U2578 (N_2578,N_2450,N_1215);
and U2579 (N_2579,N_1271,N_262);
nand U2580 (N_2580,N_645,N_1648);
xnor U2581 (N_2581,N_2167,N_1726);
nor U2582 (N_2582,N_1822,N_1888);
and U2583 (N_2583,N_1072,N_2286);
xor U2584 (N_2584,N_478,N_699);
or U2585 (N_2585,N_1277,N_1928);
or U2586 (N_2586,N_2442,N_2438);
nor U2587 (N_2587,N_2444,N_1347);
xor U2588 (N_2588,N_1755,N_637);
xor U2589 (N_2589,N_69,N_1122);
nor U2590 (N_2590,N_1832,N_1395);
xor U2591 (N_2591,N_2272,N_2488);
xor U2592 (N_2592,N_1568,N_779);
nand U2593 (N_2593,N_525,N_1467);
and U2594 (N_2594,N_350,N_469);
xor U2595 (N_2595,N_2218,N_1428);
nand U2596 (N_2596,N_2099,N_31);
or U2597 (N_2597,N_1657,N_2184);
nand U2598 (N_2598,N_1176,N_772);
xnor U2599 (N_2599,N_596,N_1642);
nand U2600 (N_2600,N_2492,N_1911);
and U2601 (N_2601,N_1152,N_2343);
xnor U2602 (N_2602,N_1967,N_1059);
xor U2603 (N_2603,N_1939,N_1011);
or U2604 (N_2604,N_210,N_448);
or U2605 (N_2605,N_1269,N_441);
nor U2606 (N_2606,N_546,N_2085);
nor U2607 (N_2607,N_1212,N_1975);
and U2608 (N_2608,N_1008,N_1044);
and U2609 (N_2609,N_1811,N_1706);
nand U2610 (N_2610,N_533,N_1079);
nor U2611 (N_2611,N_347,N_1032);
nand U2612 (N_2612,N_1944,N_2055);
xor U2613 (N_2613,N_1851,N_228);
nor U2614 (N_2614,N_1898,N_2303);
nor U2615 (N_2615,N_947,N_2297);
or U2616 (N_2616,N_1740,N_308);
and U2617 (N_2617,N_509,N_544);
nor U2618 (N_2618,N_2202,N_1159);
nor U2619 (N_2619,N_549,N_765);
and U2620 (N_2620,N_1914,N_960);
nor U2621 (N_2621,N_2191,N_1979);
nand U2622 (N_2622,N_337,N_943);
and U2623 (N_2623,N_1653,N_1093);
and U2624 (N_2624,N_1233,N_1424);
and U2625 (N_2625,N_2398,N_2389);
and U2626 (N_2626,N_975,N_2361);
nand U2627 (N_2627,N_403,N_1097);
xor U2628 (N_2628,N_1400,N_744);
and U2629 (N_2629,N_382,N_1818);
and U2630 (N_2630,N_1464,N_564);
nor U2631 (N_2631,N_2223,N_1000);
and U2632 (N_2632,N_1407,N_342);
nor U2633 (N_2633,N_298,N_1320);
nand U2634 (N_2634,N_1858,N_2125);
or U2635 (N_2635,N_2247,N_158);
xor U2636 (N_2636,N_233,N_784);
xnor U2637 (N_2637,N_1581,N_1524);
xor U2638 (N_2638,N_1106,N_2325);
or U2639 (N_2639,N_754,N_1092);
nand U2640 (N_2640,N_1804,N_1619);
or U2641 (N_2641,N_1254,N_466);
xnor U2642 (N_2642,N_1085,N_1197);
nand U2643 (N_2643,N_1909,N_1547);
and U2644 (N_2644,N_1545,N_562);
xnor U2645 (N_2645,N_2321,N_2341);
or U2646 (N_2646,N_974,N_1294);
nor U2647 (N_2647,N_603,N_419);
and U2648 (N_2648,N_1284,N_2253);
nor U2649 (N_2649,N_822,N_1463);
nand U2650 (N_2650,N_1286,N_410);
nor U2651 (N_2651,N_1190,N_20);
nand U2652 (N_2652,N_928,N_1082);
xnor U2653 (N_2653,N_1487,N_786);
or U2654 (N_2654,N_1669,N_2201);
or U2655 (N_2655,N_41,N_643);
nand U2656 (N_2656,N_36,N_748);
and U2657 (N_2657,N_207,N_1996);
nand U2658 (N_2658,N_1029,N_1980);
xnor U2659 (N_2659,N_909,N_1219);
and U2660 (N_2660,N_1250,N_163);
and U2661 (N_2661,N_2082,N_1525);
nand U2662 (N_2662,N_1054,N_250);
nand U2663 (N_2663,N_1993,N_1439);
nand U2664 (N_2664,N_2044,N_1402);
xor U2665 (N_2665,N_2344,N_833);
and U2666 (N_2666,N_1845,N_834);
nand U2667 (N_2667,N_857,N_1563);
or U2668 (N_2668,N_460,N_24);
xnor U2669 (N_2669,N_1028,N_1332);
nand U2670 (N_2670,N_502,N_2053);
xnor U2671 (N_2671,N_495,N_2470);
or U2672 (N_2672,N_984,N_204);
nor U2673 (N_2673,N_854,N_2289);
or U2674 (N_2674,N_221,N_919);
nand U2675 (N_2675,N_738,N_1815);
nand U2676 (N_2676,N_2239,N_2227);
nand U2677 (N_2677,N_97,N_622);
and U2678 (N_2678,N_1516,N_1895);
and U2679 (N_2679,N_1910,N_174);
nand U2680 (N_2680,N_176,N_1102);
and U2681 (N_2681,N_918,N_616);
or U2682 (N_2682,N_83,N_2045);
nor U2683 (N_2683,N_623,N_2021);
nor U2684 (N_2684,N_1627,N_1481);
and U2685 (N_2685,N_1352,N_1497);
and U2686 (N_2686,N_1013,N_470);
nand U2687 (N_2687,N_1398,N_240);
nand U2688 (N_2688,N_388,N_1049);
xor U2689 (N_2689,N_490,N_1929);
and U2690 (N_2690,N_1418,N_373);
and U2691 (N_2691,N_810,N_764);
nor U2692 (N_2692,N_284,N_2324);
nor U2693 (N_2693,N_1730,N_1279);
nor U2694 (N_2694,N_2187,N_1229);
xnor U2695 (N_2695,N_987,N_1668);
xor U2696 (N_2696,N_923,N_474);
xnor U2697 (N_2697,N_1884,N_387);
xor U2698 (N_2698,N_1003,N_1081);
or U2699 (N_2699,N_2296,N_1891);
xor U2700 (N_2700,N_2299,N_1399);
nor U2701 (N_2701,N_107,N_1856);
and U2702 (N_2702,N_2119,N_95);
xor U2703 (N_2703,N_1792,N_1391);
or U2704 (N_2704,N_1715,N_628);
xnor U2705 (N_2705,N_218,N_306);
and U2706 (N_2706,N_553,N_288);
or U2707 (N_2707,N_1445,N_181);
nand U2708 (N_2708,N_2261,N_885);
xor U2709 (N_2709,N_108,N_2081);
xnor U2710 (N_2710,N_1252,N_498);
nand U2711 (N_2711,N_1125,N_1088);
xor U2712 (N_2712,N_1831,N_473);
or U2713 (N_2713,N_2270,N_248);
xor U2714 (N_2714,N_2334,N_1199);
nand U2715 (N_2715,N_1060,N_2032);
or U2716 (N_2716,N_1109,N_2371);
nor U2717 (N_2717,N_1878,N_571);
nor U2718 (N_2718,N_594,N_2025);
and U2719 (N_2719,N_268,N_1577);
nor U2720 (N_2720,N_1599,N_1684);
and U2721 (N_2721,N_239,N_499);
xnor U2722 (N_2722,N_300,N_1903);
or U2723 (N_2723,N_171,N_905);
or U2724 (N_2724,N_214,N_1754);
nor U2725 (N_2725,N_2379,N_1703);
and U2726 (N_2726,N_481,N_1314);
and U2727 (N_2727,N_1103,N_1189);
xor U2728 (N_2728,N_2198,N_540);
xor U2729 (N_2729,N_1673,N_890);
nand U2730 (N_2730,N_164,N_1469);
nand U2731 (N_2731,N_2098,N_850);
or U2732 (N_2732,N_90,N_2496);
xnor U2733 (N_2733,N_914,N_156);
or U2734 (N_2734,N_820,N_2233);
and U2735 (N_2735,N_472,N_825);
nand U2736 (N_2736,N_978,N_1932);
nand U2737 (N_2737,N_1457,N_101);
nor U2738 (N_2738,N_715,N_814);
xor U2739 (N_2739,N_2476,N_231);
and U2740 (N_2740,N_582,N_1107);
nor U2741 (N_2741,N_2421,N_1223);
and U2742 (N_2742,N_677,N_88);
xor U2743 (N_2743,N_2490,N_1268);
nand U2744 (N_2744,N_949,N_657);
nor U2745 (N_2745,N_216,N_2228);
or U2746 (N_2746,N_465,N_934);
nand U2747 (N_2747,N_447,N_1786);
or U2748 (N_2748,N_1483,N_802);
or U2749 (N_2749,N_1883,N_500);
nor U2750 (N_2750,N_2388,N_2093);
and U2751 (N_2751,N_505,N_996);
nor U2752 (N_2752,N_636,N_2103);
or U2753 (N_2753,N_1071,N_1242);
nand U2754 (N_2754,N_1385,N_147);
and U2755 (N_2755,N_1685,N_567);
nand U2756 (N_2756,N_894,N_1489);
and U2757 (N_2757,N_141,N_2043);
nor U2758 (N_2758,N_1732,N_80);
nand U2759 (N_2759,N_458,N_937);
or U2760 (N_2760,N_2200,N_804);
nand U2761 (N_2761,N_613,N_2084);
nand U2762 (N_2762,N_2480,N_532);
nand U2763 (N_2763,N_1045,N_1459);
nand U2764 (N_2764,N_932,N_332);
nand U2765 (N_2765,N_1194,N_1230);
nand U2766 (N_2766,N_844,N_1037);
or U2767 (N_2767,N_1287,N_1842);
or U2768 (N_2768,N_1724,N_793);
nor U2769 (N_2769,N_2460,N_901);
nand U2770 (N_2770,N_1278,N_2205);
nand U2771 (N_2771,N_1420,N_425);
nor U2772 (N_2772,N_2306,N_476);
nand U2773 (N_2773,N_1952,N_676);
or U2774 (N_2774,N_1646,N_2072);
nor U2775 (N_2775,N_2353,N_912);
xor U2776 (N_2776,N_1589,N_2231);
and U2777 (N_2777,N_243,N_940);
or U2778 (N_2778,N_1234,N_517);
xnor U2779 (N_2779,N_698,N_1244);
nor U2780 (N_2780,N_626,N_1454);
xnor U2781 (N_2781,N_264,N_59);
nor U2782 (N_2782,N_2257,N_1628);
xnor U2783 (N_2783,N_2340,N_1440);
xnor U2784 (N_2784,N_192,N_333);
or U2785 (N_2785,N_1388,N_1203);
or U2786 (N_2786,N_1206,N_1019);
nand U2787 (N_2787,N_1473,N_2238);
nand U2788 (N_2788,N_1536,N_573);
or U2789 (N_2789,N_1246,N_1656);
xor U2790 (N_2790,N_607,N_2235);
nor U2791 (N_2791,N_2013,N_364);
or U2792 (N_2792,N_756,N_589);
nor U2793 (N_2793,N_2499,N_102);
and U2794 (N_2794,N_432,N_1309);
nand U2795 (N_2795,N_1655,N_1211);
nand U2796 (N_2796,N_187,N_873);
xor U2797 (N_2797,N_871,N_504);
nand U2798 (N_2798,N_426,N_84);
and U2799 (N_2799,N_1056,N_2335);
or U2800 (N_2800,N_2294,N_494);
nand U2801 (N_2801,N_1172,N_994);
nor U2802 (N_2802,N_1354,N_690);
nand U2803 (N_2803,N_2277,N_1185);
xnor U2804 (N_2804,N_2271,N_1120);
or U2805 (N_2805,N_979,N_1165);
and U2806 (N_2806,N_2175,N_2118);
nand U2807 (N_2807,N_1787,N_1406);
nor U2808 (N_2808,N_1774,N_1587);
nand U2809 (N_2809,N_1782,N_902);
xor U2810 (N_2810,N_1797,N_2163);
nand U2811 (N_2811,N_758,N_1617);
nor U2812 (N_2812,N_1667,N_1514);
xor U2813 (N_2813,N_1511,N_444);
xor U2814 (N_2814,N_1591,N_471);
xnor U2815 (N_2815,N_1578,N_777);
or U2816 (N_2816,N_1890,N_431);
xnor U2817 (N_2817,N_1471,N_735);
and U2818 (N_2818,N_1700,N_824);
and U2819 (N_2819,N_1258,N_1348);
or U2820 (N_2820,N_2160,N_428);
and U2821 (N_2821,N_397,N_1770);
and U2822 (N_2822,N_1969,N_184);
xnor U2823 (N_2823,N_113,N_1208);
nand U2824 (N_2824,N_1881,N_1351);
nor U2825 (N_2825,N_1790,N_801);
nand U2826 (N_2826,N_2484,N_1065);
nor U2827 (N_2827,N_980,N_212);
xor U2828 (N_2828,N_1549,N_1075);
nor U2829 (N_2829,N_278,N_19);
xnor U2830 (N_2830,N_2129,N_1339);
and U2831 (N_2831,N_1736,N_2134);
nand U2832 (N_2832,N_1341,N_1981);
or U2833 (N_2833,N_1699,N_415);
nand U2834 (N_2834,N_903,N_1350);
or U2835 (N_2835,N_719,N_746);
or U2836 (N_2836,N_989,N_487);
and U2837 (N_2837,N_531,N_1731);
xnor U2838 (N_2838,N_1989,N_370);
and U2839 (N_2839,N_1303,N_1994);
and U2840 (N_2840,N_1276,N_503);
and U2841 (N_2841,N_2087,N_860);
nand U2842 (N_2842,N_1520,N_1261);
xor U2843 (N_2843,N_1896,N_723);
or U2844 (N_2844,N_2094,N_806);
nor U2845 (N_2845,N_2383,N_1679);
xor U2846 (N_2846,N_2097,N_2137);
or U2847 (N_2847,N_2077,N_150);
nand U2848 (N_2848,N_2308,N_274);
nor U2849 (N_2849,N_2176,N_707);
nand U2850 (N_2850,N_583,N_1893);
and U2851 (N_2851,N_2188,N_1370);
xor U2852 (N_2852,N_800,N_2130);
or U2853 (N_2853,N_70,N_351);
nand U2854 (N_2854,N_2076,N_1753);
nand U2855 (N_2855,N_1630,N_841);
or U2856 (N_2856,N_2100,N_1959);
and U2857 (N_2857,N_1964,N_2375);
and U2858 (N_2858,N_1329,N_1780);
and U2859 (N_2859,N_557,N_1697);
nor U2860 (N_2860,N_577,N_1758);
or U2861 (N_2861,N_1010,N_2242);
and U2862 (N_2862,N_961,N_2126);
nor U2863 (N_2863,N_2086,N_1427);
and U2864 (N_2864,N_1323,N_2236);
nand U2865 (N_2865,N_1681,N_335);
and U2866 (N_2866,N_442,N_614);
nand U2867 (N_2867,N_111,N_1848);
nor U2868 (N_2868,N_1559,N_2158);
nor U2869 (N_2869,N_1337,N_1099);
xor U2870 (N_2870,N_563,N_796);
nand U2871 (N_2871,N_823,N_1675);
xnor U2872 (N_2872,N_1512,N_2120);
and U2873 (N_2873,N_2112,N_1048);
nand U2874 (N_2874,N_2215,N_2057);
and U2875 (N_2875,N_1196,N_1415);
nand U2876 (N_2876,N_445,N_2424);
or U2877 (N_2877,N_2357,N_2052);
or U2878 (N_2878,N_385,N_1530);
xnor U2879 (N_2879,N_1708,N_635);
and U2880 (N_2880,N_260,N_1425);
and U2881 (N_2881,N_853,N_1145);
nand U2882 (N_2882,N_1725,N_1356);
xor U2883 (N_2883,N_2454,N_2010);
and U2884 (N_2884,N_1633,N_457);
and U2885 (N_2885,N_604,N_202);
or U2886 (N_2886,N_1518,N_550);
or U2887 (N_2887,N_2473,N_2329);
or U2888 (N_2888,N_2323,N_2350);
or U2889 (N_2889,N_1158,N_87);
xnor U2890 (N_2890,N_407,N_1431);
nand U2891 (N_2891,N_527,N_1186);
nor U2892 (N_2892,N_52,N_2001);
nand U2893 (N_2893,N_2016,N_2019);
or U2894 (N_2894,N_1761,N_1776);
nand U2895 (N_2895,N_1763,N_365);
xor U2896 (N_2896,N_168,N_1950);
xnor U2897 (N_2897,N_1224,N_1873);
or U2898 (N_2898,N_2007,N_1535);
or U2899 (N_2899,N_2073,N_55);
xnor U2900 (N_2900,N_1616,N_486);
nor U2901 (N_2901,N_2387,N_1340);
nor U2902 (N_2902,N_1023,N_287);
or U2903 (N_2903,N_2177,N_1750);
xnor U2904 (N_2904,N_1519,N_390);
or U2905 (N_2905,N_2083,N_1643);
nand U2906 (N_2906,N_1868,N_378);
xnor U2907 (N_2907,N_523,N_874);
and U2908 (N_2908,N_1833,N_1798);
nor U2909 (N_2909,N_2095,N_1042);
nor U2910 (N_2910,N_2402,N_652);
nand U2911 (N_2911,N_995,N_1863);
xnor U2912 (N_2912,N_861,N_1070);
and U2913 (N_2913,N_952,N_1647);
xor U2914 (N_2914,N_526,N_552);
nand U2915 (N_2915,N_1598,N_423);
xnor U2916 (N_2916,N_1216,N_286);
xor U2917 (N_2917,N_511,N_30);
xor U2918 (N_2918,N_408,N_1249);
xor U2919 (N_2919,N_1331,N_2498);
or U2920 (N_2920,N_2209,N_2394);
nand U2921 (N_2921,N_1016,N_1275);
xnor U2922 (N_2922,N_488,N_599);
nor U2923 (N_2923,N_354,N_91);
nand U2924 (N_2924,N_2292,N_866);
and U2925 (N_2925,N_1710,N_2089);
nand U2926 (N_2926,N_1645,N_1887);
nand U2927 (N_2927,N_454,N_398);
xnor U2928 (N_2928,N_1722,N_461);
and U2929 (N_2929,N_688,N_1299);
nor U2930 (N_2930,N_658,N_631);
nand U2931 (N_2931,N_1245,N_543);
nor U2932 (N_2932,N_2135,N_965);
or U2933 (N_2933,N_931,N_1654);
nand U2934 (N_2934,N_237,N_106);
or U2935 (N_2935,N_485,N_411);
nor U2936 (N_2936,N_2298,N_1479);
nand U2937 (N_2937,N_468,N_1499);
nand U2938 (N_2938,N_1389,N_2406);
nand U2939 (N_2939,N_893,N_2070);
or U2940 (N_2940,N_1381,N_1735);
nor U2941 (N_2941,N_2168,N_681);
or U2942 (N_2942,N_740,N_1317);
and U2943 (N_2943,N_1132,N_506);
and U2944 (N_2944,N_2061,N_1584);
and U2945 (N_2945,N_334,N_1650);
or U2946 (N_2946,N_2461,N_175);
nand U2947 (N_2947,N_145,N_2312);
nand U2948 (N_2948,N_2301,N_799);
xnor U2949 (N_2949,N_1593,N_182);
nor U2950 (N_2950,N_724,N_555);
or U2951 (N_2951,N_1956,N_640);
and U2952 (N_2952,N_160,N_2342);
and U2953 (N_2953,N_2405,N_1134);
or U2954 (N_2954,N_316,N_1838);
xnor U2955 (N_2955,N_944,N_281);
nor U2956 (N_2956,N_2050,N_1235);
nor U2957 (N_2957,N_1098,N_229);
nor U2958 (N_2958,N_2445,N_1614);
and U2959 (N_2959,N_2017,N_217);
and U2960 (N_2960,N_93,N_392);
xnor U2961 (N_2961,N_1690,N_817);
nor U2962 (N_2962,N_612,N_1604);
nand U2963 (N_2963,N_2434,N_692);
and U2964 (N_2964,N_930,N_1879);
nor U2965 (N_2965,N_1948,N_263);
and U2966 (N_2966,N_2276,N_406);
and U2967 (N_2967,N_2092,N_219);
xnor U2968 (N_2968,N_1670,N_701);
xnor U2969 (N_2969,N_2469,N_1823);
nor U2970 (N_2970,N_958,N_1847);
and U2971 (N_2971,N_2249,N_665);
or U2972 (N_2972,N_1131,N_2411);
nor U2973 (N_2973,N_339,N_267);
nor U2974 (N_2974,N_1639,N_1191);
and U2975 (N_2975,N_1857,N_1934);
and U2976 (N_2976,N_1401,N_2436);
nand U2977 (N_2977,N_2128,N_2290);
nand U2978 (N_2978,N_1156,N_1442);
or U2979 (N_2979,N_1205,N_371);
xnor U2980 (N_2980,N_556,N_674);
nor U2981 (N_2981,N_811,N_2385);
or U2982 (N_2982,N_946,N_1765);
nand U2983 (N_2983,N_330,N_492);
nor U2984 (N_2984,N_282,N_1169);
or U2985 (N_2985,N_805,N_2071);
xor U2986 (N_2986,N_1579,N_170);
or U2987 (N_2987,N_2475,N_558);
xnor U2988 (N_2988,N_2154,N_16);
and U2989 (N_2989,N_1181,N_1978);
nand U2990 (N_2990,N_1917,N_166);
xor U2991 (N_2991,N_2040,N_694);
xor U2992 (N_2992,N_702,N_1241);
nor U2993 (N_2993,N_1586,N_2221);
and U2994 (N_2994,N_1933,N_2192);
and U2995 (N_2995,N_1455,N_265);
xor U2996 (N_2996,N_1338,N_1918);
and U2997 (N_2997,N_2190,N_545);
nor U2998 (N_2998,N_258,N_1262);
or U2999 (N_2999,N_2495,N_57);
nand U3000 (N_3000,N_1394,N_1253);
nand U3001 (N_3001,N_1359,N_430);
xnor U3002 (N_3002,N_1527,N_2058);
nand U3003 (N_3003,N_852,N_2074);
and U3004 (N_3004,N_1069,N_1691);
nand U3005 (N_3005,N_2448,N_1876);
or U3006 (N_3006,N_667,N_1539);
or U3007 (N_3007,N_2038,N_1324);
or U3008 (N_3008,N_418,N_1585);
and U3009 (N_3009,N_2355,N_1444);
nand U3010 (N_3010,N_882,N_956);
nand U3011 (N_3011,N_2345,N_845);
and U3012 (N_3012,N_1942,N_1756);
xor U3013 (N_3013,N_50,N_843);
nor U3014 (N_3014,N_68,N_1015);
xnor U3015 (N_3015,N_496,N_1907);
nand U3016 (N_3016,N_1239,N_1543);
and U3017 (N_3017,N_2309,N_227);
nor U3018 (N_3018,N_2356,N_935);
nor U3019 (N_3019,N_1493,N_1709);
xnor U3020 (N_3020,N_92,N_2459);
and U3021 (N_3021,N_936,N_404);
xnor U3022 (N_3022,N_396,N_1167);
or U3023 (N_3023,N_2347,N_40);
or U3024 (N_3024,N_815,N_2036);
and U3025 (N_3025,N_1438,N_1236);
xor U3026 (N_3026,N_2287,N_1507);
nor U3027 (N_3027,N_1937,N_1570);
xor U3028 (N_3028,N_1951,N_1995);
or U3029 (N_3029,N_1371,N_1773);
or U3030 (N_3030,N_1267,N_1376);
or U3031 (N_3031,N_43,N_327);
and U3032 (N_3032,N_1030,N_2273);
and U3033 (N_3033,N_1067,N_1478);
or U3034 (N_3034,N_2232,N_968);
xnor U3035 (N_3035,N_982,N_2004);
or U3036 (N_3036,N_551,N_1393);
and U3037 (N_3037,N_435,N_1812);
xor U3038 (N_3038,N_1157,N_675);
xnor U3039 (N_3039,N_2462,N_1821);
and U3040 (N_3040,N_318,N_741);
xor U3041 (N_3041,N_1280,N_292);
xor U3042 (N_3042,N_953,N_1908);
and U3043 (N_3043,N_569,N_2033);
nor U3044 (N_3044,N_346,N_1461);
nand U3045 (N_3045,N_143,N_1480);
and U3046 (N_3046,N_705,N_1177);
nor U3047 (N_3047,N_103,N_739);
nand U3048 (N_3048,N_1748,N_38);
xor U3049 (N_3049,N_2230,N_1437);
or U3050 (N_3050,N_726,N_28);
and U3051 (N_3051,N_1397,N_2468);
and U3052 (N_3052,N_641,N_336);
nor U3053 (N_3053,N_609,N_1136);
nand U3054 (N_3054,N_455,N_394);
nor U3055 (N_3055,N_2279,N_990);
xnor U3056 (N_3056,N_2489,N_1453);
nor U3057 (N_3057,N_1649,N_32);
nor U3058 (N_3058,N_1672,N_15);
nand U3059 (N_3059,N_1554,N_1550);
and U3060 (N_3060,N_1227,N_775);
xor U3061 (N_3061,N_270,N_75);
and U3062 (N_3062,N_1089,N_685);
nor U3063 (N_3063,N_2090,N_981);
nor U3064 (N_3064,N_2281,N_745);
and U3065 (N_3065,N_2440,N_2322);
nand U3066 (N_3066,N_2487,N_1882);
nand U3067 (N_3067,N_1540,N_842);
and U3068 (N_3068,N_695,N_1073);
nand U3069 (N_3069,N_269,N_475);
or U3070 (N_3070,N_2152,N_1188);
and U3071 (N_3071,N_1336,N_797);
and U3072 (N_3072,N_2478,N_1080);
or U3073 (N_3073,N_759,N_2131);
nand U3074 (N_3074,N_997,N_1410);
nor U3075 (N_3075,N_2147,N_1729);
and U3076 (N_3076,N_621,N_1778);
xnor U3077 (N_3077,N_1760,N_519);
xnor U3078 (N_3078,N_1346,N_1924);
xor U3079 (N_3079,N_1435,N_646);
or U3080 (N_3080,N_1814,N_238);
nand U3081 (N_3081,N_1068,N_312);
or U3082 (N_3082,N_283,N_1257);
or U3083 (N_3083,N_1476,N_1296);
nand U3084 (N_3084,N_177,N_74);
and U3085 (N_3085,N_1537,N_1247);
nor U3086 (N_3086,N_1844,N_778);
xor U3087 (N_3087,N_1121,N_1282);
nand U3088 (N_3088,N_1552,N_1365);
xor U3089 (N_3089,N_1496,N_528);
xor U3090 (N_3090,N_1927,N_1187);
nand U3091 (N_3091,N_1232,N_2358);
nor U3092 (N_3092,N_153,N_2337);
xnor U3093 (N_3093,N_838,N_42);
or U3094 (N_3094,N_2113,N_291);
nor U3095 (N_3095,N_1913,N_482);
nand U3096 (N_3096,N_1308,N_1641);
nor U3097 (N_3097,N_1965,N_1256);
or U3098 (N_3098,N_2193,N_1551);
or U3099 (N_3099,N_1583,N_1353);
xnor U3100 (N_3100,N_829,N_2392);
nor U3101 (N_3101,N_1429,N_1560);
nor U3102 (N_3102,N_1572,N_1521);
xor U3103 (N_3103,N_2446,N_611);
nor U3104 (N_3104,N_1573,N_285);
nor U3105 (N_3105,N_275,N_1565);
nand U3106 (N_3106,N_1138,N_89);
or U3107 (N_3107,N_1502,N_1538);
nand U3108 (N_3108,N_1047,N_1086);
nor U3109 (N_3109,N_2244,N_1031);
or U3110 (N_3110,N_576,N_131);
nand U3111 (N_3111,N_957,N_2331);
and U3112 (N_3112,N_1612,N_277);
nor U3113 (N_3113,N_1999,N_323);
and U3114 (N_3114,N_766,N_907);
nand U3115 (N_3115,N_1808,N_1624);
nor U3116 (N_3116,N_1508,N_851);
xnor U3117 (N_3117,N_2028,N_2159);
and U3118 (N_3118,N_2195,N_2156);
or U3119 (N_3119,N_1920,N_2197);
xnor U3120 (N_3120,N_2378,N_433);
and U3121 (N_3121,N_877,N_206);
or U3122 (N_3122,N_1734,N_422);
and U3123 (N_3123,N_257,N_154);
and U3124 (N_3124,N_1829,N_2136);
and U3125 (N_3125,N_1263,N_412);
nor U3126 (N_3126,N_1180,N_963);
nor U3127 (N_3127,N_96,N_1902);
or U3128 (N_3128,N_783,N_1781);
nor U3129 (N_3129,N_1039,N_383);
nor U3130 (N_3130,N_717,N_650);
xor U3131 (N_3131,N_21,N_1504);
xnor U3132 (N_3132,N_2107,N_395);
or U3133 (N_3133,N_1523,N_1307);
and U3134 (N_3134,N_2381,N_1632);
or U3135 (N_3135,N_393,N_138);
xor U3136 (N_3136,N_1607,N_280);
or U3137 (N_3137,N_651,N_1916);
xor U3138 (N_3138,N_195,N_813);
xnor U3139 (N_3139,N_917,N_134);
xnor U3140 (N_3140,N_922,N_708);
and U3141 (N_3141,N_77,N_314);
nand U3142 (N_3142,N_2397,N_2157);
xor U3143 (N_3143,N_1101,N_1557);
nand U3144 (N_3144,N_773,N_2014);
nand U3145 (N_3145,N_497,N_763);
and U3146 (N_3146,N_1413,N_1087);
nor U3147 (N_3147,N_899,N_376);
nand U3148 (N_3148,N_39,N_1243);
xnor U3149 (N_3149,N_2491,N_2054);
or U3150 (N_3150,N_194,N_1634);
nor U3151 (N_3151,N_1513,N_2284);
and U3152 (N_3152,N_2456,N_230);
nand U3153 (N_3153,N_1472,N_716);
nand U3154 (N_3154,N_2080,N_1027);
and U3155 (N_3155,N_117,N_2467);
nor U3156 (N_3156,N_855,N_2146);
or U3157 (N_3157,N_2181,N_198);
and U3158 (N_3158,N_2003,N_1609);
and U3159 (N_3159,N_81,N_1594);
or U3160 (N_3160,N_1220,N_71);
nand U3161 (N_3161,N_2285,N_584);
nand U3162 (N_3162,N_25,N_1150);
nor U3163 (N_3163,N_821,N_2295);
or U3164 (N_3164,N_2026,N_23);
and U3165 (N_3165,N_2161,N_938);
xnor U3166 (N_3166,N_1500,N_209);
xor U3167 (N_3167,N_678,N_1312);
and U3168 (N_3168,N_1610,N_1248);
xor U3169 (N_3169,N_1162,N_1007);
and U3170 (N_3170,N_180,N_234);
and U3171 (N_3171,N_374,N_326);
nand U3172 (N_3172,N_1100,N_663);
nor U3173 (N_3173,N_381,N_1225);
and U3174 (N_3174,N_2262,N_1588);
and U3175 (N_3175,N_1387,N_2332);
nand U3176 (N_3176,N_1345,N_100);
nand U3177 (N_3177,N_2225,N_2280);
nor U3178 (N_3178,N_245,N_1139);
and U3179 (N_3179,N_1702,N_99);
nor U3180 (N_3180,N_1764,N_720);
nand U3181 (N_3181,N_273,N_98);
xnor U3182 (N_3182,N_1931,N_1095);
nor U3183 (N_3183,N_515,N_518);
xnor U3184 (N_3184,N_1745,N_1528);
or U3185 (N_3185,N_197,N_1362);
xnor U3186 (N_3186,N_1129,N_1302);
nor U3187 (N_3187,N_2219,N_2267);
and U3188 (N_3188,N_1592,N_2452);
or U3189 (N_3189,N_301,N_1794);
nor U3190 (N_3190,N_2064,N_2365);
nor U3191 (N_3191,N_1448,N_185);
xnor U3192 (N_3192,N_1113,N_35);
or U3193 (N_3193,N_135,N_2148);
xnor U3194 (N_3194,N_1043,N_493);
and U3195 (N_3195,N_891,N_1123);
or U3196 (N_3196,N_1051,N_856);
and U3197 (N_3197,N_414,N_524);
xnor U3198 (N_3198,N_2439,N_307);
xnor U3199 (N_3199,N_2423,N_1374);
nand U3200 (N_3200,N_1151,N_2339);
nand U3201 (N_3201,N_615,N_1084);
or U3202 (N_3202,N_1298,N_1718);
and U3203 (N_3203,N_368,N_173);
and U3204 (N_3204,N_2494,N_998);
xnor U3205 (N_3205,N_2432,N_2463);
nand U3206 (N_3206,N_1988,N_625);
nor U3207 (N_3207,N_757,N_1562);
and U3208 (N_3208,N_1529,N_358);
or U3209 (N_3209,N_1991,N_1404);
and U3210 (N_3210,N_53,N_976);
xor U3211 (N_3211,N_2079,N_1871);
nor U3212 (N_3212,N_401,N_970);
or U3213 (N_3213,N_792,N_1947);
nor U3214 (N_3214,N_921,N_1869);
and U3215 (N_3215,N_2283,N_1485);
and U3216 (N_3216,N_1686,N_2012);
or U3217 (N_3217,N_669,N_1313);
nor U3218 (N_3218,N_247,N_2316);
and U3219 (N_3219,N_1575,N_696);
and U3220 (N_3220,N_1789,N_2186);
and U3221 (N_3221,N_2465,N_420);
nor U3222 (N_3222,N_1475,N_299);
and U3223 (N_3223,N_4,N_605);
or U3224 (N_3224,N_133,N_1854);
nor U3225 (N_3225,N_683,N_1711);
nor U3226 (N_3226,N_2170,N_1074);
or U3227 (N_3227,N_421,N_320);
nor U3228 (N_3228,N_2370,N_199);
nor U3229 (N_3229,N_1412,N_1452);
and U3230 (N_3230,N_1273,N_1677);
and U3231 (N_3231,N_1862,N_736);
or U3232 (N_3232,N_1771,N_1739);
nor U3233 (N_3233,N_1717,N_1860);
nor U3234 (N_3234,N_1310,N_1119);
xnor U3235 (N_3235,N_179,N_2060);
or U3236 (N_3236,N_73,N_737);
or U3237 (N_3237,N_155,N_1899);
nor U3238 (N_3238,N_17,N_399);
nand U3239 (N_3239,N_1315,N_2305);
or U3240 (N_3240,N_1992,N_1432);
xor U3241 (N_3241,N_172,N_2173);
and U3242 (N_3242,N_2143,N_1901);
nand U3243 (N_3243,N_1621,N_2493);
xor U3244 (N_3244,N_105,N_2234);
or U3245 (N_3245,N_634,N_464);
and U3246 (N_3246,N_372,N_1940);
nor U3247 (N_3247,N_895,N_1698);
nand U3248 (N_3248,N_1040,N_578);
xnor U3249 (N_3249,N_1997,N_352);
and U3250 (N_3250,N_959,N_2164);
nand U3251 (N_3251,N_559,N_11);
xnor U3252 (N_3252,N_380,N_1465);
xor U3253 (N_3253,N_755,N_1865);
nand U3254 (N_3254,N_27,N_120);
nor U3255 (N_3255,N_608,N_2172);
and U3256 (N_3256,N_2414,N_2179);
and U3257 (N_3257,N_1290,N_1737);
or U3258 (N_3258,N_945,N_140);
nand U3259 (N_3259,N_1174,N_1373);
or U3260 (N_3260,N_2313,N_1720);
or U3261 (N_3261,N_452,N_929);
xnor U3262 (N_3262,N_1384,N_593);
or U3263 (N_3263,N_114,N_2435);
nand U3264 (N_3264,N_598,N_1034);
or U3265 (N_3265,N_2127,N_1517);
nand U3266 (N_3266,N_2114,N_501);
nand U3267 (N_3267,N_1738,N_123);
nand U3268 (N_3268,N_142,N_863);
or U3269 (N_3269,N_1358,N_1775);
and U3270 (N_3270,N_752,N_2245);
xor U3271 (N_3271,N_2150,N_363);
xnor U3272 (N_3272,N_215,N_2155);
or U3273 (N_3273,N_343,N_110);
nand U3274 (N_3274,N_1368,N_580);
nand U3275 (N_3275,N_1721,N_2051);
and U3276 (N_3276,N_2110,N_2258);
and U3277 (N_3277,N_2049,N_1945);
xor U3278 (N_3278,N_742,N_2217);
and U3279 (N_3279,N_587,N_1386);
xnor U3280 (N_3280,N_711,N_127);
nand U3281 (N_3281,N_2318,N_627);
nand U3282 (N_3282,N_1137,N_747);
nand U3283 (N_3283,N_2075,N_293);
and U3284 (N_3284,N_1460,N_2165);
or U3285 (N_3285,N_1470,N_1785);
or U3286 (N_3286,N_529,N_328);
nand U3287 (N_3287,N_927,N_483);
and U3288 (N_3288,N_1788,N_2101);
nor U3289 (N_3289,N_2319,N_137);
nand U3290 (N_3290,N_508,N_1694);
nor U3291 (N_3291,N_242,N_220);
and U3292 (N_3292,N_1866,N_888);
nor U3293 (N_3293,N_2034,N_2210);
nand U3294 (N_3294,N_1183,N_1810);
nand U3295 (N_3295,N_1880,N_1311);
nor U3296 (N_3296,N_1281,N_542);
nand U3297 (N_3297,N_2457,N_1482);
nand U3298 (N_3298,N_2069,N_2472);
nor U3299 (N_3299,N_1665,N_2451);
nand U3300 (N_3300,N_530,N_1146);
and U3301 (N_3301,N_1597,N_2174);
or U3302 (N_3302,N_2207,N_1769);
nor U3303 (N_3303,N_1367,N_560);
nor U3304 (N_3304,N_1802,N_788);
nor U3305 (N_3305,N_565,N_1824);
and U3306 (N_3306,N_782,N_1484);
and U3307 (N_3307,N_1490,N_2189);
nor U3308 (N_3308,N_1674,N_2009);
and U3309 (N_3309,N_1421,N_1830);
and U3310 (N_3310,N_1110,N_514);
nor U3311 (N_3311,N_819,N_1226);
xnor U3312 (N_3312,N_54,N_1335);
nand U3313 (N_3313,N_1052,N_190);
xor U3314 (N_3314,N_389,N_1449);
or U3315 (N_3315,N_2023,N_1270);
nor U3316 (N_3316,N_1118,N_668);
xor U3317 (N_3317,N_129,N_730);
or U3318 (N_3318,N_513,N_986);
xnor U3319 (N_3319,N_2419,N_1874);
and U3320 (N_3320,N_1426,N_1541);
and U3321 (N_3321,N_1198,N_1548);
and U3322 (N_3322,N_1662,N_1574);
and U3323 (N_3323,N_1318,N_2417);
and U3324 (N_3324,N_1930,N_2418);
xnor U3325 (N_3325,N_876,N_2426);
xnor U3326 (N_3326,N_2483,N_79);
or U3327 (N_3327,N_1228,N_751);
or U3328 (N_3328,N_1466,N_437);
and U3329 (N_3329,N_713,N_1053);
or U3330 (N_3330,N_691,N_1938);
and U3331 (N_3331,N_2326,N_132);
nor U3332 (N_3332,N_189,N_446);
and U3333 (N_3333,N_1998,N_1837);
nand U3334 (N_3334,N_848,N_2372);
and U3335 (N_3335,N_1595,N_1784);
and U3336 (N_3336,N_1985,N_1768);
xor U3337 (N_3337,N_570,N_734);
xnor U3338 (N_3338,N_1935,N_2449);
xnor U3339 (N_3339,N_2366,N_47);
and U3340 (N_3340,N_1713,N_122);
or U3341 (N_3341,N_1231,N_579);
nor U3342 (N_3342,N_537,N_2254);
and U3343 (N_3343,N_1141,N_672);
or U3344 (N_3344,N_1260,N_1450);
nor U3345 (N_3345,N_2039,N_251);
and U3346 (N_3346,N_807,N_1569);
and U3347 (N_3347,N_1342,N_1680);
nand U3348 (N_3348,N_78,N_2011);
xnor U3349 (N_3349,N_319,N_1077);
xor U3350 (N_3350,N_1807,N_322);
nand U3351 (N_3351,N_491,N_867);
or U3352 (N_3352,N_2002,N_1556);
or U3353 (N_3353,N_416,N_1175);
xor U3354 (N_3354,N_1325,N_1705);
and U3355 (N_3355,N_362,N_167);
xor U3356 (N_3356,N_22,N_2275);
xnor U3357 (N_3357,N_2443,N_1872);
nand U3358 (N_3358,N_63,N_2124);
nor U3359 (N_3359,N_2373,N_1555);
xor U3360 (N_3360,N_1,N_1923);
xnor U3361 (N_3361,N_2393,N_790);
nor U3362 (N_3362,N_687,N_2437);
xor U3363 (N_3363,N_591,N_673);
xor U3364 (N_3364,N_2479,N_439);
nor U3365 (N_3365,N_2203,N_900);
and U3366 (N_3366,N_37,N_119);
nor U3367 (N_3367,N_2359,N_417);
or U3368 (N_3368,N_2166,N_642);
nand U3369 (N_3369,N_1293,N_659);
nor U3370 (N_3370,N_1033,N_662);
or U3371 (N_3371,N_2214,N_434);
nor U3372 (N_3372,N_1666,N_1905);
nand U3373 (N_3373,N_1783,N_951);
or U3374 (N_3374,N_2106,N_1462);
nor U3375 (N_3375,N_1972,N_2352);
and U3376 (N_3376,N_1361,N_803);
and U3377 (N_3377,N_973,N_898);
nand U3378 (N_3378,N_1446,N_2015);
xor U3379 (N_3379,N_1094,N_808);
nor U3380 (N_3380,N_205,N_706);
nand U3381 (N_3381,N_65,N_1746);
nor U3382 (N_3382,N_729,N_1143);
nor U3383 (N_3383,N_762,N_297);
nor U3384 (N_3384,N_1596,N_85);
nand U3385 (N_3385,N_964,N_880);
nor U3386 (N_3386,N_1377,N_1057);
xnor U3387 (N_3387,N_592,N_1004);
xor U3388 (N_3388,N_826,N_2441);
or U3389 (N_3389,N_2390,N_2029);
xnor U3390 (N_3390,N_1014,N_1168);
and U3391 (N_3391,N_881,N_1405);
and U3392 (N_3392,N_1611,N_1012);
nor U3393 (N_3393,N_798,N_768);
nand U3394 (N_3394,N_586,N_988);
and U3395 (N_3395,N_405,N_1217);
xnor U3396 (N_3396,N_2216,N_661);
xor U3397 (N_3397,N_1915,N_1759);
and U3398 (N_3398,N_13,N_1375);
nand U3399 (N_3399,N_235,N_1163);
nor U3400 (N_3400,N_2133,N_1801);
nor U3401 (N_3401,N_2109,N_831);
nor U3402 (N_3402,N_2425,N_1409);
xnor U3403 (N_3403,N_1291,N_955);
or U3404 (N_3404,N_566,N_1222);
xor U3405 (N_3405,N_1114,N_1943);
or U3406 (N_3406,N_1434,N_33);
or U3407 (N_3407,N_1126,N_1285);
or U3408 (N_3408,N_1364,N_130);
nor U3409 (N_3409,N_1411,N_597);
nand U3410 (N_3410,N_791,N_913);
or U3411 (N_3411,N_338,N_402);
nor U3412 (N_3412,N_1968,N_1333);
and U3413 (N_3413,N_1870,N_649);
and U3414 (N_3414,N_10,N_1436);
or U3415 (N_3415,N_1214,N_440);
nand U3416 (N_3416,N_887,N_1777);
and U3417 (N_3417,N_1076,N_2066);
nor U3418 (N_3418,N_697,N_1767);
nand U3419 (N_3419,N_1982,N_1567);
or U3420 (N_3420,N_700,N_1058);
xnor U3421 (N_3421,N_1501,N_1292);
or U3422 (N_3422,N_1441,N_2222);
nor U3423 (N_3423,N_1636,N_1055);
or U3424 (N_3424,N_324,N_151);
xnor U3425 (N_3425,N_2348,N_606);
or U3426 (N_3426,N_858,N_1322);
nor U3427 (N_3427,N_1971,N_999);
xor U3428 (N_3428,N_357,N_453);
nand U3429 (N_3429,N_1741,N_2196);
nor U3430 (N_3430,N_2268,N_1305);
nand U3431 (N_3431,N_26,N_2111);
or U3432 (N_3432,N_413,N_1600);
and U3433 (N_3433,N_1201,N_1160);
and U3434 (N_3434,N_1330,N_1061);
or U3435 (N_3435,N_1793,N_1603);
xnor U3436 (N_3436,N_725,N_732);
nand U3437 (N_3437,N_1140,N_617);
xnor U3438 (N_3438,N_1378,N_879);
nor U3439 (N_3439,N_897,N_1618);
xor U3440 (N_3440,N_1889,N_157);
nor U3441 (N_3441,N_835,N_714);
or U3442 (N_3442,N_655,N_1990);
nor U3443 (N_3443,N_1954,N_2482);
xor U3444 (N_3444,N_1629,N_2047);
nor U3445 (N_3445,N_1133,N_45);
and U3446 (N_3446,N_1192,N_789);
and U3447 (N_3447,N_1744,N_950);
xor U3448 (N_3448,N_313,N_1251);
nor U3449 (N_3449,N_2067,N_2351);
and U3450 (N_3450,N_924,N_449);
xor U3451 (N_3451,N_1062,N_1526);
and U3452 (N_3452,N_1772,N_983);
or U3453 (N_3453,N_1091,N_1921);
or U3454 (N_3454,N_1714,N_776);
and U3455 (N_3455,N_1090,N_477);
nand U3456 (N_3456,N_1659,N_2108);
and U3457 (N_3457,N_2307,N_1083);
or U3458 (N_3458,N_367,N_2455);
and U3459 (N_3459,N_317,N_1853);
xor U3460 (N_3460,N_2333,N_459);
or U3461 (N_3461,N_1986,N_967);
nor U3462 (N_3462,N_760,N_115);
and U3463 (N_3463,N_2407,N_0);
nand U3464 (N_3464,N_348,N_1799);
nand U3465 (N_3465,N_1977,N_1582);
nor U3466 (N_3466,N_2144,N_2416);
nor U3467 (N_3467,N_1828,N_1017);
nand U3468 (N_3468,N_2018,N_2132);
nor U3469 (N_3469,N_2138,N_384);
nand U3470 (N_3470,N_1984,N_1124);
or U3471 (N_3471,N_222,N_2212);
nor U3472 (N_3472,N_624,N_148);
xor U3473 (N_3473,N_391,N_256);
xor U3474 (N_3474,N_794,N_344);
or U3475 (N_3475,N_1546,N_2046);
or U3476 (N_3476,N_2458,N_1408);
xnor U3477 (N_3477,N_48,N_1941);
xnor U3478 (N_3478,N_2182,N_2062);
nand U3479 (N_3479,N_196,N_2153);
nand U3480 (N_3480,N_1606,N_1155);
or U3481 (N_3481,N_1900,N_361);
and U3482 (N_3482,N_2485,N_2349);
and U3483 (N_3483,N_864,N_1974);
nor U3484 (N_3484,N_484,N_1660);
xnor U3485 (N_3485,N_304,N_2428);
or U3486 (N_3486,N_249,N_1819);
or U3487 (N_3487,N_1447,N_1533);
and U3488 (N_3488,N_1259,N_1096);
nor U3489 (N_3489,N_355,N_1658);
or U3490 (N_3490,N_1468,N_969);
and U3491 (N_3491,N_1316,N_1623);
nor U3492 (N_3492,N_2354,N_2481);
or U3493 (N_3493,N_2430,N_1195);
or U3494 (N_3494,N_1728,N_159);
nor U3495 (N_3495,N_349,N_1178);
and U3496 (N_3496,N_769,N_585);
or U3497 (N_3497,N_2382,N_139);
and U3498 (N_3498,N_169,N_743);
xor U3499 (N_3499,N_939,N_595);
nand U3500 (N_3500,N_507,N_353);
nand U3501 (N_3501,N_2336,N_638);
nor U3502 (N_3502,N_2180,N_480);
or U3503 (N_3503,N_1166,N_1743);
nor U3504 (N_3504,N_2403,N_1663);
nand U3505 (N_3505,N_1349,N_1264);
xnor U3506 (N_3506,N_539,N_2346);
and U3507 (N_3507,N_2117,N_2096);
nor U3508 (N_3508,N_816,N_865);
or U3509 (N_3509,N_1202,N_679);
nand U3510 (N_3510,N_1474,N_731);
or U3511 (N_3511,N_232,N_653);
nor U3512 (N_3512,N_2102,N_1620);
and U3513 (N_3513,N_2246,N_1127);
or U3514 (N_3514,N_2123,N_1344);
nor U3515 (N_3515,N_82,N_375);
or U3516 (N_3516,N_568,N_223);
and U3517 (N_3517,N_1357,N_538);
nor U3518 (N_3518,N_1495,N_1886);
and U3519 (N_3519,N_2250,N_359);
nor U3520 (N_3520,N_1532,N_1038);
nand U3521 (N_3521,N_1494,N_666);
xnor U3522 (N_3522,N_1135,N_266);
nand U3523 (N_3523,N_121,N_2105);
and U3524 (N_3524,N_58,N_1300);
nand U3525 (N_3525,N_241,N_977);
nand U3526 (N_3526,N_1640,N_2241);
xnor U3527 (N_3527,N_259,N_2145);
nand U3528 (N_3528,N_1885,N_1396);
nor U3529 (N_3529,N_1622,N_2317);
nor U3530 (N_3530,N_1024,N_1961);
xor U3531 (N_3531,N_144,N_201);
nand U3532 (N_3532,N_1966,N_2194);
and U3533 (N_3533,N_2367,N_892);
or U3534 (N_3534,N_2471,N_884);
nor U3535 (N_3535,N_2464,N_954);
or U3536 (N_3536,N_2078,N_436);
or U3537 (N_3537,N_456,N_2269);
and U3538 (N_3538,N_2027,N_1651);
nor U3539 (N_3539,N_1693,N_2409);
xor U3540 (N_3540,N_2408,N_162);
nor U3541 (N_3541,N_295,N_310);
nand U3542 (N_3542,N_462,N_1723);
and U3543 (N_3543,N_1295,N_1477);
and U3544 (N_3544,N_1571,N_340);
or U3545 (N_3545,N_908,N_859);
nand U3546 (N_3546,N_1369,N_2497);
nor U3547 (N_3547,N_94,N_1383);
nor U3548 (N_3548,N_1148,N_926);
nand U3549 (N_3549,N_1171,N_1561);
nand U3550 (N_3550,N_728,N_1142);
and U3551 (N_3551,N_1973,N_118);
nand U3552 (N_3552,N_1544,N_1835);
xnor U3553 (N_3553,N_1104,N_689);
xor U3554 (N_3554,N_1751,N_165);
and U3555 (N_3555,N_1608,N_941);
and U3556 (N_3556,N_1210,N_2413);
nor U3557 (N_3557,N_1676,N_345);
nand U3558 (N_3558,N_2,N_2140);
or U3559 (N_3559,N_438,N_161);
nand U3560 (N_3560,N_2453,N_1696);
nand U3561 (N_3561,N_186,N_1355);
and U3562 (N_3562,N_18,N_610);
xor U3563 (N_3563,N_1266,N_2304);
xor U3564 (N_3564,N_572,N_1182);
or U3565 (N_3565,N_1111,N_2310);
xor U3566 (N_3566,N_561,N_1063);
and U3567 (N_3567,N_2248,N_1505);
xor U3568 (N_3568,N_261,N_451);
xnor U3569 (N_3569,N_682,N_1682);
nor U3570 (N_3570,N_427,N_489);
xnor U3571 (N_3571,N_2412,N_1392);
and U3572 (N_3572,N_581,N_787);
nand U3573 (N_3573,N_1875,N_62);
nand U3574 (N_3574,N_2206,N_2226);
and U3575 (N_3575,N_1066,N_847);
nor U3576 (N_3576,N_1002,N_1615);
xor U3577 (N_3577,N_211,N_870);
xor U3578 (N_3578,N_1173,N_1904);
and U3579 (N_3579,N_660,N_463);
nand U3580 (N_3580,N_1605,N_311);
nor U3581 (N_3581,N_1319,N_522);
xor U3582 (N_3582,N_1840,N_521);
and U3583 (N_3583,N_2330,N_836);
nor U3584 (N_3584,N_670,N_1328);
nand U3585 (N_3585,N_1626,N_1779);
nand U3586 (N_3586,N_1834,N_1046);
xnor U3587 (N_3587,N_872,N_325);
and U3588 (N_3588,N_1390,N_360);
nor U3589 (N_3589,N_920,N_224);
and U3590 (N_3590,N_2116,N_46);
and U3591 (N_3591,N_520,N_67);
nor U3592 (N_3592,N_733,N_2037);
nor U3593 (N_3593,N_686,N_1531);
xor U3594 (N_3594,N_1213,N_193);
and U3595 (N_3595,N_290,N_2427);
nor U3596 (N_3596,N_2260,N_942);
nor U3597 (N_3597,N_2386,N_1488);
nor U3598 (N_3598,N_1515,N_12);
nand U3599 (N_3599,N_44,N_86);
nand U3600 (N_3600,N_1021,N_2162);
nand U3601 (N_3601,N_588,N_254);
nor U3602 (N_3602,N_1306,N_2401);
xnor U3603 (N_3603,N_2024,N_721);
nor U3604 (N_3604,N_1704,N_1836);
xnor U3605 (N_3605,N_1707,N_1204);
nand U3606 (N_3606,N_2422,N_774);
or U3607 (N_3607,N_896,N_1380);
xor U3608 (N_3608,N_1813,N_1382);
and U3609 (N_3609,N_1843,N_146);
or U3610 (N_3610,N_1161,N_14);
and U3611 (N_3611,N_1321,N_2396);
or U3612 (N_3612,N_749,N_1001);
and U3613 (N_3613,N_1826,N_722);
xnor U3614 (N_3614,N_993,N_2252);
nand U3615 (N_3615,N_252,N_1184);
and U3616 (N_3616,N_1492,N_933);
or U3617 (N_3617,N_704,N_2169);
nor U3618 (N_3618,N_109,N_630);
and U3619 (N_3619,N_2224,N_883);
and U3620 (N_3620,N_2259,N_1638);
and U3621 (N_3621,N_910,N_1817);
or U3622 (N_3622,N_2328,N_1894);
nand U3623 (N_3623,N_2068,N_1423);
nand U3624 (N_3624,N_868,N_29);
and U3625 (N_3625,N_1064,N_5);
nand U3626 (N_3626,N_2486,N_1020);
nand U3627 (N_3627,N_1498,N_1018);
or U3628 (N_3628,N_1762,N_1825);
and U3629 (N_3629,N_1218,N_992);
and U3630 (N_3630,N_188,N_2466);
nand U3631 (N_3631,N_2363,N_2384);
and U3632 (N_3632,N_785,N_886);
nor U3633 (N_3633,N_225,N_1417);
or U3634 (N_3634,N_1334,N_315);
nor U3635 (N_3635,N_1360,N_916);
or U3636 (N_3636,N_1688,N_2376);
and U3637 (N_3637,N_2266,N_1144);
nand U3638 (N_3638,N_1564,N_124);
nor U3639 (N_3639,N_541,N_771);
or U3640 (N_3640,N_1372,N_1112);
or U3641 (N_3641,N_2048,N_656);
nor U3642 (N_3642,N_203,N_1864);
xnor U3643 (N_3643,N_1892,N_1936);
nor U3644 (N_3644,N_1796,N_2300);
nor U3645 (N_3645,N_1953,N_1238);
nand U3646 (N_3646,N_812,N_1859);
xor U3647 (N_3647,N_2364,N_2256);
nor U3648 (N_3648,N_1809,N_1922);
nand U3649 (N_3649,N_2213,N_846);
or U3650 (N_3650,N_2220,N_601);
nand U3651 (N_3651,N_535,N_1116);
or U3652 (N_3652,N_1486,N_400);
nand U3653 (N_3653,N_236,N_2237);
nand U3654 (N_3654,N_2139,N_600);
and U3655 (N_3655,N_680,N_2142);
nand U3656 (N_3656,N_837,N_1946);
nor U3657 (N_3657,N_818,N_1958);
or U3658 (N_3658,N_761,N_1255);
and U3659 (N_3659,N_632,N_246);
and U3660 (N_3660,N_479,N_1960);
or U3661 (N_3661,N_1983,N_1766);
and U3662 (N_3662,N_1602,N_309);
and U3663 (N_3663,N_1970,N_369);
nand U3664 (N_3664,N_972,N_1827);
nor U3665 (N_3665,N_602,N_971);
and U3666 (N_3666,N_9,N_76);
nand U3667 (N_3667,N_849,N_2185);
nor U3668 (N_3668,N_409,N_966);
nor U3669 (N_3669,N_1035,N_2288);
and U3670 (N_3670,N_1510,N_329);
or U3671 (N_3671,N_1506,N_1414);
nand U3672 (N_3672,N_1850,N_1747);
xnor U3673 (N_3673,N_915,N_2474);
or U3674 (N_3674,N_1326,N_1272);
or U3675 (N_3675,N_639,N_2171);
nor U3676 (N_3676,N_2338,N_1147);
or U3677 (N_3677,N_2255,N_985);
xor U3678 (N_3678,N_574,N_1301);
nor U3679 (N_3679,N_718,N_128);
or U3680 (N_3680,N_1288,N_2293);
and U3681 (N_3681,N_289,N_671);
xor U3682 (N_3682,N_548,N_149);
nor U3683 (N_3683,N_1855,N_244);
nor U3684 (N_3684,N_619,N_547);
and U3685 (N_3685,N_2377,N_2104);
nand U3686 (N_3686,N_1149,N_1661);
nand U3687 (N_3687,N_1800,N_629);
nand U3688 (N_3688,N_2065,N_2395);
nand U3689 (N_3689,N_443,N_1108);
or U3690 (N_3690,N_830,N_152);
and U3691 (N_3691,N_1601,N_1128);
and U3692 (N_3692,N_911,N_2380);
nand U3693 (N_3693,N_647,N_1816);
and U3694 (N_3694,N_750,N_1733);
or U3695 (N_3695,N_1841,N_2477);
nor U3696 (N_3696,N_2115,N_2420);
xnor U3697 (N_3697,N_3,N_2282);
or U3698 (N_3698,N_1839,N_1805);
xor U3699 (N_3699,N_2020,N_356);
xnor U3700 (N_3700,N_377,N_255);
xnor U3701 (N_3701,N_276,N_2360);
nor U3702 (N_3702,N_1613,N_1664);
or U3703 (N_3703,N_1631,N_1509);
nand U3704 (N_3704,N_2022,N_213);
xor U3705 (N_3705,N_136,N_208);
nand U3706 (N_3706,N_1867,N_862);
or U3707 (N_3707,N_2400,N_1987);
xor U3708 (N_3708,N_1209,N_1752);
nand U3709 (N_3709,N_2091,N_2030);
xnor U3710 (N_3710,N_2243,N_962);
nand U3711 (N_3711,N_1240,N_2278);
or U3712 (N_3712,N_1976,N_2404);
or U3713 (N_3713,N_2005,N_1289);
and U3714 (N_3714,N_1026,N_2274);
and U3715 (N_3715,N_2410,N_1078);
and U3716 (N_3716,N_1297,N_2006);
or U3717 (N_3717,N_948,N_828);
nor U3718 (N_3718,N_51,N_889);
or U3719 (N_3719,N_780,N_1716);
and U3720 (N_3720,N_112,N_1379);
xnor U3721 (N_3721,N_875,N_2362);
and U3722 (N_3722,N_2041,N_1366);
or U3723 (N_3723,N_1644,N_1852);
xnor U3724 (N_3724,N_1925,N_34);
xnor U3725 (N_3725,N_1919,N_191);
and U3726 (N_3726,N_709,N_1491);
nand U3727 (N_3727,N_1154,N_2151);
nor U3728 (N_3728,N_2251,N_753);
and U3729 (N_3729,N_1036,N_1283);
nand U3730 (N_3730,N_1419,N_2327);
and U3731 (N_3731,N_1451,N_61);
xnor U3732 (N_3732,N_1130,N_1534);
and U3733 (N_3733,N_703,N_2374);
nor U3734 (N_3734,N_2088,N_827);
xor U3735 (N_3735,N_1683,N_644);
nor U3736 (N_3736,N_1820,N_271);
and U3737 (N_3737,N_1962,N_253);
nor U3738 (N_3738,N_1678,N_379);
nor U3739 (N_3739,N_2183,N_832);
nor U3740 (N_3740,N_1692,N_590);
xnor U3741 (N_3741,N_467,N_2368);
and U3742 (N_3742,N_1689,N_536);
and U3743 (N_3743,N_1635,N_2429);
or U3744 (N_3744,N_450,N_183);
and U3745 (N_3745,N_1803,N_226);
xor U3746 (N_3746,N_2149,N_1422);
xor U3747 (N_3747,N_1274,N_869);
or U3748 (N_3748,N_1742,N_1795);
nor U3749 (N_3749,N_2311,N_767);
nand U3750 (N_3750,N_2391,N_2407);
and U3751 (N_3751,N_1821,N_980);
nand U3752 (N_3752,N_1428,N_6);
or U3753 (N_3753,N_2413,N_2176);
nor U3754 (N_3754,N_2167,N_2484);
and U3755 (N_3755,N_1142,N_723);
or U3756 (N_3756,N_2396,N_1837);
nor U3757 (N_3757,N_808,N_1027);
or U3758 (N_3758,N_795,N_1732);
and U3759 (N_3759,N_1898,N_843);
nor U3760 (N_3760,N_2444,N_2256);
or U3761 (N_3761,N_2231,N_617);
nor U3762 (N_3762,N_1482,N_2134);
nor U3763 (N_3763,N_2172,N_754);
and U3764 (N_3764,N_1908,N_1276);
or U3765 (N_3765,N_1672,N_165);
xnor U3766 (N_3766,N_1620,N_1164);
or U3767 (N_3767,N_43,N_1428);
or U3768 (N_3768,N_1918,N_1112);
nand U3769 (N_3769,N_693,N_1894);
and U3770 (N_3770,N_2166,N_780);
nand U3771 (N_3771,N_2383,N_526);
or U3772 (N_3772,N_2484,N_1636);
nor U3773 (N_3773,N_1077,N_1676);
nand U3774 (N_3774,N_1999,N_922);
xnor U3775 (N_3775,N_2233,N_671);
nand U3776 (N_3776,N_1101,N_606);
and U3777 (N_3777,N_1840,N_297);
xnor U3778 (N_3778,N_2404,N_1065);
xnor U3779 (N_3779,N_1782,N_2373);
or U3780 (N_3780,N_1562,N_784);
or U3781 (N_3781,N_1505,N_1617);
xor U3782 (N_3782,N_1140,N_1539);
or U3783 (N_3783,N_855,N_827);
xnor U3784 (N_3784,N_1377,N_1272);
and U3785 (N_3785,N_2077,N_23);
nand U3786 (N_3786,N_684,N_1891);
or U3787 (N_3787,N_1437,N_1693);
nand U3788 (N_3788,N_1619,N_2060);
xor U3789 (N_3789,N_2393,N_9);
and U3790 (N_3790,N_2487,N_2015);
nand U3791 (N_3791,N_786,N_2206);
nor U3792 (N_3792,N_969,N_1592);
nand U3793 (N_3793,N_407,N_993);
xnor U3794 (N_3794,N_1115,N_1247);
or U3795 (N_3795,N_791,N_1003);
and U3796 (N_3796,N_825,N_1179);
xnor U3797 (N_3797,N_1840,N_39);
xnor U3798 (N_3798,N_1696,N_2358);
nand U3799 (N_3799,N_736,N_232);
and U3800 (N_3800,N_993,N_952);
or U3801 (N_3801,N_2338,N_1695);
nor U3802 (N_3802,N_2484,N_1841);
nor U3803 (N_3803,N_683,N_1413);
and U3804 (N_3804,N_2337,N_1526);
or U3805 (N_3805,N_585,N_160);
nor U3806 (N_3806,N_1088,N_208);
nand U3807 (N_3807,N_839,N_2199);
and U3808 (N_3808,N_1069,N_1845);
nand U3809 (N_3809,N_649,N_377);
nor U3810 (N_3810,N_6,N_2004);
or U3811 (N_3811,N_1807,N_2366);
xor U3812 (N_3812,N_386,N_2360);
nor U3813 (N_3813,N_1822,N_798);
nand U3814 (N_3814,N_11,N_372);
and U3815 (N_3815,N_1450,N_632);
and U3816 (N_3816,N_431,N_851);
and U3817 (N_3817,N_223,N_1956);
or U3818 (N_3818,N_1667,N_2419);
and U3819 (N_3819,N_8,N_1229);
or U3820 (N_3820,N_669,N_1450);
xor U3821 (N_3821,N_1764,N_214);
xor U3822 (N_3822,N_1936,N_1567);
or U3823 (N_3823,N_1942,N_161);
nor U3824 (N_3824,N_2272,N_263);
xnor U3825 (N_3825,N_1387,N_1723);
nor U3826 (N_3826,N_208,N_1173);
xor U3827 (N_3827,N_589,N_1056);
xor U3828 (N_3828,N_2437,N_2350);
and U3829 (N_3829,N_1673,N_639);
xnor U3830 (N_3830,N_728,N_1623);
nand U3831 (N_3831,N_936,N_793);
and U3832 (N_3832,N_1869,N_869);
xnor U3833 (N_3833,N_2167,N_2013);
and U3834 (N_3834,N_1499,N_1991);
or U3835 (N_3835,N_1027,N_1527);
nor U3836 (N_3836,N_1948,N_259);
nand U3837 (N_3837,N_2090,N_1871);
and U3838 (N_3838,N_1967,N_930);
nand U3839 (N_3839,N_955,N_614);
and U3840 (N_3840,N_582,N_1464);
and U3841 (N_3841,N_393,N_797);
nand U3842 (N_3842,N_1747,N_1168);
nor U3843 (N_3843,N_1023,N_1755);
nor U3844 (N_3844,N_1293,N_1454);
xnor U3845 (N_3845,N_859,N_2081);
nand U3846 (N_3846,N_622,N_442);
xor U3847 (N_3847,N_1416,N_2128);
nand U3848 (N_3848,N_716,N_990);
nand U3849 (N_3849,N_842,N_1256);
xnor U3850 (N_3850,N_1807,N_450);
xnor U3851 (N_3851,N_905,N_381);
xor U3852 (N_3852,N_927,N_787);
or U3853 (N_3853,N_533,N_738);
or U3854 (N_3854,N_1314,N_851);
and U3855 (N_3855,N_693,N_213);
nand U3856 (N_3856,N_2235,N_1245);
nand U3857 (N_3857,N_622,N_827);
nand U3858 (N_3858,N_1719,N_1968);
or U3859 (N_3859,N_1345,N_1865);
or U3860 (N_3860,N_1222,N_107);
nand U3861 (N_3861,N_2481,N_608);
nand U3862 (N_3862,N_695,N_255);
nor U3863 (N_3863,N_1671,N_1712);
nor U3864 (N_3864,N_1968,N_1383);
and U3865 (N_3865,N_1273,N_123);
and U3866 (N_3866,N_1643,N_1139);
or U3867 (N_3867,N_708,N_1151);
nand U3868 (N_3868,N_1364,N_2033);
and U3869 (N_3869,N_558,N_2422);
nor U3870 (N_3870,N_1865,N_1144);
nand U3871 (N_3871,N_340,N_345);
or U3872 (N_3872,N_1500,N_2384);
nand U3873 (N_3873,N_59,N_1841);
xor U3874 (N_3874,N_1643,N_2049);
nor U3875 (N_3875,N_1397,N_1010);
nor U3876 (N_3876,N_2154,N_2183);
or U3877 (N_3877,N_1730,N_2281);
nor U3878 (N_3878,N_1229,N_1137);
and U3879 (N_3879,N_1304,N_1724);
and U3880 (N_3880,N_681,N_340);
nand U3881 (N_3881,N_404,N_746);
nor U3882 (N_3882,N_309,N_2429);
nand U3883 (N_3883,N_551,N_1239);
and U3884 (N_3884,N_829,N_469);
nand U3885 (N_3885,N_2045,N_1450);
xor U3886 (N_3886,N_1801,N_313);
xor U3887 (N_3887,N_686,N_1168);
nand U3888 (N_3888,N_2067,N_1129);
or U3889 (N_3889,N_2436,N_2394);
and U3890 (N_3890,N_408,N_2316);
nor U3891 (N_3891,N_557,N_563);
or U3892 (N_3892,N_40,N_848);
xnor U3893 (N_3893,N_2094,N_1460);
or U3894 (N_3894,N_700,N_472);
or U3895 (N_3895,N_224,N_1762);
nand U3896 (N_3896,N_57,N_1420);
nand U3897 (N_3897,N_1151,N_559);
nand U3898 (N_3898,N_1045,N_707);
and U3899 (N_3899,N_2200,N_2314);
and U3900 (N_3900,N_728,N_2154);
or U3901 (N_3901,N_1718,N_913);
nand U3902 (N_3902,N_2456,N_1611);
nor U3903 (N_3903,N_1809,N_600);
nor U3904 (N_3904,N_246,N_357);
nor U3905 (N_3905,N_1389,N_923);
and U3906 (N_3906,N_1137,N_2153);
nor U3907 (N_3907,N_905,N_1865);
or U3908 (N_3908,N_2284,N_1999);
or U3909 (N_3909,N_663,N_2291);
nand U3910 (N_3910,N_350,N_2130);
nand U3911 (N_3911,N_1897,N_1437);
xor U3912 (N_3912,N_775,N_1);
xnor U3913 (N_3913,N_2326,N_1672);
nor U3914 (N_3914,N_2229,N_982);
nor U3915 (N_3915,N_1798,N_2264);
or U3916 (N_3916,N_710,N_331);
nand U3917 (N_3917,N_1321,N_328);
and U3918 (N_3918,N_938,N_2123);
and U3919 (N_3919,N_192,N_338);
and U3920 (N_3920,N_1117,N_1023);
nor U3921 (N_3921,N_1622,N_1245);
and U3922 (N_3922,N_878,N_945);
xor U3923 (N_3923,N_23,N_2391);
nor U3924 (N_3924,N_2368,N_1613);
and U3925 (N_3925,N_1896,N_482);
xnor U3926 (N_3926,N_240,N_372);
and U3927 (N_3927,N_874,N_827);
and U3928 (N_3928,N_2401,N_1209);
xor U3929 (N_3929,N_296,N_2063);
nand U3930 (N_3930,N_188,N_1449);
nor U3931 (N_3931,N_2309,N_2077);
nand U3932 (N_3932,N_764,N_888);
nor U3933 (N_3933,N_2404,N_349);
and U3934 (N_3934,N_1306,N_1333);
xor U3935 (N_3935,N_1393,N_2106);
nand U3936 (N_3936,N_495,N_552);
nor U3937 (N_3937,N_181,N_1941);
nor U3938 (N_3938,N_501,N_382);
xnor U3939 (N_3939,N_246,N_1201);
nand U3940 (N_3940,N_181,N_587);
xor U3941 (N_3941,N_1122,N_812);
nand U3942 (N_3942,N_857,N_1725);
nor U3943 (N_3943,N_515,N_187);
xor U3944 (N_3944,N_2417,N_2233);
nor U3945 (N_3945,N_150,N_1762);
nand U3946 (N_3946,N_97,N_1305);
and U3947 (N_3947,N_1274,N_670);
or U3948 (N_3948,N_500,N_1868);
and U3949 (N_3949,N_2097,N_1469);
and U3950 (N_3950,N_2413,N_1195);
nor U3951 (N_3951,N_1947,N_1021);
nor U3952 (N_3952,N_1203,N_449);
xor U3953 (N_3953,N_1415,N_1343);
xor U3954 (N_3954,N_2293,N_166);
nor U3955 (N_3955,N_345,N_2125);
nand U3956 (N_3956,N_1061,N_321);
or U3957 (N_3957,N_674,N_888);
nor U3958 (N_3958,N_185,N_1796);
nor U3959 (N_3959,N_1196,N_1906);
nor U3960 (N_3960,N_88,N_767);
xnor U3961 (N_3961,N_1688,N_2273);
or U3962 (N_3962,N_1058,N_1255);
or U3963 (N_3963,N_256,N_1596);
nand U3964 (N_3964,N_1602,N_289);
or U3965 (N_3965,N_136,N_1749);
nand U3966 (N_3966,N_340,N_828);
xor U3967 (N_3967,N_967,N_226);
xor U3968 (N_3968,N_1032,N_1302);
or U3969 (N_3969,N_474,N_377);
nor U3970 (N_3970,N_1248,N_491);
xnor U3971 (N_3971,N_2169,N_1783);
nor U3972 (N_3972,N_1562,N_180);
xor U3973 (N_3973,N_2104,N_914);
and U3974 (N_3974,N_1228,N_2162);
and U3975 (N_3975,N_2149,N_377);
nand U3976 (N_3976,N_680,N_1980);
nor U3977 (N_3977,N_2232,N_1487);
or U3978 (N_3978,N_1854,N_1949);
nor U3979 (N_3979,N_1268,N_323);
nand U3980 (N_3980,N_1127,N_614);
nor U3981 (N_3981,N_2488,N_1242);
nand U3982 (N_3982,N_903,N_866);
xor U3983 (N_3983,N_1630,N_729);
or U3984 (N_3984,N_1953,N_710);
or U3985 (N_3985,N_964,N_2290);
and U3986 (N_3986,N_1181,N_1356);
or U3987 (N_3987,N_43,N_941);
nand U3988 (N_3988,N_48,N_1700);
nand U3989 (N_3989,N_1609,N_728);
nand U3990 (N_3990,N_243,N_906);
and U3991 (N_3991,N_356,N_104);
nor U3992 (N_3992,N_515,N_458);
nand U3993 (N_3993,N_1600,N_748);
nand U3994 (N_3994,N_156,N_978);
and U3995 (N_3995,N_2179,N_2114);
xor U3996 (N_3996,N_476,N_1006);
nor U3997 (N_3997,N_2138,N_616);
and U3998 (N_3998,N_2109,N_812);
xnor U3999 (N_3999,N_1075,N_1029);
and U4000 (N_4000,N_1068,N_1682);
or U4001 (N_4001,N_1717,N_1071);
nor U4002 (N_4002,N_2192,N_1263);
nand U4003 (N_4003,N_876,N_1150);
xor U4004 (N_4004,N_575,N_1957);
nand U4005 (N_4005,N_2240,N_293);
xnor U4006 (N_4006,N_730,N_131);
nand U4007 (N_4007,N_907,N_234);
and U4008 (N_4008,N_1951,N_1175);
or U4009 (N_4009,N_1409,N_1886);
or U4010 (N_4010,N_812,N_69);
and U4011 (N_4011,N_822,N_747);
nor U4012 (N_4012,N_1625,N_1822);
and U4013 (N_4013,N_94,N_2457);
or U4014 (N_4014,N_1910,N_957);
or U4015 (N_4015,N_568,N_740);
xnor U4016 (N_4016,N_1483,N_1481);
and U4017 (N_4017,N_2334,N_1550);
and U4018 (N_4018,N_1120,N_773);
and U4019 (N_4019,N_29,N_473);
nand U4020 (N_4020,N_717,N_654);
nand U4021 (N_4021,N_1224,N_1797);
xor U4022 (N_4022,N_883,N_2396);
nor U4023 (N_4023,N_1131,N_2336);
xnor U4024 (N_4024,N_2459,N_752);
xnor U4025 (N_4025,N_332,N_1316);
xnor U4026 (N_4026,N_116,N_837);
nand U4027 (N_4027,N_1965,N_265);
xor U4028 (N_4028,N_930,N_311);
nor U4029 (N_4029,N_1198,N_705);
xor U4030 (N_4030,N_1988,N_2489);
or U4031 (N_4031,N_2374,N_2178);
or U4032 (N_4032,N_1933,N_903);
nor U4033 (N_4033,N_2362,N_866);
nand U4034 (N_4034,N_436,N_1335);
nor U4035 (N_4035,N_661,N_2267);
nor U4036 (N_4036,N_188,N_333);
nor U4037 (N_4037,N_844,N_1508);
and U4038 (N_4038,N_975,N_907);
xnor U4039 (N_4039,N_952,N_1830);
or U4040 (N_4040,N_1961,N_1704);
nand U4041 (N_4041,N_1636,N_509);
and U4042 (N_4042,N_2404,N_123);
or U4043 (N_4043,N_753,N_1452);
nand U4044 (N_4044,N_502,N_2475);
and U4045 (N_4045,N_1102,N_718);
nand U4046 (N_4046,N_1321,N_1462);
and U4047 (N_4047,N_1695,N_722);
nand U4048 (N_4048,N_882,N_1150);
xor U4049 (N_4049,N_2346,N_2025);
and U4050 (N_4050,N_2274,N_588);
nand U4051 (N_4051,N_753,N_1629);
or U4052 (N_4052,N_1407,N_1822);
xnor U4053 (N_4053,N_1141,N_2379);
or U4054 (N_4054,N_1744,N_1185);
or U4055 (N_4055,N_51,N_1772);
nor U4056 (N_4056,N_1436,N_1759);
and U4057 (N_4057,N_1954,N_2335);
and U4058 (N_4058,N_2142,N_1467);
and U4059 (N_4059,N_2424,N_2123);
xnor U4060 (N_4060,N_521,N_64);
nor U4061 (N_4061,N_1440,N_97);
nor U4062 (N_4062,N_1443,N_1604);
xnor U4063 (N_4063,N_2067,N_1281);
nor U4064 (N_4064,N_817,N_2392);
nand U4065 (N_4065,N_285,N_1224);
nand U4066 (N_4066,N_1204,N_1097);
nand U4067 (N_4067,N_1634,N_925);
nor U4068 (N_4068,N_1607,N_1107);
and U4069 (N_4069,N_1223,N_1923);
nand U4070 (N_4070,N_520,N_961);
nand U4071 (N_4071,N_29,N_769);
and U4072 (N_4072,N_622,N_759);
xor U4073 (N_4073,N_1732,N_1475);
nor U4074 (N_4074,N_1557,N_1234);
nor U4075 (N_4075,N_744,N_1442);
nand U4076 (N_4076,N_1308,N_625);
and U4077 (N_4077,N_1784,N_2132);
xor U4078 (N_4078,N_134,N_2432);
or U4079 (N_4079,N_209,N_1589);
or U4080 (N_4080,N_1557,N_1110);
and U4081 (N_4081,N_2047,N_2420);
nor U4082 (N_4082,N_594,N_2165);
nand U4083 (N_4083,N_399,N_525);
and U4084 (N_4084,N_326,N_926);
xnor U4085 (N_4085,N_450,N_1231);
nor U4086 (N_4086,N_2377,N_1607);
nand U4087 (N_4087,N_492,N_1472);
or U4088 (N_4088,N_1364,N_859);
and U4089 (N_4089,N_2433,N_17);
and U4090 (N_4090,N_1482,N_1882);
nor U4091 (N_4091,N_1072,N_696);
xor U4092 (N_4092,N_710,N_1884);
or U4093 (N_4093,N_380,N_1493);
xnor U4094 (N_4094,N_1433,N_995);
and U4095 (N_4095,N_2284,N_276);
xor U4096 (N_4096,N_1112,N_814);
or U4097 (N_4097,N_1285,N_1095);
nand U4098 (N_4098,N_903,N_416);
xor U4099 (N_4099,N_45,N_1610);
nand U4100 (N_4100,N_1804,N_1625);
and U4101 (N_4101,N_1685,N_197);
and U4102 (N_4102,N_1418,N_660);
or U4103 (N_4103,N_2162,N_825);
and U4104 (N_4104,N_816,N_1029);
xor U4105 (N_4105,N_234,N_1798);
and U4106 (N_4106,N_100,N_2151);
nor U4107 (N_4107,N_1142,N_91);
xnor U4108 (N_4108,N_2488,N_1661);
or U4109 (N_4109,N_1115,N_1447);
nor U4110 (N_4110,N_2254,N_2020);
or U4111 (N_4111,N_881,N_677);
and U4112 (N_4112,N_1878,N_137);
nand U4113 (N_4113,N_1969,N_48);
nand U4114 (N_4114,N_242,N_2228);
and U4115 (N_4115,N_790,N_2264);
nor U4116 (N_4116,N_1448,N_1592);
xor U4117 (N_4117,N_257,N_547);
nor U4118 (N_4118,N_946,N_1783);
nand U4119 (N_4119,N_1363,N_216);
and U4120 (N_4120,N_2301,N_837);
or U4121 (N_4121,N_1647,N_2048);
nand U4122 (N_4122,N_1925,N_522);
xor U4123 (N_4123,N_1855,N_472);
nand U4124 (N_4124,N_350,N_93);
and U4125 (N_4125,N_2442,N_893);
nor U4126 (N_4126,N_581,N_1362);
or U4127 (N_4127,N_996,N_1267);
nand U4128 (N_4128,N_124,N_1903);
nand U4129 (N_4129,N_1716,N_1790);
and U4130 (N_4130,N_1944,N_922);
xor U4131 (N_4131,N_1227,N_1877);
and U4132 (N_4132,N_1503,N_1738);
nor U4133 (N_4133,N_1034,N_142);
nor U4134 (N_4134,N_1439,N_2424);
xor U4135 (N_4135,N_1443,N_2187);
xor U4136 (N_4136,N_1264,N_1623);
nand U4137 (N_4137,N_489,N_1202);
or U4138 (N_4138,N_717,N_2345);
nor U4139 (N_4139,N_167,N_1237);
xnor U4140 (N_4140,N_1794,N_2047);
and U4141 (N_4141,N_739,N_2442);
and U4142 (N_4142,N_2039,N_1996);
xnor U4143 (N_4143,N_691,N_1284);
xor U4144 (N_4144,N_2286,N_45);
and U4145 (N_4145,N_466,N_217);
or U4146 (N_4146,N_2398,N_2015);
xor U4147 (N_4147,N_235,N_1757);
xnor U4148 (N_4148,N_1868,N_2002);
xor U4149 (N_4149,N_9,N_1148);
nand U4150 (N_4150,N_1031,N_1300);
and U4151 (N_4151,N_2393,N_1960);
nor U4152 (N_4152,N_707,N_702);
nand U4153 (N_4153,N_702,N_1594);
nand U4154 (N_4154,N_2442,N_1007);
nand U4155 (N_4155,N_202,N_1454);
xor U4156 (N_4156,N_2495,N_620);
nand U4157 (N_4157,N_354,N_580);
nor U4158 (N_4158,N_1838,N_2451);
nand U4159 (N_4159,N_2304,N_1022);
and U4160 (N_4160,N_1492,N_1251);
or U4161 (N_4161,N_1656,N_1991);
or U4162 (N_4162,N_1029,N_1877);
xnor U4163 (N_4163,N_1867,N_471);
nand U4164 (N_4164,N_2066,N_12);
nor U4165 (N_4165,N_570,N_2272);
or U4166 (N_4166,N_740,N_185);
nor U4167 (N_4167,N_1047,N_111);
xnor U4168 (N_4168,N_1889,N_444);
and U4169 (N_4169,N_293,N_1636);
or U4170 (N_4170,N_421,N_1053);
nand U4171 (N_4171,N_408,N_1639);
nor U4172 (N_4172,N_481,N_380);
nor U4173 (N_4173,N_1629,N_998);
nor U4174 (N_4174,N_2018,N_2435);
xnor U4175 (N_4175,N_1827,N_106);
or U4176 (N_4176,N_1123,N_633);
nor U4177 (N_4177,N_595,N_1976);
nand U4178 (N_4178,N_2363,N_693);
or U4179 (N_4179,N_2256,N_972);
and U4180 (N_4180,N_1809,N_2472);
or U4181 (N_4181,N_1531,N_281);
and U4182 (N_4182,N_295,N_213);
and U4183 (N_4183,N_2183,N_752);
or U4184 (N_4184,N_1268,N_2313);
xor U4185 (N_4185,N_180,N_1157);
nand U4186 (N_4186,N_434,N_352);
xnor U4187 (N_4187,N_2117,N_535);
nand U4188 (N_4188,N_2274,N_1490);
or U4189 (N_4189,N_927,N_1164);
xnor U4190 (N_4190,N_558,N_1166);
nor U4191 (N_4191,N_1905,N_231);
or U4192 (N_4192,N_701,N_422);
or U4193 (N_4193,N_2069,N_2090);
nand U4194 (N_4194,N_787,N_1975);
nor U4195 (N_4195,N_549,N_1064);
or U4196 (N_4196,N_1210,N_581);
xnor U4197 (N_4197,N_1828,N_630);
xor U4198 (N_4198,N_2269,N_20);
nor U4199 (N_4199,N_1703,N_892);
or U4200 (N_4200,N_1087,N_2275);
nand U4201 (N_4201,N_280,N_2476);
nor U4202 (N_4202,N_1146,N_1052);
and U4203 (N_4203,N_267,N_62);
or U4204 (N_4204,N_1311,N_1596);
nor U4205 (N_4205,N_1524,N_93);
xnor U4206 (N_4206,N_1083,N_1571);
and U4207 (N_4207,N_1099,N_2457);
nor U4208 (N_4208,N_1117,N_856);
nand U4209 (N_4209,N_549,N_1272);
xnor U4210 (N_4210,N_2301,N_755);
nor U4211 (N_4211,N_423,N_2215);
nor U4212 (N_4212,N_1122,N_2135);
nor U4213 (N_4213,N_271,N_1819);
nor U4214 (N_4214,N_2096,N_1198);
or U4215 (N_4215,N_1813,N_1468);
xor U4216 (N_4216,N_1442,N_749);
nand U4217 (N_4217,N_1061,N_2044);
nand U4218 (N_4218,N_2115,N_2428);
nand U4219 (N_4219,N_616,N_2338);
nor U4220 (N_4220,N_1153,N_1266);
nor U4221 (N_4221,N_1373,N_948);
nor U4222 (N_4222,N_1427,N_1980);
and U4223 (N_4223,N_2461,N_660);
nor U4224 (N_4224,N_1803,N_1852);
and U4225 (N_4225,N_287,N_1897);
nor U4226 (N_4226,N_998,N_2057);
and U4227 (N_4227,N_1279,N_705);
xnor U4228 (N_4228,N_1693,N_1972);
nor U4229 (N_4229,N_467,N_199);
xnor U4230 (N_4230,N_837,N_2245);
and U4231 (N_4231,N_2232,N_870);
and U4232 (N_4232,N_1148,N_1155);
xnor U4233 (N_4233,N_2434,N_1369);
xnor U4234 (N_4234,N_646,N_2224);
xor U4235 (N_4235,N_1484,N_1116);
nand U4236 (N_4236,N_1213,N_1644);
nand U4237 (N_4237,N_2345,N_1000);
nand U4238 (N_4238,N_947,N_2120);
xnor U4239 (N_4239,N_950,N_1286);
nor U4240 (N_4240,N_108,N_1060);
nand U4241 (N_4241,N_1158,N_1741);
or U4242 (N_4242,N_2387,N_780);
or U4243 (N_4243,N_1754,N_1143);
and U4244 (N_4244,N_1595,N_1135);
and U4245 (N_4245,N_1252,N_1541);
or U4246 (N_4246,N_82,N_845);
and U4247 (N_4247,N_572,N_152);
or U4248 (N_4248,N_1479,N_1546);
or U4249 (N_4249,N_741,N_1589);
xor U4250 (N_4250,N_603,N_1669);
and U4251 (N_4251,N_579,N_1886);
nand U4252 (N_4252,N_2279,N_916);
xor U4253 (N_4253,N_574,N_1785);
nor U4254 (N_4254,N_2223,N_2393);
and U4255 (N_4255,N_2236,N_1897);
or U4256 (N_4256,N_1183,N_1066);
nand U4257 (N_4257,N_1569,N_710);
and U4258 (N_4258,N_44,N_872);
and U4259 (N_4259,N_2074,N_752);
nand U4260 (N_4260,N_2230,N_1505);
or U4261 (N_4261,N_847,N_879);
nand U4262 (N_4262,N_676,N_1311);
nor U4263 (N_4263,N_923,N_1331);
and U4264 (N_4264,N_2161,N_1876);
nor U4265 (N_4265,N_797,N_2433);
xnor U4266 (N_4266,N_2267,N_199);
and U4267 (N_4267,N_990,N_1287);
nand U4268 (N_4268,N_407,N_1967);
and U4269 (N_4269,N_1185,N_199);
or U4270 (N_4270,N_1034,N_568);
xnor U4271 (N_4271,N_1579,N_1093);
nand U4272 (N_4272,N_2418,N_2365);
nand U4273 (N_4273,N_1413,N_1097);
and U4274 (N_4274,N_750,N_613);
or U4275 (N_4275,N_941,N_1966);
or U4276 (N_4276,N_1945,N_1872);
or U4277 (N_4277,N_183,N_214);
xnor U4278 (N_4278,N_2460,N_666);
or U4279 (N_4279,N_519,N_1176);
nor U4280 (N_4280,N_2494,N_2270);
nand U4281 (N_4281,N_228,N_605);
xnor U4282 (N_4282,N_562,N_1011);
nand U4283 (N_4283,N_810,N_880);
xor U4284 (N_4284,N_2219,N_1915);
or U4285 (N_4285,N_618,N_281);
xor U4286 (N_4286,N_1714,N_2479);
nor U4287 (N_4287,N_1966,N_23);
and U4288 (N_4288,N_2205,N_893);
or U4289 (N_4289,N_2021,N_1278);
nand U4290 (N_4290,N_125,N_545);
and U4291 (N_4291,N_2377,N_1061);
nor U4292 (N_4292,N_1596,N_1675);
nor U4293 (N_4293,N_1076,N_2492);
and U4294 (N_4294,N_786,N_1220);
xor U4295 (N_4295,N_1455,N_230);
and U4296 (N_4296,N_736,N_1714);
or U4297 (N_4297,N_2392,N_112);
and U4298 (N_4298,N_768,N_1349);
and U4299 (N_4299,N_1163,N_796);
xnor U4300 (N_4300,N_1645,N_204);
or U4301 (N_4301,N_1298,N_1407);
nand U4302 (N_4302,N_891,N_985);
and U4303 (N_4303,N_854,N_1787);
xnor U4304 (N_4304,N_2088,N_2034);
nor U4305 (N_4305,N_308,N_2094);
and U4306 (N_4306,N_1410,N_129);
nor U4307 (N_4307,N_1274,N_2158);
xor U4308 (N_4308,N_931,N_1365);
and U4309 (N_4309,N_2190,N_1764);
nor U4310 (N_4310,N_1235,N_2395);
and U4311 (N_4311,N_1628,N_110);
and U4312 (N_4312,N_323,N_1543);
or U4313 (N_4313,N_1981,N_1169);
or U4314 (N_4314,N_653,N_308);
nand U4315 (N_4315,N_1553,N_365);
nor U4316 (N_4316,N_917,N_1456);
or U4317 (N_4317,N_1879,N_1989);
and U4318 (N_4318,N_190,N_2348);
or U4319 (N_4319,N_854,N_550);
and U4320 (N_4320,N_2293,N_1537);
nor U4321 (N_4321,N_1508,N_1833);
nand U4322 (N_4322,N_1342,N_1368);
nand U4323 (N_4323,N_680,N_279);
and U4324 (N_4324,N_919,N_549);
or U4325 (N_4325,N_956,N_1629);
nor U4326 (N_4326,N_2121,N_825);
nor U4327 (N_4327,N_1671,N_876);
and U4328 (N_4328,N_2019,N_802);
nor U4329 (N_4329,N_1662,N_609);
and U4330 (N_4330,N_37,N_862);
and U4331 (N_4331,N_2199,N_1586);
xnor U4332 (N_4332,N_972,N_888);
xnor U4333 (N_4333,N_344,N_635);
nor U4334 (N_4334,N_155,N_701);
xor U4335 (N_4335,N_826,N_2132);
nand U4336 (N_4336,N_273,N_264);
and U4337 (N_4337,N_2073,N_2385);
or U4338 (N_4338,N_600,N_1692);
xor U4339 (N_4339,N_1640,N_807);
and U4340 (N_4340,N_1849,N_2298);
nor U4341 (N_4341,N_1811,N_398);
nand U4342 (N_4342,N_1039,N_384);
nand U4343 (N_4343,N_904,N_1295);
or U4344 (N_4344,N_1408,N_2464);
or U4345 (N_4345,N_918,N_346);
nand U4346 (N_4346,N_2407,N_1603);
nor U4347 (N_4347,N_369,N_2101);
and U4348 (N_4348,N_290,N_2047);
and U4349 (N_4349,N_1571,N_2130);
and U4350 (N_4350,N_872,N_1568);
nand U4351 (N_4351,N_2215,N_397);
and U4352 (N_4352,N_2106,N_524);
or U4353 (N_4353,N_2357,N_1376);
xnor U4354 (N_4354,N_1328,N_129);
nor U4355 (N_4355,N_353,N_1595);
nor U4356 (N_4356,N_267,N_1437);
and U4357 (N_4357,N_547,N_2045);
nand U4358 (N_4358,N_1676,N_872);
xnor U4359 (N_4359,N_2334,N_739);
nor U4360 (N_4360,N_1683,N_371);
nor U4361 (N_4361,N_1984,N_937);
and U4362 (N_4362,N_1229,N_1209);
and U4363 (N_4363,N_2313,N_2384);
and U4364 (N_4364,N_500,N_1847);
or U4365 (N_4365,N_1569,N_1974);
or U4366 (N_4366,N_2494,N_1401);
and U4367 (N_4367,N_2139,N_2328);
nor U4368 (N_4368,N_1059,N_1979);
nor U4369 (N_4369,N_2200,N_125);
xor U4370 (N_4370,N_45,N_304);
and U4371 (N_4371,N_251,N_362);
nor U4372 (N_4372,N_326,N_425);
and U4373 (N_4373,N_934,N_2011);
or U4374 (N_4374,N_2121,N_1588);
or U4375 (N_4375,N_2317,N_476);
nand U4376 (N_4376,N_521,N_1491);
and U4377 (N_4377,N_2090,N_1227);
xor U4378 (N_4378,N_1047,N_887);
and U4379 (N_4379,N_1204,N_2051);
xor U4380 (N_4380,N_1119,N_2235);
or U4381 (N_4381,N_2339,N_1443);
and U4382 (N_4382,N_2,N_1436);
nand U4383 (N_4383,N_1987,N_1100);
or U4384 (N_4384,N_1523,N_567);
or U4385 (N_4385,N_1868,N_348);
and U4386 (N_4386,N_322,N_1467);
xor U4387 (N_4387,N_833,N_1539);
or U4388 (N_4388,N_1296,N_1214);
nor U4389 (N_4389,N_902,N_823);
nand U4390 (N_4390,N_1980,N_613);
xor U4391 (N_4391,N_1717,N_1462);
xor U4392 (N_4392,N_1087,N_1913);
or U4393 (N_4393,N_573,N_1048);
nor U4394 (N_4394,N_479,N_915);
and U4395 (N_4395,N_909,N_1932);
and U4396 (N_4396,N_117,N_2443);
nor U4397 (N_4397,N_707,N_1142);
xnor U4398 (N_4398,N_2309,N_1853);
nand U4399 (N_4399,N_71,N_489);
xnor U4400 (N_4400,N_2107,N_790);
nor U4401 (N_4401,N_2098,N_1831);
and U4402 (N_4402,N_1228,N_2067);
nand U4403 (N_4403,N_963,N_1135);
nand U4404 (N_4404,N_2297,N_1015);
nand U4405 (N_4405,N_928,N_1041);
xnor U4406 (N_4406,N_1347,N_820);
and U4407 (N_4407,N_1179,N_2);
xor U4408 (N_4408,N_216,N_362);
and U4409 (N_4409,N_2482,N_1943);
xnor U4410 (N_4410,N_2217,N_28);
xnor U4411 (N_4411,N_2068,N_288);
and U4412 (N_4412,N_1896,N_2000);
nand U4413 (N_4413,N_833,N_129);
xnor U4414 (N_4414,N_2403,N_2408);
and U4415 (N_4415,N_1781,N_2011);
nand U4416 (N_4416,N_623,N_465);
or U4417 (N_4417,N_2067,N_293);
xnor U4418 (N_4418,N_1584,N_2046);
nor U4419 (N_4419,N_919,N_322);
nor U4420 (N_4420,N_1297,N_503);
or U4421 (N_4421,N_1119,N_2301);
nor U4422 (N_4422,N_2439,N_402);
and U4423 (N_4423,N_2083,N_1983);
and U4424 (N_4424,N_2494,N_1093);
nor U4425 (N_4425,N_278,N_653);
and U4426 (N_4426,N_467,N_450);
nor U4427 (N_4427,N_2166,N_697);
and U4428 (N_4428,N_2128,N_44);
and U4429 (N_4429,N_652,N_57);
xnor U4430 (N_4430,N_757,N_1149);
and U4431 (N_4431,N_117,N_773);
xnor U4432 (N_4432,N_2311,N_1604);
or U4433 (N_4433,N_1265,N_331);
or U4434 (N_4434,N_526,N_791);
nand U4435 (N_4435,N_21,N_174);
and U4436 (N_4436,N_2012,N_1349);
and U4437 (N_4437,N_1065,N_2160);
or U4438 (N_4438,N_1864,N_2);
and U4439 (N_4439,N_2443,N_2485);
xor U4440 (N_4440,N_443,N_1328);
nor U4441 (N_4441,N_2302,N_2379);
and U4442 (N_4442,N_1021,N_2088);
or U4443 (N_4443,N_1358,N_439);
xnor U4444 (N_4444,N_1384,N_1593);
and U4445 (N_4445,N_2030,N_1118);
xnor U4446 (N_4446,N_361,N_771);
or U4447 (N_4447,N_1356,N_254);
or U4448 (N_4448,N_1983,N_1215);
xnor U4449 (N_4449,N_512,N_2013);
and U4450 (N_4450,N_1848,N_1308);
and U4451 (N_4451,N_2303,N_717);
xor U4452 (N_4452,N_1356,N_266);
nand U4453 (N_4453,N_2323,N_1830);
nand U4454 (N_4454,N_1353,N_175);
or U4455 (N_4455,N_355,N_1985);
nor U4456 (N_4456,N_540,N_2141);
nand U4457 (N_4457,N_2193,N_1939);
or U4458 (N_4458,N_384,N_1563);
xor U4459 (N_4459,N_709,N_412);
xor U4460 (N_4460,N_711,N_1834);
xor U4461 (N_4461,N_98,N_1145);
or U4462 (N_4462,N_1479,N_2483);
nor U4463 (N_4463,N_1501,N_1221);
nor U4464 (N_4464,N_1654,N_639);
or U4465 (N_4465,N_2070,N_2161);
nor U4466 (N_4466,N_637,N_1531);
or U4467 (N_4467,N_2179,N_133);
nor U4468 (N_4468,N_1098,N_113);
nor U4469 (N_4469,N_1202,N_877);
or U4470 (N_4470,N_789,N_2333);
nor U4471 (N_4471,N_2438,N_50);
xor U4472 (N_4472,N_81,N_2261);
or U4473 (N_4473,N_1472,N_2320);
xnor U4474 (N_4474,N_671,N_1462);
nand U4475 (N_4475,N_1063,N_172);
and U4476 (N_4476,N_670,N_1612);
and U4477 (N_4477,N_1087,N_354);
nor U4478 (N_4478,N_1922,N_962);
nand U4479 (N_4479,N_1664,N_1267);
nand U4480 (N_4480,N_39,N_2050);
nand U4481 (N_4481,N_1925,N_1366);
and U4482 (N_4482,N_1393,N_120);
xor U4483 (N_4483,N_285,N_903);
nand U4484 (N_4484,N_941,N_1673);
nor U4485 (N_4485,N_1917,N_2486);
or U4486 (N_4486,N_2235,N_281);
or U4487 (N_4487,N_104,N_2481);
or U4488 (N_4488,N_2497,N_2293);
nand U4489 (N_4489,N_1705,N_806);
nor U4490 (N_4490,N_867,N_1119);
and U4491 (N_4491,N_2175,N_2020);
xnor U4492 (N_4492,N_113,N_936);
xor U4493 (N_4493,N_98,N_465);
nor U4494 (N_4494,N_845,N_833);
nand U4495 (N_4495,N_817,N_508);
nor U4496 (N_4496,N_799,N_1032);
or U4497 (N_4497,N_641,N_1137);
nand U4498 (N_4498,N_989,N_1551);
xnor U4499 (N_4499,N_1802,N_1167);
and U4500 (N_4500,N_1636,N_1587);
nor U4501 (N_4501,N_2103,N_174);
or U4502 (N_4502,N_2199,N_1072);
xor U4503 (N_4503,N_879,N_2252);
and U4504 (N_4504,N_1678,N_1563);
xor U4505 (N_4505,N_153,N_1150);
and U4506 (N_4506,N_2447,N_340);
nand U4507 (N_4507,N_1723,N_837);
nor U4508 (N_4508,N_1334,N_78);
xnor U4509 (N_4509,N_902,N_660);
or U4510 (N_4510,N_45,N_1990);
nor U4511 (N_4511,N_1950,N_2114);
or U4512 (N_4512,N_1244,N_784);
and U4513 (N_4513,N_742,N_1150);
and U4514 (N_4514,N_792,N_1840);
or U4515 (N_4515,N_162,N_588);
xor U4516 (N_4516,N_2165,N_1006);
and U4517 (N_4517,N_1312,N_198);
or U4518 (N_4518,N_389,N_1959);
and U4519 (N_4519,N_1509,N_674);
xnor U4520 (N_4520,N_2423,N_310);
or U4521 (N_4521,N_310,N_29);
xnor U4522 (N_4522,N_2112,N_570);
xnor U4523 (N_4523,N_1099,N_526);
xor U4524 (N_4524,N_702,N_2277);
or U4525 (N_4525,N_2214,N_1115);
and U4526 (N_4526,N_1878,N_511);
and U4527 (N_4527,N_482,N_1133);
nor U4528 (N_4528,N_147,N_1563);
nor U4529 (N_4529,N_2247,N_1652);
nor U4530 (N_4530,N_252,N_1443);
or U4531 (N_4531,N_2391,N_1047);
xor U4532 (N_4532,N_2386,N_2015);
and U4533 (N_4533,N_183,N_1020);
or U4534 (N_4534,N_2288,N_493);
or U4535 (N_4535,N_131,N_738);
nand U4536 (N_4536,N_662,N_2185);
nor U4537 (N_4537,N_2068,N_1221);
or U4538 (N_4538,N_950,N_918);
and U4539 (N_4539,N_368,N_1412);
nor U4540 (N_4540,N_603,N_175);
and U4541 (N_4541,N_760,N_2041);
or U4542 (N_4542,N_62,N_1451);
nor U4543 (N_4543,N_2364,N_60);
xnor U4544 (N_4544,N_1309,N_435);
xnor U4545 (N_4545,N_1011,N_377);
nand U4546 (N_4546,N_1931,N_1500);
nor U4547 (N_4547,N_1963,N_83);
nor U4548 (N_4548,N_2149,N_1017);
xor U4549 (N_4549,N_2329,N_2309);
nand U4550 (N_4550,N_1847,N_1970);
nand U4551 (N_4551,N_1800,N_2097);
and U4552 (N_4552,N_1257,N_1021);
xor U4553 (N_4553,N_1736,N_1900);
and U4554 (N_4554,N_1359,N_2271);
xor U4555 (N_4555,N_1377,N_1946);
and U4556 (N_4556,N_1501,N_2160);
nor U4557 (N_4557,N_2312,N_2032);
or U4558 (N_4558,N_142,N_528);
and U4559 (N_4559,N_1013,N_344);
or U4560 (N_4560,N_2411,N_1592);
or U4561 (N_4561,N_1386,N_2415);
xor U4562 (N_4562,N_1023,N_1056);
nand U4563 (N_4563,N_406,N_2178);
nand U4564 (N_4564,N_209,N_705);
nor U4565 (N_4565,N_1520,N_349);
xnor U4566 (N_4566,N_2448,N_1848);
nor U4567 (N_4567,N_2064,N_2216);
nor U4568 (N_4568,N_2080,N_1721);
nand U4569 (N_4569,N_253,N_1389);
or U4570 (N_4570,N_1619,N_920);
and U4571 (N_4571,N_367,N_1890);
xnor U4572 (N_4572,N_1278,N_2056);
nand U4573 (N_4573,N_1112,N_1459);
and U4574 (N_4574,N_1035,N_969);
nand U4575 (N_4575,N_234,N_549);
xnor U4576 (N_4576,N_1994,N_1666);
or U4577 (N_4577,N_522,N_2441);
nand U4578 (N_4578,N_605,N_1606);
nand U4579 (N_4579,N_393,N_221);
and U4580 (N_4580,N_315,N_1387);
nor U4581 (N_4581,N_270,N_931);
nor U4582 (N_4582,N_1847,N_152);
nor U4583 (N_4583,N_1024,N_1376);
or U4584 (N_4584,N_466,N_892);
nand U4585 (N_4585,N_1020,N_194);
nand U4586 (N_4586,N_1353,N_1630);
or U4587 (N_4587,N_216,N_1795);
or U4588 (N_4588,N_749,N_2051);
xnor U4589 (N_4589,N_698,N_397);
and U4590 (N_4590,N_1901,N_1598);
and U4591 (N_4591,N_1407,N_1554);
nand U4592 (N_4592,N_1097,N_827);
nand U4593 (N_4593,N_697,N_2016);
nand U4594 (N_4594,N_1179,N_320);
or U4595 (N_4595,N_2118,N_311);
xor U4596 (N_4596,N_37,N_833);
xor U4597 (N_4597,N_1614,N_1898);
and U4598 (N_4598,N_2043,N_1133);
xnor U4599 (N_4599,N_1088,N_1579);
or U4600 (N_4600,N_1556,N_613);
or U4601 (N_4601,N_352,N_228);
xnor U4602 (N_4602,N_157,N_2094);
or U4603 (N_4603,N_776,N_722);
nand U4604 (N_4604,N_2056,N_1111);
nor U4605 (N_4605,N_1851,N_363);
xnor U4606 (N_4606,N_55,N_1420);
or U4607 (N_4607,N_2453,N_1081);
or U4608 (N_4608,N_766,N_842);
or U4609 (N_4609,N_469,N_2164);
and U4610 (N_4610,N_456,N_663);
nand U4611 (N_4611,N_1539,N_860);
xnor U4612 (N_4612,N_2141,N_1910);
or U4613 (N_4613,N_1646,N_55);
nand U4614 (N_4614,N_1068,N_813);
or U4615 (N_4615,N_1250,N_579);
nand U4616 (N_4616,N_2333,N_536);
nand U4617 (N_4617,N_1098,N_272);
and U4618 (N_4618,N_2419,N_382);
or U4619 (N_4619,N_322,N_99);
nor U4620 (N_4620,N_1547,N_1437);
and U4621 (N_4621,N_2427,N_973);
nor U4622 (N_4622,N_1702,N_796);
and U4623 (N_4623,N_740,N_1694);
and U4624 (N_4624,N_1543,N_2263);
nor U4625 (N_4625,N_1477,N_1482);
nand U4626 (N_4626,N_1317,N_486);
nor U4627 (N_4627,N_792,N_789);
nand U4628 (N_4628,N_2367,N_1160);
xor U4629 (N_4629,N_2204,N_1107);
and U4630 (N_4630,N_550,N_1252);
xor U4631 (N_4631,N_1257,N_1531);
xor U4632 (N_4632,N_2003,N_1830);
or U4633 (N_4633,N_591,N_960);
xor U4634 (N_4634,N_1540,N_512);
nor U4635 (N_4635,N_233,N_309);
and U4636 (N_4636,N_1563,N_913);
xnor U4637 (N_4637,N_347,N_946);
nor U4638 (N_4638,N_2005,N_1323);
xnor U4639 (N_4639,N_1435,N_1575);
and U4640 (N_4640,N_628,N_1797);
nand U4641 (N_4641,N_719,N_186);
nand U4642 (N_4642,N_1063,N_193);
and U4643 (N_4643,N_1009,N_264);
and U4644 (N_4644,N_1427,N_1890);
or U4645 (N_4645,N_2214,N_1944);
or U4646 (N_4646,N_1971,N_1861);
nor U4647 (N_4647,N_1838,N_1457);
nand U4648 (N_4648,N_1287,N_2247);
or U4649 (N_4649,N_2069,N_1556);
xnor U4650 (N_4650,N_716,N_2013);
xnor U4651 (N_4651,N_697,N_1434);
and U4652 (N_4652,N_60,N_1819);
and U4653 (N_4653,N_2391,N_461);
or U4654 (N_4654,N_561,N_1494);
and U4655 (N_4655,N_2331,N_588);
and U4656 (N_4656,N_782,N_1354);
nor U4657 (N_4657,N_171,N_1825);
nand U4658 (N_4658,N_1826,N_1703);
nor U4659 (N_4659,N_2092,N_390);
nand U4660 (N_4660,N_817,N_1264);
xnor U4661 (N_4661,N_1225,N_1679);
nor U4662 (N_4662,N_780,N_2247);
xnor U4663 (N_4663,N_2352,N_1194);
or U4664 (N_4664,N_346,N_554);
or U4665 (N_4665,N_961,N_2336);
nand U4666 (N_4666,N_1206,N_1244);
or U4667 (N_4667,N_2167,N_2490);
nand U4668 (N_4668,N_562,N_1540);
and U4669 (N_4669,N_2395,N_659);
or U4670 (N_4670,N_459,N_618);
or U4671 (N_4671,N_2358,N_1078);
nor U4672 (N_4672,N_1451,N_17);
or U4673 (N_4673,N_501,N_2248);
nor U4674 (N_4674,N_2435,N_1022);
and U4675 (N_4675,N_1691,N_1368);
xor U4676 (N_4676,N_2378,N_98);
and U4677 (N_4677,N_2133,N_2186);
and U4678 (N_4678,N_2278,N_712);
nor U4679 (N_4679,N_2166,N_976);
xnor U4680 (N_4680,N_1232,N_1579);
xor U4681 (N_4681,N_1702,N_2431);
xor U4682 (N_4682,N_417,N_624);
nor U4683 (N_4683,N_1849,N_153);
nand U4684 (N_4684,N_595,N_1418);
nor U4685 (N_4685,N_1274,N_459);
and U4686 (N_4686,N_2178,N_13);
xor U4687 (N_4687,N_1944,N_1337);
nand U4688 (N_4688,N_1698,N_576);
xor U4689 (N_4689,N_94,N_2338);
and U4690 (N_4690,N_2021,N_586);
xnor U4691 (N_4691,N_1472,N_499);
or U4692 (N_4692,N_1025,N_802);
xnor U4693 (N_4693,N_770,N_170);
or U4694 (N_4694,N_1683,N_1388);
xnor U4695 (N_4695,N_2347,N_2112);
and U4696 (N_4696,N_2040,N_1155);
xnor U4697 (N_4697,N_60,N_1628);
nand U4698 (N_4698,N_417,N_1788);
xnor U4699 (N_4699,N_2418,N_65);
nand U4700 (N_4700,N_325,N_1073);
xnor U4701 (N_4701,N_362,N_519);
xnor U4702 (N_4702,N_1730,N_1068);
xor U4703 (N_4703,N_1691,N_783);
xnor U4704 (N_4704,N_1168,N_1952);
nor U4705 (N_4705,N_324,N_250);
xnor U4706 (N_4706,N_2473,N_315);
nor U4707 (N_4707,N_1023,N_2482);
nand U4708 (N_4708,N_2133,N_1320);
nor U4709 (N_4709,N_218,N_1699);
or U4710 (N_4710,N_1283,N_323);
and U4711 (N_4711,N_1805,N_262);
xnor U4712 (N_4712,N_809,N_2426);
nor U4713 (N_4713,N_1452,N_1409);
nor U4714 (N_4714,N_1096,N_1578);
xnor U4715 (N_4715,N_287,N_466);
xnor U4716 (N_4716,N_423,N_1579);
or U4717 (N_4717,N_1321,N_1507);
and U4718 (N_4718,N_656,N_588);
xor U4719 (N_4719,N_2260,N_2465);
xor U4720 (N_4720,N_172,N_2490);
nor U4721 (N_4721,N_730,N_87);
or U4722 (N_4722,N_1508,N_66);
and U4723 (N_4723,N_1643,N_671);
and U4724 (N_4724,N_1584,N_526);
or U4725 (N_4725,N_1061,N_2180);
nand U4726 (N_4726,N_72,N_1216);
xnor U4727 (N_4727,N_2421,N_2425);
xnor U4728 (N_4728,N_464,N_1742);
xor U4729 (N_4729,N_1467,N_1819);
nor U4730 (N_4730,N_541,N_1891);
and U4731 (N_4731,N_1419,N_1908);
nor U4732 (N_4732,N_1022,N_1799);
nor U4733 (N_4733,N_767,N_2331);
nand U4734 (N_4734,N_2078,N_422);
nor U4735 (N_4735,N_2461,N_1089);
or U4736 (N_4736,N_2201,N_1103);
nor U4737 (N_4737,N_1501,N_2331);
nand U4738 (N_4738,N_1149,N_458);
nand U4739 (N_4739,N_263,N_226);
or U4740 (N_4740,N_789,N_868);
nor U4741 (N_4741,N_1300,N_333);
xnor U4742 (N_4742,N_177,N_1096);
nor U4743 (N_4743,N_140,N_866);
xnor U4744 (N_4744,N_760,N_1659);
or U4745 (N_4745,N_196,N_1813);
or U4746 (N_4746,N_2006,N_2064);
or U4747 (N_4747,N_675,N_1459);
nand U4748 (N_4748,N_991,N_1735);
or U4749 (N_4749,N_657,N_299);
nor U4750 (N_4750,N_1587,N_1326);
xnor U4751 (N_4751,N_1973,N_2175);
nor U4752 (N_4752,N_1478,N_711);
and U4753 (N_4753,N_2161,N_590);
xnor U4754 (N_4754,N_1107,N_1381);
nand U4755 (N_4755,N_2206,N_1262);
and U4756 (N_4756,N_868,N_403);
nand U4757 (N_4757,N_163,N_1135);
or U4758 (N_4758,N_89,N_1966);
xor U4759 (N_4759,N_2005,N_1982);
or U4760 (N_4760,N_653,N_299);
xnor U4761 (N_4761,N_1299,N_1263);
nor U4762 (N_4762,N_13,N_2358);
nand U4763 (N_4763,N_1823,N_1560);
or U4764 (N_4764,N_2170,N_1470);
nor U4765 (N_4765,N_1658,N_1729);
nand U4766 (N_4766,N_2017,N_1960);
and U4767 (N_4767,N_1558,N_471);
nor U4768 (N_4768,N_1530,N_1545);
xnor U4769 (N_4769,N_1811,N_873);
and U4770 (N_4770,N_316,N_451);
nand U4771 (N_4771,N_2438,N_1282);
and U4772 (N_4772,N_2280,N_741);
or U4773 (N_4773,N_792,N_664);
xnor U4774 (N_4774,N_1140,N_610);
or U4775 (N_4775,N_797,N_1819);
and U4776 (N_4776,N_2327,N_0);
xnor U4777 (N_4777,N_1049,N_72);
or U4778 (N_4778,N_1105,N_1111);
xnor U4779 (N_4779,N_415,N_1248);
nand U4780 (N_4780,N_701,N_1147);
or U4781 (N_4781,N_1440,N_1071);
xor U4782 (N_4782,N_1172,N_1040);
xor U4783 (N_4783,N_1391,N_2067);
and U4784 (N_4784,N_1933,N_1722);
nand U4785 (N_4785,N_1445,N_718);
and U4786 (N_4786,N_2364,N_973);
or U4787 (N_4787,N_981,N_1387);
xnor U4788 (N_4788,N_1518,N_239);
nor U4789 (N_4789,N_374,N_73);
xnor U4790 (N_4790,N_272,N_487);
xnor U4791 (N_4791,N_1029,N_312);
or U4792 (N_4792,N_1745,N_309);
nand U4793 (N_4793,N_890,N_2448);
and U4794 (N_4794,N_558,N_666);
xnor U4795 (N_4795,N_51,N_1923);
xnor U4796 (N_4796,N_473,N_2223);
nand U4797 (N_4797,N_1075,N_1);
xor U4798 (N_4798,N_2071,N_1790);
xnor U4799 (N_4799,N_1626,N_840);
or U4800 (N_4800,N_1213,N_1577);
or U4801 (N_4801,N_1122,N_141);
nor U4802 (N_4802,N_1637,N_2014);
xnor U4803 (N_4803,N_255,N_998);
xnor U4804 (N_4804,N_1834,N_673);
nor U4805 (N_4805,N_1184,N_1185);
and U4806 (N_4806,N_1797,N_717);
xnor U4807 (N_4807,N_116,N_80);
xor U4808 (N_4808,N_1022,N_1956);
nor U4809 (N_4809,N_277,N_2059);
nand U4810 (N_4810,N_423,N_876);
nand U4811 (N_4811,N_427,N_536);
nand U4812 (N_4812,N_73,N_469);
xor U4813 (N_4813,N_1993,N_507);
nand U4814 (N_4814,N_527,N_602);
nor U4815 (N_4815,N_1034,N_1294);
and U4816 (N_4816,N_496,N_170);
xnor U4817 (N_4817,N_1276,N_1065);
nor U4818 (N_4818,N_1413,N_1093);
xor U4819 (N_4819,N_1934,N_332);
or U4820 (N_4820,N_2372,N_1826);
and U4821 (N_4821,N_2391,N_1479);
nor U4822 (N_4822,N_243,N_328);
xnor U4823 (N_4823,N_1572,N_1973);
or U4824 (N_4824,N_2290,N_161);
or U4825 (N_4825,N_2240,N_933);
or U4826 (N_4826,N_1374,N_2020);
or U4827 (N_4827,N_2352,N_1316);
nor U4828 (N_4828,N_573,N_6);
and U4829 (N_4829,N_1425,N_943);
nor U4830 (N_4830,N_795,N_439);
or U4831 (N_4831,N_690,N_1789);
and U4832 (N_4832,N_1073,N_721);
xor U4833 (N_4833,N_308,N_79);
and U4834 (N_4834,N_678,N_247);
and U4835 (N_4835,N_962,N_2268);
or U4836 (N_4836,N_1673,N_2055);
nand U4837 (N_4837,N_1107,N_2120);
nor U4838 (N_4838,N_169,N_394);
nor U4839 (N_4839,N_2321,N_1484);
or U4840 (N_4840,N_1184,N_2301);
and U4841 (N_4841,N_2204,N_2424);
nor U4842 (N_4842,N_1261,N_1247);
xor U4843 (N_4843,N_2318,N_1609);
or U4844 (N_4844,N_2181,N_443);
nand U4845 (N_4845,N_766,N_962);
nand U4846 (N_4846,N_695,N_2155);
xor U4847 (N_4847,N_2029,N_91);
xor U4848 (N_4848,N_503,N_1364);
nor U4849 (N_4849,N_1452,N_2318);
nor U4850 (N_4850,N_795,N_633);
xnor U4851 (N_4851,N_1816,N_2291);
xnor U4852 (N_4852,N_2407,N_2266);
nor U4853 (N_4853,N_163,N_89);
nand U4854 (N_4854,N_39,N_378);
nand U4855 (N_4855,N_1578,N_996);
or U4856 (N_4856,N_1306,N_1528);
and U4857 (N_4857,N_2281,N_861);
nor U4858 (N_4858,N_1583,N_2113);
or U4859 (N_4859,N_1107,N_1076);
and U4860 (N_4860,N_179,N_131);
nor U4861 (N_4861,N_1041,N_1914);
and U4862 (N_4862,N_1853,N_2259);
and U4863 (N_4863,N_238,N_2183);
and U4864 (N_4864,N_1933,N_1092);
or U4865 (N_4865,N_111,N_2095);
nor U4866 (N_4866,N_406,N_930);
nor U4867 (N_4867,N_1237,N_1773);
and U4868 (N_4868,N_1065,N_1621);
nand U4869 (N_4869,N_692,N_1626);
nor U4870 (N_4870,N_1994,N_1584);
and U4871 (N_4871,N_1855,N_219);
xnor U4872 (N_4872,N_2235,N_868);
nor U4873 (N_4873,N_381,N_1775);
xor U4874 (N_4874,N_602,N_1747);
nand U4875 (N_4875,N_301,N_1327);
or U4876 (N_4876,N_23,N_368);
nor U4877 (N_4877,N_1626,N_1497);
xnor U4878 (N_4878,N_166,N_1592);
nor U4879 (N_4879,N_848,N_1804);
or U4880 (N_4880,N_1938,N_884);
nor U4881 (N_4881,N_1750,N_1848);
or U4882 (N_4882,N_498,N_559);
nand U4883 (N_4883,N_1923,N_2001);
nand U4884 (N_4884,N_2001,N_809);
xor U4885 (N_4885,N_1258,N_1261);
and U4886 (N_4886,N_859,N_3);
and U4887 (N_4887,N_2072,N_411);
nor U4888 (N_4888,N_534,N_1186);
nor U4889 (N_4889,N_1904,N_2180);
xor U4890 (N_4890,N_1931,N_2272);
and U4891 (N_4891,N_1411,N_446);
and U4892 (N_4892,N_1168,N_1834);
nor U4893 (N_4893,N_973,N_1222);
xor U4894 (N_4894,N_807,N_118);
nand U4895 (N_4895,N_755,N_553);
or U4896 (N_4896,N_1578,N_2130);
and U4897 (N_4897,N_612,N_2088);
nor U4898 (N_4898,N_1933,N_848);
nand U4899 (N_4899,N_1427,N_67);
nor U4900 (N_4900,N_1848,N_1981);
nand U4901 (N_4901,N_2151,N_1699);
xor U4902 (N_4902,N_1456,N_1111);
or U4903 (N_4903,N_1762,N_1329);
or U4904 (N_4904,N_1910,N_459);
or U4905 (N_4905,N_807,N_1296);
nand U4906 (N_4906,N_122,N_2063);
and U4907 (N_4907,N_749,N_1083);
or U4908 (N_4908,N_1154,N_1853);
xor U4909 (N_4909,N_2006,N_2075);
or U4910 (N_4910,N_566,N_1916);
or U4911 (N_4911,N_1663,N_1487);
nor U4912 (N_4912,N_503,N_2434);
and U4913 (N_4913,N_2037,N_2226);
nor U4914 (N_4914,N_2294,N_2123);
or U4915 (N_4915,N_325,N_1557);
xor U4916 (N_4916,N_584,N_527);
nand U4917 (N_4917,N_2057,N_2342);
and U4918 (N_4918,N_2367,N_2266);
xor U4919 (N_4919,N_229,N_225);
or U4920 (N_4920,N_1545,N_1227);
xnor U4921 (N_4921,N_1163,N_769);
nand U4922 (N_4922,N_543,N_1250);
and U4923 (N_4923,N_1446,N_1745);
xor U4924 (N_4924,N_811,N_979);
or U4925 (N_4925,N_969,N_510);
nor U4926 (N_4926,N_2243,N_1055);
and U4927 (N_4927,N_344,N_2396);
or U4928 (N_4928,N_655,N_2449);
and U4929 (N_4929,N_423,N_2035);
nor U4930 (N_4930,N_1497,N_1179);
or U4931 (N_4931,N_1965,N_1719);
or U4932 (N_4932,N_1325,N_1130);
or U4933 (N_4933,N_787,N_588);
or U4934 (N_4934,N_1438,N_958);
nor U4935 (N_4935,N_1469,N_1287);
nor U4936 (N_4936,N_1834,N_1570);
xnor U4937 (N_4937,N_185,N_128);
or U4938 (N_4938,N_1154,N_1279);
nor U4939 (N_4939,N_1560,N_960);
nand U4940 (N_4940,N_2436,N_739);
nor U4941 (N_4941,N_186,N_1178);
or U4942 (N_4942,N_871,N_456);
nor U4943 (N_4943,N_61,N_1577);
xor U4944 (N_4944,N_2145,N_1204);
nor U4945 (N_4945,N_1992,N_875);
nor U4946 (N_4946,N_9,N_986);
nor U4947 (N_4947,N_2315,N_1908);
nor U4948 (N_4948,N_2223,N_935);
nand U4949 (N_4949,N_1790,N_2486);
nand U4950 (N_4950,N_1153,N_486);
or U4951 (N_4951,N_1515,N_1280);
nor U4952 (N_4952,N_1723,N_172);
and U4953 (N_4953,N_866,N_1887);
nand U4954 (N_4954,N_883,N_422);
xnor U4955 (N_4955,N_1473,N_162);
nor U4956 (N_4956,N_2310,N_1900);
nor U4957 (N_4957,N_1146,N_2247);
nand U4958 (N_4958,N_2133,N_24);
xnor U4959 (N_4959,N_1752,N_247);
and U4960 (N_4960,N_660,N_2197);
xor U4961 (N_4961,N_86,N_1746);
xor U4962 (N_4962,N_1461,N_2120);
nor U4963 (N_4963,N_1470,N_1968);
or U4964 (N_4964,N_268,N_405);
nor U4965 (N_4965,N_1351,N_1801);
nand U4966 (N_4966,N_1756,N_1746);
nand U4967 (N_4967,N_18,N_1593);
xor U4968 (N_4968,N_1293,N_2417);
xnor U4969 (N_4969,N_868,N_1433);
xnor U4970 (N_4970,N_1615,N_421);
or U4971 (N_4971,N_1446,N_3);
nand U4972 (N_4972,N_1443,N_1279);
nor U4973 (N_4973,N_856,N_1703);
nand U4974 (N_4974,N_2428,N_783);
nand U4975 (N_4975,N_1003,N_871);
xnor U4976 (N_4976,N_2197,N_481);
xnor U4977 (N_4977,N_1659,N_1505);
nand U4978 (N_4978,N_427,N_308);
and U4979 (N_4979,N_800,N_598);
or U4980 (N_4980,N_2278,N_1111);
nand U4981 (N_4981,N_457,N_1065);
and U4982 (N_4982,N_2316,N_792);
nor U4983 (N_4983,N_2330,N_271);
nor U4984 (N_4984,N_2137,N_25);
xnor U4985 (N_4985,N_1111,N_358);
xor U4986 (N_4986,N_1746,N_1079);
and U4987 (N_4987,N_756,N_2449);
and U4988 (N_4988,N_2202,N_322);
xnor U4989 (N_4989,N_1973,N_1141);
and U4990 (N_4990,N_1331,N_2487);
and U4991 (N_4991,N_396,N_1492);
and U4992 (N_4992,N_2470,N_697);
nand U4993 (N_4993,N_2306,N_1485);
nand U4994 (N_4994,N_1087,N_2237);
nand U4995 (N_4995,N_1799,N_2136);
xor U4996 (N_4996,N_347,N_2353);
xnor U4997 (N_4997,N_1211,N_189);
nand U4998 (N_4998,N_759,N_269);
or U4999 (N_4999,N_1802,N_1680);
nor U5000 (N_5000,N_4950,N_3075);
nand U5001 (N_5001,N_3883,N_4038);
nor U5002 (N_5002,N_3644,N_3704);
nor U5003 (N_5003,N_4887,N_4925);
and U5004 (N_5004,N_4893,N_4010);
nand U5005 (N_5005,N_3487,N_2564);
and U5006 (N_5006,N_2532,N_4911);
and U5007 (N_5007,N_3404,N_2561);
nor U5008 (N_5008,N_3996,N_4294);
and U5009 (N_5009,N_4840,N_4259);
or U5010 (N_5010,N_2654,N_3674);
and U5011 (N_5011,N_4653,N_3223);
or U5012 (N_5012,N_4309,N_4854);
xor U5013 (N_5013,N_2830,N_3057);
nand U5014 (N_5014,N_4136,N_4710);
nand U5015 (N_5015,N_3212,N_3356);
xor U5016 (N_5016,N_4049,N_2596);
or U5017 (N_5017,N_2533,N_2949);
or U5018 (N_5018,N_4677,N_2639);
nor U5019 (N_5019,N_3975,N_4196);
nor U5020 (N_5020,N_4523,N_3537);
and U5021 (N_5021,N_4124,N_4031);
and U5022 (N_5022,N_3894,N_3747);
xor U5023 (N_5023,N_4637,N_4200);
and U5024 (N_5024,N_3655,N_2802);
or U5025 (N_5025,N_2972,N_3401);
nor U5026 (N_5026,N_2528,N_4818);
nor U5027 (N_5027,N_3776,N_2910);
and U5028 (N_5028,N_4402,N_4150);
xnor U5029 (N_5029,N_3698,N_3302);
nor U5030 (N_5030,N_2587,N_2760);
xnor U5031 (N_5031,N_4148,N_4682);
and U5032 (N_5032,N_3750,N_3526);
and U5033 (N_5033,N_3293,N_3406);
xnor U5034 (N_5034,N_2702,N_3167);
or U5035 (N_5035,N_3885,N_2772);
nand U5036 (N_5036,N_4232,N_3717);
and U5037 (N_5037,N_2676,N_3153);
nand U5038 (N_5038,N_2788,N_2745);
or U5039 (N_5039,N_3228,N_2866);
nand U5040 (N_5040,N_3496,N_4057);
nand U5041 (N_5041,N_4363,N_3659);
and U5042 (N_5042,N_3096,N_3927);
or U5043 (N_5043,N_4100,N_4012);
xnor U5044 (N_5044,N_3934,N_4505);
and U5045 (N_5045,N_4183,N_3560);
nor U5046 (N_5046,N_4502,N_3769);
xnor U5047 (N_5047,N_3594,N_3175);
nand U5048 (N_5048,N_2786,N_4310);
nand U5049 (N_5049,N_3267,N_2658);
nand U5050 (N_5050,N_3602,N_4191);
xor U5051 (N_5051,N_4387,N_3363);
nor U5052 (N_5052,N_4915,N_2579);
xor U5053 (N_5053,N_3983,N_3033);
nor U5054 (N_5054,N_4600,N_4696);
xnor U5055 (N_5055,N_4519,N_4476);
xor U5056 (N_5056,N_4233,N_4533);
or U5057 (N_5057,N_4709,N_3499);
or U5058 (N_5058,N_3206,N_4484);
xor U5059 (N_5059,N_3194,N_4611);
or U5060 (N_5060,N_3138,N_4914);
and U5061 (N_5061,N_4969,N_3669);
or U5062 (N_5062,N_4871,N_4921);
nand U5063 (N_5063,N_4406,N_2610);
xor U5064 (N_5064,N_2796,N_4493);
xor U5065 (N_5065,N_3304,N_4960);
nand U5066 (N_5066,N_4019,N_2734);
nor U5067 (N_5067,N_3082,N_2825);
nand U5068 (N_5068,N_2586,N_4572);
and U5069 (N_5069,N_4864,N_2882);
and U5070 (N_5070,N_4377,N_4464);
nor U5071 (N_5071,N_2693,N_3266);
nor U5072 (N_5072,N_4807,N_2959);
xor U5073 (N_5073,N_3347,N_4570);
nand U5074 (N_5074,N_3101,N_3572);
xor U5075 (N_5075,N_4251,N_3190);
nand U5076 (N_5076,N_2895,N_3129);
or U5077 (N_5077,N_3038,N_4959);
and U5078 (N_5078,N_2785,N_3492);
nor U5079 (N_5079,N_4895,N_4253);
or U5080 (N_5080,N_3312,N_3893);
nor U5081 (N_5081,N_3879,N_3549);
and U5082 (N_5082,N_4568,N_3865);
nand U5083 (N_5083,N_3607,N_4023);
and U5084 (N_5084,N_4112,N_3115);
and U5085 (N_5085,N_4993,N_4287);
nor U5086 (N_5086,N_3695,N_3204);
and U5087 (N_5087,N_2956,N_4545);
and U5088 (N_5088,N_3196,N_3543);
and U5089 (N_5089,N_2937,N_3703);
nand U5090 (N_5090,N_2621,N_3755);
nor U5091 (N_5091,N_3683,N_3671);
xor U5092 (N_5092,N_4546,N_2665);
or U5093 (N_5093,N_3413,N_3910);
nand U5094 (N_5094,N_3110,N_4811);
and U5095 (N_5095,N_4945,N_3801);
xnor U5096 (N_5096,N_2606,N_2574);
or U5097 (N_5097,N_3724,N_4229);
xnor U5098 (N_5098,N_3136,N_3843);
nor U5099 (N_5099,N_4783,N_2661);
or U5100 (N_5100,N_3113,N_4353);
nor U5101 (N_5101,N_4099,N_2551);
or U5102 (N_5102,N_2710,N_4935);
and U5103 (N_5103,N_4385,N_3036);
or U5104 (N_5104,N_4633,N_4567);
and U5105 (N_5105,N_3948,N_4342);
and U5106 (N_5106,N_4606,N_3920);
xnor U5107 (N_5107,N_3208,N_2752);
and U5108 (N_5108,N_3043,N_3229);
xor U5109 (N_5109,N_4890,N_4797);
nand U5110 (N_5110,N_2744,N_2504);
or U5111 (N_5111,N_4497,N_2684);
xnor U5112 (N_5112,N_3985,N_3775);
nor U5113 (N_5113,N_4375,N_3062);
and U5114 (N_5114,N_4708,N_2995);
and U5115 (N_5115,N_3818,N_3748);
nor U5116 (N_5116,N_2915,N_3445);
nand U5117 (N_5117,N_3981,N_3546);
xor U5118 (N_5118,N_3249,N_4859);
and U5119 (N_5119,N_3907,N_3783);
nand U5120 (N_5120,N_2713,N_4899);
xor U5121 (N_5121,N_4180,N_4117);
xnor U5122 (N_5122,N_2902,N_2567);
or U5123 (N_5123,N_3020,N_2926);
nor U5124 (N_5124,N_2622,N_3221);
nor U5125 (N_5125,N_3502,N_4341);
or U5126 (N_5126,N_4457,N_2728);
nand U5127 (N_5127,N_2948,N_2555);
nor U5128 (N_5128,N_3681,N_2618);
nor U5129 (N_5129,N_4860,N_4759);
nor U5130 (N_5130,N_3389,N_3651);
nand U5131 (N_5131,N_4129,N_3690);
and U5132 (N_5132,N_2843,N_2717);
nand U5133 (N_5133,N_4306,N_4033);
xnor U5134 (N_5134,N_4780,N_2731);
or U5135 (N_5135,N_2727,N_3398);
and U5136 (N_5136,N_3366,N_3309);
xnor U5137 (N_5137,N_3935,N_4867);
nor U5138 (N_5138,N_3006,N_3387);
nand U5139 (N_5139,N_4737,N_4316);
nor U5140 (N_5140,N_3003,N_3455);
xor U5141 (N_5141,N_3982,N_2633);
and U5142 (N_5142,N_3008,N_4941);
nor U5143 (N_5143,N_4805,N_4615);
and U5144 (N_5144,N_4460,N_4535);
or U5145 (N_5145,N_3552,N_2766);
and U5146 (N_5146,N_2865,N_4270);
or U5147 (N_5147,N_3545,N_4501);
and U5148 (N_5148,N_3353,N_3622);
xnor U5149 (N_5149,N_2932,N_4499);
or U5150 (N_5150,N_4444,N_3611);
nor U5151 (N_5151,N_3710,N_2847);
and U5152 (N_5152,N_2826,N_3479);
and U5153 (N_5153,N_4092,N_2550);
and U5154 (N_5154,N_3226,N_2729);
and U5155 (N_5155,N_2563,N_4734);
nand U5156 (N_5156,N_2794,N_3630);
or U5157 (N_5157,N_4120,N_3434);
or U5158 (N_5158,N_2627,N_2923);
or U5159 (N_5159,N_3000,N_4848);
nand U5160 (N_5160,N_3288,N_3351);
and U5161 (N_5161,N_2664,N_4898);
xor U5162 (N_5162,N_2749,N_4198);
nor U5163 (N_5163,N_2793,N_2867);
nor U5164 (N_5164,N_3271,N_3396);
nand U5165 (N_5165,N_2632,N_3964);
xor U5166 (N_5166,N_3149,N_2589);
xor U5167 (N_5167,N_3343,N_2540);
nand U5168 (N_5168,N_3960,N_3158);
or U5169 (N_5169,N_4826,N_4603);
nor U5170 (N_5170,N_2971,N_4711);
nand U5171 (N_5171,N_3903,N_2650);
xor U5172 (N_5172,N_4052,N_3444);
xor U5173 (N_5173,N_4624,N_2962);
and U5174 (N_5174,N_2900,N_3641);
xnor U5175 (N_5175,N_2645,N_2679);
or U5176 (N_5176,N_3744,N_2705);
xnor U5177 (N_5177,N_4176,N_3958);
and U5178 (N_5178,N_4000,N_3768);
or U5179 (N_5179,N_3119,N_2776);
nand U5180 (N_5180,N_3260,N_2741);
nand U5181 (N_5181,N_3328,N_4951);
nand U5182 (N_5182,N_4770,N_4209);
or U5183 (N_5183,N_3073,N_3160);
xor U5184 (N_5184,N_2598,N_4997);
and U5185 (N_5185,N_4383,N_3415);
xor U5186 (N_5186,N_4220,N_4018);
and U5187 (N_5187,N_4660,N_4961);
and U5188 (N_5188,N_4230,N_4108);
nor U5189 (N_5189,N_4299,N_3796);
nand U5190 (N_5190,N_4326,N_3337);
nand U5191 (N_5191,N_3254,N_4067);
nor U5192 (N_5192,N_4016,N_3074);
and U5193 (N_5193,N_2597,N_4678);
xnor U5194 (N_5194,N_4528,N_4591);
nand U5195 (N_5195,N_3700,N_3259);
xnor U5196 (N_5196,N_3086,N_2570);
nand U5197 (N_5197,N_4784,N_3891);
or U5198 (N_5198,N_2940,N_4034);
or U5199 (N_5199,N_4221,N_3418);
or U5200 (N_5200,N_2725,N_4320);
nor U5201 (N_5201,N_2828,N_4876);
and U5202 (N_5202,N_4081,N_4097);
nor U5203 (N_5203,N_3889,N_4261);
or U5204 (N_5204,N_3264,N_4837);
or U5205 (N_5205,N_2827,N_4947);
and U5206 (N_5206,N_4757,N_4690);
nand U5207 (N_5207,N_3899,N_3077);
nand U5208 (N_5208,N_2569,N_4596);
xor U5209 (N_5209,N_3999,N_4843);
or U5210 (N_5210,N_4995,N_4977);
xor U5211 (N_5211,N_3823,N_2666);
or U5212 (N_5212,N_4459,N_2851);
and U5213 (N_5213,N_3919,N_3477);
nand U5214 (N_5214,N_3466,N_3493);
nand U5215 (N_5215,N_2953,N_3811);
xnor U5216 (N_5216,N_3362,N_2817);
or U5217 (N_5217,N_3658,N_3880);
xor U5218 (N_5218,N_4906,N_3367);
nand U5219 (N_5219,N_4727,N_2980);
nor U5220 (N_5220,N_3794,N_2801);
nand U5221 (N_5221,N_3130,N_3344);
and U5222 (N_5222,N_4702,N_2719);
nor U5223 (N_5223,N_3712,N_4064);
or U5224 (N_5224,N_4247,N_3083);
nor U5225 (N_5225,N_4698,N_3861);
nand U5226 (N_5226,N_4442,N_3956);
and U5227 (N_5227,N_3048,N_3198);
xnor U5228 (N_5228,N_2892,N_2967);
xnor U5229 (N_5229,N_4269,N_3354);
nand U5230 (N_5230,N_3730,N_3318);
nand U5231 (N_5231,N_2888,N_4255);
nor U5232 (N_5232,N_2985,N_2588);
and U5233 (N_5233,N_2536,N_3649);
or U5234 (N_5234,N_3497,N_3189);
and U5235 (N_5235,N_4787,N_3623);
and U5236 (N_5236,N_4823,N_4610);
nand U5237 (N_5237,N_4612,N_2904);
and U5238 (N_5238,N_2916,N_4641);
and U5239 (N_5239,N_3433,N_4589);
and U5240 (N_5240,N_4715,N_2880);
or U5241 (N_5241,N_4729,N_3061);
nand U5242 (N_5242,N_3551,N_4892);
xor U5243 (N_5243,N_4391,N_2502);
nand U5244 (N_5244,N_4716,N_4929);
or U5245 (N_5245,N_4114,N_4365);
nor U5246 (N_5246,N_4834,N_3112);
nor U5247 (N_5247,N_4845,N_4630);
xnor U5248 (N_5248,N_4922,N_4983);
nand U5249 (N_5249,N_4468,N_3053);
xnor U5250 (N_5250,N_3871,N_3027);
nand U5251 (N_5251,N_3370,N_4152);
and U5252 (N_5252,N_3675,N_2737);
nand U5253 (N_5253,N_3952,N_3233);
nor U5254 (N_5254,N_4345,N_3106);
nand U5255 (N_5255,N_3187,N_2699);
nor U5256 (N_5256,N_4321,N_3069);
nor U5257 (N_5257,N_4467,N_4101);
or U5258 (N_5258,N_4332,N_2835);
nor U5259 (N_5259,N_4409,N_3251);
nand U5260 (N_5260,N_3248,N_4318);
nand U5261 (N_5261,N_4953,N_4404);
nor U5262 (N_5262,N_2912,N_4339);
nand U5263 (N_5263,N_4937,N_3446);
nor U5264 (N_5264,N_3253,N_3165);
nand U5265 (N_5265,N_3556,N_2829);
or U5266 (N_5266,N_3901,N_2931);
or U5267 (N_5267,N_2984,N_3781);
nand U5268 (N_5268,N_4750,N_2857);
xor U5269 (N_5269,N_3815,N_3137);
xor U5270 (N_5270,N_3122,N_3265);
nor U5271 (N_5271,N_4975,N_3408);
or U5272 (N_5272,N_4598,N_3884);
and U5273 (N_5273,N_4900,N_4087);
nor U5274 (N_5274,N_4074,N_3070);
and U5275 (N_5275,N_4273,N_3662);
nor U5276 (N_5276,N_2509,N_4752);
or U5277 (N_5277,N_4408,N_4963);
nor U5278 (N_5278,N_3574,N_3735);
nand U5279 (N_5279,N_4153,N_2993);
nand U5280 (N_5280,N_3042,N_2554);
or U5281 (N_5281,N_3682,N_2559);
and U5282 (N_5282,N_3575,N_2792);
nand U5283 (N_5283,N_3916,N_4701);
or U5284 (N_5284,N_2592,N_3887);
nand U5285 (N_5285,N_2511,N_2886);
nand U5286 (N_5286,N_2819,N_2644);
xnor U5287 (N_5287,N_3059,N_3355);
or U5288 (N_5288,N_3400,N_2909);
or U5289 (N_5289,N_4301,N_3954);
and U5290 (N_5290,N_2656,N_4262);
and U5291 (N_5291,N_4324,N_2573);
nand U5292 (N_5292,N_2769,N_2780);
nand U5293 (N_5293,N_4553,N_3830);
or U5294 (N_5294,N_3166,N_3361);
nand U5295 (N_5295,N_3617,N_4055);
and U5296 (N_5296,N_2553,N_4979);
or U5297 (N_5297,N_4987,N_4531);
and U5298 (N_5298,N_4062,N_3736);
xnor U5299 (N_5299,N_4185,N_4886);
nand U5300 (N_5300,N_3107,N_3824);
xnor U5301 (N_5301,N_4032,N_4532);
xor U5302 (N_5302,N_3842,N_2774);
and U5303 (N_5303,N_3774,N_3114);
nor U5304 (N_5304,N_4880,N_4290);
or U5305 (N_5305,N_2943,N_3500);
and U5306 (N_5306,N_3001,N_4648);
and U5307 (N_5307,N_4003,N_3613);
or U5308 (N_5308,N_3456,N_2524);
or U5309 (N_5309,N_3853,N_4395);
nor U5310 (N_5310,N_3058,N_3514);
or U5311 (N_5311,N_3384,N_3089);
nand U5312 (N_5312,N_3144,N_4158);
nor U5313 (N_5313,N_3627,N_3419);
xnor U5314 (N_5314,N_3183,N_4245);
and U5315 (N_5315,N_3834,N_3725);
nor U5316 (N_5316,N_3580,N_2535);
nand U5317 (N_5317,N_3067,N_2594);
nand U5318 (N_5318,N_4094,N_4222);
and U5319 (N_5319,N_3873,N_4265);
nor U5320 (N_5320,N_3349,N_3770);
xnor U5321 (N_5321,N_4905,N_2603);
nor U5322 (N_5322,N_3858,N_4873);
nand U5323 (N_5323,N_3732,N_4420);
and U5324 (N_5324,N_3085,N_4314);
and U5325 (N_5325,N_3459,N_3173);
xnor U5326 (N_5326,N_4902,N_3814);
nor U5327 (N_5327,N_2724,N_4122);
nor U5328 (N_5328,N_3188,N_4258);
xor U5329 (N_5329,N_3565,N_4967);
nor U5330 (N_5330,N_2784,N_4102);
and U5331 (N_5331,N_4909,N_2919);
or U5332 (N_5332,N_4990,N_4684);
nand U5333 (N_5333,N_3542,N_4449);
nand U5334 (N_5334,N_3508,N_3014);
xnor U5335 (N_5335,N_2789,N_2761);
and U5336 (N_5336,N_3892,N_3467);
and U5337 (N_5337,N_4026,N_4628);
xor U5338 (N_5338,N_2718,N_4817);
or U5339 (N_5339,N_3727,N_4792);
nand U5340 (N_5340,N_3604,N_2733);
and U5341 (N_5341,N_4942,N_4772);
nor U5342 (N_5342,N_3896,N_4439);
or U5343 (N_5343,N_3197,N_2523);
nand U5344 (N_5344,N_3561,N_3636);
nor U5345 (N_5345,N_3395,N_4056);
and U5346 (N_5346,N_2815,N_4948);
and U5347 (N_5347,N_2878,N_4853);
nand U5348 (N_5348,N_3431,N_3013);
nor U5349 (N_5349,N_4851,N_3897);
nand U5350 (N_5350,N_2500,N_4549);
nor U5351 (N_5351,N_2538,N_3481);
nor U5352 (N_5352,N_4274,N_4991);
xor U5353 (N_5353,N_4260,N_3324);
or U5354 (N_5354,N_4405,N_4025);
or U5355 (N_5355,N_4550,N_3426);
and U5356 (N_5356,N_2906,N_2743);
nand U5357 (N_5357,N_3452,N_3667);
or U5358 (N_5358,N_4986,N_4919);
and U5359 (N_5359,N_4475,N_2807);
nand U5360 (N_5360,N_4435,N_2890);
xor U5361 (N_5361,N_2611,N_4506);
and U5362 (N_5362,N_4076,N_4325);
nand U5363 (N_5363,N_4485,N_4461);
and U5364 (N_5364,N_3597,N_3177);
nand U5365 (N_5365,N_3010,N_3126);
and U5366 (N_5366,N_4021,N_4590);
nand U5367 (N_5367,N_4088,N_4812);
and U5368 (N_5368,N_4396,N_3346);
nand U5369 (N_5369,N_3258,N_3222);
nand U5370 (N_5370,N_3231,N_4355);
or U5371 (N_5371,N_2701,N_4788);
nand U5372 (N_5372,N_4650,N_4547);
or U5373 (N_5373,N_3369,N_3139);
or U5374 (N_5374,N_3749,N_3090);
xor U5375 (N_5375,N_4918,N_4370);
or U5376 (N_5376,N_4747,N_3462);
xnor U5377 (N_5377,N_3806,N_3421);
xor U5378 (N_5378,N_3079,N_4005);
or U5379 (N_5379,N_3902,N_4131);
and U5380 (N_5380,N_3143,N_2964);
or U5381 (N_5381,N_2505,N_3390);
nand U5382 (N_5382,N_3071,N_2747);
nor U5383 (N_5383,N_2883,N_4368);
and U5384 (N_5384,N_3645,N_3584);
nor U5385 (N_5385,N_3699,N_4658);
nor U5386 (N_5386,N_3157,N_3360);
nand U5387 (N_5387,N_3506,N_2837);
nand U5388 (N_5388,N_3942,N_4149);
nor U5389 (N_5389,N_4111,N_3430);
xnor U5390 (N_5390,N_3095,N_4380);
and U5391 (N_5391,N_4219,N_3184);
or U5392 (N_5392,N_4735,N_3787);
or U5393 (N_5393,N_4415,N_4394);
nand U5394 (N_5394,N_4234,N_3316);
nor U5395 (N_5395,N_3581,N_4465);
nand U5396 (N_5396,N_2929,N_3476);
xnor U5397 (N_5397,N_2615,N_4009);
and U5398 (N_5398,N_4751,N_3282);
or U5399 (N_5399,N_4344,N_2641);
nor U5400 (N_5400,N_4760,N_3837);
nand U5401 (N_5401,N_4492,N_2746);
or U5402 (N_5402,N_4237,N_3612);
nor U5403 (N_5403,N_3661,N_4469);
and U5404 (N_5404,N_3933,N_3016);
nand U5405 (N_5405,N_2759,N_4645);
or U5406 (N_5406,N_4799,N_4037);
nor U5407 (N_5407,N_4842,N_3533);
nor U5408 (N_5408,N_4719,N_3284);
nand U5409 (N_5409,N_2653,N_4418);
nand U5410 (N_5410,N_2961,N_4279);
xnor U5411 (N_5411,N_3971,N_4431);
nor U5412 (N_5412,N_3295,N_4228);
nand U5413 (N_5413,N_3980,N_3342);
nand U5414 (N_5414,N_4217,N_4609);
and U5415 (N_5415,N_4349,N_3213);
or U5416 (N_5416,N_4328,N_4125);
nor U5417 (N_5417,N_4454,N_3094);
nand U5418 (N_5418,N_3672,N_4388);
xor U5419 (N_5419,N_4187,N_3210);
or U5420 (N_5420,N_2907,N_3364);
xnor U5421 (N_5421,N_4011,N_3563);
nor U5422 (N_5422,N_2683,N_4338);
nand U5423 (N_5423,N_4730,N_3273);
and U5424 (N_5424,N_4063,N_3972);
or U5425 (N_5425,N_4095,N_4453);
nand U5426 (N_5426,N_3908,N_4171);
or U5427 (N_5427,N_4495,N_3482);
and U5428 (N_5428,N_3680,N_2680);
or U5429 (N_5429,N_4113,N_4090);
xnor U5430 (N_5430,N_3435,N_2740);
xnor U5431 (N_5431,N_2899,N_3726);
or U5432 (N_5432,N_3763,N_4578);
and U5433 (N_5433,N_4697,N_4971);
or U5434 (N_5434,N_2695,N_3737);
or U5435 (N_5435,N_3261,N_4858);
xnor U5436 (N_5436,N_2790,N_4346);
and U5437 (N_5437,N_4580,N_4661);
nand U5438 (N_5438,N_4109,N_2715);
and U5439 (N_5439,N_2501,N_4127);
and U5440 (N_5440,N_2720,N_3609);
xnor U5441 (N_5441,N_3951,N_3686);
and U5442 (N_5442,N_2670,N_3102);
nand U5443 (N_5443,N_4872,N_3518);
xor U5444 (N_5444,N_3856,N_3232);
nor U5445 (N_5445,N_4733,N_4170);
and U5446 (N_5446,N_4416,N_4278);
xnor U5447 (N_5447,N_3150,N_2686);
and U5448 (N_5448,N_4670,N_4753);
and U5449 (N_5449,N_2548,N_3962);
xnor U5450 (N_5450,N_2510,N_4266);
nand U5451 (N_5451,N_3592,N_3164);
xor U5452 (N_5452,N_4838,N_4142);
or U5453 (N_5453,N_4599,N_3386);
nand U5454 (N_5454,N_3937,N_2546);
nand U5455 (N_5455,N_4285,N_3554);
nand U5456 (N_5456,N_4717,N_3147);
or U5457 (N_5457,N_4452,N_3792);
and U5458 (N_5458,N_4704,N_3031);
xnor U5459 (N_5459,N_2934,N_3333);
or U5460 (N_5460,N_2768,N_4412);
or U5461 (N_5461,N_4808,N_2756);
nand U5462 (N_5462,N_3955,N_3977);
or U5463 (N_5463,N_4340,N_3845);
nand U5464 (N_5464,N_2873,N_3474);
nand U5465 (N_5465,N_2823,N_3844);
nor U5466 (N_5466,N_3491,N_3938);
nand U5467 (N_5467,N_4426,N_4291);
and U5468 (N_5468,N_4378,N_3297);
nor U5469 (N_5469,N_3005,N_3380);
nand U5470 (N_5470,N_4035,N_2614);
nand U5471 (N_5471,N_3803,N_3729);
and U5472 (N_5472,N_4491,N_4463);
or U5473 (N_5473,N_4223,N_2716);
nand U5474 (N_5474,N_3705,N_3782);
xnor U5475 (N_5475,N_3201,N_4466);
nand U5476 (N_5476,N_2751,N_4722);
and U5477 (N_5477,N_3241,N_3519);
xor U5478 (N_5478,N_4226,N_3132);
or U5479 (N_5479,N_3825,N_3442);
and U5480 (N_5480,N_2668,N_3802);
xnor U5481 (N_5481,N_2604,N_4559);
xor U5482 (N_5482,N_4754,N_3547);
and U5483 (N_5483,N_3940,N_3242);
xor U5484 (N_5484,N_4181,N_3986);
and U5485 (N_5485,N_3099,N_4244);
or U5486 (N_5486,N_3169,N_3936);
nand U5487 (N_5487,N_4134,N_2824);
nand U5488 (N_5488,N_4714,N_4917);
nand U5489 (N_5489,N_4264,N_4039);
xor U5490 (N_5490,N_3021,N_3917);
xor U5491 (N_5491,N_3988,N_4041);
nand U5492 (N_5492,N_3877,N_2891);
nor U5493 (N_5493,N_3812,N_4186);
and U5494 (N_5494,N_3484,N_4373);
nor U5495 (N_5495,N_4640,N_4689);
nand U5496 (N_5496,N_4930,N_4712);
or U5497 (N_5497,N_3723,N_3285);
xnor U5498 (N_5498,N_2841,N_3925);
xor U5499 (N_5499,N_3409,N_4720);
or U5500 (N_5500,N_4410,N_4800);
or U5501 (N_5501,N_3665,N_2989);
nor U5502 (N_5502,N_4128,N_3024);
nor U5503 (N_5503,N_4140,N_4583);
xor U5504 (N_5504,N_3872,N_2601);
or U5505 (N_5505,N_2879,N_3142);
nand U5506 (N_5506,N_3485,N_4820);
nand U5507 (N_5507,N_4803,N_4386);
nand U5508 (N_5508,N_4618,N_4556);
nor U5509 (N_5509,N_3034,N_2635);
nand U5510 (N_5510,N_4313,N_4796);
and U5511 (N_5511,N_3216,N_3263);
nand U5512 (N_5512,N_4841,N_3949);
or U5513 (N_5513,N_3867,N_4471);
nand U5514 (N_5514,N_4286,N_3411);
nor U5515 (N_5515,N_2897,N_3619);
or U5516 (N_5516,N_4920,N_4146);
nand U5517 (N_5517,N_4680,N_3764);
nor U5518 (N_5518,N_4307,N_2945);
and U5519 (N_5519,N_4927,N_2987);
nand U5520 (N_5520,N_3866,N_2735);
or U5521 (N_5521,N_3463,N_3578);
xnor U5522 (N_5522,N_3523,N_4746);
nand U5523 (N_5523,N_4082,N_2808);
and U5524 (N_5524,N_2875,N_4907);
xor U5525 (N_5525,N_4369,N_4544);
and U5526 (N_5526,N_3570,N_3839);
xnor U5527 (N_5527,N_4429,N_2966);
nand U5528 (N_5528,N_4357,N_3308);
nand U5529 (N_5529,N_2856,N_3785);
or U5530 (N_5530,N_2978,N_2799);
and U5531 (N_5531,N_2930,N_3895);
xor U5532 (N_5532,N_3255,N_3002);
nor U5533 (N_5533,N_4965,N_3341);
or U5534 (N_5534,N_2655,N_2714);
nand U5535 (N_5535,N_4078,N_2944);
nand U5536 (N_5536,N_4736,N_3797);
nand U5537 (N_5537,N_3162,N_2522);
nand U5538 (N_5538,N_4740,N_2896);
nor U5539 (N_5539,N_3642,N_3924);
xor U5540 (N_5540,N_4673,N_4555);
xnor U5541 (N_5541,N_3701,N_2921);
nand U5542 (N_5542,N_2730,N_4382);
and U5543 (N_5543,N_2933,N_3007);
nand U5544 (N_5544,N_4623,N_4870);
xnor U5545 (N_5545,N_4288,N_3541);
or U5546 (N_5546,N_4455,N_3301);
xnor U5547 (N_5547,N_4955,N_2690);
or U5548 (N_5548,N_4763,N_3375);
or U5549 (N_5549,N_4656,N_4077);
xor U5550 (N_5550,N_4372,N_3835);
nor U5551 (N_5551,N_3906,N_4135);
or U5552 (N_5552,N_3009,N_3449);
and U5553 (N_5553,N_4423,N_3046);
nand U5554 (N_5554,N_2810,N_3145);
nand U5555 (N_5555,N_3438,N_4436);
or U5556 (N_5556,N_4161,N_4928);
and U5557 (N_5557,N_4923,N_4621);
xor U5558 (N_5558,N_4441,N_3663);
nand U5559 (N_5559,N_4384,N_4775);
nand U5560 (N_5560,N_4322,N_3424);
xor U5561 (N_5561,N_4203,N_4104);
nand U5562 (N_5562,N_4831,N_2530);
xnor U5563 (N_5563,N_4115,N_3857);
nand U5564 (N_5564,N_3836,N_2629);
nand U5565 (N_5565,N_3326,N_3633);
and U5566 (N_5566,N_4903,N_4331);
and U5567 (N_5567,N_2549,N_4207);
nor U5568 (N_5568,N_3862,N_2764);
nand U5569 (N_5569,N_4862,N_4554);
and U5570 (N_5570,N_4894,N_3990);
nand U5571 (N_5571,N_2617,N_4427);
nand U5572 (N_5572,N_3791,N_4048);
and U5573 (N_5573,N_3041,N_4188);
xor U5574 (N_5574,N_2648,N_3281);
nor U5575 (N_5575,N_3869,N_4978);
nor U5576 (N_5576,N_4065,N_4687);
and U5577 (N_5577,N_3961,N_3553);
and U5578 (N_5578,N_4608,N_4952);
nor U5579 (N_5579,N_2624,N_4791);
and U5580 (N_5580,N_2659,N_4284);
and U5581 (N_5581,N_4276,N_3534);
nand U5582 (N_5582,N_3789,N_3929);
and U5583 (N_5583,N_3072,N_3620);
or U5584 (N_5584,N_3280,N_2578);
xnor U5585 (N_5585,N_3055,N_4173);
or U5586 (N_5586,N_3799,N_2515);
xor U5587 (N_5587,N_2512,N_4866);
xnor U5588 (N_5588,N_3595,N_3640);
xnor U5589 (N_5589,N_4249,N_2642);
and U5590 (N_5590,N_3540,N_2599);
nand U5591 (N_5591,N_2809,N_4042);
xor U5592 (N_5592,N_4085,N_3488);
nand U5593 (N_5593,N_4303,N_4364);
or U5594 (N_5594,N_3011,N_2754);
and U5595 (N_5595,N_3577,N_3694);
or U5596 (N_5596,N_4267,N_4347);
nor U5597 (N_5597,N_4806,N_3760);
and U5598 (N_5598,N_3205,N_2881);
nor U5599 (N_5599,N_2960,N_3256);
and U5600 (N_5600,N_4432,N_2869);
xnor U5601 (N_5601,N_4829,N_4411);
and U5602 (N_5602,N_4044,N_4566);
xnor U5603 (N_5603,N_4767,N_3741);
xnor U5604 (N_5604,N_3321,N_2806);
or U5605 (N_5605,N_4579,N_3203);
and U5606 (N_5606,N_2529,N_4850);
nand U5607 (N_5607,N_4327,N_4243);
nand U5608 (N_5608,N_3133,N_4739);
and U5609 (N_5609,N_2543,N_4509);
or U5610 (N_5610,N_3451,N_4766);
nor U5611 (N_5611,N_3800,N_4238);
nand U5612 (N_5612,N_4050,N_4931);
and U5613 (N_5613,N_2638,N_3300);
and U5614 (N_5614,N_3847,N_4075);
and U5615 (N_5615,N_4494,N_4257);
nand U5616 (N_5616,N_4235,N_3798);
nor U5617 (N_5617,N_2628,N_4106);
or U5618 (N_5618,N_3966,N_4329);
xnor U5619 (N_5619,N_2757,N_2750);
nor U5620 (N_5620,N_3637,N_4474);
nand U5621 (N_5621,N_4178,N_3771);
nor U5622 (N_5622,N_4014,N_4686);
xnor U5623 (N_5623,N_3176,N_4336);
nand U5624 (N_5624,N_3821,N_4472);
nand U5625 (N_5625,N_2669,N_4798);
nand U5626 (N_5626,N_4691,N_4473);
nand U5627 (N_5627,N_4479,N_4537);
and U5628 (N_5628,N_4671,N_3707);
and U5629 (N_5629,N_3155,N_3294);
and U5630 (N_5630,N_3286,N_2634);
and U5631 (N_5631,N_2816,N_3289);
or U5632 (N_5632,N_4849,N_4417);
xnor U5633 (N_5633,N_2539,N_3911);
nand U5634 (N_5634,N_4482,N_4289);
nor U5635 (N_5635,N_2791,N_3734);
xnor U5636 (N_5636,N_2694,N_3272);
xnor U5637 (N_5637,N_3262,N_3311);
nor U5638 (N_5638,N_4968,N_3779);
and U5639 (N_5639,N_3585,N_3214);
xnor U5640 (N_5640,N_3192,N_3599);
nand U5641 (N_5641,N_3146,N_3420);
and U5642 (N_5642,N_3352,N_4724);
nand U5643 (N_5643,N_2706,N_4091);
nand U5644 (N_5644,N_2758,N_3973);
nand U5645 (N_5645,N_3498,N_3848);
and U5646 (N_5646,N_2691,N_3054);
nor U5647 (N_5647,N_3720,N_3646);
and U5648 (N_5648,N_4964,N_4169);
xnor U5649 (N_5649,N_4069,N_4809);
or U5650 (N_5650,N_4976,N_3429);
nor U5651 (N_5651,N_3568,N_3820);
or U5652 (N_5652,N_2836,N_4051);
xnor U5653 (N_5653,N_4046,N_3103);
nand U5654 (N_5654,N_4522,N_4080);
nor U5655 (N_5655,N_3357,N_4123);
or U5656 (N_5656,N_3852,N_2946);
nand U5657 (N_5657,N_3600,N_2584);
and U5658 (N_5658,N_2723,N_4662);
and U5659 (N_5659,N_3606,N_3097);
nor U5660 (N_5660,N_3840,N_4597);
nand U5661 (N_5661,N_4403,N_3464);
nor U5662 (N_5662,N_3963,N_4296);
xor U5663 (N_5663,N_3296,N_4595);
xnor U5664 (N_5664,N_3524,N_4676);
or U5665 (N_5665,N_2721,N_4844);
nor U5666 (N_5666,N_3643,N_4498);
and U5667 (N_5667,N_2870,N_4450);
nor U5668 (N_5668,N_3711,N_3448);
nand U5669 (N_5669,N_4107,N_4773);
and U5670 (N_5670,N_4254,N_2698);
nor U5671 (N_5671,N_4199,N_2914);
and U5672 (N_5672,N_4548,N_4478);
or U5673 (N_5673,N_2517,N_3358);
nand U5674 (N_5674,N_4093,N_3257);
nand U5675 (N_5675,N_3047,N_3240);
xor U5676 (N_5676,N_2813,N_4263);
and U5677 (N_5677,N_3587,N_3365);
nor U5678 (N_5678,N_3076,N_3298);
xnor U5679 (N_5679,N_3808,N_4381);
and U5680 (N_5680,N_3605,N_2811);
or U5681 (N_5681,N_2685,N_4496);
or U5682 (N_5682,N_2542,N_4022);
or U5683 (N_5683,N_2545,N_2602);
or U5684 (N_5684,N_4280,N_4731);
nand U5685 (N_5685,N_2556,N_3066);
nand U5686 (N_5686,N_4958,N_3922);
nand U5687 (N_5687,N_3313,N_3065);
or U5688 (N_5688,N_3381,N_2992);
and U5689 (N_5689,N_3170,N_2547);
or U5690 (N_5690,N_4241,N_2963);
nand U5691 (N_5691,N_3290,N_3274);
nor U5692 (N_5692,N_4582,N_4588);
or U5693 (N_5693,N_3379,N_2609);
xor U5694 (N_5694,N_4527,N_4741);
or U5695 (N_5695,N_3926,N_3044);
xor U5696 (N_5696,N_3513,N_3886);
nor U5697 (N_5697,N_3615,N_3529);
and U5698 (N_5698,N_3135,N_4358);
nand U5699 (N_5699,N_2920,N_3536);
nor U5700 (N_5700,N_3080,N_3330);
or U5701 (N_5701,N_3336,N_4001);
nand U5702 (N_5702,N_4231,N_3270);
xnor U5703 (N_5703,N_3754,N_3505);
nand U5704 (N_5704,N_4825,N_4477);
xor U5705 (N_5705,N_3984,N_4934);
and U5706 (N_5706,N_3458,N_3471);
or U5707 (N_5707,N_4103,N_3527);
and U5708 (N_5708,N_2739,N_2955);
nor U5709 (N_5709,N_2541,N_2630);
or U5710 (N_5710,N_4252,N_3677);
or U5711 (N_5711,N_2647,N_3174);
or U5712 (N_5712,N_3399,N_4512);
or U5713 (N_5713,N_2986,N_2672);
nor U5714 (N_5714,N_4912,N_4305);
nor U5715 (N_5715,N_3495,N_3875);
and U5716 (N_5716,N_3697,N_3338);
and U5717 (N_5717,N_4748,N_2591);
nand U5718 (N_5718,N_4043,N_4066);
and U5719 (N_5719,N_2994,N_4271);
xor U5720 (N_5720,N_4619,N_2939);
nor U5721 (N_5721,N_4379,N_3199);
xnor U5722 (N_5722,N_4764,N_4668);
or U5723 (N_5723,N_4451,N_4027);
and U5724 (N_5724,N_3276,N_4666);
and U5725 (N_5725,N_3614,N_4836);
xnor U5726 (N_5726,N_3991,N_2506);
or U5727 (N_5727,N_2901,N_3140);
nor U5728 (N_5728,N_3522,N_3483);
xor U5729 (N_5729,N_2508,N_2674);
and U5730 (N_5730,N_3064,N_4413);
or U5731 (N_5731,N_2552,N_3220);
nand U5732 (N_5732,N_4281,N_4007);
or U5733 (N_5733,N_4503,N_3026);
xnor U5734 (N_5734,N_4652,N_4790);
and U5735 (N_5735,N_3503,N_4816);
or U5736 (N_5736,N_3100,N_3860);
nand U5737 (N_5737,N_2738,N_4534);
xor U5738 (N_5738,N_3202,N_3557);
nor U5739 (N_5739,N_3068,N_3978);
and U5740 (N_5740,N_3653,N_3217);
or U5741 (N_5741,N_4946,N_3407);
or U5742 (N_5742,N_4957,N_2795);
xnor U5743 (N_5743,N_4647,N_4639);
or U5744 (N_5744,N_3303,N_4573);
and U5745 (N_5745,N_4002,N_4794);
or U5746 (N_5746,N_2608,N_3888);
nor U5747 (N_5747,N_2582,N_3510);
nor U5748 (N_5748,N_2607,N_2585);
and U5749 (N_5749,N_3528,N_3039);
xor U5750 (N_5750,N_4520,N_4390);
and U5751 (N_5751,N_3383,N_3299);
nor U5752 (N_5752,N_4901,N_4956);
nor U5753 (N_5753,N_3291,N_3603);
xnor U5754 (N_5754,N_4246,N_4189);
or U5755 (N_5755,N_3182,N_4206);
or U5756 (N_5756,N_2703,N_3722);
nand U5757 (N_5757,N_3032,N_2709);
or U5758 (N_5758,N_3765,N_3186);
xor U5759 (N_5759,N_3323,N_3078);
xor U5760 (N_5760,N_4040,N_3904);
or U5761 (N_5761,N_4822,N_4996);
and U5762 (N_5762,N_4657,N_2814);
and U5763 (N_5763,N_3930,N_2677);
nand U5764 (N_5764,N_4193,N_3761);
nor U5765 (N_5765,N_4392,N_3416);
nor U5766 (N_5766,N_4272,N_2616);
nor U5767 (N_5767,N_2689,N_4581);
or U5768 (N_5768,N_4706,N_3287);
or U5769 (N_5769,N_3224,N_3056);
xor U5770 (N_5770,N_4462,N_2667);
nand U5771 (N_5771,N_3579,N_4397);
or U5772 (N_5772,N_4560,N_4068);
or U5773 (N_5773,N_4543,N_4334);
nor U5774 (N_5774,N_4438,N_4017);
nand U5775 (N_5775,N_4126,N_3468);
and U5776 (N_5776,N_2697,N_4605);
nor U5777 (N_5777,N_3946,N_3437);
nor U5778 (N_5778,N_4172,N_4916);
and U5779 (N_5779,N_4195,N_4810);
and U5780 (N_5780,N_4742,N_2631);
nand U5781 (N_5781,N_3247,N_3742);
or U5782 (N_5782,N_2568,N_2565);
and U5783 (N_5783,N_2681,N_4881);
and U5784 (N_5784,N_2671,N_2722);
nor U5785 (N_5785,N_4985,N_2605);
xor U5786 (N_5786,N_3152,N_4367);
and U5787 (N_5787,N_4593,N_4745);
nor U5788 (N_5788,N_3215,N_4184);
xnor U5789 (N_5789,N_3716,N_3405);
xor U5790 (N_5790,N_3976,N_2513);
nand U5791 (N_5791,N_4458,N_4197);
or U5792 (N_5792,N_2818,N_3480);
or U5793 (N_5793,N_4707,N_4456);
nor U5794 (N_5794,N_4804,N_3809);
or U5795 (N_5795,N_3944,N_4692);
nand U5796 (N_5796,N_3807,N_3037);
nand U5797 (N_5797,N_4654,N_4802);
nand U5798 (N_5798,N_2643,N_3181);
nand U5799 (N_5799,N_2526,N_3243);
nor U5800 (N_5800,N_3621,N_3269);
xnor U5801 (N_5801,N_2975,N_2707);
nand U5802 (N_5802,N_4098,N_2687);
and U5803 (N_5803,N_3562,N_3124);
or U5804 (N_5804,N_3023,N_4536);
nor U5805 (N_5805,N_2576,N_4672);
nor U5806 (N_5806,N_3591,N_4585);
or U5807 (N_5807,N_4695,N_2767);
nor U5808 (N_5808,N_3752,N_4574);
nor U5809 (N_5809,N_4744,N_2832);
nor U5810 (N_5810,N_3957,N_4824);
and U5811 (N_5811,N_2951,N_4565);
and U5812 (N_5812,N_4162,N_3520);
nor U5813 (N_5813,N_4121,N_4159);
nand U5814 (N_5814,N_4679,N_4356);
and U5815 (N_5815,N_3334,N_2507);
nor U5816 (N_5816,N_2700,N_3159);
xnor U5817 (N_5817,N_3314,N_4625);
and U5818 (N_5818,N_4539,N_3850);
nand U5819 (N_5819,N_3773,N_3882);
nor U5820 (N_5820,N_4352,N_4061);
or U5821 (N_5821,N_4157,N_2913);
and U5822 (N_5822,N_4564,N_4298);
xor U5823 (N_5823,N_4541,N_3335);
or U5824 (N_5824,N_3081,N_4586);
and U5825 (N_5825,N_2976,N_3325);
nand U5826 (N_5826,N_4999,N_4073);
xor U5827 (N_5827,N_2839,N_4275);
nor U5828 (N_5828,N_4256,N_3060);
and U5829 (N_5829,N_4422,N_3185);
nand U5830 (N_5830,N_2922,N_3525);
nand U5831 (N_5831,N_3628,N_3156);
nand U5832 (N_5832,N_4882,N_3093);
xnor U5833 (N_5833,N_4884,N_4137);
or U5834 (N_5834,N_4703,N_4242);
and U5835 (N_5835,N_3702,N_3685);
or U5836 (N_5836,N_4801,N_4828);
or U5837 (N_5837,N_3394,N_2848);
nor U5838 (N_5838,N_4086,N_4627);
nor U5839 (N_5839,N_3816,N_4194);
nor U5840 (N_5840,N_4857,N_3721);
or U5841 (N_5841,N_3987,N_3450);
nor U5842 (N_5842,N_3740,N_3501);
nor U5843 (N_5843,N_4371,N_3320);
and U5844 (N_5844,N_2755,N_4060);
nor U5845 (N_5845,N_4192,N_3486);
or U5846 (N_5846,N_3453,N_3317);
or U5847 (N_5847,N_2521,N_3631);
nor U5848 (N_5848,N_2525,N_4663);
or U5849 (N_5849,N_2531,N_3084);
and U5850 (N_5850,N_4869,N_4538);
or U5851 (N_5851,N_2777,N_4312);
xor U5852 (N_5852,N_4407,N_3461);
or U5853 (N_5853,N_3610,N_3532);
nor U5854 (N_5854,N_4913,N_3608);
nand U5855 (N_5855,N_4992,N_4562);
xor U5856 (N_5856,N_3127,N_3193);
nand U5857 (N_5857,N_4215,N_3535);
xnor U5858 (N_5858,N_3582,N_3905);
xor U5859 (N_5859,N_3322,N_2846);
and U5860 (N_5860,N_3211,N_3784);
nand U5861 (N_5861,N_4362,N_3530);
nand U5862 (N_5862,N_3195,N_4777);
nor U5863 (N_5863,N_3589,N_3624);
nor U5864 (N_5864,N_3331,N_3028);
xor U5865 (N_5865,N_4688,N_4024);
nor U5866 (N_5866,N_2863,N_2577);
nor U5867 (N_5867,N_2595,N_3278);
nand U5868 (N_5868,N_4938,N_4015);
nand U5869 (N_5869,N_4525,N_3828);
nor U5870 (N_5870,N_3225,N_4160);
or U5871 (N_5871,N_3639,N_4179);
or U5872 (N_5872,N_2763,N_2887);
or U5873 (N_5873,N_4587,N_3851);
or U5874 (N_5874,N_4227,N_4425);
xor U5875 (N_5875,N_3969,N_3777);
and U5876 (N_5876,N_4563,N_4168);
or U5877 (N_5877,N_4047,N_3583);
xnor U5878 (N_5878,N_3507,N_4830);
nor U5879 (N_5879,N_2600,N_2820);
or U5880 (N_5880,N_4944,N_2649);
nand U5881 (N_5881,N_3454,N_4428);
and U5882 (N_5882,N_3868,N_2696);
nor U5883 (N_5883,N_4138,N_2623);
xnor U5884 (N_5884,N_4302,N_3268);
nor U5885 (N_5885,N_4819,N_4721);
nor U5886 (N_5886,N_4675,N_3305);
and U5887 (N_5887,N_4283,N_3478);
xor U5888 (N_5888,N_2941,N_2620);
and U5889 (N_5889,N_3368,N_3306);
xnor U5890 (N_5890,N_3235,N_3718);
nand U5891 (N_5891,N_2970,N_4488);
nand U5892 (N_5892,N_2678,N_2742);
or U5893 (N_5893,N_4036,N_4165);
nor U5894 (N_5894,N_3945,N_4070);
nor U5895 (N_5895,N_3279,N_2908);
nand U5896 (N_5896,N_3719,N_3918);
nor U5897 (N_5897,N_4821,N_4433);
xnor U5898 (N_5898,N_2771,N_2781);
xnor U5899 (N_5899,N_3393,N_4856);
nand U5900 (N_5900,N_2868,N_3040);
xnor U5901 (N_5901,N_4163,N_4443);
or U5902 (N_5902,N_3638,N_3490);
nand U5903 (N_5903,N_3515,N_3238);
nand U5904 (N_5904,N_2988,N_2845);
xor U5905 (N_5905,N_2560,N_3465);
and U5906 (N_5906,N_4732,N_3652);
nand U5907 (N_5907,N_3632,N_4980);
or U5908 (N_5908,N_3832,N_4201);
nand U5909 (N_5909,N_3350,N_2663);
xnor U5910 (N_5910,N_4486,N_2861);
nor U5911 (N_5911,N_2990,N_4053);
xor U5912 (N_5912,N_4659,N_3239);
nand U5913 (N_5913,N_3859,N_4646);
nand U5914 (N_5914,N_3392,N_4726);
and U5915 (N_5915,N_4514,N_4348);
or U5916 (N_5916,N_3693,N_3863);
xor U5917 (N_5917,N_3810,N_3819);
nand U5918 (N_5918,N_4540,N_4414);
and U5919 (N_5919,N_4204,N_2797);
or U5920 (N_5920,N_4954,N_2911);
and U5921 (N_5921,N_4651,N_3998);
xnor U5922 (N_5922,N_4725,N_2708);
xnor U5923 (N_5923,N_4521,N_2871);
and U5924 (N_5924,N_3586,N_2519);
nand U5925 (N_5925,N_4926,N_4622);
xor U5926 (N_5926,N_4212,N_2712);
nor U5927 (N_5927,N_4932,N_2884);
and U5928 (N_5928,N_3022,N_2516);
or U5929 (N_5929,N_4989,N_3315);
nor U5930 (N_5930,N_3417,N_4604);
and U5931 (N_5931,N_4517,N_4643);
nand U5932 (N_5932,N_4755,N_4510);
nand U5933 (N_5933,N_3460,N_4139);
xnor U5934 (N_5934,N_4389,N_4962);
xor U5935 (N_5935,N_3688,N_4795);
xor U5936 (N_5936,N_2711,N_2566);
nor U5937 (N_5937,N_4008,N_4813);
nand U5938 (N_5938,N_3436,N_3414);
nand U5939 (N_5939,N_3019,N_3864);
nand U5940 (N_5940,N_2651,N_3715);
xnor U5941 (N_5941,N_4569,N_2613);
nor U5942 (N_5942,N_4424,N_3509);
or U5943 (N_5943,N_3569,N_4268);
and U5944 (N_5944,N_4214,N_4634);
nor U5945 (N_5945,N_4054,N_3706);
xor U5946 (N_5946,N_2853,N_3372);
nand U5947 (N_5947,N_2979,N_2783);
xnor U5948 (N_5948,N_3928,N_4202);
nor U5949 (N_5949,N_3826,N_4785);
nor U5950 (N_5950,N_3913,N_4470);
nor U5951 (N_5951,N_4004,N_2860);
xnor U5952 (N_5952,N_4079,N_4330);
and U5953 (N_5953,N_3841,N_2562);
and U5954 (N_5954,N_3687,N_3689);
nand U5955 (N_5955,N_3151,N_4626);
nor U5956 (N_5956,N_3345,N_4665);
or U5957 (N_5957,N_4558,N_3440);
nor U5958 (N_5958,N_3207,N_2938);
xnor U5959 (N_5959,N_3310,N_4713);
and U5960 (N_5960,N_3915,N_3531);
nor U5961 (N_5961,N_4295,N_2787);
or U5962 (N_5962,N_3373,N_2849);
and U5963 (N_5963,N_3974,N_2833);
and U5964 (N_5964,N_3425,N_2798);
nand U5965 (N_5965,N_3332,N_3870);
nand U5966 (N_5966,N_3786,N_4875);
nand U5967 (N_5967,N_2917,N_4132);
xnor U5968 (N_5968,N_4096,N_2688);
xnor U5969 (N_5969,N_2640,N_3125);
nand U5970 (N_5970,N_3374,N_4617);
nor U5971 (N_5971,N_3385,N_3025);
nand U5972 (N_5972,N_4966,N_4815);
nand U5973 (N_5973,N_2862,N_4924);
or U5974 (N_5974,N_3191,N_4116);
xor U5975 (N_5975,N_2575,N_4631);
and U5976 (N_5976,N_4594,N_4216);
or U5977 (N_5977,N_2765,N_4782);
and U5978 (N_5978,N_4743,N_3516);
nor U5979 (N_5979,N_2637,N_3558);
xor U5980 (N_5980,N_3713,N_3709);
nand U5981 (N_5981,N_3994,N_4685);
and U5982 (N_5982,N_3660,N_3029);
xnor U5983 (N_5983,N_4084,N_4511);
nor U5984 (N_5984,N_3664,N_3168);
nand U5985 (N_5985,N_3327,N_4300);
nor U5986 (N_5986,N_2969,N_2803);
and U5987 (N_5987,N_3123,N_2855);
or U5988 (N_5988,N_3993,N_3120);
nand U5989 (N_5989,N_4758,N_3831);
and U5990 (N_5990,N_3104,N_2557);
xnor U5991 (N_5991,N_2534,N_4175);
or U5992 (N_5992,N_3827,N_4250);
nand U5993 (N_5993,N_4507,N_2840);
xnor U5994 (N_5994,N_2918,N_3876);
or U5995 (N_5995,N_3423,N_3571);
nand U5996 (N_5996,N_2844,N_4655);
nor U5997 (N_5997,N_4167,N_3947);
or U5998 (N_5998,N_3469,N_3412);
and U5999 (N_5999,N_2924,N_4865);
xnor U6000 (N_6000,N_2657,N_3967);
and U6001 (N_6001,N_4632,N_2965);
or U6002 (N_6002,N_3992,N_3382);
xnor U6003 (N_6003,N_4481,N_4723);
nand U6004 (N_6004,N_3391,N_2636);
nor U6005 (N_6005,N_2947,N_3348);
nor U6006 (N_6006,N_3959,N_3941);
and U6007 (N_6007,N_2996,N_2903);
nand U6008 (N_6008,N_4374,N_2998);
nand U6009 (N_6009,N_3539,N_2876);
or U6010 (N_6010,N_4846,N_3634);
xor U6011 (N_6011,N_4445,N_3329);
nand U6012 (N_6012,N_3236,N_4904);
or U6013 (N_6013,N_2652,N_3511);
or U6014 (N_6014,N_3759,N_3489);
and U6015 (N_6015,N_3670,N_2779);
and U6016 (N_6016,N_4013,N_3377);
nor U6017 (N_6017,N_2973,N_3900);
and U6018 (N_6018,N_4045,N_2864);
and U6019 (N_6019,N_3849,N_2936);
and U6020 (N_6020,N_4399,N_3163);
nand U6021 (N_6021,N_4984,N_4896);
or U6022 (N_6022,N_4308,N_2858);
nand U6023 (N_6023,N_2619,N_4635);
nor U6024 (N_6024,N_2773,N_4835);
nand U6025 (N_6025,N_4897,N_4205);
or U6026 (N_6026,N_2626,N_4515);
nand U6027 (N_6027,N_4508,N_2520);
nand U6028 (N_6028,N_3921,N_4376);
nand U6029 (N_6029,N_4649,N_4607);
nor U6030 (N_6030,N_3544,N_3708);
nor U6031 (N_6031,N_3795,N_4852);
and U6032 (N_6032,N_3245,N_4972);
nand U6033 (N_6033,N_3105,N_4118);
nand U6034 (N_6034,N_3161,N_4949);
xor U6035 (N_6035,N_3767,N_3550);
xor U6036 (N_6036,N_2558,N_4218);
nand U6037 (N_6037,N_4440,N_3650);
or U6038 (N_6038,N_4490,N_4988);
nor U6039 (N_6039,N_4119,N_4164);
nor U6040 (N_6040,N_2778,N_3035);
nand U6041 (N_6041,N_2625,N_4059);
nor U6042 (N_6042,N_4847,N_4877);
or U6043 (N_6043,N_4940,N_3340);
xnor U6044 (N_6044,N_4674,N_2935);
or U6045 (N_6045,N_4936,N_4786);
and U6046 (N_6046,N_3931,N_3753);
nor U6047 (N_6047,N_4638,N_2958);
xor U6048 (N_6048,N_2893,N_4855);
and U6049 (N_6049,N_2673,N_2732);
xnor U6050 (N_6050,N_4883,N_2859);
nor U6051 (N_6051,N_2583,N_4489);
nor U6052 (N_6052,N_3746,N_3244);
or U6053 (N_6053,N_4781,N_3200);
and U6054 (N_6054,N_4629,N_2894);
xor U6055 (N_6055,N_3227,N_3923);
and U6056 (N_6056,N_3179,N_3970);
xor U6057 (N_6057,N_3965,N_3402);
or U6058 (N_6058,N_4561,N_4768);
xnor U6059 (N_6059,N_4236,N_4779);
nand U6060 (N_6060,N_3428,N_3088);
nor U6061 (N_6061,N_2905,N_3909);
xnor U6062 (N_6062,N_4359,N_3283);
xnor U6063 (N_6063,N_3766,N_3855);
nor U6064 (N_6064,N_3629,N_4789);
nor U6065 (N_6065,N_3098,N_4868);
xnor U6066 (N_6066,N_4350,N_4524);
nand U6067 (N_6067,N_3762,N_4614);
xor U6068 (N_6068,N_2527,N_4879);
nand U6069 (N_6069,N_2877,N_3804);
or U6070 (N_6070,N_3738,N_3275);
xnor U6071 (N_6071,N_4694,N_3230);
and U6072 (N_6072,N_4814,N_2804);
xnor U6073 (N_6073,N_3676,N_3989);
and U6074 (N_6074,N_3012,N_3050);
and U6075 (N_6075,N_3472,N_3788);
nor U6076 (N_6076,N_4878,N_3846);
or U6077 (N_6077,N_3912,N_2571);
nor U6078 (N_6078,N_4761,N_4361);
and U6079 (N_6079,N_2518,N_3692);
or U6080 (N_6080,N_4335,N_3995);
nor U6081 (N_6081,N_2831,N_3914);
and U6082 (N_6082,N_4699,N_2889);
and U6083 (N_6083,N_3397,N_3939);
and U6084 (N_6084,N_4908,N_4577);
or U6085 (N_6085,N_3154,N_2872);
and U6086 (N_6086,N_4683,N_3118);
xnor U6087 (N_6087,N_3854,N_2580);
nand U6088 (N_6088,N_2514,N_3441);
nand U6089 (N_6089,N_4154,N_4029);
or U6090 (N_6090,N_2682,N_4311);
xnor U6091 (N_6091,N_3654,N_4526);
nand U6092 (N_6092,N_4833,N_2874);
nand U6093 (N_6093,N_4446,N_3246);
xnor U6094 (N_6094,N_4292,N_2850);
nand U6095 (N_6095,N_3950,N_2590);
nand U6096 (N_6096,N_4143,N_3666);
and U6097 (N_6097,N_2537,N_3567);
or U6098 (N_6098,N_3015,N_2997);
and U6099 (N_6099,N_2675,N_2968);
xor U6100 (N_6100,N_4636,N_2762);
and U6101 (N_6101,N_3833,N_3756);
and U6102 (N_6102,N_4447,N_3171);
nand U6103 (N_6103,N_3673,N_4552);
and U6104 (N_6104,N_3475,N_3745);
xor U6105 (N_6105,N_3410,N_3758);
nand U6106 (N_6106,N_3739,N_3319);
xor U6107 (N_6107,N_3790,N_3997);
and U6108 (N_6108,N_2974,N_2838);
and U6109 (N_6109,N_3128,N_4030);
nor U6110 (N_6110,N_3793,N_3874);
and U6111 (N_6111,N_4620,N_4832);
nand U6112 (N_6112,N_4874,N_3979);
and U6113 (N_6113,N_4982,N_3439);
nor U6114 (N_6114,N_3555,N_4863);
nand U6115 (N_6115,N_2822,N_3714);
and U6116 (N_6116,N_4613,N_2854);
or U6117 (N_6117,N_2852,N_2753);
xor U6118 (N_6118,N_4939,N_3443);
nor U6119 (N_6119,N_4213,N_3134);
nand U6120 (N_6120,N_3566,N_4933);
nand U6121 (N_6121,N_4888,N_3109);
nor U6122 (N_6122,N_4576,N_2950);
nor U6123 (N_6123,N_3371,N_3219);
nor U6124 (N_6124,N_4211,N_4190);
and U6125 (N_6125,N_4616,N_4434);
nand U6126 (N_6126,N_3087,N_2885);
or U6127 (N_6127,N_4110,N_3593);
or U6128 (N_6128,N_3898,N_4400);
or U6129 (N_6129,N_2957,N_2805);
or U6130 (N_6130,N_2692,N_3422);
nand U6131 (N_6131,N_3684,N_3616);
nor U6132 (N_6132,N_2660,N_4020);
nor U6133 (N_6133,N_2812,N_2800);
nand U6134 (N_6134,N_4551,N_4974);
nor U6135 (N_6135,N_2898,N_3504);
or U6136 (N_6136,N_4343,N_3805);
nor U6137 (N_6137,N_4762,N_4174);
nor U6138 (N_6138,N_4681,N_3538);
xnor U6139 (N_6139,N_4304,N_3172);
xnor U6140 (N_6140,N_3116,N_4083);
nor U6141 (N_6141,N_4155,N_4147);
xnor U6142 (N_6142,N_4319,N_3049);
nor U6143 (N_6143,N_4973,N_3292);
xor U6144 (N_6144,N_4360,N_3890);
and U6145 (N_6145,N_3590,N_4776);
nor U6146 (N_6146,N_4718,N_2572);
xor U6147 (N_6147,N_2952,N_4765);
nand U6148 (N_6148,N_3250,N_4571);
and U6149 (N_6149,N_3601,N_3376);
xnor U6150 (N_6150,N_2704,N_3512);
or U6151 (N_6151,N_4177,N_3757);
xor U6152 (N_6152,N_3091,N_4839);
xor U6153 (N_6153,N_3813,N_3743);
xor U6154 (N_6154,N_4749,N_4518);
xnor U6155 (N_6155,N_3494,N_4667);
or U6156 (N_6156,N_4071,N_3218);
xnor U6157 (N_6157,N_3131,N_3359);
and U6158 (N_6158,N_4998,N_3878);
nand U6159 (N_6159,N_4529,N_3968);
and U6160 (N_6160,N_4669,N_4889);
and U6161 (N_6161,N_3678,N_4504);
nor U6162 (N_6162,N_4516,N_4166);
nand U6163 (N_6163,N_2581,N_3108);
xor U6164 (N_6164,N_3017,N_4058);
nor U6165 (N_6165,N_4145,N_3457);
nand U6166 (N_6166,N_4398,N_3148);
nor U6167 (N_6167,N_2544,N_3432);
or U6168 (N_6168,N_2999,N_3111);
xnor U6169 (N_6169,N_4891,N_3618);
xnor U6170 (N_6170,N_3252,N_3635);
nor U6171 (N_6171,N_4293,N_3829);
or U6172 (N_6172,N_4248,N_4130);
nor U6173 (N_6173,N_3596,N_3234);
and U6174 (N_6174,N_3817,N_4885);
and U6175 (N_6175,N_3339,N_2770);
and U6176 (N_6176,N_3772,N_3733);
or U6177 (N_6177,N_4323,N_4705);
nand U6178 (N_6178,N_3668,N_2983);
and U6179 (N_6179,N_3731,N_3052);
nand U6180 (N_6180,N_2612,N_3378);
or U6181 (N_6181,N_4693,N_4700);
xor U6182 (N_6182,N_4151,N_4225);
and U6183 (N_6183,N_3517,N_3209);
or U6184 (N_6184,N_2662,N_3403);
or U6185 (N_6185,N_4483,N_4861);
and U6186 (N_6186,N_3548,N_4778);
or U6187 (N_6187,N_3648,N_4642);
nor U6188 (N_6188,N_4644,N_3004);
and U6189 (N_6189,N_3388,N_2503);
nor U6190 (N_6190,N_4430,N_2991);
xor U6191 (N_6191,N_4393,N_4448);
or U6192 (N_6192,N_4208,N_4182);
nand U6193 (N_6193,N_3679,N_4513);
or U6194 (N_6194,N_2981,N_4437);
xor U6195 (N_6195,N_2927,N_2928);
and U6196 (N_6196,N_3559,N_2726);
nand U6197 (N_6197,N_4351,N_3473);
nor U6198 (N_6198,N_4006,N_4530);
or U6199 (N_6199,N_3881,N_3780);
nand U6200 (N_6200,N_3778,N_2646);
xnor U6201 (N_6201,N_4480,N_4141);
nand U6202 (N_6202,N_2942,N_2821);
or U6203 (N_6203,N_4664,N_3728);
and U6204 (N_6204,N_4239,N_4297);
nor U6205 (N_6205,N_4500,N_4028);
and U6206 (N_6206,N_4756,N_3751);
nor U6207 (N_6207,N_3943,N_4769);
and U6208 (N_6208,N_3141,N_3063);
nor U6209 (N_6209,N_3573,N_4317);
nand U6210 (N_6210,N_2842,N_3657);
and U6211 (N_6211,N_4575,N_3691);
nor U6212 (N_6212,N_4337,N_3237);
or U6213 (N_6213,N_4728,N_3470);
or U6214 (N_6214,N_4584,N_4771);
nor U6215 (N_6215,N_4602,N_2736);
and U6216 (N_6216,N_3045,N_4421);
and U6217 (N_6217,N_2593,N_4774);
or U6218 (N_6218,N_2748,N_3180);
and U6219 (N_6219,N_4240,N_3018);
xor U6220 (N_6220,N_4133,N_4487);
or U6221 (N_6221,N_4910,N_4943);
nand U6222 (N_6222,N_4994,N_2954);
xnor U6223 (N_6223,N_3030,N_3696);
nor U6224 (N_6224,N_3822,N_2834);
nor U6225 (N_6225,N_4156,N_3051);
xnor U6226 (N_6226,N_3521,N_3626);
xnor U6227 (N_6227,N_4738,N_3656);
nor U6228 (N_6228,N_3598,N_4354);
and U6229 (N_6229,N_3277,N_4557);
or U6230 (N_6230,N_4089,N_3564);
nand U6231 (N_6231,N_4981,N_4105);
or U6232 (N_6232,N_4333,N_4277);
or U6233 (N_6233,N_4224,N_4419);
nand U6234 (N_6234,N_4793,N_3117);
or U6235 (N_6235,N_2977,N_3588);
xnor U6236 (N_6236,N_2982,N_4144);
nand U6237 (N_6237,N_3427,N_4315);
and U6238 (N_6238,N_2782,N_4601);
nand U6239 (N_6239,N_4072,N_4210);
or U6240 (N_6240,N_4366,N_3838);
nor U6241 (N_6241,N_3178,N_4401);
xnor U6242 (N_6242,N_3092,N_3953);
nor U6243 (N_6243,N_3447,N_4282);
xnor U6244 (N_6244,N_2775,N_2925);
nand U6245 (N_6245,N_3647,N_4542);
nand U6246 (N_6246,N_4592,N_4827);
xnor U6247 (N_6247,N_4970,N_3932);
nor U6248 (N_6248,N_3576,N_3307);
xnor U6249 (N_6249,N_3625,N_3121);
and U6250 (N_6250,N_3203,N_2669);
nor U6251 (N_6251,N_4122,N_2872);
nor U6252 (N_6252,N_3829,N_4701);
xor U6253 (N_6253,N_4545,N_2525);
or U6254 (N_6254,N_2570,N_2711);
and U6255 (N_6255,N_4048,N_4931);
xor U6256 (N_6256,N_3408,N_3331);
and U6257 (N_6257,N_3040,N_4556);
and U6258 (N_6258,N_3881,N_4358);
and U6259 (N_6259,N_2916,N_3759);
nor U6260 (N_6260,N_3880,N_3474);
and U6261 (N_6261,N_3854,N_2895);
nor U6262 (N_6262,N_3318,N_3947);
nand U6263 (N_6263,N_4654,N_2674);
or U6264 (N_6264,N_3385,N_3343);
and U6265 (N_6265,N_3656,N_3110);
nand U6266 (N_6266,N_3554,N_4519);
nand U6267 (N_6267,N_2503,N_3678);
xor U6268 (N_6268,N_3792,N_3118);
or U6269 (N_6269,N_2767,N_2780);
and U6270 (N_6270,N_4073,N_4668);
nor U6271 (N_6271,N_2896,N_2522);
and U6272 (N_6272,N_4694,N_2747);
or U6273 (N_6273,N_4969,N_3769);
or U6274 (N_6274,N_4762,N_2879);
or U6275 (N_6275,N_4773,N_4787);
nor U6276 (N_6276,N_2645,N_4638);
nand U6277 (N_6277,N_3515,N_4411);
and U6278 (N_6278,N_2950,N_2635);
nor U6279 (N_6279,N_3776,N_2651);
and U6280 (N_6280,N_3235,N_3667);
nand U6281 (N_6281,N_3420,N_3624);
or U6282 (N_6282,N_4006,N_2909);
nor U6283 (N_6283,N_2633,N_3397);
xor U6284 (N_6284,N_2736,N_4182);
xor U6285 (N_6285,N_3255,N_3250);
and U6286 (N_6286,N_3697,N_3156);
nand U6287 (N_6287,N_3076,N_3212);
and U6288 (N_6288,N_3860,N_4595);
xor U6289 (N_6289,N_3766,N_4291);
nor U6290 (N_6290,N_2777,N_3283);
nor U6291 (N_6291,N_4279,N_4620);
or U6292 (N_6292,N_2515,N_3703);
nand U6293 (N_6293,N_4050,N_3182);
nand U6294 (N_6294,N_3430,N_4844);
or U6295 (N_6295,N_4258,N_3951);
xnor U6296 (N_6296,N_4848,N_4228);
nand U6297 (N_6297,N_3710,N_2517);
xor U6298 (N_6298,N_4743,N_4120);
or U6299 (N_6299,N_3196,N_2993);
nand U6300 (N_6300,N_2835,N_3247);
and U6301 (N_6301,N_2806,N_2975);
nand U6302 (N_6302,N_4467,N_2686);
or U6303 (N_6303,N_3167,N_3872);
nand U6304 (N_6304,N_3960,N_3105);
and U6305 (N_6305,N_4007,N_2966);
nor U6306 (N_6306,N_3589,N_4791);
nor U6307 (N_6307,N_2765,N_4513);
nor U6308 (N_6308,N_4862,N_3793);
or U6309 (N_6309,N_3863,N_3621);
nand U6310 (N_6310,N_3809,N_2885);
or U6311 (N_6311,N_4347,N_2915);
nor U6312 (N_6312,N_4876,N_2565);
xnor U6313 (N_6313,N_2734,N_4350);
and U6314 (N_6314,N_2514,N_2502);
nand U6315 (N_6315,N_3242,N_2692);
or U6316 (N_6316,N_4947,N_4266);
or U6317 (N_6317,N_4758,N_4731);
xnor U6318 (N_6318,N_4371,N_3154);
nand U6319 (N_6319,N_4050,N_4845);
nand U6320 (N_6320,N_2908,N_3940);
nor U6321 (N_6321,N_2986,N_4248);
nand U6322 (N_6322,N_3749,N_4336);
nor U6323 (N_6323,N_3926,N_4696);
xor U6324 (N_6324,N_3373,N_3294);
nand U6325 (N_6325,N_4935,N_3029);
and U6326 (N_6326,N_3591,N_4993);
nand U6327 (N_6327,N_3940,N_2990);
xnor U6328 (N_6328,N_4556,N_4363);
nor U6329 (N_6329,N_2800,N_3885);
xnor U6330 (N_6330,N_4151,N_4237);
and U6331 (N_6331,N_3443,N_3888);
or U6332 (N_6332,N_3570,N_2898);
xor U6333 (N_6333,N_2643,N_2605);
nor U6334 (N_6334,N_3365,N_3017);
nand U6335 (N_6335,N_4625,N_4852);
nand U6336 (N_6336,N_2500,N_3695);
nor U6337 (N_6337,N_3757,N_4566);
nor U6338 (N_6338,N_3246,N_2791);
or U6339 (N_6339,N_4223,N_4359);
nand U6340 (N_6340,N_4826,N_3159);
xnor U6341 (N_6341,N_3275,N_4182);
or U6342 (N_6342,N_3957,N_2944);
or U6343 (N_6343,N_3018,N_3990);
xnor U6344 (N_6344,N_4488,N_3487);
or U6345 (N_6345,N_4086,N_3774);
nor U6346 (N_6346,N_4731,N_4340);
xnor U6347 (N_6347,N_3099,N_4355);
and U6348 (N_6348,N_4645,N_3778);
nor U6349 (N_6349,N_4955,N_4282);
and U6350 (N_6350,N_4116,N_4976);
nand U6351 (N_6351,N_3413,N_4246);
nand U6352 (N_6352,N_4284,N_2702);
and U6353 (N_6353,N_3346,N_3507);
nor U6354 (N_6354,N_3542,N_2732);
and U6355 (N_6355,N_3170,N_2597);
or U6356 (N_6356,N_4019,N_4283);
xnor U6357 (N_6357,N_3969,N_4499);
and U6358 (N_6358,N_4646,N_4847);
xnor U6359 (N_6359,N_2906,N_4961);
nor U6360 (N_6360,N_4009,N_4489);
or U6361 (N_6361,N_3038,N_2718);
nand U6362 (N_6362,N_4754,N_2551);
xnor U6363 (N_6363,N_3524,N_4326);
or U6364 (N_6364,N_4799,N_2653);
nand U6365 (N_6365,N_2794,N_4352);
nor U6366 (N_6366,N_3597,N_2691);
xor U6367 (N_6367,N_4978,N_3426);
or U6368 (N_6368,N_4267,N_3455);
and U6369 (N_6369,N_4450,N_4538);
or U6370 (N_6370,N_4570,N_3183);
nand U6371 (N_6371,N_2776,N_3431);
xnor U6372 (N_6372,N_2612,N_4460);
or U6373 (N_6373,N_4211,N_2966);
and U6374 (N_6374,N_4473,N_4206);
or U6375 (N_6375,N_3275,N_3608);
xor U6376 (N_6376,N_2503,N_2676);
nand U6377 (N_6377,N_3947,N_2856);
nand U6378 (N_6378,N_4224,N_3892);
and U6379 (N_6379,N_2664,N_3369);
nor U6380 (N_6380,N_4536,N_3959);
xnor U6381 (N_6381,N_3676,N_4030);
nand U6382 (N_6382,N_3694,N_3533);
nand U6383 (N_6383,N_2635,N_4819);
xnor U6384 (N_6384,N_4270,N_4152);
and U6385 (N_6385,N_4193,N_4065);
or U6386 (N_6386,N_4513,N_4112);
and U6387 (N_6387,N_2640,N_3405);
xor U6388 (N_6388,N_4427,N_4299);
xor U6389 (N_6389,N_3697,N_3858);
and U6390 (N_6390,N_4765,N_3899);
xor U6391 (N_6391,N_4313,N_3799);
and U6392 (N_6392,N_2560,N_4598);
and U6393 (N_6393,N_3498,N_3712);
nor U6394 (N_6394,N_3053,N_3391);
and U6395 (N_6395,N_2878,N_3869);
or U6396 (N_6396,N_2958,N_3743);
nor U6397 (N_6397,N_2826,N_3283);
xnor U6398 (N_6398,N_2852,N_4429);
nor U6399 (N_6399,N_2859,N_2911);
nor U6400 (N_6400,N_4877,N_3397);
and U6401 (N_6401,N_2514,N_3740);
nor U6402 (N_6402,N_4625,N_2503);
or U6403 (N_6403,N_4202,N_4947);
and U6404 (N_6404,N_2939,N_4990);
nand U6405 (N_6405,N_3628,N_3813);
nand U6406 (N_6406,N_2690,N_4825);
xor U6407 (N_6407,N_3845,N_2855);
nor U6408 (N_6408,N_4349,N_4405);
and U6409 (N_6409,N_2930,N_3545);
and U6410 (N_6410,N_2552,N_4144);
or U6411 (N_6411,N_4181,N_3502);
or U6412 (N_6412,N_4517,N_3459);
nor U6413 (N_6413,N_3860,N_3186);
xor U6414 (N_6414,N_4483,N_3982);
nor U6415 (N_6415,N_2659,N_4972);
or U6416 (N_6416,N_3413,N_3779);
xor U6417 (N_6417,N_3679,N_3304);
nand U6418 (N_6418,N_3269,N_2752);
or U6419 (N_6419,N_4186,N_3868);
nor U6420 (N_6420,N_4558,N_2661);
nor U6421 (N_6421,N_4843,N_2686);
xnor U6422 (N_6422,N_3522,N_3755);
and U6423 (N_6423,N_2745,N_2743);
xnor U6424 (N_6424,N_2994,N_4839);
xnor U6425 (N_6425,N_3418,N_4573);
or U6426 (N_6426,N_4348,N_2819);
nand U6427 (N_6427,N_4183,N_3408);
xor U6428 (N_6428,N_3786,N_2515);
nand U6429 (N_6429,N_3941,N_3294);
nor U6430 (N_6430,N_3971,N_3198);
nand U6431 (N_6431,N_3367,N_4792);
nor U6432 (N_6432,N_2889,N_3118);
or U6433 (N_6433,N_3166,N_3076);
or U6434 (N_6434,N_3804,N_3586);
nand U6435 (N_6435,N_2790,N_4103);
nor U6436 (N_6436,N_3214,N_4883);
nor U6437 (N_6437,N_3805,N_4945);
nand U6438 (N_6438,N_3481,N_3486);
nand U6439 (N_6439,N_2780,N_3291);
nor U6440 (N_6440,N_3174,N_2624);
nor U6441 (N_6441,N_2761,N_3564);
and U6442 (N_6442,N_3600,N_2909);
xor U6443 (N_6443,N_3264,N_4271);
xor U6444 (N_6444,N_4359,N_4940);
or U6445 (N_6445,N_4764,N_3129);
nand U6446 (N_6446,N_4471,N_3119);
or U6447 (N_6447,N_4646,N_2698);
and U6448 (N_6448,N_4617,N_3768);
xor U6449 (N_6449,N_3895,N_3368);
xnor U6450 (N_6450,N_4607,N_2740);
xnor U6451 (N_6451,N_3840,N_3311);
and U6452 (N_6452,N_4329,N_3677);
nand U6453 (N_6453,N_4236,N_3213);
xnor U6454 (N_6454,N_4829,N_4249);
nor U6455 (N_6455,N_3078,N_3842);
and U6456 (N_6456,N_3994,N_3647);
xnor U6457 (N_6457,N_4703,N_3696);
xnor U6458 (N_6458,N_3075,N_3974);
nand U6459 (N_6459,N_3865,N_3292);
xnor U6460 (N_6460,N_4403,N_4832);
xnor U6461 (N_6461,N_4159,N_3708);
nor U6462 (N_6462,N_3274,N_2804);
xnor U6463 (N_6463,N_4184,N_4756);
or U6464 (N_6464,N_4344,N_4379);
or U6465 (N_6465,N_3352,N_2583);
nand U6466 (N_6466,N_2986,N_3834);
nor U6467 (N_6467,N_2734,N_3308);
and U6468 (N_6468,N_4222,N_3474);
xnor U6469 (N_6469,N_2598,N_3537);
or U6470 (N_6470,N_3030,N_3361);
nor U6471 (N_6471,N_3186,N_4182);
and U6472 (N_6472,N_2693,N_4922);
xor U6473 (N_6473,N_3960,N_3309);
and U6474 (N_6474,N_4176,N_3235);
xnor U6475 (N_6475,N_4180,N_2767);
or U6476 (N_6476,N_4570,N_4353);
xnor U6477 (N_6477,N_3709,N_3087);
and U6478 (N_6478,N_4393,N_3748);
nand U6479 (N_6479,N_3403,N_3056);
nand U6480 (N_6480,N_2825,N_4486);
nor U6481 (N_6481,N_4510,N_4148);
xor U6482 (N_6482,N_4981,N_3754);
and U6483 (N_6483,N_4284,N_3805);
nand U6484 (N_6484,N_4040,N_3409);
and U6485 (N_6485,N_3125,N_2955);
xnor U6486 (N_6486,N_3922,N_3274);
or U6487 (N_6487,N_2535,N_4590);
and U6488 (N_6488,N_4935,N_4584);
and U6489 (N_6489,N_2850,N_3822);
or U6490 (N_6490,N_3881,N_2947);
or U6491 (N_6491,N_4231,N_2834);
and U6492 (N_6492,N_3165,N_4917);
or U6493 (N_6493,N_3985,N_2616);
nand U6494 (N_6494,N_2544,N_3535);
nand U6495 (N_6495,N_3772,N_3591);
nand U6496 (N_6496,N_2633,N_4663);
xnor U6497 (N_6497,N_2946,N_4369);
nand U6498 (N_6498,N_3576,N_3684);
and U6499 (N_6499,N_3318,N_2733);
or U6500 (N_6500,N_3662,N_2578);
xnor U6501 (N_6501,N_3608,N_4375);
nor U6502 (N_6502,N_3057,N_4400);
nand U6503 (N_6503,N_3016,N_3969);
or U6504 (N_6504,N_3752,N_3453);
nor U6505 (N_6505,N_3486,N_2697);
xnor U6506 (N_6506,N_4578,N_2923);
or U6507 (N_6507,N_3724,N_3093);
and U6508 (N_6508,N_3669,N_4187);
xnor U6509 (N_6509,N_3300,N_3164);
nand U6510 (N_6510,N_4210,N_3245);
nand U6511 (N_6511,N_4940,N_3402);
or U6512 (N_6512,N_3214,N_2709);
and U6513 (N_6513,N_3331,N_3866);
or U6514 (N_6514,N_2914,N_4433);
xnor U6515 (N_6515,N_4187,N_3420);
or U6516 (N_6516,N_4128,N_3020);
or U6517 (N_6517,N_2660,N_3937);
or U6518 (N_6518,N_4164,N_2957);
or U6519 (N_6519,N_3849,N_3403);
nor U6520 (N_6520,N_4170,N_2638);
xor U6521 (N_6521,N_4078,N_2680);
or U6522 (N_6522,N_4088,N_3648);
xnor U6523 (N_6523,N_4734,N_2980);
nor U6524 (N_6524,N_3035,N_2813);
and U6525 (N_6525,N_4707,N_3864);
and U6526 (N_6526,N_3522,N_3829);
and U6527 (N_6527,N_4351,N_3297);
nor U6528 (N_6528,N_3546,N_3138);
and U6529 (N_6529,N_4329,N_3592);
xor U6530 (N_6530,N_3542,N_3519);
or U6531 (N_6531,N_3582,N_4735);
and U6532 (N_6532,N_4901,N_3144);
or U6533 (N_6533,N_3013,N_2790);
and U6534 (N_6534,N_4892,N_4847);
nand U6535 (N_6535,N_4011,N_3843);
or U6536 (N_6536,N_3683,N_4026);
or U6537 (N_6537,N_3046,N_3987);
xnor U6538 (N_6538,N_4380,N_3198);
and U6539 (N_6539,N_2782,N_3281);
and U6540 (N_6540,N_2560,N_4451);
nor U6541 (N_6541,N_4108,N_2580);
nand U6542 (N_6542,N_3527,N_3370);
and U6543 (N_6543,N_2663,N_4616);
nor U6544 (N_6544,N_3483,N_3109);
and U6545 (N_6545,N_3797,N_4382);
and U6546 (N_6546,N_4233,N_4375);
nand U6547 (N_6547,N_2541,N_4240);
or U6548 (N_6548,N_2904,N_3259);
nand U6549 (N_6549,N_4001,N_4733);
xor U6550 (N_6550,N_2996,N_2783);
or U6551 (N_6551,N_4377,N_3109);
nand U6552 (N_6552,N_3258,N_3061);
nor U6553 (N_6553,N_3687,N_4410);
xnor U6554 (N_6554,N_3520,N_2602);
or U6555 (N_6555,N_4941,N_3251);
and U6556 (N_6556,N_3481,N_3325);
and U6557 (N_6557,N_4717,N_3910);
xor U6558 (N_6558,N_4294,N_3571);
nand U6559 (N_6559,N_3720,N_3530);
or U6560 (N_6560,N_4631,N_3329);
and U6561 (N_6561,N_4386,N_3803);
nor U6562 (N_6562,N_3202,N_2778);
or U6563 (N_6563,N_4178,N_4280);
and U6564 (N_6564,N_4348,N_4670);
xnor U6565 (N_6565,N_3968,N_4927);
and U6566 (N_6566,N_4921,N_3041);
nand U6567 (N_6567,N_3997,N_4887);
or U6568 (N_6568,N_3235,N_4941);
or U6569 (N_6569,N_3058,N_3224);
and U6570 (N_6570,N_3954,N_3634);
xnor U6571 (N_6571,N_4863,N_4043);
xor U6572 (N_6572,N_4873,N_2632);
and U6573 (N_6573,N_4199,N_2899);
xnor U6574 (N_6574,N_2722,N_3289);
nor U6575 (N_6575,N_4506,N_3953);
nor U6576 (N_6576,N_4315,N_3630);
or U6577 (N_6577,N_4800,N_4070);
nor U6578 (N_6578,N_4605,N_4508);
nor U6579 (N_6579,N_2643,N_4922);
nand U6580 (N_6580,N_3475,N_3305);
xor U6581 (N_6581,N_4955,N_4912);
nand U6582 (N_6582,N_4962,N_4416);
xor U6583 (N_6583,N_4122,N_3318);
nand U6584 (N_6584,N_3141,N_2643);
nand U6585 (N_6585,N_2688,N_2824);
nand U6586 (N_6586,N_3105,N_4952);
or U6587 (N_6587,N_3597,N_3533);
nor U6588 (N_6588,N_4493,N_4702);
and U6589 (N_6589,N_4165,N_4452);
and U6590 (N_6590,N_4943,N_2581);
nand U6591 (N_6591,N_2636,N_4131);
xor U6592 (N_6592,N_4472,N_3818);
or U6593 (N_6593,N_3931,N_4677);
and U6594 (N_6594,N_3822,N_4974);
nand U6595 (N_6595,N_4446,N_2628);
nand U6596 (N_6596,N_3455,N_2982);
nor U6597 (N_6597,N_3065,N_2899);
or U6598 (N_6598,N_2507,N_3458);
and U6599 (N_6599,N_2509,N_4855);
and U6600 (N_6600,N_4137,N_4471);
nor U6601 (N_6601,N_4871,N_4109);
and U6602 (N_6602,N_3688,N_2568);
or U6603 (N_6603,N_4643,N_2963);
or U6604 (N_6604,N_3787,N_4586);
nand U6605 (N_6605,N_4366,N_4210);
or U6606 (N_6606,N_4562,N_3263);
and U6607 (N_6607,N_2523,N_3130);
nor U6608 (N_6608,N_4022,N_3963);
or U6609 (N_6609,N_4765,N_4378);
xnor U6610 (N_6610,N_4914,N_2867);
xnor U6611 (N_6611,N_3782,N_3370);
nand U6612 (N_6612,N_3072,N_3259);
or U6613 (N_6613,N_3608,N_2757);
nand U6614 (N_6614,N_4516,N_4788);
and U6615 (N_6615,N_4229,N_3974);
and U6616 (N_6616,N_3750,N_2699);
and U6617 (N_6617,N_2641,N_3882);
nor U6618 (N_6618,N_3623,N_3655);
nor U6619 (N_6619,N_3983,N_3758);
or U6620 (N_6620,N_4835,N_4774);
and U6621 (N_6621,N_2906,N_2896);
nor U6622 (N_6622,N_2709,N_4499);
nand U6623 (N_6623,N_4086,N_2850);
xnor U6624 (N_6624,N_3036,N_4037);
nor U6625 (N_6625,N_2566,N_3928);
nor U6626 (N_6626,N_3354,N_4585);
xor U6627 (N_6627,N_2992,N_2987);
xnor U6628 (N_6628,N_3488,N_2807);
nor U6629 (N_6629,N_2763,N_3757);
and U6630 (N_6630,N_4815,N_4563);
and U6631 (N_6631,N_4111,N_4116);
nor U6632 (N_6632,N_4632,N_4351);
and U6633 (N_6633,N_2942,N_3656);
nor U6634 (N_6634,N_3154,N_3428);
xnor U6635 (N_6635,N_2592,N_4357);
nand U6636 (N_6636,N_3469,N_3261);
or U6637 (N_6637,N_3024,N_3671);
nor U6638 (N_6638,N_3202,N_2646);
xor U6639 (N_6639,N_2943,N_3040);
nand U6640 (N_6640,N_3128,N_2951);
xnor U6641 (N_6641,N_3236,N_3040);
or U6642 (N_6642,N_4360,N_2619);
or U6643 (N_6643,N_3627,N_4893);
xor U6644 (N_6644,N_4094,N_2960);
or U6645 (N_6645,N_3095,N_2530);
or U6646 (N_6646,N_2517,N_4693);
nand U6647 (N_6647,N_4415,N_4911);
nand U6648 (N_6648,N_4019,N_3689);
or U6649 (N_6649,N_4590,N_4431);
or U6650 (N_6650,N_4651,N_3193);
nor U6651 (N_6651,N_2598,N_4383);
nand U6652 (N_6652,N_3370,N_3506);
xor U6653 (N_6653,N_3763,N_2951);
nor U6654 (N_6654,N_2647,N_3575);
xor U6655 (N_6655,N_4670,N_4683);
nor U6656 (N_6656,N_2685,N_3716);
nand U6657 (N_6657,N_4153,N_3413);
or U6658 (N_6658,N_3602,N_2680);
xnor U6659 (N_6659,N_4084,N_3407);
nand U6660 (N_6660,N_3079,N_2887);
xor U6661 (N_6661,N_2947,N_3913);
or U6662 (N_6662,N_3727,N_2992);
nor U6663 (N_6663,N_4014,N_3009);
nand U6664 (N_6664,N_3206,N_3506);
nand U6665 (N_6665,N_3965,N_4302);
and U6666 (N_6666,N_4489,N_4867);
nor U6667 (N_6667,N_3972,N_2873);
and U6668 (N_6668,N_3924,N_3028);
nand U6669 (N_6669,N_4730,N_4034);
xor U6670 (N_6670,N_4100,N_3590);
or U6671 (N_6671,N_3535,N_4826);
or U6672 (N_6672,N_4078,N_3954);
and U6673 (N_6673,N_4423,N_3097);
and U6674 (N_6674,N_4625,N_4891);
or U6675 (N_6675,N_3226,N_3836);
or U6676 (N_6676,N_3320,N_4239);
nor U6677 (N_6677,N_3919,N_4789);
xor U6678 (N_6678,N_2852,N_3988);
nor U6679 (N_6679,N_2668,N_3907);
nor U6680 (N_6680,N_3323,N_4369);
nor U6681 (N_6681,N_4980,N_2756);
xnor U6682 (N_6682,N_4078,N_4249);
or U6683 (N_6683,N_2714,N_4749);
and U6684 (N_6684,N_4397,N_4259);
xnor U6685 (N_6685,N_2577,N_2507);
nand U6686 (N_6686,N_4078,N_3559);
xnor U6687 (N_6687,N_3856,N_3870);
and U6688 (N_6688,N_4698,N_3263);
nand U6689 (N_6689,N_4204,N_4675);
nand U6690 (N_6690,N_2789,N_2688);
or U6691 (N_6691,N_4576,N_3040);
and U6692 (N_6692,N_4803,N_4072);
and U6693 (N_6693,N_3125,N_3855);
nand U6694 (N_6694,N_2744,N_2947);
or U6695 (N_6695,N_2888,N_3393);
nor U6696 (N_6696,N_2833,N_4358);
or U6697 (N_6697,N_3038,N_4467);
nand U6698 (N_6698,N_4771,N_3683);
nor U6699 (N_6699,N_4555,N_2986);
nand U6700 (N_6700,N_2836,N_4589);
or U6701 (N_6701,N_2581,N_3655);
nor U6702 (N_6702,N_4383,N_4750);
nor U6703 (N_6703,N_3499,N_3672);
nor U6704 (N_6704,N_3918,N_3621);
nor U6705 (N_6705,N_3081,N_3403);
nor U6706 (N_6706,N_4703,N_2900);
and U6707 (N_6707,N_4540,N_4957);
and U6708 (N_6708,N_3465,N_4443);
xnor U6709 (N_6709,N_3359,N_4913);
nor U6710 (N_6710,N_3841,N_2731);
or U6711 (N_6711,N_4983,N_3950);
or U6712 (N_6712,N_4224,N_3471);
and U6713 (N_6713,N_3376,N_4716);
and U6714 (N_6714,N_4992,N_2508);
xnor U6715 (N_6715,N_3832,N_3011);
or U6716 (N_6716,N_3091,N_3530);
nand U6717 (N_6717,N_3028,N_2632);
nor U6718 (N_6718,N_4553,N_2869);
xor U6719 (N_6719,N_4627,N_4353);
xor U6720 (N_6720,N_3726,N_4548);
nor U6721 (N_6721,N_4808,N_3297);
and U6722 (N_6722,N_3733,N_4796);
nand U6723 (N_6723,N_3500,N_2870);
or U6724 (N_6724,N_4194,N_4619);
and U6725 (N_6725,N_3908,N_2943);
xor U6726 (N_6726,N_3625,N_3110);
and U6727 (N_6727,N_3086,N_3343);
and U6728 (N_6728,N_4210,N_3608);
or U6729 (N_6729,N_3368,N_4305);
xnor U6730 (N_6730,N_3636,N_3353);
nand U6731 (N_6731,N_3234,N_4825);
and U6732 (N_6732,N_2543,N_4531);
xnor U6733 (N_6733,N_3677,N_4743);
xnor U6734 (N_6734,N_3185,N_4041);
nand U6735 (N_6735,N_4790,N_4197);
nor U6736 (N_6736,N_3599,N_3453);
nand U6737 (N_6737,N_4064,N_3061);
xor U6738 (N_6738,N_3163,N_3015);
or U6739 (N_6739,N_2916,N_3889);
and U6740 (N_6740,N_3685,N_2948);
xnor U6741 (N_6741,N_2538,N_3796);
nand U6742 (N_6742,N_4015,N_4384);
or U6743 (N_6743,N_2981,N_3215);
and U6744 (N_6744,N_2788,N_3132);
and U6745 (N_6745,N_3926,N_3463);
xor U6746 (N_6746,N_3611,N_4207);
and U6747 (N_6747,N_3255,N_4824);
nand U6748 (N_6748,N_3988,N_2795);
nand U6749 (N_6749,N_3125,N_3772);
nand U6750 (N_6750,N_4983,N_4575);
nand U6751 (N_6751,N_2986,N_4954);
and U6752 (N_6752,N_4287,N_4062);
and U6753 (N_6753,N_3339,N_4266);
nor U6754 (N_6754,N_3540,N_2647);
or U6755 (N_6755,N_4150,N_2702);
or U6756 (N_6756,N_2863,N_2729);
xnor U6757 (N_6757,N_4396,N_3079);
xnor U6758 (N_6758,N_4229,N_3041);
xnor U6759 (N_6759,N_3200,N_3676);
xnor U6760 (N_6760,N_3081,N_2583);
xnor U6761 (N_6761,N_3160,N_4523);
and U6762 (N_6762,N_2996,N_2734);
nor U6763 (N_6763,N_4053,N_4458);
xor U6764 (N_6764,N_3338,N_3255);
nand U6765 (N_6765,N_2741,N_3838);
and U6766 (N_6766,N_3650,N_3431);
and U6767 (N_6767,N_4190,N_4685);
nand U6768 (N_6768,N_4812,N_4106);
nand U6769 (N_6769,N_2660,N_3699);
xnor U6770 (N_6770,N_3126,N_2686);
nor U6771 (N_6771,N_4851,N_4869);
nor U6772 (N_6772,N_3109,N_3084);
or U6773 (N_6773,N_2696,N_4222);
or U6774 (N_6774,N_3614,N_4282);
or U6775 (N_6775,N_3559,N_3076);
nand U6776 (N_6776,N_3383,N_4316);
nand U6777 (N_6777,N_3209,N_4462);
or U6778 (N_6778,N_4016,N_3985);
and U6779 (N_6779,N_3153,N_2594);
and U6780 (N_6780,N_3036,N_2975);
xor U6781 (N_6781,N_4112,N_4862);
nand U6782 (N_6782,N_3603,N_3253);
nor U6783 (N_6783,N_3620,N_4500);
nand U6784 (N_6784,N_4266,N_3952);
xor U6785 (N_6785,N_4151,N_4967);
nand U6786 (N_6786,N_3346,N_3120);
xor U6787 (N_6787,N_4172,N_3263);
nor U6788 (N_6788,N_2590,N_4233);
nor U6789 (N_6789,N_4408,N_3904);
or U6790 (N_6790,N_2781,N_4872);
and U6791 (N_6791,N_4003,N_2900);
nor U6792 (N_6792,N_3289,N_4047);
or U6793 (N_6793,N_2713,N_4735);
and U6794 (N_6794,N_4203,N_2680);
nor U6795 (N_6795,N_3454,N_3351);
and U6796 (N_6796,N_3278,N_2805);
nand U6797 (N_6797,N_3414,N_3609);
nor U6798 (N_6798,N_3589,N_3055);
and U6799 (N_6799,N_3432,N_3834);
nor U6800 (N_6800,N_2983,N_3636);
nor U6801 (N_6801,N_3651,N_4973);
nor U6802 (N_6802,N_3791,N_3576);
and U6803 (N_6803,N_4144,N_3715);
nand U6804 (N_6804,N_2699,N_2972);
nand U6805 (N_6805,N_3247,N_3761);
nand U6806 (N_6806,N_4849,N_4438);
and U6807 (N_6807,N_4981,N_4349);
xnor U6808 (N_6808,N_4944,N_2969);
or U6809 (N_6809,N_3805,N_2993);
xor U6810 (N_6810,N_4703,N_3201);
and U6811 (N_6811,N_3225,N_3442);
nor U6812 (N_6812,N_4591,N_2571);
nand U6813 (N_6813,N_4935,N_4833);
and U6814 (N_6814,N_2790,N_3322);
or U6815 (N_6815,N_4700,N_3806);
or U6816 (N_6816,N_3249,N_3626);
nand U6817 (N_6817,N_4327,N_2954);
nand U6818 (N_6818,N_4939,N_2854);
or U6819 (N_6819,N_2551,N_4852);
and U6820 (N_6820,N_2558,N_3073);
nand U6821 (N_6821,N_3687,N_4098);
xor U6822 (N_6822,N_4837,N_2839);
and U6823 (N_6823,N_3673,N_4753);
xor U6824 (N_6824,N_3703,N_4316);
and U6825 (N_6825,N_2868,N_3380);
nor U6826 (N_6826,N_4294,N_3713);
xor U6827 (N_6827,N_2762,N_2618);
xnor U6828 (N_6828,N_3817,N_2601);
nor U6829 (N_6829,N_2969,N_2887);
and U6830 (N_6830,N_3653,N_3229);
nand U6831 (N_6831,N_3790,N_4159);
nor U6832 (N_6832,N_4670,N_3014);
or U6833 (N_6833,N_3965,N_2783);
xor U6834 (N_6834,N_3771,N_4031);
and U6835 (N_6835,N_3454,N_4667);
xor U6836 (N_6836,N_4200,N_3811);
and U6837 (N_6837,N_4315,N_3028);
xor U6838 (N_6838,N_4839,N_2581);
nor U6839 (N_6839,N_4762,N_2505);
nor U6840 (N_6840,N_3831,N_3355);
or U6841 (N_6841,N_3435,N_4962);
xnor U6842 (N_6842,N_3281,N_4122);
or U6843 (N_6843,N_3634,N_4206);
or U6844 (N_6844,N_3534,N_3368);
nand U6845 (N_6845,N_2946,N_3821);
xor U6846 (N_6846,N_3204,N_3621);
or U6847 (N_6847,N_3309,N_2610);
xnor U6848 (N_6848,N_4274,N_4067);
or U6849 (N_6849,N_4926,N_3137);
nand U6850 (N_6850,N_4839,N_3693);
xnor U6851 (N_6851,N_4424,N_2862);
nor U6852 (N_6852,N_2771,N_2903);
nand U6853 (N_6853,N_2543,N_4544);
or U6854 (N_6854,N_3915,N_4499);
nor U6855 (N_6855,N_4806,N_3516);
xor U6856 (N_6856,N_3259,N_3442);
nand U6857 (N_6857,N_4967,N_3865);
and U6858 (N_6858,N_2925,N_2869);
and U6859 (N_6859,N_3913,N_4912);
nor U6860 (N_6860,N_3951,N_3227);
nor U6861 (N_6861,N_2706,N_2602);
or U6862 (N_6862,N_4798,N_2724);
nor U6863 (N_6863,N_4146,N_4775);
nand U6864 (N_6864,N_2712,N_3779);
or U6865 (N_6865,N_2614,N_4278);
and U6866 (N_6866,N_4341,N_3893);
and U6867 (N_6867,N_2696,N_4285);
and U6868 (N_6868,N_4647,N_4926);
xnor U6869 (N_6869,N_4050,N_4914);
nand U6870 (N_6870,N_4101,N_2678);
nand U6871 (N_6871,N_3659,N_3963);
or U6872 (N_6872,N_3507,N_3588);
nand U6873 (N_6873,N_2565,N_3731);
and U6874 (N_6874,N_3989,N_2649);
or U6875 (N_6875,N_4927,N_2636);
xnor U6876 (N_6876,N_3321,N_4972);
or U6877 (N_6877,N_3469,N_4869);
nor U6878 (N_6878,N_2620,N_2523);
nand U6879 (N_6879,N_2512,N_3819);
nor U6880 (N_6880,N_4823,N_3202);
and U6881 (N_6881,N_2902,N_3372);
or U6882 (N_6882,N_3941,N_2958);
nand U6883 (N_6883,N_4910,N_3343);
and U6884 (N_6884,N_2884,N_2712);
xnor U6885 (N_6885,N_3419,N_4497);
or U6886 (N_6886,N_4067,N_2879);
or U6887 (N_6887,N_4804,N_3383);
xor U6888 (N_6888,N_3443,N_4795);
nor U6889 (N_6889,N_4428,N_3458);
or U6890 (N_6890,N_3987,N_4135);
nand U6891 (N_6891,N_4207,N_3957);
nor U6892 (N_6892,N_3504,N_3389);
xor U6893 (N_6893,N_4312,N_4402);
xor U6894 (N_6894,N_4689,N_2511);
nor U6895 (N_6895,N_4728,N_2646);
nand U6896 (N_6896,N_3843,N_3222);
nand U6897 (N_6897,N_4120,N_4983);
xnor U6898 (N_6898,N_4703,N_4260);
and U6899 (N_6899,N_3411,N_4907);
nor U6900 (N_6900,N_4214,N_4835);
nand U6901 (N_6901,N_3376,N_3831);
or U6902 (N_6902,N_3315,N_4830);
and U6903 (N_6903,N_4255,N_4105);
and U6904 (N_6904,N_4482,N_2724);
nand U6905 (N_6905,N_2608,N_3815);
and U6906 (N_6906,N_3256,N_3561);
nor U6907 (N_6907,N_3720,N_2979);
nor U6908 (N_6908,N_4806,N_2929);
and U6909 (N_6909,N_3079,N_4619);
nand U6910 (N_6910,N_2733,N_2646);
nand U6911 (N_6911,N_4862,N_3154);
nand U6912 (N_6912,N_4076,N_4930);
nor U6913 (N_6913,N_3617,N_3942);
and U6914 (N_6914,N_4955,N_2746);
nand U6915 (N_6915,N_3123,N_4736);
nand U6916 (N_6916,N_3773,N_2616);
or U6917 (N_6917,N_3692,N_2596);
or U6918 (N_6918,N_4869,N_4265);
xor U6919 (N_6919,N_4881,N_4516);
and U6920 (N_6920,N_2850,N_4546);
nor U6921 (N_6921,N_3339,N_4595);
or U6922 (N_6922,N_4239,N_4491);
or U6923 (N_6923,N_3765,N_4483);
or U6924 (N_6924,N_2523,N_4455);
or U6925 (N_6925,N_2741,N_3593);
nor U6926 (N_6926,N_3808,N_2934);
and U6927 (N_6927,N_3614,N_4562);
xnor U6928 (N_6928,N_4476,N_3601);
and U6929 (N_6929,N_4187,N_3865);
nand U6930 (N_6930,N_3492,N_3324);
and U6931 (N_6931,N_4089,N_3208);
and U6932 (N_6932,N_2933,N_2859);
xor U6933 (N_6933,N_3028,N_3303);
or U6934 (N_6934,N_4420,N_2929);
nand U6935 (N_6935,N_3537,N_4936);
or U6936 (N_6936,N_3904,N_2934);
or U6937 (N_6937,N_4239,N_4353);
or U6938 (N_6938,N_4528,N_3462);
xor U6939 (N_6939,N_3980,N_3125);
or U6940 (N_6940,N_3069,N_3192);
nand U6941 (N_6941,N_3022,N_4698);
xor U6942 (N_6942,N_4962,N_3783);
xnor U6943 (N_6943,N_4039,N_2512);
nand U6944 (N_6944,N_3865,N_2545);
or U6945 (N_6945,N_3854,N_3299);
or U6946 (N_6946,N_3779,N_3974);
nand U6947 (N_6947,N_2644,N_4796);
xor U6948 (N_6948,N_2916,N_3379);
and U6949 (N_6949,N_3775,N_3023);
or U6950 (N_6950,N_4041,N_4559);
and U6951 (N_6951,N_3301,N_4767);
and U6952 (N_6952,N_3110,N_2825);
xnor U6953 (N_6953,N_2752,N_4269);
nor U6954 (N_6954,N_3214,N_3546);
nor U6955 (N_6955,N_3366,N_2662);
and U6956 (N_6956,N_4871,N_3526);
or U6957 (N_6957,N_4341,N_3029);
nor U6958 (N_6958,N_4366,N_4679);
and U6959 (N_6959,N_3560,N_3989);
nor U6960 (N_6960,N_3780,N_4855);
or U6961 (N_6961,N_4946,N_3932);
and U6962 (N_6962,N_4727,N_2820);
nand U6963 (N_6963,N_4659,N_3432);
nor U6964 (N_6964,N_2616,N_4181);
nand U6965 (N_6965,N_4487,N_3589);
or U6966 (N_6966,N_2746,N_4635);
nand U6967 (N_6967,N_3245,N_3893);
nand U6968 (N_6968,N_3297,N_4926);
or U6969 (N_6969,N_3464,N_4796);
or U6970 (N_6970,N_4703,N_4121);
nor U6971 (N_6971,N_4459,N_3259);
nor U6972 (N_6972,N_2502,N_3860);
nand U6973 (N_6973,N_4442,N_4660);
or U6974 (N_6974,N_3135,N_2897);
or U6975 (N_6975,N_3268,N_3115);
or U6976 (N_6976,N_2951,N_2994);
nor U6977 (N_6977,N_4821,N_4382);
nand U6978 (N_6978,N_4524,N_4869);
or U6979 (N_6979,N_3282,N_4219);
xnor U6980 (N_6980,N_4745,N_4822);
or U6981 (N_6981,N_3588,N_3409);
or U6982 (N_6982,N_3490,N_4338);
xnor U6983 (N_6983,N_3099,N_4559);
and U6984 (N_6984,N_4423,N_3603);
nor U6985 (N_6985,N_4905,N_4922);
nor U6986 (N_6986,N_3052,N_2535);
xnor U6987 (N_6987,N_4867,N_4019);
and U6988 (N_6988,N_3138,N_3510);
nor U6989 (N_6989,N_3396,N_2734);
or U6990 (N_6990,N_4612,N_3267);
nand U6991 (N_6991,N_4310,N_2573);
nor U6992 (N_6992,N_4642,N_3740);
xor U6993 (N_6993,N_3279,N_4708);
nand U6994 (N_6994,N_4500,N_3753);
nor U6995 (N_6995,N_2551,N_3576);
and U6996 (N_6996,N_4487,N_2769);
or U6997 (N_6997,N_2877,N_3450);
nand U6998 (N_6998,N_3367,N_3565);
and U6999 (N_6999,N_3641,N_4252);
nor U7000 (N_7000,N_4106,N_3574);
and U7001 (N_7001,N_3381,N_2633);
or U7002 (N_7002,N_3466,N_3110);
nand U7003 (N_7003,N_4447,N_3961);
nand U7004 (N_7004,N_4586,N_3470);
nor U7005 (N_7005,N_4486,N_4101);
nand U7006 (N_7006,N_2982,N_3101);
nor U7007 (N_7007,N_2703,N_3416);
or U7008 (N_7008,N_4712,N_4249);
nor U7009 (N_7009,N_3393,N_4062);
and U7010 (N_7010,N_3631,N_3664);
nand U7011 (N_7011,N_4622,N_3696);
xor U7012 (N_7012,N_4763,N_3034);
nand U7013 (N_7013,N_2970,N_3711);
xnor U7014 (N_7014,N_3201,N_2656);
xor U7015 (N_7015,N_3734,N_3383);
nand U7016 (N_7016,N_2885,N_4312);
nor U7017 (N_7017,N_4100,N_2963);
nand U7018 (N_7018,N_2899,N_3010);
and U7019 (N_7019,N_2898,N_4165);
and U7020 (N_7020,N_3688,N_3970);
xor U7021 (N_7021,N_3454,N_3978);
nand U7022 (N_7022,N_4105,N_4619);
xor U7023 (N_7023,N_3600,N_4814);
xnor U7024 (N_7024,N_4086,N_4725);
xnor U7025 (N_7025,N_3368,N_2970);
xor U7026 (N_7026,N_4196,N_2552);
or U7027 (N_7027,N_4088,N_4543);
or U7028 (N_7028,N_3526,N_4886);
nor U7029 (N_7029,N_4412,N_4049);
and U7030 (N_7030,N_4299,N_3348);
and U7031 (N_7031,N_3065,N_3356);
and U7032 (N_7032,N_4049,N_2586);
or U7033 (N_7033,N_3411,N_3225);
nand U7034 (N_7034,N_4824,N_3026);
or U7035 (N_7035,N_4861,N_2584);
and U7036 (N_7036,N_4263,N_3968);
nand U7037 (N_7037,N_3246,N_2830);
and U7038 (N_7038,N_2654,N_4132);
nand U7039 (N_7039,N_3743,N_3811);
or U7040 (N_7040,N_4507,N_4594);
xnor U7041 (N_7041,N_2943,N_4337);
nor U7042 (N_7042,N_3019,N_2971);
nand U7043 (N_7043,N_4130,N_2774);
nor U7044 (N_7044,N_3987,N_3843);
and U7045 (N_7045,N_2571,N_4251);
nand U7046 (N_7046,N_4340,N_3964);
or U7047 (N_7047,N_3865,N_3066);
and U7048 (N_7048,N_4621,N_4756);
and U7049 (N_7049,N_2752,N_3576);
or U7050 (N_7050,N_4404,N_4021);
and U7051 (N_7051,N_3888,N_4847);
nor U7052 (N_7052,N_3392,N_3462);
and U7053 (N_7053,N_3941,N_3243);
xnor U7054 (N_7054,N_4643,N_3157);
nor U7055 (N_7055,N_4215,N_3337);
nand U7056 (N_7056,N_3199,N_4637);
nor U7057 (N_7057,N_3973,N_2953);
xnor U7058 (N_7058,N_4122,N_4628);
nand U7059 (N_7059,N_3138,N_2750);
nor U7060 (N_7060,N_2801,N_3400);
nand U7061 (N_7061,N_3004,N_2930);
nor U7062 (N_7062,N_3932,N_4723);
xor U7063 (N_7063,N_3946,N_3794);
and U7064 (N_7064,N_2932,N_3135);
or U7065 (N_7065,N_4867,N_2959);
nand U7066 (N_7066,N_3700,N_2980);
and U7067 (N_7067,N_3496,N_4198);
or U7068 (N_7068,N_2597,N_2939);
xor U7069 (N_7069,N_4186,N_4944);
or U7070 (N_7070,N_3449,N_3575);
xor U7071 (N_7071,N_4296,N_3742);
and U7072 (N_7072,N_3259,N_3476);
xnor U7073 (N_7073,N_4912,N_4796);
nor U7074 (N_7074,N_4410,N_2973);
nand U7075 (N_7075,N_4051,N_4774);
xnor U7076 (N_7076,N_3965,N_3952);
xnor U7077 (N_7077,N_4277,N_2523);
and U7078 (N_7078,N_3928,N_3709);
or U7079 (N_7079,N_2660,N_4697);
or U7080 (N_7080,N_2976,N_3185);
or U7081 (N_7081,N_3837,N_3756);
or U7082 (N_7082,N_2751,N_2730);
and U7083 (N_7083,N_3150,N_3448);
nand U7084 (N_7084,N_3233,N_3070);
xor U7085 (N_7085,N_4709,N_2763);
and U7086 (N_7086,N_4756,N_4793);
nor U7087 (N_7087,N_2860,N_2851);
and U7088 (N_7088,N_2985,N_2752);
nor U7089 (N_7089,N_4700,N_3135);
xor U7090 (N_7090,N_4450,N_3453);
and U7091 (N_7091,N_4123,N_2840);
xor U7092 (N_7092,N_3341,N_4913);
xnor U7093 (N_7093,N_3495,N_3112);
nor U7094 (N_7094,N_3127,N_3665);
xor U7095 (N_7095,N_4319,N_3551);
nand U7096 (N_7096,N_4792,N_3780);
and U7097 (N_7097,N_3242,N_4512);
or U7098 (N_7098,N_3521,N_3122);
nand U7099 (N_7099,N_2937,N_4247);
and U7100 (N_7100,N_4340,N_3506);
xnor U7101 (N_7101,N_3026,N_3627);
nor U7102 (N_7102,N_3313,N_3563);
nand U7103 (N_7103,N_2774,N_3592);
or U7104 (N_7104,N_2949,N_4385);
xnor U7105 (N_7105,N_3002,N_3062);
or U7106 (N_7106,N_2732,N_4787);
or U7107 (N_7107,N_3927,N_4019);
nand U7108 (N_7108,N_4902,N_3483);
and U7109 (N_7109,N_3568,N_2632);
xnor U7110 (N_7110,N_4904,N_3611);
nand U7111 (N_7111,N_3078,N_3310);
or U7112 (N_7112,N_4428,N_3918);
xor U7113 (N_7113,N_3258,N_4439);
or U7114 (N_7114,N_3198,N_4654);
nor U7115 (N_7115,N_3675,N_4835);
nand U7116 (N_7116,N_4464,N_2948);
or U7117 (N_7117,N_3995,N_2755);
or U7118 (N_7118,N_4119,N_2864);
nor U7119 (N_7119,N_2830,N_2889);
and U7120 (N_7120,N_2530,N_2855);
nand U7121 (N_7121,N_4743,N_3243);
or U7122 (N_7122,N_3220,N_3578);
nor U7123 (N_7123,N_3730,N_2779);
xor U7124 (N_7124,N_3021,N_2976);
and U7125 (N_7125,N_4104,N_3148);
xnor U7126 (N_7126,N_3621,N_3802);
nor U7127 (N_7127,N_3829,N_3651);
xnor U7128 (N_7128,N_4563,N_2520);
nand U7129 (N_7129,N_3053,N_3092);
nand U7130 (N_7130,N_4843,N_2501);
and U7131 (N_7131,N_4459,N_4058);
nor U7132 (N_7132,N_2627,N_3643);
and U7133 (N_7133,N_3170,N_2567);
nand U7134 (N_7134,N_4653,N_2605);
and U7135 (N_7135,N_4030,N_3656);
or U7136 (N_7136,N_4081,N_3983);
nor U7137 (N_7137,N_3931,N_3373);
nor U7138 (N_7138,N_4445,N_3565);
nand U7139 (N_7139,N_4624,N_4167);
xnor U7140 (N_7140,N_2833,N_2990);
nand U7141 (N_7141,N_2989,N_3866);
and U7142 (N_7142,N_2832,N_4083);
or U7143 (N_7143,N_4129,N_2830);
nor U7144 (N_7144,N_2726,N_2677);
or U7145 (N_7145,N_4572,N_3596);
and U7146 (N_7146,N_4002,N_4214);
xor U7147 (N_7147,N_2594,N_2572);
xnor U7148 (N_7148,N_4186,N_3261);
xnor U7149 (N_7149,N_3494,N_3962);
nor U7150 (N_7150,N_3207,N_2928);
and U7151 (N_7151,N_4782,N_3266);
nor U7152 (N_7152,N_4161,N_3892);
and U7153 (N_7153,N_4875,N_3026);
and U7154 (N_7154,N_4003,N_2708);
xor U7155 (N_7155,N_3890,N_2878);
nor U7156 (N_7156,N_2829,N_4800);
or U7157 (N_7157,N_3033,N_2711);
xnor U7158 (N_7158,N_4438,N_4840);
or U7159 (N_7159,N_3440,N_4802);
nor U7160 (N_7160,N_3273,N_3859);
and U7161 (N_7161,N_3024,N_2946);
xor U7162 (N_7162,N_4650,N_3251);
nand U7163 (N_7163,N_2853,N_4307);
nor U7164 (N_7164,N_3171,N_3564);
xnor U7165 (N_7165,N_4324,N_3768);
or U7166 (N_7166,N_2800,N_4771);
xor U7167 (N_7167,N_3168,N_2591);
nor U7168 (N_7168,N_3508,N_3332);
nor U7169 (N_7169,N_3564,N_4735);
nand U7170 (N_7170,N_4034,N_3999);
nand U7171 (N_7171,N_3129,N_3313);
or U7172 (N_7172,N_4409,N_3192);
and U7173 (N_7173,N_2754,N_3626);
nor U7174 (N_7174,N_4647,N_3558);
and U7175 (N_7175,N_4211,N_3820);
nor U7176 (N_7176,N_4954,N_4407);
nand U7177 (N_7177,N_4837,N_4676);
nor U7178 (N_7178,N_2766,N_4092);
and U7179 (N_7179,N_2992,N_2697);
or U7180 (N_7180,N_3750,N_3109);
xnor U7181 (N_7181,N_4355,N_4538);
nor U7182 (N_7182,N_3228,N_3989);
xor U7183 (N_7183,N_2525,N_3443);
xor U7184 (N_7184,N_4718,N_4857);
and U7185 (N_7185,N_4885,N_4343);
and U7186 (N_7186,N_3551,N_3346);
nand U7187 (N_7187,N_4848,N_3643);
and U7188 (N_7188,N_2967,N_2984);
and U7189 (N_7189,N_4808,N_4367);
and U7190 (N_7190,N_4040,N_3936);
xnor U7191 (N_7191,N_3124,N_3939);
nor U7192 (N_7192,N_3887,N_3822);
xor U7193 (N_7193,N_3803,N_3815);
xor U7194 (N_7194,N_4730,N_3966);
nor U7195 (N_7195,N_4832,N_3968);
nand U7196 (N_7196,N_3639,N_3508);
or U7197 (N_7197,N_4711,N_4338);
xor U7198 (N_7198,N_2928,N_3111);
and U7199 (N_7199,N_3786,N_3374);
nor U7200 (N_7200,N_4349,N_3080);
nor U7201 (N_7201,N_3918,N_4643);
or U7202 (N_7202,N_3824,N_3427);
xnor U7203 (N_7203,N_4380,N_3379);
or U7204 (N_7204,N_2643,N_4264);
xor U7205 (N_7205,N_2986,N_3744);
or U7206 (N_7206,N_4695,N_4569);
nor U7207 (N_7207,N_2870,N_3642);
xor U7208 (N_7208,N_3531,N_3215);
nand U7209 (N_7209,N_3056,N_3873);
xor U7210 (N_7210,N_2507,N_2928);
nor U7211 (N_7211,N_4895,N_2854);
nor U7212 (N_7212,N_3566,N_3486);
and U7213 (N_7213,N_4619,N_2907);
nand U7214 (N_7214,N_4316,N_2817);
or U7215 (N_7215,N_3000,N_4896);
xnor U7216 (N_7216,N_3263,N_4314);
nor U7217 (N_7217,N_4876,N_4789);
nor U7218 (N_7218,N_3718,N_3827);
and U7219 (N_7219,N_4699,N_4885);
nand U7220 (N_7220,N_3121,N_3923);
nand U7221 (N_7221,N_4020,N_3293);
nor U7222 (N_7222,N_2790,N_2906);
nand U7223 (N_7223,N_3052,N_3851);
and U7224 (N_7224,N_3157,N_4215);
nand U7225 (N_7225,N_4768,N_2861);
nor U7226 (N_7226,N_4646,N_4979);
and U7227 (N_7227,N_2531,N_4902);
nand U7228 (N_7228,N_4419,N_3184);
nand U7229 (N_7229,N_2731,N_3672);
or U7230 (N_7230,N_3219,N_4502);
nor U7231 (N_7231,N_3625,N_2772);
or U7232 (N_7232,N_4489,N_4290);
xor U7233 (N_7233,N_4725,N_3977);
xor U7234 (N_7234,N_4648,N_4733);
nand U7235 (N_7235,N_4164,N_2582);
nor U7236 (N_7236,N_3893,N_2526);
xnor U7237 (N_7237,N_3808,N_4233);
or U7238 (N_7238,N_4931,N_3543);
or U7239 (N_7239,N_4301,N_3060);
nand U7240 (N_7240,N_3382,N_4149);
or U7241 (N_7241,N_4757,N_3214);
xnor U7242 (N_7242,N_3035,N_4851);
or U7243 (N_7243,N_4838,N_3048);
xor U7244 (N_7244,N_3945,N_2919);
and U7245 (N_7245,N_2950,N_3378);
nand U7246 (N_7246,N_4260,N_3772);
and U7247 (N_7247,N_3669,N_2784);
nor U7248 (N_7248,N_2800,N_3243);
and U7249 (N_7249,N_2951,N_3253);
nand U7250 (N_7250,N_2835,N_4034);
or U7251 (N_7251,N_3542,N_3241);
xnor U7252 (N_7252,N_4286,N_4920);
nor U7253 (N_7253,N_3203,N_4334);
nor U7254 (N_7254,N_3989,N_3982);
nor U7255 (N_7255,N_3455,N_3387);
nand U7256 (N_7256,N_3220,N_4722);
xor U7257 (N_7257,N_3309,N_4441);
or U7258 (N_7258,N_3718,N_2543);
and U7259 (N_7259,N_4469,N_3755);
nor U7260 (N_7260,N_4751,N_2692);
and U7261 (N_7261,N_4902,N_3318);
xor U7262 (N_7262,N_3245,N_3816);
or U7263 (N_7263,N_2631,N_3686);
nand U7264 (N_7264,N_4700,N_4605);
or U7265 (N_7265,N_2974,N_3146);
or U7266 (N_7266,N_3741,N_4370);
nor U7267 (N_7267,N_3879,N_4696);
nand U7268 (N_7268,N_4929,N_3277);
and U7269 (N_7269,N_3904,N_3215);
nor U7270 (N_7270,N_3893,N_4153);
and U7271 (N_7271,N_3206,N_4234);
nand U7272 (N_7272,N_3933,N_4571);
nand U7273 (N_7273,N_3712,N_4108);
or U7274 (N_7274,N_2864,N_3508);
nand U7275 (N_7275,N_4035,N_3452);
or U7276 (N_7276,N_4689,N_4571);
and U7277 (N_7277,N_3236,N_4484);
nand U7278 (N_7278,N_4385,N_2937);
xnor U7279 (N_7279,N_3801,N_3646);
nor U7280 (N_7280,N_2843,N_4400);
or U7281 (N_7281,N_3360,N_3218);
xnor U7282 (N_7282,N_3567,N_3511);
and U7283 (N_7283,N_2687,N_4526);
or U7284 (N_7284,N_4624,N_4456);
or U7285 (N_7285,N_4957,N_3353);
nor U7286 (N_7286,N_2609,N_3909);
xnor U7287 (N_7287,N_4670,N_3556);
nor U7288 (N_7288,N_2737,N_2925);
nor U7289 (N_7289,N_2830,N_3184);
xor U7290 (N_7290,N_4176,N_4680);
nand U7291 (N_7291,N_3080,N_4759);
nor U7292 (N_7292,N_3258,N_3126);
xnor U7293 (N_7293,N_2548,N_4017);
or U7294 (N_7294,N_4278,N_3800);
xor U7295 (N_7295,N_4987,N_2913);
and U7296 (N_7296,N_4863,N_3244);
and U7297 (N_7297,N_4494,N_3055);
or U7298 (N_7298,N_4953,N_4749);
or U7299 (N_7299,N_4369,N_2781);
xnor U7300 (N_7300,N_2952,N_4818);
xor U7301 (N_7301,N_4758,N_3582);
nor U7302 (N_7302,N_3685,N_3458);
or U7303 (N_7303,N_4874,N_4881);
and U7304 (N_7304,N_3845,N_3976);
xor U7305 (N_7305,N_3768,N_3235);
and U7306 (N_7306,N_3531,N_3801);
or U7307 (N_7307,N_2745,N_4059);
xor U7308 (N_7308,N_2507,N_3556);
nand U7309 (N_7309,N_4898,N_2514);
xnor U7310 (N_7310,N_4476,N_2954);
or U7311 (N_7311,N_4401,N_2665);
nor U7312 (N_7312,N_4020,N_4917);
nand U7313 (N_7313,N_3064,N_4382);
nor U7314 (N_7314,N_3944,N_2904);
or U7315 (N_7315,N_3357,N_4965);
nor U7316 (N_7316,N_4250,N_3737);
nand U7317 (N_7317,N_3435,N_2613);
or U7318 (N_7318,N_3426,N_4180);
nand U7319 (N_7319,N_4686,N_3323);
nand U7320 (N_7320,N_4795,N_4275);
nand U7321 (N_7321,N_3998,N_3411);
or U7322 (N_7322,N_2650,N_3493);
nor U7323 (N_7323,N_3194,N_4131);
and U7324 (N_7324,N_3486,N_4233);
or U7325 (N_7325,N_2827,N_4960);
xor U7326 (N_7326,N_4327,N_4653);
or U7327 (N_7327,N_3250,N_4396);
xor U7328 (N_7328,N_4226,N_4690);
or U7329 (N_7329,N_3582,N_3707);
nand U7330 (N_7330,N_2775,N_4266);
and U7331 (N_7331,N_4178,N_4652);
xnor U7332 (N_7332,N_4268,N_4013);
and U7333 (N_7333,N_4211,N_2863);
and U7334 (N_7334,N_4607,N_4149);
xor U7335 (N_7335,N_3660,N_2705);
nor U7336 (N_7336,N_4339,N_4000);
nor U7337 (N_7337,N_4228,N_3150);
nor U7338 (N_7338,N_4291,N_3536);
xnor U7339 (N_7339,N_4826,N_2691);
or U7340 (N_7340,N_3302,N_2666);
or U7341 (N_7341,N_3141,N_2623);
nand U7342 (N_7342,N_2912,N_4826);
xnor U7343 (N_7343,N_4900,N_4007);
xor U7344 (N_7344,N_2803,N_2632);
and U7345 (N_7345,N_3946,N_2996);
xor U7346 (N_7346,N_3371,N_2659);
or U7347 (N_7347,N_3655,N_3805);
nor U7348 (N_7348,N_3492,N_3063);
nand U7349 (N_7349,N_4140,N_3372);
or U7350 (N_7350,N_4953,N_3828);
or U7351 (N_7351,N_2682,N_2631);
xor U7352 (N_7352,N_2744,N_3001);
or U7353 (N_7353,N_3076,N_3189);
nor U7354 (N_7354,N_4427,N_4938);
nand U7355 (N_7355,N_3676,N_4400);
or U7356 (N_7356,N_3418,N_3080);
and U7357 (N_7357,N_4354,N_4672);
nor U7358 (N_7358,N_4405,N_2861);
nor U7359 (N_7359,N_4497,N_4014);
and U7360 (N_7360,N_2738,N_4329);
xor U7361 (N_7361,N_3309,N_3491);
nand U7362 (N_7362,N_4539,N_3381);
and U7363 (N_7363,N_4930,N_3860);
xnor U7364 (N_7364,N_4197,N_3554);
nor U7365 (N_7365,N_4569,N_4746);
nor U7366 (N_7366,N_3656,N_4833);
and U7367 (N_7367,N_3123,N_4258);
xnor U7368 (N_7368,N_4418,N_3304);
nand U7369 (N_7369,N_3423,N_3959);
nor U7370 (N_7370,N_3606,N_2984);
nor U7371 (N_7371,N_3568,N_3690);
nand U7372 (N_7372,N_4157,N_4255);
xor U7373 (N_7373,N_3469,N_4666);
nand U7374 (N_7374,N_3069,N_3606);
nand U7375 (N_7375,N_4605,N_4906);
and U7376 (N_7376,N_2976,N_2843);
nor U7377 (N_7377,N_4023,N_3132);
and U7378 (N_7378,N_2749,N_2642);
xnor U7379 (N_7379,N_3797,N_2795);
nor U7380 (N_7380,N_2513,N_4419);
or U7381 (N_7381,N_3742,N_4552);
or U7382 (N_7382,N_4559,N_4492);
nand U7383 (N_7383,N_4076,N_4714);
nand U7384 (N_7384,N_4019,N_3578);
nand U7385 (N_7385,N_3297,N_4626);
xnor U7386 (N_7386,N_4052,N_3780);
nor U7387 (N_7387,N_4978,N_2827);
or U7388 (N_7388,N_2991,N_4317);
nor U7389 (N_7389,N_3216,N_4758);
nor U7390 (N_7390,N_2900,N_2874);
and U7391 (N_7391,N_4079,N_4511);
nand U7392 (N_7392,N_4999,N_4931);
nand U7393 (N_7393,N_3042,N_4184);
nor U7394 (N_7394,N_4170,N_3115);
xor U7395 (N_7395,N_3977,N_4991);
or U7396 (N_7396,N_3067,N_2917);
nand U7397 (N_7397,N_3710,N_4013);
xnor U7398 (N_7398,N_3425,N_4565);
or U7399 (N_7399,N_4559,N_3094);
nor U7400 (N_7400,N_3713,N_4778);
or U7401 (N_7401,N_2737,N_2899);
and U7402 (N_7402,N_3866,N_4207);
xor U7403 (N_7403,N_4713,N_4976);
nor U7404 (N_7404,N_3314,N_3808);
nor U7405 (N_7405,N_2776,N_2905);
nand U7406 (N_7406,N_3292,N_3332);
xor U7407 (N_7407,N_2790,N_4177);
or U7408 (N_7408,N_3517,N_2864);
xor U7409 (N_7409,N_3729,N_4113);
and U7410 (N_7410,N_4009,N_2781);
nor U7411 (N_7411,N_3625,N_4294);
nand U7412 (N_7412,N_2699,N_3785);
and U7413 (N_7413,N_4170,N_4694);
nand U7414 (N_7414,N_3394,N_4714);
nor U7415 (N_7415,N_3547,N_3648);
nand U7416 (N_7416,N_2643,N_4032);
and U7417 (N_7417,N_3383,N_2569);
nor U7418 (N_7418,N_4802,N_4842);
nor U7419 (N_7419,N_2889,N_3787);
nand U7420 (N_7420,N_3524,N_4020);
nand U7421 (N_7421,N_4892,N_3813);
or U7422 (N_7422,N_3568,N_2960);
nor U7423 (N_7423,N_2796,N_3212);
xor U7424 (N_7424,N_3817,N_2549);
nand U7425 (N_7425,N_3593,N_3386);
nand U7426 (N_7426,N_4933,N_2606);
and U7427 (N_7427,N_4326,N_4896);
or U7428 (N_7428,N_4753,N_2709);
nor U7429 (N_7429,N_3896,N_2592);
and U7430 (N_7430,N_3541,N_2808);
nand U7431 (N_7431,N_3361,N_3107);
nand U7432 (N_7432,N_3404,N_4864);
nor U7433 (N_7433,N_2915,N_3264);
nand U7434 (N_7434,N_4560,N_3368);
or U7435 (N_7435,N_2551,N_3996);
nor U7436 (N_7436,N_3678,N_3081);
or U7437 (N_7437,N_3754,N_3988);
nor U7438 (N_7438,N_3137,N_4911);
or U7439 (N_7439,N_3483,N_3185);
or U7440 (N_7440,N_3418,N_3385);
nor U7441 (N_7441,N_4066,N_4465);
xnor U7442 (N_7442,N_3763,N_4289);
nor U7443 (N_7443,N_3658,N_3564);
and U7444 (N_7444,N_2946,N_3861);
and U7445 (N_7445,N_3945,N_3947);
nand U7446 (N_7446,N_2839,N_4242);
xnor U7447 (N_7447,N_2593,N_3274);
xor U7448 (N_7448,N_4844,N_3502);
xor U7449 (N_7449,N_3386,N_3463);
xor U7450 (N_7450,N_4060,N_3329);
nand U7451 (N_7451,N_3941,N_2661);
xnor U7452 (N_7452,N_4528,N_3764);
xnor U7453 (N_7453,N_2534,N_2617);
and U7454 (N_7454,N_3497,N_4356);
and U7455 (N_7455,N_4357,N_2557);
xor U7456 (N_7456,N_2976,N_4403);
xnor U7457 (N_7457,N_2946,N_4668);
and U7458 (N_7458,N_4728,N_3217);
xnor U7459 (N_7459,N_2814,N_3486);
nand U7460 (N_7460,N_2835,N_3344);
nor U7461 (N_7461,N_4435,N_3417);
and U7462 (N_7462,N_4413,N_2898);
nor U7463 (N_7463,N_4839,N_2856);
nand U7464 (N_7464,N_4425,N_3561);
xnor U7465 (N_7465,N_3011,N_3793);
xor U7466 (N_7466,N_4361,N_3479);
nand U7467 (N_7467,N_4145,N_4840);
nand U7468 (N_7468,N_2943,N_3443);
nand U7469 (N_7469,N_3200,N_3443);
or U7470 (N_7470,N_2557,N_2985);
xor U7471 (N_7471,N_4235,N_4757);
or U7472 (N_7472,N_2664,N_3315);
xnor U7473 (N_7473,N_4649,N_3233);
and U7474 (N_7474,N_3204,N_4690);
nor U7475 (N_7475,N_4196,N_2605);
and U7476 (N_7476,N_4708,N_3488);
xnor U7477 (N_7477,N_3909,N_2694);
nor U7478 (N_7478,N_3844,N_4602);
nand U7479 (N_7479,N_3825,N_4780);
nor U7480 (N_7480,N_3886,N_4178);
xnor U7481 (N_7481,N_3029,N_3857);
nor U7482 (N_7482,N_4814,N_4461);
and U7483 (N_7483,N_4377,N_4426);
xnor U7484 (N_7484,N_2826,N_4415);
nand U7485 (N_7485,N_4872,N_4099);
nand U7486 (N_7486,N_3001,N_3249);
xnor U7487 (N_7487,N_2960,N_4230);
xnor U7488 (N_7488,N_2531,N_3488);
or U7489 (N_7489,N_3836,N_4436);
nor U7490 (N_7490,N_4370,N_3367);
xnor U7491 (N_7491,N_3563,N_4287);
nand U7492 (N_7492,N_2808,N_4789);
and U7493 (N_7493,N_3493,N_4879);
nand U7494 (N_7494,N_3686,N_3096);
nor U7495 (N_7495,N_4262,N_2895);
nor U7496 (N_7496,N_4453,N_2885);
nand U7497 (N_7497,N_3978,N_3471);
or U7498 (N_7498,N_2949,N_2964);
xor U7499 (N_7499,N_3975,N_4949);
and U7500 (N_7500,N_5525,N_6040);
and U7501 (N_7501,N_7102,N_5091);
nand U7502 (N_7502,N_6737,N_6326);
nor U7503 (N_7503,N_5177,N_5035);
nand U7504 (N_7504,N_5768,N_6334);
nor U7505 (N_7505,N_5910,N_7327);
xor U7506 (N_7506,N_6674,N_6841);
xnor U7507 (N_7507,N_6171,N_7272);
nor U7508 (N_7508,N_6313,N_5899);
nand U7509 (N_7509,N_7056,N_5463);
and U7510 (N_7510,N_6468,N_6542);
nand U7511 (N_7511,N_5183,N_6663);
and U7512 (N_7512,N_6933,N_5971);
or U7513 (N_7513,N_6562,N_5948);
xnor U7514 (N_7514,N_6853,N_6776);
xor U7515 (N_7515,N_6508,N_5484);
or U7516 (N_7516,N_7184,N_6805);
xnor U7517 (N_7517,N_6646,N_5278);
nor U7518 (N_7518,N_6457,N_6812);
nand U7519 (N_7519,N_7059,N_7208);
or U7520 (N_7520,N_6952,N_5606);
nor U7521 (N_7521,N_5917,N_5478);
and U7522 (N_7522,N_5189,N_5782);
xor U7523 (N_7523,N_6193,N_6125);
nand U7524 (N_7524,N_6200,N_6070);
xor U7525 (N_7525,N_5018,N_5591);
xor U7526 (N_7526,N_6099,N_5733);
xnor U7527 (N_7527,N_6860,N_7290);
nand U7528 (N_7528,N_7108,N_7177);
nand U7529 (N_7529,N_6021,N_5731);
nand U7530 (N_7530,N_6247,N_6404);
nor U7531 (N_7531,N_5653,N_6027);
nor U7532 (N_7532,N_5561,N_6991);
nand U7533 (N_7533,N_5944,N_6938);
xor U7534 (N_7534,N_6332,N_6681);
nor U7535 (N_7535,N_5406,N_6036);
and U7536 (N_7536,N_5480,N_6115);
nor U7537 (N_7537,N_6791,N_5660);
xor U7538 (N_7538,N_5119,N_5316);
and U7539 (N_7539,N_6561,N_6999);
xor U7540 (N_7540,N_6441,N_6921);
and U7541 (N_7541,N_6240,N_5643);
nand U7542 (N_7542,N_6996,N_5073);
and U7543 (N_7543,N_6611,N_5848);
xor U7544 (N_7544,N_5248,N_7380);
and U7545 (N_7545,N_6934,N_5031);
and U7546 (N_7546,N_7419,N_5900);
xnor U7547 (N_7547,N_7048,N_6594);
or U7548 (N_7548,N_6294,N_5760);
nand U7549 (N_7549,N_7231,N_5281);
nor U7550 (N_7550,N_5121,N_5855);
and U7551 (N_7551,N_5338,N_7169);
nor U7552 (N_7552,N_6945,N_7483);
or U7553 (N_7553,N_5328,N_6908);
xor U7554 (N_7554,N_6146,N_7396);
xnor U7555 (N_7555,N_6979,N_5904);
and U7556 (N_7556,N_5791,N_5418);
and U7557 (N_7557,N_6821,N_5802);
nand U7558 (N_7558,N_6721,N_5886);
nand U7559 (N_7559,N_5398,N_5505);
and U7560 (N_7560,N_7073,N_7388);
xor U7561 (N_7561,N_5599,N_6044);
xnor U7562 (N_7562,N_6621,N_5257);
or U7563 (N_7563,N_5506,N_7426);
nor U7564 (N_7564,N_5934,N_6467);
or U7565 (N_7565,N_6175,N_5079);
or U7566 (N_7566,N_6961,N_7461);
and U7567 (N_7567,N_6992,N_6768);
xnor U7568 (N_7568,N_7287,N_7174);
nor U7569 (N_7569,N_6850,N_6603);
nand U7570 (N_7570,N_6595,N_6904);
nand U7571 (N_7571,N_5265,N_6571);
xor U7572 (N_7572,N_5454,N_5854);
or U7573 (N_7573,N_5260,N_5523);
nor U7574 (N_7574,N_6394,N_5448);
nor U7575 (N_7575,N_5610,N_6723);
xor U7576 (N_7576,N_5727,N_5825);
or U7577 (N_7577,N_6453,N_5024);
xnor U7578 (N_7578,N_7376,N_5077);
nand U7579 (N_7579,N_5613,N_6731);
or U7580 (N_7580,N_7082,N_5704);
and U7581 (N_7581,N_7399,N_5542);
or U7582 (N_7582,N_5647,N_5773);
and U7583 (N_7583,N_6192,N_6652);
nand U7584 (N_7584,N_5864,N_5179);
or U7585 (N_7585,N_5047,N_7432);
nor U7586 (N_7586,N_6423,N_5284);
xnor U7587 (N_7587,N_6118,N_5043);
nand U7588 (N_7588,N_7098,N_6042);
nand U7589 (N_7589,N_7038,N_7418);
or U7590 (N_7590,N_5799,N_6108);
xnor U7591 (N_7591,N_6566,N_5269);
nor U7592 (N_7592,N_6740,N_6015);
xnor U7593 (N_7593,N_6579,N_6196);
nor U7594 (N_7594,N_6151,N_5897);
nor U7595 (N_7595,N_6228,N_6254);
nor U7596 (N_7596,N_7394,N_6762);
nor U7597 (N_7597,N_6249,N_5126);
or U7598 (N_7598,N_6225,N_5819);
xnor U7599 (N_7599,N_5710,N_7025);
xor U7600 (N_7600,N_7391,N_7349);
nand U7601 (N_7601,N_7252,N_5962);
and U7602 (N_7602,N_6823,N_5714);
or U7603 (N_7603,N_5539,N_7055);
nor U7604 (N_7604,N_6418,N_6742);
nor U7605 (N_7605,N_6414,N_7341);
and U7606 (N_7606,N_5608,N_7053);
nand U7607 (N_7607,N_6524,N_6431);
xor U7608 (N_7608,N_5258,N_6083);
xor U7609 (N_7609,N_7360,N_7157);
or U7610 (N_7610,N_5354,N_6666);
nand U7611 (N_7611,N_6887,N_6492);
and U7612 (N_7612,N_6158,N_6475);
nor U7613 (N_7613,N_6845,N_7115);
nand U7614 (N_7614,N_7223,N_5429);
and U7615 (N_7615,N_7144,N_7135);
nor U7616 (N_7616,N_6871,N_5129);
and U7617 (N_7617,N_5438,N_6459);
or U7618 (N_7618,N_5923,N_5605);
or U7619 (N_7619,N_5957,N_7482);
nor U7620 (N_7620,N_5088,N_5784);
or U7621 (N_7621,N_7291,N_6943);
or U7622 (N_7622,N_7202,N_6310);
and U7623 (N_7623,N_5026,N_6019);
or U7624 (N_7624,N_6339,N_6710);
nor U7625 (N_7625,N_5351,N_5431);
nor U7626 (N_7626,N_6064,N_6828);
xnor U7627 (N_7627,N_7337,N_6268);
nand U7628 (N_7628,N_6429,N_5973);
and U7629 (N_7629,N_6382,N_5204);
nor U7630 (N_7630,N_5102,N_5777);
and U7631 (N_7631,N_6062,N_7281);
nand U7632 (N_7632,N_5548,N_6587);
or U7633 (N_7633,N_6202,N_6329);
nand U7634 (N_7634,N_6144,N_6648);
nor U7635 (N_7635,N_6137,N_5860);
nand U7636 (N_7636,N_6642,N_5215);
xnor U7637 (N_7637,N_6834,N_7370);
and U7638 (N_7638,N_6464,N_7229);
or U7639 (N_7639,N_6609,N_5198);
nor U7640 (N_7640,N_7348,N_6435);
xnor U7641 (N_7641,N_5675,N_5672);
nand U7642 (N_7642,N_5416,N_5410);
xor U7643 (N_7643,N_5015,N_6773);
and U7644 (N_7644,N_6503,N_5585);
xor U7645 (N_7645,N_5779,N_6278);
nor U7646 (N_7646,N_6061,N_6830);
and U7647 (N_7647,N_5763,N_6803);
nand U7648 (N_7648,N_6886,N_7232);
or U7649 (N_7649,N_5786,N_7012);
nand U7650 (N_7650,N_5692,N_5130);
xor U7651 (N_7651,N_6891,N_6975);
or U7652 (N_7652,N_5170,N_7484);
nand U7653 (N_7653,N_6550,N_6946);
or U7654 (N_7654,N_5521,N_5989);
nor U7655 (N_7655,N_5063,N_5114);
and U7656 (N_7656,N_6585,N_6136);
xnor U7657 (N_7657,N_7143,N_6476);
or U7658 (N_7658,N_7270,N_5814);
xor U7659 (N_7659,N_6815,N_7475);
nor U7660 (N_7660,N_7140,N_7487);
and U7661 (N_7661,N_6427,N_6884);
xnor U7662 (N_7662,N_6460,N_5684);
or U7663 (N_7663,N_6417,N_5137);
nand U7664 (N_7664,N_5002,N_6284);
and U7665 (N_7665,N_6927,N_6638);
nor U7666 (N_7666,N_6483,N_6356);
nor U7667 (N_7667,N_7437,N_7180);
nand U7668 (N_7668,N_6288,N_5566);
nand U7669 (N_7669,N_6289,N_5845);
or U7670 (N_7670,N_6195,N_6632);
xor U7671 (N_7671,N_5027,N_6665);
nand U7672 (N_7672,N_5755,N_5742);
nor U7673 (N_7673,N_5946,N_6743);
nand U7674 (N_7674,N_5964,N_7105);
and U7675 (N_7675,N_7091,N_6543);
nand U7676 (N_7676,N_5787,N_7197);
and U7677 (N_7677,N_7317,N_6224);
or U7678 (N_7678,N_7142,N_5686);
nand U7679 (N_7679,N_5828,N_6772);
nand U7680 (N_7680,N_5912,N_5303);
xnor U7681 (N_7681,N_7479,N_7268);
nor U7682 (N_7682,N_6635,N_7468);
nand U7683 (N_7683,N_5477,N_5630);
nor U7684 (N_7684,N_5052,N_6656);
and U7685 (N_7685,N_7416,N_5430);
nand U7686 (N_7686,N_6101,N_6657);
or U7687 (N_7687,N_5370,N_5576);
nor U7688 (N_7688,N_5444,N_5364);
xnor U7689 (N_7689,N_6135,N_7440);
nand U7690 (N_7690,N_7477,N_5003);
xor U7691 (N_7691,N_6113,N_6533);
nor U7692 (N_7692,N_6563,N_6654);
or U7693 (N_7693,N_6026,N_5373);
or U7694 (N_7694,N_7023,N_5007);
nand U7695 (N_7695,N_5453,N_7490);
nor U7696 (N_7696,N_6461,N_7246);
xor U7697 (N_7697,N_6245,N_6962);
and U7698 (N_7698,N_5180,N_6680);
or U7699 (N_7699,N_5867,N_5166);
and U7700 (N_7700,N_7464,N_7068);
nor U7701 (N_7701,N_5875,N_7251);
nor U7702 (N_7702,N_6555,N_7168);
nand U7703 (N_7703,N_5276,N_5483);
nor U7704 (N_7704,N_5986,N_6341);
xor U7705 (N_7705,N_5642,N_7131);
or U7706 (N_7706,N_6170,N_6207);
nor U7707 (N_7707,N_5116,N_5876);
or U7708 (N_7708,N_5175,N_5865);
and U7709 (N_7709,N_5305,N_5626);
xnor U7710 (N_7710,N_5646,N_6520);
and U7711 (N_7711,N_5333,N_7084);
and U7712 (N_7712,N_7473,N_7271);
nand U7713 (N_7713,N_5829,N_5769);
nor U7714 (N_7714,N_6390,N_6606);
xnor U7715 (N_7715,N_5020,N_7274);
and U7716 (N_7716,N_6756,N_7412);
nand U7717 (N_7717,N_6717,N_5868);
xnor U7718 (N_7718,N_5509,N_7218);
nand U7719 (N_7719,N_6628,N_6682);
nor U7720 (N_7720,N_6451,N_7088);
xor U7721 (N_7721,N_5690,N_6159);
or U7722 (N_7722,N_7211,N_5856);
nand U7723 (N_7723,N_5176,N_5010);
or U7724 (N_7724,N_7499,N_7361);
nand U7725 (N_7725,N_6644,N_6802);
nand U7726 (N_7726,N_5174,N_5301);
xnor U7727 (N_7727,N_6400,N_6967);
xor U7728 (N_7728,N_7465,N_5913);
nand U7729 (N_7729,N_6867,N_6258);
nor U7730 (N_7730,N_5302,N_5013);
and U7731 (N_7731,N_6793,N_6735);
nor U7732 (N_7732,N_5218,N_6728);
and U7733 (N_7733,N_6795,N_6139);
nand U7734 (N_7734,N_6469,N_5232);
or U7735 (N_7735,N_5805,N_6813);
or U7736 (N_7736,N_7224,N_5665);
or U7737 (N_7737,N_7020,N_5834);
or U7738 (N_7738,N_5161,N_5901);
nand U7739 (N_7739,N_6864,N_7449);
and U7740 (N_7740,N_5261,N_7097);
nor U7741 (N_7741,N_5072,N_7421);
or U7742 (N_7742,N_6152,N_5289);
nor U7743 (N_7743,N_7233,N_6573);
nand U7744 (N_7744,N_6488,N_6715);
xor U7745 (N_7745,N_7090,N_6033);
nor U7746 (N_7746,N_5931,N_5987);
and U7747 (N_7747,N_7205,N_7194);
nand U7748 (N_7748,N_5963,N_5103);
xnor U7749 (N_7749,N_5412,N_5492);
nor U7750 (N_7750,N_6003,N_7248);
nor U7751 (N_7751,N_5649,N_6865);
xor U7752 (N_7752,N_6765,N_6279);
and U7753 (N_7753,N_5030,N_7123);
and U7754 (N_7754,N_5551,N_5751);
and U7755 (N_7755,N_6506,N_5304);
xnor U7756 (N_7756,N_7267,N_7442);
nand U7757 (N_7757,N_5283,N_5723);
xor U7758 (N_7758,N_6499,N_7052);
nor U7759 (N_7759,N_5034,N_6035);
or U7760 (N_7760,N_6025,N_6489);
and U7761 (N_7761,N_6068,N_6017);
and U7762 (N_7762,N_7235,N_5563);
and U7763 (N_7763,N_5472,N_7339);
and U7764 (N_7764,N_6174,N_5375);
and U7765 (N_7765,N_6944,N_6291);
nand U7766 (N_7766,N_7286,N_6379);
xor U7767 (N_7767,N_7301,N_5597);
nand U7768 (N_7768,N_6916,N_5350);
or U7769 (N_7769,N_5107,N_6719);
nor U7770 (N_7770,N_5253,N_5568);
and U7771 (N_7771,N_7069,N_5233);
xnor U7772 (N_7772,N_7104,N_5614);
or U7773 (N_7773,N_6712,N_7423);
nand U7774 (N_7774,N_6157,N_7334);
nor U7775 (N_7775,N_5231,N_5437);
nor U7776 (N_7776,N_5556,N_7436);
or U7777 (N_7777,N_6301,N_5244);
xnor U7778 (N_7778,N_6403,N_5889);
nor U7779 (N_7779,N_6698,N_6127);
and U7780 (N_7780,N_6620,N_6368);
nand U7781 (N_7781,N_6090,N_6650);
or U7782 (N_7782,N_6337,N_7491);
xor U7783 (N_7783,N_7403,N_5389);
or U7784 (N_7784,N_6617,N_7315);
xor U7785 (N_7785,N_7352,N_7351);
or U7786 (N_7786,N_7256,N_6187);
nor U7787 (N_7787,N_5099,N_5827);
and U7788 (N_7788,N_7458,N_6714);
or U7789 (N_7789,N_5718,N_5157);
nor U7790 (N_7790,N_6007,N_5633);
and U7791 (N_7791,N_5136,N_7381);
and U7792 (N_7792,N_6204,N_6422);
xor U7793 (N_7793,N_6747,N_5801);
and U7794 (N_7794,N_5427,N_7431);
nor U7795 (N_7795,N_5206,N_6535);
and U7796 (N_7796,N_6842,N_6761);
nor U7797 (N_7797,N_6119,N_6071);
xnor U7798 (N_7798,N_6839,N_6223);
xor U7799 (N_7799,N_5255,N_5851);
xor U7800 (N_7800,N_6325,N_5006);
nand U7801 (N_7801,N_7225,N_5458);
nand U7802 (N_7802,N_5343,N_7200);
and U7803 (N_7803,N_6079,N_5131);
and U7804 (N_7804,N_6335,N_6748);
xor U7805 (N_7805,N_6924,N_6148);
or U7806 (N_7806,N_5342,N_5312);
nor U7807 (N_7807,N_5881,N_5739);
nand U7808 (N_7808,N_5732,N_5330);
nand U7809 (N_7809,N_6643,N_5890);
xor U7810 (N_7810,N_6576,N_6804);
and U7811 (N_7811,N_5683,N_6679);
nor U7812 (N_7812,N_5325,N_7002);
nor U7813 (N_7813,N_5474,N_7398);
and U7814 (N_7814,N_6234,N_5720);
nor U7815 (N_7815,N_5520,N_6655);
nor U7816 (N_7816,N_5788,N_7463);
and U7817 (N_7817,N_6434,N_5420);
nand U7818 (N_7818,N_5981,N_6969);
nand U7819 (N_7819,N_5902,N_5296);
nor U7820 (N_7820,N_6614,N_5462);
nand U7821 (N_7821,N_5836,N_5611);
or U7822 (N_7822,N_6843,N_6676);
xor U7823 (N_7823,N_6265,N_6769);
and U7824 (N_7824,N_5128,N_7446);
and U7825 (N_7825,N_6362,N_7015);
nor U7826 (N_7826,N_6482,N_7298);
nand U7827 (N_7827,N_5122,N_6892);
nor U7828 (N_7828,N_6153,N_6527);
nand U7829 (N_7829,N_7085,N_5880);
or U7830 (N_7830,N_6080,N_5123);
nor U7831 (N_7831,N_6421,N_5673);
nand U7832 (N_7832,N_5862,N_5067);
or U7833 (N_7833,N_6906,N_7201);
xnor U7834 (N_7834,N_6531,N_5615);
nand U7835 (N_7835,N_5470,N_6093);
or U7836 (N_7836,N_6505,N_6217);
and U7837 (N_7837,N_7259,N_6824);
or U7838 (N_7838,N_6221,N_6911);
and U7839 (N_7839,N_5682,N_7365);
xor U7840 (N_7840,N_7016,N_5371);
xnor U7841 (N_7841,N_6141,N_5199);
or U7842 (N_7842,N_6704,N_5572);
or U7843 (N_7843,N_7187,N_5019);
nand U7844 (N_7844,N_6311,N_6399);
or U7845 (N_7845,N_7162,N_6833);
xnor U7846 (N_7846,N_6408,N_5691);
nand U7847 (N_7847,N_5994,N_5620);
nor U7848 (N_7848,N_6402,N_5311);
xnor U7849 (N_7849,N_5565,N_5142);
xor U7850 (N_7850,N_5824,N_5236);
xor U7851 (N_7851,N_5515,N_7347);
and U7852 (N_7852,N_7127,N_6951);
nor U7853 (N_7853,N_5885,N_7126);
and U7854 (N_7854,N_7378,N_6686);
nor U7855 (N_7855,N_6616,N_5307);
and U7856 (N_7856,N_5042,N_6495);
nor U7857 (N_7857,N_7249,N_6636);
nand U7858 (N_7858,N_5587,N_5872);
nand U7859 (N_7859,N_5830,N_7321);
and U7860 (N_7860,N_5266,N_7489);
xnor U7861 (N_7861,N_6333,N_5849);
and U7862 (N_7862,N_5400,N_5348);
nor U7863 (N_7863,N_6954,N_6602);
nor U7864 (N_7864,N_6770,N_6757);
nand U7865 (N_7865,N_7447,N_5961);
or U7866 (N_7866,N_5165,N_5703);
and U7867 (N_7867,N_5979,N_7092);
nand U7868 (N_7868,N_7471,N_5616);
nor U7869 (N_7869,N_5590,N_5071);
xor U7870 (N_7870,N_6327,N_6436);
nor U7871 (N_7871,N_7007,N_7003);
xor U7872 (N_7872,N_5436,N_5424);
or U7873 (N_7873,N_7179,N_7001);
and U7874 (N_7874,N_5972,N_5947);
or U7875 (N_7875,N_5060,N_7243);
nor U7876 (N_7876,N_7226,N_7306);
xor U7877 (N_7877,N_5861,N_5104);
nand U7878 (N_7878,N_5096,N_5816);
xnor U7879 (N_7879,N_6893,N_6560);
or U7880 (N_7880,N_6208,N_7011);
xor U7881 (N_7881,N_7428,N_7240);
nand U7882 (N_7882,N_5150,N_7032);
and U7883 (N_7883,N_6359,N_5882);
nand U7884 (N_7884,N_6835,N_6960);
nand U7885 (N_7885,N_5722,N_7217);
xnor U7886 (N_7886,N_5202,N_6558);
and U7887 (N_7887,N_5135,N_5120);
nand U7888 (N_7888,N_6182,N_5387);
and U7889 (N_7889,N_5883,N_6350);
and U7890 (N_7890,N_7216,N_7386);
nand U7891 (N_7891,N_6354,N_6425);
or U7892 (N_7892,N_6913,N_6829);
and U7893 (N_7893,N_6391,N_6696);
and U7894 (N_7894,N_6716,N_5577);
or U7895 (N_7895,N_6154,N_6898);
nor U7896 (N_7896,N_5291,N_5011);
and U7897 (N_7897,N_6971,N_5794);
nand U7898 (N_7898,N_5087,N_5347);
nand U7899 (N_7899,N_5295,N_6789);
and U7900 (N_7900,N_6599,N_5413);
nor U7901 (N_7901,N_6510,N_6570);
xnor U7902 (N_7902,N_7100,N_5967);
and U7903 (N_7903,N_5826,N_7146);
xor U7904 (N_7904,N_6037,N_5298);
or U7905 (N_7905,N_6229,N_5778);
or U7906 (N_7906,N_5871,N_7379);
xnor U7907 (N_7907,N_5776,N_5455);
or U7908 (N_7908,N_6653,N_7313);
nand U7909 (N_7909,N_7387,N_7096);
nor U7910 (N_7910,N_5532,N_5451);
nor U7911 (N_7911,N_7289,N_7439);
nand U7912 (N_7912,N_6211,N_5084);
xnor U7913 (N_7913,N_6702,N_5040);
and U7914 (N_7914,N_5155,N_5663);
nor U7915 (N_7915,N_6832,N_5894);
nor U7916 (N_7916,N_6940,N_6222);
nor U7917 (N_7917,N_7171,N_5208);
and U7918 (N_7918,N_6697,N_6197);
nand U7919 (N_7919,N_6669,N_5997);
or U7920 (N_7920,N_7415,N_6303);
and U7921 (N_7921,N_5637,N_6667);
nand U7922 (N_7922,N_6220,N_6094);
or U7923 (N_7923,N_7472,N_5671);
and U7924 (N_7924,N_5489,N_5666);
or U7925 (N_7925,N_6963,N_6377);
and U7926 (N_7926,N_7342,N_5110);
nand U7927 (N_7927,N_5391,N_6257);
and U7928 (N_7928,N_5803,N_6639);
nor U7929 (N_7929,N_5639,N_6477);
or U7930 (N_7930,N_6713,N_6156);
and U7931 (N_7931,N_6965,N_6388);
nand U7932 (N_7932,N_6078,N_6364);
or U7933 (N_7933,N_6880,N_5447);
and U7934 (N_7934,N_6130,N_7283);
xnor U7935 (N_7935,N_6371,N_6491);
nand U7936 (N_7936,N_5243,N_5239);
and U7937 (N_7937,N_5309,N_6138);
and U7938 (N_7938,N_5906,N_7039);
xor U7939 (N_7939,N_6444,N_5173);
or U7940 (N_7940,N_5212,N_5541);
nand U7941 (N_7941,N_5941,N_5094);
nor U7942 (N_7942,N_5399,N_7480);
xnor U7943 (N_7943,N_5547,N_6318);
or U7944 (N_7944,N_7116,N_6440);
and U7945 (N_7945,N_5395,N_5428);
nor U7946 (N_7946,N_7101,N_6903);
or U7947 (N_7947,N_6109,N_6816);
and U7948 (N_7948,N_5092,N_5842);
and U7949 (N_7949,N_5057,N_5196);
nand U7950 (N_7950,N_6045,N_7124);
or U7951 (N_7951,N_6057,N_5841);
nand U7952 (N_7952,N_7138,N_5262);
or U7953 (N_7953,N_5441,N_6690);
and U7954 (N_7954,N_5508,N_5440);
nand U7955 (N_7955,N_6677,N_5115);
nand U7956 (N_7956,N_5744,N_7300);
or U7957 (N_7957,N_6780,N_5640);
nor U7958 (N_7958,N_6806,N_7139);
and U7959 (N_7959,N_5061,N_6428);
or U7960 (N_7960,N_5669,N_5911);
nor U7961 (N_7961,N_6647,N_7395);
xor U7962 (N_7962,N_7408,N_7434);
nor U7963 (N_7963,N_6264,N_7114);
nor U7964 (N_7964,N_5983,N_6375);
and U7965 (N_7965,N_6072,N_6393);
xor U7966 (N_7966,N_6557,N_6866);
nor U7967 (N_7967,N_6324,N_7221);
or U7968 (N_7968,N_6395,N_5488);
or U7969 (N_7969,N_6668,N_5409);
xnor U7970 (N_7970,N_6948,N_5001);
or U7971 (N_7971,N_5661,N_5449);
xor U7972 (N_7972,N_5334,N_7329);
nor U7973 (N_7973,N_5992,N_6862);
nor U7974 (N_7974,N_6023,N_5937);
or U7975 (N_7975,N_5693,N_7081);
xnor U7976 (N_7976,N_5792,N_6902);
and U7977 (N_7977,N_5192,N_6857);
nand U7978 (N_7978,N_6352,N_6092);
and U7979 (N_7979,N_6760,N_6928);
nor U7980 (N_7980,N_5602,N_5279);
nand U7981 (N_7981,N_5461,N_7215);
and U7982 (N_7982,N_7343,N_5160);
or U7983 (N_7983,N_6013,N_6670);
xnor U7984 (N_7984,N_6994,N_7372);
nor U7985 (N_7985,N_5340,N_5594);
nor U7986 (N_7986,N_5538,N_6896);
and U7987 (N_7987,N_6047,N_5887);
nor U7988 (N_7988,N_5273,N_5632);
and U7989 (N_7989,N_5153,N_7427);
nor U7990 (N_7990,N_6889,N_6442);
nor U7991 (N_7991,N_5949,N_6559);
nand U7992 (N_7992,N_5790,N_7377);
nand U7993 (N_7993,N_5724,N_7006);
nor U7994 (N_7994,N_6840,N_5200);
nand U7995 (N_7995,N_6077,N_5361);
or U7996 (N_7996,N_6981,N_5044);
xor U7997 (N_7997,N_6116,N_5725);
nand U7998 (N_7998,N_5452,N_6122);
and U7999 (N_7999,N_5028,N_5924);
xnor U8000 (N_8000,N_6320,N_6844);
xnor U8001 (N_8001,N_7278,N_6447);
nand U8002 (N_8002,N_7155,N_6631);
and U8003 (N_8003,N_6604,N_5729);
and U8004 (N_8004,N_7266,N_7182);
xor U8005 (N_8005,N_6360,N_7474);
xnor U8006 (N_8006,N_6831,N_5815);
and U8007 (N_8007,N_6340,N_7460);
and U8008 (N_8008,N_6107,N_7459);
nor U8009 (N_8009,N_6235,N_5171);
xor U8010 (N_8010,N_6009,N_6822);
and U8011 (N_8011,N_5230,N_6104);
and U8012 (N_8012,N_6302,N_5874);
nor U8013 (N_8013,N_5764,N_6519);
nand U8014 (N_8014,N_6338,N_5918);
nand U8015 (N_8015,N_5039,N_5250);
xnor U8016 (N_8016,N_7022,N_5877);
nand U8017 (N_8017,N_5982,N_5083);
xor U8018 (N_8018,N_7156,N_5526);
xnor U8019 (N_8019,N_5132,N_6785);
nor U8020 (N_8020,N_6168,N_6878);
nand U8021 (N_8021,N_6486,N_7261);
or U8022 (N_8022,N_5498,N_5149);
nor U8023 (N_8023,N_5211,N_6194);
xnor U8024 (N_8024,N_6720,N_5184);
and U8025 (N_8025,N_6914,N_6930);
nor U8026 (N_8026,N_6688,N_5583);
nor U8027 (N_8027,N_6344,N_7080);
xor U8028 (N_8028,N_5687,N_6671);
and U8029 (N_8029,N_5465,N_7295);
xnor U8030 (N_8030,N_5810,N_6608);
or U8031 (N_8031,N_6939,N_7350);
and U8032 (N_8032,N_7078,N_6750);
nor U8033 (N_8033,N_6213,N_6724);
nor U8034 (N_8034,N_5464,N_5404);
xor U8035 (N_8035,N_7457,N_6625);
xnor U8036 (N_8036,N_7181,N_7373);
nand U8037 (N_8037,N_6272,N_5194);
nor U8038 (N_8038,N_5017,N_5268);
or U8039 (N_8039,N_6530,N_6317);
nor U8040 (N_8040,N_6416,N_6856);
nor U8041 (N_8041,N_6307,N_5708);
xnor U8042 (N_8042,N_7367,N_5152);
or U8043 (N_8043,N_5288,N_7062);
nand U8044 (N_8044,N_5306,N_5977);
or U8045 (N_8045,N_7411,N_6790);
and U8046 (N_8046,N_6184,N_5659);
nand U8047 (N_8047,N_7340,N_6985);
or U8048 (N_8048,N_7070,N_7368);
nor U8049 (N_8049,N_5806,N_6407);
xnor U8050 (N_8050,N_6389,N_6732);
nor U8051 (N_8051,N_6577,N_7335);
xor U8052 (N_8052,N_6063,N_5080);
and U8053 (N_8053,N_6711,N_7293);
xnor U8054 (N_8054,N_6465,N_5282);
nor U8055 (N_8055,N_6580,N_7450);
or U8056 (N_8056,N_5634,N_7375);
and U8057 (N_8057,N_6848,N_6398);
xnor U8058 (N_8058,N_6612,N_7405);
xor U8059 (N_8059,N_7045,N_6556);
nand U8060 (N_8060,N_7435,N_6989);
or U8061 (N_8061,N_7358,N_6528);
or U8062 (N_8062,N_5402,N_5990);
or U8063 (N_8063,N_5785,N_6574);
xor U8064 (N_8064,N_6054,N_5339);
nand U8065 (N_8065,N_6181,N_5292);
nand U8066 (N_8066,N_5263,N_6739);
and U8067 (N_8067,N_6814,N_7444);
or U8068 (N_8068,N_6176,N_7074);
xnor U8069 (N_8069,N_5113,N_5839);
and U8070 (N_8070,N_6774,N_6089);
or U8071 (N_8071,N_5726,N_5294);
nand U8072 (N_8072,N_6011,N_6238);
nor U8073 (N_8073,N_5163,N_6110);
or U8074 (N_8074,N_6727,N_5125);
or U8075 (N_8075,N_6120,N_6123);
xor U8076 (N_8076,N_6472,N_7469);
xor U8077 (N_8077,N_6256,N_6386);
nand U8078 (N_8078,N_5065,N_5059);
or U8079 (N_8079,N_7486,N_5223);
and U8080 (N_8080,N_6610,N_7150);
or U8081 (N_8081,N_6522,N_6253);
or U8082 (N_8082,N_5698,N_6237);
and U8083 (N_8083,N_6838,N_5054);
nand U8084 (N_8084,N_7441,N_7333);
xnor U8085 (N_8085,N_7401,N_6836);
xnor U8086 (N_8086,N_6296,N_6565);
xor U8087 (N_8087,N_7234,N_5535);
nand U8088 (N_8088,N_6588,N_5086);
and U8089 (N_8089,N_5368,N_6038);
and U8090 (N_8090,N_6287,N_7005);
and U8091 (N_8091,N_6149,N_7247);
or U8092 (N_8092,N_5907,N_5544);
and U8093 (N_8093,N_5490,N_7103);
xor U8094 (N_8094,N_6725,N_5823);
or U8095 (N_8095,N_7013,N_7220);
xnor U8096 (N_8096,N_7453,N_5652);
and U8097 (N_8097,N_6239,N_7004);
and U8098 (N_8098,N_7075,N_5965);
and U8099 (N_8099,N_5277,N_7303);
nor U8100 (N_8100,N_6292,N_6660);
nand U8101 (N_8101,N_5596,N_7041);
and U8102 (N_8102,N_5285,N_6298);
or U8103 (N_8103,N_5433,N_6452);
or U8104 (N_8104,N_7008,N_5380);
nand U8105 (N_8105,N_6781,N_5678);
or U8106 (N_8106,N_7410,N_7033);
nand U8107 (N_8107,N_5168,N_5497);
and U8108 (N_8108,N_7185,N_7176);
nand U8109 (N_8109,N_6179,N_6466);
xnor U8110 (N_8110,N_6605,N_7130);
nand U8111 (N_8111,N_6909,N_5247);
nor U8112 (N_8112,N_5879,N_7374);
xnor U8113 (N_8113,N_6918,N_6112);
and U8114 (N_8114,N_6269,N_6430);
or U8115 (N_8115,N_6134,N_5469);
and U8116 (N_8116,N_5164,N_7282);
nand U8117 (N_8117,N_5496,N_7346);
nor U8118 (N_8118,N_5329,N_5528);
nor U8119 (N_8119,N_5357,N_5388);
and U8120 (N_8120,N_5038,N_6968);
nand U8121 (N_8121,N_6173,N_7451);
xor U8122 (N_8122,N_7031,N_5884);
nor U8123 (N_8123,N_5870,N_5930);
and U8124 (N_8124,N_5049,N_5297);
or U8125 (N_8125,N_6384,N_5331);
and U8126 (N_8126,N_6877,N_5969);
nand U8127 (N_8127,N_7488,N_5105);
nor U8128 (N_8128,N_5378,N_5066);
nor U8129 (N_8129,N_5629,N_7154);
xor U8130 (N_8130,N_6198,N_5715);
nor U8131 (N_8131,N_6755,N_5081);
xnor U8132 (N_8132,N_7035,N_5536);
xnor U8133 (N_8133,N_7257,N_7277);
nor U8134 (N_8134,N_6846,N_7330);
or U8135 (N_8135,N_5023,N_6917);
and U8136 (N_8136,N_6095,N_5645);
nor U8137 (N_8137,N_5479,N_6568);
nor U8138 (N_8138,N_5070,N_7148);
nor U8139 (N_8139,N_5958,N_7445);
and U8140 (N_8140,N_7417,N_6032);
nand U8141 (N_8141,N_5656,N_7244);
nand U8142 (N_8142,N_5486,N_5550);
xor U8143 (N_8143,N_6615,N_6281);
nor U8144 (N_8144,N_6741,N_7354);
or U8145 (N_8145,N_5355,N_6800);
nor U8146 (N_8146,N_6041,N_6280);
or U8147 (N_8147,N_5697,N_5021);
xnor U8148 (N_8148,N_5314,N_6881);
or U8149 (N_8149,N_6870,N_7325);
and U8150 (N_8150,N_5909,N_5322);
and U8151 (N_8151,N_5111,N_5758);
xor U8152 (N_8152,N_7057,N_6075);
nand U8153 (N_8153,N_7496,N_6598);
nand U8154 (N_8154,N_5360,N_7170);
and U8155 (N_8155,N_6882,N_6872);
xnor U8156 (N_8156,N_7280,N_5689);
nand U8157 (N_8157,N_6706,N_6111);
xnor U8158 (N_8158,N_6596,N_5271);
xnor U8159 (N_8159,N_7492,N_7141);
nand U8160 (N_8160,N_5197,N_5517);
xnor U8161 (N_8161,N_5607,N_7058);
xor U8162 (N_8162,N_5817,N_5182);
and U8163 (N_8163,N_6067,N_6066);
and U8164 (N_8164,N_7302,N_7328);
or U8165 (N_8165,N_7385,N_5628);
or U8166 (N_8166,N_5151,N_6474);
nor U8167 (N_8167,N_6912,N_7047);
or U8168 (N_8168,N_5774,N_5959);
xor U8169 (N_8169,N_6733,N_5975);
or U8170 (N_8170,N_7369,N_6369);
nor U8171 (N_8171,N_5873,N_6549);
nor U8172 (N_8172,N_6973,N_7151);
nand U8173 (N_8173,N_6189,N_5796);
xor U8174 (N_8174,N_5140,N_5188);
nand U8175 (N_8175,N_5349,N_5252);
nand U8176 (N_8176,N_5621,N_5390);
xnor U8177 (N_8177,N_5978,N_6784);
nand U8178 (N_8178,N_5224,N_6295);
nand U8179 (N_8179,N_5878,N_6448);
or U8180 (N_8180,N_6777,N_7429);
or U8181 (N_8181,N_6513,N_7192);
nor U8182 (N_8182,N_6746,N_6458);
xnor U8183 (N_8183,N_6165,N_6409);
nor U8184 (N_8184,N_6500,N_6942);
xor U8185 (N_8185,N_5863,N_5529);
nor U8186 (N_8186,N_5275,N_6536);
nor U8187 (N_8187,N_6512,N_6250);
nor U8188 (N_8188,N_6100,N_5857);
xor U8189 (N_8189,N_5064,N_7046);
or U8190 (N_8190,N_6766,N_6226);
nor U8191 (N_8191,N_6055,N_6787);
xor U8192 (N_8192,N_6521,N_7265);
and U8193 (N_8193,N_6385,N_6433);
xnor U8194 (N_8194,N_5504,N_5800);
or U8195 (N_8195,N_5240,N_5951);
nand U8196 (N_8196,N_5552,N_6754);
nand U8197 (N_8197,N_5299,N_5953);
and U8198 (N_8198,N_7119,N_6412);
xor U8199 (N_8199,N_5382,N_6374);
nand U8200 (N_8200,N_5226,N_5524);
nand U8201 (N_8201,N_5310,N_5270);
and U8202 (N_8202,N_5564,N_5569);
xor U8203 (N_8203,N_6672,N_6734);
nor U8204 (N_8204,N_6783,N_6357);
nand U8205 (N_8205,N_6048,N_6103);
or U8206 (N_8206,N_6964,N_7199);
nand U8207 (N_8207,N_6583,N_6949);
nor U8208 (N_8208,N_6345,N_7028);
nand U8209 (N_8209,N_6796,N_6129);
and U8210 (N_8210,N_6082,N_7118);
nand U8211 (N_8211,N_5510,N_5358);
nand U8212 (N_8212,N_5216,N_6172);
or U8213 (N_8213,N_5553,N_6336);
xor U8214 (N_8214,N_5187,N_5012);
nor U8215 (N_8215,N_5976,N_7054);
or U8216 (N_8216,N_7413,N_6518);
nand U8217 (N_8217,N_5935,N_6051);
nand U8218 (N_8218,N_5631,N_6309);
and U8219 (N_8219,N_7424,N_5812);
and U8220 (N_8220,N_7178,N_5933);
nor U8221 (N_8221,N_5869,N_6970);
and U8222 (N_8222,N_6487,N_7064);
and U8223 (N_8223,N_7134,N_6935);
nor U8224 (N_8224,N_7371,N_7207);
or U8225 (N_8225,N_5750,N_6695);
or U8226 (N_8226,N_6347,N_7422);
or U8227 (N_8227,N_5558,N_7345);
nor U8228 (N_8228,N_5798,N_5336);
nor U8229 (N_8229,N_5118,N_5319);
nor U8230 (N_8230,N_5098,N_5112);
and U8231 (N_8231,N_6383,N_6456);
xnor U8232 (N_8232,N_6545,N_5567);
or U8233 (N_8233,N_6002,N_6694);
or U8234 (N_8234,N_5009,N_5481);
or U8235 (N_8235,N_6798,N_5308);
and U8236 (N_8236,N_5385,N_6358);
or U8237 (N_8237,N_6321,N_5335);
xor U8238 (N_8238,N_5468,N_6879);
nand U8239 (N_8239,N_5148,N_5426);
and U8240 (N_8240,N_5144,N_6410);
xnor U8241 (N_8241,N_6764,N_6745);
nand U8242 (N_8242,N_6662,N_5650);
nor U8243 (N_8243,N_5679,N_5866);
and U8244 (N_8244,N_7238,N_7077);
xor U8245 (N_8245,N_5905,N_5891);
and U8246 (N_8246,N_5540,N_7136);
xor U8247 (N_8247,N_6312,N_5456);
and U8248 (N_8248,N_7263,N_5657);
or U8249 (N_8249,N_5757,N_6018);
xnor U8250 (N_8250,N_6020,N_7036);
xor U8251 (N_8251,N_5041,N_7183);
nand U8252 (N_8252,N_5076,N_6300);
and U8253 (N_8253,N_7305,N_6397);
nor U8254 (N_8254,N_5571,N_5185);
and U8255 (N_8255,N_7042,N_5575);
nand U8256 (N_8256,N_6630,N_6275);
or U8257 (N_8257,N_7279,N_5068);
nor U8258 (N_8258,N_5033,N_6890);
xor U8259 (N_8259,N_5254,N_6365);
xor U8260 (N_8260,N_7275,N_6618);
or U8261 (N_8261,N_6983,N_5022);
nor U8262 (N_8262,N_6230,N_5818);
and U8263 (N_8263,N_6186,N_6366);
nand U8264 (N_8264,N_6753,N_6699);
or U8265 (N_8265,N_7260,N_5085);
xnor U8266 (N_8266,N_6150,N_7120);
and U8267 (N_8267,N_6263,N_6241);
and U8268 (N_8268,N_5705,N_7087);
or U8269 (N_8269,N_6147,N_5352);
or U8270 (N_8270,N_7160,N_5892);
or U8271 (N_8271,N_6178,N_5220);
and U8272 (N_8272,N_6140,N_6304);
xnor U8273 (N_8273,N_6290,N_5154);
nor U8274 (N_8274,N_7355,N_5651);
nand U8275 (N_8275,N_5648,N_6897);
xnor U8276 (N_8276,N_6490,N_6161);
and U8277 (N_8277,N_6936,N_6972);
and U8278 (N_8278,N_7203,N_7024);
or U8279 (N_8279,N_5264,N_6809);
nand U8280 (N_8280,N_6105,N_5921);
xor U8281 (N_8281,N_6693,N_6861);
or U8282 (N_8282,N_6718,N_6923);
nor U8283 (N_8283,N_5407,N_7173);
nand U8284 (N_8284,N_6794,N_7359);
and U8285 (N_8285,N_5968,N_7111);
nand U8286 (N_8286,N_7175,N_6306);
xor U8287 (N_8287,N_6589,N_5888);
nor U8288 (N_8288,N_6008,N_5417);
xor U8289 (N_8289,N_5475,N_5274);
nor U8290 (N_8290,N_5376,N_5593);
or U8291 (N_8291,N_7297,N_5696);
and U8292 (N_8292,N_5770,N_7132);
nor U8293 (N_8293,N_6214,N_6001);
nor U8294 (N_8294,N_6124,N_5414);
nor U8295 (N_8295,N_6274,N_5709);
xnor U8296 (N_8296,N_6010,N_5405);
or U8297 (N_8297,N_5939,N_5090);
nand U8298 (N_8298,N_6484,N_6515);
nand U8299 (N_8299,N_5457,N_5914);
or U8300 (N_8300,N_6346,N_7245);
nor U8301 (N_8301,N_6959,N_7066);
nand U8302 (N_8302,N_6859,N_6299);
xor U8303 (N_8303,N_6552,N_5609);
nand U8304 (N_8304,N_5980,N_5831);
nor U8305 (N_8305,N_7237,N_5156);
xnor U8306 (N_8306,N_7362,N_5527);
and U8307 (N_8307,N_6937,N_5095);
xnor U8308 (N_8308,N_5807,N_6622);
xnor U8309 (N_8309,N_6343,N_6855);
nand U8310 (N_8310,N_7498,N_6895);
and U8311 (N_8311,N_7198,N_6439);
and U8312 (N_8312,N_6056,N_6016);
or U8313 (N_8313,N_5363,N_6445);
or U8314 (N_8314,N_5403,N_6597);
and U8315 (N_8315,N_6212,N_5627);
xor U8316 (N_8316,N_7420,N_5728);
or U8317 (N_8317,N_5676,N_5537);
and U8318 (N_8318,N_7172,N_6209);
and U8319 (N_8319,N_6349,N_5191);
xor U8320 (N_8320,N_6759,N_7083);
nand U8321 (N_8321,N_6591,N_5499);
nand U8322 (N_8322,N_6998,N_6956);
xor U8323 (N_8323,N_5482,N_6203);
and U8324 (N_8324,N_6950,N_6818);
xnor U8325 (N_8325,N_5487,N_5317);
xor U8326 (N_8326,N_6328,N_5612);
xor U8327 (N_8327,N_7095,N_7364);
nand U8328 (N_8328,N_6875,N_5207);
and U8329 (N_8329,N_7443,N_6132);
and U8330 (N_8330,N_7196,N_6091);
nor U8331 (N_8331,N_6958,N_5234);
xor U8332 (N_8332,N_5466,N_7089);
and U8333 (N_8333,N_7214,N_6126);
and U8334 (N_8334,N_6849,N_5927);
or U8335 (N_8335,N_5203,N_5512);
nand U8336 (N_8336,N_6160,N_5272);
nor U8337 (N_8337,N_5300,N_6128);
nand U8338 (N_8338,N_5383,N_5765);
and U8339 (N_8339,N_5147,N_7455);
nor U8340 (N_8340,N_5323,N_5635);
nor U8341 (N_8341,N_7400,N_5032);
and U8342 (N_8342,N_5922,N_5681);
nor U8343 (N_8343,N_5711,N_5622);
and U8344 (N_8344,N_7456,N_7476);
and U8345 (N_8345,N_5749,N_6907);
and U8346 (N_8346,N_5736,N_5960);
xor U8347 (N_8347,N_6167,N_5996);
or U8348 (N_8348,N_7288,N_6437);
or U8349 (N_8349,N_5600,N_6684);
or U8350 (N_8350,N_6233,N_7230);
nor U8351 (N_8351,N_6744,N_7110);
nor U8352 (N_8352,N_6114,N_5835);
and U8353 (N_8353,N_7285,N_7497);
nor U8354 (N_8354,N_6478,N_5623);
nor U8355 (N_8355,N_5713,N_7309);
xnor U8356 (N_8356,N_6501,N_6285);
and U8357 (N_8357,N_6569,N_6984);
xor U8358 (N_8358,N_6086,N_5053);
xor U8359 (N_8359,N_5062,N_6629);
and U8360 (N_8360,N_5397,N_6191);
and U8361 (N_8361,N_6858,N_5337);
xor U8362 (N_8362,N_5586,N_5222);
or U8363 (N_8363,N_6392,N_6634);
nor U8364 (N_8364,N_5242,N_5025);
or U8365 (N_8365,N_5707,N_6758);
or U8366 (N_8366,N_6455,N_5181);
and U8367 (N_8367,N_7210,N_5752);
or U8368 (N_8368,N_7438,N_5895);
nand U8369 (N_8369,N_6446,N_7026);
or U8370 (N_8370,N_6541,N_7152);
and U8371 (N_8371,N_7310,N_6164);
xor U8372 (N_8372,N_5327,N_5641);
xnor U8373 (N_8373,N_5346,N_7478);
and U8374 (N_8374,N_5259,N_6043);
or U8375 (N_8375,N_6899,N_7072);
and U8376 (N_8376,N_6641,N_5078);
and U8377 (N_8377,N_5780,N_5048);
or U8378 (N_8378,N_5326,N_5293);
nor U8379 (N_8379,N_5117,N_5225);
and U8380 (N_8380,N_5562,N_5759);
xor U8381 (N_8381,N_6869,N_5644);
nand U8382 (N_8382,N_5636,N_5267);
nor U8383 (N_8383,N_5050,N_5443);
and U8384 (N_8384,N_5813,N_6243);
and U8385 (N_8385,N_5853,N_5936);
or U8386 (N_8386,N_5392,N_7106);
xor U8387 (N_8387,N_6449,N_6633);
xor U8388 (N_8388,N_6673,N_7467);
or U8389 (N_8389,N_6029,N_6205);
nor U8390 (N_8390,N_5139,N_7000);
or U8391 (N_8391,N_5945,N_5745);
nand U8392 (N_8392,N_5205,N_5201);
nand U8393 (N_8393,N_6069,N_6982);
or U8394 (N_8394,N_6000,N_6919);
or U8395 (N_8395,N_6236,N_6990);
nor U8396 (N_8396,N_6977,N_7425);
nand U8397 (N_8397,N_7363,N_6323);
xnor U8398 (N_8398,N_7113,N_6651);
nor U8399 (N_8399,N_7149,N_7406);
nand U8400 (N_8400,N_6022,N_6685);
or U8401 (N_8401,N_6030,N_6883);
nand U8402 (N_8402,N_5700,N_5169);
and U8403 (N_8403,N_7494,N_7167);
xnor U8404 (N_8404,N_6251,N_5459);
nor U8405 (N_8405,N_6854,N_5762);
and U8406 (N_8406,N_6925,N_6380);
and U8407 (N_8407,N_5738,N_6319);
and U8408 (N_8408,N_5579,N_5442);
and U8409 (N_8409,N_6065,N_7397);
nand U8410 (N_8410,N_5502,N_7336);
nand U8411 (N_8411,N_7485,N_6480);
xor U8412 (N_8412,N_6847,N_6282);
and U8413 (N_8413,N_6687,N_6548);
xor U8414 (N_8414,N_6645,N_5743);
and U8415 (N_8415,N_5313,N_5256);
nor U8416 (N_8416,N_6145,N_5186);
nand U8417 (N_8417,N_5625,N_6424);
xnor U8418 (N_8418,N_5401,N_5051);
and U8419 (N_8419,N_5804,N_7189);
nor U8420 (N_8420,N_6511,N_5747);
or U8421 (N_8421,N_7145,N_5530);
nand U8422 (N_8422,N_7222,N_5920);
xnor U8423 (N_8423,N_6537,N_5766);
nor U8424 (N_8424,N_6988,N_5513);
nand U8425 (N_8425,N_6053,N_6322);
or U8426 (N_8426,N_5925,N_6081);
nor U8427 (N_8427,N_5503,N_7017);
nor U8428 (N_8428,N_5158,N_7112);
nor U8429 (N_8429,N_5321,N_6028);
or U8430 (N_8430,N_7014,N_6572);
nor U8431 (N_8431,N_5471,N_5445);
xor U8432 (N_8432,N_6097,N_6997);
xor U8433 (N_8433,N_5374,N_5193);
xor U8434 (N_8434,N_7404,N_7393);
nand U8435 (N_8435,N_5809,N_5100);
or U8436 (N_8436,N_6810,N_6305);
xnor U8437 (N_8437,N_7311,N_5658);
nand U8438 (N_8438,N_6797,N_7076);
nand U8439 (N_8439,N_6637,N_5246);
xor U8440 (N_8440,N_6691,N_5999);
and U8441 (N_8441,N_5966,N_6707);
or U8442 (N_8442,N_7255,N_5219);
nor U8443 (N_8443,N_6098,N_5667);
nor U8444 (N_8444,N_5514,N_7284);
nand U8445 (N_8445,N_5746,N_6507);
and U8446 (N_8446,N_7159,N_7319);
and U8447 (N_8447,N_7079,N_6496);
and U8448 (N_8448,N_7063,N_5235);
nand U8449 (N_8449,N_5393,N_5356);
and U8450 (N_8450,N_5756,N_5280);
nand U8451 (N_8451,N_5435,N_5993);
and U8452 (N_8452,N_7050,N_7109);
xnor U8453 (N_8453,N_6005,N_6102);
xnor U8454 (N_8454,N_6231,N_6540);
xor U8455 (N_8455,N_6664,N_6014);
xor U8456 (N_8456,N_6624,N_6060);
nand U8457 (N_8457,N_7296,N_6544);
nand U8458 (N_8458,N_7433,N_6438);
nand U8459 (N_8459,N_5516,N_7250);
nor U8460 (N_8460,N_5167,N_7357);
nand U8461 (N_8461,N_5735,N_6376);
nor U8462 (N_8462,N_6941,N_7332);
xnor U8463 (N_8463,N_6926,N_5938);
nand U8464 (N_8464,N_7462,N_5668);
or U8465 (N_8465,N_6050,N_6260);
nand U8466 (N_8466,N_6752,N_6297);
nor U8467 (N_8467,N_5574,N_5141);
and U8468 (N_8468,N_6405,N_5701);
nor U8469 (N_8469,N_5775,N_7227);
nand U8470 (N_8470,N_5699,N_6538);
xnor U8471 (N_8471,N_6590,N_6957);
nand U8472 (N_8472,N_6771,N_5037);
or U8473 (N_8473,N_6826,N_7452);
nand U8474 (N_8474,N_7186,N_7212);
or U8475 (N_8475,N_6155,N_6980);
nor U8476 (N_8476,N_7125,N_5859);
nor U8477 (N_8477,N_6308,N_6216);
xnor U8478 (N_8478,N_6266,N_6786);
nand U8479 (N_8479,N_6169,N_7344);
or U8480 (N_8480,N_7389,N_5162);
and U8481 (N_8481,N_6481,N_6498);
nand U8482 (N_8482,N_6729,N_7307);
and U8483 (N_8483,N_6348,N_6316);
and U8484 (N_8484,N_6443,N_7158);
nor U8485 (N_8485,N_7209,N_7122);
nand U8486 (N_8486,N_6782,N_6463);
or U8487 (N_8487,N_5014,N_7353);
xnor U8488 (N_8488,N_5518,N_6039);
nand U8489 (N_8489,N_6888,N_6413);
nand U8490 (N_8490,N_6966,N_6703);
nand U8491 (N_8491,N_6373,N_5511);
xnor U8492 (N_8492,N_6539,N_6974);
xor U8493 (N_8493,N_6252,N_6227);
xor U8494 (N_8494,N_5476,N_7414);
and U8495 (N_8495,N_7430,N_7190);
nand U8496 (N_8496,N_5324,N_5493);
and U8497 (N_8497,N_5955,N_6534);
and U8498 (N_8498,N_5446,N_7034);
and U8499 (N_8499,N_6142,N_6087);
or U8500 (N_8500,N_6450,N_7292);
nor U8501 (N_8501,N_7273,N_7402);
xor U8502 (N_8502,N_5005,N_6567);
nor U8503 (N_8503,N_5677,N_5075);
or U8504 (N_8504,N_5101,N_5228);
or U8505 (N_8505,N_6471,N_6689);
xor U8506 (N_8506,N_5833,N_7094);
and U8507 (N_8507,N_5377,N_6736);
nand U8508 (N_8508,N_5573,N_5932);
xor U8509 (N_8509,N_5008,N_6901);
and U8510 (N_8510,N_6331,N_7448);
and U8511 (N_8511,N_6659,N_5821);
xor U8512 (N_8512,N_6432,N_6162);
nand U8513 (N_8513,N_6792,N_6199);
nand U8514 (N_8514,N_5929,N_7161);
and U8515 (N_8515,N_6700,N_7060);
nor U8516 (N_8516,N_5089,N_6976);
xnor U8517 (N_8517,N_6485,N_7299);
xnor U8518 (N_8518,N_5808,N_6370);
or U8519 (N_8519,N_6947,N_5016);
nand U8520 (N_8520,N_7366,N_5741);
nand U8521 (N_8521,N_5721,N_6166);
or U8522 (N_8522,N_5694,N_5379);
or U8523 (N_8523,N_5146,N_6031);
nor U8524 (N_8524,N_5719,N_5422);
and U8525 (N_8525,N_6932,N_6683);
nor U8526 (N_8526,N_7166,N_6851);
and U8527 (N_8527,N_6502,N_7193);
xor U8528 (N_8528,N_5662,N_6905);
and U8529 (N_8529,N_6915,N_6827);
nand U8530 (N_8530,N_5494,N_6931);
and U8531 (N_8531,N_6271,N_6526);
nor U8532 (N_8532,N_5245,N_5767);
nand U8533 (N_8533,N_6188,N_6351);
and U8534 (N_8534,N_6286,N_5108);
nand U8535 (N_8535,N_6363,N_5315);
and U8536 (N_8536,N_5781,N_6708);
xnor U8537 (N_8537,N_5985,N_6076);
nor U8538 (N_8538,N_5501,N_5036);
nor U8539 (N_8539,N_5772,N_7128);
and U8540 (N_8540,N_6387,N_5695);
or U8541 (N_8541,N_5332,N_6807);
nand U8542 (N_8542,N_6920,N_6529);
or U8543 (N_8543,N_6426,N_7236);
or U8544 (N_8544,N_6586,N_6473);
and U8545 (N_8545,N_6248,N_5603);
xnor U8546 (N_8546,N_6701,N_6396);
and U8547 (N_8547,N_5345,N_5367);
or U8548 (N_8548,N_5974,N_5287);
and U8549 (N_8549,N_5366,N_7037);
nor U8550 (N_8550,N_6658,N_5227);
nor U8551 (N_8551,N_7165,N_5097);
and U8552 (N_8552,N_6049,N_5178);
xnor U8553 (N_8553,N_5793,N_7051);
or U8554 (N_8554,N_5143,N_6692);
xor U8555 (N_8555,N_5852,N_5190);
nor U8556 (N_8556,N_5439,N_6868);
nor U8557 (N_8557,N_5533,N_5903);
nand U8558 (N_8558,N_6283,N_7093);
or U8559 (N_8559,N_6837,N_5598);
or U8560 (N_8560,N_7067,N_5491);
nor U8561 (N_8561,N_5580,N_5789);
or U8562 (N_8562,N_5408,N_5421);
and U8563 (N_8563,N_6678,N_6661);
nor U8564 (N_8564,N_6900,N_5838);
and U8565 (N_8565,N_6218,N_7314);
and U8566 (N_8566,N_5970,N_5559);
or U8567 (N_8567,N_5432,N_5926);
nor U8568 (N_8568,N_5029,N_7383);
nand U8569 (N_8569,N_6177,N_5217);
and U8570 (N_8570,N_6052,N_5858);
and U8571 (N_8571,N_7276,N_5545);
nand U8572 (N_8572,N_6046,N_7086);
nand U8573 (N_8573,N_6012,N_6084);
and U8574 (N_8574,N_7061,N_7071);
xor U8575 (N_8575,N_6406,N_5820);
or U8576 (N_8576,N_5919,N_6709);
xor U8577 (N_8577,N_6874,N_6314);
nand U8578 (N_8578,N_6986,N_6401);
nor U8579 (N_8579,N_5106,N_7382);
xnor U8580 (N_8580,N_5717,N_7228);
and U8581 (N_8581,N_5229,N_6355);
and U8582 (N_8582,N_6262,N_5069);
and U8583 (N_8583,N_6497,N_5716);
nand U8584 (N_8584,N_5450,N_5467);
and U8585 (N_8585,N_5685,N_6361);
nor U8586 (N_8586,N_6059,N_6378);
nor U8587 (N_8587,N_6987,N_7318);
nand U8588 (N_8588,N_5844,N_6004);
and U8589 (N_8589,N_6330,N_6261);
or U8590 (N_8590,N_5004,N_5386);
or U8591 (N_8591,N_5619,N_6722);
xnor U8592 (N_8592,N_7204,N_5940);
nand U8593 (N_8593,N_7030,N_5344);
nand U8594 (N_8594,N_5740,N_5209);
or U8595 (N_8595,N_5127,N_6185);
nand U8596 (N_8596,N_7320,N_7493);
xnor U8597 (N_8597,N_5214,N_5952);
nand U8598 (N_8598,N_5341,N_6619);
or U8599 (N_8599,N_5734,N_6372);
nand U8600 (N_8600,N_7495,N_6546);
xnor U8601 (N_8601,N_7326,N_5210);
nand U8602 (N_8602,N_5372,N_5172);
xnor U8603 (N_8603,N_5159,N_6799);
nor U8604 (N_8604,N_7019,N_7304);
nor U8605 (N_8605,N_5584,N_5359);
nand U8606 (N_8606,N_5915,N_5943);
nand U8607 (N_8607,N_6885,N_5840);
or U8608 (N_8608,N_6415,N_7009);
and U8609 (N_8609,N_5251,N_6600);
nand U8610 (N_8610,N_6564,N_5353);
or U8611 (N_8611,N_5618,N_5434);
and U8612 (N_8612,N_6581,N_6929);
nand U8613 (N_8613,N_5832,N_7323);
or U8614 (N_8614,N_5145,N_7043);
nor U8615 (N_8615,N_5850,N_5237);
or U8616 (N_8616,N_7324,N_6088);
and U8617 (N_8617,N_6470,N_5589);
and U8618 (N_8618,N_5688,N_6726);
or U8619 (N_8619,N_7195,N_7331);
xor U8620 (N_8620,N_7409,N_6738);
nand U8621 (N_8621,N_6894,N_5134);
and U8622 (N_8622,N_6675,N_6183);
or U8623 (N_8623,N_6244,N_5592);
and U8624 (N_8624,N_6509,N_5241);
xnor U8625 (N_8625,N_5195,N_6215);
xor U8626 (N_8626,N_6532,N_5500);
xnor U8627 (N_8627,N_6121,N_5507);
xnor U8628 (N_8628,N_6514,N_6627);
nor U8629 (N_8629,N_6601,N_7322);
or U8630 (N_8630,N_5557,N_5046);
xnor U8631 (N_8631,N_6232,N_5595);
and U8632 (N_8632,N_6006,N_7065);
nand U8633 (N_8633,N_6554,N_5419);
nand U8634 (N_8634,N_5893,N_6293);
and U8635 (N_8635,N_5582,N_5549);
xor U8636 (N_8636,N_6705,N_5730);
nor U8637 (N_8637,N_7133,N_6163);
nand U8638 (N_8638,N_5950,N_6493);
or U8639 (N_8639,N_5588,N_6767);
nand U8640 (N_8640,N_7107,N_5843);
and U8641 (N_8641,N_6751,N_5423);
nor U8642 (N_8642,N_6582,N_6270);
nor U8643 (N_8643,N_5045,N_6411);
and U8644 (N_8644,N_6024,N_6516);
or U8645 (N_8645,N_7312,N_7264);
nor U8646 (N_8646,N_5754,N_7219);
nor U8647 (N_8647,N_6259,N_5531);
or U8648 (N_8648,N_6315,N_5654);
and U8649 (N_8649,N_5286,N_6034);
nor U8650 (N_8650,N_7044,N_5984);
and U8651 (N_8651,N_6381,N_7117);
or U8652 (N_8652,N_5221,N_6276);
or U8653 (N_8653,N_6592,N_6993);
nand U8654 (N_8654,N_5394,N_7129);
xnor U8655 (N_8655,N_6808,N_5058);
and U8656 (N_8656,N_7040,N_5473);
and U8657 (N_8657,N_5570,N_6190);
nor U8658 (N_8658,N_5249,N_6978);
nand U8659 (N_8659,N_6267,N_6547);
or U8660 (N_8660,N_7470,N_7384);
nand U8661 (N_8661,N_6073,N_5495);
nand U8662 (N_8662,N_6210,N_6420);
xnor U8663 (N_8663,N_7466,N_5680);
or U8664 (N_8664,N_5093,N_7407);
nand U8665 (N_8665,N_5638,N_7294);
and U8666 (N_8666,N_6242,N_7163);
nand U8667 (N_8667,N_5578,N_7188);
or U8668 (N_8668,N_6953,N_6106);
xor U8669 (N_8669,N_5822,N_7308);
and U8670 (N_8670,N_6180,N_6593);
nand U8671 (N_8671,N_7021,N_5771);
and U8672 (N_8672,N_5795,N_6523);
nor U8673 (N_8673,N_7137,N_5365);
nor U8674 (N_8674,N_5898,N_5604);
and U8675 (N_8675,N_6353,N_6607);
or U8676 (N_8676,N_7481,N_5783);
nand U8677 (N_8677,N_5124,N_5753);
nor U8678 (N_8678,N_5460,N_5074);
and U8679 (N_8679,N_5995,N_5674);
xnor U8680 (N_8680,N_5664,N_5837);
xor U8681 (N_8681,N_5617,N_7239);
or U8682 (N_8682,N_6623,N_5133);
and U8683 (N_8683,N_6255,N_5213);
and U8684 (N_8684,N_6811,N_6995);
nor U8685 (N_8685,N_6575,N_5624);
nand U8686 (N_8686,N_6626,N_7029);
nor U8687 (N_8687,N_5396,N_6219);
or U8688 (N_8688,N_7269,N_6763);
xor U8689 (N_8689,N_5702,N_7213);
nand U8690 (N_8690,N_5082,N_6922);
nand U8691 (N_8691,N_7242,N_5381);
nor U8692 (N_8692,N_5411,N_7316);
nand U8693 (N_8693,N_7241,N_6910);
xnor U8694 (N_8694,N_5543,N_5415);
xor U8695 (N_8695,N_5485,N_6133);
nand U8696 (N_8696,N_5555,N_6649);
nand U8697 (N_8697,N_6479,N_5748);
or U8698 (N_8698,N_6342,N_5055);
or U8699 (N_8699,N_6640,N_5712);
xnor U8700 (N_8700,N_5320,N_6578);
nand U8701 (N_8701,N_6277,N_5896);
and U8702 (N_8702,N_7018,N_5384);
xnor U8703 (N_8703,N_6819,N_6749);
or U8704 (N_8704,N_5655,N_5811);
nor U8705 (N_8705,N_6117,N_6143);
or U8706 (N_8706,N_5546,N_6820);
nand U8707 (N_8707,N_5847,N_6462);
nand U8708 (N_8708,N_5369,N_7099);
xor U8709 (N_8709,N_7191,N_5601);
or U8710 (N_8710,N_6825,N_6096);
and U8711 (N_8711,N_5988,N_7392);
xnor U8712 (N_8712,N_7254,N_6553);
nor U8713 (N_8713,N_5534,N_6504);
nand U8714 (N_8714,N_5056,N_7164);
or U8715 (N_8715,N_7010,N_5991);
or U8716 (N_8716,N_7390,N_7153);
or U8717 (N_8717,N_5670,N_6525);
nand U8718 (N_8718,N_7262,N_5362);
xor U8719 (N_8719,N_6788,N_5706);
nand U8720 (N_8720,N_6613,N_5318);
xnor U8721 (N_8721,N_5761,N_5797);
xnor U8722 (N_8722,N_6517,N_7027);
and U8723 (N_8723,N_5954,N_5138);
nor U8724 (N_8724,N_6206,N_5846);
nand U8725 (N_8725,N_7121,N_6873);
and U8726 (N_8726,N_7338,N_6058);
and U8727 (N_8727,N_7049,N_7356);
or U8728 (N_8728,N_6494,N_5522);
nand U8729 (N_8729,N_7253,N_5554);
and U8730 (N_8730,N_6201,N_5290);
nor U8731 (N_8731,N_6454,N_6584);
and U8732 (N_8732,N_6551,N_5737);
and U8733 (N_8733,N_7454,N_6074);
and U8734 (N_8734,N_6863,N_5998);
or U8735 (N_8735,N_7258,N_6131);
nand U8736 (N_8736,N_5928,N_5942);
or U8737 (N_8737,N_6779,N_6367);
nand U8738 (N_8738,N_6085,N_6852);
xnor U8739 (N_8739,N_6273,N_5000);
nand U8740 (N_8740,N_6817,N_6246);
nand U8741 (N_8741,N_6730,N_5908);
and U8742 (N_8742,N_5956,N_5916);
xnor U8743 (N_8743,N_5425,N_6876);
and U8744 (N_8744,N_5581,N_5560);
or U8745 (N_8745,N_6775,N_5519);
nor U8746 (N_8746,N_6778,N_6801);
and U8747 (N_8747,N_6955,N_5109);
xnor U8748 (N_8748,N_5238,N_7206);
and U8749 (N_8749,N_6419,N_7147);
or U8750 (N_8750,N_5878,N_7387);
and U8751 (N_8751,N_7309,N_7304);
and U8752 (N_8752,N_7458,N_7144);
and U8753 (N_8753,N_5865,N_5471);
nand U8754 (N_8754,N_6149,N_5436);
nand U8755 (N_8755,N_5219,N_6712);
nor U8756 (N_8756,N_7319,N_5179);
nand U8757 (N_8757,N_5316,N_7317);
xnor U8758 (N_8758,N_7418,N_5496);
xor U8759 (N_8759,N_6724,N_6209);
nand U8760 (N_8760,N_5775,N_6472);
and U8761 (N_8761,N_5998,N_6188);
nand U8762 (N_8762,N_5667,N_6652);
or U8763 (N_8763,N_7307,N_6466);
nor U8764 (N_8764,N_6102,N_5007);
nand U8765 (N_8765,N_6815,N_6470);
nor U8766 (N_8766,N_6548,N_6849);
nand U8767 (N_8767,N_5210,N_6112);
xor U8768 (N_8768,N_6978,N_5459);
or U8769 (N_8769,N_7392,N_5211);
nand U8770 (N_8770,N_6225,N_6063);
nand U8771 (N_8771,N_6365,N_6632);
nand U8772 (N_8772,N_7338,N_6047);
and U8773 (N_8773,N_6956,N_7414);
nor U8774 (N_8774,N_7190,N_5447);
nor U8775 (N_8775,N_6288,N_6366);
or U8776 (N_8776,N_6358,N_7077);
and U8777 (N_8777,N_6919,N_6741);
nor U8778 (N_8778,N_5932,N_6407);
or U8779 (N_8779,N_5159,N_6687);
nor U8780 (N_8780,N_5267,N_7391);
nor U8781 (N_8781,N_7467,N_6503);
xor U8782 (N_8782,N_5891,N_6221);
nor U8783 (N_8783,N_5553,N_7275);
nand U8784 (N_8784,N_5804,N_5426);
nor U8785 (N_8785,N_6479,N_5714);
and U8786 (N_8786,N_6775,N_5074);
nor U8787 (N_8787,N_6509,N_6589);
or U8788 (N_8788,N_6102,N_6341);
nor U8789 (N_8789,N_6709,N_7218);
xor U8790 (N_8790,N_6358,N_6389);
nor U8791 (N_8791,N_6968,N_5193);
or U8792 (N_8792,N_7409,N_7283);
or U8793 (N_8793,N_7298,N_7299);
or U8794 (N_8794,N_7175,N_7249);
xnor U8795 (N_8795,N_6925,N_6462);
and U8796 (N_8796,N_5454,N_7419);
xnor U8797 (N_8797,N_7488,N_5258);
xor U8798 (N_8798,N_5334,N_5704);
nor U8799 (N_8799,N_6906,N_6919);
xnor U8800 (N_8800,N_5991,N_7456);
or U8801 (N_8801,N_6081,N_5915);
nand U8802 (N_8802,N_5877,N_6018);
or U8803 (N_8803,N_7291,N_5320);
xor U8804 (N_8804,N_5212,N_7219);
xor U8805 (N_8805,N_5060,N_6321);
nor U8806 (N_8806,N_6802,N_7415);
nand U8807 (N_8807,N_5006,N_6462);
or U8808 (N_8808,N_5307,N_7128);
xor U8809 (N_8809,N_6542,N_6775);
nor U8810 (N_8810,N_6738,N_6032);
nand U8811 (N_8811,N_7411,N_5849);
and U8812 (N_8812,N_7150,N_5936);
nor U8813 (N_8813,N_7443,N_5376);
or U8814 (N_8814,N_6051,N_7126);
nand U8815 (N_8815,N_6623,N_7302);
nand U8816 (N_8816,N_7301,N_5328);
nand U8817 (N_8817,N_6539,N_7166);
and U8818 (N_8818,N_5371,N_6808);
xnor U8819 (N_8819,N_5455,N_5218);
xnor U8820 (N_8820,N_5100,N_5736);
and U8821 (N_8821,N_7240,N_6364);
and U8822 (N_8822,N_5409,N_5228);
nand U8823 (N_8823,N_5439,N_6250);
and U8824 (N_8824,N_7439,N_7044);
nor U8825 (N_8825,N_5385,N_6303);
or U8826 (N_8826,N_5674,N_5067);
or U8827 (N_8827,N_6710,N_6436);
nor U8828 (N_8828,N_6554,N_5915);
xor U8829 (N_8829,N_5723,N_5630);
nor U8830 (N_8830,N_5710,N_6951);
or U8831 (N_8831,N_7144,N_6294);
and U8832 (N_8832,N_6709,N_6363);
nand U8833 (N_8833,N_6036,N_6467);
and U8834 (N_8834,N_7173,N_6097);
nand U8835 (N_8835,N_5578,N_5446);
xor U8836 (N_8836,N_7006,N_5788);
and U8837 (N_8837,N_7140,N_6172);
nand U8838 (N_8838,N_5642,N_7268);
or U8839 (N_8839,N_6647,N_7233);
nor U8840 (N_8840,N_7087,N_6394);
or U8841 (N_8841,N_5915,N_6136);
and U8842 (N_8842,N_7447,N_5430);
nor U8843 (N_8843,N_7070,N_6875);
nor U8844 (N_8844,N_6932,N_5736);
nor U8845 (N_8845,N_6180,N_6066);
nand U8846 (N_8846,N_6555,N_5574);
nand U8847 (N_8847,N_7158,N_6196);
nand U8848 (N_8848,N_7103,N_7469);
and U8849 (N_8849,N_6266,N_5307);
xor U8850 (N_8850,N_6146,N_5935);
nor U8851 (N_8851,N_6361,N_6260);
xnor U8852 (N_8852,N_7469,N_5406);
and U8853 (N_8853,N_5415,N_7272);
or U8854 (N_8854,N_5292,N_5559);
or U8855 (N_8855,N_6156,N_5353);
or U8856 (N_8856,N_7299,N_6781);
nand U8857 (N_8857,N_7374,N_6510);
nand U8858 (N_8858,N_5002,N_7282);
xor U8859 (N_8859,N_6698,N_5487);
xnor U8860 (N_8860,N_7304,N_5365);
xnor U8861 (N_8861,N_5499,N_7428);
nor U8862 (N_8862,N_6254,N_6878);
nand U8863 (N_8863,N_6010,N_5611);
and U8864 (N_8864,N_6891,N_5471);
nor U8865 (N_8865,N_7171,N_5164);
or U8866 (N_8866,N_6155,N_5625);
nand U8867 (N_8867,N_5419,N_5445);
nand U8868 (N_8868,N_7243,N_6627);
or U8869 (N_8869,N_6422,N_7392);
nand U8870 (N_8870,N_5259,N_5419);
nand U8871 (N_8871,N_6024,N_5824);
or U8872 (N_8872,N_6779,N_6657);
xor U8873 (N_8873,N_6734,N_5143);
nand U8874 (N_8874,N_7227,N_7238);
and U8875 (N_8875,N_5307,N_5491);
and U8876 (N_8876,N_7098,N_6014);
and U8877 (N_8877,N_5820,N_5280);
or U8878 (N_8878,N_6038,N_5032);
nor U8879 (N_8879,N_6428,N_5315);
or U8880 (N_8880,N_7086,N_5975);
or U8881 (N_8881,N_5990,N_7217);
nor U8882 (N_8882,N_5221,N_5907);
or U8883 (N_8883,N_6421,N_6133);
nand U8884 (N_8884,N_6653,N_5575);
nor U8885 (N_8885,N_7420,N_5056);
and U8886 (N_8886,N_6963,N_6462);
nor U8887 (N_8887,N_5075,N_7229);
xor U8888 (N_8888,N_6237,N_5302);
nand U8889 (N_8889,N_5531,N_6406);
nand U8890 (N_8890,N_7484,N_6675);
or U8891 (N_8891,N_7400,N_6715);
nor U8892 (N_8892,N_7274,N_5621);
nor U8893 (N_8893,N_6330,N_6337);
and U8894 (N_8894,N_6923,N_7345);
and U8895 (N_8895,N_5488,N_6253);
xor U8896 (N_8896,N_5433,N_7114);
nor U8897 (N_8897,N_5596,N_5098);
or U8898 (N_8898,N_6487,N_5612);
and U8899 (N_8899,N_5678,N_6775);
xnor U8900 (N_8900,N_5041,N_5724);
nor U8901 (N_8901,N_5118,N_5801);
nor U8902 (N_8902,N_7127,N_6009);
and U8903 (N_8903,N_5957,N_6241);
nor U8904 (N_8904,N_5902,N_6906);
nand U8905 (N_8905,N_5781,N_6721);
nand U8906 (N_8906,N_7347,N_6514);
and U8907 (N_8907,N_7042,N_5404);
xnor U8908 (N_8908,N_6103,N_7024);
nand U8909 (N_8909,N_5100,N_7296);
or U8910 (N_8910,N_7070,N_5276);
and U8911 (N_8911,N_5656,N_7196);
nor U8912 (N_8912,N_5024,N_5057);
and U8913 (N_8913,N_6231,N_7425);
nand U8914 (N_8914,N_6495,N_5712);
nand U8915 (N_8915,N_6276,N_5420);
nor U8916 (N_8916,N_7382,N_6851);
or U8917 (N_8917,N_7250,N_6286);
or U8918 (N_8918,N_6555,N_6854);
or U8919 (N_8919,N_6068,N_6822);
nor U8920 (N_8920,N_5065,N_7236);
or U8921 (N_8921,N_6318,N_7057);
nand U8922 (N_8922,N_6707,N_6528);
nor U8923 (N_8923,N_6383,N_7094);
nand U8924 (N_8924,N_5044,N_6544);
nand U8925 (N_8925,N_7221,N_6843);
xnor U8926 (N_8926,N_6775,N_6805);
and U8927 (N_8927,N_5525,N_5765);
or U8928 (N_8928,N_5304,N_5068);
xor U8929 (N_8929,N_6953,N_7047);
and U8930 (N_8930,N_7356,N_5469);
nand U8931 (N_8931,N_7210,N_5481);
nand U8932 (N_8932,N_7120,N_5074);
xnor U8933 (N_8933,N_7026,N_5126);
nand U8934 (N_8934,N_5442,N_7051);
nor U8935 (N_8935,N_7029,N_5066);
xnor U8936 (N_8936,N_5943,N_6335);
and U8937 (N_8937,N_6293,N_6653);
nand U8938 (N_8938,N_6377,N_6422);
and U8939 (N_8939,N_7018,N_5920);
and U8940 (N_8940,N_6389,N_6883);
nor U8941 (N_8941,N_6367,N_6060);
nand U8942 (N_8942,N_5098,N_5748);
xor U8943 (N_8943,N_6641,N_5792);
and U8944 (N_8944,N_6772,N_6192);
xnor U8945 (N_8945,N_6383,N_5098);
xor U8946 (N_8946,N_6107,N_6452);
nor U8947 (N_8947,N_6230,N_5181);
and U8948 (N_8948,N_6459,N_5746);
or U8949 (N_8949,N_6002,N_6250);
and U8950 (N_8950,N_7398,N_6762);
xnor U8951 (N_8951,N_5465,N_5537);
or U8952 (N_8952,N_6465,N_5700);
nor U8953 (N_8953,N_6634,N_5216);
and U8954 (N_8954,N_6107,N_5221);
nor U8955 (N_8955,N_5573,N_6228);
nand U8956 (N_8956,N_5675,N_7336);
and U8957 (N_8957,N_6836,N_5369);
nand U8958 (N_8958,N_7449,N_5637);
nand U8959 (N_8959,N_5345,N_6245);
nand U8960 (N_8960,N_5076,N_6882);
nor U8961 (N_8961,N_6161,N_7081);
or U8962 (N_8962,N_6730,N_5290);
and U8963 (N_8963,N_7469,N_6364);
nor U8964 (N_8964,N_6632,N_5341);
xnor U8965 (N_8965,N_6011,N_5755);
or U8966 (N_8966,N_6332,N_6860);
and U8967 (N_8967,N_5443,N_6223);
xnor U8968 (N_8968,N_6183,N_7216);
xor U8969 (N_8969,N_7298,N_6512);
xor U8970 (N_8970,N_5044,N_5406);
or U8971 (N_8971,N_6929,N_7331);
or U8972 (N_8972,N_6537,N_6883);
nand U8973 (N_8973,N_7231,N_5191);
or U8974 (N_8974,N_6029,N_6452);
and U8975 (N_8975,N_6282,N_6189);
nor U8976 (N_8976,N_5874,N_5555);
xor U8977 (N_8977,N_7230,N_7192);
nand U8978 (N_8978,N_6777,N_5497);
and U8979 (N_8979,N_7498,N_7424);
nor U8980 (N_8980,N_5806,N_5076);
and U8981 (N_8981,N_6458,N_6486);
and U8982 (N_8982,N_5186,N_6834);
or U8983 (N_8983,N_5537,N_5830);
and U8984 (N_8984,N_5764,N_6232);
or U8985 (N_8985,N_6742,N_6474);
nor U8986 (N_8986,N_6693,N_5727);
or U8987 (N_8987,N_7399,N_7332);
and U8988 (N_8988,N_6191,N_5559);
or U8989 (N_8989,N_7215,N_7087);
or U8990 (N_8990,N_7284,N_6346);
or U8991 (N_8991,N_5057,N_7119);
nand U8992 (N_8992,N_7064,N_5145);
nand U8993 (N_8993,N_5708,N_5498);
nand U8994 (N_8994,N_5047,N_6973);
and U8995 (N_8995,N_5228,N_6072);
and U8996 (N_8996,N_6653,N_6076);
or U8997 (N_8997,N_7334,N_6988);
xor U8998 (N_8998,N_5737,N_6840);
nand U8999 (N_8999,N_6847,N_5981);
nand U9000 (N_9000,N_5409,N_5669);
nand U9001 (N_9001,N_6688,N_5725);
xor U9002 (N_9002,N_6005,N_5350);
and U9003 (N_9003,N_6404,N_5054);
and U9004 (N_9004,N_5257,N_6117);
nand U9005 (N_9005,N_5479,N_6437);
and U9006 (N_9006,N_5714,N_6595);
xnor U9007 (N_9007,N_7279,N_6910);
nor U9008 (N_9008,N_5903,N_6514);
and U9009 (N_9009,N_6982,N_6659);
nor U9010 (N_9010,N_6671,N_6304);
xor U9011 (N_9011,N_6930,N_6802);
or U9012 (N_9012,N_5573,N_7052);
or U9013 (N_9013,N_7487,N_6688);
and U9014 (N_9014,N_6398,N_7128);
xnor U9015 (N_9015,N_6838,N_7183);
nor U9016 (N_9016,N_7167,N_5885);
nand U9017 (N_9017,N_6050,N_6513);
or U9018 (N_9018,N_5654,N_5466);
nor U9019 (N_9019,N_7386,N_5931);
xor U9020 (N_9020,N_6670,N_6520);
and U9021 (N_9021,N_7119,N_6459);
nor U9022 (N_9022,N_6862,N_6329);
or U9023 (N_9023,N_5536,N_6831);
nor U9024 (N_9024,N_6818,N_5855);
nor U9025 (N_9025,N_6017,N_6246);
nand U9026 (N_9026,N_6446,N_6331);
and U9027 (N_9027,N_5861,N_7139);
nand U9028 (N_9028,N_5336,N_6512);
and U9029 (N_9029,N_7122,N_5561);
xnor U9030 (N_9030,N_5540,N_5332);
and U9031 (N_9031,N_7314,N_5972);
nor U9032 (N_9032,N_7163,N_6746);
and U9033 (N_9033,N_7203,N_5037);
xnor U9034 (N_9034,N_5516,N_6410);
or U9035 (N_9035,N_5038,N_6283);
nand U9036 (N_9036,N_6571,N_6657);
nor U9037 (N_9037,N_5085,N_6522);
and U9038 (N_9038,N_7099,N_5144);
or U9039 (N_9039,N_5989,N_7434);
nand U9040 (N_9040,N_6121,N_6855);
and U9041 (N_9041,N_6051,N_5091);
nor U9042 (N_9042,N_5754,N_6154);
xor U9043 (N_9043,N_5301,N_5470);
xnor U9044 (N_9044,N_5593,N_7229);
nand U9045 (N_9045,N_7090,N_7431);
or U9046 (N_9046,N_7194,N_7481);
and U9047 (N_9047,N_5456,N_5410);
nand U9048 (N_9048,N_6707,N_7473);
nor U9049 (N_9049,N_7084,N_6343);
nor U9050 (N_9050,N_7084,N_5938);
or U9051 (N_9051,N_6015,N_6350);
nand U9052 (N_9052,N_6191,N_7135);
and U9053 (N_9053,N_6528,N_7011);
and U9054 (N_9054,N_5380,N_5962);
nand U9055 (N_9055,N_5933,N_7122);
xor U9056 (N_9056,N_5108,N_5817);
nand U9057 (N_9057,N_6043,N_5524);
or U9058 (N_9058,N_5039,N_7254);
xnor U9059 (N_9059,N_6096,N_6451);
or U9060 (N_9060,N_7076,N_7430);
xor U9061 (N_9061,N_6065,N_5171);
nand U9062 (N_9062,N_6709,N_6638);
nand U9063 (N_9063,N_5554,N_7400);
or U9064 (N_9064,N_6175,N_7403);
nor U9065 (N_9065,N_6912,N_5123);
or U9066 (N_9066,N_6086,N_5937);
and U9067 (N_9067,N_6431,N_6511);
nor U9068 (N_9068,N_6618,N_7120);
xor U9069 (N_9069,N_6156,N_5250);
nor U9070 (N_9070,N_6167,N_6850);
or U9071 (N_9071,N_6515,N_6811);
nor U9072 (N_9072,N_6824,N_5600);
and U9073 (N_9073,N_7090,N_7115);
nor U9074 (N_9074,N_5967,N_5908);
nand U9075 (N_9075,N_5540,N_6642);
and U9076 (N_9076,N_6285,N_5769);
or U9077 (N_9077,N_5804,N_5486);
or U9078 (N_9078,N_5385,N_6892);
nor U9079 (N_9079,N_7313,N_6718);
and U9080 (N_9080,N_5807,N_6923);
nor U9081 (N_9081,N_5788,N_6653);
nor U9082 (N_9082,N_6420,N_5886);
and U9083 (N_9083,N_6196,N_6493);
and U9084 (N_9084,N_6635,N_5143);
and U9085 (N_9085,N_6573,N_7289);
xor U9086 (N_9086,N_6875,N_7450);
nor U9087 (N_9087,N_7342,N_5738);
xor U9088 (N_9088,N_6682,N_6660);
or U9089 (N_9089,N_7098,N_5393);
and U9090 (N_9090,N_5527,N_7004);
nor U9091 (N_9091,N_6798,N_5565);
xnor U9092 (N_9092,N_6952,N_7107);
nand U9093 (N_9093,N_5829,N_5950);
and U9094 (N_9094,N_5145,N_7090);
and U9095 (N_9095,N_5202,N_5754);
or U9096 (N_9096,N_7223,N_7262);
nor U9097 (N_9097,N_5268,N_7162);
nor U9098 (N_9098,N_5713,N_5290);
nor U9099 (N_9099,N_6115,N_5536);
or U9100 (N_9100,N_6715,N_6635);
and U9101 (N_9101,N_5739,N_5887);
nor U9102 (N_9102,N_5839,N_7120);
nand U9103 (N_9103,N_5850,N_5562);
and U9104 (N_9104,N_6450,N_6299);
or U9105 (N_9105,N_7422,N_5366);
xor U9106 (N_9106,N_7198,N_7161);
and U9107 (N_9107,N_6990,N_7218);
and U9108 (N_9108,N_7274,N_5882);
nor U9109 (N_9109,N_7287,N_5487);
nand U9110 (N_9110,N_5321,N_6991);
nor U9111 (N_9111,N_5205,N_5399);
or U9112 (N_9112,N_6997,N_7469);
xor U9113 (N_9113,N_7091,N_6634);
xnor U9114 (N_9114,N_6149,N_6259);
nor U9115 (N_9115,N_6153,N_6789);
and U9116 (N_9116,N_5647,N_6484);
nand U9117 (N_9117,N_7419,N_5879);
and U9118 (N_9118,N_6237,N_6459);
nor U9119 (N_9119,N_6569,N_5098);
or U9120 (N_9120,N_6605,N_5436);
xnor U9121 (N_9121,N_6796,N_7492);
xor U9122 (N_9122,N_6066,N_6848);
and U9123 (N_9123,N_7084,N_5991);
nand U9124 (N_9124,N_7117,N_5974);
nor U9125 (N_9125,N_5328,N_5639);
xnor U9126 (N_9126,N_6806,N_5579);
nand U9127 (N_9127,N_5376,N_6806);
nor U9128 (N_9128,N_6468,N_5813);
nor U9129 (N_9129,N_6618,N_7383);
nor U9130 (N_9130,N_7153,N_5621);
or U9131 (N_9131,N_5286,N_7214);
or U9132 (N_9132,N_6422,N_6065);
xor U9133 (N_9133,N_6692,N_5660);
and U9134 (N_9134,N_7111,N_6483);
nor U9135 (N_9135,N_6690,N_5398);
nand U9136 (N_9136,N_6889,N_7007);
or U9137 (N_9137,N_6970,N_5919);
nand U9138 (N_9138,N_6179,N_6481);
xor U9139 (N_9139,N_7185,N_6535);
and U9140 (N_9140,N_5246,N_7496);
nor U9141 (N_9141,N_5263,N_7224);
nor U9142 (N_9142,N_5977,N_6700);
nor U9143 (N_9143,N_5466,N_5237);
and U9144 (N_9144,N_6360,N_6107);
nor U9145 (N_9145,N_5187,N_5853);
nor U9146 (N_9146,N_6243,N_5510);
and U9147 (N_9147,N_5286,N_6887);
and U9148 (N_9148,N_6444,N_5642);
and U9149 (N_9149,N_7273,N_6247);
and U9150 (N_9150,N_7095,N_5863);
xor U9151 (N_9151,N_6612,N_6308);
or U9152 (N_9152,N_6117,N_6760);
nor U9153 (N_9153,N_6390,N_5131);
and U9154 (N_9154,N_5945,N_5662);
nor U9155 (N_9155,N_5253,N_6797);
or U9156 (N_9156,N_5979,N_6149);
or U9157 (N_9157,N_6259,N_5008);
and U9158 (N_9158,N_6528,N_6656);
and U9159 (N_9159,N_5701,N_5650);
nor U9160 (N_9160,N_5462,N_6107);
nor U9161 (N_9161,N_5409,N_6163);
nand U9162 (N_9162,N_7262,N_5675);
and U9163 (N_9163,N_5966,N_5741);
nor U9164 (N_9164,N_5999,N_5419);
nor U9165 (N_9165,N_6284,N_5003);
nor U9166 (N_9166,N_6662,N_6358);
or U9167 (N_9167,N_7301,N_5259);
xnor U9168 (N_9168,N_6382,N_6990);
nor U9169 (N_9169,N_7373,N_6560);
and U9170 (N_9170,N_5910,N_5447);
nor U9171 (N_9171,N_5753,N_6416);
and U9172 (N_9172,N_7086,N_7015);
xor U9173 (N_9173,N_6570,N_6748);
xor U9174 (N_9174,N_7355,N_5716);
nor U9175 (N_9175,N_6802,N_5647);
and U9176 (N_9176,N_7392,N_7052);
nand U9177 (N_9177,N_5644,N_7051);
nor U9178 (N_9178,N_6659,N_5050);
nand U9179 (N_9179,N_5901,N_6648);
nand U9180 (N_9180,N_6079,N_6769);
xor U9181 (N_9181,N_6488,N_5715);
and U9182 (N_9182,N_5631,N_7131);
nand U9183 (N_9183,N_6644,N_6420);
nor U9184 (N_9184,N_6767,N_6555);
and U9185 (N_9185,N_7155,N_6636);
and U9186 (N_9186,N_7376,N_6161);
nor U9187 (N_9187,N_7427,N_7394);
or U9188 (N_9188,N_5739,N_6897);
nand U9189 (N_9189,N_5131,N_5373);
xnor U9190 (N_9190,N_5743,N_6794);
nand U9191 (N_9191,N_6148,N_5266);
nand U9192 (N_9192,N_7361,N_6744);
and U9193 (N_9193,N_5538,N_6095);
xnor U9194 (N_9194,N_5141,N_7334);
and U9195 (N_9195,N_6759,N_5025);
nand U9196 (N_9196,N_7277,N_6030);
nor U9197 (N_9197,N_6707,N_7366);
xor U9198 (N_9198,N_5636,N_6072);
and U9199 (N_9199,N_6037,N_7341);
and U9200 (N_9200,N_7214,N_5688);
or U9201 (N_9201,N_5321,N_7055);
nand U9202 (N_9202,N_6509,N_5475);
and U9203 (N_9203,N_6593,N_5629);
nor U9204 (N_9204,N_6209,N_6181);
nor U9205 (N_9205,N_6680,N_7292);
or U9206 (N_9206,N_7052,N_5821);
xor U9207 (N_9207,N_6879,N_7052);
and U9208 (N_9208,N_6605,N_5776);
nand U9209 (N_9209,N_5575,N_5718);
xor U9210 (N_9210,N_6193,N_5489);
nor U9211 (N_9211,N_7308,N_5666);
xnor U9212 (N_9212,N_6664,N_6606);
nand U9213 (N_9213,N_5163,N_6912);
nor U9214 (N_9214,N_5391,N_6703);
or U9215 (N_9215,N_5649,N_6780);
and U9216 (N_9216,N_5298,N_6566);
nand U9217 (N_9217,N_5853,N_6763);
xor U9218 (N_9218,N_5263,N_6242);
nand U9219 (N_9219,N_5036,N_5321);
xnor U9220 (N_9220,N_6448,N_6192);
nor U9221 (N_9221,N_6933,N_6461);
and U9222 (N_9222,N_6981,N_6070);
nand U9223 (N_9223,N_5256,N_6137);
nand U9224 (N_9224,N_7146,N_5226);
nor U9225 (N_9225,N_6292,N_5844);
xor U9226 (N_9226,N_6386,N_6587);
xnor U9227 (N_9227,N_6812,N_7391);
xor U9228 (N_9228,N_7084,N_5901);
nand U9229 (N_9229,N_5477,N_5230);
nand U9230 (N_9230,N_6024,N_5219);
nand U9231 (N_9231,N_5167,N_5055);
and U9232 (N_9232,N_6015,N_5309);
nor U9233 (N_9233,N_5713,N_6468);
xor U9234 (N_9234,N_7424,N_6221);
nand U9235 (N_9235,N_6842,N_6508);
or U9236 (N_9236,N_7239,N_5538);
and U9237 (N_9237,N_7411,N_5334);
nor U9238 (N_9238,N_7343,N_7077);
nor U9239 (N_9239,N_6759,N_5481);
nor U9240 (N_9240,N_6843,N_7430);
nand U9241 (N_9241,N_5757,N_7353);
nand U9242 (N_9242,N_6930,N_5640);
nand U9243 (N_9243,N_6739,N_7295);
and U9244 (N_9244,N_5815,N_5208);
nand U9245 (N_9245,N_6109,N_5623);
nand U9246 (N_9246,N_6024,N_7126);
nor U9247 (N_9247,N_6273,N_6115);
and U9248 (N_9248,N_5120,N_5020);
or U9249 (N_9249,N_5582,N_6536);
xor U9250 (N_9250,N_5116,N_5747);
or U9251 (N_9251,N_6572,N_5762);
xor U9252 (N_9252,N_7343,N_6403);
xnor U9253 (N_9253,N_5466,N_5844);
nand U9254 (N_9254,N_6979,N_6388);
nand U9255 (N_9255,N_5328,N_7166);
or U9256 (N_9256,N_5782,N_6647);
nand U9257 (N_9257,N_5545,N_5731);
or U9258 (N_9258,N_5236,N_7309);
xor U9259 (N_9259,N_6548,N_5632);
nand U9260 (N_9260,N_6575,N_6480);
nand U9261 (N_9261,N_5673,N_5998);
and U9262 (N_9262,N_5883,N_7355);
xor U9263 (N_9263,N_5190,N_5783);
nor U9264 (N_9264,N_5614,N_6607);
nor U9265 (N_9265,N_7173,N_5741);
nand U9266 (N_9266,N_6136,N_5301);
nor U9267 (N_9267,N_6149,N_7336);
and U9268 (N_9268,N_5461,N_6085);
or U9269 (N_9269,N_6219,N_6833);
xor U9270 (N_9270,N_6969,N_7427);
nor U9271 (N_9271,N_5664,N_7041);
nand U9272 (N_9272,N_5076,N_6113);
and U9273 (N_9273,N_5889,N_5351);
nand U9274 (N_9274,N_7206,N_6508);
nand U9275 (N_9275,N_5985,N_5575);
xnor U9276 (N_9276,N_6688,N_5497);
nand U9277 (N_9277,N_7070,N_7214);
nor U9278 (N_9278,N_5889,N_6688);
nor U9279 (N_9279,N_5112,N_6584);
or U9280 (N_9280,N_6468,N_5802);
nand U9281 (N_9281,N_5655,N_6875);
and U9282 (N_9282,N_6007,N_7388);
or U9283 (N_9283,N_5437,N_6294);
nor U9284 (N_9284,N_6119,N_6955);
and U9285 (N_9285,N_6108,N_5679);
and U9286 (N_9286,N_5958,N_6408);
nand U9287 (N_9287,N_6618,N_6465);
nor U9288 (N_9288,N_6365,N_5679);
and U9289 (N_9289,N_6197,N_7194);
xnor U9290 (N_9290,N_6686,N_6143);
nand U9291 (N_9291,N_6720,N_7477);
nand U9292 (N_9292,N_7490,N_5330);
or U9293 (N_9293,N_5274,N_7238);
nor U9294 (N_9294,N_5626,N_5904);
and U9295 (N_9295,N_6550,N_6062);
and U9296 (N_9296,N_7154,N_5172);
nand U9297 (N_9297,N_6398,N_5764);
or U9298 (N_9298,N_7190,N_7182);
nand U9299 (N_9299,N_5841,N_6717);
or U9300 (N_9300,N_7220,N_5476);
xor U9301 (N_9301,N_6417,N_5236);
nand U9302 (N_9302,N_7000,N_5642);
xnor U9303 (N_9303,N_5482,N_6671);
or U9304 (N_9304,N_6302,N_5893);
nand U9305 (N_9305,N_6854,N_7480);
or U9306 (N_9306,N_6698,N_5794);
nand U9307 (N_9307,N_6683,N_5884);
xnor U9308 (N_9308,N_7345,N_5215);
or U9309 (N_9309,N_5278,N_7443);
and U9310 (N_9310,N_6378,N_5569);
and U9311 (N_9311,N_6759,N_7156);
nand U9312 (N_9312,N_7051,N_6680);
or U9313 (N_9313,N_6737,N_7265);
and U9314 (N_9314,N_5049,N_5302);
nand U9315 (N_9315,N_6565,N_5311);
and U9316 (N_9316,N_6813,N_5860);
nor U9317 (N_9317,N_5300,N_5514);
xnor U9318 (N_9318,N_6487,N_5553);
xor U9319 (N_9319,N_5813,N_6978);
xnor U9320 (N_9320,N_5422,N_5490);
and U9321 (N_9321,N_6433,N_6431);
or U9322 (N_9322,N_6966,N_7409);
nand U9323 (N_9323,N_5909,N_7036);
xnor U9324 (N_9324,N_6106,N_6886);
nand U9325 (N_9325,N_6811,N_5982);
nand U9326 (N_9326,N_6073,N_7325);
xor U9327 (N_9327,N_7002,N_5515);
or U9328 (N_9328,N_6184,N_5604);
nor U9329 (N_9329,N_5130,N_6463);
nand U9330 (N_9330,N_7143,N_6998);
xnor U9331 (N_9331,N_6976,N_7320);
nand U9332 (N_9332,N_6978,N_5556);
nand U9333 (N_9333,N_6298,N_5775);
xnor U9334 (N_9334,N_5853,N_6867);
nand U9335 (N_9335,N_5586,N_5214);
nand U9336 (N_9336,N_5142,N_5000);
and U9337 (N_9337,N_7066,N_6318);
or U9338 (N_9338,N_7032,N_5600);
nor U9339 (N_9339,N_6696,N_5546);
nand U9340 (N_9340,N_6669,N_7297);
and U9341 (N_9341,N_5804,N_6550);
nand U9342 (N_9342,N_6652,N_6897);
and U9343 (N_9343,N_7287,N_7363);
nor U9344 (N_9344,N_6599,N_6983);
and U9345 (N_9345,N_6227,N_6150);
xnor U9346 (N_9346,N_6086,N_5765);
xnor U9347 (N_9347,N_6238,N_6404);
and U9348 (N_9348,N_6313,N_5852);
xnor U9349 (N_9349,N_6519,N_7246);
nor U9350 (N_9350,N_5194,N_6452);
nand U9351 (N_9351,N_5078,N_5783);
or U9352 (N_9352,N_7376,N_5369);
nor U9353 (N_9353,N_5129,N_6104);
nor U9354 (N_9354,N_5982,N_5587);
xnor U9355 (N_9355,N_5104,N_6243);
and U9356 (N_9356,N_7262,N_6644);
or U9357 (N_9357,N_5046,N_5570);
xnor U9358 (N_9358,N_5279,N_5109);
nand U9359 (N_9359,N_6486,N_6277);
xor U9360 (N_9360,N_5742,N_5398);
nor U9361 (N_9361,N_5205,N_5740);
nand U9362 (N_9362,N_6542,N_7319);
nand U9363 (N_9363,N_7136,N_6381);
xor U9364 (N_9364,N_7099,N_5764);
and U9365 (N_9365,N_6665,N_5456);
and U9366 (N_9366,N_6206,N_6637);
xnor U9367 (N_9367,N_7350,N_7409);
xor U9368 (N_9368,N_6589,N_6583);
nand U9369 (N_9369,N_5395,N_5869);
and U9370 (N_9370,N_7350,N_5404);
or U9371 (N_9371,N_7453,N_6436);
nand U9372 (N_9372,N_6066,N_5102);
xnor U9373 (N_9373,N_5302,N_6022);
or U9374 (N_9374,N_5234,N_5235);
nor U9375 (N_9375,N_6412,N_6714);
and U9376 (N_9376,N_7265,N_6782);
xnor U9377 (N_9377,N_5050,N_5209);
xor U9378 (N_9378,N_7357,N_5839);
or U9379 (N_9379,N_6342,N_5672);
xor U9380 (N_9380,N_7114,N_7158);
nor U9381 (N_9381,N_6689,N_7374);
and U9382 (N_9382,N_5914,N_5819);
or U9383 (N_9383,N_5813,N_5145);
and U9384 (N_9384,N_5174,N_7036);
and U9385 (N_9385,N_6420,N_5171);
or U9386 (N_9386,N_5296,N_6755);
nand U9387 (N_9387,N_7453,N_6569);
and U9388 (N_9388,N_6752,N_7471);
and U9389 (N_9389,N_5314,N_5199);
xnor U9390 (N_9390,N_6449,N_5400);
xnor U9391 (N_9391,N_5536,N_6333);
nand U9392 (N_9392,N_5032,N_7110);
or U9393 (N_9393,N_6628,N_5787);
xnor U9394 (N_9394,N_7002,N_6772);
xor U9395 (N_9395,N_7458,N_6765);
xor U9396 (N_9396,N_5457,N_6387);
nand U9397 (N_9397,N_5850,N_6602);
xor U9398 (N_9398,N_6727,N_5097);
xnor U9399 (N_9399,N_7327,N_6450);
or U9400 (N_9400,N_7109,N_5076);
and U9401 (N_9401,N_6510,N_7011);
xnor U9402 (N_9402,N_7083,N_5492);
xnor U9403 (N_9403,N_6065,N_7164);
and U9404 (N_9404,N_5047,N_7344);
nor U9405 (N_9405,N_5760,N_6507);
and U9406 (N_9406,N_5617,N_5098);
nand U9407 (N_9407,N_5663,N_5492);
nand U9408 (N_9408,N_5912,N_6912);
nor U9409 (N_9409,N_6821,N_7232);
or U9410 (N_9410,N_5790,N_5840);
nor U9411 (N_9411,N_7061,N_5224);
and U9412 (N_9412,N_5311,N_5718);
or U9413 (N_9413,N_5896,N_5223);
and U9414 (N_9414,N_5603,N_5009);
nand U9415 (N_9415,N_5315,N_6774);
nor U9416 (N_9416,N_6502,N_5530);
nand U9417 (N_9417,N_5452,N_5280);
xor U9418 (N_9418,N_7377,N_5865);
and U9419 (N_9419,N_7442,N_7299);
or U9420 (N_9420,N_5922,N_6751);
nand U9421 (N_9421,N_5027,N_6852);
nor U9422 (N_9422,N_5578,N_5012);
nand U9423 (N_9423,N_6430,N_5309);
xor U9424 (N_9424,N_6703,N_6393);
xnor U9425 (N_9425,N_5218,N_6891);
xnor U9426 (N_9426,N_5141,N_6369);
nor U9427 (N_9427,N_5657,N_5973);
or U9428 (N_9428,N_6573,N_7308);
nand U9429 (N_9429,N_5117,N_6110);
or U9430 (N_9430,N_7043,N_5708);
or U9431 (N_9431,N_5536,N_5839);
nand U9432 (N_9432,N_6522,N_5853);
xnor U9433 (N_9433,N_6995,N_5626);
nand U9434 (N_9434,N_7489,N_6044);
nor U9435 (N_9435,N_6873,N_5733);
and U9436 (N_9436,N_6535,N_6091);
nand U9437 (N_9437,N_6956,N_5134);
and U9438 (N_9438,N_7276,N_7148);
xnor U9439 (N_9439,N_6092,N_7401);
nand U9440 (N_9440,N_7369,N_5772);
or U9441 (N_9441,N_6110,N_6681);
or U9442 (N_9442,N_5567,N_5160);
and U9443 (N_9443,N_7352,N_6905);
nor U9444 (N_9444,N_5745,N_6680);
nor U9445 (N_9445,N_7367,N_5415);
xor U9446 (N_9446,N_6576,N_6932);
xnor U9447 (N_9447,N_5464,N_6156);
or U9448 (N_9448,N_6178,N_5498);
nand U9449 (N_9449,N_5143,N_5287);
and U9450 (N_9450,N_6025,N_6095);
or U9451 (N_9451,N_6193,N_5538);
xor U9452 (N_9452,N_5551,N_6441);
nor U9453 (N_9453,N_5149,N_6443);
nor U9454 (N_9454,N_5708,N_7222);
xnor U9455 (N_9455,N_5213,N_6620);
xnor U9456 (N_9456,N_5595,N_5410);
xor U9457 (N_9457,N_6274,N_6653);
and U9458 (N_9458,N_6764,N_7116);
nand U9459 (N_9459,N_6597,N_6842);
or U9460 (N_9460,N_7044,N_6710);
or U9461 (N_9461,N_6810,N_5158);
and U9462 (N_9462,N_6767,N_5476);
or U9463 (N_9463,N_6196,N_6917);
or U9464 (N_9464,N_5073,N_6609);
or U9465 (N_9465,N_6251,N_5173);
or U9466 (N_9466,N_5589,N_6831);
nand U9467 (N_9467,N_5965,N_5320);
or U9468 (N_9468,N_6214,N_6153);
nand U9469 (N_9469,N_5091,N_7496);
or U9470 (N_9470,N_6143,N_6420);
or U9471 (N_9471,N_7174,N_7474);
and U9472 (N_9472,N_5461,N_5555);
and U9473 (N_9473,N_5177,N_5594);
or U9474 (N_9474,N_5835,N_6270);
nand U9475 (N_9475,N_5693,N_6174);
or U9476 (N_9476,N_6039,N_5326);
or U9477 (N_9477,N_6234,N_5334);
nand U9478 (N_9478,N_7337,N_6040);
xnor U9479 (N_9479,N_6922,N_7347);
nor U9480 (N_9480,N_7176,N_5740);
xnor U9481 (N_9481,N_6393,N_6474);
nor U9482 (N_9482,N_5790,N_5426);
or U9483 (N_9483,N_7002,N_5658);
nand U9484 (N_9484,N_6101,N_7132);
nor U9485 (N_9485,N_5540,N_6274);
xor U9486 (N_9486,N_5499,N_6991);
nand U9487 (N_9487,N_5287,N_6095);
and U9488 (N_9488,N_6436,N_6653);
nor U9489 (N_9489,N_5308,N_5507);
nand U9490 (N_9490,N_5125,N_5790);
xnor U9491 (N_9491,N_5944,N_6384);
nor U9492 (N_9492,N_6377,N_7204);
nand U9493 (N_9493,N_5410,N_5638);
xnor U9494 (N_9494,N_5648,N_6276);
or U9495 (N_9495,N_7425,N_5013);
xor U9496 (N_9496,N_5538,N_5530);
and U9497 (N_9497,N_5189,N_6812);
or U9498 (N_9498,N_5715,N_5930);
xnor U9499 (N_9499,N_7382,N_6513);
nand U9500 (N_9500,N_5453,N_6244);
or U9501 (N_9501,N_5805,N_7124);
nor U9502 (N_9502,N_5542,N_5135);
nand U9503 (N_9503,N_7000,N_7202);
nand U9504 (N_9504,N_5156,N_5480);
nor U9505 (N_9505,N_5292,N_6296);
or U9506 (N_9506,N_7075,N_6543);
or U9507 (N_9507,N_5243,N_6388);
and U9508 (N_9508,N_6446,N_5626);
or U9509 (N_9509,N_6153,N_6977);
and U9510 (N_9510,N_7290,N_6492);
nand U9511 (N_9511,N_6250,N_5937);
and U9512 (N_9512,N_5997,N_5975);
nand U9513 (N_9513,N_6566,N_5123);
xor U9514 (N_9514,N_6945,N_5966);
and U9515 (N_9515,N_7485,N_7386);
nand U9516 (N_9516,N_6424,N_6681);
or U9517 (N_9517,N_5486,N_6450);
xnor U9518 (N_9518,N_7039,N_6282);
nand U9519 (N_9519,N_6049,N_6506);
or U9520 (N_9520,N_6782,N_6775);
nor U9521 (N_9521,N_5201,N_6751);
or U9522 (N_9522,N_5988,N_6232);
nor U9523 (N_9523,N_6632,N_5775);
or U9524 (N_9524,N_5476,N_5450);
xor U9525 (N_9525,N_7266,N_7110);
nor U9526 (N_9526,N_7449,N_7048);
and U9527 (N_9527,N_6907,N_6631);
xor U9528 (N_9528,N_5350,N_6787);
nand U9529 (N_9529,N_5823,N_6420);
nor U9530 (N_9530,N_5796,N_6886);
or U9531 (N_9531,N_6619,N_7075);
nor U9532 (N_9532,N_5123,N_6307);
or U9533 (N_9533,N_5673,N_6145);
or U9534 (N_9534,N_7241,N_6399);
xnor U9535 (N_9535,N_5797,N_6875);
nor U9536 (N_9536,N_5220,N_5152);
nand U9537 (N_9537,N_6534,N_6537);
xnor U9538 (N_9538,N_5885,N_5056);
or U9539 (N_9539,N_5559,N_5728);
xor U9540 (N_9540,N_6759,N_6650);
or U9541 (N_9541,N_6464,N_6662);
xnor U9542 (N_9542,N_6221,N_6756);
xnor U9543 (N_9543,N_5450,N_5238);
xnor U9544 (N_9544,N_5397,N_5887);
nand U9545 (N_9545,N_6996,N_5992);
and U9546 (N_9546,N_6828,N_6140);
nand U9547 (N_9547,N_5521,N_6607);
and U9548 (N_9548,N_6023,N_5949);
or U9549 (N_9549,N_6480,N_6119);
and U9550 (N_9550,N_5721,N_6075);
or U9551 (N_9551,N_5180,N_6648);
and U9552 (N_9552,N_6532,N_6259);
and U9553 (N_9553,N_6796,N_5534);
nand U9554 (N_9554,N_5020,N_6901);
nor U9555 (N_9555,N_6218,N_5537);
or U9556 (N_9556,N_5038,N_6545);
nand U9557 (N_9557,N_6009,N_6846);
xor U9558 (N_9558,N_5748,N_6942);
nor U9559 (N_9559,N_7375,N_5285);
and U9560 (N_9560,N_7211,N_7190);
xnor U9561 (N_9561,N_7148,N_6290);
xor U9562 (N_9562,N_5225,N_5768);
nor U9563 (N_9563,N_6136,N_6679);
xnor U9564 (N_9564,N_6843,N_7088);
or U9565 (N_9565,N_7405,N_5244);
or U9566 (N_9566,N_5701,N_6091);
nand U9567 (N_9567,N_5342,N_6515);
xnor U9568 (N_9568,N_6740,N_5501);
nand U9569 (N_9569,N_5799,N_7320);
xnor U9570 (N_9570,N_6453,N_5562);
and U9571 (N_9571,N_5943,N_6818);
xnor U9572 (N_9572,N_7161,N_7435);
nor U9573 (N_9573,N_6167,N_6694);
and U9574 (N_9574,N_6384,N_6024);
nand U9575 (N_9575,N_6919,N_6556);
nor U9576 (N_9576,N_5559,N_6856);
and U9577 (N_9577,N_5422,N_6925);
xnor U9578 (N_9578,N_5306,N_7230);
or U9579 (N_9579,N_6429,N_7393);
xnor U9580 (N_9580,N_5962,N_6415);
nor U9581 (N_9581,N_6583,N_6905);
nor U9582 (N_9582,N_7291,N_7304);
or U9583 (N_9583,N_6529,N_6007);
xnor U9584 (N_9584,N_6194,N_6577);
xor U9585 (N_9585,N_5720,N_6931);
nand U9586 (N_9586,N_5705,N_5664);
xor U9587 (N_9587,N_6853,N_7470);
xor U9588 (N_9588,N_6313,N_5637);
and U9589 (N_9589,N_5800,N_6199);
xnor U9590 (N_9590,N_5619,N_6741);
xor U9591 (N_9591,N_6226,N_5574);
nor U9592 (N_9592,N_5324,N_5136);
nand U9593 (N_9593,N_6658,N_6207);
or U9594 (N_9594,N_7101,N_7382);
nor U9595 (N_9595,N_6395,N_6418);
nor U9596 (N_9596,N_6145,N_6598);
or U9597 (N_9597,N_5893,N_5175);
or U9598 (N_9598,N_6972,N_7137);
and U9599 (N_9599,N_5841,N_6207);
or U9600 (N_9600,N_6756,N_6886);
nor U9601 (N_9601,N_6622,N_6798);
xor U9602 (N_9602,N_7014,N_6955);
nor U9603 (N_9603,N_5874,N_5408);
xnor U9604 (N_9604,N_7065,N_5343);
nand U9605 (N_9605,N_6212,N_7042);
nand U9606 (N_9606,N_5939,N_6571);
nor U9607 (N_9607,N_7185,N_5984);
nor U9608 (N_9608,N_6610,N_5054);
nand U9609 (N_9609,N_6927,N_5306);
nand U9610 (N_9610,N_5682,N_5570);
nand U9611 (N_9611,N_7097,N_6123);
and U9612 (N_9612,N_6537,N_6726);
and U9613 (N_9613,N_7312,N_6466);
or U9614 (N_9614,N_6018,N_6691);
nand U9615 (N_9615,N_7163,N_6945);
nand U9616 (N_9616,N_6281,N_5780);
or U9617 (N_9617,N_5524,N_7088);
nand U9618 (N_9618,N_5241,N_5567);
nand U9619 (N_9619,N_7170,N_5718);
nor U9620 (N_9620,N_6774,N_5307);
xor U9621 (N_9621,N_5447,N_5523);
nand U9622 (N_9622,N_5848,N_6887);
xnor U9623 (N_9623,N_6935,N_5767);
nand U9624 (N_9624,N_7098,N_6882);
nand U9625 (N_9625,N_6550,N_6564);
or U9626 (N_9626,N_6870,N_6608);
nand U9627 (N_9627,N_6089,N_7253);
nand U9628 (N_9628,N_6935,N_6243);
xor U9629 (N_9629,N_7066,N_6970);
nor U9630 (N_9630,N_7067,N_5871);
nand U9631 (N_9631,N_5314,N_7051);
and U9632 (N_9632,N_6515,N_5579);
nor U9633 (N_9633,N_7371,N_7083);
xor U9634 (N_9634,N_6645,N_5028);
nor U9635 (N_9635,N_5519,N_5390);
or U9636 (N_9636,N_6346,N_6693);
or U9637 (N_9637,N_7103,N_6865);
or U9638 (N_9638,N_6381,N_6749);
xor U9639 (N_9639,N_6402,N_6507);
nand U9640 (N_9640,N_7147,N_7264);
or U9641 (N_9641,N_5466,N_5707);
xor U9642 (N_9642,N_5235,N_7007);
xor U9643 (N_9643,N_5804,N_6924);
xor U9644 (N_9644,N_7415,N_6163);
and U9645 (N_9645,N_6285,N_7128);
nand U9646 (N_9646,N_6350,N_6709);
nand U9647 (N_9647,N_5455,N_5130);
xor U9648 (N_9648,N_6873,N_6753);
xnor U9649 (N_9649,N_5857,N_6335);
xor U9650 (N_9650,N_5872,N_6822);
and U9651 (N_9651,N_5421,N_5060);
and U9652 (N_9652,N_5788,N_5921);
or U9653 (N_9653,N_6339,N_7015);
and U9654 (N_9654,N_5245,N_5661);
and U9655 (N_9655,N_5706,N_6430);
and U9656 (N_9656,N_5667,N_5635);
or U9657 (N_9657,N_5797,N_6239);
nand U9658 (N_9658,N_6471,N_5167);
or U9659 (N_9659,N_7360,N_5075);
and U9660 (N_9660,N_5871,N_5738);
nand U9661 (N_9661,N_7440,N_6362);
or U9662 (N_9662,N_6901,N_5189);
xor U9663 (N_9663,N_6795,N_6808);
and U9664 (N_9664,N_5976,N_5825);
nand U9665 (N_9665,N_7370,N_7170);
or U9666 (N_9666,N_5378,N_6864);
or U9667 (N_9667,N_5142,N_6650);
or U9668 (N_9668,N_7394,N_5788);
or U9669 (N_9669,N_6400,N_6001);
nand U9670 (N_9670,N_6426,N_5839);
nand U9671 (N_9671,N_5280,N_5970);
xor U9672 (N_9672,N_6889,N_6956);
and U9673 (N_9673,N_6762,N_6414);
nor U9674 (N_9674,N_6692,N_7009);
and U9675 (N_9675,N_5597,N_7083);
and U9676 (N_9676,N_6405,N_6757);
or U9677 (N_9677,N_6130,N_6508);
or U9678 (N_9678,N_5968,N_6135);
and U9679 (N_9679,N_7338,N_6633);
nor U9680 (N_9680,N_6457,N_5609);
xor U9681 (N_9681,N_5234,N_5972);
nor U9682 (N_9682,N_5460,N_6528);
nor U9683 (N_9683,N_7496,N_7102);
nor U9684 (N_9684,N_5620,N_5357);
nand U9685 (N_9685,N_5689,N_7488);
nand U9686 (N_9686,N_7152,N_5054);
nand U9687 (N_9687,N_7438,N_7080);
and U9688 (N_9688,N_6727,N_5347);
or U9689 (N_9689,N_5890,N_6744);
nand U9690 (N_9690,N_7107,N_5134);
or U9691 (N_9691,N_5199,N_6082);
or U9692 (N_9692,N_7170,N_6253);
and U9693 (N_9693,N_5061,N_5701);
xor U9694 (N_9694,N_6978,N_6937);
xor U9695 (N_9695,N_7120,N_6474);
nand U9696 (N_9696,N_5599,N_5174);
nand U9697 (N_9697,N_6568,N_6732);
nand U9698 (N_9698,N_6886,N_5413);
and U9699 (N_9699,N_7133,N_5172);
nor U9700 (N_9700,N_7030,N_6366);
xor U9701 (N_9701,N_7377,N_5817);
nand U9702 (N_9702,N_6001,N_6867);
or U9703 (N_9703,N_6572,N_6185);
or U9704 (N_9704,N_5163,N_7374);
nor U9705 (N_9705,N_7279,N_7321);
nor U9706 (N_9706,N_7061,N_5239);
and U9707 (N_9707,N_6271,N_6167);
xnor U9708 (N_9708,N_6006,N_5070);
xor U9709 (N_9709,N_6347,N_7195);
nor U9710 (N_9710,N_5288,N_5671);
nor U9711 (N_9711,N_6408,N_5982);
nand U9712 (N_9712,N_6015,N_7400);
xor U9713 (N_9713,N_6269,N_5058);
nand U9714 (N_9714,N_6106,N_7375);
nand U9715 (N_9715,N_6586,N_6653);
or U9716 (N_9716,N_6781,N_6362);
nand U9717 (N_9717,N_7079,N_6498);
nor U9718 (N_9718,N_6210,N_7292);
and U9719 (N_9719,N_5040,N_6747);
nand U9720 (N_9720,N_5324,N_5860);
and U9721 (N_9721,N_6802,N_6782);
xnor U9722 (N_9722,N_5961,N_5803);
and U9723 (N_9723,N_5796,N_6885);
or U9724 (N_9724,N_6700,N_6934);
xor U9725 (N_9725,N_5270,N_7076);
or U9726 (N_9726,N_7014,N_7292);
xor U9727 (N_9727,N_6847,N_6135);
xnor U9728 (N_9728,N_6766,N_7488);
or U9729 (N_9729,N_7337,N_6129);
nand U9730 (N_9730,N_7475,N_5126);
and U9731 (N_9731,N_6193,N_6792);
xnor U9732 (N_9732,N_6622,N_6026);
nor U9733 (N_9733,N_6871,N_6255);
nand U9734 (N_9734,N_6205,N_6325);
nor U9735 (N_9735,N_5286,N_7094);
nand U9736 (N_9736,N_5094,N_6199);
or U9737 (N_9737,N_7264,N_6022);
nand U9738 (N_9738,N_5402,N_5909);
and U9739 (N_9739,N_5389,N_6222);
nor U9740 (N_9740,N_6702,N_6779);
and U9741 (N_9741,N_5646,N_5156);
nand U9742 (N_9742,N_5714,N_6301);
or U9743 (N_9743,N_5050,N_5354);
xnor U9744 (N_9744,N_5978,N_6216);
and U9745 (N_9745,N_6994,N_5883);
nor U9746 (N_9746,N_7339,N_5285);
nand U9747 (N_9747,N_5173,N_5382);
nor U9748 (N_9748,N_5674,N_5212);
nand U9749 (N_9749,N_7249,N_5646);
xor U9750 (N_9750,N_5443,N_6164);
xnor U9751 (N_9751,N_7319,N_5660);
nand U9752 (N_9752,N_5417,N_5138);
nor U9753 (N_9753,N_6778,N_6898);
and U9754 (N_9754,N_6344,N_7438);
nor U9755 (N_9755,N_6758,N_5413);
nand U9756 (N_9756,N_6994,N_6361);
nor U9757 (N_9757,N_5752,N_5841);
or U9758 (N_9758,N_5864,N_6125);
or U9759 (N_9759,N_5428,N_7261);
or U9760 (N_9760,N_7358,N_5623);
and U9761 (N_9761,N_5429,N_6409);
or U9762 (N_9762,N_6019,N_6566);
xor U9763 (N_9763,N_6358,N_6223);
and U9764 (N_9764,N_5917,N_7328);
or U9765 (N_9765,N_5418,N_6726);
xor U9766 (N_9766,N_5483,N_5418);
or U9767 (N_9767,N_6002,N_5013);
nor U9768 (N_9768,N_5034,N_7405);
nor U9769 (N_9769,N_5383,N_6770);
nor U9770 (N_9770,N_6463,N_5133);
or U9771 (N_9771,N_6596,N_6091);
and U9772 (N_9772,N_6045,N_6913);
nor U9773 (N_9773,N_5581,N_5272);
nand U9774 (N_9774,N_6234,N_6618);
and U9775 (N_9775,N_7213,N_6361);
and U9776 (N_9776,N_6860,N_6196);
and U9777 (N_9777,N_6532,N_7375);
nor U9778 (N_9778,N_6321,N_5815);
or U9779 (N_9779,N_5921,N_6402);
or U9780 (N_9780,N_5211,N_7461);
or U9781 (N_9781,N_6539,N_7476);
xor U9782 (N_9782,N_5814,N_7252);
or U9783 (N_9783,N_5393,N_5972);
or U9784 (N_9784,N_6473,N_6284);
nor U9785 (N_9785,N_6715,N_6561);
nor U9786 (N_9786,N_7212,N_5549);
nor U9787 (N_9787,N_5030,N_7298);
and U9788 (N_9788,N_5392,N_5946);
and U9789 (N_9789,N_5924,N_5002);
and U9790 (N_9790,N_6903,N_6115);
and U9791 (N_9791,N_6868,N_6815);
and U9792 (N_9792,N_6496,N_6755);
xor U9793 (N_9793,N_5653,N_7177);
nand U9794 (N_9794,N_6058,N_5155);
and U9795 (N_9795,N_6830,N_6092);
nand U9796 (N_9796,N_6836,N_6899);
or U9797 (N_9797,N_5468,N_5657);
and U9798 (N_9798,N_6492,N_6661);
or U9799 (N_9799,N_5470,N_6934);
xor U9800 (N_9800,N_6342,N_6797);
or U9801 (N_9801,N_6526,N_5405);
and U9802 (N_9802,N_6706,N_5052);
xor U9803 (N_9803,N_5560,N_7192);
or U9804 (N_9804,N_5652,N_5351);
xnor U9805 (N_9805,N_5589,N_5681);
xnor U9806 (N_9806,N_5947,N_6097);
nor U9807 (N_9807,N_7492,N_6859);
and U9808 (N_9808,N_5780,N_5335);
or U9809 (N_9809,N_6452,N_6697);
xor U9810 (N_9810,N_6794,N_7471);
or U9811 (N_9811,N_5480,N_6641);
xnor U9812 (N_9812,N_5064,N_7425);
nor U9813 (N_9813,N_5880,N_5264);
nor U9814 (N_9814,N_6670,N_5114);
nor U9815 (N_9815,N_5802,N_6699);
or U9816 (N_9816,N_6374,N_5602);
or U9817 (N_9817,N_5114,N_7103);
and U9818 (N_9818,N_5512,N_5535);
or U9819 (N_9819,N_5077,N_5906);
or U9820 (N_9820,N_7190,N_5592);
or U9821 (N_9821,N_6381,N_6185);
nor U9822 (N_9822,N_5758,N_6753);
xnor U9823 (N_9823,N_6351,N_6604);
xor U9824 (N_9824,N_7430,N_5257);
nor U9825 (N_9825,N_5133,N_6186);
and U9826 (N_9826,N_6997,N_6918);
or U9827 (N_9827,N_5657,N_6611);
and U9828 (N_9828,N_6947,N_5347);
nor U9829 (N_9829,N_5007,N_5470);
and U9830 (N_9830,N_6867,N_6317);
nand U9831 (N_9831,N_5848,N_7324);
or U9832 (N_9832,N_6233,N_5897);
and U9833 (N_9833,N_6158,N_6163);
nand U9834 (N_9834,N_6298,N_5496);
nand U9835 (N_9835,N_6203,N_7167);
nand U9836 (N_9836,N_5015,N_6349);
or U9837 (N_9837,N_7355,N_6483);
nor U9838 (N_9838,N_6168,N_6129);
nor U9839 (N_9839,N_5755,N_7266);
xor U9840 (N_9840,N_5110,N_5065);
and U9841 (N_9841,N_5020,N_5418);
and U9842 (N_9842,N_6832,N_5114);
or U9843 (N_9843,N_7175,N_5983);
nor U9844 (N_9844,N_7240,N_6496);
and U9845 (N_9845,N_6068,N_7248);
and U9846 (N_9846,N_6191,N_6949);
nand U9847 (N_9847,N_5845,N_5248);
nor U9848 (N_9848,N_6714,N_6292);
and U9849 (N_9849,N_7498,N_5021);
xor U9850 (N_9850,N_5388,N_5104);
and U9851 (N_9851,N_6658,N_5666);
nand U9852 (N_9852,N_6466,N_5443);
or U9853 (N_9853,N_5761,N_5407);
nand U9854 (N_9854,N_6053,N_5915);
or U9855 (N_9855,N_5249,N_5636);
and U9856 (N_9856,N_6863,N_7046);
or U9857 (N_9857,N_6689,N_7446);
or U9858 (N_9858,N_6805,N_6281);
xnor U9859 (N_9859,N_7180,N_5381);
nand U9860 (N_9860,N_7279,N_5640);
nand U9861 (N_9861,N_5407,N_6324);
or U9862 (N_9862,N_7318,N_5143);
nand U9863 (N_9863,N_7056,N_5999);
nand U9864 (N_9864,N_6475,N_5963);
or U9865 (N_9865,N_5085,N_5482);
xor U9866 (N_9866,N_5717,N_7032);
nand U9867 (N_9867,N_5377,N_6112);
or U9868 (N_9868,N_6756,N_5108);
and U9869 (N_9869,N_6284,N_5677);
nand U9870 (N_9870,N_6540,N_7488);
nor U9871 (N_9871,N_5008,N_6225);
nor U9872 (N_9872,N_7125,N_6043);
nor U9873 (N_9873,N_5107,N_6465);
and U9874 (N_9874,N_6706,N_7006);
or U9875 (N_9875,N_6115,N_5336);
nand U9876 (N_9876,N_5732,N_6149);
nand U9877 (N_9877,N_7450,N_6330);
nand U9878 (N_9878,N_6190,N_7174);
nand U9879 (N_9879,N_5832,N_7222);
and U9880 (N_9880,N_5802,N_7197);
nand U9881 (N_9881,N_6585,N_7035);
or U9882 (N_9882,N_5764,N_6252);
nand U9883 (N_9883,N_7457,N_7459);
nand U9884 (N_9884,N_6356,N_7015);
or U9885 (N_9885,N_7490,N_5305);
and U9886 (N_9886,N_6941,N_5554);
nor U9887 (N_9887,N_5962,N_6549);
nor U9888 (N_9888,N_6359,N_5177);
or U9889 (N_9889,N_5415,N_5928);
nand U9890 (N_9890,N_5661,N_6900);
xnor U9891 (N_9891,N_5876,N_5948);
nor U9892 (N_9892,N_7258,N_5643);
nand U9893 (N_9893,N_5189,N_6896);
and U9894 (N_9894,N_5633,N_5050);
xnor U9895 (N_9895,N_7167,N_7188);
or U9896 (N_9896,N_5217,N_5161);
nor U9897 (N_9897,N_7438,N_6061);
and U9898 (N_9898,N_7490,N_5071);
or U9899 (N_9899,N_5572,N_6556);
nand U9900 (N_9900,N_5651,N_6162);
nand U9901 (N_9901,N_5417,N_7136);
or U9902 (N_9902,N_6935,N_5746);
nor U9903 (N_9903,N_5916,N_7480);
or U9904 (N_9904,N_6176,N_5072);
nor U9905 (N_9905,N_5699,N_5313);
nor U9906 (N_9906,N_5377,N_5250);
nand U9907 (N_9907,N_5394,N_6493);
nor U9908 (N_9908,N_5104,N_5712);
nand U9909 (N_9909,N_5650,N_5186);
or U9910 (N_9910,N_6694,N_5669);
xor U9911 (N_9911,N_6048,N_5466);
and U9912 (N_9912,N_7385,N_6042);
and U9913 (N_9913,N_6363,N_6490);
or U9914 (N_9914,N_6406,N_5037);
nand U9915 (N_9915,N_6552,N_6615);
xor U9916 (N_9916,N_5832,N_6551);
nand U9917 (N_9917,N_7407,N_6645);
or U9918 (N_9918,N_7030,N_5710);
and U9919 (N_9919,N_6611,N_5358);
xor U9920 (N_9920,N_5076,N_5208);
xnor U9921 (N_9921,N_7091,N_5812);
or U9922 (N_9922,N_6295,N_7489);
nand U9923 (N_9923,N_6662,N_6745);
xnor U9924 (N_9924,N_5415,N_6123);
or U9925 (N_9925,N_6658,N_7199);
and U9926 (N_9926,N_6628,N_5511);
or U9927 (N_9927,N_6529,N_5948);
nand U9928 (N_9928,N_5423,N_7194);
nor U9929 (N_9929,N_6390,N_6583);
and U9930 (N_9930,N_6018,N_5836);
nor U9931 (N_9931,N_7387,N_5142);
or U9932 (N_9932,N_6066,N_7278);
xor U9933 (N_9933,N_6350,N_6309);
xnor U9934 (N_9934,N_5183,N_5189);
or U9935 (N_9935,N_5993,N_6351);
nor U9936 (N_9936,N_5993,N_6902);
and U9937 (N_9937,N_7057,N_6076);
nand U9938 (N_9938,N_6480,N_6660);
nor U9939 (N_9939,N_7417,N_6995);
and U9940 (N_9940,N_5467,N_5671);
nor U9941 (N_9941,N_5735,N_5732);
and U9942 (N_9942,N_5369,N_6136);
xor U9943 (N_9943,N_6584,N_7011);
nand U9944 (N_9944,N_5726,N_6055);
nor U9945 (N_9945,N_5084,N_6321);
xnor U9946 (N_9946,N_5423,N_6825);
xor U9947 (N_9947,N_6580,N_5847);
and U9948 (N_9948,N_7336,N_5699);
nand U9949 (N_9949,N_6068,N_6390);
or U9950 (N_9950,N_7056,N_5264);
nand U9951 (N_9951,N_7417,N_6692);
and U9952 (N_9952,N_5326,N_6472);
nand U9953 (N_9953,N_5086,N_5435);
nor U9954 (N_9954,N_6842,N_6102);
nor U9955 (N_9955,N_5352,N_6991);
and U9956 (N_9956,N_5390,N_7432);
nor U9957 (N_9957,N_6916,N_6227);
xnor U9958 (N_9958,N_5661,N_6537);
or U9959 (N_9959,N_5019,N_6292);
nand U9960 (N_9960,N_6125,N_5839);
and U9961 (N_9961,N_5468,N_6134);
or U9962 (N_9962,N_6820,N_6259);
or U9963 (N_9963,N_6137,N_7474);
or U9964 (N_9964,N_5317,N_5496);
nand U9965 (N_9965,N_6899,N_6884);
or U9966 (N_9966,N_7444,N_5369);
or U9967 (N_9967,N_5755,N_7046);
nand U9968 (N_9968,N_6749,N_6209);
nand U9969 (N_9969,N_5404,N_5505);
nand U9970 (N_9970,N_6396,N_5533);
and U9971 (N_9971,N_6120,N_6807);
xnor U9972 (N_9972,N_5009,N_5303);
nand U9973 (N_9973,N_6698,N_5379);
and U9974 (N_9974,N_6352,N_6564);
nor U9975 (N_9975,N_6613,N_7032);
or U9976 (N_9976,N_7204,N_6074);
xnor U9977 (N_9977,N_5188,N_5339);
xnor U9978 (N_9978,N_6827,N_6118);
nor U9979 (N_9979,N_6410,N_5503);
nand U9980 (N_9980,N_6554,N_6012);
or U9981 (N_9981,N_6324,N_7026);
nor U9982 (N_9982,N_6685,N_6878);
nand U9983 (N_9983,N_5193,N_5597);
nand U9984 (N_9984,N_5220,N_6145);
xnor U9985 (N_9985,N_5061,N_7106);
nor U9986 (N_9986,N_7286,N_6977);
and U9987 (N_9987,N_6834,N_7113);
and U9988 (N_9988,N_6103,N_7457);
and U9989 (N_9989,N_5708,N_6683);
nor U9990 (N_9990,N_5810,N_5149);
nand U9991 (N_9991,N_7143,N_5678);
nand U9992 (N_9992,N_6233,N_7249);
nand U9993 (N_9993,N_7227,N_5550);
and U9994 (N_9994,N_5912,N_6691);
nor U9995 (N_9995,N_7194,N_5589);
nand U9996 (N_9996,N_6325,N_7351);
and U9997 (N_9997,N_5125,N_5681);
xor U9998 (N_9998,N_5968,N_7208);
or U9999 (N_9999,N_6453,N_6455);
nor UO_0 (O_0,N_8304,N_8685);
and UO_1 (O_1,N_7572,N_7820);
and UO_2 (O_2,N_8284,N_8738);
nand UO_3 (O_3,N_9150,N_8130);
nor UO_4 (O_4,N_8034,N_8122);
nor UO_5 (O_5,N_8949,N_7748);
nand UO_6 (O_6,N_9620,N_7678);
and UO_7 (O_7,N_8927,N_9487);
nor UO_8 (O_8,N_9198,N_9878);
nor UO_9 (O_9,N_9762,N_9016);
xnor UO_10 (O_10,N_8178,N_8361);
xnor UO_11 (O_11,N_9910,N_9873);
and UO_12 (O_12,N_9583,N_7622);
nor UO_13 (O_13,N_7721,N_8409);
nand UO_14 (O_14,N_7999,N_8423);
nand UO_15 (O_15,N_9596,N_9521);
nand UO_16 (O_16,N_7755,N_7992);
or UO_17 (O_17,N_8978,N_9166);
nand UO_18 (O_18,N_8394,N_8355);
and UO_19 (O_19,N_7576,N_9268);
or UO_20 (O_20,N_7639,N_7938);
nand UO_21 (O_21,N_8031,N_8369);
nand UO_22 (O_22,N_8958,N_8070);
xnor UO_23 (O_23,N_8838,N_9880);
and UO_24 (O_24,N_9509,N_8216);
nor UO_25 (O_25,N_9669,N_9142);
nand UO_26 (O_26,N_9301,N_7757);
and UO_27 (O_27,N_7777,N_8297);
and UO_28 (O_28,N_8853,N_8990);
xor UO_29 (O_29,N_9175,N_8789);
nand UO_30 (O_30,N_9074,N_7890);
nor UO_31 (O_31,N_8171,N_7824);
nand UO_32 (O_32,N_8426,N_8454);
xor UO_33 (O_33,N_8580,N_8940);
and UO_34 (O_34,N_7926,N_7706);
or UO_35 (O_35,N_9203,N_8002);
xnor UO_36 (O_36,N_9085,N_8107);
xor UO_37 (O_37,N_9305,N_8470);
or UO_38 (O_38,N_9356,N_8415);
and UO_39 (O_39,N_8448,N_8189);
and UO_40 (O_40,N_7832,N_9946);
nand UO_41 (O_41,N_8324,N_8869);
nand UO_42 (O_42,N_7607,N_9050);
nand UO_43 (O_43,N_8167,N_8101);
or UO_44 (O_44,N_8310,N_9424);
or UO_45 (O_45,N_9133,N_9205);
or UO_46 (O_46,N_9459,N_8153);
or UO_47 (O_47,N_8270,N_8972);
xnor UO_48 (O_48,N_8053,N_9429);
nor UO_49 (O_49,N_7863,N_8458);
nor UO_50 (O_50,N_9895,N_8278);
nand UO_51 (O_51,N_9299,N_9963);
nor UO_52 (O_52,N_8022,N_9649);
or UO_53 (O_53,N_9043,N_9850);
and UO_54 (O_54,N_8911,N_7972);
xnor UO_55 (O_55,N_8509,N_7809);
and UO_56 (O_56,N_8992,N_8987);
nand UO_57 (O_57,N_9026,N_9921);
and UO_58 (O_58,N_7531,N_7903);
and UO_59 (O_59,N_8997,N_7897);
nand UO_60 (O_60,N_9892,N_9093);
nor UO_61 (O_61,N_8678,N_8281);
nor UO_62 (O_62,N_9621,N_7973);
nand UO_63 (O_63,N_8691,N_7808);
or UO_64 (O_64,N_9506,N_9474);
nand UO_65 (O_65,N_9564,N_8896);
xnor UO_66 (O_66,N_9397,N_8555);
or UO_67 (O_67,N_8761,N_7889);
or UO_68 (O_68,N_8592,N_8707);
and UO_69 (O_69,N_9333,N_8457);
xor UO_70 (O_70,N_8325,N_9049);
nor UO_71 (O_71,N_8844,N_8276);
nor UO_72 (O_72,N_7806,N_8078);
nor UO_73 (O_73,N_8859,N_9494);
nor UO_74 (O_74,N_8784,N_7522);
xnor UO_75 (O_75,N_9661,N_9915);
or UO_76 (O_76,N_8037,N_8337);
xor UO_77 (O_77,N_9064,N_8421);
and UO_78 (O_78,N_9469,N_8792);
nor UO_79 (O_79,N_9541,N_7759);
nor UO_80 (O_80,N_7770,N_9911);
nand UO_81 (O_81,N_8488,N_8150);
or UO_82 (O_82,N_9224,N_7711);
and UO_83 (O_83,N_9995,N_8957);
and UO_84 (O_84,N_8058,N_9556);
xor UO_85 (O_85,N_9206,N_7909);
nor UO_86 (O_86,N_7570,N_7830);
xor UO_87 (O_87,N_9088,N_9319);
nor UO_88 (O_88,N_9035,N_7841);
xor UO_89 (O_89,N_8025,N_9839);
and UO_90 (O_90,N_8030,N_9815);
nor UO_91 (O_91,N_9394,N_7730);
nand UO_92 (O_92,N_8502,N_8866);
or UO_93 (O_93,N_9021,N_8397);
xnor UO_94 (O_94,N_8287,N_7693);
and UO_95 (O_95,N_9633,N_9650);
nor UO_96 (O_96,N_9821,N_9163);
xor UO_97 (O_97,N_7971,N_9859);
nor UO_98 (O_98,N_8767,N_9270);
or UO_99 (O_99,N_8254,N_9691);
nand UO_100 (O_100,N_7778,N_8191);
xnor UO_101 (O_101,N_7835,N_8802);
or UO_102 (O_102,N_9876,N_8431);
nor UO_103 (O_103,N_8809,N_7612);
nor UO_104 (O_104,N_9410,N_8614);
nor UO_105 (O_105,N_8755,N_7557);
nand UO_106 (O_106,N_9265,N_9605);
or UO_107 (O_107,N_8742,N_9342);
nor UO_108 (O_108,N_9664,N_7794);
or UO_109 (O_109,N_8634,N_9805);
or UO_110 (O_110,N_7661,N_8664);
nor UO_111 (O_111,N_8979,N_8406);
and UO_112 (O_112,N_9518,N_9368);
or UO_113 (O_113,N_7705,N_9577);
nor UO_114 (O_114,N_9007,N_9926);
and UO_115 (O_115,N_7514,N_8237);
xnor UO_116 (O_116,N_9532,N_8001);
nand UO_117 (O_117,N_7967,N_8206);
or UO_118 (O_118,N_8374,N_8495);
or UO_119 (O_119,N_9369,N_9412);
or UO_120 (O_120,N_7513,N_7630);
or UO_121 (O_121,N_7592,N_8141);
nand UO_122 (O_122,N_8465,N_7923);
nor UO_123 (O_123,N_9399,N_8888);
or UO_124 (O_124,N_9787,N_9783);
nor UO_125 (O_125,N_8964,N_9826);
and UO_126 (O_126,N_9699,N_9767);
nand UO_127 (O_127,N_9427,N_9546);
nand UO_128 (O_128,N_8551,N_7985);
nand UO_129 (O_129,N_9652,N_8225);
nor UO_130 (O_130,N_8667,N_8959);
or UO_131 (O_131,N_8754,N_8375);
xnor UO_132 (O_132,N_9452,N_8867);
or UO_133 (O_133,N_9670,N_9889);
xnor UO_134 (O_134,N_8379,N_8647);
nand UO_135 (O_135,N_9219,N_9632);
nand UO_136 (O_136,N_9200,N_8644);
xnor UO_137 (O_137,N_7609,N_7663);
or UO_138 (O_138,N_7523,N_7695);
or UO_139 (O_139,N_8516,N_9920);
nand UO_140 (O_140,N_8079,N_7605);
xor UO_141 (O_141,N_8852,N_7520);
xnor UO_142 (O_142,N_8346,N_9018);
and UO_143 (O_143,N_8383,N_8921);
nor UO_144 (O_144,N_7907,N_9025);
nand UO_145 (O_145,N_9400,N_8474);
and UO_146 (O_146,N_8995,N_9491);
or UO_147 (O_147,N_8967,N_8543);
or UO_148 (O_148,N_8919,N_8800);
or UO_149 (O_149,N_7602,N_9638);
and UO_150 (O_150,N_9948,N_7785);
xor UO_151 (O_151,N_7656,N_8719);
nand UO_152 (O_152,N_9854,N_7707);
and UO_153 (O_153,N_7957,N_8968);
xor UO_154 (O_154,N_9260,N_9773);
nor UO_155 (O_155,N_7593,N_8412);
xnor UO_156 (O_156,N_8468,N_7944);
or UO_157 (O_157,N_9599,N_8271);
nand UO_158 (O_158,N_9906,N_8904);
and UO_159 (O_159,N_9257,N_8347);
nor UO_160 (O_160,N_8290,N_9034);
nand UO_161 (O_161,N_8732,N_9337);
nor UO_162 (O_162,N_9078,N_7750);
and UO_163 (O_163,N_8633,N_7573);
nor UO_164 (O_164,N_9625,N_9969);
nand UO_165 (O_165,N_9418,N_7819);
or UO_166 (O_166,N_9919,N_9843);
xnor UO_167 (O_167,N_9982,N_9330);
nand UO_168 (O_168,N_8105,N_7638);
xor UO_169 (O_169,N_9352,N_9197);
nand UO_170 (O_170,N_9309,N_7702);
and UO_171 (O_171,N_7932,N_9362);
xnor UO_172 (O_172,N_9724,N_9637);
xor UO_173 (O_173,N_7584,N_7600);
nand UO_174 (O_174,N_8492,N_8672);
nor UO_175 (O_175,N_9833,N_9101);
nand UO_176 (O_176,N_8577,N_7905);
xnor UO_177 (O_177,N_8975,N_8392);
nand UO_178 (O_178,N_9108,N_7917);
or UO_179 (O_179,N_7502,N_8293);
nand UO_180 (O_180,N_8386,N_8926);
and UO_181 (O_181,N_9832,N_7552);
nor UO_182 (O_182,N_7990,N_9312);
nor UO_183 (O_183,N_8452,N_9540);
and UO_184 (O_184,N_8675,N_8778);
xor UO_185 (O_185,N_8521,N_9485);
xor UO_186 (O_186,N_9226,N_8823);
nor UO_187 (O_187,N_7623,N_8545);
nor UO_188 (O_188,N_8760,N_7618);
or UO_189 (O_189,N_8312,N_9775);
xor UO_190 (O_190,N_9945,N_9811);
xor UO_191 (O_191,N_7673,N_8475);
nor UO_192 (O_192,N_8028,N_9283);
and UO_193 (O_193,N_8810,N_8948);
xnor UO_194 (O_194,N_7931,N_9961);
xnor UO_195 (O_195,N_7590,N_9313);
nor UO_196 (O_196,N_7616,N_7766);
nor UO_197 (O_197,N_9514,N_8039);
or UO_198 (O_198,N_7625,N_8011);
nand UO_199 (O_199,N_9598,N_9236);
and UO_200 (O_200,N_8095,N_7549);
nor UO_201 (O_201,N_7644,N_9128);
nand UO_202 (O_202,N_8944,N_8131);
or UO_203 (O_203,N_8624,N_7976);
xor UO_204 (O_204,N_7955,N_7634);
nand UO_205 (O_205,N_8352,N_7613);
nand UO_206 (O_206,N_9076,N_8531);
and UO_207 (O_207,N_9765,N_8885);
or UO_208 (O_208,N_9998,N_8152);
or UO_209 (O_209,N_7746,N_8725);
and UO_210 (O_210,N_8828,N_9324);
nand UO_211 (O_211,N_7650,N_8519);
or UO_212 (O_212,N_7936,N_8289);
nor UO_213 (O_213,N_8467,N_9974);
xnor UO_214 (O_214,N_8752,N_9111);
or UO_215 (O_215,N_7838,N_9851);
and UO_216 (O_216,N_8372,N_9802);
nor UO_217 (O_217,N_8963,N_8980);
nor UO_218 (O_218,N_7627,N_8422);
and UO_219 (O_219,N_8071,N_7945);
or UO_220 (O_220,N_7881,N_9067);
or UO_221 (O_221,N_8140,N_7561);
and UO_222 (O_222,N_9774,N_9992);
xor UO_223 (O_223,N_8656,N_9387);
nor UO_224 (O_224,N_9759,N_7655);
or UO_225 (O_225,N_7548,N_8484);
and UO_226 (O_226,N_9189,N_8326);
and UO_227 (O_227,N_8183,N_9462);
and UO_228 (O_228,N_7813,N_9803);
nand UO_229 (O_229,N_9655,N_9061);
xor UO_230 (O_230,N_7833,N_9897);
nand UO_231 (O_231,N_9235,N_8127);
xnor UO_232 (O_232,N_9210,N_9502);
nor UO_233 (O_233,N_9934,N_9334);
and UO_234 (O_234,N_7620,N_9628);
nand UO_235 (O_235,N_7534,N_9555);
nor UO_236 (O_236,N_8747,N_8512);
and UO_237 (O_237,N_8774,N_9698);
nand UO_238 (O_238,N_8615,N_8523);
xnor UO_239 (O_239,N_9656,N_7736);
or UO_240 (O_240,N_7867,N_7647);
nor UO_241 (O_241,N_9003,N_8597);
and UO_242 (O_242,N_8089,N_9580);
and UO_243 (O_243,N_8564,N_7871);
or UO_244 (O_244,N_7503,N_7798);
xor UO_245 (O_245,N_8834,N_9329);
and UO_246 (O_246,N_9073,N_9392);
and UO_247 (O_247,N_9592,N_8817);
xnor UO_248 (O_248,N_7743,N_8873);
xor UO_249 (O_249,N_8662,N_9668);
nor UO_250 (O_250,N_9456,N_9865);
nand UO_251 (O_251,N_8331,N_9090);
xnor UO_252 (O_252,N_9493,N_7723);
nand UO_253 (O_253,N_8323,N_8504);
or UO_254 (O_254,N_9616,N_7575);
nor UO_255 (O_255,N_8874,N_8164);
nand UO_256 (O_256,N_9228,N_9962);
or UO_257 (O_257,N_8500,N_8910);
xnor UO_258 (O_258,N_9708,N_9022);
or UO_259 (O_259,N_9856,N_7924);
nand UO_260 (O_260,N_9243,N_7574);
or UO_261 (O_261,N_7529,N_7551);
or UO_262 (O_262,N_9601,N_7733);
nand UO_263 (O_263,N_9534,N_8812);
nand UO_264 (O_264,N_7793,N_8762);
nor UO_265 (O_265,N_9574,N_8381);
nand UO_266 (O_266,N_8441,N_9566);
nor UO_267 (O_267,N_8632,N_8993);
or UO_268 (O_268,N_9320,N_9626);
nand UO_269 (O_269,N_7546,N_9173);
and UO_270 (O_270,N_8858,N_8234);
nor UO_271 (O_271,N_7828,N_9586);
nand UO_272 (O_272,N_8338,N_9565);
nand UO_273 (O_273,N_8170,N_7658);
xor UO_274 (O_274,N_8414,N_9239);
or UO_275 (O_275,N_7868,N_9692);
nand UO_276 (O_276,N_8538,N_8473);
nand UO_277 (O_277,N_8236,N_8768);
and UO_278 (O_278,N_9147,N_9100);
xor UO_279 (O_279,N_8906,N_7856);
nor UO_280 (O_280,N_9488,N_8539);
nor UO_281 (O_281,N_9285,N_8951);
and UO_282 (O_282,N_8933,N_9933);
and UO_283 (O_283,N_8086,N_9808);
or UO_284 (O_284,N_9753,N_9547);
and UO_285 (O_285,N_8791,N_9827);
nand UO_286 (O_286,N_9249,N_9001);
nand UO_287 (O_287,N_8845,N_8224);
nand UO_288 (O_288,N_9654,N_7904);
nor UO_289 (O_289,N_8561,N_8076);
nand UO_290 (O_290,N_9807,N_8110);
xor UO_291 (O_291,N_9194,N_8333);
nand UO_292 (O_292,N_7640,N_8388);
or UO_293 (O_293,N_7553,N_9868);
nor UO_294 (O_294,N_7862,N_8830);
nor UO_295 (O_295,N_8116,N_9888);
and UO_296 (O_296,N_9641,N_9983);
or UO_297 (O_297,N_8973,N_9593);
nor UO_298 (O_298,N_8204,N_8961);
or UO_299 (O_299,N_9501,N_9784);
and UO_300 (O_300,N_8166,N_9780);
xor UO_301 (O_301,N_7914,N_9582);
nor UO_302 (O_302,N_9894,N_9776);
or UO_303 (O_303,N_9202,N_9195);
or UO_304 (O_304,N_9576,N_9955);
nor UO_305 (O_305,N_7847,N_8720);
or UO_306 (O_306,N_7949,N_7802);
xnor UO_307 (O_307,N_8291,N_9719);
nand UO_308 (O_308,N_8090,N_8908);
and UO_309 (O_309,N_8981,N_8102);
nand UO_310 (O_310,N_9575,N_8407);
nand UO_311 (O_311,N_8833,N_8600);
or UO_312 (O_312,N_7935,N_8553);
or UO_313 (O_313,N_9823,N_7884);
nor UO_314 (O_314,N_8175,N_7900);
or UO_315 (O_315,N_8064,N_7950);
nand UO_316 (O_316,N_7933,N_9401);
and UO_317 (O_317,N_8401,N_7906);
and UO_318 (O_318,N_9156,N_9107);
or UO_319 (O_319,N_9659,N_8499);
nor UO_320 (O_320,N_7696,N_9588);
or UO_321 (O_321,N_9788,N_8408);
nand UO_322 (O_322,N_7916,N_9375);
and UO_323 (O_323,N_9937,N_9237);
and UO_324 (O_324,N_7727,N_9717);
or UO_325 (O_325,N_9267,N_8772);
nor UO_326 (O_326,N_9099,N_7921);
or UO_327 (O_327,N_7713,N_9480);
or UO_328 (O_328,N_8112,N_7586);
nor UO_329 (O_329,N_7687,N_8654);
and UO_330 (O_330,N_8673,N_9131);
nand UO_331 (O_331,N_8097,N_9662);
xnor UO_332 (O_332,N_8280,N_9567);
nand UO_333 (O_333,N_8188,N_8999);
nor UO_334 (O_334,N_9077,N_9928);
or UO_335 (O_335,N_7788,N_9442);
nand UO_336 (O_336,N_9478,N_8616);
or UO_337 (O_337,N_8410,N_8480);
xor UO_338 (O_338,N_9380,N_9475);
and UO_339 (O_339,N_9943,N_9302);
and UO_340 (O_340,N_9858,N_7734);
nor UO_341 (O_341,N_7568,N_9936);
nand UO_342 (O_342,N_7751,N_7608);
nor UO_343 (O_343,N_8962,N_8229);
and UO_344 (O_344,N_9510,N_8850);
nand UO_345 (O_345,N_8937,N_9680);
and UO_346 (O_346,N_8350,N_9054);
or UO_347 (O_347,N_8862,N_9371);
nor UO_348 (O_348,N_8142,N_7827);
and UO_349 (O_349,N_7732,N_9706);
and UO_350 (O_350,N_8455,N_8946);
nor UO_351 (O_351,N_9749,N_9490);
nand UO_352 (O_352,N_9709,N_8730);
and UO_353 (O_353,N_8416,N_7922);
xnor UO_354 (O_354,N_8476,N_9941);
nand UO_355 (O_355,N_8221,N_8590);
nor UO_356 (O_356,N_9460,N_9673);
and UO_357 (O_357,N_8340,N_8210);
or UO_358 (O_358,N_9925,N_9213);
and UO_359 (O_359,N_8514,N_7510);
nor UO_360 (O_360,N_9603,N_9682);
or UO_361 (O_361,N_8542,N_9527);
nand UO_362 (O_362,N_9095,N_8046);
nor UO_363 (O_363,N_8126,N_8601);
nand UO_364 (O_364,N_8299,N_8843);
nand UO_365 (O_365,N_9814,N_9700);
or UO_366 (O_366,N_8393,N_8091);
xnor UO_367 (O_367,N_9732,N_9996);
xnor UO_368 (O_368,N_8356,N_9451);
nor UO_369 (O_369,N_9120,N_8955);
nor UO_370 (O_370,N_7840,N_9848);
xor UO_371 (O_371,N_8629,N_9028);
nand UO_372 (O_372,N_8695,N_9862);
or UO_373 (O_373,N_9322,N_8207);
nor UO_374 (O_374,N_9595,N_9884);
and UO_375 (O_375,N_8200,N_9137);
and UO_376 (O_376,N_7594,N_9176);
xor UO_377 (O_377,N_9763,N_9572);
nor UO_378 (O_378,N_8118,N_8739);
or UO_379 (O_379,N_8439,N_9458);
nand UO_380 (O_380,N_9300,N_8839);
and UO_381 (O_381,N_8264,N_8971);
and UO_382 (O_382,N_9644,N_8851);
nor UO_383 (O_383,N_9461,N_9799);
xnor UO_384 (O_384,N_7920,N_7895);
nor UO_385 (O_385,N_8345,N_8259);
or UO_386 (O_386,N_9917,N_9123);
nand UO_387 (O_387,N_9689,N_9964);
nand UO_388 (O_388,N_7708,N_9870);
and UO_389 (O_389,N_9331,N_7740);
nor UO_390 (O_390,N_7589,N_9648);
and UO_391 (O_391,N_8365,N_9338);
or UO_392 (O_392,N_8686,N_7671);
or UO_393 (O_393,N_9005,N_7679);
xnor UO_394 (O_394,N_9531,N_8004);
nand UO_395 (O_395,N_9871,N_7547);
or UO_396 (O_396,N_8181,N_9845);
nand UO_397 (O_397,N_8428,N_8505);
nand UO_398 (O_398,N_8918,N_7617);
or UO_399 (O_399,N_9428,N_7857);
xnor UO_400 (O_400,N_9039,N_9242);
nor UO_401 (O_401,N_9256,N_8119);
nor UO_402 (O_402,N_7891,N_9558);
nand UO_403 (O_403,N_7698,N_9087);
xnor UO_404 (O_404,N_8821,N_9498);
nor UO_405 (O_405,N_8041,N_9212);
and UO_406 (O_406,N_7754,N_8782);
nand UO_407 (O_407,N_9341,N_8103);
and UO_408 (O_408,N_9466,N_8045);
nor UO_409 (O_409,N_9742,N_9473);
nor UO_410 (O_410,N_9161,N_9116);
and UO_411 (O_411,N_8773,N_9201);
or UO_412 (O_412,N_9144,N_7662);
nor UO_413 (O_413,N_9048,N_9070);
or UO_414 (O_414,N_8783,N_8787);
xnor UO_415 (O_415,N_8320,N_8696);
or UO_416 (O_416,N_8020,N_8708);
nand UO_417 (O_417,N_8035,N_7507);
nor UO_418 (O_418,N_9336,N_7980);
xnor UO_419 (O_419,N_8718,N_9752);
xor UO_420 (O_420,N_8269,N_8043);
and UO_421 (O_421,N_8947,N_9191);
and UO_422 (O_422,N_9777,N_7683);
nand UO_423 (O_423,N_8429,N_9993);
and UO_424 (O_424,N_8055,N_8630);
nor UO_425 (O_425,N_8871,N_9045);
or UO_426 (O_426,N_9126,N_7649);
xor UO_427 (O_427,N_8771,N_9011);
xor UO_428 (O_428,N_8576,N_9903);
xor UO_429 (O_429,N_8029,N_8316);
and UO_430 (O_430,N_7610,N_8628);
nor UO_431 (O_431,N_8741,N_9844);
xor UO_432 (O_432,N_9530,N_7844);
nand UO_433 (O_433,N_8935,N_7875);
xor UO_434 (O_434,N_8794,N_9609);
and UO_435 (O_435,N_8308,N_8536);
nand UO_436 (O_436,N_7714,N_9440);
and UO_437 (O_437,N_7697,N_7874);
nor UO_438 (O_438,N_8498,N_8256);
nand UO_439 (O_439,N_8349,N_8518);
or UO_440 (O_440,N_8060,N_9830);
nand UO_441 (O_441,N_9170,N_7816);
xnor UO_442 (O_442,N_8230,N_8641);
nor UO_443 (O_443,N_8905,N_7962);
nand UO_444 (O_444,N_8700,N_8884);
nor UO_445 (O_445,N_8405,N_9622);
xnor UO_446 (O_446,N_9952,N_8788);
xor UO_447 (O_447,N_8016,N_9817);
nor UO_448 (O_448,N_9745,N_9446);
nand UO_449 (O_449,N_9796,N_8562);
or UO_450 (O_450,N_8075,N_8477);
nand UO_451 (O_451,N_9232,N_7769);
nand UO_452 (O_452,N_8398,N_8625);
and UO_453 (O_453,N_8438,N_9340);
nand UO_454 (O_454,N_8286,N_9389);
or UO_455 (O_455,N_9711,N_8887);
nand UO_456 (O_456,N_7814,N_8436);
nand UO_457 (O_457,N_9317,N_9849);
nand UO_458 (O_458,N_9207,N_9524);
or UO_459 (O_459,N_9127,N_9764);
xnor UO_460 (O_460,N_8966,N_7684);
or UO_461 (O_461,N_9059,N_9396);
nand UO_462 (O_462,N_8334,N_7633);
or UO_463 (O_463,N_7850,N_8322);
and UO_464 (O_464,N_9979,N_8568);
xor UO_465 (O_465,N_9130,N_8098);
or UO_466 (O_466,N_9406,N_9223);
nand UO_467 (O_467,N_8440,N_7719);
nand UO_468 (O_468,N_7533,N_8595);
nor UO_469 (O_469,N_8668,N_8786);
nand UO_470 (O_470,N_7582,N_9227);
and UO_471 (O_471,N_7953,N_8897);
nor UO_472 (O_472,N_7578,N_9407);
or UO_473 (O_473,N_8367,N_9046);
or UO_474 (O_474,N_9104,N_9914);
xor UO_475 (O_475,N_7978,N_9657);
nor UO_476 (O_476,N_9877,N_8898);
xor UO_477 (O_477,N_8734,N_7887);
nor UO_478 (O_478,N_7803,N_7645);
xor UO_479 (O_479,N_8010,N_8424);
nor UO_480 (O_480,N_7970,N_7927);
or UO_481 (O_481,N_8915,N_8007);
or UO_482 (O_482,N_9768,N_8715);
xor UO_483 (O_483,N_8589,N_9949);
nand UO_484 (O_484,N_8649,N_9082);
nor UO_485 (O_485,N_9052,N_9636);
nor UO_486 (O_486,N_8261,N_8247);
xor UO_487 (O_487,N_8479,N_8879);
or UO_488 (O_488,N_8507,N_8177);
or UO_489 (O_489,N_8450,N_9879);
xor UO_490 (O_490,N_8661,N_9584);
xnor UO_491 (O_491,N_8396,N_9697);
or UO_492 (O_492,N_8218,N_9015);
nor UO_493 (O_493,N_8371,N_9756);
nor UO_494 (O_494,N_8681,N_8084);
xnor UO_495 (O_495,N_7739,N_9525);
or UO_496 (O_496,N_9716,N_8798);
xnor UO_497 (O_497,N_7928,N_7991);
xnor UO_498 (O_498,N_8960,N_8669);
and UO_499 (O_499,N_9307,N_8241);
nand UO_500 (O_500,N_9991,N_8179);
or UO_501 (O_501,N_9869,N_9994);
and UO_502 (O_502,N_9363,N_8108);
xnor UO_503 (O_503,N_9157,N_8954);
and UO_504 (O_504,N_7762,N_9890);
nor UO_505 (O_505,N_8330,N_9694);
xnor UO_506 (O_506,N_7982,N_8709);
nor UO_507 (O_507,N_8793,N_8377);
or UO_508 (O_508,N_8257,N_8307);
nand UO_509 (O_509,N_7526,N_8402);
nor UO_510 (O_510,N_9985,N_8242);
nand UO_511 (O_511,N_9225,N_7579);
or UO_512 (O_512,N_9276,N_8573);
xnor UO_513 (O_513,N_9684,N_9570);
or UO_514 (O_514,N_8743,N_9230);
nor UO_515 (O_515,N_7604,N_9448);
or UO_516 (O_516,N_7758,N_8087);
nor UO_517 (O_517,N_8113,N_7654);
and UO_518 (O_518,N_7699,N_9281);
or UO_519 (O_519,N_9613,N_9721);
and UO_520 (O_520,N_7675,N_9304);
nor UO_521 (O_521,N_8217,N_8511);
nand UO_522 (O_522,N_9036,N_9997);
xor UO_523 (O_523,N_7682,N_9678);
nor UO_524 (O_524,N_7641,N_9187);
and UO_525 (O_525,N_7786,N_9071);
nand UO_526 (O_526,N_8750,N_8129);
nor UO_527 (O_527,N_9326,N_8052);
nor UO_528 (O_528,N_9735,N_8014);
nor UO_529 (O_529,N_9450,N_9186);
nand UO_530 (O_530,N_9980,N_9190);
nand UO_531 (O_531,N_8248,N_8391);
or UO_532 (O_532,N_7524,N_8985);
xnor UO_533 (O_533,N_8796,N_9172);
nor UO_534 (O_534,N_8635,N_7521);
or UO_535 (O_535,N_7815,N_8889);
nor UO_536 (O_536,N_9477,N_8094);
xnor UO_537 (O_537,N_7930,N_9792);
and UO_538 (O_538,N_7587,N_7911);
and UO_539 (O_539,N_8418,N_8593);
nor UO_540 (O_540,N_8917,N_8048);
and UO_541 (O_541,N_8849,N_7776);
or UO_542 (O_542,N_8565,N_8305);
nor UO_543 (O_543,N_8588,N_8827);
nand UO_544 (O_544,N_9439,N_8988);
xnor UO_545 (O_545,N_8584,N_8653);
nand UO_546 (O_546,N_8881,N_8132);
and UO_547 (O_547,N_9838,N_8120);
or UO_548 (O_548,N_9351,N_8213);
xor UO_549 (O_549,N_7948,N_8517);
nand UO_550 (O_550,N_8180,N_7729);
and UO_551 (O_551,N_7525,N_8527);
and UO_552 (O_552,N_8702,N_9081);
xor UO_553 (O_553,N_8779,N_9885);
nand UO_554 (O_554,N_8503,N_8366);
and UO_555 (O_555,N_7724,N_8706);
xor UO_556 (O_556,N_8157,N_9350);
nand UO_557 (O_557,N_7913,N_9132);
xor UO_558 (O_558,N_9437,N_9967);
and UO_559 (O_559,N_9492,N_8042);
or UO_560 (O_560,N_8886,N_7753);
or UO_561 (O_561,N_8655,N_8268);
xor UO_562 (O_562,N_9316,N_7961);
nor UO_563 (O_563,N_7792,N_9470);
xnor UO_564 (O_564,N_9275,N_9159);
xor UO_565 (O_565,N_9989,N_8574);
nand UO_566 (O_566,N_8541,N_9271);
and UO_567 (O_567,N_8883,N_8209);
and UO_568 (O_568,N_9748,N_8425);
nand UO_569 (O_569,N_9481,N_8208);
nor UO_570 (O_570,N_8831,N_8697);
nor UO_571 (O_571,N_9155,N_8930);
or UO_572 (O_572,N_8463,N_9743);
nand UO_573 (O_573,N_8748,N_8876);
nor UO_574 (O_574,N_8701,N_9602);
xnor UO_575 (O_575,N_8544,N_9209);
nor UO_576 (O_576,N_8343,N_8163);
nor UO_577 (O_577,N_9710,N_9794);
xnor UO_578 (O_578,N_8563,N_9381);
xnor UO_579 (O_579,N_7852,N_7888);
or UO_580 (O_580,N_8901,N_7709);
nand UO_581 (O_581,N_8059,N_8515);
and UO_582 (O_582,N_9266,N_7508);
xnor UO_583 (O_583,N_9391,N_7883);
xor UO_584 (O_584,N_9364,N_7989);
xor UO_585 (O_585,N_9746,N_9800);
xor UO_586 (O_586,N_8795,N_7519);
and UO_587 (O_587,N_9965,N_7628);
nand UO_588 (O_588,N_9672,N_8018);
nor UO_589 (O_589,N_8722,N_9578);
xor UO_590 (O_590,N_7756,N_8818);
xnor UO_591 (O_591,N_9589,N_7943);
nor UO_592 (O_592,N_9294,N_8645);
or UO_593 (O_593,N_7642,N_9703);
and UO_594 (O_594,N_8914,N_9809);
xor UO_595 (O_595,N_9479,N_8050);
xor UO_596 (O_596,N_7692,N_8162);
nor UO_597 (O_597,N_8279,N_9904);
nand UO_598 (O_598,N_8459,N_8219);
xor UO_599 (O_599,N_8262,N_8533);
nand UO_600 (O_600,N_8606,N_8596);
or UO_601 (O_601,N_7912,N_7870);
or UO_602 (O_602,N_7563,N_9528);
nor UO_603 (O_603,N_8857,N_9246);
nor UO_604 (O_604,N_8864,N_7660);
nand UO_605 (O_605,N_7763,N_8952);
nor UO_606 (O_606,N_8547,N_8165);
and UO_607 (O_607,N_8688,N_7865);
nor UO_608 (O_608,N_7836,N_8865);
or UO_609 (O_609,N_9519,N_8860);
and UO_610 (O_610,N_8769,N_8203);
and UO_611 (O_611,N_8199,N_9109);
nand UO_612 (O_612,N_8353,N_9030);
xor UO_613 (O_613,N_8520,N_9353);
nor UO_614 (O_614,N_9679,N_9426);
or UO_615 (O_615,N_9563,N_9922);
nor UO_616 (O_616,N_8038,N_9660);
xnor UO_617 (O_617,N_7860,N_9058);
nand UO_618 (O_618,N_9504,N_8335);
and UO_619 (O_619,N_8724,N_7528);
nand UO_620 (O_620,N_9083,N_9515);
and UO_621 (O_621,N_8665,N_8639);
nor UO_622 (O_622,N_8348,N_8583);
nor UO_623 (O_623,N_9215,N_8658);
nand UO_624 (O_624,N_9629,N_9663);
nand UO_625 (O_625,N_7672,N_7918);
and UO_626 (O_626,N_8689,N_9931);
nand UO_627 (O_627,N_7861,N_9395);
or UO_628 (O_628,N_9112,N_8902);
nor UO_629 (O_629,N_8462,N_9486);
nor UO_630 (O_630,N_9913,N_8451);
nand UO_631 (O_631,N_9413,N_8676);
nand UO_632 (O_632,N_9269,N_9549);
nand UO_633 (O_633,N_9117,N_8273);
nor UO_634 (O_634,N_8481,N_8840);
nor UO_635 (O_635,N_7540,N_9483);
nor UO_636 (O_636,N_7542,N_9600);
or UO_637 (O_637,N_8413,N_8005);
xnor UO_638 (O_638,N_8690,N_8073);
xor UO_639 (O_639,N_8938,N_8526);
and UO_640 (O_640,N_7843,N_9024);
nand UO_641 (O_641,N_7984,N_9402);
or UO_642 (O_642,N_7772,N_8560);
nor UO_643 (O_643,N_9542,N_9094);
nand UO_644 (O_644,N_9292,N_9944);
nand UO_645 (O_645,N_9345,N_7700);
nor UO_646 (O_646,N_9523,N_8461);
or UO_647 (O_647,N_9614,N_8556);
nand UO_648 (O_648,N_8378,N_9141);
xor UO_649 (O_649,N_9562,N_8442);
and UO_650 (O_650,N_9444,N_8096);
and UO_651 (O_651,N_8244,N_9261);
nand UO_652 (O_652,N_8106,N_8026);
nor UO_653 (O_653,N_8220,N_8837);
nand UO_654 (O_654,N_9503,N_8801);
or UO_655 (O_655,N_8699,N_8671);
and UO_656 (O_656,N_7664,N_9891);
or UO_657 (O_657,N_9465,N_9376);
nor UO_658 (O_658,N_9177,N_8023);
or UO_659 (O_659,N_7738,N_7580);
or UO_660 (O_660,N_9781,N_8846);
and UO_661 (O_661,N_7761,N_8184);
and UO_662 (O_662,N_8161,N_8117);
nand UO_663 (O_663,N_8296,N_8913);
nand UO_664 (O_664,N_7960,N_7747);
nand UO_665 (O_665,N_8427,N_8306);
or UO_666 (O_666,N_9947,N_7799);
xor UO_667 (O_667,N_9548,N_8744);
xnor UO_668 (O_668,N_9702,N_7516);
or UO_669 (O_669,N_8493,N_8233);
and UO_670 (O_670,N_9537,N_8693);
nor UO_671 (O_671,N_8925,N_8956);
nor UO_672 (O_672,N_9386,N_8626);
nand UO_673 (O_673,N_8047,N_8197);
and UO_674 (O_674,N_7968,N_7822);
or UO_675 (O_675,N_8820,N_9611);
or UO_676 (O_676,N_8751,N_8186);
or UO_677 (O_677,N_7670,N_7997);
nor UO_678 (O_678,N_8790,N_9725);
and UO_679 (O_679,N_9545,N_9184);
or UO_680 (O_680,N_9357,N_7939);
xnor UO_681 (O_681,N_8922,N_9647);
nand UO_682 (O_682,N_8524,N_7725);
xnor UO_683 (O_683,N_9896,N_8062);
nand UO_684 (O_684,N_9347,N_9365);
and UO_685 (O_685,N_7872,N_8613);
and UO_686 (O_686,N_8258,N_8471);
xor UO_687 (O_687,N_7996,N_9612);
or UO_688 (O_688,N_9244,N_7964);
and UO_689 (O_689,N_9060,N_8781);
nand UO_690 (O_690,N_9430,N_8737);
and UO_691 (O_691,N_8530,N_8943);
nor UO_692 (O_692,N_8728,N_7876);
xnor UO_693 (O_693,N_7742,N_7937);
and UO_694 (O_694,N_9252,N_9097);
xor UO_695 (O_695,N_9771,N_7681);
nand UO_696 (O_696,N_8315,N_9960);
and UO_697 (O_697,N_9355,N_7790);
xor UO_698 (O_698,N_8021,N_9069);
and UO_699 (O_699,N_7886,N_8109);
nand UO_700 (O_700,N_7998,N_7812);
and UO_701 (O_701,N_9758,N_8115);
or UO_702 (O_702,N_8970,N_9075);
xor UO_703 (O_703,N_8637,N_9000);
xnor UO_704 (O_704,N_9544,N_8721);
nand UO_705 (O_705,N_8942,N_9907);
nor UO_706 (O_706,N_9033,N_7779);
or UO_707 (O_707,N_9431,N_8100);
xnor UO_708 (O_708,N_9383,N_8483);
nand UO_709 (O_709,N_8766,N_9199);
nor UO_710 (O_710,N_7637,N_9066);
and UO_711 (O_711,N_8074,N_8239);
xor UO_712 (O_712,N_8912,N_7784);
or UO_713 (O_713,N_9790,N_9935);
or UO_714 (O_714,N_9306,N_9938);
nor UO_715 (O_715,N_8657,N_9831);
nand UO_716 (O_716,N_8627,N_9146);
xor UO_717 (O_717,N_8806,N_8138);
nor UO_718 (O_718,N_8878,N_9522);
xnor UO_719 (O_719,N_7532,N_7885);
and UO_720 (O_720,N_9220,N_9010);
or UO_721 (O_721,N_8160,N_9538);
or UO_722 (O_722,N_8246,N_9640);
and UO_723 (O_723,N_9388,N_8133);
or UO_724 (O_724,N_7715,N_7818);
nand UO_725 (O_725,N_9398,N_7577);
or UO_726 (O_726,N_8068,N_9866);
xor UO_727 (O_727,N_7983,N_8085);
or UO_728 (O_728,N_9273,N_7596);
and UO_729 (O_729,N_8128,N_9098);
xor UO_730 (O_730,N_9860,N_9986);
nor UO_731 (O_731,N_8674,N_9651);
nor UO_732 (O_732,N_9118,N_8599);
nor UO_733 (O_733,N_9789,N_8240);
and UO_734 (O_734,N_8227,N_9667);
and UO_735 (O_735,N_7652,N_8077);
xor UO_736 (O_736,N_9553,N_8013);
or UO_737 (O_737,N_7800,N_9032);
nor UO_738 (O_738,N_7512,N_8569);
and UO_739 (O_739,N_8469,N_9134);
nor UO_740 (O_740,N_7690,N_9733);
nor UO_741 (O_741,N_7873,N_7804);
nor UO_742 (O_742,N_8648,N_9886);
and UO_743 (O_743,N_7544,N_9349);
nor UO_744 (O_744,N_8618,N_9004);
nand UO_745 (O_745,N_7538,N_8650);
nor UO_746 (O_746,N_9560,N_7810);
xnor UO_747 (O_747,N_8733,N_8067);
or UO_748 (O_748,N_9722,N_9581);
nand UO_749 (O_749,N_7632,N_7974);
xor UO_750 (O_750,N_8003,N_8591);
nand UO_751 (O_751,N_8159,N_9436);
xor UO_752 (O_752,N_8698,N_8072);
xnor UO_753 (O_753,N_7929,N_9231);
xnor UO_754 (O_754,N_7554,N_9348);
and UO_755 (O_755,N_8757,N_9314);
or UO_756 (O_756,N_8249,N_9325);
and UO_757 (O_757,N_9536,N_8567);
nor UO_758 (O_758,N_8359,N_9852);
and UO_759 (O_759,N_9976,N_7829);
and UO_760 (O_760,N_8735,N_9009);
or UO_761 (O_761,N_8890,N_8403);
xor UO_762 (O_762,N_8855,N_7817);
nor UO_763 (O_763,N_8172,N_8252);
nor UO_764 (O_764,N_9042,N_8581);
xnor UO_765 (O_765,N_8430,N_8080);
nand UO_766 (O_766,N_9115,N_8151);
nor UO_767 (O_767,N_9853,N_8065);
and UO_768 (O_768,N_8711,N_7560);
xor UO_769 (O_769,N_8731,N_8342);
nand UO_770 (O_770,N_9624,N_9013);
nor UO_771 (O_771,N_9533,N_8033);
or UO_772 (O_772,N_9740,N_9898);
nand UO_773 (O_773,N_9056,N_7774);
xor UO_774 (O_774,N_9438,N_9234);
and UO_775 (O_775,N_8525,N_9551);
nor UO_776 (O_776,N_8063,N_9723);
and UO_777 (O_777,N_9152,N_9623);
nor UO_778 (O_778,N_7963,N_8929);
nand UO_779 (O_779,N_8907,N_9591);
or UO_780 (O_780,N_8336,N_9443);
or UO_781 (O_781,N_8989,N_8198);
or UO_782 (O_782,N_8222,N_7855);
and UO_783 (O_783,N_7651,N_8449);
xnor UO_784 (O_784,N_8621,N_9818);
nor UO_785 (O_785,N_9044,N_7966);
and UO_786 (O_786,N_8548,N_7559);
nor UO_787 (O_787,N_8327,N_7601);
nor UO_788 (O_788,N_8288,N_7737);
xnor UO_789 (O_789,N_8099,N_9950);
or UO_790 (O_790,N_9053,N_9286);
and UO_791 (O_791,N_8807,N_9323);
nor UO_792 (O_792,N_7694,N_8494);
or UO_793 (O_793,N_9883,N_9008);
nand UO_794 (O_794,N_8243,N_9359);
and UO_795 (O_795,N_8532,N_8417);
xor UO_796 (O_796,N_9403,N_9966);
or UO_797 (O_797,N_9959,N_8093);
or UO_798 (O_798,N_8704,N_8826);
and UO_799 (O_799,N_9597,N_9747);
nand UO_800 (O_800,N_9810,N_8255);
nor UO_801 (O_801,N_7643,N_8124);
xnor UO_802 (O_802,N_9124,N_8996);
and UO_803 (O_803,N_7501,N_7537);
nand UO_804 (O_804,N_8104,N_9881);
and UO_805 (O_805,N_7915,N_9148);
xnor UO_806 (O_806,N_7745,N_8508);
or UO_807 (O_807,N_7511,N_8684);
or UO_808 (O_808,N_8158,N_7946);
nor UO_809 (O_809,N_9457,N_8575);
nand UO_810 (O_810,N_8554,N_9739);
or UO_811 (O_811,N_8585,N_9579);
nor UO_812 (O_812,N_7987,N_9425);
and UO_813 (O_813,N_9264,N_9068);
or UO_814 (O_814,N_9610,N_8017);
xnor UO_815 (O_815,N_8566,N_8620);
nand UO_816 (O_816,N_7635,N_8842);
nand UO_817 (O_817,N_8559,N_8212);
or UO_818 (O_818,N_9916,N_9842);
nor UO_819 (O_819,N_8856,N_9315);
nor UO_820 (O_820,N_8603,N_7712);
nand UO_821 (O_821,N_9185,N_9728);
xor UO_822 (O_822,N_9918,N_8998);
xor UO_823 (O_823,N_7826,N_9585);
or UO_824 (O_824,N_8491,N_8156);
xnor UO_825 (O_825,N_7752,N_7898);
and UO_826 (O_826,N_7947,N_8266);
nor UO_827 (O_827,N_9681,N_8182);
or UO_828 (O_828,N_8265,N_7995);
nor UO_829 (O_829,N_9954,N_8420);
xor UO_830 (O_830,N_9183,N_9683);
and UO_831 (O_831,N_8572,N_9408);
or UO_832 (O_832,N_8019,N_8344);
nand UO_833 (O_833,N_9837,N_9151);
or UO_834 (O_834,N_8253,N_7823);
nand UO_835 (O_835,N_8008,N_7615);
and UO_836 (O_836,N_9674,N_9893);
or UO_837 (O_837,N_9715,N_8916);
or UO_838 (O_838,N_9639,N_7956);
nor UO_839 (O_839,N_9455,N_9779);
nor UO_840 (O_840,N_7965,N_8765);
and UO_841 (O_841,N_9037,N_9454);
or UO_842 (O_842,N_7564,N_9245);
and UO_843 (O_843,N_7717,N_9816);
nor UO_844 (O_844,N_8804,N_8753);
nand UO_845 (O_845,N_9409,N_9686);
nand UO_846 (O_846,N_8066,N_7530);
nor UO_847 (O_847,N_7731,N_7811);
xnor UO_848 (O_848,N_9824,N_7864);
nor UO_849 (O_849,N_9882,N_7515);
nor UO_850 (O_850,N_9114,N_9987);
and UO_851 (O_851,N_8594,N_9806);
xor UO_852 (O_852,N_8139,N_9978);
nor UO_853 (O_853,N_8135,N_8749);
nor UO_854 (O_854,N_8623,N_8622);
nor UO_855 (O_855,N_7767,N_9182);
or UO_856 (O_856,N_8435,N_8612);
nor UO_857 (O_857,N_8051,N_9813);
and UO_858 (O_858,N_9463,N_9511);
and UO_859 (O_859,N_7506,N_7545);
and UO_860 (O_860,N_8535,N_8380);
or UO_861 (O_861,N_8144,N_9778);
nand UO_862 (O_862,N_9750,N_8797);
nand UO_863 (O_863,N_7680,N_7787);
or UO_864 (O_864,N_8302,N_8587);
or UO_865 (O_865,N_7934,N_9772);
and UO_866 (O_866,N_8364,N_9559);
xnor UO_867 (O_867,N_8666,N_7969);
and UO_868 (O_868,N_8598,N_8301);
nor UO_869 (O_869,N_8756,N_8083);
xnor UO_870 (O_870,N_8939,N_7773);
xnor UO_871 (O_871,N_8329,N_9432);
nand UO_872 (O_872,N_9366,N_7597);
and UO_873 (O_873,N_7704,N_9180);
nor UO_874 (O_874,N_9761,N_9981);
nand UO_875 (O_875,N_9404,N_8211);
and UO_876 (O_876,N_9179,N_8444);
nor UO_877 (O_877,N_9296,N_9687);
and UO_878 (O_878,N_8683,N_9160);
xor UO_879 (O_879,N_9631,N_9496);
xor UO_880 (O_880,N_7646,N_9607);
or UO_881 (O_881,N_9119,N_8608);
nor UO_882 (O_882,N_9367,N_8282);
and UO_883 (O_883,N_9887,N_9378);
or UO_884 (O_884,N_9630,N_8892);
nand UO_885 (O_885,N_8125,N_8486);
or UO_886 (O_886,N_9384,N_9358);
or UO_887 (O_887,N_9619,N_9744);
nand UO_888 (O_888,N_7569,N_9754);
nor UO_889 (O_889,N_8389,N_7555);
or UO_890 (O_890,N_8456,N_9422);
and UO_891 (O_891,N_9178,N_9932);
nand UO_892 (O_892,N_9247,N_9958);
xor UO_893 (O_893,N_8447,N_9217);
nand UO_894 (O_894,N_8991,N_7797);
nand UO_895 (O_895,N_9984,N_9293);
and UO_896 (O_896,N_9701,N_9676);
nand UO_897 (O_897,N_8149,N_8311);
nor UO_898 (O_898,N_9909,N_8318);
or UO_899 (O_899,N_7741,N_8799);
nand UO_900 (O_900,N_9704,N_9828);
or UO_901 (O_901,N_9819,N_8640);
nand UO_902 (O_902,N_8636,N_7866);
nand UO_903 (O_903,N_7701,N_7505);
nor UO_904 (O_904,N_7676,N_7849);
and UO_905 (O_905,N_9760,N_8351);
xor UO_906 (O_906,N_9712,N_7626);
and UO_907 (O_907,N_8974,N_8716);
nand UO_908 (O_908,N_8169,N_9321);
or UO_909 (O_909,N_7710,N_9973);
nand UO_910 (O_910,N_7993,N_9797);
nand UO_911 (O_911,N_7581,N_9901);
nor UO_912 (O_912,N_7703,N_9730);
nand UO_913 (O_913,N_9867,N_9872);
nor UO_914 (O_914,N_9065,N_9096);
xor UO_915 (O_915,N_9214,N_9568);
or UO_916 (O_916,N_7896,N_7979);
and UO_917 (O_917,N_7839,N_8872);
xor UO_918 (O_918,N_8054,N_8358);
nor UO_919 (O_919,N_7614,N_8829);
xnor UO_920 (O_920,N_9604,N_8482);
or UO_921 (O_921,N_8832,N_7735);
nand UO_922 (O_922,N_8920,N_8670);
nand UO_923 (O_923,N_9014,N_9335);
nand UO_924 (O_924,N_9646,N_9497);
nor UO_925 (O_925,N_7893,N_9900);
and UO_926 (O_926,N_8819,N_8522);
and UO_927 (O_927,N_9829,N_8501);
or UO_928 (O_928,N_9310,N_8437);
nor UO_929 (O_929,N_7795,N_9635);
or UO_930 (O_930,N_7831,N_8317);
or UO_931 (O_931,N_9343,N_8745);
nand UO_932 (O_932,N_9606,N_8434);
and UO_933 (O_933,N_8808,N_7940);
nand UO_934 (O_934,N_7556,N_7571);
nand UO_935 (O_935,N_9047,N_8868);
nor UO_936 (O_936,N_9543,N_7674);
and UO_937 (O_937,N_9433,N_9379);
or UO_938 (O_938,N_8215,N_9507);
nand UO_939 (O_939,N_9370,N_8936);
nor UO_940 (O_940,N_9573,N_9218);
xnor UO_941 (O_941,N_8009,N_8703);
or UO_942 (O_942,N_8609,N_8319);
xnor UO_943 (O_943,N_9940,N_8663);
and UO_944 (O_944,N_9972,N_7668);
or UO_945 (O_945,N_8238,N_9766);
and UO_946 (O_946,N_8506,N_8057);
xor UO_947 (O_947,N_9377,N_7859);
or UO_948 (O_948,N_8148,N_8231);
nand UO_949 (O_949,N_7858,N_8710);
nor UO_950 (O_950,N_9658,N_8891);
nand UO_951 (O_951,N_9467,N_9221);
and UO_952 (O_952,N_9726,N_7869);
xor UO_953 (O_953,N_8466,N_8726);
and UO_954 (O_954,N_8578,N_7942);
xor UO_955 (O_955,N_7728,N_8549);
nor UO_956 (O_956,N_7718,N_8321);
and UO_957 (O_957,N_7853,N_9590);
xnor UO_958 (O_958,N_9287,N_8770);
and UO_959 (O_959,N_9529,N_9405);
xor UO_960 (O_960,N_8400,N_8376);
xor UO_961 (O_961,N_8899,N_9103);
nor UO_962 (O_962,N_7951,N_9977);
or UO_963 (O_963,N_8646,N_9012);
nand UO_964 (O_964,N_7854,N_8540);
xor UO_965 (O_965,N_9279,N_8740);
xnor UO_966 (O_966,N_8373,N_9923);
xnor UO_967 (O_967,N_9645,N_8309);
or UO_968 (O_968,N_9499,N_8677);
nand UO_969 (O_969,N_8478,N_9145);
xor UO_970 (O_970,N_7583,N_8485);
nand UO_971 (O_971,N_9617,N_8195);
xnor UO_972 (O_972,N_9193,N_7603);
or UO_973 (O_973,N_9263,N_9516);
nand UO_974 (O_974,N_9262,N_7821);
xnor UO_975 (O_975,N_8300,N_8777);
and UO_976 (O_976,N_8994,N_9091);
nor UO_977 (O_977,N_9168,N_8387);
nand UO_978 (O_978,N_9255,N_9360);
and UO_979 (O_979,N_7726,N_9027);
nand UO_980 (O_980,N_9693,N_9204);
nand UO_981 (O_981,N_9079,N_9453);
xor UO_982 (O_982,N_9902,N_8283);
nor UO_983 (O_983,N_8419,N_8193);
or UO_984 (O_984,N_9734,N_8953);
nor UO_985 (O_985,N_8497,N_8510);
xor UO_986 (O_986,N_7606,N_7877);
or UO_987 (O_987,N_7902,N_9258);
xnor UO_988 (O_988,N_9642,N_8235);
nand UO_989 (O_989,N_7848,N_7958);
and UO_990 (O_990,N_8390,N_7517);
xor UO_991 (O_991,N_9957,N_9930);
or UO_992 (O_992,N_7901,N_8605);
xor UO_993 (O_993,N_8489,N_7621);
xor UO_994 (O_994,N_9653,N_7975);
xor UO_995 (O_995,N_8875,N_9062);
or UO_996 (O_996,N_8529,N_8679);
and UO_997 (O_997,N_7768,N_9627);
and UO_998 (O_998,N_7686,N_9970);
nand UO_999 (O_999,N_8550,N_8713);
and UO_1000 (O_1000,N_9441,N_7539);
and UO_1001 (O_1001,N_9738,N_9372);
xor UO_1002 (O_1002,N_8443,N_8969);
xnor UO_1003 (O_1003,N_9041,N_9092);
or UO_1004 (O_1004,N_9484,N_9513);
nor UO_1005 (O_1005,N_9741,N_7988);
nor UO_1006 (O_1006,N_7925,N_8123);
nand UO_1007 (O_1007,N_9690,N_8805);
nor UO_1008 (O_1008,N_8174,N_8934);
or UO_1009 (O_1009,N_8145,N_9956);
nor UO_1010 (O_1010,N_9415,N_7631);
nand UO_1011 (O_1011,N_9770,N_9374);
or UO_1012 (O_1012,N_7845,N_8931);
nand UO_1013 (O_1013,N_9373,N_9019);
nor UO_1014 (O_1014,N_8558,N_8362);
nand UO_1015 (O_1015,N_9786,N_8205);
nand UO_1016 (O_1016,N_9587,N_8012);
nor UO_1017 (O_1017,N_7527,N_8006);
nand UO_1018 (O_1018,N_8775,N_9793);
nor UO_1019 (O_1019,N_7807,N_7892);
nand UO_1020 (O_1020,N_8736,N_8490);
xor UO_1021 (O_1021,N_8764,N_8354);
xor UO_1022 (O_1022,N_7882,N_7994);
and UO_1023 (O_1023,N_9526,N_9393);
and UO_1024 (O_1024,N_9951,N_7880);
nor UO_1025 (O_1025,N_9594,N_7760);
nor UO_1026 (O_1026,N_8863,N_8617);
or UO_1027 (O_1027,N_9251,N_7744);
and UO_1028 (O_1028,N_9705,N_8395);
or UO_1029 (O_1029,N_8909,N_8638);
nor UO_1030 (O_1030,N_7624,N_9971);
and UO_1031 (O_1031,N_8313,N_8976);
xor UO_1032 (O_1032,N_9057,N_8445);
or UO_1033 (O_1033,N_8134,N_9905);
xor UO_1034 (O_1034,N_9086,N_9102);
xnor UO_1035 (O_1035,N_7567,N_9822);
xnor UO_1036 (O_1036,N_9924,N_7591);
or UO_1037 (O_1037,N_8604,N_7691);
and UO_1038 (O_1038,N_8399,N_9846);
nand UO_1039 (O_1039,N_7598,N_8571);
nand UO_1040 (O_1040,N_8295,N_8557);
xor UO_1041 (O_1041,N_8176,N_8611);
or UO_1042 (O_1042,N_8277,N_8586);
or UO_1043 (O_1043,N_8232,N_9332);
and UO_1044 (O_1044,N_7941,N_9927);
and UO_1045 (O_1045,N_8651,N_8294);
nor UO_1046 (O_1046,N_9051,N_8496);
xnor UO_1047 (O_1047,N_8056,N_8924);
nor UO_1048 (O_1048,N_9464,N_9942);
nor UO_1049 (O_1049,N_9233,N_8986);
and UO_1050 (O_1050,N_8245,N_7796);
xor UO_1051 (O_1051,N_9171,N_9106);
nand UO_1052 (O_1052,N_7535,N_7749);
and UO_1053 (O_1053,N_9755,N_7986);
nand UO_1054 (O_1054,N_8895,N_8552);
or UO_1055 (O_1055,N_9571,N_8723);
nor UO_1056 (O_1056,N_9288,N_8835);
or UO_1057 (O_1057,N_8214,N_9143);
nand UO_1058 (O_1058,N_8061,N_9411);
nand UO_1059 (O_1059,N_8652,N_8848);
nor UO_1060 (O_1060,N_7782,N_9423);
and UO_1061 (O_1061,N_8088,N_8404);
nand UO_1062 (O_1062,N_9713,N_8446);
or UO_1063 (O_1063,N_8111,N_8759);
nand UO_1064 (O_1064,N_9714,N_9737);
nor UO_1065 (O_1065,N_8570,N_8460);
nor UO_1066 (O_1066,N_9471,N_9278);
xor UO_1067 (O_1067,N_8758,N_9346);
nor UO_1068 (O_1068,N_8928,N_8032);
nand UO_1069 (O_1069,N_9089,N_7837);
nand UO_1070 (O_1070,N_9677,N_9517);
and UO_1071 (O_1071,N_9181,N_8274);
xnor UO_1072 (O_1072,N_9855,N_8965);
nor UO_1073 (O_1073,N_8984,N_9561);
nor UO_1074 (O_1074,N_9718,N_8729);
or UO_1075 (O_1075,N_8870,N_9736);
xnor UO_1076 (O_1076,N_8015,N_9836);
xnor UO_1077 (O_1077,N_7666,N_8487);
xnor UO_1078 (O_1078,N_9554,N_9825);
nor UO_1079 (O_1079,N_7765,N_8841);
nor UO_1080 (O_1080,N_7780,N_7834);
nor UO_1081 (O_1081,N_8411,N_8785);
or UO_1082 (O_1082,N_9557,N_8339);
or UO_1083 (O_1083,N_7894,N_8546);
or UO_1084 (O_1084,N_9216,N_8121);
nor UO_1085 (O_1085,N_8223,N_8537);
or UO_1086 (O_1086,N_8082,N_8154);
nand UO_1087 (O_1087,N_9248,N_9552);
and UO_1088 (O_1088,N_8534,N_7977);
xnor UO_1089 (O_1089,N_8528,N_9149);
nand UO_1090 (O_1090,N_8024,N_9472);
nor UO_1091 (O_1091,N_9291,N_9311);
and UO_1092 (O_1092,N_7899,N_7783);
and UO_1093 (O_1093,N_7541,N_8298);
or UO_1094 (O_1094,N_8822,N_7716);
or UO_1095 (O_1095,N_8187,N_7509);
or UO_1096 (O_1096,N_8602,N_9158);
or UO_1097 (O_1097,N_8464,N_9055);
xnor UO_1098 (O_1098,N_7775,N_8982);
nand UO_1099 (O_1099,N_9500,N_9318);
and UO_1100 (O_1100,N_7665,N_9449);
or UO_1101 (O_1101,N_9820,N_9020);
nor UO_1102 (O_1102,N_8582,N_7504);
and UO_1103 (O_1103,N_7669,N_8267);
or UO_1104 (O_1104,N_8824,N_9468);
xnor UO_1105 (O_1105,N_8854,N_8341);
nor UO_1106 (O_1106,N_8923,N_7908);
xor UO_1107 (O_1107,N_9153,N_8146);
nand UO_1108 (O_1108,N_7952,N_9259);
xor UO_1109 (O_1109,N_9666,N_9414);
nand UO_1110 (O_1110,N_7959,N_9696);
nand UO_1111 (O_1111,N_8660,N_9953);
nand UO_1112 (O_1112,N_8137,N_9801);
and UO_1113 (O_1113,N_8303,N_8983);
nor UO_1114 (O_1114,N_7565,N_9720);
and UO_1115 (O_1115,N_9512,N_8363);
or UO_1116 (O_1116,N_8292,N_9295);
nand UO_1117 (O_1117,N_9508,N_8977);
or UO_1118 (O_1118,N_9912,N_9282);
nand UO_1119 (O_1119,N_9447,N_9272);
nor UO_1120 (O_1120,N_8894,N_9361);
xnor UO_1121 (O_1121,N_8000,N_8780);
or UO_1122 (O_1122,N_9121,N_9382);
xnor UO_1123 (O_1123,N_8357,N_9834);
or UO_1124 (O_1124,N_8114,N_7689);
nand UO_1125 (O_1125,N_9421,N_9841);
nand UO_1126 (O_1126,N_8285,N_8275);
and UO_1127 (O_1127,N_7878,N_9253);
xnor UO_1128 (O_1128,N_8714,N_9795);
nand UO_1129 (O_1129,N_7566,N_9135);
nor UO_1130 (O_1130,N_8368,N_7518);
and UO_1131 (O_1131,N_9812,N_8027);
nand UO_1132 (O_1132,N_9241,N_8717);
or UO_1133 (O_1133,N_9274,N_9290);
or UO_1134 (O_1134,N_7720,N_9634);
nand UO_1135 (O_1135,N_8360,N_9804);
xnor UO_1136 (O_1136,N_9875,N_9847);
nor UO_1137 (O_1137,N_8816,N_9791);
and UO_1138 (O_1138,N_7789,N_9729);
or UO_1139 (O_1139,N_8384,N_7550);
or UO_1140 (O_1140,N_8190,N_8069);
xnor UO_1141 (O_1141,N_9419,N_8903);
and UO_1142 (O_1142,N_7842,N_9999);
or UO_1143 (O_1143,N_9857,N_8776);
nand UO_1144 (O_1144,N_7619,N_9136);
nand UO_1145 (O_1145,N_9861,N_8185);
or UO_1146 (O_1146,N_9476,N_8049);
nand UO_1147 (O_1147,N_7910,N_8836);
nor UO_1148 (O_1148,N_7851,N_8155);
nor UO_1149 (O_1149,N_9864,N_8950);
xor UO_1150 (O_1150,N_9250,N_9615);
and UO_1151 (O_1151,N_9238,N_8932);
or UO_1152 (O_1152,N_9113,N_9038);
nand UO_1153 (O_1153,N_9297,N_9167);
nand UO_1154 (O_1154,N_9988,N_7648);
and UO_1155 (O_1155,N_8472,N_8202);
and UO_1156 (O_1156,N_9874,N_9328);
xnor UO_1157 (O_1157,N_9782,N_9188);
xnor UO_1158 (O_1158,N_9863,N_8382);
or UO_1159 (O_1159,N_7585,N_8705);
and UO_1160 (O_1160,N_7500,N_9229);
and UO_1161 (O_1161,N_9608,N_7825);
nand UO_1162 (O_1162,N_7879,N_9665);
or UO_1163 (O_1163,N_8260,N_9105);
xor UO_1164 (O_1164,N_8201,N_8513);
xor UO_1165 (O_1165,N_9435,N_9174);
nand UO_1166 (O_1166,N_7919,N_8147);
xor UO_1167 (O_1167,N_9929,N_7599);
nand UO_1168 (O_1168,N_9169,N_9339);
or UO_1169 (O_1169,N_9284,N_9416);
nor UO_1170 (O_1170,N_9125,N_7558);
nand UO_1171 (O_1171,N_7685,N_9769);
and UO_1172 (O_1172,N_9618,N_9489);
nor UO_1173 (O_1173,N_9192,N_8036);
nor UO_1174 (O_1174,N_7791,N_8228);
nor UO_1175 (O_1175,N_8811,N_7688);
nor UO_1176 (O_1176,N_9162,N_8194);
nor UO_1177 (O_1177,N_7981,N_9550);
nand UO_1178 (O_1178,N_9417,N_8941);
nand UO_1179 (O_1179,N_8814,N_9505);
nor UO_1180 (O_1180,N_9727,N_9434);
and UO_1181 (O_1181,N_8880,N_9344);
xnor UO_1182 (O_1182,N_9165,N_8370);
or UO_1183 (O_1183,N_8813,N_9327);
or UO_1184 (O_1184,N_9196,N_8196);
xnor UO_1185 (O_1185,N_8694,N_8803);
nor UO_1186 (O_1186,N_9240,N_9643);
nor UO_1187 (O_1187,N_8680,N_7801);
nand UO_1188 (O_1188,N_9006,N_8040);
xnor UO_1189 (O_1189,N_9899,N_7536);
nand UO_1190 (O_1190,N_7629,N_9569);
or UO_1191 (O_1191,N_8092,N_9110);
and UO_1192 (O_1192,N_7667,N_8081);
nor UO_1193 (O_1193,N_9688,N_7954);
xor UO_1194 (O_1194,N_8847,N_9695);
xor UO_1195 (O_1195,N_8619,N_9445);
and UO_1196 (O_1196,N_8861,N_9029);
nor UO_1197 (O_1197,N_9154,N_9390);
xor UO_1198 (O_1198,N_7677,N_9539);
xnor UO_1199 (O_1199,N_9798,N_8825);
nor UO_1200 (O_1200,N_9040,N_7543);
or UO_1201 (O_1201,N_9208,N_9254);
nor UO_1202 (O_1202,N_7805,N_8272);
xor UO_1203 (O_1203,N_8250,N_9731);
and UO_1204 (O_1204,N_8877,N_9002);
or UO_1205 (O_1205,N_9280,N_7722);
nor UO_1206 (O_1206,N_9685,N_8692);
nor UO_1207 (O_1207,N_9671,N_8251);
nand UO_1208 (O_1208,N_9140,N_9482);
xor UO_1209 (O_1209,N_7659,N_9975);
nand UO_1210 (O_1210,N_9990,N_8882);
nor UO_1211 (O_1211,N_9751,N_7764);
or UO_1212 (O_1212,N_8727,N_8746);
nor UO_1213 (O_1213,N_9298,N_9084);
nor UO_1214 (O_1214,N_9211,N_7653);
or UO_1215 (O_1215,N_8893,N_8610);
nand UO_1216 (O_1216,N_8044,N_8643);
and UO_1217 (O_1217,N_9031,N_9495);
nor UO_1218 (O_1218,N_9420,N_8453);
nand UO_1219 (O_1219,N_7562,N_8385);
nor UO_1220 (O_1220,N_8642,N_9080);
and UO_1221 (O_1221,N_8143,N_9063);
nor UO_1222 (O_1222,N_8226,N_8263);
or UO_1223 (O_1223,N_8173,N_8314);
and UO_1224 (O_1224,N_9908,N_9277);
nand UO_1225 (O_1225,N_8945,N_9675);
and UO_1226 (O_1226,N_9385,N_9222);
nor UO_1227 (O_1227,N_8168,N_8332);
xor UO_1228 (O_1228,N_9535,N_9939);
nor UO_1229 (O_1229,N_7611,N_7781);
and UO_1230 (O_1230,N_9785,N_8631);
xor UO_1231 (O_1231,N_7771,N_9520);
nand UO_1232 (O_1232,N_9138,N_8607);
and UO_1233 (O_1233,N_9840,N_9164);
nand UO_1234 (O_1234,N_9968,N_8900);
nor UO_1235 (O_1235,N_9129,N_9122);
nor UO_1236 (O_1236,N_8815,N_8433);
or UO_1237 (O_1237,N_9303,N_8682);
nand UO_1238 (O_1238,N_9707,N_9139);
nand UO_1239 (O_1239,N_9835,N_8328);
nand UO_1240 (O_1240,N_7595,N_7846);
or UO_1241 (O_1241,N_8763,N_9289);
nand UO_1242 (O_1242,N_8659,N_7588);
nor UO_1243 (O_1243,N_8687,N_9354);
xor UO_1244 (O_1244,N_9023,N_7657);
or UO_1245 (O_1245,N_7636,N_8192);
and UO_1246 (O_1246,N_9072,N_8136);
and UO_1247 (O_1247,N_9308,N_9757);
nor UO_1248 (O_1248,N_9017,N_8579);
nor UO_1249 (O_1249,N_8432,N_8712);
and UO_1250 (O_1250,N_9885,N_7646);
nor UO_1251 (O_1251,N_8748,N_7504);
and UO_1252 (O_1252,N_7787,N_8703);
nand UO_1253 (O_1253,N_7864,N_9133);
and UO_1254 (O_1254,N_8892,N_9185);
xor UO_1255 (O_1255,N_8583,N_8367);
or UO_1256 (O_1256,N_9276,N_9462);
and UO_1257 (O_1257,N_8039,N_9059);
or UO_1258 (O_1258,N_9835,N_7920);
xnor UO_1259 (O_1259,N_9368,N_7549);
nand UO_1260 (O_1260,N_7783,N_8997);
xnor UO_1261 (O_1261,N_7777,N_8909);
and UO_1262 (O_1262,N_7596,N_7550);
nand UO_1263 (O_1263,N_8853,N_9776);
and UO_1264 (O_1264,N_9836,N_8642);
and UO_1265 (O_1265,N_7878,N_9496);
nor UO_1266 (O_1266,N_9809,N_8182);
xor UO_1267 (O_1267,N_8115,N_8097);
or UO_1268 (O_1268,N_7697,N_8162);
and UO_1269 (O_1269,N_7733,N_7968);
xnor UO_1270 (O_1270,N_9703,N_9363);
and UO_1271 (O_1271,N_8684,N_9897);
and UO_1272 (O_1272,N_8617,N_9056);
xnor UO_1273 (O_1273,N_8787,N_8193);
and UO_1274 (O_1274,N_9955,N_9404);
nand UO_1275 (O_1275,N_8365,N_8247);
nor UO_1276 (O_1276,N_7666,N_8166);
nand UO_1277 (O_1277,N_9266,N_9428);
and UO_1278 (O_1278,N_9815,N_8588);
nor UO_1279 (O_1279,N_9892,N_8703);
and UO_1280 (O_1280,N_9389,N_8730);
xor UO_1281 (O_1281,N_9238,N_9913);
and UO_1282 (O_1282,N_9726,N_8125);
and UO_1283 (O_1283,N_8043,N_9244);
xnor UO_1284 (O_1284,N_9479,N_9217);
and UO_1285 (O_1285,N_9811,N_8339);
or UO_1286 (O_1286,N_8176,N_7948);
nand UO_1287 (O_1287,N_9505,N_8443);
and UO_1288 (O_1288,N_9571,N_7959);
nor UO_1289 (O_1289,N_9026,N_9670);
or UO_1290 (O_1290,N_8110,N_9420);
nand UO_1291 (O_1291,N_8795,N_8031);
and UO_1292 (O_1292,N_8103,N_9059);
xor UO_1293 (O_1293,N_7905,N_9160);
or UO_1294 (O_1294,N_7600,N_8148);
and UO_1295 (O_1295,N_9166,N_8920);
and UO_1296 (O_1296,N_7737,N_8968);
nor UO_1297 (O_1297,N_8662,N_9703);
xnor UO_1298 (O_1298,N_8473,N_8772);
and UO_1299 (O_1299,N_7695,N_8656);
and UO_1300 (O_1300,N_7510,N_9481);
and UO_1301 (O_1301,N_8719,N_8787);
nor UO_1302 (O_1302,N_9915,N_8949);
or UO_1303 (O_1303,N_8398,N_9902);
or UO_1304 (O_1304,N_8397,N_9888);
nand UO_1305 (O_1305,N_8482,N_7872);
nor UO_1306 (O_1306,N_8383,N_9535);
nand UO_1307 (O_1307,N_9165,N_8012);
or UO_1308 (O_1308,N_8200,N_9128);
xnor UO_1309 (O_1309,N_8322,N_8173);
nor UO_1310 (O_1310,N_8397,N_8212);
or UO_1311 (O_1311,N_8476,N_7596);
nand UO_1312 (O_1312,N_7596,N_8121);
nand UO_1313 (O_1313,N_9577,N_9517);
nor UO_1314 (O_1314,N_7958,N_9686);
xor UO_1315 (O_1315,N_8674,N_8247);
nor UO_1316 (O_1316,N_8539,N_8770);
nor UO_1317 (O_1317,N_9669,N_9368);
and UO_1318 (O_1318,N_9206,N_7591);
xor UO_1319 (O_1319,N_9750,N_9125);
nor UO_1320 (O_1320,N_8977,N_9634);
nor UO_1321 (O_1321,N_9923,N_9675);
nor UO_1322 (O_1322,N_9947,N_9723);
or UO_1323 (O_1323,N_9951,N_8633);
nor UO_1324 (O_1324,N_8854,N_9637);
or UO_1325 (O_1325,N_9852,N_7742);
nand UO_1326 (O_1326,N_9160,N_8982);
nor UO_1327 (O_1327,N_8291,N_8517);
nor UO_1328 (O_1328,N_8551,N_9337);
xnor UO_1329 (O_1329,N_7977,N_8450);
xor UO_1330 (O_1330,N_8004,N_7801);
and UO_1331 (O_1331,N_8939,N_8410);
nor UO_1332 (O_1332,N_9283,N_8215);
or UO_1333 (O_1333,N_7975,N_9202);
xor UO_1334 (O_1334,N_8899,N_9722);
and UO_1335 (O_1335,N_9357,N_9445);
xnor UO_1336 (O_1336,N_8176,N_9965);
nor UO_1337 (O_1337,N_9453,N_7846);
and UO_1338 (O_1338,N_7807,N_8278);
nor UO_1339 (O_1339,N_8334,N_8795);
or UO_1340 (O_1340,N_9759,N_7548);
nand UO_1341 (O_1341,N_8150,N_8516);
and UO_1342 (O_1342,N_9644,N_8963);
or UO_1343 (O_1343,N_8019,N_9736);
and UO_1344 (O_1344,N_7841,N_9897);
nor UO_1345 (O_1345,N_9130,N_7658);
or UO_1346 (O_1346,N_8446,N_9535);
nor UO_1347 (O_1347,N_8732,N_8294);
nor UO_1348 (O_1348,N_8081,N_9344);
nor UO_1349 (O_1349,N_9976,N_9315);
or UO_1350 (O_1350,N_8039,N_8017);
nand UO_1351 (O_1351,N_9402,N_8859);
and UO_1352 (O_1352,N_9745,N_9217);
xor UO_1353 (O_1353,N_8218,N_9068);
nor UO_1354 (O_1354,N_7567,N_8359);
nor UO_1355 (O_1355,N_8241,N_7530);
nor UO_1356 (O_1356,N_7677,N_9951);
and UO_1357 (O_1357,N_9501,N_7588);
xor UO_1358 (O_1358,N_9680,N_9762);
nor UO_1359 (O_1359,N_7610,N_9188);
xor UO_1360 (O_1360,N_8728,N_8928);
or UO_1361 (O_1361,N_8788,N_7844);
nor UO_1362 (O_1362,N_8398,N_7902);
or UO_1363 (O_1363,N_7721,N_9077);
or UO_1364 (O_1364,N_8579,N_9070);
nor UO_1365 (O_1365,N_8095,N_7509);
and UO_1366 (O_1366,N_8596,N_7931);
nand UO_1367 (O_1367,N_9083,N_8369);
nor UO_1368 (O_1368,N_8261,N_8954);
nor UO_1369 (O_1369,N_9417,N_8620);
xnor UO_1370 (O_1370,N_8325,N_8664);
or UO_1371 (O_1371,N_8185,N_8475);
nor UO_1372 (O_1372,N_9234,N_8035);
or UO_1373 (O_1373,N_9929,N_7786);
nor UO_1374 (O_1374,N_9953,N_8307);
and UO_1375 (O_1375,N_8280,N_8814);
and UO_1376 (O_1376,N_7682,N_7972);
xor UO_1377 (O_1377,N_9032,N_9582);
xnor UO_1378 (O_1378,N_9782,N_8803);
xor UO_1379 (O_1379,N_9879,N_8257);
nand UO_1380 (O_1380,N_9397,N_7975);
or UO_1381 (O_1381,N_8271,N_8038);
or UO_1382 (O_1382,N_8654,N_7532);
and UO_1383 (O_1383,N_9660,N_9882);
or UO_1384 (O_1384,N_7986,N_9715);
or UO_1385 (O_1385,N_9115,N_8766);
and UO_1386 (O_1386,N_8178,N_8035);
or UO_1387 (O_1387,N_9780,N_9272);
and UO_1388 (O_1388,N_9616,N_8140);
nand UO_1389 (O_1389,N_9548,N_7963);
or UO_1390 (O_1390,N_9010,N_8081);
or UO_1391 (O_1391,N_8331,N_7529);
or UO_1392 (O_1392,N_8552,N_9679);
or UO_1393 (O_1393,N_9051,N_7817);
nand UO_1394 (O_1394,N_8319,N_9057);
or UO_1395 (O_1395,N_8284,N_7925);
and UO_1396 (O_1396,N_9445,N_7572);
or UO_1397 (O_1397,N_9570,N_9874);
nor UO_1398 (O_1398,N_9992,N_9649);
xor UO_1399 (O_1399,N_7762,N_8646);
nor UO_1400 (O_1400,N_9079,N_8981);
nor UO_1401 (O_1401,N_8055,N_8988);
nor UO_1402 (O_1402,N_9821,N_9813);
nand UO_1403 (O_1403,N_7733,N_8864);
and UO_1404 (O_1404,N_9026,N_8229);
nor UO_1405 (O_1405,N_8663,N_8181);
or UO_1406 (O_1406,N_8447,N_8775);
xnor UO_1407 (O_1407,N_8023,N_9778);
nand UO_1408 (O_1408,N_9795,N_9595);
nand UO_1409 (O_1409,N_8152,N_9820);
nand UO_1410 (O_1410,N_8673,N_7832);
and UO_1411 (O_1411,N_9172,N_8893);
nand UO_1412 (O_1412,N_8505,N_9145);
nor UO_1413 (O_1413,N_8752,N_8715);
nand UO_1414 (O_1414,N_8973,N_7824);
xor UO_1415 (O_1415,N_8763,N_8271);
xnor UO_1416 (O_1416,N_8020,N_7581);
nand UO_1417 (O_1417,N_7581,N_8497);
nand UO_1418 (O_1418,N_7874,N_9119);
or UO_1419 (O_1419,N_9339,N_8802);
and UO_1420 (O_1420,N_8858,N_9341);
or UO_1421 (O_1421,N_8190,N_9237);
nand UO_1422 (O_1422,N_9842,N_8808);
or UO_1423 (O_1423,N_8523,N_9316);
nor UO_1424 (O_1424,N_9483,N_8967);
nand UO_1425 (O_1425,N_8852,N_8141);
nor UO_1426 (O_1426,N_8994,N_8063);
nand UO_1427 (O_1427,N_7572,N_9410);
nand UO_1428 (O_1428,N_9789,N_8863);
nor UO_1429 (O_1429,N_8141,N_8792);
nand UO_1430 (O_1430,N_9936,N_9003);
and UO_1431 (O_1431,N_7589,N_8083);
xnor UO_1432 (O_1432,N_9909,N_9834);
or UO_1433 (O_1433,N_9736,N_8058);
nand UO_1434 (O_1434,N_7928,N_8338);
nor UO_1435 (O_1435,N_7948,N_9451);
nand UO_1436 (O_1436,N_9141,N_9544);
nor UO_1437 (O_1437,N_7851,N_9176);
and UO_1438 (O_1438,N_8969,N_9321);
or UO_1439 (O_1439,N_7798,N_9437);
or UO_1440 (O_1440,N_8438,N_7674);
nand UO_1441 (O_1441,N_7716,N_7537);
xnor UO_1442 (O_1442,N_9908,N_9086);
or UO_1443 (O_1443,N_8422,N_9627);
xor UO_1444 (O_1444,N_9390,N_7561);
nor UO_1445 (O_1445,N_8246,N_9244);
or UO_1446 (O_1446,N_9512,N_9650);
xor UO_1447 (O_1447,N_8424,N_9598);
nor UO_1448 (O_1448,N_8369,N_9620);
nor UO_1449 (O_1449,N_8311,N_8771);
nor UO_1450 (O_1450,N_8738,N_9916);
or UO_1451 (O_1451,N_7627,N_9825);
and UO_1452 (O_1452,N_7717,N_9100);
nand UO_1453 (O_1453,N_9171,N_8715);
and UO_1454 (O_1454,N_9323,N_8507);
nand UO_1455 (O_1455,N_7560,N_8419);
or UO_1456 (O_1456,N_7954,N_9573);
or UO_1457 (O_1457,N_8258,N_7928);
xnor UO_1458 (O_1458,N_9462,N_9003);
nand UO_1459 (O_1459,N_7770,N_7894);
nor UO_1460 (O_1460,N_7610,N_9038);
nor UO_1461 (O_1461,N_9848,N_7849);
nand UO_1462 (O_1462,N_7518,N_9400);
xor UO_1463 (O_1463,N_9490,N_8764);
and UO_1464 (O_1464,N_9254,N_7596);
nand UO_1465 (O_1465,N_8844,N_8339);
nand UO_1466 (O_1466,N_7755,N_8949);
nor UO_1467 (O_1467,N_9065,N_9163);
or UO_1468 (O_1468,N_8941,N_9188);
xnor UO_1469 (O_1469,N_9654,N_8688);
and UO_1470 (O_1470,N_8641,N_8171);
and UO_1471 (O_1471,N_7940,N_8540);
nand UO_1472 (O_1472,N_8258,N_8229);
nand UO_1473 (O_1473,N_9914,N_8881);
and UO_1474 (O_1474,N_8888,N_9717);
or UO_1475 (O_1475,N_9259,N_7824);
nand UO_1476 (O_1476,N_7551,N_7957);
xor UO_1477 (O_1477,N_7886,N_7843);
nand UO_1478 (O_1478,N_9117,N_7825);
or UO_1479 (O_1479,N_8441,N_9298);
or UO_1480 (O_1480,N_9116,N_9261);
and UO_1481 (O_1481,N_7749,N_8673);
nor UO_1482 (O_1482,N_9174,N_9669);
nand UO_1483 (O_1483,N_8607,N_7655);
and UO_1484 (O_1484,N_9347,N_9120);
or UO_1485 (O_1485,N_7662,N_7675);
nand UO_1486 (O_1486,N_9133,N_7653);
nand UO_1487 (O_1487,N_7642,N_7871);
nand UO_1488 (O_1488,N_7891,N_9443);
and UO_1489 (O_1489,N_9555,N_8244);
nor UO_1490 (O_1490,N_9309,N_9352);
nand UO_1491 (O_1491,N_9652,N_8545);
or UO_1492 (O_1492,N_7993,N_9924);
nand UO_1493 (O_1493,N_9257,N_7902);
xor UO_1494 (O_1494,N_8412,N_9582);
nor UO_1495 (O_1495,N_7778,N_8239);
xnor UO_1496 (O_1496,N_7823,N_8993);
or UO_1497 (O_1497,N_8727,N_8182);
or UO_1498 (O_1498,N_9713,N_9265);
nand UO_1499 (O_1499,N_8213,N_8881);
endmodule