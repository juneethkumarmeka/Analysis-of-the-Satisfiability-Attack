module basic_2000_20000_2500_50_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
and U0 (N_0,In_1085,In_803);
nand U1 (N_1,In_720,In_395);
and U2 (N_2,In_340,In_876);
xnor U3 (N_3,In_1467,In_813);
xor U4 (N_4,In_1028,In_1519);
xnor U5 (N_5,In_1144,In_424);
nand U6 (N_6,In_1379,In_236);
or U7 (N_7,In_899,In_1751);
or U8 (N_8,In_1084,In_1096);
nor U9 (N_9,In_1732,In_1559);
and U10 (N_10,In_452,In_621);
or U11 (N_11,In_515,In_1564);
and U12 (N_12,In_1723,In_1216);
nand U13 (N_13,In_1730,In_276);
and U14 (N_14,In_1582,In_506);
or U15 (N_15,In_1907,In_956);
nand U16 (N_16,In_1572,In_687);
or U17 (N_17,In_1857,In_1166);
nor U18 (N_18,In_192,In_40);
nand U19 (N_19,In_1703,In_1674);
xnor U20 (N_20,In_1836,In_894);
and U21 (N_21,In_841,In_309);
and U22 (N_22,In_1460,In_1081);
and U23 (N_23,In_485,In_835);
and U24 (N_24,In_405,In_1055);
xnor U25 (N_25,In_130,In_298);
nand U26 (N_26,In_187,In_1910);
nor U27 (N_27,In_241,In_102);
or U28 (N_28,In_1710,In_1009);
and U29 (N_29,In_781,In_863);
nor U30 (N_30,In_1265,In_42);
xnor U31 (N_31,In_1436,In_1391);
nor U32 (N_32,In_618,In_1491);
and U33 (N_33,In_604,In_29);
and U34 (N_34,In_944,In_1626);
xor U35 (N_35,In_1652,In_231);
nor U36 (N_36,In_567,In_1145);
nand U37 (N_37,In_1715,In_126);
xnor U38 (N_38,In_1845,In_1252);
nand U39 (N_39,In_305,In_287);
and U40 (N_40,In_80,In_250);
xor U41 (N_41,In_1134,In_1059);
xnor U42 (N_42,In_145,In_1975);
and U43 (N_43,In_908,In_1697);
or U44 (N_44,In_367,In_638);
xor U45 (N_45,In_1686,In_1414);
nor U46 (N_46,In_1413,In_1895);
nand U47 (N_47,In_437,In_1048);
and U48 (N_48,In_408,In_232);
and U49 (N_49,In_693,In_1945);
nor U50 (N_50,In_1223,In_1879);
xor U51 (N_51,In_1184,In_1397);
nand U52 (N_52,In_186,In_1533);
nor U53 (N_53,In_691,In_1405);
nor U54 (N_54,In_1797,In_1357);
nor U55 (N_55,In_1555,In_632);
or U56 (N_56,In_627,In_1725);
or U57 (N_57,In_1951,In_1329);
or U58 (N_58,In_643,In_449);
nand U59 (N_59,In_1146,In_1658);
nor U60 (N_60,In_1936,In_1767);
nand U61 (N_61,In_740,In_1347);
or U62 (N_62,In_1915,In_1562);
xor U63 (N_63,In_312,In_25);
and U64 (N_64,In_1129,In_1455);
or U65 (N_65,In_936,In_1692);
nor U66 (N_66,In_226,In_353);
and U67 (N_67,In_1181,In_1236);
xnor U68 (N_68,In_1113,In_158);
nand U69 (N_69,In_205,In_1257);
and U70 (N_70,In_37,In_1416);
and U71 (N_71,In_1976,In_496);
nand U72 (N_72,In_1784,In_216);
and U73 (N_73,In_734,In_1142);
nor U74 (N_74,In_1655,In_923);
and U75 (N_75,In_1735,In_1040);
xor U76 (N_76,In_1380,In_625);
nor U77 (N_77,In_749,In_297);
and U78 (N_78,In_934,In_1523);
xnor U79 (N_79,In_1728,In_458);
or U80 (N_80,In_1809,In_922);
and U81 (N_81,In_724,In_1622);
xnor U82 (N_82,In_817,In_262);
nand U83 (N_83,In_1140,In_255);
nand U84 (N_84,In_1638,In_417);
or U85 (N_85,In_436,In_1851);
nor U86 (N_86,In_1322,In_1624);
xor U87 (N_87,In_1772,In_1100);
xnor U88 (N_88,In_704,In_514);
or U89 (N_89,In_958,In_1004);
and U90 (N_90,In_845,In_1822);
xnor U91 (N_91,In_1923,In_1516);
nand U92 (N_92,In_731,In_1779);
nor U93 (N_93,In_1326,In_1891);
and U94 (N_94,In_591,In_1813);
nor U95 (N_95,In_628,In_359);
or U96 (N_96,In_131,In_717);
or U97 (N_97,In_669,In_681);
nor U98 (N_98,In_872,In_1886);
nor U99 (N_99,In_1261,In_1003);
and U100 (N_100,In_1046,In_679);
or U101 (N_101,In_1878,In_185);
nor U102 (N_102,In_1761,In_50);
xor U103 (N_103,In_1849,In_398);
xnor U104 (N_104,In_107,In_1745);
xor U105 (N_105,In_479,In_1187);
xor U106 (N_106,In_1883,In_204);
and U107 (N_107,In_1429,In_1830);
xor U108 (N_108,In_1959,In_1587);
and U109 (N_109,In_1272,In_896);
or U110 (N_110,In_1071,In_751);
nand U111 (N_111,In_1487,In_1873);
or U112 (N_112,In_60,In_482);
xor U113 (N_113,In_774,In_1597);
xnor U114 (N_114,In_1253,In_912);
nand U115 (N_115,In_597,In_1447);
nand U116 (N_116,In_1837,In_1631);
xnor U117 (N_117,In_1325,In_371);
xor U118 (N_118,In_474,In_1916);
or U119 (N_119,In_31,In_1358);
nor U120 (N_120,In_1589,In_1546);
nand U121 (N_121,In_1355,In_1296);
and U122 (N_122,In_1995,In_1561);
xnor U123 (N_123,In_619,In_215);
xnor U124 (N_124,In_252,In_1557);
nor U125 (N_125,In_650,In_832);
xnor U126 (N_126,In_2,In_162);
and U127 (N_127,In_560,In_744);
nand U128 (N_128,In_23,In_1766);
or U129 (N_129,In_1966,In_1527);
nand U130 (N_130,In_1424,In_315);
nor U131 (N_131,In_492,In_667);
nand U132 (N_132,In_675,In_265);
nor U133 (N_133,In_502,In_380);
or U134 (N_134,In_759,In_880);
xor U135 (N_135,In_1262,In_1408);
nand U136 (N_136,In_1160,In_1250);
nor U137 (N_137,In_569,In_1102);
and U138 (N_138,In_1339,In_200);
nand U139 (N_139,In_1578,In_777);
nand U140 (N_140,In_392,In_1406);
and U141 (N_141,In_1498,In_1741);
or U142 (N_142,In_286,In_1471);
xnor U143 (N_143,In_1522,In_1600);
nor U144 (N_144,In_225,In_83);
or U145 (N_145,In_127,In_873);
nor U146 (N_146,In_132,In_583);
or U147 (N_147,In_1468,In_1073);
and U148 (N_148,In_797,In_1792);
nand U149 (N_149,In_199,In_1651);
nor U150 (N_150,In_123,In_1904);
or U151 (N_151,In_188,In_768);
xor U152 (N_152,In_955,In_840);
nand U153 (N_153,In_946,In_1202);
xor U154 (N_154,In_1137,In_52);
or U155 (N_155,In_1785,In_1815);
nor U156 (N_156,In_966,In_489);
xnor U157 (N_157,In_1530,In_1679);
nor U158 (N_158,In_0,In_882);
or U159 (N_159,In_584,In_1281);
nor U160 (N_160,In_1094,In_1621);
xor U161 (N_161,In_1955,In_463);
nor U162 (N_162,In_240,In_1299);
and U163 (N_163,In_1421,In_1057);
xor U164 (N_164,In_495,In_1536);
and U165 (N_165,In_670,In_1075);
xor U166 (N_166,In_1362,In_441);
xnor U167 (N_167,In_257,In_1049);
or U168 (N_168,In_1008,In_652);
xnor U169 (N_169,In_1591,In_657);
and U170 (N_170,In_1343,In_376);
or U171 (N_171,In_366,In_1105);
and U172 (N_172,In_626,In_1011);
nand U173 (N_173,In_674,In_1366);
and U174 (N_174,In_86,In_645);
or U175 (N_175,In_293,In_1518);
and U176 (N_176,In_1595,In_369);
or U177 (N_177,In_1588,In_1940);
xor U178 (N_178,In_1855,In_728);
nor U179 (N_179,In_1378,In_1159);
nand U180 (N_180,In_1614,In_27);
xnor U181 (N_181,In_1338,In_112);
xnor U182 (N_182,In_600,In_1107);
and U183 (N_183,In_725,In_1782);
or U184 (N_184,In_277,In_1095);
and U185 (N_185,In_1332,In_808);
xnor U186 (N_186,In_1086,In_430);
xor U187 (N_187,In_1573,In_124);
nand U188 (N_188,In_1714,In_406);
xor U189 (N_189,In_846,In_971);
or U190 (N_190,In_136,In_1946);
and U191 (N_191,In_1979,In_1806);
and U192 (N_192,In_1585,In_1412);
or U193 (N_193,In_6,In_1163);
nor U194 (N_194,In_95,In_1620);
and U195 (N_195,In_1278,In_227);
nand U196 (N_196,In_1865,In_651);
nand U197 (N_197,In_1842,In_1705);
nand U198 (N_198,In_382,In_1393);
or U199 (N_199,In_160,In_636);
or U200 (N_200,In_1742,In_1906);
and U201 (N_201,In_1420,In_1079);
xor U202 (N_202,In_1151,In_524);
nand U203 (N_203,In_76,In_1774);
or U204 (N_204,In_105,In_1549);
or U205 (N_205,In_1122,In_1777);
xnor U206 (N_206,In_1069,In_1520);
and U207 (N_207,In_209,In_874);
xnor U208 (N_208,In_530,In_1570);
nand U209 (N_209,In_1033,In_892);
or U210 (N_210,In_178,In_1941);
nor U211 (N_211,In_247,In_374);
nand U212 (N_212,In_1512,In_824);
xnor U213 (N_213,In_1470,In_1641);
and U214 (N_214,In_196,In_1409);
xnor U215 (N_215,In_688,In_664);
xor U216 (N_216,In_1970,In_919);
nor U217 (N_217,In_1690,In_341);
and U218 (N_218,In_1068,In_828);
nor U219 (N_219,In_542,In_1490);
nor U220 (N_220,In_680,In_1313);
xor U221 (N_221,In_985,In_601);
or U222 (N_222,In_1628,In_311);
or U223 (N_223,In_1133,In_450);
or U224 (N_224,In_1706,In_1182);
and U225 (N_225,In_1427,In_1876);
nand U226 (N_226,In_1604,In_306);
nor U227 (N_227,In_1275,In_411);
nand U228 (N_228,In_272,In_1623);
and U229 (N_229,In_1213,In_454);
nor U230 (N_230,In_1024,In_19);
nor U231 (N_231,In_1067,In_1365);
xor U232 (N_232,In_1880,In_939);
and U233 (N_233,In_219,In_822);
xnor U234 (N_234,In_1466,In_960);
nand U235 (N_235,In_302,In_319);
xnor U236 (N_236,In_948,In_1568);
nor U237 (N_237,In_1882,In_533);
xnor U238 (N_238,In_1045,In_684);
nor U239 (N_239,In_1759,In_891);
nor U240 (N_240,In_662,In_488);
nor U241 (N_241,In_1256,In_238);
and U242 (N_242,In_602,In_703);
or U243 (N_243,In_1270,In_1808);
and U244 (N_244,In_501,In_1973);
nor U245 (N_245,In_363,In_859);
nand U246 (N_246,In_1639,In_1579);
and U247 (N_247,In_1481,In_1884);
nor U248 (N_248,In_468,In_320);
xnor U249 (N_249,In_1968,In_228);
nand U250 (N_250,In_1248,In_1221);
xnor U251 (N_251,In_1287,In_47);
nand U252 (N_252,In_1663,In_1678);
or U253 (N_253,In_1529,In_345);
and U254 (N_254,In_1346,In_504);
nor U255 (N_255,In_1241,In_282);
xor U256 (N_256,In_1435,In_498);
and U257 (N_257,In_494,In_1673);
and U258 (N_258,In_356,In_739);
nor U259 (N_259,In_798,In_1061);
or U260 (N_260,In_1453,In_169);
or U261 (N_261,In_387,In_950);
xnor U262 (N_262,In_1769,In_1610);
nand U263 (N_263,In_661,In_1254);
xor U264 (N_264,In_1999,In_576);
nor U265 (N_265,In_1051,In_935);
nor U266 (N_266,In_1099,In_1727);
and U267 (N_267,In_1169,In_1064);
nand U268 (N_268,In_75,In_1348);
or U269 (N_269,In_1312,In_975);
or U270 (N_270,In_1188,In_1890);
and U271 (N_271,In_548,In_596);
and U272 (N_272,In_1041,In_85);
or U273 (N_273,In_1023,In_696);
or U274 (N_274,In_409,In_544);
nand U275 (N_275,In_1080,In_1027);
and U276 (N_276,In_1164,In_1775);
nand U277 (N_277,In_141,In_1643);
or U278 (N_278,In_1255,In_1709);
nor U279 (N_279,In_237,In_708);
or U280 (N_280,In_244,In_1249);
nand U281 (N_281,In_1634,In_108);
nand U282 (N_282,In_1239,In_729);
nor U283 (N_283,In_710,In_1994);
nor U284 (N_284,In_1874,In_1576);
nor U285 (N_285,In_1243,In_599);
and U286 (N_286,In_1486,In_967);
nand U287 (N_287,In_1392,In_91);
nand U288 (N_288,In_1565,In_806);
xnor U289 (N_289,In_968,In_1893);
or U290 (N_290,In_55,In_1078);
or U291 (N_291,In_159,In_1200);
xnor U292 (N_292,In_243,In_1308);
and U293 (N_293,In_1850,In_285);
nand U294 (N_294,In_1083,In_1060);
xor U295 (N_295,In_1500,In_44);
nand U296 (N_296,In_1238,In_799);
or U297 (N_297,In_368,In_1802);
and U298 (N_298,In_1980,In_695);
nand U299 (N_299,In_522,In_994);
xnor U300 (N_300,In_1509,In_555);
or U301 (N_301,In_1052,In_954);
xor U302 (N_302,In_475,In_1488);
and U303 (N_303,In_713,In_997);
nand U304 (N_304,In_333,In_1629);
and U305 (N_305,In_156,In_1738);
xor U306 (N_306,In_827,In_572);
nor U307 (N_307,In_462,In_590);
nor U308 (N_308,In_1345,In_1801);
nor U309 (N_309,In_1349,In_1625);
nand U310 (N_310,In_1841,In_1538);
and U311 (N_311,In_969,In_1387);
nor U312 (N_312,In_16,In_897);
and U313 (N_313,In_1297,In_1171);
nand U314 (N_314,In_1583,In_1958);
or U315 (N_315,In_1909,In_191);
and U316 (N_316,In_261,In_668);
and U317 (N_317,In_1503,In_1260);
and U318 (N_318,In_217,In_917);
xor U319 (N_319,In_1885,In_523);
nand U320 (N_320,In_271,In_608);
nor U321 (N_321,In_1875,In_1581);
nand U322 (N_322,In_1547,In_1903);
xor U323 (N_323,In_748,In_115);
nand U324 (N_324,In_1938,In_1092);
and U325 (N_325,In_1704,In_1943);
xor U326 (N_326,In_157,In_1445);
and U327 (N_327,In_230,In_940);
or U328 (N_328,In_46,In_1110);
nor U329 (N_329,In_864,In_1524);
nor U330 (N_330,In_268,In_1315);
nor U331 (N_331,In_466,In_1920);
and U332 (N_332,In_1031,In_539);
or U333 (N_333,In_1267,In_587);
and U334 (N_334,In_71,In_1505);
nand U335 (N_335,In_1111,In_151);
or U336 (N_336,In_819,In_1395);
and U337 (N_337,In_1103,In_229);
xor U338 (N_338,In_1337,In_811);
and U339 (N_339,In_1063,In_1988);
xnor U340 (N_340,In_1043,In_578);
nor U341 (N_341,In_113,In_1090);
nor U342 (N_342,In_1832,In_12);
or U343 (N_343,In_1234,In_78);
xnor U344 (N_344,In_1981,In_508);
xor U345 (N_345,In_878,In_672);
and U346 (N_346,In_1795,In_794);
or U347 (N_347,In_352,In_883);
and U348 (N_348,In_427,In_1077);
and U349 (N_349,In_1402,In_1310);
and U350 (N_350,In_1450,In_1716);
xor U351 (N_351,In_1844,In_7);
xnor U352 (N_352,In_1864,In_220);
and U353 (N_353,In_766,In_1448);
or U354 (N_354,In_577,In_1755);
xnor U355 (N_355,In_1054,In_982);
nand U356 (N_356,In_1037,In_1957);
nor U357 (N_357,In_1168,In_1502);
xnor U358 (N_358,In_378,In_1719);
nand U359 (N_359,In_1619,In_182);
and U360 (N_360,In_754,In_732);
or U361 (N_361,In_1953,In_1605);
or U362 (N_362,In_581,In_941);
nand U363 (N_363,In_1177,In_1758);
or U364 (N_364,In_1676,In_1611);
nand U365 (N_365,In_48,In_416);
xor U366 (N_366,In_152,In_1929);
nand U367 (N_367,In_1584,In_646);
and U368 (N_368,In_278,In_771);
xnor U369 (N_369,In_254,In_476);
or U370 (N_370,In_1756,In_556);
or U371 (N_371,In_1781,In_4);
and U372 (N_372,In_336,In_1172);
nor U373 (N_373,In_1788,In_1765);
or U374 (N_374,In_21,In_327);
nand U375 (N_375,In_365,In_1660);
and U376 (N_376,In_1749,In_1464);
nand U377 (N_377,In_213,In_1298);
xor U378 (N_378,In_87,In_149);
and U379 (N_379,In_1590,In_588);
or U380 (N_380,In_1062,In_170);
nor U381 (N_381,In_313,In_924);
nand U382 (N_382,In_142,In_1018);
xnor U383 (N_383,In_1242,In_1135);
and U384 (N_384,In_837,In_1411);
nand U385 (N_385,In_493,In_1125);
nor U386 (N_386,In_1517,In_443);
or U387 (N_387,In_527,In_1131);
or U388 (N_388,In_154,In_849);
nand U389 (N_389,In_1862,In_839);
or U390 (N_390,In_1456,In_89);
and U391 (N_391,In_33,In_726);
and U392 (N_392,In_535,In_623);
and U393 (N_393,In_1457,In_1846);
xor U394 (N_394,In_1065,In_1693);
or U395 (N_395,In_100,In_1971);
nand U396 (N_396,In_516,In_913);
nand U397 (N_397,In_1602,In_594);
nor U398 (N_398,In_825,In_723);
or U399 (N_399,In_915,In_9);
nor U400 (N_400,In_782,In_429);
nand U401 (N_401,In_1148,In_889);
nand U402 (N_402,In_148,N_332);
and U403 (N_403,N_61,N_161);
xnor U404 (N_404,In_1374,In_316);
nor U405 (N_405,In_875,N_388);
xnor U406 (N_406,N_29,In_778);
xor U407 (N_407,In_67,N_212);
or U408 (N_408,In_467,In_1757);
xnor U409 (N_409,In_1661,In_991);
nand U410 (N_410,In_1196,In_1930);
nor U411 (N_411,In_1389,In_41);
or U412 (N_412,N_285,In_1117);
nor U413 (N_413,In_1665,In_995);
or U414 (N_414,N_153,In_925);
nand U415 (N_415,In_370,In_1542);
or U416 (N_416,In_1101,N_235);
and U417 (N_417,In_421,In_1185);
or U418 (N_418,In_1963,N_94);
xnor U419 (N_419,In_1972,In_264);
or U420 (N_420,In_1178,In_472);
nor U421 (N_421,N_274,In_1410);
xor U422 (N_422,N_4,In_559);
and U423 (N_423,In_1934,In_558);
or U424 (N_424,N_65,In_1274);
xor U425 (N_425,In_972,In_1088);
or U426 (N_426,In_99,In_1922);
and U427 (N_427,In_869,In_1089);
and U428 (N_428,In_1367,In_914);
nand U429 (N_429,In_364,In_323);
xnor U430 (N_430,In_757,In_208);
xor U431 (N_431,In_815,N_96);
or U432 (N_432,In_1513,In_1219);
or U433 (N_433,In_1123,In_1768);
or U434 (N_434,N_345,In_762);
and U435 (N_435,In_1917,In_775);
xor U436 (N_436,In_884,In_1269);
nand U437 (N_437,N_352,In_893);
and U438 (N_438,In_129,In_10);
xnor U439 (N_439,In_92,In_988);
nor U440 (N_440,In_1599,In_1961);
and U441 (N_441,In_769,In_1082);
or U442 (N_442,In_1294,N_249);
nor U443 (N_443,In_699,In_28);
or U444 (N_444,In_742,In_1831);
and U445 (N_445,In_1442,In_1982);
xnor U446 (N_446,In_1038,In_270);
and U447 (N_447,In_415,In_1376);
nand U448 (N_448,In_1925,In_362);
nor U449 (N_449,In_246,In_1724);
and U450 (N_450,In_890,In_836);
and U451 (N_451,In_790,N_315);
and U452 (N_452,In_996,N_177);
and U453 (N_453,In_1321,N_142);
nand U454 (N_454,N_256,In_1330);
or U455 (N_455,In_634,In_607);
nor U456 (N_456,In_546,N_99);
nand U457 (N_457,In_177,In_773);
or U458 (N_458,N_181,In_509);
xor U459 (N_459,In_1580,In_871);
nand U460 (N_460,N_183,N_150);
xnor U461 (N_461,In_1544,In_1452);
or U462 (N_462,In_655,N_397);
nor U463 (N_463,In_1829,N_147);
or U464 (N_464,N_133,In_1942);
or U465 (N_465,In_792,N_174);
nor U466 (N_466,In_414,N_382);
xnor U467 (N_467,N_22,N_329);
nand U468 (N_468,N_314,N_32);
or U469 (N_469,In_848,In_1556);
nand U470 (N_470,In_34,N_351);
nor U471 (N_471,In_22,In_258);
or U472 (N_472,N_160,In_1283);
or U473 (N_473,In_1615,In_1462);
and U474 (N_474,In_595,In_350);
xnor U475 (N_475,In_557,N_272);
or U476 (N_476,In_1566,In_776);
xnor U477 (N_477,In_1288,In_1016);
and U478 (N_478,In_1306,In_1649);
xnor U479 (N_479,N_343,In_1762);
xor U480 (N_480,In_163,In_1926);
nor U481 (N_481,In_155,In_563);
and U482 (N_482,N_144,In_1786);
or U483 (N_483,N_36,In_1335);
nor U484 (N_484,In_1819,In_1150);
nor U485 (N_485,N_267,N_44);
or U486 (N_486,N_166,N_126);
or U487 (N_487,In_1199,In_585);
nor U488 (N_488,N_38,In_635);
or U489 (N_489,In_1746,In_1425);
nor U490 (N_490,N_21,In_752);
or U491 (N_491,In_580,In_964);
nor U492 (N_492,N_10,In_1228);
and U493 (N_493,In_1694,In_656);
and U494 (N_494,In_61,In_1702);
and U495 (N_495,N_110,In_1403);
nor U496 (N_496,In_1,N_318);
xor U497 (N_497,In_1685,N_245);
xnor U498 (N_498,In_1292,N_39);
xnor U499 (N_499,N_116,In_1531);
or U500 (N_500,In_1752,In_1737);
xor U501 (N_501,In_1480,In_1005);
xnor U502 (N_502,In_1644,In_420);
nand U503 (N_503,In_1800,N_367);
nor U504 (N_504,In_862,In_1956);
nand U505 (N_505,In_911,In_181);
or U506 (N_506,In_1141,In_334);
nand U507 (N_507,In_709,In_1478);
or U508 (N_508,In_1807,In_317);
or U509 (N_509,In_1637,N_252);
or U510 (N_510,In_483,In_690);
xnor U511 (N_511,N_180,In_1682);
xor U512 (N_512,In_1721,In_1695);
nor U513 (N_513,In_391,N_107);
nand U514 (N_514,In_1495,In_1672);
xnor U515 (N_515,N_326,N_119);
or U516 (N_516,In_1317,N_234);
nand U517 (N_517,In_357,In_1858);
nand U518 (N_518,In_1273,In_1974);
and U519 (N_519,In_404,N_375);
and U520 (N_520,In_622,N_254);
or U521 (N_521,In_1340,In_106);
xnor U522 (N_522,In_360,N_394);
xnor U523 (N_523,In_1303,In_990);
and U524 (N_524,In_1571,In_1108);
nor U525 (N_525,In_1648,In_963);
nand U526 (N_526,In_461,In_45);
and U527 (N_527,In_1139,In_1548);
or U528 (N_528,In_343,In_1120);
nand U529 (N_529,N_233,N_125);
and U530 (N_530,In_1032,N_349);
nor U531 (N_531,In_1494,In_1540);
nand U532 (N_532,N_106,In_1754);
xnor U533 (N_533,In_1118,In_867);
nor U534 (N_534,In_685,In_1838);
and U535 (N_535,In_918,N_275);
nor U536 (N_536,In_283,In_456);
and U537 (N_537,In_428,In_1010);
xnor U538 (N_538,In_457,In_1305);
xnor U539 (N_539,In_300,In_1699);
xnor U540 (N_540,In_54,N_73);
and U541 (N_541,N_227,In_1119);
xor U542 (N_542,N_264,In_961);
or U543 (N_543,In_1871,In_714);
nor U544 (N_544,In_1567,In_1247);
or U545 (N_545,In_738,N_263);
and U546 (N_546,In_1276,In_281);
nor U547 (N_547,In_294,In_66);
and U548 (N_548,In_1908,In_1763);
nand U549 (N_549,In_109,In_484);
and U550 (N_550,In_1251,In_1984);
nand U551 (N_551,N_286,In_1316);
nand U552 (N_552,In_465,In_1231);
nor U553 (N_553,In_1433,In_259);
xnor U554 (N_554,In_1645,In_442);
xnor U555 (N_555,N_373,In_932);
nor U556 (N_556,In_868,In_571);
nand U557 (N_557,In_70,In_1889);
xor U558 (N_558,In_234,N_294);
or U559 (N_559,In_540,In_712);
and U560 (N_560,In_1415,In_1683);
nand U561 (N_561,N_13,In_295);
or U562 (N_562,In_324,N_221);
and U563 (N_563,In_552,In_280);
or U564 (N_564,In_1816,In_1439);
and U565 (N_565,N_386,N_43);
nor U566 (N_566,N_84,N_389);
nand U567 (N_567,N_64,In_1776);
nor U568 (N_568,N_355,N_317);
nor U569 (N_569,In_470,In_1399);
nor U570 (N_570,N_51,In_1047);
nor U571 (N_571,In_444,In_447);
nor U572 (N_572,In_1091,N_209);
xnor U573 (N_573,N_100,In_931);
xnor U574 (N_574,N_82,N_139);
nor U575 (N_575,In_322,In_347);
and U576 (N_576,In_1821,In_1654);
xor U577 (N_577,In_1847,In_613);
and U578 (N_578,In_586,N_269);
and U579 (N_579,In_1905,In_1212);
nor U580 (N_580,In_1861,In_1803);
nand U581 (N_581,N_193,In_1898);
nor U582 (N_582,In_663,In_642);
or U583 (N_583,In_735,In_1224);
nor U584 (N_584,In_84,In_1577);
xnor U585 (N_585,In_861,N_384);
nor U586 (N_586,In_511,In_1000);
and U587 (N_587,In_814,In_1190);
nand U588 (N_588,In_500,In_355);
xnor U589 (N_589,In_1537,N_333);
or U590 (N_590,In_1112,N_134);
nor U591 (N_591,N_101,In_1967);
nor U592 (N_592,N_276,In_536);
xor U593 (N_593,In_1701,N_309);
nor U594 (N_594,In_1007,In_886);
nand U595 (N_595,In_1474,In_144);
nor U596 (N_596,In_553,In_1368);
nor U597 (N_597,In_1783,N_371);
xor U598 (N_598,In_266,N_87);
nor U599 (N_599,In_1461,In_1302);
nand U600 (N_600,In_1382,In_486);
nor U601 (N_601,In_561,N_184);
xor U602 (N_602,In_1469,In_133);
nor U603 (N_603,In_1240,In_1863);
and U604 (N_604,In_14,In_1760);
xnor U605 (N_605,In_1650,N_146);
nor U606 (N_606,N_205,In_1342);
nor U607 (N_607,In_801,N_80);
or U608 (N_608,In_658,N_369);
and U609 (N_609,In_248,N_336);
xnor U610 (N_610,In_385,In_1286);
nand U611 (N_611,In_1021,In_1824);
or U612 (N_612,N_224,In_1939);
nand U613 (N_613,N_208,In_730);
xnor U614 (N_614,In_1827,In_1384);
or U615 (N_615,In_1044,In_1400);
nor U616 (N_616,In_394,N_41);
nand U617 (N_617,In_1662,In_1736);
or U618 (N_618,In_694,In_1508);
nand U619 (N_619,In_682,In_1388);
or U620 (N_620,In_1116,N_232);
nor U621 (N_621,In_137,N_97);
or U622 (N_622,In_1264,N_26);
xnor U623 (N_623,In_1501,In_1372);
nor U624 (N_624,In_1526,In_1545);
nand U625 (N_625,N_25,In_823);
nor U626 (N_626,In_497,In_1770);
or U627 (N_627,N_313,In_1237);
nor U628 (N_628,In_747,In_1271);
or U629 (N_629,N_72,N_176);
and U630 (N_630,In_933,In_1843);
or U631 (N_631,In_1790,N_47);
or U632 (N_632,In_856,In_1076);
xor U633 (N_633,In_1896,N_93);
nor U634 (N_634,In_292,In_168);
and U635 (N_635,In_910,In_953);
nand U636 (N_636,N_364,In_987);
and U637 (N_637,In_852,N_277);
xor U638 (N_638,In_1293,In_617);
xor U639 (N_639,N_159,In_614);
xnor U640 (N_640,In_1473,In_620);
xnor U641 (N_641,In_410,In_32);
or U642 (N_642,In_1352,In_1691);
nor U643 (N_643,In_180,In_120);
and U644 (N_644,In_1205,In_397);
nor U645 (N_645,In_755,In_1978);
and U646 (N_646,In_1066,In_3);
nor U647 (N_647,In_779,In_857);
nand U648 (N_648,In_1050,N_148);
or U649 (N_649,N_88,In_1711);
or U650 (N_650,In_473,In_741);
or U651 (N_651,N_168,N_213);
nor U652 (N_652,In_1295,In_629);
xnor U653 (N_653,In_818,N_165);
xnor U654 (N_654,In_1226,In_1543);
and U655 (N_655,N_145,In_1750);
xnor U656 (N_656,In_1872,In_1586);
and U657 (N_657,In_72,N_300);
nand U658 (N_658,N_280,N_356);
xor U659 (N_659,In_235,In_711);
nor U660 (N_660,In_1035,N_250);
xnor U661 (N_661,In_464,In_1284);
nor U662 (N_662,In_906,In_1475);
xnor U663 (N_663,In_1818,In_787);
and U664 (N_664,In_612,In_1318);
or U665 (N_665,In_885,In_1592);
nand U666 (N_666,In_1124,In_1020);
xor U667 (N_667,In_1437,In_901);
or U668 (N_668,In_1675,N_23);
and U669 (N_669,In_1446,In_1359);
and U670 (N_670,In_565,In_653);
nor U671 (N_671,In_318,In_1477);
nor U672 (N_672,In_611,In_1289);
nand U673 (N_673,N_71,In_1132);
xnor U674 (N_674,N_130,N_74);
nor U675 (N_675,In_1952,In_937);
and U676 (N_676,N_311,In_407);
nor U677 (N_677,N_218,In_448);
or U678 (N_678,N_138,N_378);
or U679 (N_679,In_1176,In_758);
nor U680 (N_680,In_321,In_881);
and U681 (N_681,N_261,In_631);
or U682 (N_682,In_1598,In_800);
nor U683 (N_683,In_93,In_1646);
or U684 (N_684,In_1630,In_1390);
and U685 (N_685,In_745,In_426);
or U686 (N_686,In_399,N_135);
and U687 (N_687,N_358,In_1817);
and U688 (N_688,In_1375,In_1778);
or U689 (N_689,N_298,In_77);
nor U690 (N_690,In_210,In_1230);
nand U691 (N_691,N_340,In_945);
xor U692 (N_692,In_1911,N_225);
nor U693 (N_693,In_677,N_3);
and U694 (N_694,N_1,In_1152);
and U695 (N_695,In_1426,N_290);
and U696 (N_696,In_1423,In_1833);
nor U697 (N_697,In_403,In_666);
and U698 (N_698,In_753,In_1733);
xnor U699 (N_699,In_26,In_290);
or U700 (N_700,In_1991,In_633);
or U701 (N_701,In_1794,In_1364);
or U702 (N_702,In_659,In_134);
or U703 (N_703,In_38,In_505);
nor U704 (N_704,In_289,In_65);
xor U705 (N_705,In_1174,In_1350);
and U706 (N_706,In_1354,In_1902);
xor U707 (N_707,In_175,N_308);
xnor U708 (N_708,N_238,N_127);
and U709 (N_709,In_1812,In_1647);
or U710 (N_710,In_1900,In_1244);
nor U711 (N_711,In_1506,N_237);
or U712 (N_712,In_1493,In_1233);
nor U713 (N_713,In_951,N_360);
and U714 (N_714,In_1324,N_366);
and U715 (N_715,In_1668,N_376);
nor U716 (N_716,In_384,In_1948);
or U717 (N_717,In_1791,N_132);
nand U718 (N_718,In_525,N_310);
nand U719 (N_719,In_926,In_1987);
xnor U720 (N_720,N_344,In_784);
and U721 (N_721,N_391,In_249);
nand U722 (N_722,In_1341,In_1601);
and U723 (N_723,N_78,N_9);
and U724 (N_724,N_170,In_820);
xnor U725 (N_725,In_1158,N_341);
or U726 (N_726,In_379,N_219);
and U727 (N_727,In_1204,In_1640);
nor U728 (N_728,In_1279,In_301);
nand U729 (N_729,In_550,In_589);
nor U730 (N_730,In_959,In_1700);
or U731 (N_731,N_6,In_1371);
xor U732 (N_732,N_103,In_432);
xor U733 (N_733,In_1183,In_1194);
nand U734 (N_734,In_1353,In_487);
nor U735 (N_735,N_327,N_200);
or U736 (N_736,In_1613,N_299);
xnor U737 (N_737,In_1157,In_1499);
xnor U738 (N_738,In_1868,N_350);
nor U739 (N_739,In_1927,In_854);
or U740 (N_740,In_331,In_1671);
xnor U741 (N_741,In_1225,N_291);
nand U742 (N_742,In_1866,In_1729);
nand U743 (N_743,In_396,In_640);
and U744 (N_744,In_510,In_992);
and U745 (N_745,In_1432,In_1401);
nand U746 (N_746,In_838,In_190);
xor U747 (N_747,N_31,In_698);
nand U748 (N_748,In_870,In_1147);
nor U749 (N_749,N_151,In_1377);
and U750 (N_750,In_1162,In_952);
nand U751 (N_751,In_1430,In_1965);
xor U752 (N_752,N_279,In_702);
nand U753 (N_753,In_763,N_204);
and U754 (N_754,In_1206,In_434);
and U755 (N_755,In_1138,In_30);
nand U756 (N_756,In_164,In_843);
xor U757 (N_757,In_260,N_136);
xor U758 (N_758,In_1707,In_1541);
xor U759 (N_759,In_1214,In_1642);
nor U760 (N_760,In_1459,In_593);
nand U761 (N_761,In_1924,N_258);
xnor U762 (N_762,N_175,In_1428);
nand U763 (N_763,In_440,In_851);
nand U764 (N_764,In_224,In_176);
xor U765 (N_765,In_328,N_186);
nand U766 (N_766,In_445,In_807);
nor U767 (N_767,In_103,N_178);
nor U768 (N_768,In_1825,N_57);
or U769 (N_769,N_223,In_1489);
xnor U770 (N_770,N_271,In_789);
nor U771 (N_771,N_48,In_1627);
and U772 (N_772,In_947,N_42);
xor U773 (N_773,In_513,In_207);
nor U774 (N_774,N_342,In_760);
xnor U775 (N_775,In_929,In_1793);
nor U776 (N_776,N_77,In_733);
xnor U777 (N_777,In_1155,N_288);
nor U778 (N_778,N_262,N_283);
or U779 (N_779,In_203,N_24);
or U780 (N_780,In_1810,N_270);
and U781 (N_781,In_1657,In_736);
nor U782 (N_782,N_381,N_15);
xnor U783 (N_783,In_1300,In_833);
nor U784 (N_784,In_812,In_1259);
nor U785 (N_785,N_312,In_805);
nand U786 (N_786,In_346,In_592);
nand U787 (N_787,In_1515,In_62);
xnor U788 (N_788,In_1195,N_244);
or U789 (N_789,N_18,In_24);
or U790 (N_790,In_212,In_795);
and U791 (N_791,In_1042,In_480);
nor U792 (N_792,N_137,In_853);
nor U793 (N_793,N_295,In_1282);
or U794 (N_794,In_110,N_60);
xor U795 (N_795,In_1307,In_150);
xnor U796 (N_796,N_377,N_173);
nor U797 (N_797,In_18,In_1173);
xor U798 (N_798,N_196,In_381);
and U799 (N_799,N_81,N_253);
xnor U800 (N_800,N_420,In_1484);
nor U801 (N_801,In_202,In_1419);
or U802 (N_802,N_30,N_716);
nor U803 (N_803,N_172,N_201);
or U804 (N_804,In_339,In_957);
nand U805 (N_805,N_167,N_687);
or U806 (N_806,In_1839,In_446);
and U807 (N_807,In_1156,In_986);
xor U808 (N_808,In_1684,In_1208);
xor U809 (N_809,In_858,In_1314);
xnor U810 (N_810,N_566,N_169);
nand U811 (N_811,In_1070,In_332);
nor U812 (N_812,N_645,In_1291);
nor U813 (N_813,In_1708,In_737);
and U814 (N_814,In_201,N_659);
xnor U815 (N_815,N_111,N_605);
and U816 (N_816,In_116,In_491);
xor U817 (N_817,In_1804,In_942);
or U818 (N_818,In_727,N_535);
nor U819 (N_819,In_1997,In_1290);
or U820 (N_820,N_383,In_1859);
or U821 (N_821,In_388,N_756);
xor U822 (N_822,N_638,In_564);
nor U823 (N_823,N_556,In_358);
and U824 (N_824,N_502,N_762);
or U825 (N_825,In_1596,N_534);
or U826 (N_826,N_636,N_243);
xnor U827 (N_827,N_574,In_700);
and U828 (N_828,In_905,In_1937);
nand U829 (N_829,N_37,N_675);
and U830 (N_830,In_15,In_1036);
or U831 (N_831,In_273,N_622);
or U832 (N_832,N_484,In_1417);
nand U833 (N_833,In_68,N_567);
or U834 (N_834,N_319,In_1653);
nand U835 (N_835,N_706,In_1796);
xnor U836 (N_836,In_245,In_1483);
and U837 (N_837,In_844,In_143);
nand U838 (N_838,In_1022,In_433);
nor U839 (N_839,In_1492,N_594);
nand U840 (N_840,In_1193,N_790);
and U841 (N_841,In_907,In_88);
xor U842 (N_842,N_668,N_422);
nand U843 (N_843,N_331,N_739);
and U844 (N_844,N_494,N_189);
or U845 (N_845,N_697,N_715);
or U846 (N_846,N_650,N_749);
nor U847 (N_847,N_320,In_1990);
or U848 (N_848,In_984,In_118);
xor U849 (N_849,In_128,In_111);
or U850 (N_850,N_782,N_708);
or U851 (N_851,In_1327,In_1688);
or U852 (N_852,N_129,N_686);
nor U853 (N_853,In_308,In_279);
nand U854 (N_854,N_630,In_1914);
and U855 (N_855,N_602,In_1258);
xnor U856 (N_856,N_152,N_491);
or U857 (N_857,In_1820,N_598);
xor U858 (N_858,In_393,In_36);
xor U859 (N_859,N_575,In_377);
nand U860 (N_860,N_187,In_1894);
nor U861 (N_861,N_287,N_568);
or U862 (N_862,N_455,N_7);
and U863 (N_863,N_55,N_486);
and U864 (N_864,N_581,In_816);
nor U865 (N_865,In_11,In_1369);
and U866 (N_866,N_216,In_1229);
nor U867 (N_867,N_518,In_1006);
nor U868 (N_868,In_1074,N_414);
nor U869 (N_869,N_462,N_619);
xor U870 (N_870,In_1569,N_440);
xnor U871 (N_871,In_1747,N_562);
nand U872 (N_872,N_599,N_433);
and U873 (N_873,In_722,In_977);
and U874 (N_874,N_413,In_520);
or U875 (N_875,N_657,N_418);
or U876 (N_876,In_98,In_1121);
nand U877 (N_877,In_1510,N_485);
nand U878 (N_878,In_1201,N_541);
nor U879 (N_879,In_1235,In_1731);
xnor U880 (N_880,In_1950,In_903);
nor U881 (N_881,In_1441,N_328);
or U882 (N_882,N_467,N_691);
nand U883 (N_883,N_117,In_1463);
and U884 (N_884,In_299,In_829);
nand U885 (N_885,N_334,In_888);
xor U886 (N_886,In_1521,In_1539);
nand U887 (N_887,In_499,N_392);
nor U888 (N_888,In_1454,N_520);
or U889 (N_889,In_970,N_437);
or U890 (N_890,In_1149,In_810);
nand U891 (N_891,N_769,In_974);
nor U892 (N_892,In_654,N_289);
xor U893 (N_893,In_1192,In_1479);
or U894 (N_894,In_610,In_786);
or U895 (N_895,N_563,In_1888);
and U896 (N_896,In_1370,N_778);
nor U897 (N_897,N_236,N_610);
and U898 (N_898,N_661,N_52);
and U899 (N_899,In_222,N_703);
nor U900 (N_900,In_1633,In_507);
and U901 (N_901,N_625,N_307);
nand U902 (N_902,N_601,In_166);
and U903 (N_903,In_1098,In_1947);
and U904 (N_904,In_1422,N_595);
or U905 (N_905,N_463,In_1443);
xnor U906 (N_906,In_1932,In_419);
nor U907 (N_907,In_1867,In_5);
or U908 (N_908,In_743,In_1025);
xor U909 (N_909,N_596,N_717);
and U910 (N_910,N_248,N_785);
and U911 (N_911,N_228,In_877);
or U912 (N_912,N_398,N_191);
nor U913 (N_913,In_697,N_611);
or U914 (N_914,In_459,In_979);
or U915 (N_915,In_389,N_108);
nand U916 (N_916,N_431,In_660);
or U917 (N_917,In_706,N_202);
nor U918 (N_918,N_363,In_1143);
or U919 (N_919,In_314,In_1949);
or U920 (N_920,In_97,N_614);
nand U921 (N_921,In_425,N_514);
xor U922 (N_922,N_663,N_466);
nor U923 (N_923,In_689,N_740);
nor U924 (N_924,In_1528,N_58);
or U925 (N_925,N_63,In_1386);
xnor U926 (N_926,N_546,In_1856);
and U927 (N_927,In_1277,In_1617);
xor U928 (N_928,N_712,N_642);
xnor U929 (N_929,In_750,N_603);
or U930 (N_930,In_671,In_1954);
nor U931 (N_931,In_8,N_629);
nor U932 (N_932,N_488,In_1336);
or U933 (N_933,N_316,In_1280);
nand U934 (N_934,In_1748,In_267);
and U935 (N_935,In_74,N_203);
xor U936 (N_936,In_1680,N_210);
and U937 (N_937,In_402,N_580);
nand U938 (N_938,In_1334,In_767);
nor U939 (N_939,N_772,In_310);
and U940 (N_940,In_785,In_1960);
and U941 (N_941,N_481,In_1309);
nand U942 (N_942,In_949,N_199);
xnor U943 (N_943,N_627,In_1798);
xnor U944 (N_944,In_1805,In_1853);
nor U945 (N_945,N_660,N_572);
xor U946 (N_946,N_164,N_620);
or U947 (N_947,N_695,N_408);
nand U948 (N_948,N_509,N_434);
xnor U949 (N_949,In_1186,N_724);
nor U950 (N_950,In_1560,N_530);
nor U951 (N_951,In_401,In_534);
and U952 (N_952,N_587,In_770);
nor U953 (N_953,In_834,N_729);
nor U954 (N_954,In_1203,N_539);
or U955 (N_955,N_646,N_696);
and U956 (N_956,N_421,In_1167);
nor U957 (N_957,N_643,N_564);
and U958 (N_958,In_981,In_1670);
or U959 (N_959,N_430,In_251);
xor U960 (N_960,In_547,In_1899);
nand U961 (N_961,In_1161,N_616);
nand U962 (N_962,In_1396,N_56);
nor U963 (N_963,In_1356,N_190);
or U964 (N_964,In_354,N_393);
or U965 (N_965,In_1739,In_980);
nand U966 (N_966,In_1983,In_788);
and U967 (N_967,In_847,In_1713);
or U968 (N_968,N_524,In_1053);
xor U969 (N_969,In_195,N_365);
nor U970 (N_970,N_551,In_64);
or U971 (N_971,In_337,N_435);
and U972 (N_972,N_405,N_53);
nand U973 (N_973,In_198,N_34);
nor U974 (N_974,In_554,In_531);
nor U975 (N_975,In_275,In_1319);
xnor U976 (N_976,N_678,N_427);
nor U977 (N_977,N_89,In_1811);
and U978 (N_978,In_183,N_694);
and U979 (N_979,In_418,In_521);
and U980 (N_980,N_33,N_538);
and U981 (N_981,N_733,N_665);
nor U982 (N_982,N_444,N_593);
nor U983 (N_983,N_278,In_351);
or U984 (N_984,N_469,In_673);
nand U985 (N_985,In_1532,In_528);
and U986 (N_986,In_928,In_239);
or U987 (N_987,N_497,N_579);
nor U988 (N_988,N_265,N_69);
or U989 (N_989,In_1127,In_361);
nor U990 (N_990,N_19,In_1535);
xor U991 (N_991,In_104,In_1734);
and U992 (N_992,In_1210,In_221);
or U993 (N_993,N_109,In_503);
xnor U994 (N_994,N_423,N_396);
xnor U995 (N_995,N_465,N_399);
nor U996 (N_996,In_1928,N_20);
xnor U997 (N_997,In_637,In_1227);
nand U998 (N_998,In_1935,In_998);
or U999 (N_999,In_1245,N_492);
or U1000 (N_1000,In_1266,N_516);
nand U1001 (N_1001,N_472,In_63);
nor U1002 (N_1002,N_692,In_1189);
and U1003 (N_1003,In_1087,In_1002);
nand U1004 (N_1004,N_527,In_1834);
nand U1005 (N_1005,In_1511,In_850);
nand U1006 (N_1006,In_615,N_368);
xnor U1007 (N_1007,N_493,In_117);
nor U1008 (N_1008,In_1328,N_11);
xnor U1009 (N_1009,In_73,In_344);
or U1010 (N_1010,N_504,N_2);
and U1011 (N_1011,N_158,In_598);
or U1012 (N_1012,In_373,In_1773);
nor U1013 (N_1013,N_450,N_732);
nand U1014 (N_1014,In_1093,N_255);
nand U1015 (N_1015,N_325,In_1383);
nor U1016 (N_1016,In_647,In_1128);
xor U1017 (N_1017,N_105,In_1222);
nor U1018 (N_1018,N_222,N_512);
or U1019 (N_1019,N_788,In_372);
nand U1020 (N_1020,In_1398,In_335);
and U1021 (N_1021,In_639,In_1551);
or U1022 (N_1022,In_1722,In_342);
or U1023 (N_1023,N_140,N_45);
nor U1024 (N_1024,N_521,In_82);
xnor U1025 (N_1025,In_1301,N_669);
xnor U1026 (N_1026,N_592,In_138);
nor U1027 (N_1027,N_401,N_744);
nor U1028 (N_1028,In_90,N_549);
xnor U1029 (N_1029,N_380,In_1504);
or U1030 (N_1030,N_634,In_1323);
xor U1031 (N_1031,In_543,N_330);
and U1032 (N_1032,In_1618,N_505);
nand U1033 (N_1033,In_551,In_455);
nor U1034 (N_1034,N_640,In_1636);
and U1035 (N_1035,In_451,N_452);
and U1036 (N_1036,In_140,In_284);
nor U1037 (N_1037,In_469,N_540);
nor U1038 (N_1038,In_274,N_303);
nand U1039 (N_1039,In_174,N_429);
and U1040 (N_1040,In_1977,In_1351);
nor U1041 (N_1041,N_722,In_916);
xor U1042 (N_1042,In_570,N_447);
xnor U1043 (N_1043,N_454,N_390);
xor U1044 (N_1044,N_428,N_475);
or U1045 (N_1045,N_537,In_549);
nand U1046 (N_1046,N_682,In_1320);
nor U1047 (N_1047,In_1363,In_976);
xnor U1048 (N_1048,N_424,N_557);
nor U1049 (N_1049,In_973,N_171);
and U1050 (N_1050,N_730,N_789);
xnor U1051 (N_1051,N_552,N_515);
xor U1052 (N_1052,In_676,N_768);
or U1053 (N_1053,In_153,In_1612);
nor U1054 (N_1054,N_719,In_1013);
or U1055 (N_1055,In_1743,N_115);
nand U1056 (N_1056,N_500,In_1019);
nand U1057 (N_1057,In_325,N_647);
or U1058 (N_1058,In_253,In_1969);
nor U1059 (N_1059,In_490,In_167);
nor U1060 (N_1060,N_12,In_921);
xnor U1061 (N_1061,N_720,N_482);
nand U1062 (N_1062,In_218,N_305);
nor U1063 (N_1063,In_1656,N_128);
xor U1064 (N_1064,In_1563,N_155);
and U1065 (N_1065,In_993,In_288);
nor U1066 (N_1066,In_1431,N_583);
xnor U1067 (N_1067,N_584,In_1593);
nor U1068 (N_1068,In_644,N_306);
xnor U1069 (N_1069,N_569,In_1607);
nand U1070 (N_1070,In_96,In_184);
or U1071 (N_1071,N_461,N_302);
nor U1072 (N_1072,N_76,In_1407);
nor U1073 (N_1073,In_865,N_704);
nand U1074 (N_1074,In_1017,In_1918);
xnor U1075 (N_1075,N_501,N_419);
xnor U1076 (N_1076,N_489,N_644);
nand U1077 (N_1077,N_617,In_1897);
nor U1078 (N_1078,In_303,In_1712);
or U1079 (N_1079,In_1246,In_830);
nor U1080 (N_1080,N_761,In_1718);
nor U1081 (N_1081,In_400,In_1854);
nor U1082 (N_1082,N_671,N_652);
nor U1083 (N_1083,In_1418,In_1687);
or U1084 (N_1084,N_215,N_259);
nor U1085 (N_1085,In_1444,N_728);
and U1086 (N_1086,In_965,N_618);
nand U1087 (N_1087,N_738,N_532);
or U1088 (N_1088,N_693,N_195);
nand U1089 (N_1089,In_1666,N_543);
or U1090 (N_1090,In_197,N_755);
nor U1091 (N_1091,N_585,In_1698);
nand U1092 (N_1092,In_43,N_759);
and U1093 (N_1093,N_590,In_1740);
nor U1094 (N_1094,N_400,N_672);
nand U1095 (N_1095,N_667,N_359);
and U1096 (N_1096,N_448,N_623);
or U1097 (N_1097,In_1554,In_1575);
xnor U1098 (N_1098,In_1344,N_66);
xnor U1099 (N_1099,N_586,N_774);
nand U1100 (N_1100,N_185,In_538);
or U1101 (N_1101,N_754,N_457);
or U1102 (N_1102,N_550,N_241);
and U1103 (N_1103,N_214,In_909);
nand U1104 (N_1104,In_1594,In_1681);
or U1105 (N_1105,In_1482,N_685);
nor U1106 (N_1106,N_104,In_1385);
nor U1107 (N_1107,N_102,In_900);
nor U1108 (N_1108,N_680,In_1449);
and U1109 (N_1109,In_1534,N_416);
and U1110 (N_1110,In_606,N_773);
and U1111 (N_1111,N_179,In_1485);
nor U1112 (N_1112,N_597,N_470);
nor U1113 (N_1113,N_323,In_1848);
nor U1114 (N_1114,N_395,In_518);
and U1115 (N_1115,In_678,N_783);
nand U1116 (N_1116,In_119,N_75);
or U1117 (N_1117,N_217,In_1331);
xnor U1118 (N_1118,N_736,In_193);
and U1119 (N_1119,In_1126,N_439);
nand U1120 (N_1120,N_27,N_626);
xnor U1121 (N_1121,N_91,N_677);
xnor U1122 (N_1122,In_791,N_483);
xnor U1123 (N_1123,N_559,N_528);
xnor U1124 (N_1124,In_1609,In_1826);
and U1125 (N_1125,N_468,In_1550);
nand U1126 (N_1126,N_348,In_431);
xor U1127 (N_1127,In_1215,In_804);
nand U1128 (N_1128,In_938,N_674);
nor U1129 (N_1129,In_1153,N_745);
xor U1130 (N_1130,In_1434,In_1472);
or U1131 (N_1131,In_1012,N_449);
nor U1132 (N_1132,N_379,N_231);
nand U1133 (N_1133,In_1373,In_1852);
xor U1134 (N_1134,N_709,N_487);
and U1135 (N_1135,N_517,In_173);
nand U1136 (N_1136,In_263,In_59);
nor U1137 (N_1137,N_510,N_711);
nand U1138 (N_1138,N_544,N_673);
and U1139 (N_1139,N_339,In_1211);
and U1140 (N_1140,N_304,N_409);
nor U1141 (N_1141,N_632,In_304);
or U1142 (N_1142,In_962,N_781);
and U1143 (N_1143,In_423,N_16);
and U1144 (N_1144,In_1507,N_743);
and U1145 (N_1145,N_40,N_473);
and U1146 (N_1146,In_1029,N_471);
and U1147 (N_1147,In_517,In_20);
or U1148 (N_1148,In_1451,N_479);
or U1149 (N_1149,In_1677,N_321);
xnor U1150 (N_1150,In_1465,In_1753);
nand U1151 (N_1151,N_426,N_425);
nor U1152 (N_1152,N_666,N_796);
xnor U1153 (N_1153,N_456,N_731);
and U1154 (N_1154,N_545,N_609);
and U1155 (N_1155,In_383,N_725);
and U1156 (N_1156,N_681,In_1696);
xor U1157 (N_1157,N_795,In_1901);
nor U1158 (N_1158,N_404,N_67);
nor U1159 (N_1159,N_784,N_742);
xor U1160 (N_1160,In_453,N_770);
nor U1161 (N_1161,N_372,N_760);
nor U1162 (N_1162,N_297,N_411);
nand U1163 (N_1163,N_727,N_588);
and U1164 (N_1164,In_989,In_1440);
or U1165 (N_1165,N_600,In_1814);
nand U1166 (N_1166,N_387,In_1114);
and U1167 (N_1167,In_471,N_50);
or U1168 (N_1168,In_1993,N_741);
and U1169 (N_1169,In_1130,In_624);
nand U1170 (N_1170,N_747,N_143);
or U1171 (N_1171,In_809,N_591);
nand U1172 (N_1172,N_460,In_630);
nor U1173 (N_1173,In_1603,N_542);
nand U1174 (N_1174,In_179,N_641);
and U1175 (N_1175,N_794,N_679);
nor U1176 (N_1176,N_120,N_558);
and U1177 (N_1177,N_123,In_1931);
and U1178 (N_1178,In_920,N_451);
or U1179 (N_1179,N_604,N_792);
nand U1180 (N_1180,In_1870,In_1001);
nand U1181 (N_1181,N_737,In_1058);
nand U1182 (N_1182,N_220,N_8);
and U1183 (N_1183,N_266,In_1608);
and U1184 (N_1184,In_705,N_664);
and U1185 (N_1185,In_566,In_930);
xor U1186 (N_1186,N_257,In_842);
or U1187 (N_1187,N_357,N_702);
nor U1188 (N_1188,In_171,N_633);
or U1189 (N_1189,N_607,N_251);
and U1190 (N_1190,N_141,N_734);
nor U1191 (N_1191,In_53,N_296);
or U1192 (N_1192,In_1996,N_529);
nand U1193 (N_1193,N_284,N_337);
nand U1194 (N_1194,In_1191,In_526);
xor U1195 (N_1195,N_506,In_1198);
nor U1196 (N_1196,N_656,N_779);
or U1197 (N_1197,N_608,In_422);
or U1198 (N_1198,In_821,N_648);
nand U1199 (N_1199,N_459,N_85);
and U1200 (N_1200,N_1015,N_746);
and U1201 (N_1201,N_1162,In_125);
nand U1202 (N_1202,In_1207,N_121);
nor U1203 (N_1203,N_944,In_1106);
xnor U1204 (N_1204,N_1072,In_562);
or U1205 (N_1205,N_873,In_1154);
xnor U1206 (N_1206,N_301,N_282);
nor U1207 (N_1207,N_118,N_1177);
nand U1208 (N_1208,N_1031,N_927);
and U1209 (N_1209,N_1181,In_802);
and U1210 (N_1210,N_1057,N_908);
or U1211 (N_1211,N_1078,N_1000);
xnor U1212 (N_1212,N_163,N_939);
and U1213 (N_1213,N_982,N_157);
xnor U1214 (N_1214,N_1139,N_887);
xor U1215 (N_1215,N_1130,N_1083);
or U1216 (N_1216,N_1192,N_960);
nand U1217 (N_1217,N_941,N_480);
xor U1218 (N_1218,N_936,N_1086);
and U1219 (N_1219,N_1146,N_1186);
nand U1220 (N_1220,N_577,N_840);
and U1221 (N_1221,N_923,N_893);
and U1222 (N_1222,In_330,N_1178);
xnor U1223 (N_1223,N_1063,N_834);
nor U1224 (N_1224,In_242,N_854);
nand U1225 (N_1225,N_1007,N_753);
nand U1226 (N_1226,In_1458,N_62);
or U1227 (N_1227,N_816,N_942);
xnor U1228 (N_1228,N_635,N_182);
nor U1229 (N_1229,N_1096,N_777);
xor U1230 (N_1230,N_1009,N_714);
and U1231 (N_1231,N_1075,N_1138);
or U1232 (N_1232,N_293,N_1107);
or U1233 (N_1233,In_1869,N_751);
and U1234 (N_1234,N_862,N_606);
and U1235 (N_1235,In_135,N_1058);
nor U1236 (N_1236,N_1189,N_1050);
xor U1237 (N_1237,In_1616,In_541);
nand U1238 (N_1238,In_17,In_1285);
xnor U1239 (N_1239,N_670,N_848);
nand U1240 (N_1240,N_819,N_1169);
or U1241 (N_1241,In_927,N_833);
xnor U1242 (N_1242,N_1128,In_902);
xnor U1243 (N_1243,N_943,N_843);
nor U1244 (N_1244,In_386,In_51);
and U1245 (N_1245,N_857,In_307);
xor U1246 (N_1246,N_1191,N_490);
and U1247 (N_1247,N_1092,N_90);
xnor U1248 (N_1248,N_850,N_273);
and U1249 (N_1249,N_1125,N_835);
nand U1250 (N_1250,N_969,N_830);
and U1251 (N_1251,In_1218,N_949);
and U1252 (N_1252,N_820,N_86);
nand U1253 (N_1253,N_1098,N_1028);
nand U1254 (N_1254,In_716,N_1190);
nor U1255 (N_1255,N_844,In_58);
and U1256 (N_1256,N_932,In_256);
nor U1257 (N_1257,In_390,In_1039);
nand U1258 (N_1258,In_983,N_1155);
nor U1259 (N_1259,N_1019,In_649);
nor U1260 (N_1260,In_1771,N_1095);
and U1261 (N_1261,In_1717,N_748);
xnor U1262 (N_1262,N_547,N_1116);
and U1263 (N_1263,N_976,In_1220);
xnor U1264 (N_1264,In_605,N_870);
and U1265 (N_1265,N_1118,N_247);
nor U1266 (N_1266,In_1962,N_821);
or U1267 (N_1267,N_1187,In_1175);
nand U1268 (N_1268,N_825,N_1018);
nor U1269 (N_1269,N_1064,N_507);
xnor U1270 (N_1270,N_68,N_441);
nand U1271 (N_1271,N_881,N_533);
nand U1272 (N_1272,N_767,N_0);
or U1273 (N_1273,N_683,In_233);
xor U1274 (N_1274,In_147,N_324);
or U1275 (N_1275,N_1011,N_735);
or U1276 (N_1276,In_114,N_947);
and U1277 (N_1277,N_860,N_855);
nor U1278 (N_1278,In_999,In_1789);
or U1279 (N_1279,N_1194,N_1151);
or U1280 (N_1280,N_1029,In_1964);
xnor U1281 (N_1281,N_1049,N_897);
xnor U1282 (N_1282,In_49,N_987);
and U1283 (N_1283,N_14,N_957);
nor U1284 (N_1284,In_793,N_757);
nand U1285 (N_1285,N_1126,N_953);
xnor U1286 (N_1286,In_56,In_438);
nor U1287 (N_1287,N_554,N_1102);
nand U1288 (N_1288,In_609,N_917);
and U1289 (N_1289,N_827,N_883);
nand U1290 (N_1290,N_1154,N_994);
or U1291 (N_1291,In_1170,In_1992);
xnor U1292 (N_1292,N_1068,N_1005);
and U1293 (N_1293,In_413,In_575);
xnor U1294 (N_1294,N_1048,N_1043);
or U1295 (N_1295,In_146,In_898);
xnor U1296 (N_1296,N_710,N_335);
xnor U1297 (N_1297,N_1120,In_519);
or U1298 (N_1298,N_197,N_1183);
or U1299 (N_1299,N_1145,N_1073);
or U1300 (N_1300,N_1110,In_435);
or U1301 (N_1301,N_445,In_121);
xor U1302 (N_1302,N_1091,N_1088);
and U1303 (N_1303,In_582,N_752);
nor U1304 (N_1304,N_845,In_1115);
or U1305 (N_1305,N_412,N_1106);
and U1306 (N_1306,In_122,N_194);
and U1307 (N_1307,N_713,N_322);
or U1308 (N_1308,In_94,N_904);
and U1309 (N_1309,N_1180,N_851);
xnor U1310 (N_1310,N_1079,N_1143);
nand U1311 (N_1311,N_1193,N_684);
or U1312 (N_1312,In_1933,N_292);
or U1313 (N_1313,N_839,N_1195);
or U1314 (N_1314,N_1042,N_1127);
or U1315 (N_1315,In_338,N_1117);
nand U1316 (N_1316,N_1158,N_999);
nor U1317 (N_1317,In_79,N_879);
or U1318 (N_1318,N_763,N_112);
xor U1319 (N_1319,N_1023,In_375);
nor U1320 (N_1320,N_1173,N_5);
or U1321 (N_1321,N_511,N_407);
nor U1322 (N_1322,In_1881,In_866);
xor U1323 (N_1323,In_579,N_1069);
xor U1324 (N_1324,In_1034,In_349);
nand U1325 (N_1325,In_1197,In_326);
and U1326 (N_1326,In_1209,N_866);
or U1327 (N_1327,N_347,N_526);
xor U1328 (N_1328,N_1131,In_1632);
or U1329 (N_1329,In_532,N_79);
or U1330 (N_1330,N_959,N_226);
and U1331 (N_1331,N_900,N_938);
nand U1332 (N_1332,N_912,In_1552);
and U1333 (N_1333,N_829,In_1497);
nor U1334 (N_1334,N_899,In_194);
and U1335 (N_1335,N_1123,N_156);
xnor U1336 (N_1336,N_565,N_971);
xnor U1337 (N_1337,N_1199,N_1051);
nand U1338 (N_1338,N_867,N_1089);
nand U1339 (N_1339,N_980,In_545);
nand U1340 (N_1340,N_817,In_1986);
xnor U1341 (N_1341,In_904,N_974);
and U1342 (N_1342,N_909,In_101);
xnor U1343 (N_1343,N_436,N_346);
or U1344 (N_1344,N_1164,N_446);
or U1345 (N_1345,N_898,In_1669);
nor U1346 (N_1346,N_992,N_998);
nor U1347 (N_1347,N_246,N_924);
nand U1348 (N_1348,N_1001,N_1046);
nand U1349 (N_1349,In_206,N_1080);
and U1350 (N_1350,N_496,N_750);
nand U1351 (N_1351,N_838,In_1268);
nor U1352 (N_1352,N_1124,N_919);
nand U1353 (N_1353,N_499,In_460);
xor U1354 (N_1354,N_955,In_887);
xor U1355 (N_1355,N_807,N_824);
xnor U1356 (N_1356,N_442,N_403);
nand U1357 (N_1357,N_361,N_991);
xor U1358 (N_1358,In_715,N_229);
nand U1359 (N_1359,N_1006,In_701);
and U1360 (N_1360,N_951,N_122);
nor U1361 (N_1361,N_805,N_1185);
xor U1362 (N_1362,N_869,In_481);
or U1363 (N_1363,In_81,In_1496);
xnor U1364 (N_1364,In_412,N_918);
or U1365 (N_1365,N_1122,N_966);
xor U1366 (N_1366,N_458,N_874);
and U1367 (N_1367,N_811,N_410);
or U1368 (N_1368,N_649,N_766);
and U1369 (N_1369,N_802,In_1635);
nor U1370 (N_1370,N_415,N_950);
or U1371 (N_1371,N_1133,N_1174);
and U1372 (N_1372,N_1025,N_891);
nor U1373 (N_1373,N_1012,N_793);
and U1374 (N_1374,In_1360,N_192);
or U1375 (N_1375,N_1157,N_986);
or U1376 (N_1376,N_814,N_965);
nor U1377 (N_1377,N_718,N_878);
nand U1378 (N_1378,N_1170,In_1726);
xnor U1379 (N_1379,N_1103,N_1165);
or U1380 (N_1380,N_990,N_374);
and U1381 (N_1381,N_1197,In_1333);
and U1382 (N_1382,N_836,N_1160);
nor U1383 (N_1383,N_1032,N_70);
nor U1384 (N_1384,N_1188,N_997);
or U1385 (N_1385,In_1887,N_49);
nor U1386 (N_1386,N_613,N_1036);
nor U1387 (N_1387,N_1059,N_954);
nand U1388 (N_1388,N_863,N_35);
nor U1389 (N_1389,N_653,In_1667);
and U1390 (N_1390,N_615,In_39);
xnor U1391 (N_1391,N_1097,N_498);
and U1392 (N_1392,N_1040,In_1165);
and U1393 (N_1393,N_1137,N_676);
nor U1394 (N_1394,In_761,N_628);
or U1395 (N_1395,In_692,N_786);
or U1396 (N_1396,N_1112,N_1087);
and U1397 (N_1397,N_662,In_1072);
and U1398 (N_1398,N_1047,N_1175);
or U1399 (N_1399,In_1180,N_1141);
xnor U1400 (N_1400,N_922,N_871);
nand U1401 (N_1401,N_1115,N_892);
nand U1402 (N_1402,In_1985,In_707);
nand U1403 (N_1403,In_329,In_57);
xor U1404 (N_1404,N_1152,N_859);
and U1405 (N_1405,N_1172,N_826);
nand U1406 (N_1406,N_385,N_1027);
xnor U1407 (N_1407,In_765,N_903);
nor U1408 (N_1408,N_1037,In_746);
and U1409 (N_1409,N_765,N_995);
and U1410 (N_1410,N_1082,N_525);
or U1411 (N_1411,N_578,In_512);
xnor U1412 (N_1412,N_495,In_1014);
xnor U1413 (N_1413,N_230,In_1919);
and U1414 (N_1414,N_443,In_855);
nor U1415 (N_1415,N_890,N_813);
and U1416 (N_1416,In_764,N_905);
nand U1417 (N_1417,N_868,N_721);
or U1418 (N_1418,N_929,N_952);
or U1419 (N_1419,N_797,N_281);
xor U1420 (N_1420,N_1034,N_846);
nor U1421 (N_1421,N_370,N_700);
nor U1422 (N_1422,N_937,N_1026);
nand U1423 (N_1423,In_665,N_1142);
or U1424 (N_1424,N_979,N_1176);
and U1425 (N_1425,N_989,N_690);
or U1426 (N_1426,N_1074,N_885);
nand U1427 (N_1427,In_1217,N_988);
or U1428 (N_1428,In_13,N_1093);
xnor U1429 (N_1429,N_985,N_453);
xnor U1430 (N_1430,N_149,N_1168);
nor U1431 (N_1431,N_570,In_537);
or U1432 (N_1432,N_612,In_1136);
nand U1433 (N_1433,N_895,In_1944);
xnor U1434 (N_1434,N_1144,In_269);
or U1435 (N_1435,N_967,N_726);
nor U1436 (N_1436,N_1184,N_925);
nand U1437 (N_1437,N_1010,N_916);
nor U1438 (N_1438,N_1140,In_1553);
nor U1439 (N_1439,N_972,N_798);
xor U1440 (N_1440,N_961,N_1022);
nor U1441 (N_1441,N_1070,In_1764);
and U1442 (N_1442,In_1823,N_474);
and U1443 (N_1443,N_1148,N_639);
nor U1444 (N_1444,N_476,N_1163);
or U1445 (N_1445,In_1438,N_1114);
nand U1446 (N_1446,N_1038,N_915);
nor U1447 (N_1447,In_831,N_1013);
nor U1448 (N_1448,N_1071,N_806);
nor U1449 (N_1449,N_1159,N_865);
xor U1450 (N_1450,N_791,N_1135);
nand U1451 (N_1451,N_242,N_92);
nand U1452 (N_1452,N_338,N_884);
nor U1453 (N_1453,N_1109,N_114);
xor U1454 (N_1454,In_1744,N_975);
and U1455 (N_1455,N_131,In_1913);
and U1456 (N_1456,In_895,N_926);
nand U1457 (N_1457,N_1101,N_856);
nand U1458 (N_1458,N_621,In_1476);
and U1459 (N_1459,N_933,In_783);
xor U1460 (N_1460,N_582,N_17);
and U1461 (N_1461,N_818,N_503);
xor U1462 (N_1462,N_508,N_1066);
nand U1463 (N_1463,In_211,N_1044);
or U1464 (N_1464,N_432,In_1381);
nor U1465 (N_1465,In_1311,In_1525);
nor U1466 (N_1466,In_616,N_651);
nor U1467 (N_1467,In_1659,In_1840);
nor U1468 (N_1468,In_1912,N_699);
xnor U1469 (N_1469,N_1105,N_852);
and U1470 (N_1470,N_1052,In_1056);
nand U1471 (N_1471,N_1108,N_832);
nor U1472 (N_1472,N_438,In_1104);
xor U1473 (N_1473,In_1835,In_296);
nand U1474 (N_1474,In_1998,N_211);
and U1475 (N_1475,In_603,N_1053);
or U1476 (N_1476,N_809,N_808);
xor U1477 (N_1477,N_1014,N_519);
nand U1478 (N_1478,N_1084,In_477);
nand U1479 (N_1479,In_1828,N_901);
nand U1480 (N_1480,In_529,N_701);
and U1481 (N_1481,N_902,In_189);
nor U1482 (N_1482,N_98,In_860);
or U1483 (N_1483,N_658,In_165);
and U1484 (N_1484,N_984,In_1877);
xnor U1485 (N_1485,In_641,N_935);
nand U1486 (N_1486,N_95,N_560);
or U1487 (N_1487,N_631,N_354);
and U1488 (N_1488,In_573,N_1017);
and U1489 (N_1489,In_721,N_803);
nor U1490 (N_1490,In_1989,N_406);
and U1491 (N_1491,N_1004,In_719);
nand U1492 (N_1492,N_771,N_1166);
or U1493 (N_1493,In_1097,In_686);
or U1494 (N_1494,N_1198,N_841);
xnor U1495 (N_1495,In_1689,N_931);
nand U1496 (N_1496,In_568,N_1067);
and U1497 (N_1497,N_815,N_973);
nor U1498 (N_1498,In_796,N_1196);
nor U1499 (N_1499,N_548,N_571);
nor U1500 (N_1500,In_69,In_772);
and U1501 (N_1501,N_402,N_698);
xor U1502 (N_1502,N_847,N_523);
and U1503 (N_1503,N_822,N_764);
nand U1504 (N_1504,N_799,N_637);
and U1505 (N_1505,N_1021,In_1394);
nand U1506 (N_1506,N_896,N_894);
xnor U1507 (N_1507,In_1558,N_983);
nand U1508 (N_1508,N_1156,N_46);
and U1509 (N_1509,N_1171,N_758);
or U1510 (N_1510,N_707,N_1045);
and U1511 (N_1511,N_522,N_787);
and U1512 (N_1512,N_776,N_207);
or U1513 (N_1513,In_1015,N_1119);
nand U1514 (N_1514,In_223,N_1003);
xnor U1515 (N_1515,In_1232,In_756);
and U1516 (N_1516,In_683,N_1076);
and U1517 (N_1517,N_968,In_348);
nand U1518 (N_1518,N_536,N_842);
xnor U1519 (N_1519,In_1304,N_1085);
nand U1520 (N_1520,N_1147,N_858);
nand U1521 (N_1521,N_907,N_59);
nor U1522 (N_1522,N_801,N_478);
nand U1523 (N_1523,N_28,N_1056);
xnor U1524 (N_1524,N_240,In_826);
xor U1525 (N_1525,In_1921,N_124);
xnor U1526 (N_1526,N_555,In_1361);
nor U1527 (N_1527,N_1062,N_1065);
or U1528 (N_1528,In_574,N_464);
nand U1529 (N_1529,N_849,N_268);
xnor U1530 (N_1530,In_478,N_1182);
xor U1531 (N_1531,N_906,N_940);
or U1532 (N_1532,N_83,N_958);
and U1533 (N_1533,In_1109,N_723);
nor U1534 (N_1534,N_1132,N_688);
and U1535 (N_1535,N_239,In_1664);
and U1536 (N_1536,In_1787,N_877);
or U1537 (N_1537,N_1008,In_1030);
or U1538 (N_1538,N_861,N_54);
nand U1539 (N_1539,In_1263,N_1179);
nor U1540 (N_1540,In_1606,N_928);
nand U1541 (N_1541,N_188,N_996);
and U1542 (N_1542,N_705,N_800);
nand U1543 (N_1543,In_1799,N_780);
nor U1544 (N_1544,N_1041,In_718);
xor U1545 (N_1545,N_880,N_823);
nand U1546 (N_1546,N_1121,N_876);
nor U1547 (N_1547,In_1026,N_353);
xor U1548 (N_1548,N_553,N_1100);
xor U1549 (N_1549,N_993,In_1514);
xnor U1550 (N_1550,In_35,In_1179);
nand U1551 (N_1551,N_962,N_804);
and U1552 (N_1552,In_978,N_1111);
or U1553 (N_1553,N_775,N_970);
nand U1554 (N_1554,In_161,N_978);
or U1555 (N_1555,N_886,N_1090);
nand U1556 (N_1556,N_964,N_1054);
nand U1557 (N_1557,N_1002,N_946);
or U1558 (N_1558,N_477,In_439);
and U1559 (N_1559,N_154,N_1033);
or U1560 (N_1560,N_362,In_943);
nor U1561 (N_1561,In_139,N_1039);
and U1562 (N_1562,N_1099,N_573);
and U1563 (N_1563,N_977,N_934);
and U1564 (N_1564,N_1129,N_1150);
and U1565 (N_1565,N_828,N_206);
xnor U1566 (N_1566,N_1134,N_589);
nand U1567 (N_1567,N_981,N_910);
nor U1568 (N_1568,N_1136,In_214);
nand U1569 (N_1569,N_654,N_1020);
or U1570 (N_1570,N_913,N_875);
or U1571 (N_1571,In_1574,N_914);
nand U1572 (N_1572,N_1077,N_689);
and U1573 (N_1573,N_831,In_780);
and U1574 (N_1574,N_513,N_911);
xnor U1575 (N_1575,N_655,In_1892);
or U1576 (N_1576,N_888,In_648);
xnor U1577 (N_1577,N_417,N_260);
or U1578 (N_1578,N_853,N_920);
xnor U1579 (N_1579,N_1149,N_930);
nand U1580 (N_1580,In_172,N_837);
nor U1581 (N_1581,N_956,N_561);
nand U1582 (N_1582,In_1860,N_1024);
nand U1583 (N_1583,N_624,N_531);
nand U1584 (N_1584,N_1113,N_1094);
nor U1585 (N_1585,N_963,N_1153);
xor U1586 (N_1586,N_162,N_1055);
nand U1587 (N_1587,N_1030,N_872);
and U1588 (N_1588,N_921,In_1780);
nor U1589 (N_1589,N_882,N_113);
nor U1590 (N_1590,N_1167,N_1161);
and U1591 (N_1591,In_879,N_576);
xnor U1592 (N_1592,In_1404,N_1081);
xnor U1593 (N_1593,N_948,N_889);
and U1594 (N_1594,N_1104,In_291);
and U1595 (N_1595,N_864,N_810);
nand U1596 (N_1596,N_198,N_1035);
or U1597 (N_1597,In_1720,N_1016);
or U1598 (N_1598,N_945,N_812);
or U1599 (N_1599,N_1061,N_1060);
and U1600 (N_1600,N_1405,N_1531);
and U1601 (N_1601,N_1249,N_1539);
or U1602 (N_1602,N_1592,N_1217);
nand U1603 (N_1603,N_1513,N_1346);
and U1604 (N_1604,N_1447,N_1481);
or U1605 (N_1605,N_1548,N_1480);
or U1606 (N_1606,N_1272,N_1216);
xor U1607 (N_1607,N_1428,N_1468);
or U1608 (N_1608,N_1223,N_1577);
nand U1609 (N_1609,N_1341,N_1459);
nand U1610 (N_1610,N_1330,N_1427);
nand U1611 (N_1611,N_1415,N_1448);
and U1612 (N_1612,N_1358,N_1474);
and U1613 (N_1613,N_1209,N_1324);
nor U1614 (N_1614,N_1311,N_1434);
nand U1615 (N_1615,N_1425,N_1560);
or U1616 (N_1616,N_1570,N_1335);
or U1617 (N_1617,N_1452,N_1408);
nand U1618 (N_1618,N_1483,N_1536);
or U1619 (N_1619,N_1544,N_1521);
nand U1620 (N_1620,N_1527,N_1348);
or U1621 (N_1621,N_1492,N_1437);
nand U1622 (N_1622,N_1368,N_1477);
xnor U1623 (N_1623,N_1522,N_1310);
and U1624 (N_1624,N_1239,N_1430);
nand U1625 (N_1625,N_1424,N_1248);
xnor U1626 (N_1626,N_1562,N_1420);
xnor U1627 (N_1627,N_1479,N_1302);
or U1628 (N_1628,N_1457,N_1396);
xor U1629 (N_1629,N_1213,N_1581);
nand U1630 (N_1630,N_1529,N_1506);
or U1631 (N_1631,N_1391,N_1332);
nand U1632 (N_1632,N_1493,N_1557);
or U1633 (N_1633,N_1262,N_1319);
and U1634 (N_1634,N_1289,N_1345);
xnor U1635 (N_1635,N_1431,N_1490);
nor U1636 (N_1636,N_1453,N_1378);
xor U1637 (N_1637,N_1300,N_1407);
xnor U1638 (N_1638,N_1467,N_1259);
nor U1639 (N_1639,N_1224,N_1393);
nand U1640 (N_1640,N_1422,N_1261);
or U1641 (N_1641,N_1251,N_1443);
xor U1642 (N_1642,N_1372,N_1244);
and U1643 (N_1643,N_1387,N_1250);
xnor U1644 (N_1644,N_1455,N_1450);
xnor U1645 (N_1645,N_1414,N_1571);
nand U1646 (N_1646,N_1350,N_1576);
nor U1647 (N_1647,N_1351,N_1280);
xor U1648 (N_1648,N_1207,N_1556);
nor U1649 (N_1649,N_1215,N_1287);
nand U1650 (N_1650,N_1419,N_1542);
and U1651 (N_1651,N_1361,N_1456);
nor U1652 (N_1652,N_1336,N_1582);
xor U1653 (N_1653,N_1395,N_1356);
or U1654 (N_1654,N_1200,N_1380);
nor U1655 (N_1655,N_1555,N_1487);
xor U1656 (N_1656,N_1375,N_1565);
nor U1657 (N_1657,N_1242,N_1333);
and U1658 (N_1658,N_1511,N_1354);
and U1659 (N_1659,N_1518,N_1231);
and U1660 (N_1660,N_1211,N_1284);
and U1661 (N_1661,N_1476,N_1340);
xor U1662 (N_1662,N_1495,N_1291);
nand U1663 (N_1663,N_1334,N_1499);
nand U1664 (N_1664,N_1279,N_1464);
and U1665 (N_1665,N_1446,N_1488);
xor U1666 (N_1666,N_1507,N_1233);
nand U1667 (N_1667,N_1253,N_1377);
nand U1668 (N_1668,N_1293,N_1505);
nor U1669 (N_1669,N_1598,N_1440);
xor U1670 (N_1670,N_1264,N_1219);
xor U1671 (N_1671,N_1460,N_1410);
and U1672 (N_1672,N_1339,N_1463);
or U1673 (N_1673,N_1385,N_1486);
and U1674 (N_1674,N_1500,N_1386);
or U1675 (N_1675,N_1260,N_1374);
xor U1676 (N_1676,N_1212,N_1337);
nand U1677 (N_1677,N_1305,N_1470);
or U1678 (N_1678,N_1277,N_1344);
nand U1679 (N_1679,N_1338,N_1573);
nor U1680 (N_1680,N_1303,N_1388);
or U1681 (N_1681,N_1312,N_1404);
and U1682 (N_1682,N_1390,N_1578);
xnor U1683 (N_1683,N_1235,N_1237);
nor U1684 (N_1684,N_1389,N_1588);
and U1685 (N_1685,N_1376,N_1533);
nor U1686 (N_1686,N_1530,N_1412);
and U1687 (N_1687,N_1553,N_1423);
xnor U1688 (N_1688,N_1301,N_1281);
and U1689 (N_1689,N_1201,N_1502);
or U1690 (N_1690,N_1269,N_1439);
nor U1691 (N_1691,N_1204,N_1245);
nand U1692 (N_1692,N_1534,N_1275);
nand U1693 (N_1693,N_1561,N_1567);
nor U1694 (N_1694,N_1206,N_1417);
and U1695 (N_1695,N_1568,N_1230);
xnor U1696 (N_1696,N_1329,N_1541);
or U1697 (N_1697,N_1421,N_1469);
nand U1698 (N_1698,N_1247,N_1366);
nor U1699 (N_1699,N_1579,N_1528);
nand U1700 (N_1700,N_1296,N_1360);
nor U1701 (N_1701,N_1315,N_1263);
nand U1702 (N_1702,N_1400,N_1401);
nor U1703 (N_1703,N_1535,N_1229);
xor U1704 (N_1704,N_1294,N_1347);
or U1705 (N_1705,N_1236,N_1501);
nand U1706 (N_1706,N_1586,N_1429);
and U1707 (N_1707,N_1478,N_1595);
or U1708 (N_1708,N_1257,N_1325);
nor U1709 (N_1709,N_1357,N_1308);
and U1710 (N_1710,N_1270,N_1292);
and U1711 (N_1711,N_1526,N_1540);
and U1712 (N_1712,N_1362,N_1210);
nor U1713 (N_1713,N_1432,N_1594);
nor U1714 (N_1714,N_1299,N_1295);
nand U1715 (N_1715,N_1218,N_1278);
and U1716 (N_1716,N_1545,N_1441);
and U1717 (N_1717,N_1413,N_1323);
nand U1718 (N_1718,N_1208,N_1491);
nand U1719 (N_1719,N_1398,N_1596);
and U1720 (N_1720,N_1583,N_1273);
nand U1721 (N_1721,N_1267,N_1328);
and U1722 (N_1722,N_1551,N_1549);
and U1723 (N_1723,N_1520,N_1317);
xor U1724 (N_1724,N_1355,N_1574);
xor U1725 (N_1725,N_1271,N_1364);
xor U1726 (N_1726,N_1519,N_1472);
nand U1727 (N_1727,N_1494,N_1537);
xor U1728 (N_1728,N_1409,N_1369);
nor U1729 (N_1729,N_1489,N_1297);
or U1730 (N_1730,N_1203,N_1550);
xor U1731 (N_1731,N_1254,N_1285);
xor U1732 (N_1732,N_1418,N_1381);
xnor U1733 (N_1733,N_1482,N_1438);
nor U1734 (N_1734,N_1523,N_1454);
nand U1735 (N_1735,N_1384,N_1307);
xnor U1736 (N_1736,N_1282,N_1363);
nand U1737 (N_1737,N_1298,N_1205);
xnor U1738 (N_1738,N_1462,N_1485);
and U1739 (N_1739,N_1266,N_1498);
and U1740 (N_1740,N_1322,N_1225);
or U1741 (N_1741,N_1584,N_1406);
nor U1742 (N_1742,N_1274,N_1590);
and U1743 (N_1743,N_1559,N_1475);
xor U1744 (N_1744,N_1371,N_1327);
or U1745 (N_1745,N_1442,N_1290);
and U1746 (N_1746,N_1503,N_1445);
xor U1747 (N_1747,N_1397,N_1265);
xor U1748 (N_1748,N_1509,N_1349);
and U1749 (N_1749,N_1394,N_1226);
or U1750 (N_1750,N_1228,N_1246);
or U1751 (N_1751,N_1403,N_1546);
nand U1752 (N_1752,N_1370,N_1365);
and U1753 (N_1753,N_1321,N_1458);
xor U1754 (N_1754,N_1352,N_1286);
nand U1755 (N_1755,N_1342,N_1416);
xor U1756 (N_1756,N_1558,N_1240);
or U1757 (N_1757,N_1238,N_1320);
and U1758 (N_1758,N_1484,N_1359);
nor U1759 (N_1759,N_1524,N_1504);
xor U1760 (N_1760,N_1563,N_1451);
and U1761 (N_1761,N_1326,N_1268);
nand U1762 (N_1762,N_1575,N_1471);
nand U1763 (N_1763,N_1473,N_1580);
or U1764 (N_1764,N_1465,N_1532);
xnor U1765 (N_1765,N_1569,N_1497);
or U1766 (N_1766,N_1516,N_1367);
nand U1767 (N_1767,N_1564,N_1309);
xnor U1768 (N_1768,N_1202,N_1318);
xor U1769 (N_1769,N_1515,N_1435);
nand U1770 (N_1770,N_1597,N_1543);
and U1771 (N_1771,N_1313,N_1258);
or U1772 (N_1772,N_1566,N_1392);
or U1773 (N_1773,N_1221,N_1283);
nor U1774 (N_1774,N_1517,N_1538);
or U1775 (N_1775,N_1402,N_1214);
nand U1776 (N_1776,N_1234,N_1383);
nand U1777 (N_1777,N_1426,N_1232);
or U1778 (N_1778,N_1316,N_1304);
and U1779 (N_1779,N_1449,N_1466);
and U1780 (N_1780,N_1255,N_1525);
nor U1781 (N_1781,N_1373,N_1591);
and U1782 (N_1782,N_1288,N_1514);
xnor U1783 (N_1783,N_1508,N_1585);
and U1784 (N_1784,N_1256,N_1382);
or U1785 (N_1785,N_1587,N_1461);
xnor U1786 (N_1786,N_1220,N_1599);
or U1787 (N_1787,N_1241,N_1589);
xor U1788 (N_1788,N_1554,N_1547);
nand U1789 (N_1789,N_1314,N_1343);
and U1790 (N_1790,N_1411,N_1444);
xor U1791 (N_1791,N_1243,N_1227);
xnor U1792 (N_1792,N_1433,N_1379);
and U1793 (N_1793,N_1399,N_1572);
xor U1794 (N_1794,N_1252,N_1276);
xnor U1795 (N_1795,N_1496,N_1222);
and U1796 (N_1796,N_1593,N_1552);
xnor U1797 (N_1797,N_1510,N_1353);
and U1798 (N_1798,N_1512,N_1331);
nor U1799 (N_1799,N_1436,N_1306);
and U1800 (N_1800,N_1256,N_1444);
nor U1801 (N_1801,N_1386,N_1460);
xor U1802 (N_1802,N_1356,N_1260);
xnor U1803 (N_1803,N_1550,N_1234);
nor U1804 (N_1804,N_1560,N_1288);
xor U1805 (N_1805,N_1246,N_1521);
xor U1806 (N_1806,N_1522,N_1318);
and U1807 (N_1807,N_1380,N_1433);
xor U1808 (N_1808,N_1359,N_1517);
nor U1809 (N_1809,N_1223,N_1490);
nand U1810 (N_1810,N_1364,N_1307);
and U1811 (N_1811,N_1271,N_1343);
nand U1812 (N_1812,N_1430,N_1449);
xor U1813 (N_1813,N_1346,N_1307);
nand U1814 (N_1814,N_1220,N_1478);
or U1815 (N_1815,N_1318,N_1536);
and U1816 (N_1816,N_1543,N_1482);
and U1817 (N_1817,N_1446,N_1316);
nor U1818 (N_1818,N_1569,N_1589);
and U1819 (N_1819,N_1213,N_1380);
or U1820 (N_1820,N_1398,N_1307);
xor U1821 (N_1821,N_1277,N_1428);
xnor U1822 (N_1822,N_1580,N_1235);
and U1823 (N_1823,N_1464,N_1363);
or U1824 (N_1824,N_1220,N_1366);
or U1825 (N_1825,N_1348,N_1378);
and U1826 (N_1826,N_1420,N_1332);
or U1827 (N_1827,N_1363,N_1370);
nor U1828 (N_1828,N_1322,N_1463);
and U1829 (N_1829,N_1360,N_1415);
and U1830 (N_1830,N_1429,N_1367);
xor U1831 (N_1831,N_1341,N_1362);
nor U1832 (N_1832,N_1579,N_1556);
xor U1833 (N_1833,N_1573,N_1547);
and U1834 (N_1834,N_1276,N_1323);
xor U1835 (N_1835,N_1257,N_1267);
and U1836 (N_1836,N_1541,N_1298);
xor U1837 (N_1837,N_1271,N_1379);
nand U1838 (N_1838,N_1592,N_1483);
xor U1839 (N_1839,N_1204,N_1313);
nand U1840 (N_1840,N_1509,N_1286);
nor U1841 (N_1841,N_1562,N_1587);
xnor U1842 (N_1842,N_1254,N_1278);
xnor U1843 (N_1843,N_1496,N_1270);
xor U1844 (N_1844,N_1354,N_1373);
and U1845 (N_1845,N_1235,N_1566);
or U1846 (N_1846,N_1227,N_1363);
xor U1847 (N_1847,N_1421,N_1347);
nand U1848 (N_1848,N_1256,N_1462);
nand U1849 (N_1849,N_1515,N_1406);
or U1850 (N_1850,N_1365,N_1437);
and U1851 (N_1851,N_1264,N_1431);
nor U1852 (N_1852,N_1291,N_1224);
nor U1853 (N_1853,N_1307,N_1507);
nand U1854 (N_1854,N_1412,N_1248);
xor U1855 (N_1855,N_1270,N_1441);
nand U1856 (N_1856,N_1423,N_1541);
or U1857 (N_1857,N_1317,N_1215);
nand U1858 (N_1858,N_1207,N_1335);
and U1859 (N_1859,N_1399,N_1377);
or U1860 (N_1860,N_1507,N_1477);
nor U1861 (N_1861,N_1478,N_1418);
and U1862 (N_1862,N_1457,N_1337);
xor U1863 (N_1863,N_1592,N_1274);
and U1864 (N_1864,N_1460,N_1478);
nor U1865 (N_1865,N_1292,N_1308);
nor U1866 (N_1866,N_1298,N_1317);
nand U1867 (N_1867,N_1434,N_1361);
nand U1868 (N_1868,N_1317,N_1515);
nand U1869 (N_1869,N_1248,N_1446);
nand U1870 (N_1870,N_1228,N_1385);
nand U1871 (N_1871,N_1491,N_1252);
nor U1872 (N_1872,N_1212,N_1498);
xnor U1873 (N_1873,N_1364,N_1250);
nand U1874 (N_1874,N_1393,N_1283);
and U1875 (N_1875,N_1359,N_1535);
or U1876 (N_1876,N_1200,N_1216);
or U1877 (N_1877,N_1296,N_1218);
nor U1878 (N_1878,N_1503,N_1205);
and U1879 (N_1879,N_1358,N_1498);
nor U1880 (N_1880,N_1320,N_1387);
or U1881 (N_1881,N_1588,N_1438);
nor U1882 (N_1882,N_1540,N_1570);
and U1883 (N_1883,N_1499,N_1547);
xor U1884 (N_1884,N_1246,N_1254);
xor U1885 (N_1885,N_1489,N_1436);
or U1886 (N_1886,N_1305,N_1582);
nor U1887 (N_1887,N_1255,N_1484);
nand U1888 (N_1888,N_1298,N_1415);
nand U1889 (N_1889,N_1506,N_1533);
nor U1890 (N_1890,N_1391,N_1566);
or U1891 (N_1891,N_1469,N_1525);
or U1892 (N_1892,N_1478,N_1292);
and U1893 (N_1893,N_1370,N_1594);
or U1894 (N_1894,N_1360,N_1506);
and U1895 (N_1895,N_1486,N_1209);
xnor U1896 (N_1896,N_1419,N_1568);
xnor U1897 (N_1897,N_1504,N_1282);
nand U1898 (N_1898,N_1516,N_1246);
or U1899 (N_1899,N_1597,N_1593);
and U1900 (N_1900,N_1243,N_1263);
nor U1901 (N_1901,N_1472,N_1312);
nor U1902 (N_1902,N_1440,N_1322);
nor U1903 (N_1903,N_1390,N_1537);
or U1904 (N_1904,N_1538,N_1440);
or U1905 (N_1905,N_1380,N_1458);
nand U1906 (N_1906,N_1341,N_1443);
nor U1907 (N_1907,N_1214,N_1397);
and U1908 (N_1908,N_1388,N_1362);
nand U1909 (N_1909,N_1522,N_1445);
nor U1910 (N_1910,N_1466,N_1566);
nor U1911 (N_1911,N_1572,N_1354);
nand U1912 (N_1912,N_1307,N_1229);
or U1913 (N_1913,N_1262,N_1271);
xor U1914 (N_1914,N_1494,N_1320);
xnor U1915 (N_1915,N_1201,N_1243);
nand U1916 (N_1916,N_1379,N_1377);
and U1917 (N_1917,N_1393,N_1293);
or U1918 (N_1918,N_1349,N_1326);
nor U1919 (N_1919,N_1488,N_1406);
or U1920 (N_1920,N_1208,N_1262);
nand U1921 (N_1921,N_1543,N_1328);
nor U1922 (N_1922,N_1345,N_1481);
nor U1923 (N_1923,N_1207,N_1539);
or U1924 (N_1924,N_1263,N_1326);
and U1925 (N_1925,N_1337,N_1304);
nand U1926 (N_1926,N_1580,N_1484);
xnor U1927 (N_1927,N_1209,N_1251);
nor U1928 (N_1928,N_1488,N_1439);
xnor U1929 (N_1929,N_1597,N_1591);
and U1930 (N_1930,N_1513,N_1275);
nand U1931 (N_1931,N_1409,N_1514);
xnor U1932 (N_1932,N_1331,N_1383);
xnor U1933 (N_1933,N_1543,N_1473);
or U1934 (N_1934,N_1581,N_1448);
nand U1935 (N_1935,N_1483,N_1242);
nor U1936 (N_1936,N_1558,N_1410);
xnor U1937 (N_1937,N_1533,N_1236);
and U1938 (N_1938,N_1465,N_1276);
nor U1939 (N_1939,N_1557,N_1255);
nor U1940 (N_1940,N_1549,N_1382);
or U1941 (N_1941,N_1378,N_1306);
nand U1942 (N_1942,N_1230,N_1398);
xnor U1943 (N_1943,N_1559,N_1484);
nor U1944 (N_1944,N_1553,N_1322);
or U1945 (N_1945,N_1519,N_1582);
or U1946 (N_1946,N_1218,N_1402);
or U1947 (N_1947,N_1495,N_1429);
nor U1948 (N_1948,N_1459,N_1357);
and U1949 (N_1949,N_1326,N_1211);
nor U1950 (N_1950,N_1395,N_1585);
xnor U1951 (N_1951,N_1506,N_1256);
xor U1952 (N_1952,N_1424,N_1457);
nand U1953 (N_1953,N_1367,N_1340);
nand U1954 (N_1954,N_1241,N_1507);
nor U1955 (N_1955,N_1489,N_1534);
nand U1956 (N_1956,N_1571,N_1502);
and U1957 (N_1957,N_1541,N_1324);
nand U1958 (N_1958,N_1201,N_1310);
nor U1959 (N_1959,N_1568,N_1242);
or U1960 (N_1960,N_1566,N_1542);
and U1961 (N_1961,N_1502,N_1508);
nor U1962 (N_1962,N_1380,N_1237);
xor U1963 (N_1963,N_1470,N_1593);
nand U1964 (N_1964,N_1290,N_1299);
xnor U1965 (N_1965,N_1208,N_1209);
or U1966 (N_1966,N_1380,N_1447);
nand U1967 (N_1967,N_1208,N_1564);
nor U1968 (N_1968,N_1319,N_1271);
or U1969 (N_1969,N_1251,N_1416);
nor U1970 (N_1970,N_1300,N_1305);
or U1971 (N_1971,N_1477,N_1265);
xnor U1972 (N_1972,N_1423,N_1309);
and U1973 (N_1973,N_1474,N_1450);
and U1974 (N_1974,N_1240,N_1436);
and U1975 (N_1975,N_1209,N_1287);
or U1976 (N_1976,N_1514,N_1507);
or U1977 (N_1977,N_1496,N_1275);
xor U1978 (N_1978,N_1507,N_1218);
nand U1979 (N_1979,N_1229,N_1503);
or U1980 (N_1980,N_1201,N_1466);
and U1981 (N_1981,N_1516,N_1243);
xnor U1982 (N_1982,N_1590,N_1207);
nand U1983 (N_1983,N_1262,N_1432);
and U1984 (N_1984,N_1288,N_1465);
and U1985 (N_1985,N_1239,N_1277);
nor U1986 (N_1986,N_1418,N_1420);
xnor U1987 (N_1987,N_1348,N_1430);
and U1988 (N_1988,N_1584,N_1466);
nand U1989 (N_1989,N_1253,N_1290);
xnor U1990 (N_1990,N_1599,N_1352);
or U1991 (N_1991,N_1595,N_1322);
nand U1992 (N_1992,N_1454,N_1267);
nor U1993 (N_1993,N_1341,N_1385);
nor U1994 (N_1994,N_1268,N_1332);
nor U1995 (N_1995,N_1559,N_1418);
or U1996 (N_1996,N_1468,N_1570);
nand U1997 (N_1997,N_1380,N_1423);
or U1998 (N_1998,N_1500,N_1414);
nand U1999 (N_1999,N_1537,N_1257);
xnor U2000 (N_2000,N_1802,N_1831);
nand U2001 (N_2001,N_1862,N_1806);
xor U2002 (N_2002,N_1746,N_1638);
nand U2003 (N_2003,N_1763,N_1827);
nor U2004 (N_2004,N_1602,N_1899);
xnor U2005 (N_2005,N_1679,N_1909);
nor U2006 (N_2006,N_1817,N_1907);
xor U2007 (N_2007,N_1896,N_1803);
and U2008 (N_2008,N_1610,N_1676);
and U2009 (N_2009,N_1799,N_1880);
or U2010 (N_2010,N_1953,N_1965);
nor U2011 (N_2011,N_1925,N_1888);
nand U2012 (N_2012,N_1689,N_1807);
xor U2013 (N_2013,N_1667,N_1875);
and U2014 (N_2014,N_1708,N_1723);
and U2015 (N_2015,N_1881,N_1669);
and U2016 (N_2016,N_1765,N_1865);
or U2017 (N_2017,N_1911,N_1663);
and U2018 (N_2018,N_1857,N_1939);
nand U2019 (N_2019,N_1915,N_1717);
nor U2020 (N_2020,N_1617,N_1928);
nor U2021 (N_2021,N_1790,N_1760);
nor U2022 (N_2022,N_1824,N_1737);
nor U2023 (N_2023,N_1890,N_1812);
and U2024 (N_2024,N_1701,N_1629);
and U2025 (N_2025,N_1601,N_1715);
nor U2026 (N_2026,N_1963,N_1945);
nand U2027 (N_2027,N_1794,N_1600);
nor U2028 (N_2028,N_1648,N_1886);
nand U2029 (N_2029,N_1929,N_1635);
and U2030 (N_2030,N_1613,N_1959);
xor U2031 (N_2031,N_1835,N_1893);
nor U2032 (N_2032,N_1946,N_1797);
nand U2033 (N_2033,N_1722,N_1764);
xor U2034 (N_2034,N_1816,N_1993);
nand U2035 (N_2035,N_1735,N_1690);
and U2036 (N_2036,N_1672,N_1762);
nand U2037 (N_2037,N_1604,N_1673);
nand U2038 (N_2038,N_1988,N_1871);
nor U2039 (N_2039,N_1826,N_1664);
and U2040 (N_2040,N_1661,N_1620);
nor U2041 (N_2041,N_1718,N_1753);
xor U2042 (N_2042,N_1720,N_1640);
nor U2043 (N_2043,N_1754,N_1972);
xor U2044 (N_2044,N_1630,N_1996);
xnor U2045 (N_2045,N_1631,N_1736);
xor U2046 (N_2046,N_1651,N_1784);
and U2047 (N_2047,N_1788,N_1787);
or U2048 (N_2048,N_1655,N_1728);
xor U2049 (N_2049,N_1952,N_1776);
and U2050 (N_2050,N_1639,N_1800);
nor U2051 (N_2051,N_1713,N_1805);
and U2052 (N_2052,N_1964,N_1666);
xnor U2053 (N_2053,N_1898,N_1727);
nor U2054 (N_2054,N_1724,N_1742);
nand U2055 (N_2055,N_1744,N_1912);
xnor U2056 (N_2056,N_1984,N_1821);
or U2057 (N_2057,N_1968,N_1844);
xor U2058 (N_2058,N_1948,N_1632);
xnor U2059 (N_2059,N_1813,N_1641);
or U2060 (N_2060,N_1808,N_1756);
and U2061 (N_2061,N_1927,N_1955);
and U2062 (N_2062,N_1726,N_1654);
nand U2063 (N_2063,N_1677,N_1643);
xnor U2064 (N_2064,N_1774,N_1627);
nand U2065 (N_2065,N_1652,N_1766);
nand U2066 (N_2066,N_1930,N_1628);
or U2067 (N_2067,N_1660,N_1646);
xnor U2068 (N_2068,N_1851,N_1889);
or U2069 (N_2069,N_1947,N_1850);
or U2070 (N_2070,N_1789,N_1819);
xor U2071 (N_2071,N_1608,N_1810);
nand U2072 (N_2072,N_1804,N_1860);
xnor U2073 (N_2073,N_1868,N_1864);
and U2074 (N_2074,N_1838,N_1693);
xor U2075 (N_2075,N_1759,N_1944);
nand U2076 (N_2076,N_1801,N_1607);
and U2077 (N_2077,N_1791,N_1874);
nand U2078 (N_2078,N_1936,N_1606);
and U2079 (N_2079,N_1935,N_1702);
nor U2080 (N_2080,N_1998,N_1994);
nor U2081 (N_2081,N_1719,N_1872);
or U2082 (N_2082,N_1616,N_1782);
nand U2083 (N_2083,N_1894,N_1703);
nor U2084 (N_2084,N_1849,N_1924);
and U2085 (N_2085,N_1839,N_1665);
xnor U2086 (N_2086,N_1992,N_1709);
and U2087 (N_2087,N_1873,N_1603);
nand U2088 (N_2088,N_1721,N_1657);
nor U2089 (N_2089,N_1882,N_1830);
nor U2090 (N_2090,N_1979,N_1637);
and U2091 (N_2091,N_1969,N_1623);
and U2092 (N_2092,N_1842,N_1745);
or U2093 (N_2093,N_1732,N_1985);
and U2094 (N_2094,N_1908,N_1956);
and U2095 (N_2095,N_1662,N_1642);
and U2096 (N_2096,N_1751,N_1905);
and U2097 (N_2097,N_1783,N_1738);
nand U2098 (N_2098,N_1752,N_1919);
xor U2099 (N_2099,N_1845,N_1768);
and U2100 (N_2100,N_1761,N_1855);
and U2101 (N_2101,N_1901,N_1618);
and U2102 (N_2102,N_1622,N_1699);
nor U2103 (N_2103,N_1983,N_1913);
and U2104 (N_2104,N_1614,N_1989);
or U2105 (N_2105,N_1695,N_1793);
and U2106 (N_2106,N_1926,N_1848);
nand U2107 (N_2107,N_1685,N_1931);
nor U2108 (N_2108,N_1981,N_1974);
xor U2109 (N_2109,N_1743,N_1692);
or U2110 (N_2110,N_1971,N_1841);
xor U2111 (N_2111,N_1770,N_1859);
or U2112 (N_2112,N_1847,N_1694);
or U2113 (N_2113,N_1649,N_1858);
xor U2114 (N_2114,N_1854,N_1633);
xor U2115 (N_2115,N_1885,N_1786);
nand U2116 (N_2116,N_1906,N_1798);
nand U2117 (N_2117,N_1796,N_1834);
nand U2118 (N_2118,N_1653,N_1837);
nor U2119 (N_2119,N_1914,N_1611);
and U2120 (N_2120,N_1659,N_1895);
nor U2121 (N_2121,N_1686,N_1792);
nand U2122 (N_2122,N_1769,N_1741);
and U2123 (N_2123,N_1892,N_1684);
and U2124 (N_2124,N_1777,N_1619);
nor U2125 (N_2125,N_1973,N_1934);
or U2126 (N_2126,N_1887,N_1867);
xnor U2127 (N_2127,N_1932,N_1997);
nor U2128 (N_2128,N_1883,N_1832);
xnor U2129 (N_2129,N_1605,N_1878);
xor U2130 (N_2130,N_1877,N_1903);
xnor U2131 (N_2131,N_1897,N_1902);
nand U2132 (N_2132,N_1975,N_1626);
xor U2133 (N_2133,N_1706,N_1986);
nor U2134 (N_2134,N_1815,N_1836);
nor U2135 (N_2135,N_1863,N_1683);
or U2136 (N_2136,N_1818,N_1962);
or U2137 (N_2137,N_1977,N_1991);
or U2138 (N_2138,N_1904,N_1705);
nor U2139 (N_2139,N_1829,N_1682);
and U2140 (N_2140,N_1814,N_1866);
xor U2141 (N_2141,N_1711,N_1978);
nand U2142 (N_2142,N_1757,N_1938);
or U2143 (N_2143,N_1670,N_1917);
nor U2144 (N_2144,N_1671,N_1876);
xor U2145 (N_2145,N_1731,N_1729);
and U2146 (N_2146,N_1976,N_1923);
and U2147 (N_2147,N_1809,N_1748);
and U2148 (N_2148,N_1674,N_1823);
and U2149 (N_2149,N_1767,N_1922);
or U2150 (N_2150,N_1716,N_1987);
or U2151 (N_2151,N_1843,N_1749);
or U2152 (N_2152,N_1697,N_1937);
nor U2153 (N_2153,N_1636,N_1696);
and U2154 (N_2154,N_1698,N_1691);
nand U2155 (N_2155,N_1950,N_1921);
and U2156 (N_2156,N_1949,N_1750);
nand U2157 (N_2157,N_1621,N_1733);
or U2158 (N_2158,N_1833,N_1775);
xnor U2159 (N_2159,N_1852,N_1811);
xor U2160 (N_2160,N_1758,N_1933);
nor U2161 (N_2161,N_1943,N_1778);
nand U2162 (N_2162,N_1980,N_1918);
nor U2163 (N_2163,N_1870,N_1781);
nand U2164 (N_2164,N_1967,N_1700);
xor U2165 (N_2165,N_1785,N_1970);
nand U2166 (N_2166,N_1916,N_1707);
nand U2167 (N_2167,N_1658,N_1725);
nand U2168 (N_2168,N_1644,N_1820);
nor U2169 (N_2169,N_1966,N_1856);
nand U2170 (N_2170,N_1675,N_1624);
nand U2171 (N_2171,N_1957,N_1941);
nand U2172 (N_2172,N_1999,N_1954);
nand U2173 (N_2173,N_1747,N_1704);
or U2174 (N_2174,N_1740,N_1958);
and U2175 (N_2175,N_1840,N_1739);
xnor U2176 (N_2176,N_1609,N_1861);
xnor U2177 (N_2177,N_1714,N_1634);
xnor U2178 (N_2178,N_1712,N_1884);
and U2179 (N_2179,N_1645,N_1853);
and U2180 (N_2180,N_1772,N_1940);
xor U2181 (N_2181,N_1647,N_1982);
and U2182 (N_2182,N_1656,N_1942);
and U2183 (N_2183,N_1773,N_1734);
nor U2184 (N_2184,N_1795,N_1961);
nor U2185 (N_2185,N_1612,N_1825);
nor U2186 (N_2186,N_1900,N_1680);
nor U2187 (N_2187,N_1668,N_1920);
and U2188 (N_2188,N_1625,N_1678);
and U2189 (N_2189,N_1846,N_1780);
xor U2190 (N_2190,N_1688,N_1779);
nor U2191 (N_2191,N_1990,N_1995);
xnor U2192 (N_2192,N_1650,N_1730);
and U2193 (N_2193,N_1879,N_1910);
and U2194 (N_2194,N_1869,N_1960);
nor U2195 (N_2195,N_1710,N_1822);
or U2196 (N_2196,N_1615,N_1828);
nor U2197 (N_2197,N_1681,N_1951);
and U2198 (N_2198,N_1771,N_1755);
and U2199 (N_2199,N_1891,N_1687);
nand U2200 (N_2200,N_1758,N_1727);
nor U2201 (N_2201,N_1629,N_1792);
nand U2202 (N_2202,N_1701,N_1870);
nor U2203 (N_2203,N_1711,N_1848);
xnor U2204 (N_2204,N_1859,N_1939);
xnor U2205 (N_2205,N_1663,N_1704);
nor U2206 (N_2206,N_1928,N_1615);
and U2207 (N_2207,N_1860,N_1771);
nor U2208 (N_2208,N_1710,N_1934);
and U2209 (N_2209,N_1681,N_1840);
xor U2210 (N_2210,N_1605,N_1806);
or U2211 (N_2211,N_1896,N_1845);
and U2212 (N_2212,N_1813,N_1925);
xnor U2213 (N_2213,N_1736,N_1801);
nand U2214 (N_2214,N_1731,N_1931);
and U2215 (N_2215,N_1718,N_1789);
nand U2216 (N_2216,N_1656,N_1874);
xnor U2217 (N_2217,N_1700,N_1604);
nor U2218 (N_2218,N_1811,N_1678);
xnor U2219 (N_2219,N_1857,N_1657);
or U2220 (N_2220,N_1626,N_1909);
nor U2221 (N_2221,N_1746,N_1930);
or U2222 (N_2222,N_1907,N_1880);
nor U2223 (N_2223,N_1895,N_1870);
and U2224 (N_2224,N_1798,N_1633);
xor U2225 (N_2225,N_1693,N_1725);
nand U2226 (N_2226,N_1982,N_1807);
and U2227 (N_2227,N_1996,N_1927);
and U2228 (N_2228,N_1881,N_1687);
xor U2229 (N_2229,N_1609,N_1653);
or U2230 (N_2230,N_1642,N_1851);
xnor U2231 (N_2231,N_1953,N_1905);
nor U2232 (N_2232,N_1833,N_1630);
and U2233 (N_2233,N_1705,N_1605);
xor U2234 (N_2234,N_1978,N_1983);
or U2235 (N_2235,N_1817,N_1911);
or U2236 (N_2236,N_1763,N_1741);
xor U2237 (N_2237,N_1666,N_1972);
or U2238 (N_2238,N_1943,N_1996);
and U2239 (N_2239,N_1978,N_1847);
nand U2240 (N_2240,N_1855,N_1618);
nand U2241 (N_2241,N_1881,N_1625);
nor U2242 (N_2242,N_1844,N_1988);
xor U2243 (N_2243,N_1808,N_1769);
or U2244 (N_2244,N_1672,N_1830);
and U2245 (N_2245,N_1961,N_1991);
and U2246 (N_2246,N_1636,N_1786);
and U2247 (N_2247,N_1822,N_1790);
xor U2248 (N_2248,N_1972,N_1689);
nor U2249 (N_2249,N_1863,N_1857);
nor U2250 (N_2250,N_1663,N_1628);
nand U2251 (N_2251,N_1773,N_1607);
nor U2252 (N_2252,N_1869,N_1922);
or U2253 (N_2253,N_1669,N_1832);
nor U2254 (N_2254,N_1697,N_1970);
nand U2255 (N_2255,N_1830,N_1619);
nor U2256 (N_2256,N_1639,N_1935);
and U2257 (N_2257,N_1855,N_1706);
nor U2258 (N_2258,N_1658,N_1804);
and U2259 (N_2259,N_1727,N_1875);
xor U2260 (N_2260,N_1626,N_1771);
nand U2261 (N_2261,N_1898,N_1821);
nor U2262 (N_2262,N_1791,N_1631);
nor U2263 (N_2263,N_1860,N_1687);
or U2264 (N_2264,N_1617,N_1657);
xor U2265 (N_2265,N_1980,N_1602);
nand U2266 (N_2266,N_1878,N_1688);
nand U2267 (N_2267,N_1845,N_1945);
and U2268 (N_2268,N_1708,N_1769);
or U2269 (N_2269,N_1839,N_1820);
or U2270 (N_2270,N_1807,N_1691);
xor U2271 (N_2271,N_1802,N_1716);
or U2272 (N_2272,N_1974,N_1979);
or U2273 (N_2273,N_1660,N_1653);
and U2274 (N_2274,N_1604,N_1835);
or U2275 (N_2275,N_1739,N_1886);
nand U2276 (N_2276,N_1663,N_1646);
and U2277 (N_2277,N_1912,N_1885);
nand U2278 (N_2278,N_1747,N_1701);
or U2279 (N_2279,N_1608,N_1614);
or U2280 (N_2280,N_1639,N_1749);
nor U2281 (N_2281,N_1872,N_1877);
nand U2282 (N_2282,N_1943,N_1771);
nand U2283 (N_2283,N_1894,N_1949);
and U2284 (N_2284,N_1698,N_1920);
or U2285 (N_2285,N_1807,N_1960);
xnor U2286 (N_2286,N_1954,N_1754);
nor U2287 (N_2287,N_1665,N_1929);
nand U2288 (N_2288,N_1775,N_1786);
or U2289 (N_2289,N_1848,N_1615);
nand U2290 (N_2290,N_1904,N_1992);
nor U2291 (N_2291,N_1726,N_1763);
or U2292 (N_2292,N_1943,N_1805);
nand U2293 (N_2293,N_1901,N_1783);
and U2294 (N_2294,N_1814,N_1848);
or U2295 (N_2295,N_1679,N_1763);
nor U2296 (N_2296,N_1682,N_1988);
nor U2297 (N_2297,N_1610,N_1924);
xnor U2298 (N_2298,N_1669,N_1639);
xor U2299 (N_2299,N_1745,N_1932);
nor U2300 (N_2300,N_1607,N_1966);
or U2301 (N_2301,N_1639,N_1787);
xor U2302 (N_2302,N_1885,N_1748);
or U2303 (N_2303,N_1729,N_1703);
nand U2304 (N_2304,N_1894,N_1757);
nor U2305 (N_2305,N_1720,N_1705);
and U2306 (N_2306,N_1869,N_1976);
xor U2307 (N_2307,N_1827,N_1769);
nand U2308 (N_2308,N_1974,N_1712);
nand U2309 (N_2309,N_1654,N_1732);
nor U2310 (N_2310,N_1790,N_1750);
xnor U2311 (N_2311,N_1934,N_1702);
and U2312 (N_2312,N_1606,N_1683);
nor U2313 (N_2313,N_1605,N_1975);
xor U2314 (N_2314,N_1617,N_1703);
and U2315 (N_2315,N_1940,N_1897);
or U2316 (N_2316,N_1830,N_1842);
or U2317 (N_2317,N_1920,N_1751);
nor U2318 (N_2318,N_1678,N_1729);
xor U2319 (N_2319,N_1630,N_1969);
and U2320 (N_2320,N_1965,N_1972);
xnor U2321 (N_2321,N_1865,N_1759);
nor U2322 (N_2322,N_1998,N_1632);
nor U2323 (N_2323,N_1632,N_1756);
nor U2324 (N_2324,N_1756,N_1679);
or U2325 (N_2325,N_1732,N_1735);
and U2326 (N_2326,N_1607,N_1723);
and U2327 (N_2327,N_1793,N_1713);
xnor U2328 (N_2328,N_1871,N_1827);
nand U2329 (N_2329,N_1745,N_1665);
or U2330 (N_2330,N_1734,N_1858);
and U2331 (N_2331,N_1833,N_1634);
nand U2332 (N_2332,N_1852,N_1922);
nor U2333 (N_2333,N_1883,N_1775);
or U2334 (N_2334,N_1940,N_1941);
nor U2335 (N_2335,N_1662,N_1987);
and U2336 (N_2336,N_1736,N_1888);
or U2337 (N_2337,N_1756,N_1914);
xnor U2338 (N_2338,N_1817,N_1709);
nand U2339 (N_2339,N_1681,N_1999);
nand U2340 (N_2340,N_1926,N_1654);
and U2341 (N_2341,N_1784,N_1638);
or U2342 (N_2342,N_1769,N_1876);
nand U2343 (N_2343,N_1714,N_1734);
and U2344 (N_2344,N_1859,N_1745);
or U2345 (N_2345,N_1842,N_1648);
or U2346 (N_2346,N_1807,N_1849);
nor U2347 (N_2347,N_1630,N_1767);
and U2348 (N_2348,N_1841,N_1774);
nor U2349 (N_2349,N_1838,N_1632);
xor U2350 (N_2350,N_1670,N_1612);
or U2351 (N_2351,N_1758,N_1934);
xnor U2352 (N_2352,N_1955,N_1740);
xor U2353 (N_2353,N_1798,N_1614);
nand U2354 (N_2354,N_1829,N_1707);
xnor U2355 (N_2355,N_1916,N_1640);
nor U2356 (N_2356,N_1621,N_1937);
and U2357 (N_2357,N_1880,N_1894);
nand U2358 (N_2358,N_1642,N_1944);
and U2359 (N_2359,N_1923,N_1889);
nand U2360 (N_2360,N_1992,N_1921);
nand U2361 (N_2361,N_1726,N_1602);
nand U2362 (N_2362,N_1797,N_1917);
and U2363 (N_2363,N_1891,N_1770);
xnor U2364 (N_2364,N_1727,N_1966);
xnor U2365 (N_2365,N_1863,N_1901);
nor U2366 (N_2366,N_1797,N_1836);
nand U2367 (N_2367,N_1842,N_1802);
and U2368 (N_2368,N_1721,N_1678);
nor U2369 (N_2369,N_1775,N_1972);
xnor U2370 (N_2370,N_1925,N_1765);
or U2371 (N_2371,N_1964,N_1903);
nand U2372 (N_2372,N_1649,N_1667);
nor U2373 (N_2373,N_1759,N_1877);
xor U2374 (N_2374,N_1965,N_1934);
and U2375 (N_2375,N_1838,N_1801);
or U2376 (N_2376,N_1863,N_1785);
and U2377 (N_2377,N_1993,N_1872);
xor U2378 (N_2378,N_1771,N_1846);
or U2379 (N_2379,N_1606,N_1816);
nor U2380 (N_2380,N_1682,N_1879);
xor U2381 (N_2381,N_1710,N_1614);
nand U2382 (N_2382,N_1686,N_1715);
nor U2383 (N_2383,N_1640,N_1976);
nor U2384 (N_2384,N_1989,N_1894);
nor U2385 (N_2385,N_1871,N_1726);
xor U2386 (N_2386,N_1632,N_1685);
or U2387 (N_2387,N_1799,N_1980);
xnor U2388 (N_2388,N_1682,N_1841);
or U2389 (N_2389,N_1648,N_1692);
and U2390 (N_2390,N_1850,N_1718);
or U2391 (N_2391,N_1761,N_1997);
nor U2392 (N_2392,N_1775,N_1688);
or U2393 (N_2393,N_1927,N_1828);
nor U2394 (N_2394,N_1701,N_1611);
xor U2395 (N_2395,N_1929,N_1699);
and U2396 (N_2396,N_1653,N_1944);
or U2397 (N_2397,N_1917,N_1632);
or U2398 (N_2398,N_1737,N_1608);
or U2399 (N_2399,N_1725,N_1665);
and U2400 (N_2400,N_2300,N_2095);
xnor U2401 (N_2401,N_2206,N_2200);
nand U2402 (N_2402,N_2335,N_2060);
and U2403 (N_2403,N_2086,N_2058);
nor U2404 (N_2404,N_2395,N_2314);
or U2405 (N_2405,N_2178,N_2032);
xor U2406 (N_2406,N_2091,N_2366);
nand U2407 (N_2407,N_2145,N_2329);
or U2408 (N_2408,N_2350,N_2320);
xnor U2409 (N_2409,N_2168,N_2182);
nand U2410 (N_2410,N_2349,N_2049);
nand U2411 (N_2411,N_2284,N_2343);
or U2412 (N_2412,N_2215,N_2194);
or U2413 (N_2413,N_2275,N_2212);
nor U2414 (N_2414,N_2204,N_2156);
nand U2415 (N_2415,N_2279,N_2238);
or U2416 (N_2416,N_2175,N_2179);
nor U2417 (N_2417,N_2181,N_2353);
and U2418 (N_2418,N_2149,N_2323);
or U2419 (N_2419,N_2365,N_2102);
xnor U2420 (N_2420,N_2271,N_2030);
xor U2421 (N_2421,N_2332,N_2360);
nor U2422 (N_2422,N_2059,N_2305);
and U2423 (N_2423,N_2199,N_2042);
and U2424 (N_2424,N_2210,N_2381);
and U2425 (N_2425,N_2027,N_2240);
xnor U2426 (N_2426,N_2039,N_2174);
nand U2427 (N_2427,N_2347,N_2070);
xnor U2428 (N_2428,N_2148,N_2159);
nor U2429 (N_2429,N_2304,N_2112);
and U2430 (N_2430,N_2376,N_2163);
nand U2431 (N_2431,N_2348,N_2139);
or U2432 (N_2432,N_2268,N_2031);
xor U2433 (N_2433,N_2235,N_2056);
and U2434 (N_2434,N_2161,N_2385);
xor U2435 (N_2435,N_2114,N_2044);
nor U2436 (N_2436,N_2016,N_2263);
nor U2437 (N_2437,N_2355,N_2183);
and U2438 (N_2438,N_2080,N_2184);
nand U2439 (N_2439,N_2101,N_2333);
xnor U2440 (N_2440,N_2371,N_2264);
nor U2441 (N_2441,N_2144,N_2386);
and U2442 (N_2442,N_2007,N_2189);
xor U2443 (N_2443,N_2010,N_2265);
nor U2444 (N_2444,N_2171,N_2246);
nor U2445 (N_2445,N_2379,N_2047);
or U2446 (N_2446,N_2363,N_2219);
or U2447 (N_2447,N_2104,N_2025);
xor U2448 (N_2448,N_2142,N_2046);
nand U2449 (N_2449,N_2336,N_2354);
and U2450 (N_2450,N_2261,N_2085);
and U2451 (N_2451,N_2321,N_2307);
xnor U2452 (N_2452,N_2232,N_2244);
and U2453 (N_2453,N_2170,N_2327);
nand U2454 (N_2454,N_2002,N_2029);
nand U2455 (N_2455,N_2198,N_2176);
and U2456 (N_2456,N_2055,N_2223);
and U2457 (N_2457,N_2021,N_2151);
nand U2458 (N_2458,N_2356,N_2377);
nor U2459 (N_2459,N_2153,N_2328);
and U2460 (N_2460,N_2285,N_2064);
nand U2461 (N_2461,N_2172,N_2270);
and U2462 (N_2462,N_2069,N_2276);
or U2463 (N_2463,N_2146,N_2015);
nor U2464 (N_2464,N_2083,N_2193);
nor U2465 (N_2465,N_2001,N_2211);
and U2466 (N_2466,N_2259,N_2107);
nand U2467 (N_2467,N_2318,N_2378);
and U2468 (N_2468,N_2008,N_2322);
or U2469 (N_2469,N_2130,N_2018);
nand U2470 (N_2470,N_2037,N_2158);
xnor U2471 (N_2471,N_2117,N_2187);
nand U2472 (N_2472,N_2242,N_2196);
nand U2473 (N_2473,N_2294,N_2207);
or U2474 (N_2474,N_2118,N_2399);
nor U2475 (N_2475,N_2397,N_2387);
nand U2476 (N_2476,N_2293,N_2043);
and U2477 (N_2477,N_2124,N_2197);
nand U2478 (N_2478,N_2132,N_2071);
xnor U2479 (N_2479,N_2267,N_2133);
and U2480 (N_2480,N_2334,N_2023);
or U2481 (N_2481,N_2262,N_2088);
nand U2482 (N_2482,N_2359,N_2241);
or U2483 (N_2483,N_2020,N_2109);
and U2484 (N_2484,N_2251,N_2165);
nor U2485 (N_2485,N_2269,N_2077);
nor U2486 (N_2486,N_2121,N_2105);
nand U2487 (N_2487,N_2250,N_2066);
or U2488 (N_2488,N_2249,N_2330);
nand U2489 (N_2489,N_2167,N_2160);
xnor U2490 (N_2490,N_2134,N_2177);
or U2491 (N_2491,N_2218,N_2191);
nor U2492 (N_2492,N_2340,N_2203);
xor U2493 (N_2493,N_2384,N_2110);
and U2494 (N_2494,N_2103,N_2051);
nor U2495 (N_2495,N_2122,N_2342);
or U2496 (N_2496,N_2052,N_2111);
xor U2497 (N_2497,N_2119,N_2065);
xnor U2498 (N_2498,N_2048,N_2033);
nor U2499 (N_2499,N_2396,N_2392);
and U2500 (N_2500,N_2050,N_2147);
or U2501 (N_2501,N_2097,N_2005);
and U2502 (N_2502,N_2014,N_2099);
or U2503 (N_2503,N_2310,N_2131);
nand U2504 (N_2504,N_2315,N_2312);
nand U2505 (N_2505,N_2282,N_2098);
and U2506 (N_2506,N_2063,N_2388);
nor U2507 (N_2507,N_2129,N_2141);
and U2508 (N_2508,N_2361,N_2108);
and U2509 (N_2509,N_2185,N_2054);
nor U2510 (N_2510,N_2120,N_2209);
xnor U2511 (N_2511,N_2036,N_2180);
or U2512 (N_2512,N_2389,N_2061);
or U2513 (N_2513,N_2226,N_2319);
or U2514 (N_2514,N_2192,N_2345);
xnor U2515 (N_2515,N_2123,N_2143);
nand U2516 (N_2516,N_2011,N_2306);
or U2517 (N_2517,N_2201,N_2140);
nand U2518 (N_2518,N_2081,N_2228);
xnor U2519 (N_2519,N_2311,N_2162);
xnor U2520 (N_2520,N_2222,N_2325);
and U2521 (N_2521,N_2324,N_2257);
or U2522 (N_2522,N_2231,N_2357);
nor U2523 (N_2523,N_2213,N_2073);
xnor U2524 (N_2524,N_2346,N_2034);
nor U2525 (N_2525,N_2173,N_2372);
and U2526 (N_2526,N_2224,N_2000);
or U2527 (N_2527,N_2094,N_2035);
nor U2528 (N_2528,N_2188,N_2286);
and U2529 (N_2529,N_2038,N_2338);
nand U2530 (N_2530,N_2138,N_2126);
and U2531 (N_2531,N_2398,N_2079);
xor U2532 (N_2532,N_2277,N_2026);
xnor U2533 (N_2533,N_2009,N_2078);
nand U2534 (N_2534,N_2362,N_2100);
and U2535 (N_2535,N_2006,N_2341);
or U2536 (N_2536,N_2195,N_2316);
nand U2537 (N_2537,N_2374,N_2237);
and U2538 (N_2538,N_2125,N_2243);
and U2539 (N_2539,N_2280,N_2288);
nand U2540 (N_2540,N_2290,N_2115);
and U2541 (N_2541,N_2164,N_2375);
nor U2542 (N_2542,N_2239,N_2067);
nor U2543 (N_2543,N_2383,N_2352);
nand U2544 (N_2544,N_2296,N_2373);
nand U2545 (N_2545,N_2295,N_2155);
nand U2546 (N_2546,N_2041,N_2152);
nor U2547 (N_2547,N_2202,N_2394);
and U2548 (N_2548,N_2260,N_2245);
nand U2549 (N_2549,N_2057,N_2278);
or U2550 (N_2550,N_2358,N_2116);
and U2551 (N_2551,N_2072,N_2283);
nor U2552 (N_2552,N_2331,N_2012);
nor U2553 (N_2553,N_2106,N_2344);
nor U2554 (N_2554,N_2028,N_2302);
and U2555 (N_2555,N_2214,N_2281);
or U2556 (N_2556,N_2113,N_2254);
or U2557 (N_2557,N_2393,N_2253);
xor U2558 (N_2558,N_2364,N_2370);
nand U2559 (N_2559,N_2013,N_2003);
xor U2560 (N_2560,N_2225,N_2084);
nor U2561 (N_2561,N_2157,N_2258);
xnor U2562 (N_2562,N_2289,N_2220);
nand U2563 (N_2563,N_2303,N_2248);
nand U2564 (N_2564,N_2136,N_2298);
or U2565 (N_2565,N_2390,N_2208);
xnor U2566 (N_2566,N_2292,N_2040);
nor U2567 (N_2567,N_2150,N_2093);
nand U2568 (N_2568,N_2089,N_2272);
nand U2569 (N_2569,N_2380,N_2154);
and U2570 (N_2570,N_2221,N_2337);
xnor U2571 (N_2571,N_2339,N_2287);
nand U2572 (N_2572,N_2266,N_2247);
nor U2573 (N_2573,N_2062,N_2082);
and U2574 (N_2574,N_2368,N_2309);
or U2575 (N_2575,N_2127,N_2186);
nor U2576 (N_2576,N_2190,N_2166);
xor U2577 (N_2577,N_2128,N_2205);
xnor U2578 (N_2578,N_2255,N_2299);
and U2579 (N_2579,N_2137,N_2024);
nand U2580 (N_2580,N_2087,N_2092);
nand U2581 (N_2581,N_2053,N_2068);
nand U2582 (N_2582,N_2216,N_2297);
or U2583 (N_2583,N_2004,N_2022);
or U2584 (N_2584,N_2169,N_2090);
or U2585 (N_2585,N_2317,N_2308);
nand U2586 (N_2586,N_2234,N_2301);
nand U2587 (N_2587,N_2230,N_2274);
nand U2588 (N_2588,N_2096,N_2229);
xor U2589 (N_2589,N_2017,N_2291);
or U2590 (N_2590,N_2391,N_2019);
nand U2591 (N_2591,N_2045,N_2217);
or U2592 (N_2592,N_2326,N_2256);
xor U2593 (N_2593,N_2227,N_2382);
or U2594 (N_2594,N_2313,N_2076);
or U2595 (N_2595,N_2074,N_2252);
and U2596 (N_2596,N_2369,N_2236);
nand U2597 (N_2597,N_2351,N_2135);
nor U2598 (N_2598,N_2273,N_2367);
nand U2599 (N_2599,N_2233,N_2075);
and U2600 (N_2600,N_2213,N_2312);
nor U2601 (N_2601,N_2332,N_2068);
xor U2602 (N_2602,N_2370,N_2119);
nand U2603 (N_2603,N_2394,N_2052);
and U2604 (N_2604,N_2089,N_2111);
xnor U2605 (N_2605,N_2056,N_2033);
or U2606 (N_2606,N_2350,N_2306);
nand U2607 (N_2607,N_2380,N_2275);
xnor U2608 (N_2608,N_2319,N_2169);
and U2609 (N_2609,N_2133,N_2110);
and U2610 (N_2610,N_2198,N_2233);
nor U2611 (N_2611,N_2129,N_2025);
nor U2612 (N_2612,N_2084,N_2141);
and U2613 (N_2613,N_2118,N_2036);
nor U2614 (N_2614,N_2139,N_2174);
nand U2615 (N_2615,N_2305,N_2295);
xnor U2616 (N_2616,N_2266,N_2012);
nor U2617 (N_2617,N_2019,N_2288);
nor U2618 (N_2618,N_2002,N_2246);
xor U2619 (N_2619,N_2074,N_2010);
xor U2620 (N_2620,N_2205,N_2035);
and U2621 (N_2621,N_2187,N_2158);
nor U2622 (N_2622,N_2253,N_2215);
xnor U2623 (N_2623,N_2225,N_2331);
xnor U2624 (N_2624,N_2349,N_2034);
or U2625 (N_2625,N_2336,N_2086);
nor U2626 (N_2626,N_2073,N_2088);
xnor U2627 (N_2627,N_2080,N_2279);
xor U2628 (N_2628,N_2175,N_2061);
nor U2629 (N_2629,N_2384,N_2378);
xnor U2630 (N_2630,N_2228,N_2243);
xnor U2631 (N_2631,N_2206,N_2099);
xor U2632 (N_2632,N_2201,N_2172);
nand U2633 (N_2633,N_2054,N_2288);
or U2634 (N_2634,N_2250,N_2084);
and U2635 (N_2635,N_2317,N_2306);
and U2636 (N_2636,N_2289,N_2184);
nand U2637 (N_2637,N_2223,N_2054);
and U2638 (N_2638,N_2397,N_2174);
and U2639 (N_2639,N_2148,N_2033);
and U2640 (N_2640,N_2211,N_2380);
nor U2641 (N_2641,N_2262,N_2282);
and U2642 (N_2642,N_2253,N_2352);
nor U2643 (N_2643,N_2042,N_2020);
nor U2644 (N_2644,N_2215,N_2237);
nor U2645 (N_2645,N_2145,N_2030);
and U2646 (N_2646,N_2313,N_2110);
nand U2647 (N_2647,N_2073,N_2117);
or U2648 (N_2648,N_2158,N_2000);
nand U2649 (N_2649,N_2379,N_2385);
and U2650 (N_2650,N_2094,N_2004);
nor U2651 (N_2651,N_2272,N_2156);
and U2652 (N_2652,N_2259,N_2308);
or U2653 (N_2653,N_2245,N_2052);
or U2654 (N_2654,N_2067,N_2131);
and U2655 (N_2655,N_2147,N_2207);
xor U2656 (N_2656,N_2079,N_2326);
nand U2657 (N_2657,N_2189,N_2330);
nand U2658 (N_2658,N_2332,N_2361);
nor U2659 (N_2659,N_2042,N_2237);
nor U2660 (N_2660,N_2240,N_2278);
nor U2661 (N_2661,N_2224,N_2329);
and U2662 (N_2662,N_2124,N_2070);
nand U2663 (N_2663,N_2010,N_2055);
xor U2664 (N_2664,N_2148,N_2031);
xor U2665 (N_2665,N_2164,N_2351);
and U2666 (N_2666,N_2175,N_2260);
and U2667 (N_2667,N_2124,N_2046);
xnor U2668 (N_2668,N_2181,N_2109);
or U2669 (N_2669,N_2021,N_2351);
nor U2670 (N_2670,N_2288,N_2244);
or U2671 (N_2671,N_2354,N_2351);
nor U2672 (N_2672,N_2327,N_2188);
and U2673 (N_2673,N_2286,N_2019);
nor U2674 (N_2674,N_2041,N_2369);
xnor U2675 (N_2675,N_2372,N_2385);
xor U2676 (N_2676,N_2040,N_2290);
nor U2677 (N_2677,N_2379,N_2363);
and U2678 (N_2678,N_2144,N_2112);
or U2679 (N_2679,N_2023,N_2097);
nand U2680 (N_2680,N_2178,N_2245);
nand U2681 (N_2681,N_2211,N_2372);
or U2682 (N_2682,N_2093,N_2354);
nor U2683 (N_2683,N_2378,N_2008);
xor U2684 (N_2684,N_2142,N_2334);
nand U2685 (N_2685,N_2357,N_2334);
nor U2686 (N_2686,N_2280,N_2325);
xor U2687 (N_2687,N_2393,N_2155);
and U2688 (N_2688,N_2159,N_2039);
xor U2689 (N_2689,N_2372,N_2075);
or U2690 (N_2690,N_2266,N_2287);
nor U2691 (N_2691,N_2057,N_2075);
nor U2692 (N_2692,N_2377,N_2242);
xnor U2693 (N_2693,N_2036,N_2100);
and U2694 (N_2694,N_2302,N_2257);
nor U2695 (N_2695,N_2148,N_2267);
xor U2696 (N_2696,N_2017,N_2387);
and U2697 (N_2697,N_2233,N_2076);
xnor U2698 (N_2698,N_2165,N_2309);
or U2699 (N_2699,N_2092,N_2016);
or U2700 (N_2700,N_2336,N_2153);
and U2701 (N_2701,N_2038,N_2287);
nand U2702 (N_2702,N_2376,N_2267);
and U2703 (N_2703,N_2337,N_2354);
xor U2704 (N_2704,N_2274,N_2018);
xor U2705 (N_2705,N_2227,N_2219);
xnor U2706 (N_2706,N_2123,N_2072);
xnor U2707 (N_2707,N_2146,N_2032);
nand U2708 (N_2708,N_2138,N_2211);
nand U2709 (N_2709,N_2007,N_2067);
xor U2710 (N_2710,N_2024,N_2138);
nand U2711 (N_2711,N_2082,N_2163);
xnor U2712 (N_2712,N_2394,N_2390);
and U2713 (N_2713,N_2266,N_2141);
nand U2714 (N_2714,N_2345,N_2171);
nor U2715 (N_2715,N_2239,N_2362);
nand U2716 (N_2716,N_2398,N_2259);
and U2717 (N_2717,N_2156,N_2320);
nand U2718 (N_2718,N_2080,N_2240);
xor U2719 (N_2719,N_2284,N_2017);
nand U2720 (N_2720,N_2123,N_2057);
and U2721 (N_2721,N_2026,N_2355);
and U2722 (N_2722,N_2221,N_2300);
and U2723 (N_2723,N_2194,N_2328);
and U2724 (N_2724,N_2267,N_2310);
xor U2725 (N_2725,N_2201,N_2156);
nand U2726 (N_2726,N_2258,N_2142);
nand U2727 (N_2727,N_2312,N_2078);
nand U2728 (N_2728,N_2023,N_2117);
or U2729 (N_2729,N_2206,N_2109);
nand U2730 (N_2730,N_2216,N_2002);
nor U2731 (N_2731,N_2089,N_2266);
or U2732 (N_2732,N_2295,N_2136);
xor U2733 (N_2733,N_2373,N_2232);
or U2734 (N_2734,N_2021,N_2341);
nor U2735 (N_2735,N_2190,N_2374);
nor U2736 (N_2736,N_2236,N_2384);
xnor U2737 (N_2737,N_2064,N_2381);
or U2738 (N_2738,N_2321,N_2275);
xnor U2739 (N_2739,N_2214,N_2034);
xnor U2740 (N_2740,N_2376,N_2055);
nor U2741 (N_2741,N_2217,N_2158);
and U2742 (N_2742,N_2060,N_2358);
xor U2743 (N_2743,N_2291,N_2268);
xor U2744 (N_2744,N_2275,N_2335);
nor U2745 (N_2745,N_2225,N_2074);
and U2746 (N_2746,N_2249,N_2298);
or U2747 (N_2747,N_2362,N_2399);
xnor U2748 (N_2748,N_2212,N_2358);
or U2749 (N_2749,N_2070,N_2325);
nor U2750 (N_2750,N_2052,N_2008);
nand U2751 (N_2751,N_2283,N_2013);
or U2752 (N_2752,N_2137,N_2103);
and U2753 (N_2753,N_2050,N_2224);
nand U2754 (N_2754,N_2121,N_2259);
and U2755 (N_2755,N_2094,N_2055);
nand U2756 (N_2756,N_2187,N_2150);
and U2757 (N_2757,N_2045,N_2152);
or U2758 (N_2758,N_2149,N_2244);
nor U2759 (N_2759,N_2002,N_2237);
xnor U2760 (N_2760,N_2211,N_2266);
and U2761 (N_2761,N_2074,N_2196);
or U2762 (N_2762,N_2039,N_2007);
or U2763 (N_2763,N_2110,N_2243);
nor U2764 (N_2764,N_2261,N_2200);
and U2765 (N_2765,N_2358,N_2354);
nor U2766 (N_2766,N_2286,N_2251);
nor U2767 (N_2767,N_2236,N_2074);
nor U2768 (N_2768,N_2348,N_2239);
nor U2769 (N_2769,N_2175,N_2170);
xor U2770 (N_2770,N_2391,N_2152);
and U2771 (N_2771,N_2109,N_2255);
and U2772 (N_2772,N_2147,N_2307);
nor U2773 (N_2773,N_2113,N_2109);
nor U2774 (N_2774,N_2196,N_2149);
and U2775 (N_2775,N_2163,N_2320);
or U2776 (N_2776,N_2229,N_2387);
or U2777 (N_2777,N_2310,N_2189);
nand U2778 (N_2778,N_2253,N_2017);
nor U2779 (N_2779,N_2075,N_2078);
or U2780 (N_2780,N_2256,N_2305);
xnor U2781 (N_2781,N_2109,N_2002);
and U2782 (N_2782,N_2108,N_2257);
and U2783 (N_2783,N_2387,N_2378);
and U2784 (N_2784,N_2022,N_2275);
xor U2785 (N_2785,N_2256,N_2128);
and U2786 (N_2786,N_2042,N_2027);
or U2787 (N_2787,N_2140,N_2224);
nor U2788 (N_2788,N_2278,N_2191);
or U2789 (N_2789,N_2197,N_2233);
nor U2790 (N_2790,N_2005,N_2192);
nor U2791 (N_2791,N_2201,N_2049);
nand U2792 (N_2792,N_2091,N_2174);
or U2793 (N_2793,N_2347,N_2290);
xor U2794 (N_2794,N_2058,N_2037);
xnor U2795 (N_2795,N_2101,N_2121);
xor U2796 (N_2796,N_2269,N_2170);
nor U2797 (N_2797,N_2255,N_2231);
nor U2798 (N_2798,N_2208,N_2321);
nand U2799 (N_2799,N_2010,N_2232);
and U2800 (N_2800,N_2448,N_2549);
xnor U2801 (N_2801,N_2669,N_2670);
and U2802 (N_2802,N_2445,N_2744);
nand U2803 (N_2803,N_2601,N_2593);
xnor U2804 (N_2804,N_2679,N_2544);
xnor U2805 (N_2805,N_2492,N_2529);
and U2806 (N_2806,N_2729,N_2757);
and U2807 (N_2807,N_2415,N_2466);
and U2808 (N_2808,N_2478,N_2768);
nand U2809 (N_2809,N_2701,N_2759);
nand U2810 (N_2810,N_2778,N_2659);
or U2811 (N_2811,N_2600,N_2416);
nand U2812 (N_2812,N_2766,N_2428);
nor U2813 (N_2813,N_2716,N_2740);
and U2814 (N_2814,N_2675,N_2621);
nand U2815 (N_2815,N_2489,N_2450);
and U2816 (N_2816,N_2686,N_2779);
nand U2817 (N_2817,N_2585,N_2646);
and U2818 (N_2818,N_2524,N_2725);
and U2819 (N_2819,N_2718,N_2470);
or U2820 (N_2820,N_2697,N_2534);
and U2821 (N_2821,N_2571,N_2685);
nor U2822 (N_2822,N_2695,N_2795);
nand U2823 (N_2823,N_2407,N_2682);
nand U2824 (N_2824,N_2707,N_2656);
and U2825 (N_2825,N_2561,N_2565);
xnor U2826 (N_2826,N_2581,N_2611);
nor U2827 (N_2827,N_2752,N_2566);
nor U2828 (N_2828,N_2727,N_2617);
or U2829 (N_2829,N_2780,N_2404);
xor U2830 (N_2830,N_2429,N_2750);
nor U2831 (N_2831,N_2641,N_2764);
or U2832 (N_2832,N_2777,N_2487);
and U2833 (N_2833,N_2755,N_2511);
or U2834 (N_2834,N_2642,N_2664);
xnor U2835 (N_2835,N_2484,N_2710);
or U2836 (N_2836,N_2523,N_2420);
xor U2837 (N_2837,N_2556,N_2770);
nand U2838 (N_2838,N_2479,N_2721);
or U2839 (N_2839,N_2475,N_2781);
xnor U2840 (N_2840,N_2403,N_2618);
nand U2841 (N_2841,N_2596,N_2735);
or U2842 (N_2842,N_2666,N_2599);
nor U2843 (N_2843,N_2513,N_2771);
nand U2844 (N_2844,N_2486,N_2602);
nor U2845 (N_2845,N_2567,N_2594);
nor U2846 (N_2846,N_2606,N_2713);
and U2847 (N_2847,N_2432,N_2538);
nor U2848 (N_2848,N_2765,N_2608);
or U2849 (N_2849,N_2461,N_2418);
nand U2850 (N_2850,N_2742,N_2442);
nor U2851 (N_2851,N_2712,N_2510);
or U2852 (N_2852,N_2463,N_2604);
xnor U2853 (N_2853,N_2465,N_2541);
or U2854 (N_2854,N_2493,N_2748);
and U2855 (N_2855,N_2451,N_2532);
nand U2856 (N_2856,N_2681,N_2661);
nor U2857 (N_2857,N_2494,N_2434);
and U2858 (N_2858,N_2413,N_2526);
and U2859 (N_2859,N_2546,N_2405);
nand U2860 (N_2860,N_2414,N_2772);
nor U2861 (N_2861,N_2690,N_2460);
nor U2862 (N_2862,N_2654,N_2512);
and U2863 (N_2863,N_2563,N_2663);
nand U2864 (N_2864,N_2425,N_2570);
nand U2865 (N_2865,N_2427,N_2540);
nand U2866 (N_2866,N_2467,N_2530);
xnor U2867 (N_2867,N_2422,N_2635);
xnor U2868 (N_2868,N_2706,N_2788);
xor U2869 (N_2869,N_2495,N_2631);
and U2870 (N_2870,N_2753,N_2717);
or U2871 (N_2871,N_2746,N_2726);
or U2872 (N_2872,N_2651,N_2782);
xor U2873 (N_2873,N_2569,N_2722);
nand U2874 (N_2874,N_2678,N_2609);
nand U2875 (N_2875,N_2630,N_2649);
and U2876 (N_2876,N_2481,N_2503);
xnor U2877 (N_2877,N_2736,N_2688);
or U2878 (N_2878,N_2591,N_2568);
and U2879 (N_2879,N_2551,N_2446);
nand U2880 (N_2880,N_2714,N_2547);
nand U2881 (N_2881,N_2756,N_2402);
and U2882 (N_2882,N_2444,N_2424);
or U2883 (N_2883,N_2514,N_2471);
nor U2884 (N_2884,N_2528,N_2576);
xor U2885 (N_2885,N_2455,N_2555);
and U2886 (N_2886,N_2474,N_2454);
and U2887 (N_2887,N_2578,N_2462);
or U2888 (N_2888,N_2623,N_2767);
nand U2889 (N_2889,N_2728,N_2739);
and U2890 (N_2890,N_2655,N_2419);
xor U2891 (N_2891,N_2439,N_2527);
nor U2892 (N_2892,N_2790,N_2586);
and U2893 (N_2893,N_2411,N_2457);
nand U2894 (N_2894,N_2580,N_2592);
or U2895 (N_2895,N_2558,N_2639);
xor U2896 (N_2896,N_2708,N_2662);
nand U2897 (N_2897,N_2562,N_2693);
or U2898 (N_2898,N_2734,N_2644);
xor U2899 (N_2899,N_2436,N_2437);
and U2900 (N_2900,N_2412,N_2543);
and U2901 (N_2901,N_2583,N_2498);
and U2902 (N_2902,N_2535,N_2438);
xor U2903 (N_2903,N_2637,N_2521);
xnor U2904 (N_2904,N_2776,N_2645);
and U2905 (N_2905,N_2536,N_2473);
nor U2906 (N_2906,N_2579,N_2539);
and U2907 (N_2907,N_2783,N_2762);
nor U2908 (N_2908,N_2440,N_2650);
nor U2909 (N_2909,N_2560,N_2658);
or U2910 (N_2910,N_2632,N_2501);
nor U2911 (N_2911,N_2469,N_2441);
xnor U2912 (N_2912,N_2497,N_2763);
and U2913 (N_2913,N_2785,N_2667);
xor U2914 (N_2914,N_2731,N_2557);
and U2915 (N_2915,N_2577,N_2515);
or U2916 (N_2916,N_2542,N_2499);
and U2917 (N_2917,N_2452,N_2468);
nor U2918 (N_2918,N_2786,N_2505);
xor U2919 (N_2919,N_2629,N_2423);
nand U2920 (N_2920,N_2737,N_2624);
nand U2921 (N_2921,N_2491,N_2531);
or U2922 (N_2922,N_2643,N_2680);
xor U2923 (N_2923,N_2789,N_2724);
nand U2924 (N_2924,N_2622,N_2673);
and U2925 (N_2925,N_2456,N_2715);
nor U2926 (N_2926,N_2464,N_2598);
nand U2927 (N_2927,N_2657,N_2545);
xnor U2928 (N_2928,N_2709,N_2426);
xnor U2929 (N_2929,N_2733,N_2496);
nor U2930 (N_2930,N_2677,N_2694);
and U2931 (N_2931,N_2537,N_2751);
nand U2932 (N_2932,N_2435,N_2612);
xor U2933 (N_2933,N_2689,N_2408);
and U2934 (N_2934,N_2758,N_2640);
and U2935 (N_2935,N_2747,N_2406);
nor U2936 (N_2936,N_2760,N_2738);
or U2937 (N_2937,N_2485,N_2614);
and U2938 (N_2938,N_2589,N_2626);
xnor U2939 (N_2939,N_2732,N_2647);
nand U2940 (N_2940,N_2449,N_2787);
and U2941 (N_2941,N_2648,N_2684);
and U2942 (N_2942,N_2665,N_2443);
xnor U2943 (N_2943,N_2769,N_2720);
and U2944 (N_2944,N_2794,N_2401);
and U2945 (N_2945,N_2638,N_2683);
nand U2946 (N_2946,N_2796,N_2517);
nand U2947 (N_2947,N_2605,N_2610);
or U2948 (N_2948,N_2433,N_2775);
and U2949 (N_2949,N_2552,N_2711);
or U2950 (N_2950,N_2588,N_2516);
nor U2951 (N_2951,N_2702,N_2421);
nor U2952 (N_2952,N_2525,N_2410);
and U2953 (N_2953,N_2483,N_2573);
nand U2954 (N_2954,N_2575,N_2730);
xnor U2955 (N_2955,N_2533,N_2507);
and U2956 (N_2956,N_2792,N_2799);
and U2957 (N_2957,N_2672,N_2550);
xnor U2958 (N_2958,N_2797,N_2453);
xnor U2959 (N_2959,N_2636,N_2696);
xnor U2960 (N_2960,N_2773,N_2480);
and U2961 (N_2961,N_2628,N_2504);
nand U2962 (N_2962,N_2502,N_2459);
nor U2963 (N_2963,N_2687,N_2477);
and U2964 (N_2964,N_2447,N_2625);
and U2965 (N_2965,N_2572,N_2653);
and U2966 (N_2966,N_2703,N_2400);
and U2967 (N_2967,N_2472,N_2409);
or U2968 (N_2968,N_2698,N_2509);
and U2969 (N_2969,N_2616,N_2520);
nor U2970 (N_2970,N_2613,N_2692);
and U2971 (N_2971,N_2798,N_2761);
nand U2972 (N_2972,N_2417,N_2634);
nand U2973 (N_2973,N_2518,N_2582);
nand U2974 (N_2974,N_2488,N_2482);
nand U2975 (N_2975,N_2793,N_2741);
nand U2976 (N_2976,N_2676,N_2522);
nor U2977 (N_2977,N_2705,N_2619);
xnor U2978 (N_2978,N_2704,N_2548);
nor U2979 (N_2979,N_2691,N_2674);
nor U2980 (N_2980,N_2458,N_2745);
nand U2981 (N_2981,N_2723,N_2564);
xnor U2982 (N_2982,N_2791,N_2506);
xnor U2983 (N_2983,N_2633,N_2607);
nor U2984 (N_2984,N_2500,N_2587);
xor U2985 (N_2985,N_2652,N_2671);
or U2986 (N_2986,N_2699,N_2584);
nor U2987 (N_2987,N_2660,N_2519);
xor U2988 (N_2988,N_2597,N_2700);
nor U2989 (N_2989,N_2620,N_2743);
and U2990 (N_2990,N_2749,N_2603);
nand U2991 (N_2991,N_2754,N_2719);
or U2992 (N_2992,N_2430,N_2574);
nand U2993 (N_2993,N_2784,N_2774);
nor U2994 (N_2994,N_2595,N_2553);
xor U2995 (N_2995,N_2668,N_2559);
nor U2996 (N_2996,N_2615,N_2627);
xnor U2997 (N_2997,N_2508,N_2431);
and U2998 (N_2998,N_2554,N_2590);
or U2999 (N_2999,N_2490,N_2476);
xor U3000 (N_3000,N_2642,N_2554);
or U3001 (N_3001,N_2470,N_2417);
nor U3002 (N_3002,N_2734,N_2643);
xnor U3003 (N_3003,N_2579,N_2440);
nand U3004 (N_3004,N_2441,N_2572);
nand U3005 (N_3005,N_2685,N_2744);
and U3006 (N_3006,N_2636,N_2562);
xnor U3007 (N_3007,N_2627,N_2634);
xor U3008 (N_3008,N_2584,N_2622);
nand U3009 (N_3009,N_2504,N_2559);
or U3010 (N_3010,N_2666,N_2474);
nand U3011 (N_3011,N_2623,N_2667);
nand U3012 (N_3012,N_2697,N_2430);
and U3013 (N_3013,N_2666,N_2772);
xnor U3014 (N_3014,N_2528,N_2545);
or U3015 (N_3015,N_2585,N_2796);
nor U3016 (N_3016,N_2794,N_2767);
nand U3017 (N_3017,N_2697,N_2498);
nand U3018 (N_3018,N_2470,N_2484);
and U3019 (N_3019,N_2447,N_2743);
xnor U3020 (N_3020,N_2446,N_2532);
nand U3021 (N_3021,N_2514,N_2627);
nor U3022 (N_3022,N_2600,N_2509);
nor U3023 (N_3023,N_2417,N_2452);
and U3024 (N_3024,N_2402,N_2608);
and U3025 (N_3025,N_2669,N_2514);
nor U3026 (N_3026,N_2551,N_2792);
or U3027 (N_3027,N_2417,N_2675);
nand U3028 (N_3028,N_2790,N_2647);
or U3029 (N_3029,N_2424,N_2749);
and U3030 (N_3030,N_2726,N_2531);
and U3031 (N_3031,N_2787,N_2580);
and U3032 (N_3032,N_2781,N_2635);
or U3033 (N_3033,N_2723,N_2660);
or U3034 (N_3034,N_2495,N_2665);
nor U3035 (N_3035,N_2492,N_2512);
and U3036 (N_3036,N_2514,N_2567);
xor U3037 (N_3037,N_2679,N_2686);
nand U3038 (N_3038,N_2660,N_2569);
nor U3039 (N_3039,N_2687,N_2533);
nand U3040 (N_3040,N_2733,N_2661);
xor U3041 (N_3041,N_2528,N_2718);
nor U3042 (N_3042,N_2457,N_2732);
nor U3043 (N_3043,N_2723,N_2535);
xor U3044 (N_3044,N_2566,N_2678);
nand U3045 (N_3045,N_2419,N_2456);
nor U3046 (N_3046,N_2630,N_2769);
nand U3047 (N_3047,N_2402,N_2420);
or U3048 (N_3048,N_2723,N_2604);
xor U3049 (N_3049,N_2571,N_2548);
nand U3050 (N_3050,N_2502,N_2453);
or U3051 (N_3051,N_2568,N_2742);
or U3052 (N_3052,N_2752,N_2648);
or U3053 (N_3053,N_2583,N_2631);
nor U3054 (N_3054,N_2514,N_2647);
and U3055 (N_3055,N_2564,N_2523);
and U3056 (N_3056,N_2684,N_2528);
nand U3057 (N_3057,N_2667,N_2714);
or U3058 (N_3058,N_2605,N_2635);
or U3059 (N_3059,N_2584,N_2511);
nor U3060 (N_3060,N_2656,N_2786);
xor U3061 (N_3061,N_2784,N_2649);
or U3062 (N_3062,N_2476,N_2573);
or U3063 (N_3063,N_2785,N_2481);
nor U3064 (N_3064,N_2665,N_2605);
nor U3065 (N_3065,N_2628,N_2527);
xor U3066 (N_3066,N_2506,N_2464);
nand U3067 (N_3067,N_2433,N_2643);
nand U3068 (N_3068,N_2724,N_2494);
xnor U3069 (N_3069,N_2526,N_2650);
nand U3070 (N_3070,N_2412,N_2440);
or U3071 (N_3071,N_2521,N_2732);
nand U3072 (N_3072,N_2597,N_2601);
xor U3073 (N_3073,N_2567,N_2408);
nor U3074 (N_3074,N_2723,N_2587);
and U3075 (N_3075,N_2676,N_2488);
xnor U3076 (N_3076,N_2484,N_2444);
nor U3077 (N_3077,N_2609,N_2665);
nor U3078 (N_3078,N_2541,N_2568);
nand U3079 (N_3079,N_2453,N_2628);
and U3080 (N_3080,N_2495,N_2796);
and U3081 (N_3081,N_2741,N_2644);
nor U3082 (N_3082,N_2489,N_2431);
nand U3083 (N_3083,N_2507,N_2489);
and U3084 (N_3084,N_2413,N_2664);
or U3085 (N_3085,N_2585,N_2560);
and U3086 (N_3086,N_2708,N_2765);
or U3087 (N_3087,N_2771,N_2403);
and U3088 (N_3088,N_2733,N_2764);
nor U3089 (N_3089,N_2738,N_2538);
nor U3090 (N_3090,N_2441,N_2750);
nor U3091 (N_3091,N_2520,N_2416);
or U3092 (N_3092,N_2607,N_2576);
and U3093 (N_3093,N_2794,N_2554);
nand U3094 (N_3094,N_2502,N_2452);
nor U3095 (N_3095,N_2705,N_2573);
and U3096 (N_3096,N_2424,N_2715);
nand U3097 (N_3097,N_2570,N_2472);
nand U3098 (N_3098,N_2517,N_2734);
xor U3099 (N_3099,N_2494,N_2619);
xor U3100 (N_3100,N_2768,N_2734);
or U3101 (N_3101,N_2799,N_2433);
nor U3102 (N_3102,N_2719,N_2501);
nand U3103 (N_3103,N_2444,N_2562);
nand U3104 (N_3104,N_2469,N_2758);
nor U3105 (N_3105,N_2705,N_2755);
xnor U3106 (N_3106,N_2504,N_2493);
nor U3107 (N_3107,N_2503,N_2729);
or U3108 (N_3108,N_2680,N_2417);
or U3109 (N_3109,N_2492,N_2498);
xnor U3110 (N_3110,N_2779,N_2581);
or U3111 (N_3111,N_2613,N_2622);
and U3112 (N_3112,N_2511,N_2551);
nor U3113 (N_3113,N_2564,N_2781);
xnor U3114 (N_3114,N_2624,N_2703);
and U3115 (N_3115,N_2581,N_2513);
or U3116 (N_3116,N_2481,N_2508);
and U3117 (N_3117,N_2638,N_2554);
xnor U3118 (N_3118,N_2615,N_2425);
nor U3119 (N_3119,N_2419,N_2401);
or U3120 (N_3120,N_2540,N_2451);
xor U3121 (N_3121,N_2724,N_2796);
nand U3122 (N_3122,N_2762,N_2509);
xor U3123 (N_3123,N_2580,N_2674);
nor U3124 (N_3124,N_2725,N_2718);
and U3125 (N_3125,N_2781,N_2498);
nor U3126 (N_3126,N_2506,N_2560);
nand U3127 (N_3127,N_2441,N_2653);
nor U3128 (N_3128,N_2484,N_2441);
xnor U3129 (N_3129,N_2630,N_2480);
nor U3130 (N_3130,N_2650,N_2680);
and U3131 (N_3131,N_2670,N_2702);
nor U3132 (N_3132,N_2469,N_2615);
nand U3133 (N_3133,N_2592,N_2586);
and U3134 (N_3134,N_2640,N_2725);
xnor U3135 (N_3135,N_2493,N_2776);
xor U3136 (N_3136,N_2622,N_2522);
nand U3137 (N_3137,N_2659,N_2705);
nor U3138 (N_3138,N_2592,N_2550);
and U3139 (N_3139,N_2601,N_2685);
nor U3140 (N_3140,N_2599,N_2472);
xor U3141 (N_3141,N_2677,N_2641);
nand U3142 (N_3142,N_2577,N_2581);
nand U3143 (N_3143,N_2752,N_2721);
nor U3144 (N_3144,N_2512,N_2663);
nor U3145 (N_3145,N_2439,N_2685);
or U3146 (N_3146,N_2744,N_2457);
and U3147 (N_3147,N_2571,N_2663);
or U3148 (N_3148,N_2725,N_2606);
xnor U3149 (N_3149,N_2753,N_2465);
or U3150 (N_3150,N_2503,N_2414);
nand U3151 (N_3151,N_2641,N_2557);
and U3152 (N_3152,N_2415,N_2692);
nand U3153 (N_3153,N_2692,N_2765);
or U3154 (N_3154,N_2663,N_2424);
and U3155 (N_3155,N_2553,N_2527);
and U3156 (N_3156,N_2449,N_2688);
xnor U3157 (N_3157,N_2567,N_2547);
xnor U3158 (N_3158,N_2417,N_2703);
and U3159 (N_3159,N_2461,N_2785);
and U3160 (N_3160,N_2753,N_2503);
nor U3161 (N_3161,N_2418,N_2630);
or U3162 (N_3162,N_2660,N_2503);
or U3163 (N_3163,N_2560,N_2421);
or U3164 (N_3164,N_2639,N_2773);
nand U3165 (N_3165,N_2622,N_2417);
xor U3166 (N_3166,N_2520,N_2721);
xor U3167 (N_3167,N_2607,N_2513);
xor U3168 (N_3168,N_2537,N_2701);
or U3169 (N_3169,N_2763,N_2640);
nand U3170 (N_3170,N_2481,N_2698);
nand U3171 (N_3171,N_2469,N_2495);
nor U3172 (N_3172,N_2551,N_2626);
nand U3173 (N_3173,N_2476,N_2462);
xnor U3174 (N_3174,N_2400,N_2663);
and U3175 (N_3175,N_2410,N_2713);
and U3176 (N_3176,N_2732,N_2433);
nand U3177 (N_3177,N_2679,N_2548);
and U3178 (N_3178,N_2772,N_2549);
and U3179 (N_3179,N_2722,N_2492);
or U3180 (N_3180,N_2514,N_2493);
nand U3181 (N_3181,N_2539,N_2718);
nand U3182 (N_3182,N_2544,N_2706);
nor U3183 (N_3183,N_2716,N_2436);
and U3184 (N_3184,N_2612,N_2444);
or U3185 (N_3185,N_2502,N_2471);
xnor U3186 (N_3186,N_2481,N_2781);
or U3187 (N_3187,N_2592,N_2748);
and U3188 (N_3188,N_2736,N_2559);
xor U3189 (N_3189,N_2477,N_2402);
nand U3190 (N_3190,N_2691,N_2764);
or U3191 (N_3191,N_2497,N_2623);
or U3192 (N_3192,N_2462,N_2756);
and U3193 (N_3193,N_2789,N_2773);
or U3194 (N_3194,N_2793,N_2552);
xnor U3195 (N_3195,N_2523,N_2517);
nand U3196 (N_3196,N_2759,N_2705);
nand U3197 (N_3197,N_2438,N_2626);
nand U3198 (N_3198,N_2466,N_2690);
or U3199 (N_3199,N_2700,N_2701);
xor U3200 (N_3200,N_3070,N_2904);
nor U3201 (N_3201,N_3113,N_2842);
xnor U3202 (N_3202,N_3132,N_2822);
or U3203 (N_3203,N_3146,N_3148);
nand U3204 (N_3204,N_3053,N_2941);
nand U3205 (N_3205,N_3024,N_2869);
or U3206 (N_3206,N_3011,N_2866);
nor U3207 (N_3207,N_3119,N_3176);
and U3208 (N_3208,N_3134,N_3032);
and U3209 (N_3209,N_2848,N_3072);
or U3210 (N_3210,N_2908,N_2909);
and U3211 (N_3211,N_2997,N_3107);
nor U3212 (N_3212,N_3108,N_3057);
xor U3213 (N_3213,N_3085,N_3142);
and U3214 (N_3214,N_2993,N_2979);
xor U3215 (N_3215,N_2964,N_3105);
and U3216 (N_3216,N_2934,N_3028);
xor U3217 (N_3217,N_3060,N_3138);
xnor U3218 (N_3218,N_2931,N_3094);
nand U3219 (N_3219,N_3124,N_3062);
nand U3220 (N_3220,N_3144,N_2870);
or U3221 (N_3221,N_3069,N_3130);
and U3222 (N_3222,N_3123,N_2973);
or U3223 (N_3223,N_3087,N_2975);
and U3224 (N_3224,N_3080,N_2896);
nor U3225 (N_3225,N_2922,N_2855);
or U3226 (N_3226,N_3161,N_2968);
and U3227 (N_3227,N_3005,N_2877);
and U3228 (N_3228,N_2950,N_3051);
or U3229 (N_3229,N_3003,N_2906);
xor U3230 (N_3230,N_2803,N_2923);
and U3231 (N_3231,N_3008,N_3115);
nor U3232 (N_3232,N_3137,N_3031);
nand U3233 (N_3233,N_2834,N_3125);
nor U3234 (N_3234,N_3101,N_3086);
and U3235 (N_3235,N_2804,N_2945);
nor U3236 (N_3236,N_3066,N_3061);
or U3237 (N_3237,N_3166,N_2988);
nor U3238 (N_3238,N_2971,N_2925);
nand U3239 (N_3239,N_3191,N_3155);
xnor U3240 (N_3240,N_2930,N_2825);
or U3241 (N_3241,N_2985,N_2903);
nor U3242 (N_3242,N_3180,N_2990);
nor U3243 (N_3243,N_3199,N_2991);
nor U3244 (N_3244,N_2876,N_3065);
nand U3245 (N_3245,N_3012,N_3126);
nand U3246 (N_3246,N_3046,N_2847);
and U3247 (N_3247,N_2940,N_2829);
xor U3248 (N_3248,N_3077,N_3095);
nand U3249 (N_3249,N_2826,N_3047);
xnor U3250 (N_3250,N_3170,N_3045);
xnor U3251 (N_3251,N_3078,N_2886);
nor U3252 (N_3252,N_3151,N_2806);
xor U3253 (N_3253,N_3135,N_3149);
nor U3254 (N_3254,N_2958,N_2969);
xnor U3255 (N_3255,N_3136,N_2933);
or U3256 (N_3256,N_3145,N_3091);
or U3257 (N_3257,N_2824,N_2998);
nor U3258 (N_3258,N_2860,N_2924);
nor U3259 (N_3259,N_2843,N_2862);
nand U3260 (N_3260,N_2844,N_3006);
and U3261 (N_3261,N_2871,N_3165);
xor U3262 (N_3262,N_2918,N_2872);
nor U3263 (N_3263,N_3073,N_3188);
nand U3264 (N_3264,N_2852,N_3088);
or U3265 (N_3265,N_2984,N_2819);
nand U3266 (N_3266,N_3030,N_3168);
and U3267 (N_3267,N_2817,N_2816);
xor U3268 (N_3268,N_2957,N_2944);
or U3269 (N_3269,N_3017,N_2890);
nand U3270 (N_3270,N_3139,N_2987);
and U3271 (N_3271,N_3037,N_2912);
nor U3272 (N_3272,N_2888,N_3043);
nor U3273 (N_3273,N_3153,N_2881);
nand U3274 (N_3274,N_2823,N_2996);
xor U3275 (N_3275,N_2821,N_3158);
nor U3276 (N_3276,N_2902,N_2937);
nor U3277 (N_3277,N_3027,N_2899);
nand U3278 (N_3278,N_2995,N_3175);
nand U3279 (N_3279,N_3067,N_2884);
and U3280 (N_3280,N_3118,N_3013);
nor U3281 (N_3281,N_2838,N_2856);
and U3282 (N_3282,N_2915,N_2895);
nand U3283 (N_3283,N_2916,N_2893);
and U3284 (N_3284,N_2809,N_2959);
nor U3285 (N_3285,N_3172,N_3100);
nand U3286 (N_3286,N_3058,N_3019);
nand U3287 (N_3287,N_2882,N_2919);
or U3288 (N_3288,N_2837,N_3016);
nor U3289 (N_3289,N_3103,N_2976);
or U3290 (N_3290,N_3127,N_3049);
and U3291 (N_3291,N_2850,N_3198);
xor U3292 (N_3292,N_3015,N_2974);
nand U3293 (N_3293,N_3026,N_2952);
and U3294 (N_3294,N_2875,N_3143);
nand U3295 (N_3295,N_2857,N_2867);
nor U3296 (N_3296,N_3002,N_3154);
and U3297 (N_3297,N_3162,N_2831);
or U3298 (N_3298,N_2808,N_2914);
nand U3299 (N_3299,N_2865,N_3193);
and U3300 (N_3300,N_3056,N_2929);
xor U3301 (N_3301,N_2948,N_2953);
nand U3302 (N_3302,N_3014,N_2994);
nand U3303 (N_3303,N_3152,N_3197);
nor U3304 (N_3304,N_3048,N_3018);
or U3305 (N_3305,N_3004,N_3141);
nor U3306 (N_3306,N_2943,N_2961);
and U3307 (N_3307,N_3114,N_2807);
or U3308 (N_3308,N_3074,N_2849);
nand U3309 (N_3309,N_2839,N_3010);
xor U3310 (N_3310,N_3167,N_2854);
xnor U3311 (N_3311,N_3092,N_3187);
xnor U3312 (N_3312,N_2917,N_2840);
and U3313 (N_3313,N_2954,N_2983);
and U3314 (N_3314,N_3147,N_3076);
xnor U3315 (N_3315,N_2980,N_2853);
xor U3316 (N_3316,N_3068,N_2960);
and U3317 (N_3317,N_3038,N_2981);
and U3318 (N_3318,N_3097,N_2939);
nor U3319 (N_3319,N_2861,N_3116);
and U3320 (N_3320,N_3042,N_3110);
nor U3321 (N_3321,N_3009,N_3156);
xor U3322 (N_3322,N_2898,N_2805);
and U3323 (N_3323,N_3102,N_3163);
nand U3324 (N_3324,N_3173,N_3007);
nor U3325 (N_3325,N_2815,N_3195);
nor U3326 (N_3326,N_2999,N_3071);
and U3327 (N_3327,N_3196,N_2935);
nor U3328 (N_3328,N_2818,N_3020);
and U3329 (N_3329,N_2835,N_2977);
nor U3330 (N_3330,N_3169,N_3157);
or U3331 (N_3331,N_2830,N_3025);
and U3332 (N_3332,N_2962,N_3039);
nand U3333 (N_3333,N_2863,N_2810);
or U3334 (N_3334,N_2883,N_3186);
nand U3335 (N_3335,N_3178,N_2900);
nor U3336 (N_3336,N_3079,N_2972);
and U3337 (N_3337,N_2905,N_2947);
xor U3338 (N_3338,N_2928,N_2942);
nand U3339 (N_3339,N_3159,N_2966);
and U3340 (N_3340,N_2967,N_2926);
nand U3341 (N_3341,N_3112,N_3096);
or U3342 (N_3342,N_2913,N_2949);
nor U3343 (N_3343,N_2868,N_2874);
or U3344 (N_3344,N_3098,N_2992);
xnor U3345 (N_3345,N_2921,N_2907);
and U3346 (N_3346,N_2878,N_3104);
xor U3347 (N_3347,N_3109,N_2978);
and U3348 (N_3348,N_2827,N_3117);
xnor U3349 (N_3349,N_3160,N_2811);
nor U3350 (N_3350,N_2970,N_3050);
xnor U3351 (N_3351,N_3099,N_3082);
nand U3352 (N_3352,N_2946,N_3185);
nor U3353 (N_3353,N_3052,N_2833);
and U3354 (N_3354,N_3059,N_3192);
xor U3355 (N_3355,N_3184,N_2832);
nand U3356 (N_3356,N_3083,N_2891);
and U3357 (N_3357,N_3111,N_3022);
xor U3358 (N_3358,N_3063,N_2956);
nand U3359 (N_3359,N_3120,N_3189);
or U3360 (N_3360,N_2820,N_3190);
xnor U3361 (N_3361,N_3121,N_3122);
nor U3362 (N_3362,N_3023,N_3000);
nand U3363 (N_3363,N_2814,N_3064);
xor U3364 (N_3364,N_3093,N_3001);
xnor U3365 (N_3365,N_3054,N_3182);
xnor U3366 (N_3366,N_2879,N_3131);
xor U3367 (N_3367,N_3133,N_2936);
nand U3368 (N_3368,N_2965,N_2841);
and U3369 (N_3369,N_2864,N_2800);
or U3370 (N_3370,N_3129,N_3035);
nor U3371 (N_3371,N_2836,N_2938);
nand U3372 (N_3372,N_2801,N_3171);
nand U3373 (N_3373,N_2927,N_3174);
nand U3374 (N_3374,N_2894,N_3090);
nor U3375 (N_3375,N_2897,N_2846);
and U3376 (N_3376,N_2873,N_2858);
nor U3377 (N_3377,N_2955,N_2880);
and U3378 (N_3378,N_3106,N_2911);
nand U3379 (N_3379,N_3179,N_2910);
nor U3380 (N_3380,N_3177,N_2982);
xor U3381 (N_3381,N_3150,N_2963);
and U3382 (N_3382,N_3029,N_2812);
and U3383 (N_3383,N_2813,N_3081);
or U3384 (N_3384,N_3089,N_2986);
and U3385 (N_3385,N_3055,N_2887);
nand U3386 (N_3386,N_3021,N_2851);
and U3387 (N_3387,N_2885,N_3041);
xnor U3388 (N_3388,N_3034,N_2932);
nand U3389 (N_3389,N_2920,N_2802);
nor U3390 (N_3390,N_3075,N_3140);
or U3391 (N_3391,N_2889,N_2892);
nand U3392 (N_3392,N_3044,N_3040);
nor U3393 (N_3393,N_3164,N_3036);
and U3394 (N_3394,N_2901,N_3033);
nand U3395 (N_3395,N_3181,N_3194);
or U3396 (N_3396,N_3183,N_3084);
nor U3397 (N_3397,N_3128,N_2859);
xnor U3398 (N_3398,N_2951,N_2828);
and U3399 (N_3399,N_2845,N_2989);
xor U3400 (N_3400,N_2868,N_3199);
and U3401 (N_3401,N_2837,N_3002);
xor U3402 (N_3402,N_3009,N_3172);
nor U3403 (N_3403,N_2957,N_3122);
or U3404 (N_3404,N_2970,N_2936);
or U3405 (N_3405,N_3165,N_2870);
and U3406 (N_3406,N_2941,N_3156);
and U3407 (N_3407,N_3013,N_3070);
or U3408 (N_3408,N_2891,N_2801);
or U3409 (N_3409,N_3103,N_2894);
or U3410 (N_3410,N_2878,N_2835);
xor U3411 (N_3411,N_3000,N_2830);
nor U3412 (N_3412,N_3056,N_3186);
nor U3413 (N_3413,N_3092,N_2947);
nand U3414 (N_3414,N_2973,N_2926);
nor U3415 (N_3415,N_2874,N_2934);
xnor U3416 (N_3416,N_2854,N_3134);
nor U3417 (N_3417,N_2910,N_2902);
and U3418 (N_3418,N_2860,N_2866);
xor U3419 (N_3419,N_3014,N_2962);
and U3420 (N_3420,N_2979,N_3050);
xor U3421 (N_3421,N_3112,N_2994);
and U3422 (N_3422,N_2989,N_2833);
and U3423 (N_3423,N_2918,N_2947);
or U3424 (N_3424,N_2911,N_3014);
xnor U3425 (N_3425,N_2999,N_3131);
xor U3426 (N_3426,N_2822,N_2942);
and U3427 (N_3427,N_3106,N_2945);
nand U3428 (N_3428,N_3142,N_3063);
nor U3429 (N_3429,N_2968,N_3024);
nor U3430 (N_3430,N_2847,N_3193);
xor U3431 (N_3431,N_3001,N_3123);
xnor U3432 (N_3432,N_2962,N_2957);
nand U3433 (N_3433,N_3040,N_3196);
xor U3434 (N_3434,N_3152,N_2992);
nand U3435 (N_3435,N_2980,N_3041);
nand U3436 (N_3436,N_3117,N_2970);
xnor U3437 (N_3437,N_2945,N_3028);
nor U3438 (N_3438,N_3155,N_2821);
nor U3439 (N_3439,N_3071,N_3185);
xor U3440 (N_3440,N_2994,N_2825);
xor U3441 (N_3441,N_2938,N_3177);
nand U3442 (N_3442,N_3056,N_2924);
and U3443 (N_3443,N_3197,N_2835);
nor U3444 (N_3444,N_2856,N_3087);
nor U3445 (N_3445,N_2926,N_3159);
nand U3446 (N_3446,N_2906,N_2864);
or U3447 (N_3447,N_2873,N_3069);
and U3448 (N_3448,N_2998,N_2818);
nor U3449 (N_3449,N_2826,N_2844);
or U3450 (N_3450,N_2924,N_3030);
xnor U3451 (N_3451,N_3012,N_2832);
nand U3452 (N_3452,N_3187,N_3077);
xor U3453 (N_3453,N_2806,N_3042);
and U3454 (N_3454,N_2940,N_2957);
or U3455 (N_3455,N_3121,N_2820);
xnor U3456 (N_3456,N_3191,N_3139);
or U3457 (N_3457,N_2900,N_3168);
xor U3458 (N_3458,N_3024,N_2865);
and U3459 (N_3459,N_2985,N_3175);
and U3460 (N_3460,N_3157,N_3150);
and U3461 (N_3461,N_3013,N_2806);
and U3462 (N_3462,N_3109,N_2997);
nor U3463 (N_3463,N_3168,N_2843);
and U3464 (N_3464,N_3143,N_2963);
and U3465 (N_3465,N_2863,N_3070);
xnor U3466 (N_3466,N_2972,N_3085);
or U3467 (N_3467,N_3079,N_3163);
or U3468 (N_3468,N_3037,N_3160);
and U3469 (N_3469,N_3185,N_3172);
nor U3470 (N_3470,N_3053,N_3156);
and U3471 (N_3471,N_3116,N_2842);
and U3472 (N_3472,N_2800,N_3090);
and U3473 (N_3473,N_2899,N_2856);
nand U3474 (N_3474,N_3037,N_3015);
nand U3475 (N_3475,N_3118,N_3010);
nor U3476 (N_3476,N_3101,N_2911);
xor U3477 (N_3477,N_3157,N_3109);
nor U3478 (N_3478,N_3099,N_2991);
or U3479 (N_3479,N_3071,N_3091);
nand U3480 (N_3480,N_3151,N_2890);
and U3481 (N_3481,N_3006,N_3120);
and U3482 (N_3482,N_3176,N_2980);
and U3483 (N_3483,N_2804,N_3021);
nor U3484 (N_3484,N_2821,N_2941);
nor U3485 (N_3485,N_2832,N_2927);
and U3486 (N_3486,N_2935,N_2995);
and U3487 (N_3487,N_2877,N_3137);
xor U3488 (N_3488,N_3072,N_2989);
and U3489 (N_3489,N_2865,N_2873);
xnor U3490 (N_3490,N_2948,N_3047);
nor U3491 (N_3491,N_3038,N_2991);
or U3492 (N_3492,N_3046,N_3174);
nand U3493 (N_3493,N_3011,N_2811);
or U3494 (N_3494,N_2925,N_2898);
or U3495 (N_3495,N_2829,N_3128);
xnor U3496 (N_3496,N_2998,N_2942);
nand U3497 (N_3497,N_3014,N_3142);
and U3498 (N_3498,N_3121,N_2817);
nor U3499 (N_3499,N_2816,N_2877);
nor U3500 (N_3500,N_2960,N_2903);
and U3501 (N_3501,N_2918,N_2955);
nor U3502 (N_3502,N_2916,N_3043);
and U3503 (N_3503,N_3155,N_3084);
nor U3504 (N_3504,N_2965,N_2954);
nor U3505 (N_3505,N_3112,N_2903);
nand U3506 (N_3506,N_3174,N_2850);
nand U3507 (N_3507,N_3168,N_3145);
xnor U3508 (N_3508,N_3016,N_2920);
and U3509 (N_3509,N_2910,N_2812);
nand U3510 (N_3510,N_3060,N_2866);
nor U3511 (N_3511,N_2947,N_3007);
and U3512 (N_3512,N_3099,N_3160);
nor U3513 (N_3513,N_3190,N_3093);
and U3514 (N_3514,N_3049,N_3055);
or U3515 (N_3515,N_2919,N_3059);
xnor U3516 (N_3516,N_3044,N_3161);
and U3517 (N_3517,N_3173,N_2855);
and U3518 (N_3518,N_2881,N_2848);
and U3519 (N_3519,N_2877,N_3123);
nand U3520 (N_3520,N_2979,N_3110);
nand U3521 (N_3521,N_2912,N_2814);
nor U3522 (N_3522,N_3187,N_2941);
or U3523 (N_3523,N_3086,N_3196);
xnor U3524 (N_3524,N_2870,N_2944);
nand U3525 (N_3525,N_3150,N_2946);
and U3526 (N_3526,N_2983,N_3100);
xor U3527 (N_3527,N_2843,N_3029);
or U3528 (N_3528,N_3085,N_3185);
and U3529 (N_3529,N_3161,N_2868);
xor U3530 (N_3530,N_2971,N_3170);
or U3531 (N_3531,N_2903,N_2935);
xor U3532 (N_3532,N_2833,N_3169);
nand U3533 (N_3533,N_3125,N_2876);
nand U3534 (N_3534,N_3165,N_3017);
nor U3535 (N_3535,N_2853,N_2801);
nand U3536 (N_3536,N_2989,N_2995);
or U3537 (N_3537,N_2921,N_3150);
nor U3538 (N_3538,N_3101,N_3075);
or U3539 (N_3539,N_3199,N_2849);
nand U3540 (N_3540,N_2940,N_2950);
nand U3541 (N_3541,N_2916,N_2985);
xor U3542 (N_3542,N_3164,N_3028);
nand U3543 (N_3543,N_3147,N_3065);
nand U3544 (N_3544,N_3078,N_3006);
nand U3545 (N_3545,N_3152,N_2920);
nor U3546 (N_3546,N_3001,N_3071);
and U3547 (N_3547,N_2836,N_2902);
xor U3548 (N_3548,N_2877,N_3114);
nor U3549 (N_3549,N_3174,N_3157);
nand U3550 (N_3550,N_3164,N_3132);
nor U3551 (N_3551,N_3160,N_2876);
and U3552 (N_3552,N_2913,N_2839);
nand U3553 (N_3553,N_3141,N_2949);
and U3554 (N_3554,N_2857,N_2869);
nand U3555 (N_3555,N_3157,N_3076);
nand U3556 (N_3556,N_3091,N_2910);
xor U3557 (N_3557,N_2970,N_2823);
nor U3558 (N_3558,N_2914,N_2960);
nand U3559 (N_3559,N_3046,N_3108);
and U3560 (N_3560,N_2920,N_2931);
or U3561 (N_3561,N_3162,N_2970);
xnor U3562 (N_3562,N_3066,N_3166);
or U3563 (N_3563,N_2833,N_3084);
or U3564 (N_3564,N_2952,N_3160);
and U3565 (N_3565,N_3093,N_3128);
or U3566 (N_3566,N_3049,N_3101);
and U3567 (N_3567,N_3198,N_2921);
xnor U3568 (N_3568,N_3034,N_2952);
xor U3569 (N_3569,N_3125,N_2829);
and U3570 (N_3570,N_2843,N_2821);
and U3571 (N_3571,N_2902,N_2985);
or U3572 (N_3572,N_2950,N_2931);
nand U3573 (N_3573,N_3149,N_3162);
xor U3574 (N_3574,N_2892,N_3016);
or U3575 (N_3575,N_2985,N_2930);
xnor U3576 (N_3576,N_2873,N_3098);
or U3577 (N_3577,N_2995,N_2881);
xnor U3578 (N_3578,N_3029,N_3104);
or U3579 (N_3579,N_2845,N_3197);
nor U3580 (N_3580,N_2968,N_2807);
nor U3581 (N_3581,N_2917,N_3146);
xor U3582 (N_3582,N_2873,N_3015);
nand U3583 (N_3583,N_3034,N_2942);
and U3584 (N_3584,N_3128,N_2968);
nor U3585 (N_3585,N_2923,N_2965);
nand U3586 (N_3586,N_3193,N_2808);
and U3587 (N_3587,N_2934,N_3098);
nand U3588 (N_3588,N_3065,N_2817);
and U3589 (N_3589,N_3148,N_2990);
and U3590 (N_3590,N_2998,N_3100);
and U3591 (N_3591,N_3068,N_2999);
nor U3592 (N_3592,N_2812,N_2858);
xor U3593 (N_3593,N_3094,N_2944);
nor U3594 (N_3594,N_3122,N_3058);
xor U3595 (N_3595,N_3116,N_3168);
or U3596 (N_3596,N_3129,N_2880);
or U3597 (N_3597,N_3113,N_3063);
xnor U3598 (N_3598,N_2995,N_3105);
xor U3599 (N_3599,N_3047,N_3178);
and U3600 (N_3600,N_3371,N_3234);
nor U3601 (N_3601,N_3301,N_3389);
nor U3602 (N_3602,N_3463,N_3481);
or U3603 (N_3603,N_3358,N_3265);
nor U3604 (N_3604,N_3317,N_3528);
nand U3605 (N_3605,N_3202,N_3263);
xor U3606 (N_3606,N_3342,N_3491);
or U3607 (N_3607,N_3309,N_3414);
and U3608 (N_3608,N_3323,N_3589);
xor U3609 (N_3609,N_3211,N_3538);
nor U3610 (N_3610,N_3270,N_3258);
and U3611 (N_3611,N_3210,N_3478);
or U3612 (N_3612,N_3483,N_3432);
or U3613 (N_3613,N_3386,N_3373);
xnor U3614 (N_3614,N_3369,N_3430);
nand U3615 (N_3615,N_3391,N_3570);
nor U3616 (N_3616,N_3372,N_3330);
nor U3617 (N_3617,N_3361,N_3470);
and U3618 (N_3618,N_3465,N_3446);
nor U3619 (N_3619,N_3366,N_3542);
or U3620 (N_3620,N_3579,N_3501);
xor U3621 (N_3621,N_3339,N_3338);
nor U3622 (N_3622,N_3474,N_3255);
or U3623 (N_3623,N_3215,N_3519);
nand U3624 (N_3624,N_3375,N_3468);
nor U3625 (N_3625,N_3547,N_3283);
xor U3626 (N_3626,N_3572,N_3537);
nand U3627 (N_3627,N_3569,N_3487);
nor U3628 (N_3628,N_3354,N_3295);
and U3629 (N_3629,N_3401,N_3461);
nand U3630 (N_3630,N_3298,N_3237);
and U3631 (N_3631,N_3521,N_3477);
or U3632 (N_3632,N_3525,N_3396);
and U3633 (N_3633,N_3213,N_3314);
nor U3634 (N_3634,N_3239,N_3208);
nand U3635 (N_3635,N_3412,N_3480);
or U3636 (N_3636,N_3229,N_3260);
xor U3637 (N_3637,N_3225,N_3413);
nand U3638 (N_3638,N_3290,N_3273);
and U3639 (N_3639,N_3293,N_3532);
nand U3640 (N_3640,N_3495,N_3454);
xnor U3641 (N_3641,N_3559,N_3421);
nor U3642 (N_3642,N_3564,N_3233);
and U3643 (N_3643,N_3466,N_3580);
nand U3644 (N_3644,N_3508,N_3425);
nand U3645 (N_3645,N_3246,N_3464);
and U3646 (N_3646,N_3378,N_3485);
or U3647 (N_3647,N_3302,N_3400);
or U3648 (N_3648,N_3226,N_3434);
nand U3649 (N_3649,N_3367,N_3287);
nor U3650 (N_3650,N_3571,N_3545);
or U3651 (N_3651,N_3451,N_3303);
nand U3652 (N_3652,N_3473,N_3512);
or U3653 (N_3653,N_3388,N_3384);
nand U3654 (N_3654,N_3513,N_3475);
xor U3655 (N_3655,N_3201,N_3274);
xor U3656 (N_3656,N_3341,N_3228);
or U3657 (N_3657,N_3348,N_3533);
xor U3658 (N_3658,N_3447,N_3516);
and U3659 (N_3659,N_3522,N_3460);
xnor U3660 (N_3660,N_3279,N_3422);
nor U3661 (N_3661,N_3574,N_3515);
and U3662 (N_3662,N_3312,N_3257);
xnor U3663 (N_3663,N_3252,N_3449);
or U3664 (N_3664,N_3536,N_3504);
or U3665 (N_3665,N_3462,N_3418);
nor U3666 (N_3666,N_3482,N_3558);
xnor U3667 (N_3667,N_3242,N_3496);
or U3668 (N_3668,N_3444,N_3346);
and U3669 (N_3669,N_3299,N_3500);
nand U3670 (N_3670,N_3221,N_3588);
or U3671 (N_3671,N_3356,N_3514);
xnor U3672 (N_3672,N_3230,N_3305);
nand U3673 (N_3673,N_3380,N_3429);
nand U3674 (N_3674,N_3292,N_3256);
or U3675 (N_3675,N_3546,N_3435);
or U3676 (N_3676,N_3405,N_3506);
or U3677 (N_3677,N_3592,N_3551);
or U3678 (N_3678,N_3486,N_3324);
or U3679 (N_3679,N_3370,N_3236);
and U3680 (N_3680,N_3300,N_3423);
nand U3681 (N_3681,N_3565,N_3336);
nor U3682 (N_3682,N_3499,N_3296);
nor U3683 (N_3683,N_3539,N_3549);
xor U3684 (N_3684,N_3280,N_3355);
nand U3685 (N_3685,N_3598,N_3523);
nor U3686 (N_3686,N_3593,N_3448);
or U3687 (N_3687,N_3254,N_3411);
and U3688 (N_3688,N_3526,N_3288);
nand U3689 (N_3689,N_3364,N_3212);
xor U3690 (N_3690,N_3219,N_3489);
or U3691 (N_3691,N_3584,N_3245);
or U3692 (N_3692,N_3479,N_3507);
nand U3693 (N_3693,N_3352,N_3382);
xnor U3694 (N_3694,N_3315,N_3232);
and U3695 (N_3695,N_3222,N_3224);
and U3696 (N_3696,N_3417,N_3471);
or U3697 (N_3697,N_3320,N_3248);
xor U3698 (N_3698,N_3575,N_3573);
and U3699 (N_3699,N_3281,N_3376);
nor U3700 (N_3700,N_3262,N_3377);
nand U3701 (N_3701,N_3307,N_3502);
nand U3702 (N_3702,N_3490,N_3328);
xnor U3703 (N_3703,N_3428,N_3277);
nand U3704 (N_3704,N_3326,N_3431);
nor U3705 (N_3705,N_3553,N_3294);
or U3706 (N_3706,N_3310,N_3445);
and U3707 (N_3707,N_3319,N_3590);
xor U3708 (N_3708,N_3583,N_3455);
xnor U3709 (N_3709,N_3531,N_3567);
xnor U3710 (N_3710,N_3443,N_3472);
nor U3711 (N_3711,N_3476,N_3505);
and U3712 (N_3712,N_3322,N_3340);
nand U3713 (N_3713,N_3209,N_3544);
xor U3714 (N_3714,N_3568,N_3581);
nor U3715 (N_3715,N_3407,N_3497);
xor U3716 (N_3716,N_3267,N_3206);
nor U3717 (N_3717,N_3214,N_3420);
xor U3718 (N_3718,N_3241,N_3408);
and U3719 (N_3719,N_3395,N_3333);
or U3720 (N_3720,N_3488,N_3363);
nand U3721 (N_3721,N_3510,N_3562);
nand U3722 (N_3722,N_3393,N_3403);
nor U3723 (N_3723,N_3387,N_3596);
or U3724 (N_3724,N_3253,N_3509);
and U3725 (N_3725,N_3344,N_3394);
or U3726 (N_3726,N_3285,N_3441);
and U3727 (N_3727,N_3313,N_3207);
or U3728 (N_3728,N_3304,N_3216);
and U3729 (N_3729,N_3535,N_3306);
xor U3730 (N_3730,N_3297,N_3453);
and U3731 (N_3731,N_3351,N_3227);
xor U3732 (N_3732,N_3249,N_3238);
nand U3733 (N_3733,N_3534,N_3576);
nand U3734 (N_3734,N_3436,N_3540);
nor U3735 (N_3735,N_3467,N_3345);
and U3736 (N_3736,N_3511,N_3275);
or U3737 (N_3737,N_3282,N_3362);
nor U3738 (N_3738,N_3349,N_3360);
and U3739 (N_3739,N_3554,N_3374);
xnor U3740 (N_3740,N_3289,N_3577);
xnor U3741 (N_3741,N_3585,N_3550);
nor U3742 (N_3742,N_3334,N_3271);
nor U3743 (N_3743,N_3368,N_3347);
xor U3744 (N_3744,N_3442,N_3243);
nand U3745 (N_3745,N_3205,N_3259);
xor U3746 (N_3746,N_3484,N_3518);
nand U3747 (N_3747,N_3591,N_3269);
nor U3748 (N_3748,N_3231,N_3251);
xor U3749 (N_3749,N_3332,N_3308);
nor U3750 (N_3750,N_3566,N_3220);
nand U3751 (N_3751,N_3335,N_3548);
or U3752 (N_3752,N_3286,N_3557);
nand U3753 (N_3753,N_3582,N_3452);
nand U3754 (N_3754,N_3529,N_3530);
or U3755 (N_3755,N_3524,N_3527);
xor U3756 (N_3756,N_3594,N_3469);
and U3757 (N_3757,N_3331,N_3498);
nor U3758 (N_3758,N_3398,N_3321);
or U3759 (N_3759,N_3586,N_3433);
nand U3760 (N_3760,N_3311,N_3240);
or U3761 (N_3761,N_3494,N_3204);
nand U3762 (N_3762,N_3459,N_3595);
or U3763 (N_3763,N_3217,N_3385);
nor U3764 (N_3764,N_3415,N_3250);
xnor U3765 (N_3765,N_3218,N_3560);
nand U3766 (N_3766,N_3223,N_3284);
nor U3767 (N_3767,N_3404,N_3261);
xor U3768 (N_3768,N_3440,N_3555);
nor U3769 (N_3769,N_3278,N_3397);
or U3770 (N_3770,N_3457,N_3235);
nor U3771 (N_3771,N_3543,N_3424);
and U3772 (N_3772,N_3552,N_3383);
or U3773 (N_3773,N_3556,N_3327);
or U3774 (N_3774,N_3325,N_3439);
or U3775 (N_3775,N_3563,N_3357);
or U3776 (N_3776,N_3438,N_3247);
or U3777 (N_3777,N_3587,N_3541);
nor U3778 (N_3778,N_3276,N_3406);
and U3779 (N_3779,N_3493,N_3343);
nor U3780 (N_3780,N_3203,N_3561);
and U3781 (N_3781,N_3492,N_3291);
or U3782 (N_3782,N_3200,N_3458);
xnor U3783 (N_3783,N_3392,N_3318);
or U3784 (N_3784,N_3410,N_3419);
xnor U3785 (N_3785,N_3599,N_3329);
or U3786 (N_3786,N_3365,N_3337);
nand U3787 (N_3787,N_3268,N_3520);
and U3788 (N_3788,N_3450,N_3437);
xor U3789 (N_3789,N_3578,N_3402);
and U3790 (N_3790,N_3426,N_3244);
xnor U3791 (N_3791,N_3399,N_3390);
and U3792 (N_3792,N_3353,N_3381);
nand U3793 (N_3793,N_3427,N_3416);
nor U3794 (N_3794,N_3316,N_3359);
xnor U3795 (N_3795,N_3379,N_3503);
nor U3796 (N_3796,N_3409,N_3456);
xor U3797 (N_3797,N_3266,N_3264);
nand U3798 (N_3798,N_3272,N_3350);
nand U3799 (N_3799,N_3517,N_3597);
nor U3800 (N_3800,N_3250,N_3397);
nand U3801 (N_3801,N_3247,N_3525);
and U3802 (N_3802,N_3255,N_3398);
nand U3803 (N_3803,N_3506,N_3259);
nor U3804 (N_3804,N_3525,N_3441);
or U3805 (N_3805,N_3461,N_3326);
xor U3806 (N_3806,N_3323,N_3401);
nand U3807 (N_3807,N_3498,N_3452);
or U3808 (N_3808,N_3214,N_3408);
xnor U3809 (N_3809,N_3210,N_3562);
xnor U3810 (N_3810,N_3435,N_3389);
xor U3811 (N_3811,N_3488,N_3247);
or U3812 (N_3812,N_3582,N_3449);
nor U3813 (N_3813,N_3598,N_3551);
nor U3814 (N_3814,N_3510,N_3227);
xnor U3815 (N_3815,N_3282,N_3342);
xnor U3816 (N_3816,N_3390,N_3254);
nor U3817 (N_3817,N_3568,N_3427);
nand U3818 (N_3818,N_3305,N_3428);
or U3819 (N_3819,N_3308,N_3279);
nand U3820 (N_3820,N_3492,N_3211);
and U3821 (N_3821,N_3519,N_3585);
or U3822 (N_3822,N_3361,N_3527);
nand U3823 (N_3823,N_3402,N_3256);
nand U3824 (N_3824,N_3206,N_3328);
nor U3825 (N_3825,N_3486,N_3345);
or U3826 (N_3826,N_3337,N_3217);
nand U3827 (N_3827,N_3510,N_3408);
and U3828 (N_3828,N_3241,N_3393);
xnor U3829 (N_3829,N_3466,N_3568);
and U3830 (N_3830,N_3224,N_3357);
or U3831 (N_3831,N_3394,N_3378);
and U3832 (N_3832,N_3330,N_3548);
xor U3833 (N_3833,N_3484,N_3338);
and U3834 (N_3834,N_3464,N_3592);
nand U3835 (N_3835,N_3271,N_3426);
nor U3836 (N_3836,N_3492,N_3512);
and U3837 (N_3837,N_3598,N_3480);
or U3838 (N_3838,N_3285,N_3578);
nand U3839 (N_3839,N_3506,N_3352);
and U3840 (N_3840,N_3235,N_3376);
xor U3841 (N_3841,N_3242,N_3545);
or U3842 (N_3842,N_3465,N_3278);
or U3843 (N_3843,N_3578,N_3555);
xor U3844 (N_3844,N_3492,N_3550);
xnor U3845 (N_3845,N_3361,N_3598);
nor U3846 (N_3846,N_3522,N_3232);
or U3847 (N_3847,N_3319,N_3492);
nor U3848 (N_3848,N_3293,N_3522);
xor U3849 (N_3849,N_3422,N_3580);
nand U3850 (N_3850,N_3504,N_3200);
or U3851 (N_3851,N_3510,N_3419);
and U3852 (N_3852,N_3412,N_3531);
xnor U3853 (N_3853,N_3532,N_3318);
or U3854 (N_3854,N_3371,N_3570);
nor U3855 (N_3855,N_3577,N_3457);
or U3856 (N_3856,N_3302,N_3421);
and U3857 (N_3857,N_3486,N_3453);
nand U3858 (N_3858,N_3463,N_3506);
xor U3859 (N_3859,N_3413,N_3458);
nand U3860 (N_3860,N_3451,N_3358);
xor U3861 (N_3861,N_3484,N_3331);
and U3862 (N_3862,N_3446,N_3412);
xor U3863 (N_3863,N_3565,N_3583);
nand U3864 (N_3864,N_3229,N_3240);
nor U3865 (N_3865,N_3480,N_3546);
or U3866 (N_3866,N_3261,N_3564);
and U3867 (N_3867,N_3241,N_3579);
nor U3868 (N_3868,N_3346,N_3376);
or U3869 (N_3869,N_3488,N_3477);
xor U3870 (N_3870,N_3330,N_3233);
xor U3871 (N_3871,N_3250,N_3319);
and U3872 (N_3872,N_3321,N_3272);
xor U3873 (N_3873,N_3266,N_3551);
or U3874 (N_3874,N_3579,N_3306);
xnor U3875 (N_3875,N_3551,N_3330);
nand U3876 (N_3876,N_3416,N_3352);
nand U3877 (N_3877,N_3252,N_3477);
nor U3878 (N_3878,N_3511,N_3514);
nor U3879 (N_3879,N_3487,N_3316);
nand U3880 (N_3880,N_3569,N_3392);
xor U3881 (N_3881,N_3408,N_3349);
and U3882 (N_3882,N_3387,N_3504);
xor U3883 (N_3883,N_3419,N_3489);
and U3884 (N_3884,N_3328,N_3407);
or U3885 (N_3885,N_3344,N_3480);
or U3886 (N_3886,N_3363,N_3598);
nor U3887 (N_3887,N_3420,N_3542);
and U3888 (N_3888,N_3350,N_3529);
and U3889 (N_3889,N_3353,N_3554);
xnor U3890 (N_3890,N_3252,N_3304);
and U3891 (N_3891,N_3516,N_3309);
and U3892 (N_3892,N_3295,N_3584);
nand U3893 (N_3893,N_3516,N_3452);
nor U3894 (N_3894,N_3516,N_3301);
nand U3895 (N_3895,N_3248,N_3223);
or U3896 (N_3896,N_3563,N_3242);
or U3897 (N_3897,N_3562,N_3211);
nand U3898 (N_3898,N_3344,N_3513);
nor U3899 (N_3899,N_3594,N_3428);
xor U3900 (N_3900,N_3321,N_3314);
nor U3901 (N_3901,N_3243,N_3231);
xnor U3902 (N_3902,N_3588,N_3572);
and U3903 (N_3903,N_3356,N_3523);
nand U3904 (N_3904,N_3271,N_3340);
nand U3905 (N_3905,N_3328,N_3262);
or U3906 (N_3906,N_3354,N_3575);
or U3907 (N_3907,N_3492,N_3347);
and U3908 (N_3908,N_3564,N_3520);
xor U3909 (N_3909,N_3340,N_3214);
and U3910 (N_3910,N_3353,N_3428);
nand U3911 (N_3911,N_3266,N_3356);
nor U3912 (N_3912,N_3247,N_3561);
or U3913 (N_3913,N_3343,N_3446);
xor U3914 (N_3914,N_3430,N_3215);
nor U3915 (N_3915,N_3340,N_3344);
and U3916 (N_3916,N_3306,N_3571);
and U3917 (N_3917,N_3343,N_3218);
nor U3918 (N_3918,N_3289,N_3494);
nand U3919 (N_3919,N_3298,N_3223);
nand U3920 (N_3920,N_3418,N_3351);
nor U3921 (N_3921,N_3337,N_3599);
or U3922 (N_3922,N_3358,N_3396);
and U3923 (N_3923,N_3207,N_3509);
nand U3924 (N_3924,N_3236,N_3599);
or U3925 (N_3925,N_3391,N_3246);
nand U3926 (N_3926,N_3593,N_3555);
nor U3927 (N_3927,N_3517,N_3242);
nand U3928 (N_3928,N_3539,N_3371);
or U3929 (N_3929,N_3510,N_3386);
xnor U3930 (N_3930,N_3486,N_3515);
nor U3931 (N_3931,N_3274,N_3572);
nor U3932 (N_3932,N_3200,N_3492);
nor U3933 (N_3933,N_3320,N_3341);
nor U3934 (N_3934,N_3485,N_3211);
nand U3935 (N_3935,N_3596,N_3512);
xnor U3936 (N_3936,N_3513,N_3353);
and U3937 (N_3937,N_3200,N_3574);
xor U3938 (N_3938,N_3575,N_3595);
nor U3939 (N_3939,N_3483,N_3381);
nor U3940 (N_3940,N_3402,N_3525);
nand U3941 (N_3941,N_3313,N_3397);
xor U3942 (N_3942,N_3203,N_3490);
nand U3943 (N_3943,N_3438,N_3570);
or U3944 (N_3944,N_3480,N_3475);
nand U3945 (N_3945,N_3592,N_3537);
or U3946 (N_3946,N_3382,N_3364);
xor U3947 (N_3947,N_3277,N_3324);
nor U3948 (N_3948,N_3245,N_3211);
nor U3949 (N_3949,N_3400,N_3541);
xnor U3950 (N_3950,N_3394,N_3478);
or U3951 (N_3951,N_3340,N_3264);
xnor U3952 (N_3952,N_3544,N_3301);
and U3953 (N_3953,N_3477,N_3262);
and U3954 (N_3954,N_3357,N_3404);
and U3955 (N_3955,N_3217,N_3468);
nand U3956 (N_3956,N_3595,N_3281);
nor U3957 (N_3957,N_3504,N_3240);
nand U3958 (N_3958,N_3247,N_3545);
xnor U3959 (N_3959,N_3386,N_3329);
nor U3960 (N_3960,N_3240,N_3299);
xnor U3961 (N_3961,N_3486,N_3279);
nor U3962 (N_3962,N_3410,N_3590);
or U3963 (N_3963,N_3423,N_3447);
or U3964 (N_3964,N_3348,N_3206);
nor U3965 (N_3965,N_3592,N_3201);
nor U3966 (N_3966,N_3272,N_3425);
and U3967 (N_3967,N_3474,N_3337);
nor U3968 (N_3968,N_3541,N_3495);
xor U3969 (N_3969,N_3331,N_3404);
nand U3970 (N_3970,N_3493,N_3206);
xnor U3971 (N_3971,N_3226,N_3424);
nor U3972 (N_3972,N_3586,N_3397);
or U3973 (N_3973,N_3275,N_3283);
nand U3974 (N_3974,N_3560,N_3356);
or U3975 (N_3975,N_3457,N_3395);
and U3976 (N_3976,N_3396,N_3535);
nor U3977 (N_3977,N_3589,N_3414);
xor U3978 (N_3978,N_3375,N_3236);
xnor U3979 (N_3979,N_3407,N_3289);
nor U3980 (N_3980,N_3269,N_3276);
nor U3981 (N_3981,N_3497,N_3552);
nand U3982 (N_3982,N_3239,N_3405);
or U3983 (N_3983,N_3544,N_3499);
xor U3984 (N_3984,N_3318,N_3443);
nor U3985 (N_3985,N_3528,N_3367);
nand U3986 (N_3986,N_3522,N_3416);
xnor U3987 (N_3987,N_3493,N_3225);
and U3988 (N_3988,N_3364,N_3278);
nor U3989 (N_3989,N_3494,N_3288);
nor U3990 (N_3990,N_3432,N_3257);
xnor U3991 (N_3991,N_3305,N_3573);
nand U3992 (N_3992,N_3580,N_3565);
nand U3993 (N_3993,N_3290,N_3307);
or U3994 (N_3994,N_3331,N_3213);
and U3995 (N_3995,N_3538,N_3568);
and U3996 (N_3996,N_3534,N_3285);
xor U3997 (N_3997,N_3543,N_3406);
nor U3998 (N_3998,N_3291,N_3237);
and U3999 (N_3999,N_3589,N_3539);
and U4000 (N_4000,N_3740,N_3925);
nand U4001 (N_4001,N_3616,N_3812);
nor U4002 (N_4002,N_3663,N_3782);
or U4003 (N_4003,N_3694,N_3698);
xnor U4004 (N_4004,N_3672,N_3714);
nand U4005 (N_4005,N_3987,N_3828);
nand U4006 (N_4006,N_3945,N_3977);
nand U4007 (N_4007,N_3783,N_3781);
nand U4008 (N_4008,N_3708,N_3767);
nand U4009 (N_4009,N_3723,N_3742);
or U4010 (N_4010,N_3696,N_3879);
nor U4011 (N_4011,N_3825,N_3632);
nand U4012 (N_4012,N_3900,N_3736);
xor U4013 (N_4013,N_3950,N_3711);
nor U4014 (N_4014,N_3805,N_3936);
or U4015 (N_4015,N_3821,N_3756);
xnor U4016 (N_4016,N_3874,N_3615);
nor U4017 (N_4017,N_3791,N_3833);
xnor U4018 (N_4018,N_3610,N_3735);
nor U4019 (N_4019,N_3636,N_3885);
nor U4020 (N_4020,N_3707,N_3916);
xor U4021 (N_4021,N_3606,N_3892);
xor U4022 (N_4022,N_3769,N_3882);
xnor U4023 (N_4023,N_3932,N_3975);
xor U4024 (N_4024,N_3952,N_3854);
nor U4025 (N_4025,N_3989,N_3710);
xor U4026 (N_4026,N_3773,N_3832);
nand U4027 (N_4027,N_3751,N_3661);
and U4028 (N_4028,N_3691,N_3956);
and U4029 (N_4029,N_3968,N_3686);
xor U4030 (N_4030,N_3944,N_3884);
or U4031 (N_4031,N_3917,N_3820);
and U4032 (N_4032,N_3867,N_3847);
xnor U4033 (N_4033,N_3886,N_3704);
nor U4034 (N_4034,N_3701,N_3843);
nand U4035 (N_4035,N_3607,N_3969);
nor U4036 (N_4036,N_3953,N_3644);
and U4037 (N_4037,N_3753,N_3868);
nand U4038 (N_4038,N_3862,N_3901);
nor U4039 (N_4039,N_3961,N_3873);
or U4040 (N_4040,N_3613,N_3717);
and U4041 (N_4041,N_3739,N_3889);
and U4042 (N_4042,N_3846,N_3938);
nand U4043 (N_4043,N_3796,N_3991);
nand U4044 (N_4044,N_3729,N_3815);
xnor U4045 (N_4045,N_3934,N_3859);
and U4046 (N_4046,N_3979,N_3744);
xnor U4047 (N_4047,N_3904,N_3774);
nor U4048 (N_4048,N_3806,N_3699);
nand U4049 (N_4049,N_3721,N_3697);
nand U4050 (N_4050,N_3647,N_3864);
xor U4051 (N_4051,N_3972,N_3845);
or U4052 (N_4052,N_3660,N_3921);
nor U4053 (N_4053,N_3780,N_3706);
or U4054 (N_4054,N_3622,N_3920);
and U4055 (N_4055,N_3702,N_3871);
and U4056 (N_4056,N_3861,N_3662);
nand U4057 (N_4057,N_3899,N_3981);
and U4058 (N_4058,N_3928,N_3683);
or U4059 (N_4059,N_3974,N_3960);
and U4060 (N_4060,N_3824,N_3954);
xnor U4061 (N_4061,N_3652,N_3830);
and U4062 (N_4062,N_3638,N_3645);
and U4063 (N_4063,N_3999,N_3840);
xnor U4064 (N_4064,N_3687,N_3651);
nand U4065 (N_4065,N_3643,N_3911);
nand U4066 (N_4066,N_3878,N_3787);
nand U4067 (N_4067,N_3620,N_3967);
xor U4068 (N_4068,N_3988,N_3675);
nand U4069 (N_4069,N_3848,N_3748);
nand U4070 (N_4070,N_3640,N_3775);
and U4071 (N_4071,N_3619,N_3978);
and U4072 (N_4072,N_3665,N_3757);
nor U4073 (N_4073,N_3895,N_3658);
or U4074 (N_4074,N_3947,N_3724);
nor U4075 (N_4075,N_3865,N_3631);
nand U4076 (N_4076,N_3726,N_3679);
and U4077 (N_4077,N_3926,N_3997);
nand U4078 (N_4078,N_3754,N_3689);
nand U4079 (N_4079,N_3839,N_3604);
xor U4080 (N_4080,N_3678,N_3809);
and U4081 (N_4081,N_3800,N_3940);
nand U4082 (N_4082,N_3677,N_3994);
and U4083 (N_4083,N_3762,N_3628);
xnor U4084 (N_4084,N_3908,N_3746);
nand U4085 (N_4085,N_3693,N_3804);
and U4086 (N_4086,N_3627,N_3760);
or U4087 (N_4087,N_3849,N_3870);
or U4088 (N_4088,N_3692,N_3655);
and U4089 (N_4089,N_3603,N_3635);
and U4090 (N_4090,N_3747,N_3612);
and U4091 (N_4091,N_3887,N_3770);
and U4092 (N_4092,N_3629,N_3772);
nor U4093 (N_4093,N_3637,N_3819);
or U4094 (N_4094,N_3798,N_3690);
or U4095 (N_4095,N_3850,N_3803);
xor U4096 (N_4096,N_3778,N_3618);
or U4097 (N_4097,N_3958,N_3810);
or U4098 (N_4098,N_3793,N_3881);
or U4099 (N_4099,N_3785,N_3777);
nor U4100 (N_4100,N_3822,N_3984);
nor U4101 (N_4101,N_3814,N_3924);
nor U4102 (N_4102,N_3856,N_3933);
or U4103 (N_4103,N_3676,N_3688);
and U4104 (N_4104,N_3943,N_3722);
or U4105 (N_4105,N_3682,N_3712);
nor U4106 (N_4106,N_3851,N_3980);
or U4107 (N_4107,N_3869,N_3951);
xor U4108 (N_4108,N_3650,N_3919);
or U4109 (N_4109,N_3728,N_3937);
and U4110 (N_4110,N_3799,N_3903);
and U4111 (N_4111,N_3853,N_3835);
and U4112 (N_4112,N_3966,N_3811);
nor U4113 (N_4113,N_3674,N_3891);
or U4114 (N_4114,N_3836,N_3653);
xnor U4115 (N_4115,N_3641,N_3808);
or U4116 (N_4116,N_3971,N_3909);
xnor U4117 (N_4117,N_3858,N_3719);
xnor U4118 (N_4118,N_3755,N_3827);
or U4119 (N_4119,N_3654,N_3930);
nor U4120 (N_4120,N_3965,N_3976);
or U4121 (N_4121,N_3749,N_3709);
or U4122 (N_4122,N_3905,N_3941);
nor U4123 (N_4123,N_3703,N_3992);
nand U4124 (N_4124,N_3888,N_3818);
xor U4125 (N_4125,N_3964,N_3841);
nor U4126 (N_4126,N_3914,N_3982);
nand U4127 (N_4127,N_3970,N_3601);
xnor U4128 (N_4128,N_3877,N_3621);
xor U4129 (N_4129,N_3743,N_3996);
and U4130 (N_4130,N_3948,N_3838);
xor U4131 (N_4131,N_3718,N_3918);
nor U4132 (N_4132,N_3890,N_3670);
and U4133 (N_4133,N_3639,N_3893);
or U4134 (N_4134,N_3614,N_3779);
nand U4135 (N_4135,N_3831,N_3942);
xor U4136 (N_4136,N_3922,N_3912);
xor U4137 (N_4137,N_3725,N_3720);
nand U4138 (N_4138,N_3829,N_3759);
nor U4139 (N_4139,N_3957,N_3986);
nand U4140 (N_4140,N_3673,N_3750);
nand U4141 (N_4141,N_3765,N_3766);
and U4142 (N_4142,N_3605,N_3855);
nand U4143 (N_4143,N_3752,N_3656);
or U4144 (N_4144,N_3642,N_3741);
and U4145 (N_4145,N_3983,N_3897);
nor U4146 (N_4146,N_3801,N_3768);
nor U4147 (N_4147,N_3666,N_3738);
or U4148 (N_4148,N_3617,N_3931);
or U4149 (N_4149,N_3949,N_3648);
or U4150 (N_4150,N_3915,N_3737);
and U4151 (N_4151,N_3758,N_3705);
nor U4152 (N_4152,N_3913,N_3894);
nand U4153 (N_4153,N_3816,N_3667);
xor U4154 (N_4154,N_3863,N_3630);
nor U4155 (N_4155,N_3763,N_3876);
nor U4156 (N_4156,N_3633,N_3624);
and U4157 (N_4157,N_3985,N_3784);
xnor U4158 (N_4158,N_3962,N_3929);
nand U4159 (N_4159,N_3896,N_3802);
and U4160 (N_4160,N_3935,N_3727);
or U4161 (N_4161,N_3883,N_3764);
or U4162 (N_4162,N_3795,N_3713);
or U4163 (N_4163,N_3730,N_3734);
nor U4164 (N_4164,N_3646,N_3649);
nand U4165 (N_4165,N_3681,N_3963);
nand U4166 (N_4166,N_3625,N_3745);
and U4167 (N_4167,N_3837,N_3789);
xnor U4168 (N_4168,N_3866,N_3680);
and U4169 (N_4169,N_3844,N_3823);
or U4170 (N_4170,N_3995,N_3700);
or U4171 (N_4171,N_3813,N_3715);
nor U4172 (N_4172,N_3669,N_3955);
xnor U4173 (N_4173,N_3664,N_3716);
nor U4174 (N_4174,N_3990,N_3826);
and U4175 (N_4175,N_3685,N_3939);
and U4176 (N_4176,N_3608,N_3761);
and U4177 (N_4177,N_3790,N_3732);
xnor U4178 (N_4178,N_3733,N_3684);
xnor U4179 (N_4179,N_3852,N_3634);
xnor U4180 (N_4180,N_3910,N_3842);
nor U4181 (N_4181,N_3907,N_3797);
nor U4182 (N_4182,N_3834,N_3998);
xnor U4183 (N_4183,N_3659,N_3872);
xnor U4184 (N_4184,N_3898,N_3792);
nor U4185 (N_4185,N_3671,N_3973);
xor U4186 (N_4186,N_3626,N_3776);
and U4187 (N_4187,N_3609,N_3993);
xor U4188 (N_4188,N_3657,N_3771);
and U4189 (N_4189,N_3695,N_3923);
and U4190 (N_4190,N_3623,N_3902);
or U4191 (N_4191,N_3807,N_3875);
xnor U4192 (N_4192,N_3959,N_3602);
and U4193 (N_4193,N_3906,N_3731);
or U4194 (N_4194,N_3786,N_3794);
nor U4195 (N_4195,N_3668,N_3880);
nor U4196 (N_4196,N_3600,N_3788);
and U4197 (N_4197,N_3817,N_3860);
or U4198 (N_4198,N_3611,N_3927);
nand U4199 (N_4199,N_3857,N_3946);
nand U4200 (N_4200,N_3767,N_3918);
nor U4201 (N_4201,N_3873,N_3716);
and U4202 (N_4202,N_3802,N_3983);
and U4203 (N_4203,N_3857,N_3977);
nor U4204 (N_4204,N_3729,N_3753);
nand U4205 (N_4205,N_3954,N_3946);
nand U4206 (N_4206,N_3643,N_3738);
xor U4207 (N_4207,N_3803,N_3784);
xnor U4208 (N_4208,N_3602,N_3610);
and U4209 (N_4209,N_3867,N_3747);
and U4210 (N_4210,N_3606,N_3998);
or U4211 (N_4211,N_3922,N_3740);
or U4212 (N_4212,N_3810,N_3918);
nor U4213 (N_4213,N_3758,N_3637);
and U4214 (N_4214,N_3852,N_3643);
or U4215 (N_4215,N_3882,N_3941);
or U4216 (N_4216,N_3938,N_3759);
and U4217 (N_4217,N_3931,N_3895);
nor U4218 (N_4218,N_3888,N_3956);
and U4219 (N_4219,N_3901,N_3875);
nand U4220 (N_4220,N_3900,N_3785);
xnor U4221 (N_4221,N_3676,N_3722);
or U4222 (N_4222,N_3711,N_3999);
nand U4223 (N_4223,N_3891,N_3772);
xnor U4224 (N_4224,N_3788,N_3921);
nand U4225 (N_4225,N_3722,N_3635);
and U4226 (N_4226,N_3771,N_3628);
or U4227 (N_4227,N_3644,N_3715);
xnor U4228 (N_4228,N_3862,N_3954);
and U4229 (N_4229,N_3752,N_3877);
and U4230 (N_4230,N_3950,N_3854);
and U4231 (N_4231,N_3965,N_3651);
nand U4232 (N_4232,N_3987,N_3871);
or U4233 (N_4233,N_3652,N_3852);
xor U4234 (N_4234,N_3686,N_3825);
nand U4235 (N_4235,N_3923,N_3979);
nor U4236 (N_4236,N_3993,N_3956);
nor U4237 (N_4237,N_3820,N_3719);
or U4238 (N_4238,N_3879,N_3969);
and U4239 (N_4239,N_3938,N_3620);
and U4240 (N_4240,N_3774,N_3721);
and U4241 (N_4241,N_3659,N_3645);
or U4242 (N_4242,N_3898,N_3625);
nand U4243 (N_4243,N_3690,N_3867);
nor U4244 (N_4244,N_3919,N_3971);
nor U4245 (N_4245,N_3656,N_3865);
xnor U4246 (N_4246,N_3940,N_3658);
and U4247 (N_4247,N_3990,N_3921);
nor U4248 (N_4248,N_3623,N_3905);
nand U4249 (N_4249,N_3807,N_3730);
or U4250 (N_4250,N_3826,N_3900);
xnor U4251 (N_4251,N_3869,N_3913);
and U4252 (N_4252,N_3883,N_3775);
nand U4253 (N_4253,N_3624,N_3815);
and U4254 (N_4254,N_3656,N_3947);
nand U4255 (N_4255,N_3944,N_3992);
nor U4256 (N_4256,N_3882,N_3984);
and U4257 (N_4257,N_3645,N_3662);
nand U4258 (N_4258,N_3700,N_3921);
xnor U4259 (N_4259,N_3740,N_3608);
and U4260 (N_4260,N_3634,N_3834);
or U4261 (N_4261,N_3635,N_3690);
nand U4262 (N_4262,N_3685,N_3893);
or U4263 (N_4263,N_3769,N_3696);
and U4264 (N_4264,N_3906,N_3983);
nor U4265 (N_4265,N_3854,N_3786);
nand U4266 (N_4266,N_3986,N_3843);
nor U4267 (N_4267,N_3700,N_3803);
nand U4268 (N_4268,N_3645,N_3739);
nor U4269 (N_4269,N_3979,N_3894);
xnor U4270 (N_4270,N_3731,N_3665);
xnor U4271 (N_4271,N_3748,N_3804);
xor U4272 (N_4272,N_3706,N_3731);
xor U4273 (N_4273,N_3743,N_3769);
nor U4274 (N_4274,N_3701,N_3667);
xnor U4275 (N_4275,N_3613,N_3658);
or U4276 (N_4276,N_3851,N_3660);
xor U4277 (N_4277,N_3939,N_3795);
or U4278 (N_4278,N_3632,N_3622);
xor U4279 (N_4279,N_3797,N_3836);
and U4280 (N_4280,N_3912,N_3955);
xor U4281 (N_4281,N_3669,N_3708);
xnor U4282 (N_4282,N_3678,N_3836);
and U4283 (N_4283,N_3641,N_3670);
nor U4284 (N_4284,N_3787,N_3908);
nand U4285 (N_4285,N_3833,N_3769);
and U4286 (N_4286,N_3784,N_3742);
xor U4287 (N_4287,N_3714,N_3740);
nand U4288 (N_4288,N_3883,N_3840);
or U4289 (N_4289,N_3807,N_3861);
nand U4290 (N_4290,N_3970,N_3933);
or U4291 (N_4291,N_3774,N_3696);
and U4292 (N_4292,N_3912,N_3987);
xor U4293 (N_4293,N_3671,N_3636);
or U4294 (N_4294,N_3706,N_3955);
nand U4295 (N_4295,N_3914,N_3732);
and U4296 (N_4296,N_3676,N_3689);
or U4297 (N_4297,N_3978,N_3667);
nand U4298 (N_4298,N_3752,N_3946);
xor U4299 (N_4299,N_3937,N_3663);
nor U4300 (N_4300,N_3649,N_3822);
and U4301 (N_4301,N_3753,N_3759);
nor U4302 (N_4302,N_3808,N_3959);
nand U4303 (N_4303,N_3799,N_3909);
or U4304 (N_4304,N_3869,N_3917);
nor U4305 (N_4305,N_3773,N_3847);
nand U4306 (N_4306,N_3866,N_3920);
xnor U4307 (N_4307,N_3856,N_3746);
nor U4308 (N_4308,N_3795,N_3673);
and U4309 (N_4309,N_3742,N_3801);
nand U4310 (N_4310,N_3743,N_3944);
nand U4311 (N_4311,N_3880,N_3828);
nand U4312 (N_4312,N_3954,N_3916);
nor U4313 (N_4313,N_3668,N_3915);
or U4314 (N_4314,N_3999,N_3824);
or U4315 (N_4315,N_3655,N_3768);
xor U4316 (N_4316,N_3905,N_3664);
xnor U4317 (N_4317,N_3914,N_3740);
nand U4318 (N_4318,N_3944,N_3667);
nand U4319 (N_4319,N_3905,N_3717);
and U4320 (N_4320,N_3874,N_3649);
xor U4321 (N_4321,N_3709,N_3780);
and U4322 (N_4322,N_3657,N_3979);
and U4323 (N_4323,N_3787,N_3954);
xor U4324 (N_4324,N_3677,N_3879);
or U4325 (N_4325,N_3780,N_3769);
nor U4326 (N_4326,N_3978,N_3604);
or U4327 (N_4327,N_3914,N_3639);
nor U4328 (N_4328,N_3879,N_3767);
nor U4329 (N_4329,N_3976,N_3848);
or U4330 (N_4330,N_3848,N_3741);
or U4331 (N_4331,N_3631,N_3811);
nand U4332 (N_4332,N_3855,N_3901);
or U4333 (N_4333,N_3834,N_3896);
and U4334 (N_4334,N_3809,N_3663);
nor U4335 (N_4335,N_3606,N_3796);
nor U4336 (N_4336,N_3880,N_3817);
xnor U4337 (N_4337,N_3959,N_3749);
or U4338 (N_4338,N_3634,N_3716);
nand U4339 (N_4339,N_3845,N_3663);
xor U4340 (N_4340,N_3826,N_3607);
nor U4341 (N_4341,N_3706,N_3879);
or U4342 (N_4342,N_3769,N_3879);
and U4343 (N_4343,N_3994,N_3649);
nand U4344 (N_4344,N_3668,N_3698);
xnor U4345 (N_4345,N_3954,N_3897);
nand U4346 (N_4346,N_3869,N_3859);
nor U4347 (N_4347,N_3700,N_3645);
or U4348 (N_4348,N_3934,N_3809);
or U4349 (N_4349,N_3910,N_3818);
or U4350 (N_4350,N_3771,N_3703);
xnor U4351 (N_4351,N_3898,N_3751);
and U4352 (N_4352,N_3851,N_3652);
nand U4353 (N_4353,N_3833,N_3795);
xor U4354 (N_4354,N_3770,N_3882);
or U4355 (N_4355,N_3956,N_3647);
nor U4356 (N_4356,N_3885,N_3720);
nand U4357 (N_4357,N_3615,N_3728);
or U4358 (N_4358,N_3607,N_3723);
xor U4359 (N_4359,N_3976,N_3752);
xnor U4360 (N_4360,N_3726,N_3994);
nor U4361 (N_4361,N_3654,N_3899);
or U4362 (N_4362,N_3812,N_3729);
nor U4363 (N_4363,N_3663,N_3707);
xor U4364 (N_4364,N_3947,N_3948);
xnor U4365 (N_4365,N_3823,N_3825);
xnor U4366 (N_4366,N_3800,N_3970);
nor U4367 (N_4367,N_3855,N_3759);
nor U4368 (N_4368,N_3914,N_3638);
xor U4369 (N_4369,N_3854,N_3974);
nor U4370 (N_4370,N_3770,N_3909);
nor U4371 (N_4371,N_3919,N_3644);
xor U4372 (N_4372,N_3663,N_3873);
nand U4373 (N_4373,N_3825,N_3973);
nand U4374 (N_4374,N_3665,N_3717);
nand U4375 (N_4375,N_3740,N_3721);
nor U4376 (N_4376,N_3676,N_3681);
nand U4377 (N_4377,N_3660,N_3941);
xnor U4378 (N_4378,N_3695,N_3977);
nand U4379 (N_4379,N_3651,N_3731);
xnor U4380 (N_4380,N_3920,N_3838);
or U4381 (N_4381,N_3860,N_3805);
or U4382 (N_4382,N_3924,N_3602);
or U4383 (N_4383,N_3639,N_3798);
and U4384 (N_4384,N_3640,N_3941);
or U4385 (N_4385,N_3830,N_3992);
and U4386 (N_4386,N_3859,N_3819);
nor U4387 (N_4387,N_3660,N_3995);
nand U4388 (N_4388,N_3804,N_3683);
nand U4389 (N_4389,N_3895,N_3676);
xor U4390 (N_4390,N_3943,N_3614);
and U4391 (N_4391,N_3667,N_3728);
xor U4392 (N_4392,N_3766,N_3809);
nor U4393 (N_4393,N_3976,N_3637);
xor U4394 (N_4394,N_3895,N_3608);
or U4395 (N_4395,N_3853,N_3874);
nor U4396 (N_4396,N_3618,N_3845);
xnor U4397 (N_4397,N_3717,N_3957);
nor U4398 (N_4398,N_3851,N_3623);
nand U4399 (N_4399,N_3993,N_3963);
xnor U4400 (N_4400,N_4223,N_4270);
nor U4401 (N_4401,N_4238,N_4128);
nand U4402 (N_4402,N_4379,N_4289);
nor U4403 (N_4403,N_4229,N_4315);
nor U4404 (N_4404,N_4393,N_4391);
and U4405 (N_4405,N_4095,N_4222);
xnor U4406 (N_4406,N_4039,N_4085);
or U4407 (N_4407,N_4332,N_4213);
xnor U4408 (N_4408,N_4299,N_4322);
nor U4409 (N_4409,N_4247,N_4338);
nand U4410 (N_4410,N_4250,N_4044);
xnor U4411 (N_4411,N_4113,N_4127);
xor U4412 (N_4412,N_4178,N_4145);
xnor U4413 (N_4413,N_4397,N_4183);
xor U4414 (N_4414,N_4094,N_4370);
nand U4415 (N_4415,N_4168,N_4045);
nand U4416 (N_4416,N_4252,N_4034);
or U4417 (N_4417,N_4186,N_4268);
or U4418 (N_4418,N_4243,N_4233);
and U4419 (N_4419,N_4033,N_4376);
or U4420 (N_4420,N_4217,N_4021);
xnor U4421 (N_4421,N_4240,N_4333);
and U4422 (N_4422,N_4148,N_4203);
xnor U4423 (N_4423,N_4334,N_4141);
or U4424 (N_4424,N_4142,N_4272);
nor U4425 (N_4425,N_4019,N_4116);
or U4426 (N_4426,N_4262,N_4326);
nand U4427 (N_4427,N_4339,N_4149);
nor U4428 (N_4428,N_4248,N_4392);
xnor U4429 (N_4429,N_4080,N_4253);
nand U4430 (N_4430,N_4235,N_4308);
nor U4431 (N_4431,N_4353,N_4239);
xor U4432 (N_4432,N_4209,N_4053);
nor U4433 (N_4433,N_4181,N_4138);
nand U4434 (N_4434,N_4271,N_4121);
or U4435 (N_4435,N_4016,N_4398);
and U4436 (N_4436,N_4193,N_4263);
or U4437 (N_4437,N_4096,N_4088);
and U4438 (N_4438,N_4241,N_4075);
nor U4439 (N_4439,N_4010,N_4300);
xnor U4440 (N_4440,N_4295,N_4329);
nor U4441 (N_4441,N_4067,N_4399);
nor U4442 (N_4442,N_4356,N_4109);
or U4443 (N_4443,N_4182,N_4218);
or U4444 (N_4444,N_4390,N_4364);
nand U4445 (N_4445,N_4294,N_4012);
xor U4446 (N_4446,N_4282,N_4082);
nor U4447 (N_4447,N_4154,N_4389);
or U4448 (N_4448,N_4062,N_4291);
nand U4449 (N_4449,N_4003,N_4144);
nand U4450 (N_4450,N_4384,N_4107);
nor U4451 (N_4451,N_4216,N_4171);
xnor U4452 (N_4452,N_4074,N_4279);
xnor U4453 (N_4453,N_4157,N_4265);
xnor U4454 (N_4454,N_4049,N_4084);
and U4455 (N_4455,N_4340,N_4172);
nand U4456 (N_4456,N_4076,N_4207);
or U4457 (N_4457,N_4023,N_4382);
xor U4458 (N_4458,N_4320,N_4038);
and U4459 (N_4459,N_4132,N_4347);
and U4460 (N_4460,N_4006,N_4395);
xnor U4461 (N_4461,N_4285,N_4007);
or U4462 (N_4462,N_4324,N_4287);
nand U4463 (N_4463,N_4026,N_4114);
nand U4464 (N_4464,N_4000,N_4350);
nor U4465 (N_4465,N_4345,N_4052);
or U4466 (N_4466,N_4120,N_4072);
nand U4467 (N_4467,N_4343,N_4115);
xnor U4468 (N_4468,N_4099,N_4331);
or U4469 (N_4469,N_4090,N_4337);
and U4470 (N_4470,N_4089,N_4314);
xor U4471 (N_4471,N_4081,N_4009);
nor U4472 (N_4472,N_4043,N_4064);
xor U4473 (N_4473,N_4086,N_4255);
and U4474 (N_4474,N_4002,N_4312);
nor U4475 (N_4475,N_4208,N_4274);
nand U4476 (N_4476,N_4280,N_4360);
nand U4477 (N_4477,N_4122,N_4221);
xnor U4478 (N_4478,N_4042,N_4169);
or U4479 (N_4479,N_4079,N_4231);
or U4480 (N_4480,N_4134,N_4219);
or U4481 (N_4481,N_4131,N_4202);
nor U4482 (N_4482,N_4244,N_4123);
nand U4483 (N_4483,N_4194,N_4143);
nand U4484 (N_4484,N_4078,N_4355);
nand U4485 (N_4485,N_4286,N_4147);
nor U4486 (N_4486,N_4166,N_4112);
nand U4487 (N_4487,N_4190,N_4199);
and U4488 (N_4488,N_4028,N_4097);
and U4489 (N_4489,N_4001,N_4319);
nand U4490 (N_4490,N_4210,N_4346);
nand U4491 (N_4491,N_4187,N_4302);
or U4492 (N_4492,N_4054,N_4377);
and U4493 (N_4493,N_4069,N_4325);
nor U4494 (N_4494,N_4290,N_4163);
xnor U4495 (N_4495,N_4108,N_4066);
or U4496 (N_4496,N_4179,N_4191);
or U4497 (N_4497,N_4125,N_4124);
nand U4498 (N_4498,N_4091,N_4386);
nor U4499 (N_4499,N_4254,N_4304);
or U4500 (N_4500,N_4361,N_4301);
xnor U4501 (N_4501,N_4024,N_4373);
nor U4502 (N_4502,N_4071,N_4351);
xnor U4503 (N_4503,N_4061,N_4160);
or U4504 (N_4504,N_4206,N_4046);
and U4505 (N_4505,N_4135,N_4103);
nor U4506 (N_4506,N_4011,N_4365);
nand U4507 (N_4507,N_4368,N_4032);
nor U4508 (N_4508,N_4111,N_4242);
or U4509 (N_4509,N_4344,N_4256);
nand U4510 (N_4510,N_4381,N_4152);
and U4511 (N_4511,N_4318,N_4087);
nand U4512 (N_4512,N_4110,N_4065);
nand U4513 (N_4513,N_4167,N_4305);
xor U4514 (N_4514,N_4330,N_4374);
nand U4515 (N_4515,N_4060,N_4059);
or U4516 (N_4516,N_4129,N_4165);
nand U4517 (N_4517,N_4378,N_4161);
or U4518 (N_4518,N_4195,N_4246);
or U4519 (N_4519,N_4278,N_4041);
xor U4520 (N_4520,N_4215,N_4375);
and U4521 (N_4521,N_4101,N_4245);
xnor U4522 (N_4522,N_4047,N_4269);
and U4523 (N_4523,N_4303,N_4385);
or U4524 (N_4524,N_4335,N_4357);
nor U4525 (N_4525,N_4232,N_4146);
xnor U4526 (N_4526,N_4212,N_4328);
nand U4527 (N_4527,N_4098,N_4017);
xnor U4528 (N_4528,N_4366,N_4159);
nor U4529 (N_4529,N_4077,N_4236);
nor U4530 (N_4530,N_4055,N_4174);
xnor U4531 (N_4531,N_4180,N_4175);
xor U4532 (N_4532,N_4369,N_4133);
xnor U4533 (N_4533,N_4100,N_4367);
xnor U4534 (N_4534,N_4197,N_4352);
nor U4535 (N_4535,N_4383,N_4018);
nor U4536 (N_4536,N_4068,N_4293);
or U4537 (N_4537,N_4056,N_4192);
or U4538 (N_4538,N_4310,N_4237);
xnor U4539 (N_4539,N_4226,N_4029);
nand U4540 (N_4540,N_4025,N_4104);
xnor U4541 (N_4541,N_4057,N_4030);
or U4542 (N_4542,N_4092,N_4119);
and U4543 (N_4543,N_4297,N_4150);
and U4544 (N_4544,N_4048,N_4258);
nor U4545 (N_4545,N_4266,N_4151);
nor U4546 (N_4546,N_4380,N_4277);
and U4547 (N_4547,N_4083,N_4189);
nand U4548 (N_4548,N_4249,N_4176);
nand U4549 (N_4549,N_4372,N_4118);
nand U4550 (N_4550,N_4227,N_4275);
xor U4551 (N_4551,N_4284,N_4220);
nor U4552 (N_4552,N_4309,N_4014);
xnor U4553 (N_4553,N_4158,N_4396);
and U4554 (N_4554,N_4363,N_4117);
nor U4555 (N_4555,N_4214,N_4153);
or U4556 (N_4556,N_4204,N_4008);
or U4557 (N_4557,N_4020,N_4257);
and U4558 (N_4558,N_4205,N_4273);
nand U4559 (N_4559,N_4311,N_4281);
nor U4560 (N_4560,N_4225,N_4070);
xor U4561 (N_4561,N_4316,N_4349);
xor U4562 (N_4562,N_4261,N_4102);
nor U4563 (N_4563,N_4040,N_4198);
xnor U4564 (N_4564,N_4251,N_4185);
nor U4565 (N_4565,N_4387,N_4177);
or U4566 (N_4566,N_4359,N_4354);
nor U4567 (N_4567,N_4105,N_4296);
and U4568 (N_4568,N_4276,N_4234);
or U4569 (N_4569,N_4317,N_4200);
and U4570 (N_4570,N_4307,N_4037);
xnor U4571 (N_4571,N_4036,N_4005);
nor U4572 (N_4572,N_4288,N_4031);
nor U4573 (N_4573,N_4050,N_4358);
nor U4574 (N_4574,N_4156,N_4298);
or U4575 (N_4575,N_4371,N_4348);
xor U4576 (N_4576,N_4267,N_4292);
nand U4577 (N_4577,N_4162,N_4015);
nor U4578 (N_4578,N_4211,N_4362);
xor U4579 (N_4579,N_4130,N_4184);
nand U4580 (N_4580,N_4224,N_4228);
nand U4581 (N_4581,N_4137,N_4260);
or U4582 (N_4582,N_4164,N_4058);
xnor U4583 (N_4583,N_4013,N_4259);
nand U4584 (N_4584,N_4139,N_4196);
and U4585 (N_4585,N_4035,N_4341);
or U4586 (N_4586,N_4027,N_4004);
and U4587 (N_4587,N_4394,N_4306);
xor U4588 (N_4588,N_4323,N_4140);
or U4589 (N_4589,N_4051,N_4170);
nor U4590 (N_4590,N_4126,N_4022);
nand U4591 (N_4591,N_4264,N_4321);
xor U4592 (N_4592,N_4342,N_4327);
nand U4593 (N_4593,N_4201,N_4313);
nand U4594 (N_4594,N_4173,N_4283);
nor U4595 (N_4595,N_4230,N_4155);
and U4596 (N_4596,N_4093,N_4063);
or U4597 (N_4597,N_4136,N_4073);
and U4598 (N_4598,N_4388,N_4106);
and U4599 (N_4599,N_4188,N_4336);
nor U4600 (N_4600,N_4075,N_4211);
or U4601 (N_4601,N_4287,N_4254);
nor U4602 (N_4602,N_4155,N_4120);
or U4603 (N_4603,N_4219,N_4018);
nand U4604 (N_4604,N_4168,N_4103);
or U4605 (N_4605,N_4061,N_4303);
and U4606 (N_4606,N_4241,N_4064);
or U4607 (N_4607,N_4220,N_4257);
xor U4608 (N_4608,N_4296,N_4027);
nor U4609 (N_4609,N_4273,N_4347);
xnor U4610 (N_4610,N_4189,N_4055);
and U4611 (N_4611,N_4282,N_4312);
and U4612 (N_4612,N_4171,N_4083);
and U4613 (N_4613,N_4059,N_4213);
nand U4614 (N_4614,N_4169,N_4226);
xnor U4615 (N_4615,N_4126,N_4016);
or U4616 (N_4616,N_4155,N_4103);
nand U4617 (N_4617,N_4380,N_4232);
and U4618 (N_4618,N_4162,N_4098);
and U4619 (N_4619,N_4384,N_4002);
nand U4620 (N_4620,N_4254,N_4031);
xor U4621 (N_4621,N_4143,N_4314);
nor U4622 (N_4622,N_4323,N_4136);
xor U4623 (N_4623,N_4028,N_4084);
nand U4624 (N_4624,N_4075,N_4109);
or U4625 (N_4625,N_4319,N_4209);
or U4626 (N_4626,N_4134,N_4012);
nand U4627 (N_4627,N_4323,N_4237);
and U4628 (N_4628,N_4392,N_4006);
nor U4629 (N_4629,N_4332,N_4387);
nor U4630 (N_4630,N_4398,N_4165);
or U4631 (N_4631,N_4042,N_4105);
xnor U4632 (N_4632,N_4064,N_4306);
nor U4633 (N_4633,N_4140,N_4302);
xnor U4634 (N_4634,N_4381,N_4347);
nand U4635 (N_4635,N_4016,N_4212);
and U4636 (N_4636,N_4248,N_4124);
or U4637 (N_4637,N_4319,N_4000);
and U4638 (N_4638,N_4331,N_4027);
or U4639 (N_4639,N_4229,N_4237);
nand U4640 (N_4640,N_4271,N_4274);
nand U4641 (N_4641,N_4216,N_4385);
nor U4642 (N_4642,N_4355,N_4385);
and U4643 (N_4643,N_4291,N_4265);
xor U4644 (N_4644,N_4380,N_4061);
nor U4645 (N_4645,N_4291,N_4184);
and U4646 (N_4646,N_4028,N_4313);
and U4647 (N_4647,N_4108,N_4358);
xor U4648 (N_4648,N_4253,N_4374);
and U4649 (N_4649,N_4327,N_4091);
or U4650 (N_4650,N_4318,N_4377);
nand U4651 (N_4651,N_4002,N_4215);
xnor U4652 (N_4652,N_4304,N_4344);
nor U4653 (N_4653,N_4189,N_4336);
xnor U4654 (N_4654,N_4330,N_4149);
and U4655 (N_4655,N_4286,N_4353);
nor U4656 (N_4656,N_4115,N_4255);
xnor U4657 (N_4657,N_4395,N_4060);
or U4658 (N_4658,N_4371,N_4235);
and U4659 (N_4659,N_4390,N_4372);
or U4660 (N_4660,N_4130,N_4215);
or U4661 (N_4661,N_4372,N_4333);
nor U4662 (N_4662,N_4016,N_4115);
nor U4663 (N_4663,N_4382,N_4042);
nor U4664 (N_4664,N_4217,N_4189);
nand U4665 (N_4665,N_4055,N_4383);
xor U4666 (N_4666,N_4345,N_4355);
xnor U4667 (N_4667,N_4297,N_4219);
nand U4668 (N_4668,N_4385,N_4376);
and U4669 (N_4669,N_4384,N_4305);
nand U4670 (N_4670,N_4236,N_4357);
or U4671 (N_4671,N_4166,N_4190);
or U4672 (N_4672,N_4143,N_4175);
nand U4673 (N_4673,N_4224,N_4394);
or U4674 (N_4674,N_4258,N_4332);
or U4675 (N_4675,N_4102,N_4199);
nand U4676 (N_4676,N_4366,N_4261);
nor U4677 (N_4677,N_4109,N_4085);
nand U4678 (N_4678,N_4078,N_4242);
xor U4679 (N_4679,N_4180,N_4308);
and U4680 (N_4680,N_4301,N_4026);
xnor U4681 (N_4681,N_4086,N_4076);
xor U4682 (N_4682,N_4318,N_4037);
and U4683 (N_4683,N_4140,N_4124);
nand U4684 (N_4684,N_4057,N_4326);
nand U4685 (N_4685,N_4144,N_4336);
or U4686 (N_4686,N_4068,N_4326);
nand U4687 (N_4687,N_4173,N_4115);
and U4688 (N_4688,N_4117,N_4045);
or U4689 (N_4689,N_4394,N_4061);
or U4690 (N_4690,N_4012,N_4266);
nor U4691 (N_4691,N_4058,N_4136);
nand U4692 (N_4692,N_4353,N_4168);
nand U4693 (N_4693,N_4230,N_4187);
or U4694 (N_4694,N_4293,N_4045);
or U4695 (N_4695,N_4273,N_4341);
nand U4696 (N_4696,N_4161,N_4062);
xor U4697 (N_4697,N_4185,N_4392);
and U4698 (N_4698,N_4054,N_4361);
and U4699 (N_4699,N_4244,N_4192);
xnor U4700 (N_4700,N_4050,N_4161);
nor U4701 (N_4701,N_4330,N_4365);
and U4702 (N_4702,N_4016,N_4342);
nor U4703 (N_4703,N_4036,N_4350);
nor U4704 (N_4704,N_4126,N_4391);
or U4705 (N_4705,N_4082,N_4197);
xor U4706 (N_4706,N_4337,N_4012);
nand U4707 (N_4707,N_4328,N_4153);
nor U4708 (N_4708,N_4051,N_4227);
or U4709 (N_4709,N_4049,N_4359);
nor U4710 (N_4710,N_4023,N_4133);
xnor U4711 (N_4711,N_4227,N_4297);
nand U4712 (N_4712,N_4067,N_4217);
nor U4713 (N_4713,N_4110,N_4213);
or U4714 (N_4714,N_4178,N_4300);
or U4715 (N_4715,N_4015,N_4147);
and U4716 (N_4716,N_4336,N_4102);
and U4717 (N_4717,N_4157,N_4203);
nor U4718 (N_4718,N_4041,N_4241);
and U4719 (N_4719,N_4379,N_4114);
xor U4720 (N_4720,N_4274,N_4088);
or U4721 (N_4721,N_4299,N_4197);
or U4722 (N_4722,N_4173,N_4084);
or U4723 (N_4723,N_4294,N_4337);
xor U4724 (N_4724,N_4198,N_4136);
nor U4725 (N_4725,N_4208,N_4199);
nor U4726 (N_4726,N_4206,N_4184);
nor U4727 (N_4727,N_4180,N_4154);
and U4728 (N_4728,N_4312,N_4059);
nand U4729 (N_4729,N_4310,N_4001);
xnor U4730 (N_4730,N_4064,N_4187);
and U4731 (N_4731,N_4148,N_4174);
and U4732 (N_4732,N_4110,N_4178);
and U4733 (N_4733,N_4175,N_4281);
and U4734 (N_4734,N_4230,N_4026);
and U4735 (N_4735,N_4310,N_4085);
or U4736 (N_4736,N_4293,N_4372);
xnor U4737 (N_4737,N_4072,N_4152);
and U4738 (N_4738,N_4240,N_4326);
nor U4739 (N_4739,N_4206,N_4298);
nor U4740 (N_4740,N_4255,N_4347);
xor U4741 (N_4741,N_4358,N_4248);
and U4742 (N_4742,N_4206,N_4176);
and U4743 (N_4743,N_4387,N_4287);
xnor U4744 (N_4744,N_4109,N_4282);
xnor U4745 (N_4745,N_4092,N_4318);
and U4746 (N_4746,N_4197,N_4237);
nor U4747 (N_4747,N_4066,N_4251);
xnor U4748 (N_4748,N_4169,N_4005);
xor U4749 (N_4749,N_4160,N_4174);
and U4750 (N_4750,N_4085,N_4191);
or U4751 (N_4751,N_4142,N_4009);
or U4752 (N_4752,N_4041,N_4222);
or U4753 (N_4753,N_4165,N_4177);
nor U4754 (N_4754,N_4236,N_4071);
and U4755 (N_4755,N_4238,N_4186);
nand U4756 (N_4756,N_4161,N_4294);
nand U4757 (N_4757,N_4000,N_4013);
and U4758 (N_4758,N_4399,N_4347);
and U4759 (N_4759,N_4174,N_4188);
or U4760 (N_4760,N_4191,N_4164);
nor U4761 (N_4761,N_4036,N_4171);
xor U4762 (N_4762,N_4235,N_4134);
and U4763 (N_4763,N_4103,N_4392);
and U4764 (N_4764,N_4388,N_4337);
and U4765 (N_4765,N_4184,N_4101);
xor U4766 (N_4766,N_4010,N_4347);
nor U4767 (N_4767,N_4065,N_4191);
or U4768 (N_4768,N_4192,N_4317);
xor U4769 (N_4769,N_4143,N_4376);
nand U4770 (N_4770,N_4323,N_4041);
or U4771 (N_4771,N_4027,N_4375);
nor U4772 (N_4772,N_4195,N_4141);
or U4773 (N_4773,N_4033,N_4001);
and U4774 (N_4774,N_4148,N_4275);
or U4775 (N_4775,N_4094,N_4325);
and U4776 (N_4776,N_4040,N_4268);
nand U4777 (N_4777,N_4125,N_4000);
xor U4778 (N_4778,N_4056,N_4184);
nand U4779 (N_4779,N_4143,N_4154);
xor U4780 (N_4780,N_4099,N_4283);
nand U4781 (N_4781,N_4205,N_4233);
xor U4782 (N_4782,N_4352,N_4252);
and U4783 (N_4783,N_4365,N_4096);
nor U4784 (N_4784,N_4052,N_4149);
and U4785 (N_4785,N_4394,N_4229);
nor U4786 (N_4786,N_4165,N_4046);
nor U4787 (N_4787,N_4264,N_4368);
nand U4788 (N_4788,N_4351,N_4318);
xor U4789 (N_4789,N_4311,N_4105);
and U4790 (N_4790,N_4202,N_4274);
nor U4791 (N_4791,N_4251,N_4353);
nor U4792 (N_4792,N_4102,N_4200);
and U4793 (N_4793,N_4005,N_4060);
xor U4794 (N_4794,N_4098,N_4072);
xor U4795 (N_4795,N_4247,N_4186);
nor U4796 (N_4796,N_4186,N_4291);
or U4797 (N_4797,N_4094,N_4228);
and U4798 (N_4798,N_4142,N_4049);
xnor U4799 (N_4799,N_4287,N_4285);
and U4800 (N_4800,N_4496,N_4562);
nor U4801 (N_4801,N_4466,N_4481);
and U4802 (N_4802,N_4548,N_4634);
nor U4803 (N_4803,N_4565,N_4546);
nand U4804 (N_4804,N_4514,N_4429);
nor U4805 (N_4805,N_4601,N_4411);
nand U4806 (N_4806,N_4589,N_4604);
or U4807 (N_4807,N_4662,N_4799);
or U4808 (N_4808,N_4409,N_4449);
nand U4809 (N_4809,N_4478,N_4573);
and U4810 (N_4810,N_4581,N_4720);
nand U4811 (N_4811,N_4443,N_4650);
nand U4812 (N_4812,N_4733,N_4461);
nor U4813 (N_4813,N_4760,N_4682);
nor U4814 (N_4814,N_4557,N_4631);
and U4815 (N_4815,N_4757,N_4642);
nand U4816 (N_4816,N_4783,N_4564);
xnor U4817 (N_4817,N_4651,N_4453);
or U4818 (N_4818,N_4539,N_4714);
or U4819 (N_4819,N_4612,N_4775);
nor U4820 (N_4820,N_4521,N_4704);
or U4821 (N_4821,N_4438,N_4495);
or U4822 (N_4822,N_4587,N_4559);
nor U4823 (N_4823,N_4415,N_4728);
nor U4824 (N_4824,N_4743,N_4763);
nand U4825 (N_4825,N_4724,N_4554);
and U4826 (N_4826,N_4759,N_4576);
nand U4827 (N_4827,N_4540,N_4505);
or U4828 (N_4828,N_4476,N_4711);
nand U4829 (N_4829,N_4566,N_4645);
or U4830 (N_4830,N_4499,N_4452);
nand U4831 (N_4831,N_4717,N_4652);
nand U4832 (N_4832,N_4590,N_4709);
or U4833 (N_4833,N_4598,N_4765);
or U4834 (N_4834,N_4406,N_4713);
or U4835 (N_4835,N_4518,N_4686);
nor U4836 (N_4836,N_4700,N_4427);
nor U4837 (N_4837,N_4618,N_4577);
nand U4838 (N_4838,N_4440,N_4542);
or U4839 (N_4839,N_4788,N_4431);
or U4840 (N_4840,N_4501,N_4517);
or U4841 (N_4841,N_4571,N_4699);
or U4842 (N_4842,N_4669,N_4663);
xnor U4843 (N_4843,N_4718,N_4430);
xnor U4844 (N_4844,N_4653,N_4485);
and U4845 (N_4845,N_4472,N_4617);
nand U4846 (N_4846,N_4417,N_4660);
and U4847 (N_4847,N_4616,N_4607);
xor U4848 (N_4848,N_4531,N_4677);
and U4849 (N_4849,N_4420,N_4407);
nor U4850 (N_4850,N_4667,N_4639);
nor U4851 (N_4851,N_4730,N_4405);
xnor U4852 (N_4852,N_4796,N_4620);
or U4853 (N_4853,N_4769,N_4413);
nor U4854 (N_4854,N_4551,N_4640);
nand U4855 (N_4855,N_4649,N_4490);
nor U4856 (N_4856,N_4793,N_4786);
or U4857 (N_4857,N_4725,N_4456);
and U4858 (N_4858,N_4585,N_4544);
nor U4859 (N_4859,N_4568,N_4575);
xor U4860 (N_4860,N_4673,N_4526);
and U4861 (N_4861,N_4421,N_4648);
xnor U4862 (N_4862,N_4690,N_4753);
xnor U4863 (N_4863,N_4668,N_4722);
or U4864 (N_4864,N_4735,N_4402);
or U4865 (N_4865,N_4549,N_4547);
nor U4866 (N_4866,N_4470,N_4614);
xnor U4867 (N_4867,N_4696,N_4458);
nor U4868 (N_4868,N_4474,N_4468);
nand U4869 (N_4869,N_4570,N_4615);
nand U4870 (N_4870,N_4644,N_4770);
and U4871 (N_4871,N_4777,N_4408);
and U4872 (N_4872,N_4773,N_4630);
nor U4873 (N_4873,N_4567,N_4675);
and U4874 (N_4874,N_4707,N_4513);
and U4875 (N_4875,N_4659,N_4623);
or U4876 (N_4876,N_4493,N_4439);
xor U4877 (N_4877,N_4782,N_4797);
and U4878 (N_4878,N_4738,N_4688);
and U4879 (N_4879,N_4475,N_4586);
nand U4880 (N_4880,N_4610,N_4619);
nand U4881 (N_4881,N_4766,N_4625);
nor U4882 (N_4882,N_4758,N_4503);
nor U4883 (N_4883,N_4694,N_4723);
and U4884 (N_4884,N_4779,N_4418);
nor U4885 (N_4885,N_4787,N_4477);
or U4886 (N_4886,N_4498,N_4778);
or U4887 (N_4887,N_4502,N_4741);
xor U4888 (N_4888,N_4596,N_4454);
xnor U4889 (N_4889,N_4422,N_4448);
nor U4890 (N_4890,N_4479,N_4712);
nor U4891 (N_4891,N_4425,N_4670);
nand U4892 (N_4892,N_4543,N_4444);
xnor U4893 (N_4893,N_4523,N_4462);
nor U4894 (N_4894,N_4595,N_4791);
nor U4895 (N_4895,N_4473,N_4463);
and U4896 (N_4896,N_4767,N_4522);
nor U4897 (N_4897,N_4583,N_4538);
and U4898 (N_4898,N_4574,N_4552);
nand U4899 (N_4899,N_4592,N_4622);
and U4900 (N_4900,N_4533,N_4762);
nand U4901 (N_4901,N_4572,N_4729);
nor U4902 (N_4902,N_4768,N_4613);
and U4903 (N_4903,N_4437,N_4746);
nor U4904 (N_4904,N_4751,N_4776);
and U4905 (N_4905,N_4494,N_4654);
nand U4906 (N_4906,N_4608,N_4484);
xnor U4907 (N_4907,N_4764,N_4795);
and U4908 (N_4908,N_4721,N_4752);
nor U4909 (N_4909,N_4433,N_4747);
xnor U4910 (N_4910,N_4482,N_4451);
nand U4911 (N_4911,N_4404,N_4748);
nand U4912 (N_4912,N_4727,N_4516);
xnor U4913 (N_4913,N_4671,N_4792);
nor U4914 (N_4914,N_4602,N_4750);
or U4915 (N_4915,N_4628,N_4605);
or U4916 (N_4916,N_4504,N_4664);
and U4917 (N_4917,N_4563,N_4794);
xnor U4918 (N_4918,N_4680,N_4627);
xor U4919 (N_4919,N_4582,N_4447);
and U4920 (N_4920,N_4656,N_4491);
nor U4921 (N_4921,N_4611,N_4455);
nand U4922 (N_4922,N_4459,N_4591);
nor U4923 (N_4923,N_4467,N_4637);
nand U4924 (N_4924,N_4665,N_4500);
xor U4925 (N_4925,N_4460,N_4629);
or U4926 (N_4926,N_4436,N_4534);
and U4927 (N_4927,N_4784,N_4441);
xor U4928 (N_4928,N_4550,N_4509);
or U4929 (N_4929,N_4695,N_4511);
nand U4930 (N_4930,N_4600,N_4633);
nand U4931 (N_4931,N_4772,N_4755);
nor U4932 (N_4932,N_4703,N_4488);
and U4933 (N_4933,N_4715,N_4465);
nand U4934 (N_4934,N_4558,N_4744);
nor U4935 (N_4935,N_4506,N_4497);
xor U4936 (N_4936,N_4781,N_4754);
nor U4937 (N_4937,N_4643,N_4412);
and U4938 (N_4938,N_4681,N_4701);
and U4939 (N_4939,N_4646,N_4731);
and U4940 (N_4940,N_4535,N_4520);
and U4941 (N_4941,N_4512,N_4636);
xnor U4942 (N_4942,N_4737,N_4674);
and U4943 (N_4943,N_4706,N_4756);
nor U4944 (N_4944,N_4626,N_4486);
or U4945 (N_4945,N_4556,N_4528);
nor U4946 (N_4946,N_4403,N_4527);
nor U4947 (N_4947,N_4692,N_4432);
nand U4948 (N_4948,N_4658,N_4597);
and U4949 (N_4949,N_4489,N_4685);
and U4950 (N_4950,N_4569,N_4426);
and U4951 (N_4951,N_4732,N_4492);
nand U4952 (N_4952,N_4632,N_4471);
nor U4953 (N_4953,N_4419,N_4410);
nand U4954 (N_4954,N_4529,N_4584);
xnor U4955 (N_4955,N_4736,N_4442);
xnor U4956 (N_4956,N_4423,N_4693);
xor U4957 (N_4957,N_4469,N_4638);
xor U4958 (N_4958,N_4553,N_4678);
nand U4959 (N_4959,N_4698,N_4641);
xnor U4960 (N_4960,N_4726,N_4537);
and U4961 (N_4961,N_4416,N_4624);
and U4962 (N_4962,N_4603,N_4401);
nor U4963 (N_4963,N_4508,N_4519);
or U4964 (N_4964,N_4464,N_4530);
and U4965 (N_4965,N_4483,N_4697);
or U4966 (N_4966,N_4515,N_4739);
nor U4967 (N_4967,N_4734,N_4434);
nand U4968 (N_4968,N_4719,N_4774);
nor U4969 (N_4969,N_4525,N_4740);
nand U4970 (N_4970,N_4536,N_4435);
xor U4971 (N_4971,N_4400,N_4705);
or U4972 (N_4972,N_4661,N_4789);
nand U4973 (N_4973,N_4510,N_4621);
and U4974 (N_4974,N_4672,N_4785);
nand U4975 (N_4975,N_4414,N_4749);
or U4976 (N_4976,N_4702,N_4524);
and U4977 (N_4977,N_4742,N_4507);
or U4978 (N_4978,N_4691,N_4606);
or U4979 (N_4979,N_4424,N_4647);
xnor U4980 (N_4980,N_4716,N_4450);
nand U4981 (N_4981,N_4561,N_4790);
nand U4982 (N_4982,N_4655,N_4560);
or U4983 (N_4983,N_4771,N_4689);
nor U4984 (N_4984,N_4545,N_4593);
xor U4985 (N_4985,N_4532,N_4457);
nand U4986 (N_4986,N_4594,N_4761);
and U4987 (N_4987,N_4666,N_4710);
nand U4988 (N_4988,N_4541,N_4684);
nand U4989 (N_4989,N_4780,N_4555);
or U4990 (N_4990,N_4446,N_4657);
and U4991 (N_4991,N_4578,N_4798);
xnor U4992 (N_4992,N_4683,N_4588);
nor U4993 (N_4993,N_4676,N_4579);
or U4994 (N_4994,N_4687,N_4445);
xnor U4995 (N_4995,N_4428,N_4679);
xnor U4996 (N_4996,N_4580,N_4635);
and U4997 (N_4997,N_4609,N_4708);
and U4998 (N_4998,N_4480,N_4487);
xor U4999 (N_4999,N_4599,N_4745);
or U5000 (N_5000,N_4532,N_4769);
and U5001 (N_5001,N_4615,N_4501);
nand U5002 (N_5002,N_4455,N_4594);
or U5003 (N_5003,N_4728,N_4632);
or U5004 (N_5004,N_4714,N_4751);
nor U5005 (N_5005,N_4738,N_4724);
or U5006 (N_5006,N_4498,N_4631);
nand U5007 (N_5007,N_4433,N_4628);
or U5008 (N_5008,N_4479,N_4547);
and U5009 (N_5009,N_4660,N_4476);
xnor U5010 (N_5010,N_4698,N_4474);
nor U5011 (N_5011,N_4647,N_4611);
and U5012 (N_5012,N_4556,N_4629);
nand U5013 (N_5013,N_4777,N_4507);
xnor U5014 (N_5014,N_4716,N_4708);
xnor U5015 (N_5015,N_4562,N_4581);
and U5016 (N_5016,N_4402,N_4647);
and U5017 (N_5017,N_4465,N_4696);
xnor U5018 (N_5018,N_4562,N_4647);
xor U5019 (N_5019,N_4675,N_4731);
xnor U5020 (N_5020,N_4428,N_4469);
nand U5021 (N_5021,N_4506,N_4609);
or U5022 (N_5022,N_4425,N_4603);
nand U5023 (N_5023,N_4720,N_4513);
xnor U5024 (N_5024,N_4565,N_4449);
or U5025 (N_5025,N_4484,N_4697);
or U5026 (N_5026,N_4714,N_4616);
nand U5027 (N_5027,N_4701,N_4724);
and U5028 (N_5028,N_4438,N_4602);
nor U5029 (N_5029,N_4438,N_4745);
xor U5030 (N_5030,N_4625,N_4640);
xnor U5031 (N_5031,N_4715,N_4793);
and U5032 (N_5032,N_4733,N_4403);
and U5033 (N_5033,N_4497,N_4712);
or U5034 (N_5034,N_4592,N_4562);
nand U5035 (N_5035,N_4792,N_4765);
nand U5036 (N_5036,N_4580,N_4601);
xor U5037 (N_5037,N_4416,N_4761);
and U5038 (N_5038,N_4583,N_4520);
nor U5039 (N_5039,N_4451,N_4484);
xnor U5040 (N_5040,N_4753,N_4579);
and U5041 (N_5041,N_4559,N_4663);
and U5042 (N_5042,N_4610,N_4670);
or U5043 (N_5043,N_4736,N_4417);
or U5044 (N_5044,N_4525,N_4483);
or U5045 (N_5045,N_4745,N_4521);
nor U5046 (N_5046,N_4630,N_4615);
nand U5047 (N_5047,N_4569,N_4797);
and U5048 (N_5048,N_4585,N_4468);
or U5049 (N_5049,N_4513,N_4538);
nand U5050 (N_5050,N_4517,N_4792);
nand U5051 (N_5051,N_4701,N_4752);
nor U5052 (N_5052,N_4577,N_4489);
and U5053 (N_5053,N_4551,N_4752);
or U5054 (N_5054,N_4518,N_4730);
xnor U5055 (N_5055,N_4497,N_4722);
xor U5056 (N_5056,N_4557,N_4721);
nand U5057 (N_5057,N_4429,N_4704);
nor U5058 (N_5058,N_4680,N_4704);
nor U5059 (N_5059,N_4626,N_4439);
xor U5060 (N_5060,N_4695,N_4537);
nand U5061 (N_5061,N_4628,N_4536);
and U5062 (N_5062,N_4658,N_4604);
and U5063 (N_5063,N_4459,N_4683);
nor U5064 (N_5064,N_4556,N_4787);
nor U5065 (N_5065,N_4762,N_4680);
and U5066 (N_5066,N_4508,N_4664);
or U5067 (N_5067,N_4542,N_4431);
or U5068 (N_5068,N_4694,N_4576);
nor U5069 (N_5069,N_4686,N_4570);
or U5070 (N_5070,N_4541,N_4525);
nor U5071 (N_5071,N_4412,N_4764);
or U5072 (N_5072,N_4760,N_4443);
nand U5073 (N_5073,N_4668,N_4525);
xor U5074 (N_5074,N_4576,N_4417);
xor U5075 (N_5075,N_4560,N_4525);
xnor U5076 (N_5076,N_4653,N_4770);
or U5077 (N_5077,N_4662,N_4469);
nor U5078 (N_5078,N_4547,N_4591);
nand U5079 (N_5079,N_4531,N_4488);
nor U5080 (N_5080,N_4652,N_4649);
xnor U5081 (N_5081,N_4503,N_4588);
or U5082 (N_5082,N_4561,N_4746);
nor U5083 (N_5083,N_4696,N_4478);
nor U5084 (N_5084,N_4415,N_4764);
xnor U5085 (N_5085,N_4686,N_4766);
nor U5086 (N_5086,N_4472,N_4727);
nand U5087 (N_5087,N_4624,N_4631);
or U5088 (N_5088,N_4551,N_4521);
xnor U5089 (N_5089,N_4682,N_4734);
xnor U5090 (N_5090,N_4400,N_4579);
and U5091 (N_5091,N_4778,N_4708);
nor U5092 (N_5092,N_4594,N_4792);
nor U5093 (N_5093,N_4760,N_4406);
nor U5094 (N_5094,N_4659,N_4601);
xnor U5095 (N_5095,N_4778,N_4697);
or U5096 (N_5096,N_4692,N_4700);
nor U5097 (N_5097,N_4468,N_4553);
xnor U5098 (N_5098,N_4471,N_4432);
xor U5099 (N_5099,N_4619,N_4468);
nand U5100 (N_5100,N_4741,N_4600);
or U5101 (N_5101,N_4617,N_4506);
nor U5102 (N_5102,N_4795,N_4563);
nor U5103 (N_5103,N_4650,N_4414);
xor U5104 (N_5104,N_4445,N_4764);
and U5105 (N_5105,N_4737,N_4643);
nand U5106 (N_5106,N_4633,N_4622);
or U5107 (N_5107,N_4673,N_4716);
nor U5108 (N_5108,N_4539,N_4577);
nand U5109 (N_5109,N_4406,N_4435);
nor U5110 (N_5110,N_4412,N_4709);
xor U5111 (N_5111,N_4650,N_4457);
and U5112 (N_5112,N_4683,N_4714);
or U5113 (N_5113,N_4442,N_4682);
xor U5114 (N_5114,N_4705,N_4789);
and U5115 (N_5115,N_4641,N_4697);
nor U5116 (N_5116,N_4626,N_4631);
nor U5117 (N_5117,N_4482,N_4470);
xor U5118 (N_5118,N_4488,N_4715);
xor U5119 (N_5119,N_4673,N_4455);
and U5120 (N_5120,N_4562,N_4693);
nand U5121 (N_5121,N_4774,N_4680);
xor U5122 (N_5122,N_4511,N_4561);
nor U5123 (N_5123,N_4730,N_4457);
nand U5124 (N_5124,N_4508,N_4513);
nand U5125 (N_5125,N_4675,N_4615);
nor U5126 (N_5126,N_4689,N_4650);
nor U5127 (N_5127,N_4712,N_4487);
nand U5128 (N_5128,N_4585,N_4694);
and U5129 (N_5129,N_4607,N_4569);
nand U5130 (N_5130,N_4525,N_4447);
and U5131 (N_5131,N_4747,N_4531);
and U5132 (N_5132,N_4481,N_4650);
nor U5133 (N_5133,N_4739,N_4429);
and U5134 (N_5134,N_4652,N_4534);
and U5135 (N_5135,N_4457,N_4624);
xor U5136 (N_5136,N_4533,N_4449);
or U5137 (N_5137,N_4611,N_4475);
and U5138 (N_5138,N_4553,N_4410);
and U5139 (N_5139,N_4432,N_4704);
nor U5140 (N_5140,N_4410,N_4566);
xor U5141 (N_5141,N_4533,N_4461);
or U5142 (N_5142,N_4467,N_4542);
nand U5143 (N_5143,N_4631,N_4620);
or U5144 (N_5144,N_4721,N_4765);
nor U5145 (N_5145,N_4539,N_4740);
xnor U5146 (N_5146,N_4685,N_4730);
and U5147 (N_5147,N_4678,N_4732);
xnor U5148 (N_5148,N_4588,N_4666);
nor U5149 (N_5149,N_4400,N_4772);
xor U5150 (N_5150,N_4529,N_4707);
nor U5151 (N_5151,N_4635,N_4741);
nor U5152 (N_5152,N_4566,N_4546);
nand U5153 (N_5153,N_4578,N_4505);
xor U5154 (N_5154,N_4603,N_4667);
or U5155 (N_5155,N_4712,N_4757);
or U5156 (N_5156,N_4748,N_4602);
and U5157 (N_5157,N_4439,N_4798);
nand U5158 (N_5158,N_4794,N_4437);
and U5159 (N_5159,N_4797,N_4507);
nor U5160 (N_5160,N_4773,N_4546);
nand U5161 (N_5161,N_4729,N_4496);
and U5162 (N_5162,N_4682,N_4681);
nand U5163 (N_5163,N_4746,N_4425);
nor U5164 (N_5164,N_4746,N_4552);
or U5165 (N_5165,N_4575,N_4517);
xnor U5166 (N_5166,N_4681,N_4707);
and U5167 (N_5167,N_4481,N_4729);
nand U5168 (N_5168,N_4662,N_4650);
nand U5169 (N_5169,N_4700,N_4704);
and U5170 (N_5170,N_4460,N_4718);
or U5171 (N_5171,N_4520,N_4444);
nor U5172 (N_5172,N_4621,N_4444);
or U5173 (N_5173,N_4753,N_4477);
and U5174 (N_5174,N_4639,N_4738);
or U5175 (N_5175,N_4417,N_4543);
nor U5176 (N_5176,N_4787,N_4602);
nor U5177 (N_5177,N_4594,N_4437);
xor U5178 (N_5178,N_4585,N_4500);
or U5179 (N_5179,N_4533,N_4736);
nand U5180 (N_5180,N_4448,N_4634);
nor U5181 (N_5181,N_4608,N_4589);
xor U5182 (N_5182,N_4611,N_4593);
or U5183 (N_5183,N_4733,N_4762);
nand U5184 (N_5184,N_4428,N_4500);
or U5185 (N_5185,N_4613,N_4401);
xor U5186 (N_5186,N_4401,N_4441);
xor U5187 (N_5187,N_4532,N_4449);
nor U5188 (N_5188,N_4726,N_4626);
nor U5189 (N_5189,N_4602,N_4416);
nor U5190 (N_5190,N_4632,N_4578);
nand U5191 (N_5191,N_4716,N_4594);
or U5192 (N_5192,N_4772,N_4520);
nor U5193 (N_5193,N_4684,N_4581);
nand U5194 (N_5194,N_4635,N_4481);
xnor U5195 (N_5195,N_4699,N_4426);
xor U5196 (N_5196,N_4639,N_4506);
nor U5197 (N_5197,N_4661,N_4584);
nand U5198 (N_5198,N_4482,N_4429);
xnor U5199 (N_5199,N_4657,N_4459);
and U5200 (N_5200,N_4940,N_4980);
and U5201 (N_5201,N_4813,N_4983);
nor U5202 (N_5202,N_5037,N_4965);
or U5203 (N_5203,N_5132,N_4915);
or U5204 (N_5204,N_4853,N_4852);
and U5205 (N_5205,N_4814,N_4962);
and U5206 (N_5206,N_4874,N_4892);
nand U5207 (N_5207,N_4829,N_4803);
xor U5208 (N_5208,N_4947,N_4968);
xnor U5209 (N_5209,N_4828,N_4825);
xnor U5210 (N_5210,N_5087,N_4954);
nor U5211 (N_5211,N_4952,N_4903);
nor U5212 (N_5212,N_4864,N_5008);
and U5213 (N_5213,N_5133,N_4811);
xnor U5214 (N_5214,N_5131,N_4946);
nor U5215 (N_5215,N_4970,N_4887);
nor U5216 (N_5216,N_4847,N_5102);
xor U5217 (N_5217,N_4821,N_4950);
nor U5218 (N_5218,N_5091,N_4808);
nand U5219 (N_5219,N_5177,N_5136);
nand U5220 (N_5220,N_5085,N_5140);
and U5221 (N_5221,N_4839,N_4804);
nor U5222 (N_5222,N_4832,N_4870);
and U5223 (N_5223,N_4920,N_4926);
or U5224 (N_5224,N_4949,N_4942);
xnor U5225 (N_5225,N_5105,N_4869);
nand U5226 (N_5226,N_5005,N_4816);
nor U5227 (N_5227,N_5064,N_4830);
and U5228 (N_5228,N_4921,N_4898);
xnor U5229 (N_5229,N_5072,N_5106);
xnor U5230 (N_5230,N_5029,N_4939);
nor U5231 (N_5231,N_5184,N_4857);
nand U5232 (N_5232,N_4871,N_4851);
and U5233 (N_5233,N_4937,N_4990);
xnor U5234 (N_5234,N_5180,N_5117);
and U5235 (N_5235,N_5161,N_4979);
nand U5236 (N_5236,N_4998,N_5048);
nor U5237 (N_5237,N_4985,N_5081);
or U5238 (N_5238,N_4890,N_5188);
nand U5239 (N_5239,N_5014,N_4823);
nand U5240 (N_5240,N_4882,N_4809);
nand U5241 (N_5241,N_4900,N_5063);
nand U5242 (N_5242,N_4880,N_4984);
or U5243 (N_5243,N_4810,N_4910);
nand U5244 (N_5244,N_4817,N_5069);
or U5245 (N_5245,N_4815,N_4833);
nor U5246 (N_5246,N_4895,N_5032);
nand U5247 (N_5247,N_5114,N_5143);
nand U5248 (N_5248,N_4917,N_4801);
and U5249 (N_5249,N_5027,N_4888);
nor U5250 (N_5250,N_5192,N_5185);
or U5251 (N_5251,N_4836,N_5183);
nand U5252 (N_5252,N_5111,N_4842);
or U5253 (N_5253,N_4835,N_5138);
nor U5254 (N_5254,N_5078,N_5066);
nor U5255 (N_5255,N_4807,N_5084);
nor U5256 (N_5256,N_5057,N_4924);
or U5257 (N_5257,N_4894,N_4974);
nand U5258 (N_5258,N_5196,N_5083);
nand U5259 (N_5259,N_5122,N_4916);
xor U5260 (N_5260,N_4805,N_4971);
or U5261 (N_5261,N_5082,N_5047);
nand U5262 (N_5262,N_5011,N_4841);
and U5263 (N_5263,N_5017,N_4854);
xor U5264 (N_5264,N_5164,N_5067);
nor U5265 (N_5265,N_4929,N_4928);
nand U5266 (N_5266,N_4893,N_5059);
xnor U5267 (N_5267,N_5071,N_5109);
or U5268 (N_5268,N_5086,N_4992);
nor U5269 (N_5269,N_5018,N_5137);
and U5270 (N_5270,N_4879,N_4850);
or U5271 (N_5271,N_5034,N_4849);
or U5272 (N_5272,N_4914,N_5156);
xor U5273 (N_5273,N_5020,N_4820);
nand U5274 (N_5274,N_5186,N_4867);
and U5275 (N_5275,N_5075,N_5160);
or U5276 (N_5276,N_5182,N_5135);
and U5277 (N_5277,N_5147,N_5033);
xnor U5278 (N_5278,N_5049,N_4886);
nor U5279 (N_5279,N_5019,N_5159);
xnor U5280 (N_5280,N_5103,N_4905);
and U5281 (N_5281,N_4997,N_4812);
and U5282 (N_5282,N_4961,N_4945);
nand U5283 (N_5283,N_5062,N_4936);
xor U5284 (N_5284,N_4846,N_4856);
xnor U5285 (N_5285,N_5098,N_5054);
or U5286 (N_5286,N_5190,N_5024);
and U5287 (N_5287,N_4902,N_4875);
and U5288 (N_5288,N_5055,N_4931);
nand U5289 (N_5289,N_4911,N_5139);
nor U5290 (N_5290,N_5058,N_4987);
and U5291 (N_5291,N_4938,N_5129);
and U5292 (N_5292,N_4935,N_4858);
and U5293 (N_5293,N_5036,N_4933);
xor U5294 (N_5294,N_5007,N_4883);
nand U5295 (N_5295,N_5187,N_4824);
nand U5296 (N_5296,N_4923,N_5130);
xor U5297 (N_5297,N_4963,N_5015);
and U5298 (N_5298,N_5070,N_4843);
or U5299 (N_5299,N_4845,N_5004);
nand U5300 (N_5300,N_5068,N_5176);
nor U5301 (N_5301,N_4904,N_4969);
or U5302 (N_5302,N_4927,N_4891);
and U5303 (N_5303,N_5197,N_5128);
or U5304 (N_5304,N_5031,N_5028);
or U5305 (N_5305,N_5169,N_4860);
or U5306 (N_5306,N_4982,N_5120);
or U5307 (N_5307,N_5096,N_5170);
nor U5308 (N_5308,N_5149,N_5000);
nor U5309 (N_5309,N_5021,N_5056);
nor U5310 (N_5310,N_5151,N_4944);
or U5311 (N_5311,N_5181,N_5023);
nand U5312 (N_5312,N_4848,N_5089);
nand U5313 (N_5313,N_5010,N_5094);
or U5314 (N_5314,N_4958,N_5107);
and U5315 (N_5315,N_4876,N_4953);
xnor U5316 (N_5316,N_5154,N_4827);
nand U5317 (N_5317,N_4932,N_4906);
or U5318 (N_5318,N_5061,N_5092);
xor U5319 (N_5319,N_4918,N_5053);
nor U5320 (N_5320,N_4806,N_5003);
and U5321 (N_5321,N_5100,N_4988);
xnor U5322 (N_5322,N_4896,N_5039);
or U5323 (N_5323,N_5041,N_4959);
nand U5324 (N_5324,N_4951,N_4802);
nand U5325 (N_5325,N_5127,N_5150);
nand U5326 (N_5326,N_5171,N_5108);
xor U5327 (N_5327,N_5157,N_5097);
nor U5328 (N_5328,N_4855,N_4826);
xnor U5329 (N_5329,N_4975,N_5162);
nand U5330 (N_5330,N_5142,N_5088);
and U5331 (N_5331,N_5166,N_4819);
xnor U5332 (N_5332,N_5141,N_5099);
and U5333 (N_5333,N_5040,N_4863);
and U5334 (N_5334,N_5101,N_4955);
nand U5335 (N_5335,N_5153,N_5022);
xor U5336 (N_5336,N_5026,N_5126);
xor U5337 (N_5337,N_4877,N_5052);
and U5338 (N_5338,N_4925,N_5110);
and U5339 (N_5339,N_5165,N_5112);
nand U5340 (N_5340,N_5191,N_4866);
nor U5341 (N_5341,N_5194,N_5045);
and U5342 (N_5342,N_5178,N_4919);
xor U5343 (N_5343,N_4859,N_5198);
or U5344 (N_5344,N_5044,N_4834);
or U5345 (N_5345,N_4930,N_4999);
nand U5346 (N_5346,N_4948,N_5043);
nor U5347 (N_5347,N_4899,N_4818);
and U5348 (N_5348,N_4861,N_4994);
or U5349 (N_5349,N_4986,N_4981);
xor U5350 (N_5350,N_5042,N_5175);
and U5351 (N_5351,N_4862,N_5155);
or U5352 (N_5352,N_4956,N_4881);
xnor U5353 (N_5353,N_5076,N_5013);
nand U5354 (N_5354,N_5104,N_4996);
or U5355 (N_5355,N_5125,N_5124);
or U5356 (N_5356,N_4964,N_5060);
xor U5357 (N_5357,N_5118,N_4977);
nand U5358 (N_5358,N_5025,N_5030);
xor U5359 (N_5359,N_5195,N_4943);
or U5360 (N_5360,N_5035,N_5199);
xor U5361 (N_5361,N_4907,N_4976);
and U5362 (N_5362,N_4884,N_4957);
or U5363 (N_5363,N_4865,N_5115);
xnor U5364 (N_5364,N_5189,N_4901);
or U5365 (N_5365,N_4934,N_5095);
nor U5366 (N_5366,N_4973,N_5038);
and U5367 (N_5367,N_5134,N_4837);
xnor U5368 (N_5368,N_5051,N_4831);
and U5369 (N_5369,N_5174,N_4912);
xor U5370 (N_5370,N_5116,N_4967);
nand U5371 (N_5371,N_4897,N_5001);
and U5372 (N_5372,N_4993,N_4991);
and U5373 (N_5373,N_5090,N_5093);
or U5374 (N_5374,N_5119,N_5113);
nand U5375 (N_5375,N_4885,N_4989);
or U5376 (N_5376,N_5050,N_4941);
nand U5377 (N_5377,N_5179,N_5073);
or U5378 (N_5378,N_4873,N_4889);
and U5379 (N_5379,N_5163,N_5065);
and U5380 (N_5380,N_4978,N_4800);
or U5381 (N_5381,N_4844,N_5167);
and U5382 (N_5382,N_5148,N_5009);
and U5383 (N_5383,N_4909,N_5121);
xor U5384 (N_5384,N_4972,N_4838);
or U5385 (N_5385,N_5012,N_4922);
and U5386 (N_5386,N_5006,N_5077);
nand U5387 (N_5387,N_4908,N_5173);
nand U5388 (N_5388,N_4878,N_5172);
nand U5389 (N_5389,N_5080,N_5079);
or U5390 (N_5390,N_5002,N_5145);
xor U5391 (N_5391,N_4913,N_5123);
nand U5392 (N_5392,N_5146,N_5046);
xnor U5393 (N_5393,N_4872,N_5152);
xor U5394 (N_5394,N_5074,N_4868);
and U5395 (N_5395,N_4840,N_4822);
or U5396 (N_5396,N_4995,N_5168);
and U5397 (N_5397,N_5193,N_4960);
nor U5398 (N_5398,N_5158,N_5016);
nand U5399 (N_5399,N_4966,N_5144);
nand U5400 (N_5400,N_4967,N_4998);
or U5401 (N_5401,N_4855,N_5187);
nor U5402 (N_5402,N_5008,N_4826);
and U5403 (N_5403,N_5026,N_4816);
nor U5404 (N_5404,N_4912,N_5168);
nand U5405 (N_5405,N_4846,N_4957);
nand U5406 (N_5406,N_5120,N_5143);
xnor U5407 (N_5407,N_5146,N_4992);
or U5408 (N_5408,N_4965,N_5168);
and U5409 (N_5409,N_4801,N_5162);
nand U5410 (N_5410,N_4846,N_4928);
nand U5411 (N_5411,N_5183,N_4870);
xor U5412 (N_5412,N_5036,N_5095);
nand U5413 (N_5413,N_4991,N_4941);
or U5414 (N_5414,N_4886,N_4941);
and U5415 (N_5415,N_5126,N_5146);
nand U5416 (N_5416,N_4858,N_4827);
or U5417 (N_5417,N_5184,N_4914);
and U5418 (N_5418,N_4856,N_5091);
xor U5419 (N_5419,N_5128,N_4872);
nor U5420 (N_5420,N_5030,N_5105);
xnor U5421 (N_5421,N_5063,N_4958);
and U5422 (N_5422,N_5013,N_5051);
or U5423 (N_5423,N_4946,N_5065);
nand U5424 (N_5424,N_4802,N_4910);
nand U5425 (N_5425,N_5114,N_5052);
nand U5426 (N_5426,N_4970,N_4842);
xor U5427 (N_5427,N_4892,N_5117);
or U5428 (N_5428,N_5145,N_5067);
nand U5429 (N_5429,N_5142,N_4999);
or U5430 (N_5430,N_5124,N_5192);
xnor U5431 (N_5431,N_4956,N_5097);
nand U5432 (N_5432,N_4925,N_5112);
xor U5433 (N_5433,N_4828,N_4802);
and U5434 (N_5434,N_4990,N_4870);
or U5435 (N_5435,N_5073,N_4907);
nor U5436 (N_5436,N_5051,N_5042);
nand U5437 (N_5437,N_5031,N_4816);
or U5438 (N_5438,N_5022,N_5122);
nor U5439 (N_5439,N_5039,N_4910);
nor U5440 (N_5440,N_5102,N_4823);
nor U5441 (N_5441,N_5150,N_5194);
nor U5442 (N_5442,N_5103,N_5141);
nor U5443 (N_5443,N_5066,N_4877);
or U5444 (N_5444,N_5139,N_4842);
or U5445 (N_5445,N_5134,N_5031);
xor U5446 (N_5446,N_5148,N_5045);
nand U5447 (N_5447,N_5172,N_5187);
or U5448 (N_5448,N_4843,N_4831);
or U5449 (N_5449,N_4970,N_5091);
or U5450 (N_5450,N_5004,N_4885);
nor U5451 (N_5451,N_5142,N_5166);
or U5452 (N_5452,N_4957,N_5108);
nand U5453 (N_5453,N_5175,N_5154);
nand U5454 (N_5454,N_5115,N_5019);
xnor U5455 (N_5455,N_4883,N_5131);
or U5456 (N_5456,N_5169,N_4822);
xor U5457 (N_5457,N_5099,N_4839);
and U5458 (N_5458,N_5000,N_4977);
xnor U5459 (N_5459,N_4870,N_4962);
or U5460 (N_5460,N_5176,N_4963);
nor U5461 (N_5461,N_5059,N_5176);
or U5462 (N_5462,N_4900,N_4811);
nand U5463 (N_5463,N_5166,N_4833);
or U5464 (N_5464,N_4936,N_5165);
or U5465 (N_5465,N_4890,N_5057);
or U5466 (N_5466,N_5005,N_4974);
or U5467 (N_5467,N_5065,N_5023);
nand U5468 (N_5468,N_5087,N_4950);
nand U5469 (N_5469,N_4831,N_5081);
nand U5470 (N_5470,N_4902,N_5074);
or U5471 (N_5471,N_5070,N_5120);
nor U5472 (N_5472,N_4925,N_4954);
nand U5473 (N_5473,N_5116,N_5003);
nand U5474 (N_5474,N_4935,N_5199);
xnor U5475 (N_5475,N_5042,N_4849);
nand U5476 (N_5476,N_4981,N_4966);
nor U5477 (N_5477,N_5091,N_4836);
or U5478 (N_5478,N_4873,N_5108);
and U5479 (N_5479,N_5093,N_4838);
and U5480 (N_5480,N_5035,N_5107);
or U5481 (N_5481,N_5029,N_5031);
nand U5482 (N_5482,N_5106,N_5007);
nand U5483 (N_5483,N_5070,N_5011);
xnor U5484 (N_5484,N_5126,N_5164);
nand U5485 (N_5485,N_5101,N_4817);
nand U5486 (N_5486,N_5020,N_5035);
nor U5487 (N_5487,N_4829,N_5076);
nand U5488 (N_5488,N_4906,N_5006);
nor U5489 (N_5489,N_4836,N_5003);
nand U5490 (N_5490,N_4902,N_4949);
and U5491 (N_5491,N_5139,N_5022);
and U5492 (N_5492,N_5120,N_4867);
or U5493 (N_5493,N_5175,N_4898);
xor U5494 (N_5494,N_5138,N_5148);
and U5495 (N_5495,N_5176,N_5131);
nor U5496 (N_5496,N_4985,N_4939);
xor U5497 (N_5497,N_5121,N_5020);
nand U5498 (N_5498,N_5133,N_4908);
or U5499 (N_5499,N_5193,N_4842);
nor U5500 (N_5500,N_4926,N_5005);
or U5501 (N_5501,N_5045,N_5159);
xor U5502 (N_5502,N_4969,N_4823);
nor U5503 (N_5503,N_5122,N_4947);
nand U5504 (N_5504,N_5018,N_4937);
xor U5505 (N_5505,N_4858,N_4855);
nor U5506 (N_5506,N_4944,N_5077);
xor U5507 (N_5507,N_4829,N_5196);
nor U5508 (N_5508,N_4897,N_5069);
or U5509 (N_5509,N_4967,N_5073);
and U5510 (N_5510,N_4863,N_5193);
or U5511 (N_5511,N_4928,N_4847);
nor U5512 (N_5512,N_5090,N_4884);
and U5513 (N_5513,N_4930,N_5168);
and U5514 (N_5514,N_5013,N_5193);
xor U5515 (N_5515,N_4864,N_4987);
nand U5516 (N_5516,N_4960,N_5078);
and U5517 (N_5517,N_4824,N_4920);
and U5518 (N_5518,N_4967,N_4993);
nand U5519 (N_5519,N_5027,N_4818);
and U5520 (N_5520,N_5036,N_4917);
nor U5521 (N_5521,N_4870,N_4918);
xnor U5522 (N_5522,N_4816,N_4997);
xor U5523 (N_5523,N_4907,N_5055);
nand U5524 (N_5524,N_5191,N_4961);
nand U5525 (N_5525,N_4952,N_5079);
nor U5526 (N_5526,N_5087,N_4963);
xor U5527 (N_5527,N_5169,N_5041);
nand U5528 (N_5528,N_5044,N_4921);
and U5529 (N_5529,N_4955,N_5009);
and U5530 (N_5530,N_5095,N_5062);
nor U5531 (N_5531,N_4941,N_4994);
or U5532 (N_5532,N_4949,N_5031);
or U5533 (N_5533,N_5106,N_4912);
nand U5534 (N_5534,N_4852,N_5019);
nand U5535 (N_5535,N_4882,N_4914);
and U5536 (N_5536,N_5008,N_4828);
nand U5537 (N_5537,N_5179,N_5072);
nor U5538 (N_5538,N_5168,N_5059);
nor U5539 (N_5539,N_4920,N_4892);
and U5540 (N_5540,N_4878,N_5020);
xnor U5541 (N_5541,N_4853,N_5162);
xnor U5542 (N_5542,N_4891,N_5117);
xnor U5543 (N_5543,N_5182,N_4924);
or U5544 (N_5544,N_5085,N_5078);
xor U5545 (N_5545,N_5016,N_5021);
nor U5546 (N_5546,N_5090,N_5179);
or U5547 (N_5547,N_5055,N_4875);
nand U5548 (N_5548,N_5162,N_5001);
and U5549 (N_5549,N_5092,N_5151);
nand U5550 (N_5550,N_4807,N_4871);
nor U5551 (N_5551,N_5124,N_4891);
and U5552 (N_5552,N_5052,N_5097);
nor U5553 (N_5553,N_5110,N_4814);
or U5554 (N_5554,N_5039,N_5146);
and U5555 (N_5555,N_5175,N_4962);
nor U5556 (N_5556,N_5036,N_5114);
nor U5557 (N_5557,N_4804,N_4924);
nand U5558 (N_5558,N_4876,N_4881);
and U5559 (N_5559,N_4880,N_5119);
or U5560 (N_5560,N_4926,N_4800);
nor U5561 (N_5561,N_4966,N_4832);
xnor U5562 (N_5562,N_4847,N_5157);
xnor U5563 (N_5563,N_4976,N_4998);
or U5564 (N_5564,N_4939,N_5068);
nand U5565 (N_5565,N_4856,N_4853);
nor U5566 (N_5566,N_5056,N_5130);
or U5567 (N_5567,N_5113,N_4866);
xnor U5568 (N_5568,N_4890,N_4943);
xnor U5569 (N_5569,N_5056,N_4839);
nor U5570 (N_5570,N_4893,N_4896);
or U5571 (N_5571,N_5032,N_4985);
nand U5572 (N_5572,N_4831,N_4938);
xnor U5573 (N_5573,N_4890,N_5090);
and U5574 (N_5574,N_4876,N_5093);
or U5575 (N_5575,N_4815,N_4963);
xnor U5576 (N_5576,N_4895,N_5037);
or U5577 (N_5577,N_5182,N_4969);
nand U5578 (N_5578,N_4956,N_5086);
xnor U5579 (N_5579,N_5082,N_5127);
or U5580 (N_5580,N_5186,N_4869);
or U5581 (N_5581,N_4958,N_4957);
nand U5582 (N_5582,N_5075,N_4862);
nand U5583 (N_5583,N_4835,N_4804);
nand U5584 (N_5584,N_4810,N_4981);
nand U5585 (N_5585,N_5116,N_5026);
or U5586 (N_5586,N_5127,N_5010);
xor U5587 (N_5587,N_5134,N_5164);
and U5588 (N_5588,N_5011,N_4958);
nand U5589 (N_5589,N_4903,N_5140);
or U5590 (N_5590,N_4894,N_4982);
nor U5591 (N_5591,N_4941,N_4900);
xnor U5592 (N_5592,N_5193,N_4907);
nor U5593 (N_5593,N_4960,N_4802);
or U5594 (N_5594,N_5084,N_4939);
or U5595 (N_5595,N_4902,N_4939);
xnor U5596 (N_5596,N_4864,N_5139);
xor U5597 (N_5597,N_5072,N_5060);
and U5598 (N_5598,N_4911,N_5105);
or U5599 (N_5599,N_5029,N_5175);
and U5600 (N_5600,N_5367,N_5463);
or U5601 (N_5601,N_5396,N_5250);
and U5602 (N_5602,N_5405,N_5215);
and U5603 (N_5603,N_5425,N_5269);
nor U5604 (N_5604,N_5502,N_5442);
and U5605 (N_5605,N_5232,N_5468);
or U5606 (N_5606,N_5544,N_5496);
nor U5607 (N_5607,N_5323,N_5289);
nor U5608 (N_5608,N_5589,N_5572);
or U5609 (N_5609,N_5492,N_5374);
and U5610 (N_5610,N_5504,N_5590);
xor U5611 (N_5611,N_5552,N_5527);
and U5612 (N_5612,N_5252,N_5313);
nand U5613 (N_5613,N_5387,N_5267);
nor U5614 (N_5614,N_5228,N_5320);
or U5615 (N_5615,N_5414,N_5540);
nand U5616 (N_5616,N_5460,N_5231);
nand U5617 (N_5617,N_5211,N_5410);
xnor U5618 (N_5618,N_5408,N_5562);
nor U5619 (N_5619,N_5518,N_5418);
nand U5620 (N_5620,N_5413,N_5517);
and U5621 (N_5621,N_5435,N_5475);
nor U5622 (N_5622,N_5542,N_5292);
nand U5623 (N_5623,N_5419,N_5343);
nand U5624 (N_5624,N_5240,N_5402);
or U5625 (N_5625,N_5275,N_5516);
nor U5626 (N_5626,N_5422,N_5317);
xnor U5627 (N_5627,N_5281,N_5441);
xor U5628 (N_5628,N_5263,N_5308);
nand U5629 (N_5629,N_5225,N_5278);
nand U5630 (N_5630,N_5213,N_5244);
nor U5631 (N_5631,N_5327,N_5285);
and U5632 (N_5632,N_5365,N_5484);
xor U5633 (N_5633,N_5479,N_5537);
or U5634 (N_5634,N_5257,N_5530);
nor U5635 (N_5635,N_5322,N_5245);
nor U5636 (N_5636,N_5533,N_5432);
or U5637 (N_5637,N_5597,N_5534);
nor U5638 (N_5638,N_5394,N_5403);
nor U5639 (N_5639,N_5349,N_5337);
xor U5640 (N_5640,N_5456,N_5575);
or U5641 (N_5641,N_5401,N_5581);
and U5642 (N_5642,N_5279,N_5598);
and U5643 (N_5643,N_5525,N_5453);
nand U5644 (N_5644,N_5406,N_5353);
nor U5645 (N_5645,N_5212,N_5461);
xor U5646 (N_5646,N_5264,N_5217);
and U5647 (N_5647,N_5248,N_5481);
and U5648 (N_5648,N_5336,N_5272);
nand U5649 (N_5649,N_5535,N_5591);
xnor U5650 (N_5650,N_5407,N_5478);
nor U5651 (N_5651,N_5316,N_5383);
nor U5652 (N_5652,N_5446,N_5315);
nor U5653 (N_5653,N_5411,N_5564);
nor U5654 (N_5654,N_5362,N_5208);
nor U5655 (N_5655,N_5237,N_5295);
nor U5656 (N_5656,N_5233,N_5444);
nor U5657 (N_5657,N_5288,N_5437);
nand U5658 (N_5658,N_5369,N_5393);
or U5659 (N_5659,N_5286,N_5273);
xor U5660 (N_5660,N_5451,N_5270);
or U5661 (N_5661,N_5338,N_5253);
nor U5662 (N_5662,N_5366,N_5464);
nand U5663 (N_5663,N_5235,N_5522);
and U5664 (N_5664,N_5205,N_5566);
or U5665 (N_5665,N_5238,N_5578);
or U5666 (N_5666,N_5465,N_5459);
nor U5667 (N_5667,N_5571,N_5259);
or U5668 (N_5668,N_5584,N_5548);
and U5669 (N_5669,N_5471,N_5384);
xor U5670 (N_5670,N_5326,N_5551);
nor U5671 (N_5671,N_5271,N_5420);
nor U5672 (N_5672,N_5200,N_5489);
xor U5673 (N_5673,N_5351,N_5380);
and U5674 (N_5674,N_5251,N_5427);
nor U5675 (N_5675,N_5358,N_5550);
and U5676 (N_5676,N_5477,N_5574);
xor U5677 (N_5677,N_5226,N_5487);
and U5678 (N_5678,N_5538,N_5221);
nor U5679 (N_5679,N_5577,N_5543);
or U5680 (N_5680,N_5368,N_5529);
xnor U5681 (N_5681,N_5519,N_5301);
nand U5682 (N_5682,N_5229,N_5547);
nor U5683 (N_5683,N_5483,N_5379);
and U5684 (N_5684,N_5596,N_5284);
nand U5685 (N_5685,N_5207,N_5470);
nor U5686 (N_5686,N_5400,N_5583);
nand U5687 (N_5687,N_5390,N_5310);
nor U5688 (N_5688,N_5595,N_5412);
nor U5689 (N_5689,N_5234,N_5239);
and U5690 (N_5690,N_5485,N_5559);
and U5691 (N_5691,N_5436,N_5345);
nor U5692 (N_5692,N_5227,N_5206);
and U5693 (N_5693,N_5523,N_5386);
nor U5694 (N_5694,N_5311,N_5563);
or U5695 (N_5695,N_5218,N_5256);
xor U5696 (N_5696,N_5261,N_5415);
nor U5697 (N_5697,N_5399,N_5381);
and U5698 (N_5698,N_5296,N_5568);
and U5699 (N_5699,N_5291,N_5507);
and U5700 (N_5700,N_5495,N_5569);
and U5701 (N_5701,N_5486,N_5354);
or U5702 (N_5702,N_5204,N_5341);
or U5703 (N_5703,N_5222,N_5249);
and U5704 (N_5704,N_5472,N_5498);
nand U5705 (N_5705,N_5500,N_5283);
or U5706 (N_5706,N_5364,N_5579);
nor U5707 (N_5707,N_5265,N_5546);
or U5708 (N_5708,N_5592,N_5305);
nor U5709 (N_5709,N_5333,N_5255);
nor U5710 (N_5710,N_5560,N_5545);
and U5711 (N_5711,N_5203,N_5306);
and U5712 (N_5712,N_5541,N_5309);
or U5713 (N_5713,N_5321,N_5230);
and U5714 (N_5714,N_5329,N_5359);
nor U5715 (N_5715,N_5312,N_5440);
nand U5716 (N_5716,N_5377,N_5428);
xnor U5717 (N_5717,N_5580,N_5268);
or U5718 (N_5718,N_5335,N_5370);
and U5719 (N_5719,N_5332,N_5448);
xnor U5720 (N_5720,N_5392,N_5431);
and U5721 (N_5721,N_5356,N_5473);
or U5722 (N_5722,N_5357,N_5509);
or U5723 (N_5723,N_5299,N_5493);
nand U5724 (N_5724,N_5482,N_5450);
nand U5725 (N_5725,N_5494,N_5382);
or U5726 (N_5726,N_5378,N_5346);
or U5727 (N_5727,N_5219,N_5404);
nor U5728 (N_5728,N_5355,N_5416);
or U5729 (N_5729,N_5554,N_5524);
xor U5730 (N_5730,N_5304,N_5510);
and U5731 (N_5731,N_5526,N_5202);
nand U5732 (N_5732,N_5254,N_5302);
nand U5733 (N_5733,N_5576,N_5503);
nand U5734 (N_5734,N_5434,N_5521);
nor U5735 (N_5735,N_5558,N_5508);
and U5736 (N_5736,N_5247,N_5389);
or U5737 (N_5737,N_5277,N_5449);
or U5738 (N_5738,N_5445,N_5290);
nand U5739 (N_5739,N_5447,N_5314);
nor U5740 (N_5740,N_5586,N_5458);
xor U5741 (N_5741,N_5474,N_5201);
or U5742 (N_5742,N_5438,N_5488);
nand U5743 (N_5743,N_5512,N_5505);
xnor U5744 (N_5744,N_5328,N_5210);
xor U5745 (N_5745,N_5433,N_5531);
nand U5746 (N_5746,N_5209,N_5398);
and U5747 (N_5747,N_5424,N_5466);
nand U5748 (N_5748,N_5395,N_5397);
xor U5749 (N_5749,N_5452,N_5565);
and U5750 (N_5750,N_5480,N_5599);
xor U5751 (N_5751,N_5266,N_5243);
xnor U5752 (N_5752,N_5573,N_5375);
nand U5753 (N_5753,N_5372,N_5506);
and U5754 (N_5754,N_5443,N_5262);
nor U5755 (N_5755,N_5342,N_5439);
xnor U5756 (N_5756,N_5258,N_5348);
nor U5757 (N_5757,N_5499,N_5567);
nand U5758 (N_5758,N_5319,N_5347);
and U5759 (N_5759,N_5360,N_5553);
or U5760 (N_5760,N_5287,N_5469);
and U5761 (N_5761,N_5555,N_5462);
nor U5762 (N_5762,N_5339,N_5330);
and U5763 (N_5763,N_5260,N_5220);
xor U5764 (N_5764,N_5388,N_5371);
xnor U5765 (N_5765,N_5421,N_5497);
xor U5766 (N_5766,N_5280,N_5491);
xnor U5767 (N_5767,N_5556,N_5385);
xor U5768 (N_5768,N_5476,N_5361);
nor U5769 (N_5769,N_5511,N_5587);
and U5770 (N_5770,N_5223,N_5536);
and U5771 (N_5771,N_5561,N_5246);
nand U5772 (N_5772,N_5298,N_5303);
and U5773 (N_5773,N_5430,N_5455);
nor U5774 (N_5774,N_5318,N_5514);
nor U5775 (N_5775,N_5300,N_5373);
and U5776 (N_5776,N_5376,N_5334);
nor U5777 (N_5777,N_5352,N_5423);
nor U5778 (N_5778,N_5350,N_5588);
and U5779 (N_5779,N_5539,N_5593);
or U5780 (N_5780,N_5331,N_5417);
nor U5781 (N_5781,N_5467,N_5363);
nor U5782 (N_5782,N_5294,N_5513);
or U5783 (N_5783,N_5214,N_5520);
nor U5784 (N_5784,N_5282,N_5236);
and U5785 (N_5785,N_5325,N_5241);
nor U5786 (N_5786,N_5549,N_5570);
or U5787 (N_5787,N_5391,N_5293);
xor U5788 (N_5788,N_5324,N_5515);
or U5789 (N_5789,N_5501,N_5557);
or U5790 (N_5790,N_5344,N_5224);
nand U5791 (N_5791,N_5340,N_5307);
nand U5792 (N_5792,N_5409,N_5426);
and U5793 (N_5793,N_5429,N_5216);
and U5794 (N_5794,N_5582,N_5297);
or U5795 (N_5795,N_5585,N_5276);
nor U5796 (N_5796,N_5490,N_5594);
and U5797 (N_5797,N_5457,N_5532);
or U5798 (N_5798,N_5242,N_5274);
nand U5799 (N_5799,N_5454,N_5528);
xor U5800 (N_5800,N_5551,N_5576);
or U5801 (N_5801,N_5519,N_5545);
and U5802 (N_5802,N_5474,N_5475);
and U5803 (N_5803,N_5300,N_5591);
nor U5804 (N_5804,N_5386,N_5262);
and U5805 (N_5805,N_5358,N_5300);
nor U5806 (N_5806,N_5201,N_5392);
nand U5807 (N_5807,N_5355,N_5224);
nand U5808 (N_5808,N_5251,N_5516);
nor U5809 (N_5809,N_5325,N_5240);
and U5810 (N_5810,N_5417,N_5325);
xnor U5811 (N_5811,N_5589,N_5555);
or U5812 (N_5812,N_5227,N_5598);
and U5813 (N_5813,N_5341,N_5244);
xnor U5814 (N_5814,N_5523,N_5435);
or U5815 (N_5815,N_5317,N_5591);
nor U5816 (N_5816,N_5230,N_5485);
nand U5817 (N_5817,N_5290,N_5557);
and U5818 (N_5818,N_5577,N_5303);
or U5819 (N_5819,N_5215,N_5312);
nor U5820 (N_5820,N_5266,N_5521);
nor U5821 (N_5821,N_5223,N_5278);
nand U5822 (N_5822,N_5482,N_5249);
xnor U5823 (N_5823,N_5373,N_5386);
and U5824 (N_5824,N_5337,N_5358);
and U5825 (N_5825,N_5543,N_5373);
nand U5826 (N_5826,N_5387,N_5270);
nand U5827 (N_5827,N_5511,N_5583);
and U5828 (N_5828,N_5299,N_5237);
xnor U5829 (N_5829,N_5370,N_5347);
xor U5830 (N_5830,N_5273,N_5207);
and U5831 (N_5831,N_5515,N_5575);
xnor U5832 (N_5832,N_5568,N_5486);
and U5833 (N_5833,N_5384,N_5450);
nand U5834 (N_5834,N_5594,N_5565);
or U5835 (N_5835,N_5516,N_5574);
and U5836 (N_5836,N_5402,N_5338);
or U5837 (N_5837,N_5213,N_5239);
xor U5838 (N_5838,N_5333,N_5525);
and U5839 (N_5839,N_5204,N_5295);
and U5840 (N_5840,N_5217,N_5350);
nand U5841 (N_5841,N_5237,N_5270);
nor U5842 (N_5842,N_5218,N_5555);
xor U5843 (N_5843,N_5509,N_5306);
and U5844 (N_5844,N_5497,N_5309);
xor U5845 (N_5845,N_5200,N_5569);
nand U5846 (N_5846,N_5534,N_5300);
xnor U5847 (N_5847,N_5270,N_5293);
nand U5848 (N_5848,N_5233,N_5273);
nor U5849 (N_5849,N_5404,N_5565);
xnor U5850 (N_5850,N_5236,N_5208);
nand U5851 (N_5851,N_5326,N_5320);
nand U5852 (N_5852,N_5350,N_5586);
xor U5853 (N_5853,N_5544,N_5428);
nor U5854 (N_5854,N_5217,N_5421);
and U5855 (N_5855,N_5589,N_5523);
and U5856 (N_5856,N_5396,N_5459);
xor U5857 (N_5857,N_5520,N_5515);
or U5858 (N_5858,N_5263,N_5480);
nor U5859 (N_5859,N_5589,N_5467);
or U5860 (N_5860,N_5478,N_5239);
nand U5861 (N_5861,N_5499,N_5389);
and U5862 (N_5862,N_5333,N_5345);
nand U5863 (N_5863,N_5473,N_5591);
and U5864 (N_5864,N_5552,N_5221);
or U5865 (N_5865,N_5415,N_5471);
nand U5866 (N_5866,N_5301,N_5528);
nand U5867 (N_5867,N_5250,N_5263);
or U5868 (N_5868,N_5496,N_5525);
nand U5869 (N_5869,N_5524,N_5582);
xor U5870 (N_5870,N_5412,N_5431);
xor U5871 (N_5871,N_5518,N_5272);
nand U5872 (N_5872,N_5583,N_5273);
and U5873 (N_5873,N_5356,N_5244);
nand U5874 (N_5874,N_5487,N_5300);
xor U5875 (N_5875,N_5418,N_5382);
nor U5876 (N_5876,N_5348,N_5235);
xor U5877 (N_5877,N_5564,N_5443);
nand U5878 (N_5878,N_5446,N_5289);
nor U5879 (N_5879,N_5590,N_5381);
xor U5880 (N_5880,N_5252,N_5518);
xor U5881 (N_5881,N_5411,N_5596);
xnor U5882 (N_5882,N_5297,N_5262);
nand U5883 (N_5883,N_5347,N_5311);
xor U5884 (N_5884,N_5338,N_5209);
or U5885 (N_5885,N_5352,N_5226);
and U5886 (N_5886,N_5202,N_5384);
or U5887 (N_5887,N_5402,N_5396);
or U5888 (N_5888,N_5219,N_5547);
xnor U5889 (N_5889,N_5354,N_5504);
xnor U5890 (N_5890,N_5592,N_5425);
and U5891 (N_5891,N_5515,N_5217);
nand U5892 (N_5892,N_5506,N_5366);
nor U5893 (N_5893,N_5484,N_5491);
nor U5894 (N_5894,N_5204,N_5462);
or U5895 (N_5895,N_5366,N_5521);
nor U5896 (N_5896,N_5313,N_5230);
nand U5897 (N_5897,N_5483,N_5239);
nand U5898 (N_5898,N_5260,N_5445);
nor U5899 (N_5899,N_5385,N_5537);
xnor U5900 (N_5900,N_5212,N_5484);
nor U5901 (N_5901,N_5322,N_5264);
nor U5902 (N_5902,N_5424,N_5243);
and U5903 (N_5903,N_5327,N_5486);
nor U5904 (N_5904,N_5540,N_5557);
and U5905 (N_5905,N_5225,N_5466);
xor U5906 (N_5906,N_5471,N_5500);
xnor U5907 (N_5907,N_5590,N_5463);
nand U5908 (N_5908,N_5464,N_5330);
nor U5909 (N_5909,N_5569,N_5578);
xnor U5910 (N_5910,N_5292,N_5293);
or U5911 (N_5911,N_5262,N_5558);
xnor U5912 (N_5912,N_5339,N_5372);
or U5913 (N_5913,N_5541,N_5580);
or U5914 (N_5914,N_5326,N_5547);
nand U5915 (N_5915,N_5510,N_5396);
and U5916 (N_5916,N_5262,N_5377);
nor U5917 (N_5917,N_5519,N_5495);
xor U5918 (N_5918,N_5466,N_5461);
xnor U5919 (N_5919,N_5429,N_5225);
nor U5920 (N_5920,N_5374,N_5460);
and U5921 (N_5921,N_5218,N_5597);
xnor U5922 (N_5922,N_5263,N_5235);
nand U5923 (N_5923,N_5522,N_5226);
and U5924 (N_5924,N_5465,N_5454);
xor U5925 (N_5925,N_5251,N_5336);
or U5926 (N_5926,N_5463,N_5454);
nor U5927 (N_5927,N_5215,N_5509);
nor U5928 (N_5928,N_5319,N_5354);
xor U5929 (N_5929,N_5400,N_5286);
and U5930 (N_5930,N_5350,N_5341);
and U5931 (N_5931,N_5442,N_5567);
nor U5932 (N_5932,N_5547,N_5557);
xnor U5933 (N_5933,N_5238,N_5518);
xor U5934 (N_5934,N_5218,N_5248);
xnor U5935 (N_5935,N_5332,N_5512);
or U5936 (N_5936,N_5280,N_5276);
nor U5937 (N_5937,N_5242,N_5460);
nor U5938 (N_5938,N_5445,N_5492);
xor U5939 (N_5939,N_5445,N_5382);
or U5940 (N_5940,N_5448,N_5239);
and U5941 (N_5941,N_5351,N_5488);
nand U5942 (N_5942,N_5454,N_5506);
nor U5943 (N_5943,N_5279,N_5542);
and U5944 (N_5944,N_5381,N_5502);
xor U5945 (N_5945,N_5555,N_5312);
xnor U5946 (N_5946,N_5322,N_5405);
or U5947 (N_5947,N_5373,N_5446);
and U5948 (N_5948,N_5342,N_5375);
and U5949 (N_5949,N_5479,N_5520);
nor U5950 (N_5950,N_5517,N_5262);
nand U5951 (N_5951,N_5445,N_5268);
and U5952 (N_5952,N_5295,N_5552);
nand U5953 (N_5953,N_5273,N_5332);
xor U5954 (N_5954,N_5521,N_5341);
xor U5955 (N_5955,N_5385,N_5423);
or U5956 (N_5956,N_5332,N_5266);
and U5957 (N_5957,N_5386,N_5591);
or U5958 (N_5958,N_5438,N_5363);
nor U5959 (N_5959,N_5546,N_5495);
or U5960 (N_5960,N_5570,N_5362);
nor U5961 (N_5961,N_5261,N_5389);
and U5962 (N_5962,N_5316,N_5320);
or U5963 (N_5963,N_5455,N_5341);
or U5964 (N_5964,N_5562,N_5275);
xnor U5965 (N_5965,N_5247,N_5445);
nand U5966 (N_5966,N_5308,N_5453);
nand U5967 (N_5967,N_5595,N_5489);
and U5968 (N_5968,N_5388,N_5593);
nor U5969 (N_5969,N_5202,N_5530);
nand U5970 (N_5970,N_5454,N_5428);
nor U5971 (N_5971,N_5430,N_5517);
or U5972 (N_5972,N_5417,N_5537);
xnor U5973 (N_5973,N_5441,N_5351);
xnor U5974 (N_5974,N_5429,N_5299);
or U5975 (N_5975,N_5218,N_5489);
nand U5976 (N_5976,N_5565,N_5481);
or U5977 (N_5977,N_5292,N_5551);
nand U5978 (N_5978,N_5535,N_5207);
nor U5979 (N_5979,N_5486,N_5299);
and U5980 (N_5980,N_5277,N_5222);
nor U5981 (N_5981,N_5416,N_5356);
xor U5982 (N_5982,N_5468,N_5305);
nor U5983 (N_5983,N_5582,N_5375);
xnor U5984 (N_5984,N_5516,N_5597);
xnor U5985 (N_5985,N_5354,N_5200);
nor U5986 (N_5986,N_5547,N_5489);
xnor U5987 (N_5987,N_5568,N_5278);
nor U5988 (N_5988,N_5219,N_5247);
xor U5989 (N_5989,N_5202,N_5428);
and U5990 (N_5990,N_5593,N_5577);
nor U5991 (N_5991,N_5592,N_5342);
xnor U5992 (N_5992,N_5548,N_5235);
xor U5993 (N_5993,N_5340,N_5391);
xnor U5994 (N_5994,N_5202,N_5445);
nand U5995 (N_5995,N_5565,N_5368);
nor U5996 (N_5996,N_5516,N_5438);
or U5997 (N_5997,N_5436,N_5518);
nand U5998 (N_5998,N_5526,N_5464);
nor U5999 (N_5999,N_5549,N_5362);
nand U6000 (N_6000,N_5918,N_5715);
and U6001 (N_6001,N_5938,N_5789);
or U6002 (N_6002,N_5945,N_5620);
nand U6003 (N_6003,N_5639,N_5985);
xnor U6004 (N_6004,N_5832,N_5726);
nand U6005 (N_6005,N_5681,N_5793);
and U6006 (N_6006,N_5716,N_5728);
nor U6007 (N_6007,N_5643,N_5846);
or U6008 (N_6008,N_5827,N_5625);
xor U6009 (N_6009,N_5676,N_5954);
xnor U6010 (N_6010,N_5952,N_5914);
and U6011 (N_6011,N_5934,N_5656);
nand U6012 (N_6012,N_5764,N_5910);
or U6013 (N_6013,N_5919,N_5750);
or U6014 (N_6014,N_5886,N_5966);
nand U6015 (N_6015,N_5733,N_5790);
or U6016 (N_6016,N_5937,N_5761);
xnor U6017 (N_6017,N_5927,N_5714);
nor U6018 (N_6018,N_5976,N_5612);
and U6019 (N_6019,N_5654,N_5608);
xnor U6020 (N_6020,N_5932,N_5663);
and U6021 (N_6021,N_5812,N_5863);
nand U6022 (N_6022,N_5775,N_5951);
nand U6023 (N_6023,N_5783,N_5967);
nor U6024 (N_6024,N_5854,N_5978);
or U6025 (N_6025,N_5893,N_5792);
and U6026 (N_6026,N_5756,N_5707);
or U6027 (N_6027,N_5963,N_5920);
xor U6028 (N_6028,N_5653,N_5844);
or U6029 (N_6029,N_5680,N_5923);
and U6030 (N_6030,N_5641,N_5839);
xnor U6031 (N_6031,N_5852,N_5767);
and U6032 (N_6032,N_5743,N_5867);
nand U6033 (N_6033,N_5644,N_5701);
or U6034 (N_6034,N_5662,N_5755);
nor U6035 (N_6035,N_5882,N_5618);
nand U6036 (N_6036,N_5787,N_5794);
or U6037 (N_6037,N_5982,N_5878);
nor U6038 (N_6038,N_5961,N_5947);
nor U6039 (N_6039,N_5980,N_5725);
nand U6040 (N_6040,N_5722,N_5710);
nand U6041 (N_6041,N_5779,N_5685);
xnor U6042 (N_6042,N_5753,N_5697);
xnor U6043 (N_6043,N_5890,N_5774);
nor U6044 (N_6044,N_5782,N_5666);
or U6045 (N_6045,N_5968,N_5816);
xor U6046 (N_6046,N_5862,N_5994);
nand U6047 (N_6047,N_5781,N_5622);
xor U6048 (N_6048,N_5823,N_5996);
and U6049 (N_6049,N_5704,N_5788);
nand U6050 (N_6050,N_5702,N_5671);
or U6051 (N_6051,N_5944,N_5640);
or U6052 (N_6052,N_5721,N_5977);
nand U6053 (N_6053,N_5864,N_5695);
nor U6054 (N_6054,N_5965,N_5845);
xor U6055 (N_6055,N_5684,N_5858);
or U6056 (N_6056,N_5892,N_5732);
nand U6057 (N_6057,N_5989,N_5628);
and U6058 (N_6058,N_5931,N_5830);
nand U6059 (N_6059,N_5807,N_5682);
nand U6060 (N_6060,N_5942,N_5616);
and U6061 (N_6061,N_5703,N_5757);
xnor U6062 (N_6062,N_5777,N_5820);
nand U6063 (N_6063,N_5879,N_5896);
xnor U6064 (N_6064,N_5635,N_5804);
and U6065 (N_6065,N_5699,N_5999);
or U6066 (N_6066,N_5948,N_5691);
xnor U6067 (N_6067,N_5835,N_5751);
xor U6068 (N_6068,N_5766,N_5650);
and U6069 (N_6069,N_5621,N_5953);
xnor U6070 (N_6070,N_5856,N_5669);
nand U6071 (N_6071,N_5667,N_5773);
and U6072 (N_6072,N_5799,N_5609);
nand U6073 (N_6073,N_5670,N_5824);
and U6074 (N_6074,N_5984,N_5649);
nor U6075 (N_6075,N_5801,N_5747);
and U6076 (N_6076,N_5729,N_5655);
xnor U6077 (N_6077,N_5922,N_5795);
nand U6078 (N_6078,N_5958,N_5611);
nor U6079 (N_6079,N_5717,N_5735);
and U6080 (N_6080,N_5908,N_5836);
and U6081 (N_6081,N_5632,N_5797);
and U6082 (N_6082,N_5855,N_5642);
nor U6083 (N_6083,N_5638,N_5817);
or U6084 (N_6084,N_5819,N_5913);
or U6085 (N_6085,N_5897,N_5689);
or U6086 (N_6086,N_5739,N_5969);
and U6087 (N_6087,N_5939,N_5718);
or U6088 (N_6088,N_5905,N_5708);
or U6089 (N_6089,N_5636,N_5730);
or U6090 (N_6090,N_5902,N_5615);
and U6091 (N_6091,N_5860,N_5895);
nand U6092 (N_6092,N_5724,N_5916);
nand U6093 (N_6093,N_5623,N_5674);
nor U6094 (N_6094,N_5678,N_5917);
nand U6095 (N_6095,N_5759,N_5872);
nor U6096 (N_6096,N_5894,N_5776);
xor U6097 (N_6097,N_5601,N_5745);
and U6098 (N_6098,N_5847,N_5972);
xnor U6099 (N_6099,N_5613,N_5979);
xor U6100 (N_6100,N_5758,N_5778);
nor U6101 (N_6101,N_5696,N_5837);
or U6102 (N_6102,N_5749,N_5617);
nor U6103 (N_6103,N_5828,N_5687);
and U6104 (N_6104,N_5762,N_5626);
and U6105 (N_6105,N_5677,N_5970);
or U6106 (N_6106,N_5850,N_5711);
nand U6107 (N_6107,N_5734,N_5990);
nand U6108 (N_6108,N_5698,N_5813);
and U6109 (N_6109,N_5898,N_5818);
and U6110 (N_6110,N_5763,N_5881);
xor U6111 (N_6111,N_5808,N_5851);
and U6112 (N_6112,N_5853,N_5675);
or U6113 (N_6113,N_5815,N_5974);
xnor U6114 (N_6114,N_5859,N_5690);
or U6115 (N_6115,N_5796,N_5809);
or U6116 (N_6116,N_5993,N_5936);
or U6117 (N_6117,N_5800,N_5912);
xnor U6118 (N_6118,N_5737,N_5605);
or U6119 (N_6119,N_5805,N_5709);
and U6120 (N_6120,N_5744,N_5803);
xnor U6121 (N_6121,N_5873,N_5814);
nor U6122 (N_6122,N_5768,N_5903);
nor U6123 (N_6123,N_5700,N_5624);
nor U6124 (N_6124,N_5991,N_5838);
nand U6125 (N_6125,N_5810,N_5772);
xnor U6126 (N_6126,N_5664,N_5825);
or U6127 (N_6127,N_5865,N_5712);
nor U6128 (N_6128,N_5652,N_5998);
xnor U6129 (N_6129,N_5741,N_5798);
nor U6130 (N_6130,N_5889,N_5926);
nand U6131 (N_6131,N_5885,N_5975);
or U6132 (N_6132,N_5651,N_5658);
xor U6133 (N_6133,N_5752,N_5771);
or U6134 (N_6134,N_5887,N_5986);
and U6135 (N_6135,N_5940,N_5962);
or U6136 (N_6136,N_5811,N_5871);
and U6137 (N_6137,N_5627,N_5740);
and U6138 (N_6138,N_5924,N_5769);
xnor U6139 (N_6139,N_5992,N_5604);
nand U6140 (N_6140,N_5935,N_5692);
xnor U6141 (N_6141,N_5907,N_5848);
xor U6142 (N_6142,N_5672,N_5802);
nand U6143 (N_6143,N_5899,N_5876);
nand U6144 (N_6144,N_5949,N_5706);
xor U6145 (N_6145,N_5646,N_5875);
xor U6146 (N_6146,N_5600,N_5720);
and U6147 (N_6147,N_5874,N_5660);
or U6148 (N_6148,N_5693,N_5806);
and U6149 (N_6149,N_5956,N_5833);
or U6150 (N_6150,N_5665,N_5971);
xor U6151 (N_6151,N_5957,N_5668);
and U6152 (N_6152,N_5888,N_5713);
and U6153 (N_6153,N_5880,N_5904);
xnor U6154 (N_6154,N_5857,N_5829);
xor U6155 (N_6155,N_5964,N_5821);
and U6156 (N_6156,N_5661,N_5941);
nor U6157 (N_6157,N_5633,N_5987);
and U6158 (N_6158,N_5694,N_5784);
or U6159 (N_6159,N_5915,N_5770);
or U6160 (N_6160,N_5955,N_5647);
or U6161 (N_6161,N_5765,N_5719);
xnor U6162 (N_6162,N_5929,N_5849);
nor U6163 (N_6163,N_5603,N_5826);
xor U6164 (N_6164,N_5995,N_5925);
and U6165 (N_6165,N_5909,N_5731);
and U6166 (N_6166,N_5883,N_5746);
nand U6167 (N_6167,N_5629,N_5610);
nor U6168 (N_6168,N_5866,N_5631);
nor U6169 (N_6169,N_5831,N_5997);
or U6170 (N_6170,N_5602,N_5921);
and U6171 (N_6171,N_5841,N_5900);
or U6172 (N_6172,N_5630,N_5933);
nand U6173 (N_6173,N_5614,N_5748);
nand U6174 (N_6174,N_5843,N_5869);
nor U6175 (N_6175,N_5679,N_5760);
and U6176 (N_6176,N_5657,N_5950);
xnor U6177 (N_6177,N_5930,N_5928);
and U6178 (N_6178,N_5959,N_5705);
or U6179 (N_6179,N_5637,N_5736);
or U6180 (N_6180,N_5983,N_5988);
nor U6181 (N_6181,N_5911,N_5981);
nand U6182 (N_6182,N_5742,N_5786);
xnor U6183 (N_6183,N_5738,N_5973);
nor U6184 (N_6184,N_5884,N_5688);
and U6185 (N_6185,N_5607,N_5891);
nand U6186 (N_6186,N_5606,N_5946);
or U6187 (N_6187,N_5842,N_5870);
and U6188 (N_6188,N_5785,N_5901);
nand U6189 (N_6189,N_5906,N_5791);
xnor U6190 (N_6190,N_5754,N_5861);
and U6191 (N_6191,N_5673,N_5960);
nand U6192 (N_6192,N_5943,N_5877);
nor U6193 (N_6193,N_5723,N_5822);
or U6194 (N_6194,N_5868,N_5780);
and U6195 (N_6195,N_5834,N_5645);
xnor U6196 (N_6196,N_5686,N_5840);
or U6197 (N_6197,N_5727,N_5683);
nand U6198 (N_6198,N_5659,N_5648);
nor U6199 (N_6199,N_5634,N_5619);
or U6200 (N_6200,N_5744,N_5828);
or U6201 (N_6201,N_5657,N_5809);
nand U6202 (N_6202,N_5957,N_5989);
xor U6203 (N_6203,N_5925,N_5816);
nor U6204 (N_6204,N_5738,N_5777);
and U6205 (N_6205,N_5856,N_5664);
xnor U6206 (N_6206,N_5873,N_5902);
nand U6207 (N_6207,N_5980,N_5606);
nand U6208 (N_6208,N_5815,N_5716);
xnor U6209 (N_6209,N_5656,N_5791);
xnor U6210 (N_6210,N_5712,N_5994);
nor U6211 (N_6211,N_5904,N_5615);
or U6212 (N_6212,N_5664,N_5635);
nor U6213 (N_6213,N_5648,N_5958);
nor U6214 (N_6214,N_5703,N_5943);
nor U6215 (N_6215,N_5723,N_5954);
nand U6216 (N_6216,N_5873,N_5669);
and U6217 (N_6217,N_5843,N_5649);
nand U6218 (N_6218,N_5677,N_5781);
and U6219 (N_6219,N_5902,N_5820);
xor U6220 (N_6220,N_5703,N_5889);
nand U6221 (N_6221,N_5997,N_5865);
nor U6222 (N_6222,N_5624,N_5965);
or U6223 (N_6223,N_5688,N_5965);
nor U6224 (N_6224,N_5710,N_5655);
nand U6225 (N_6225,N_5968,N_5991);
nand U6226 (N_6226,N_5907,N_5884);
xnor U6227 (N_6227,N_5723,N_5646);
nor U6228 (N_6228,N_5838,N_5743);
nand U6229 (N_6229,N_5859,N_5993);
nand U6230 (N_6230,N_5652,N_5960);
or U6231 (N_6231,N_5769,N_5980);
and U6232 (N_6232,N_5870,N_5888);
or U6233 (N_6233,N_5980,N_5696);
and U6234 (N_6234,N_5719,N_5891);
nor U6235 (N_6235,N_5949,N_5649);
nand U6236 (N_6236,N_5604,N_5954);
and U6237 (N_6237,N_5751,N_5729);
nor U6238 (N_6238,N_5628,N_5631);
nand U6239 (N_6239,N_5646,N_5823);
and U6240 (N_6240,N_5815,N_5623);
and U6241 (N_6241,N_5798,N_5619);
nand U6242 (N_6242,N_5964,N_5626);
nor U6243 (N_6243,N_5967,N_5855);
or U6244 (N_6244,N_5934,N_5827);
nand U6245 (N_6245,N_5969,N_5789);
nand U6246 (N_6246,N_5770,N_5828);
nand U6247 (N_6247,N_5678,N_5612);
nand U6248 (N_6248,N_5634,N_5890);
and U6249 (N_6249,N_5772,N_5850);
and U6250 (N_6250,N_5819,N_5635);
nand U6251 (N_6251,N_5660,N_5624);
and U6252 (N_6252,N_5951,N_5815);
xnor U6253 (N_6253,N_5751,N_5756);
nand U6254 (N_6254,N_5626,N_5610);
xor U6255 (N_6255,N_5977,N_5745);
nand U6256 (N_6256,N_5680,N_5709);
xor U6257 (N_6257,N_5813,N_5677);
nand U6258 (N_6258,N_5675,N_5791);
nand U6259 (N_6259,N_5876,N_5910);
nor U6260 (N_6260,N_5709,N_5886);
nand U6261 (N_6261,N_5769,N_5925);
nand U6262 (N_6262,N_5939,N_5620);
and U6263 (N_6263,N_5978,N_5666);
nor U6264 (N_6264,N_5648,N_5953);
nor U6265 (N_6265,N_5630,N_5760);
xor U6266 (N_6266,N_5930,N_5612);
or U6267 (N_6267,N_5770,N_5820);
nor U6268 (N_6268,N_5810,N_5823);
or U6269 (N_6269,N_5600,N_5630);
nor U6270 (N_6270,N_5709,N_5751);
and U6271 (N_6271,N_5773,N_5672);
or U6272 (N_6272,N_5721,N_5867);
nand U6273 (N_6273,N_5735,N_5984);
nor U6274 (N_6274,N_5856,N_5831);
nand U6275 (N_6275,N_5877,N_5803);
or U6276 (N_6276,N_5955,N_5632);
and U6277 (N_6277,N_5609,N_5994);
or U6278 (N_6278,N_5645,N_5930);
or U6279 (N_6279,N_5763,N_5756);
and U6280 (N_6280,N_5707,N_5603);
or U6281 (N_6281,N_5631,N_5683);
nand U6282 (N_6282,N_5675,N_5768);
or U6283 (N_6283,N_5938,N_5864);
or U6284 (N_6284,N_5824,N_5765);
and U6285 (N_6285,N_5832,N_5676);
nor U6286 (N_6286,N_5723,N_5933);
xor U6287 (N_6287,N_5603,N_5851);
or U6288 (N_6288,N_5650,N_5710);
and U6289 (N_6289,N_5642,N_5643);
nand U6290 (N_6290,N_5803,N_5970);
nor U6291 (N_6291,N_5712,N_5680);
nand U6292 (N_6292,N_5859,N_5898);
nand U6293 (N_6293,N_5741,N_5643);
xor U6294 (N_6294,N_5990,N_5994);
or U6295 (N_6295,N_5881,N_5740);
xnor U6296 (N_6296,N_5924,N_5968);
or U6297 (N_6297,N_5611,N_5725);
nor U6298 (N_6298,N_5636,N_5783);
xor U6299 (N_6299,N_5830,N_5969);
and U6300 (N_6300,N_5991,N_5696);
nor U6301 (N_6301,N_5867,N_5672);
xor U6302 (N_6302,N_5667,N_5988);
nor U6303 (N_6303,N_5727,N_5967);
and U6304 (N_6304,N_5679,N_5891);
or U6305 (N_6305,N_5870,N_5875);
xor U6306 (N_6306,N_5911,N_5719);
or U6307 (N_6307,N_5852,N_5961);
or U6308 (N_6308,N_5989,N_5842);
xnor U6309 (N_6309,N_5757,N_5815);
or U6310 (N_6310,N_5879,N_5981);
or U6311 (N_6311,N_5705,N_5600);
and U6312 (N_6312,N_5990,N_5613);
nor U6313 (N_6313,N_5900,N_5970);
nor U6314 (N_6314,N_5973,N_5682);
xor U6315 (N_6315,N_5856,N_5791);
nor U6316 (N_6316,N_5864,N_5933);
nor U6317 (N_6317,N_5620,N_5608);
or U6318 (N_6318,N_5668,N_5697);
or U6319 (N_6319,N_5763,N_5918);
or U6320 (N_6320,N_5941,N_5870);
or U6321 (N_6321,N_5821,N_5850);
xor U6322 (N_6322,N_5698,N_5968);
nand U6323 (N_6323,N_5822,N_5767);
nor U6324 (N_6324,N_5615,N_5759);
or U6325 (N_6325,N_5781,N_5745);
nor U6326 (N_6326,N_5712,N_5693);
xnor U6327 (N_6327,N_5887,N_5821);
nor U6328 (N_6328,N_5900,N_5960);
nor U6329 (N_6329,N_5795,N_5796);
nor U6330 (N_6330,N_5679,N_5852);
nand U6331 (N_6331,N_5639,N_5938);
nor U6332 (N_6332,N_5981,N_5901);
nand U6333 (N_6333,N_5708,N_5639);
nand U6334 (N_6334,N_5628,N_5867);
xor U6335 (N_6335,N_5748,N_5705);
or U6336 (N_6336,N_5848,N_5965);
and U6337 (N_6337,N_5740,N_5977);
nor U6338 (N_6338,N_5750,N_5698);
nand U6339 (N_6339,N_5654,N_5704);
or U6340 (N_6340,N_5968,N_5691);
nor U6341 (N_6341,N_5741,N_5810);
or U6342 (N_6342,N_5688,N_5863);
xor U6343 (N_6343,N_5863,N_5740);
and U6344 (N_6344,N_5907,N_5952);
and U6345 (N_6345,N_5651,N_5676);
and U6346 (N_6346,N_5943,N_5947);
or U6347 (N_6347,N_5816,N_5769);
nand U6348 (N_6348,N_5989,N_5790);
xor U6349 (N_6349,N_5989,N_5777);
nor U6350 (N_6350,N_5742,N_5912);
nor U6351 (N_6351,N_5952,N_5786);
or U6352 (N_6352,N_5664,N_5621);
nand U6353 (N_6353,N_5853,N_5719);
and U6354 (N_6354,N_5904,N_5791);
xnor U6355 (N_6355,N_5764,N_5619);
or U6356 (N_6356,N_5777,N_5727);
xor U6357 (N_6357,N_5653,N_5805);
nand U6358 (N_6358,N_5874,N_5855);
xor U6359 (N_6359,N_5781,N_5820);
nand U6360 (N_6360,N_5736,N_5859);
xnor U6361 (N_6361,N_5939,N_5850);
or U6362 (N_6362,N_5952,N_5855);
nor U6363 (N_6363,N_5888,N_5656);
nand U6364 (N_6364,N_5730,N_5715);
and U6365 (N_6365,N_5983,N_5721);
xor U6366 (N_6366,N_5669,N_5708);
or U6367 (N_6367,N_5855,N_5727);
nand U6368 (N_6368,N_5640,N_5822);
and U6369 (N_6369,N_5869,N_5929);
or U6370 (N_6370,N_5690,N_5831);
nand U6371 (N_6371,N_5857,N_5684);
nand U6372 (N_6372,N_5893,N_5610);
nand U6373 (N_6373,N_5754,N_5794);
nand U6374 (N_6374,N_5603,N_5706);
or U6375 (N_6375,N_5701,N_5758);
or U6376 (N_6376,N_5624,N_5913);
and U6377 (N_6377,N_5998,N_5630);
and U6378 (N_6378,N_5791,N_5690);
nor U6379 (N_6379,N_5644,N_5967);
or U6380 (N_6380,N_5679,N_5771);
or U6381 (N_6381,N_5712,N_5797);
xnor U6382 (N_6382,N_5701,N_5926);
xor U6383 (N_6383,N_5914,N_5902);
nand U6384 (N_6384,N_5969,N_5708);
nor U6385 (N_6385,N_5696,N_5761);
nand U6386 (N_6386,N_5600,N_5803);
nor U6387 (N_6387,N_5979,N_5625);
or U6388 (N_6388,N_5864,N_5903);
and U6389 (N_6389,N_5683,N_5853);
nor U6390 (N_6390,N_5895,N_5631);
nor U6391 (N_6391,N_5817,N_5715);
xnor U6392 (N_6392,N_5647,N_5839);
nor U6393 (N_6393,N_5862,N_5817);
xnor U6394 (N_6394,N_5675,N_5700);
xor U6395 (N_6395,N_5719,N_5908);
xor U6396 (N_6396,N_5771,N_5616);
and U6397 (N_6397,N_5813,N_5955);
xor U6398 (N_6398,N_5753,N_5835);
or U6399 (N_6399,N_5843,N_5815);
nand U6400 (N_6400,N_6223,N_6160);
xnor U6401 (N_6401,N_6140,N_6288);
or U6402 (N_6402,N_6343,N_6182);
nor U6403 (N_6403,N_6279,N_6185);
nand U6404 (N_6404,N_6148,N_6016);
nor U6405 (N_6405,N_6026,N_6013);
and U6406 (N_6406,N_6225,N_6335);
nor U6407 (N_6407,N_6123,N_6001);
nor U6408 (N_6408,N_6040,N_6371);
and U6409 (N_6409,N_6051,N_6125);
and U6410 (N_6410,N_6360,N_6150);
and U6411 (N_6411,N_6075,N_6263);
xnor U6412 (N_6412,N_6242,N_6137);
xor U6413 (N_6413,N_6029,N_6337);
xor U6414 (N_6414,N_6107,N_6091);
or U6415 (N_6415,N_6264,N_6329);
and U6416 (N_6416,N_6277,N_6077);
xnor U6417 (N_6417,N_6196,N_6094);
or U6418 (N_6418,N_6060,N_6308);
xor U6419 (N_6419,N_6202,N_6230);
or U6420 (N_6420,N_6383,N_6267);
nand U6421 (N_6421,N_6227,N_6188);
xnor U6422 (N_6422,N_6251,N_6324);
or U6423 (N_6423,N_6216,N_6306);
xnor U6424 (N_6424,N_6376,N_6278);
and U6425 (N_6425,N_6393,N_6276);
and U6426 (N_6426,N_6363,N_6214);
and U6427 (N_6427,N_6255,N_6061);
or U6428 (N_6428,N_6020,N_6390);
nand U6429 (N_6429,N_6133,N_6023);
nand U6430 (N_6430,N_6378,N_6240);
or U6431 (N_6431,N_6028,N_6122);
nor U6432 (N_6432,N_6351,N_6395);
and U6433 (N_6433,N_6114,N_6284);
and U6434 (N_6434,N_6187,N_6340);
or U6435 (N_6435,N_6300,N_6036);
nor U6436 (N_6436,N_6174,N_6008);
nor U6437 (N_6437,N_6256,N_6235);
xnor U6438 (N_6438,N_6167,N_6101);
or U6439 (N_6439,N_6171,N_6043);
nor U6440 (N_6440,N_6072,N_6195);
or U6441 (N_6441,N_6206,N_6283);
xnor U6442 (N_6442,N_6233,N_6361);
nand U6443 (N_6443,N_6117,N_6321);
or U6444 (N_6444,N_6076,N_6350);
and U6445 (N_6445,N_6213,N_6247);
and U6446 (N_6446,N_6204,N_6320);
or U6447 (N_6447,N_6323,N_6170);
nor U6448 (N_6448,N_6069,N_6012);
or U6449 (N_6449,N_6237,N_6151);
xor U6450 (N_6450,N_6319,N_6241);
and U6451 (N_6451,N_6193,N_6175);
and U6452 (N_6452,N_6358,N_6136);
or U6453 (N_6453,N_6146,N_6292);
xnor U6454 (N_6454,N_6038,N_6231);
or U6455 (N_6455,N_6302,N_6249);
xor U6456 (N_6456,N_6134,N_6236);
nor U6457 (N_6457,N_6070,N_6342);
or U6458 (N_6458,N_6352,N_6131);
and U6459 (N_6459,N_6368,N_6312);
nor U6460 (N_6460,N_6296,N_6304);
xnor U6461 (N_6461,N_6111,N_6128);
nand U6462 (N_6462,N_6387,N_6041);
xor U6463 (N_6463,N_6313,N_6258);
xnor U6464 (N_6464,N_6156,N_6215);
xor U6465 (N_6465,N_6092,N_6135);
nand U6466 (N_6466,N_6210,N_6115);
or U6467 (N_6467,N_6021,N_6058);
nand U6468 (N_6468,N_6341,N_6275);
nor U6469 (N_6469,N_6222,N_6373);
xor U6470 (N_6470,N_6093,N_6142);
nor U6471 (N_6471,N_6253,N_6153);
nand U6472 (N_6472,N_6130,N_6050);
nor U6473 (N_6473,N_6157,N_6095);
nor U6474 (N_6474,N_6143,N_6113);
nand U6475 (N_6475,N_6310,N_6207);
nand U6476 (N_6476,N_6318,N_6333);
or U6477 (N_6477,N_6252,N_6208);
xnor U6478 (N_6478,N_6190,N_6357);
xor U6479 (N_6479,N_6211,N_6392);
nand U6480 (N_6480,N_6014,N_6224);
and U6481 (N_6481,N_6099,N_6010);
xnor U6482 (N_6482,N_6067,N_6221);
nand U6483 (N_6483,N_6019,N_6355);
nor U6484 (N_6484,N_6159,N_6141);
xnor U6485 (N_6485,N_6299,N_6062);
or U6486 (N_6486,N_6078,N_6248);
xnor U6487 (N_6487,N_6176,N_6068);
nor U6488 (N_6488,N_6180,N_6003);
and U6489 (N_6489,N_6025,N_6367);
and U6490 (N_6490,N_6163,N_6269);
xnor U6491 (N_6491,N_6109,N_6005);
nand U6492 (N_6492,N_6042,N_6152);
xor U6493 (N_6493,N_6045,N_6246);
nor U6494 (N_6494,N_6239,N_6178);
nand U6495 (N_6495,N_6238,N_6369);
or U6496 (N_6496,N_6126,N_6127);
nor U6497 (N_6497,N_6243,N_6348);
nor U6498 (N_6498,N_6226,N_6098);
or U6499 (N_6499,N_6183,N_6086);
and U6500 (N_6500,N_6220,N_6089);
xor U6501 (N_6501,N_6106,N_6017);
nor U6502 (N_6502,N_6228,N_6200);
nand U6503 (N_6503,N_6124,N_6071);
or U6504 (N_6504,N_6262,N_6347);
nor U6505 (N_6505,N_6203,N_6388);
nor U6506 (N_6506,N_6100,N_6311);
nor U6507 (N_6507,N_6389,N_6194);
nand U6508 (N_6508,N_6287,N_6108);
or U6509 (N_6509,N_6049,N_6359);
xnor U6510 (N_6510,N_6129,N_6336);
or U6511 (N_6511,N_6011,N_6074);
nor U6512 (N_6512,N_6334,N_6059);
xor U6513 (N_6513,N_6349,N_6365);
and U6514 (N_6514,N_6166,N_6007);
xnor U6515 (N_6515,N_6332,N_6268);
xnor U6516 (N_6516,N_6346,N_6073);
and U6517 (N_6517,N_6305,N_6046);
xnor U6518 (N_6518,N_6328,N_6009);
nand U6519 (N_6519,N_6186,N_6102);
nor U6520 (N_6520,N_6118,N_6282);
xnor U6521 (N_6521,N_6285,N_6055);
and U6522 (N_6522,N_6212,N_6172);
and U6523 (N_6523,N_6066,N_6165);
xor U6524 (N_6524,N_6197,N_6006);
nand U6525 (N_6525,N_6034,N_6381);
or U6526 (N_6526,N_6022,N_6338);
nand U6527 (N_6527,N_6382,N_6398);
nor U6528 (N_6528,N_6030,N_6104);
xor U6529 (N_6529,N_6326,N_6037);
or U6530 (N_6530,N_6052,N_6158);
xor U6531 (N_6531,N_6265,N_6177);
xor U6532 (N_6532,N_6139,N_6082);
xnor U6533 (N_6533,N_6274,N_6260);
nand U6534 (N_6534,N_6110,N_6027);
nor U6535 (N_6535,N_6147,N_6144);
or U6536 (N_6536,N_6374,N_6096);
nand U6537 (N_6537,N_6002,N_6353);
and U6538 (N_6538,N_6257,N_6377);
nand U6539 (N_6539,N_6245,N_6372);
or U6540 (N_6540,N_6386,N_6391);
xor U6541 (N_6541,N_6217,N_6132);
nand U6542 (N_6542,N_6314,N_6331);
and U6543 (N_6543,N_6293,N_6081);
nand U6544 (N_6544,N_6024,N_6344);
xnor U6545 (N_6545,N_6219,N_6315);
nand U6546 (N_6546,N_6063,N_6205);
nor U6547 (N_6547,N_6270,N_6317);
nand U6548 (N_6548,N_6362,N_6339);
or U6549 (N_6549,N_6281,N_6154);
xnor U6550 (N_6550,N_6032,N_6090);
and U6551 (N_6551,N_6120,N_6316);
nor U6552 (N_6552,N_6057,N_6149);
nand U6553 (N_6553,N_6330,N_6250);
xor U6554 (N_6554,N_6015,N_6162);
or U6555 (N_6555,N_6356,N_6272);
or U6556 (N_6556,N_6198,N_6087);
xnor U6557 (N_6557,N_6169,N_6004);
and U6558 (N_6558,N_6181,N_6105);
and U6559 (N_6559,N_6103,N_6271);
and U6560 (N_6560,N_6201,N_6121);
xnor U6561 (N_6561,N_6192,N_6083);
nor U6562 (N_6562,N_6259,N_6327);
xor U6563 (N_6563,N_6385,N_6053);
nand U6564 (N_6564,N_6065,N_6218);
or U6565 (N_6565,N_6261,N_6097);
and U6566 (N_6566,N_6375,N_6229);
xnor U6567 (N_6567,N_6379,N_6184);
or U6568 (N_6568,N_6085,N_6254);
nor U6569 (N_6569,N_6384,N_6039);
or U6570 (N_6570,N_6168,N_6345);
and U6571 (N_6571,N_6084,N_6088);
or U6572 (N_6572,N_6054,N_6145);
and U6573 (N_6573,N_6179,N_6380);
xnor U6574 (N_6574,N_6164,N_6370);
or U6575 (N_6575,N_6294,N_6394);
xor U6576 (N_6576,N_6119,N_6286);
or U6577 (N_6577,N_6232,N_6366);
nor U6578 (N_6578,N_6325,N_6301);
nor U6579 (N_6579,N_6161,N_6033);
or U6580 (N_6580,N_6173,N_6018);
and U6581 (N_6581,N_6116,N_6399);
nor U6582 (N_6582,N_6189,N_6079);
and U6583 (N_6583,N_6322,N_6191);
or U6584 (N_6584,N_6298,N_6199);
or U6585 (N_6585,N_6266,N_6396);
or U6586 (N_6586,N_6234,N_6397);
nor U6587 (N_6587,N_6354,N_6047);
and U6588 (N_6588,N_6295,N_6290);
xnor U6589 (N_6589,N_6307,N_6273);
nor U6590 (N_6590,N_6138,N_6244);
or U6591 (N_6591,N_6080,N_6297);
nor U6592 (N_6592,N_6031,N_6280);
or U6593 (N_6593,N_6056,N_6155);
nand U6594 (N_6594,N_6064,N_6000);
nor U6595 (N_6595,N_6364,N_6048);
xnor U6596 (N_6596,N_6303,N_6309);
or U6597 (N_6597,N_6112,N_6209);
and U6598 (N_6598,N_6291,N_6044);
nand U6599 (N_6599,N_6035,N_6289);
nor U6600 (N_6600,N_6062,N_6378);
xor U6601 (N_6601,N_6061,N_6064);
and U6602 (N_6602,N_6301,N_6156);
nor U6603 (N_6603,N_6087,N_6186);
or U6604 (N_6604,N_6050,N_6029);
or U6605 (N_6605,N_6224,N_6255);
or U6606 (N_6606,N_6252,N_6356);
nand U6607 (N_6607,N_6056,N_6342);
or U6608 (N_6608,N_6068,N_6251);
or U6609 (N_6609,N_6186,N_6161);
nand U6610 (N_6610,N_6257,N_6032);
or U6611 (N_6611,N_6277,N_6315);
nor U6612 (N_6612,N_6306,N_6322);
nand U6613 (N_6613,N_6199,N_6321);
nor U6614 (N_6614,N_6017,N_6244);
nor U6615 (N_6615,N_6076,N_6255);
nor U6616 (N_6616,N_6376,N_6079);
nand U6617 (N_6617,N_6208,N_6071);
nor U6618 (N_6618,N_6196,N_6356);
or U6619 (N_6619,N_6205,N_6316);
or U6620 (N_6620,N_6254,N_6174);
xnor U6621 (N_6621,N_6085,N_6228);
and U6622 (N_6622,N_6380,N_6214);
nor U6623 (N_6623,N_6081,N_6134);
and U6624 (N_6624,N_6030,N_6006);
or U6625 (N_6625,N_6119,N_6126);
nor U6626 (N_6626,N_6244,N_6127);
nand U6627 (N_6627,N_6039,N_6011);
or U6628 (N_6628,N_6125,N_6197);
nor U6629 (N_6629,N_6140,N_6317);
nor U6630 (N_6630,N_6244,N_6137);
nor U6631 (N_6631,N_6384,N_6234);
nand U6632 (N_6632,N_6180,N_6368);
and U6633 (N_6633,N_6254,N_6388);
xor U6634 (N_6634,N_6160,N_6398);
and U6635 (N_6635,N_6187,N_6335);
or U6636 (N_6636,N_6310,N_6007);
nor U6637 (N_6637,N_6014,N_6106);
xnor U6638 (N_6638,N_6262,N_6142);
and U6639 (N_6639,N_6286,N_6125);
or U6640 (N_6640,N_6094,N_6209);
xnor U6641 (N_6641,N_6070,N_6101);
nor U6642 (N_6642,N_6286,N_6037);
nor U6643 (N_6643,N_6216,N_6013);
or U6644 (N_6644,N_6121,N_6085);
nor U6645 (N_6645,N_6135,N_6057);
and U6646 (N_6646,N_6017,N_6115);
xor U6647 (N_6647,N_6219,N_6015);
xor U6648 (N_6648,N_6257,N_6388);
and U6649 (N_6649,N_6365,N_6078);
nand U6650 (N_6650,N_6126,N_6363);
xor U6651 (N_6651,N_6114,N_6232);
xnor U6652 (N_6652,N_6202,N_6098);
and U6653 (N_6653,N_6278,N_6093);
or U6654 (N_6654,N_6362,N_6174);
nand U6655 (N_6655,N_6125,N_6131);
or U6656 (N_6656,N_6103,N_6291);
xor U6657 (N_6657,N_6368,N_6378);
or U6658 (N_6658,N_6009,N_6284);
and U6659 (N_6659,N_6394,N_6276);
or U6660 (N_6660,N_6049,N_6050);
nor U6661 (N_6661,N_6270,N_6243);
and U6662 (N_6662,N_6385,N_6191);
xor U6663 (N_6663,N_6312,N_6290);
nor U6664 (N_6664,N_6027,N_6284);
nor U6665 (N_6665,N_6261,N_6229);
and U6666 (N_6666,N_6316,N_6162);
or U6667 (N_6667,N_6019,N_6008);
nand U6668 (N_6668,N_6094,N_6358);
nor U6669 (N_6669,N_6188,N_6230);
nor U6670 (N_6670,N_6111,N_6199);
xnor U6671 (N_6671,N_6196,N_6335);
and U6672 (N_6672,N_6394,N_6283);
or U6673 (N_6673,N_6246,N_6295);
nand U6674 (N_6674,N_6249,N_6123);
nand U6675 (N_6675,N_6169,N_6319);
or U6676 (N_6676,N_6184,N_6143);
nand U6677 (N_6677,N_6214,N_6343);
xnor U6678 (N_6678,N_6147,N_6367);
and U6679 (N_6679,N_6335,N_6347);
nor U6680 (N_6680,N_6388,N_6110);
and U6681 (N_6681,N_6293,N_6023);
nor U6682 (N_6682,N_6099,N_6398);
xor U6683 (N_6683,N_6153,N_6048);
or U6684 (N_6684,N_6205,N_6177);
nand U6685 (N_6685,N_6006,N_6176);
xor U6686 (N_6686,N_6236,N_6347);
xnor U6687 (N_6687,N_6171,N_6374);
xor U6688 (N_6688,N_6090,N_6010);
and U6689 (N_6689,N_6300,N_6195);
nand U6690 (N_6690,N_6142,N_6228);
nand U6691 (N_6691,N_6161,N_6088);
xor U6692 (N_6692,N_6084,N_6031);
xor U6693 (N_6693,N_6098,N_6087);
and U6694 (N_6694,N_6218,N_6164);
xor U6695 (N_6695,N_6229,N_6135);
nor U6696 (N_6696,N_6057,N_6201);
nor U6697 (N_6697,N_6356,N_6206);
nand U6698 (N_6698,N_6039,N_6179);
and U6699 (N_6699,N_6260,N_6235);
nand U6700 (N_6700,N_6311,N_6324);
and U6701 (N_6701,N_6374,N_6343);
nor U6702 (N_6702,N_6291,N_6060);
nor U6703 (N_6703,N_6327,N_6320);
nor U6704 (N_6704,N_6021,N_6282);
or U6705 (N_6705,N_6203,N_6353);
and U6706 (N_6706,N_6315,N_6269);
nand U6707 (N_6707,N_6163,N_6176);
nor U6708 (N_6708,N_6380,N_6109);
or U6709 (N_6709,N_6149,N_6223);
nand U6710 (N_6710,N_6154,N_6203);
and U6711 (N_6711,N_6056,N_6225);
or U6712 (N_6712,N_6255,N_6289);
or U6713 (N_6713,N_6218,N_6279);
xor U6714 (N_6714,N_6010,N_6065);
nand U6715 (N_6715,N_6075,N_6086);
xnor U6716 (N_6716,N_6306,N_6235);
and U6717 (N_6717,N_6156,N_6102);
and U6718 (N_6718,N_6210,N_6212);
and U6719 (N_6719,N_6121,N_6224);
or U6720 (N_6720,N_6121,N_6286);
nor U6721 (N_6721,N_6349,N_6015);
or U6722 (N_6722,N_6185,N_6104);
nor U6723 (N_6723,N_6271,N_6228);
nand U6724 (N_6724,N_6305,N_6110);
nor U6725 (N_6725,N_6183,N_6267);
nand U6726 (N_6726,N_6392,N_6090);
nor U6727 (N_6727,N_6008,N_6394);
and U6728 (N_6728,N_6002,N_6271);
or U6729 (N_6729,N_6051,N_6130);
nor U6730 (N_6730,N_6025,N_6018);
and U6731 (N_6731,N_6391,N_6009);
and U6732 (N_6732,N_6040,N_6049);
xnor U6733 (N_6733,N_6197,N_6002);
xnor U6734 (N_6734,N_6387,N_6166);
xnor U6735 (N_6735,N_6298,N_6136);
nor U6736 (N_6736,N_6267,N_6173);
nand U6737 (N_6737,N_6087,N_6232);
nor U6738 (N_6738,N_6010,N_6305);
or U6739 (N_6739,N_6091,N_6266);
xor U6740 (N_6740,N_6342,N_6286);
and U6741 (N_6741,N_6088,N_6054);
nor U6742 (N_6742,N_6200,N_6113);
xor U6743 (N_6743,N_6385,N_6131);
nor U6744 (N_6744,N_6329,N_6056);
and U6745 (N_6745,N_6245,N_6311);
nand U6746 (N_6746,N_6227,N_6159);
nand U6747 (N_6747,N_6341,N_6090);
xnor U6748 (N_6748,N_6040,N_6382);
xor U6749 (N_6749,N_6237,N_6147);
nor U6750 (N_6750,N_6013,N_6355);
and U6751 (N_6751,N_6261,N_6179);
nor U6752 (N_6752,N_6211,N_6353);
xor U6753 (N_6753,N_6087,N_6163);
nand U6754 (N_6754,N_6351,N_6249);
or U6755 (N_6755,N_6399,N_6253);
and U6756 (N_6756,N_6145,N_6327);
or U6757 (N_6757,N_6380,N_6012);
or U6758 (N_6758,N_6250,N_6335);
nor U6759 (N_6759,N_6105,N_6111);
nor U6760 (N_6760,N_6308,N_6158);
xor U6761 (N_6761,N_6184,N_6139);
nor U6762 (N_6762,N_6066,N_6141);
nand U6763 (N_6763,N_6341,N_6210);
nor U6764 (N_6764,N_6038,N_6315);
nand U6765 (N_6765,N_6197,N_6360);
nand U6766 (N_6766,N_6099,N_6359);
and U6767 (N_6767,N_6252,N_6391);
nand U6768 (N_6768,N_6074,N_6378);
nand U6769 (N_6769,N_6110,N_6063);
and U6770 (N_6770,N_6242,N_6380);
or U6771 (N_6771,N_6180,N_6127);
nor U6772 (N_6772,N_6279,N_6337);
and U6773 (N_6773,N_6162,N_6036);
or U6774 (N_6774,N_6192,N_6147);
and U6775 (N_6775,N_6329,N_6112);
nor U6776 (N_6776,N_6163,N_6302);
xnor U6777 (N_6777,N_6158,N_6260);
xnor U6778 (N_6778,N_6163,N_6001);
xnor U6779 (N_6779,N_6259,N_6373);
and U6780 (N_6780,N_6287,N_6215);
and U6781 (N_6781,N_6273,N_6126);
xnor U6782 (N_6782,N_6156,N_6390);
nor U6783 (N_6783,N_6059,N_6205);
nand U6784 (N_6784,N_6173,N_6119);
xnor U6785 (N_6785,N_6324,N_6353);
or U6786 (N_6786,N_6296,N_6221);
nor U6787 (N_6787,N_6169,N_6389);
nand U6788 (N_6788,N_6365,N_6250);
nand U6789 (N_6789,N_6122,N_6186);
nand U6790 (N_6790,N_6046,N_6294);
nor U6791 (N_6791,N_6035,N_6013);
nand U6792 (N_6792,N_6029,N_6098);
or U6793 (N_6793,N_6258,N_6025);
nor U6794 (N_6794,N_6188,N_6240);
nor U6795 (N_6795,N_6213,N_6051);
and U6796 (N_6796,N_6360,N_6257);
xnor U6797 (N_6797,N_6145,N_6334);
and U6798 (N_6798,N_6340,N_6339);
nand U6799 (N_6799,N_6162,N_6189);
or U6800 (N_6800,N_6585,N_6753);
and U6801 (N_6801,N_6519,N_6759);
or U6802 (N_6802,N_6506,N_6429);
and U6803 (N_6803,N_6775,N_6613);
nor U6804 (N_6804,N_6442,N_6448);
nand U6805 (N_6805,N_6450,N_6610);
nor U6806 (N_6806,N_6544,N_6594);
nand U6807 (N_6807,N_6618,N_6560);
nor U6808 (N_6808,N_6491,N_6572);
xnor U6809 (N_6809,N_6559,N_6466);
xor U6810 (N_6810,N_6454,N_6521);
or U6811 (N_6811,N_6583,N_6698);
and U6812 (N_6812,N_6561,N_6414);
nand U6813 (N_6813,N_6680,N_6716);
and U6814 (N_6814,N_6413,N_6638);
nand U6815 (N_6815,N_6453,N_6714);
or U6816 (N_6816,N_6776,N_6552);
xnor U6817 (N_6817,N_6432,N_6791);
nand U6818 (N_6818,N_6730,N_6732);
nor U6819 (N_6819,N_6734,N_6721);
and U6820 (N_6820,N_6640,N_6408);
or U6821 (N_6821,N_6459,N_6428);
or U6822 (N_6822,N_6611,N_6565);
nand U6823 (N_6823,N_6627,N_6783);
nor U6824 (N_6824,N_6757,N_6761);
or U6825 (N_6825,N_6515,N_6481);
nor U6826 (N_6826,N_6601,N_6449);
xnor U6827 (N_6827,N_6599,N_6503);
and U6828 (N_6828,N_6616,N_6542);
and U6829 (N_6829,N_6778,N_6670);
or U6830 (N_6830,N_6467,N_6743);
and U6831 (N_6831,N_6646,N_6703);
nand U6832 (N_6832,N_6742,N_6693);
xor U6833 (N_6833,N_6694,N_6705);
xor U6834 (N_6834,N_6751,N_6617);
xnor U6835 (N_6835,N_6674,N_6756);
and U6836 (N_6836,N_6592,N_6427);
and U6837 (N_6837,N_6451,N_6685);
or U6838 (N_6838,N_6792,N_6483);
nor U6839 (N_6839,N_6400,N_6660);
xor U6840 (N_6840,N_6486,N_6725);
and U6841 (N_6841,N_6666,N_6456);
and U6842 (N_6842,N_6538,N_6492);
nand U6843 (N_6843,N_6562,N_6747);
or U6844 (N_6844,N_6551,N_6582);
nor U6845 (N_6845,N_6619,N_6591);
and U6846 (N_6846,N_6508,N_6794);
or U6847 (N_6847,N_6425,N_6471);
or U6848 (N_6848,N_6423,N_6493);
xor U6849 (N_6849,N_6411,N_6487);
xor U6850 (N_6850,N_6779,N_6692);
nand U6851 (N_6851,N_6782,N_6419);
or U6852 (N_6852,N_6505,N_6550);
nor U6853 (N_6853,N_6718,N_6630);
xor U6854 (N_6854,N_6607,N_6696);
or U6855 (N_6855,N_6490,N_6580);
and U6856 (N_6856,N_6426,N_6679);
xor U6857 (N_6857,N_6785,N_6780);
xor U6858 (N_6858,N_6765,N_6665);
nand U6859 (N_6859,N_6633,N_6479);
nor U6860 (N_6860,N_6641,N_6590);
xnor U6861 (N_6861,N_6691,N_6689);
and U6862 (N_6862,N_6533,N_6474);
or U6863 (N_6863,N_6570,N_6539);
nand U6864 (N_6864,N_6628,N_6526);
nor U6865 (N_6865,N_6573,N_6702);
nand U6866 (N_6866,N_6612,N_6568);
nor U6867 (N_6867,N_6522,N_6536);
or U6868 (N_6868,N_6763,N_6738);
nand U6869 (N_6869,N_6784,N_6623);
or U6870 (N_6870,N_6494,N_6445);
nand U6871 (N_6871,N_6553,N_6748);
or U6872 (N_6872,N_6476,N_6754);
xor U6873 (N_6873,N_6710,N_6566);
xor U6874 (N_6874,N_6488,N_6571);
or U6875 (N_6875,N_6787,N_6403);
nor U6876 (N_6876,N_6407,N_6688);
nand U6877 (N_6877,N_6774,N_6600);
or U6878 (N_6878,N_6405,N_6699);
and U6879 (N_6879,N_6762,N_6657);
xor U6880 (N_6880,N_6659,N_6460);
nand U6881 (N_6881,N_6681,N_6537);
xnor U6882 (N_6882,N_6736,N_6713);
nor U6883 (N_6883,N_6579,N_6706);
and U6884 (N_6884,N_6437,N_6789);
nor U6885 (N_6885,N_6447,N_6667);
nand U6886 (N_6886,N_6418,N_6675);
nand U6887 (N_6887,N_6661,N_6457);
and U6888 (N_6888,N_6575,N_6722);
and U6889 (N_6889,N_6620,N_6412);
and U6890 (N_6890,N_6707,N_6768);
or U6891 (N_6891,N_6602,N_6655);
or U6892 (N_6892,N_6438,N_6529);
nand U6893 (N_6893,N_6523,N_6647);
nand U6894 (N_6894,N_6518,N_6712);
or U6895 (N_6895,N_6605,N_6656);
nor U6896 (N_6896,N_6576,N_6773);
and U6897 (N_6897,N_6643,N_6547);
xor U6898 (N_6898,N_6593,N_6540);
or U6899 (N_6899,N_6462,N_6777);
and U6900 (N_6900,N_6439,N_6767);
nand U6901 (N_6901,N_6682,N_6567);
and U6902 (N_6902,N_6589,N_6475);
and U6903 (N_6903,N_6744,N_6788);
or U6904 (N_6904,N_6501,N_6634);
xnor U6905 (N_6905,N_6598,N_6435);
and U6906 (N_6906,N_6420,N_6458);
nand U6907 (N_6907,N_6772,N_6662);
xnor U6908 (N_6908,N_6527,N_6709);
nor U6909 (N_6909,N_6422,N_6524);
and U6910 (N_6910,N_6671,N_6648);
xor U6911 (N_6911,N_6401,N_6549);
and U6912 (N_6912,N_6745,N_6650);
or U6913 (N_6913,N_6644,N_6786);
nor U6914 (N_6914,N_6433,N_6677);
nor U6915 (N_6915,N_6581,N_6797);
nor U6916 (N_6916,N_6584,N_6404);
or U6917 (N_6917,N_6497,N_6793);
nor U6918 (N_6918,N_6629,N_6781);
nor U6919 (N_6919,N_6444,N_6517);
nor U6920 (N_6920,N_6402,N_6525);
xnor U6921 (N_6921,N_6502,N_6556);
nand U6922 (N_6922,N_6637,N_6755);
nand U6923 (N_6923,N_6597,N_6764);
or U6924 (N_6924,N_6625,N_6749);
nor U6925 (N_6925,N_6690,N_6760);
nand U6926 (N_6926,N_6608,N_6520);
or U6927 (N_6927,N_6558,N_6727);
or U6928 (N_6928,N_6739,N_6541);
nand U6929 (N_6929,N_6511,N_6635);
nand U6930 (N_6930,N_6431,N_6498);
xnor U6931 (N_6931,N_6606,N_6489);
xnor U6932 (N_6932,N_6672,N_6455);
xor U6933 (N_6933,N_6771,N_6614);
and U6934 (N_6934,N_6711,N_6639);
or U6935 (N_6935,N_6726,N_6532);
nand U6936 (N_6936,N_6642,N_6704);
xnor U6937 (N_6937,N_6470,N_6545);
and U6938 (N_6938,N_6577,N_6441);
nand U6939 (N_6939,N_6557,N_6632);
nand U6940 (N_6940,N_6495,N_6622);
xnor U6941 (N_6941,N_6669,N_6430);
or U6942 (N_6942,N_6509,N_6609);
xor U6943 (N_6943,N_6443,N_6478);
and U6944 (N_6944,N_6741,N_6651);
or U6945 (N_6945,N_6687,N_6452);
xor U6946 (N_6946,N_6416,N_6735);
nand U6947 (N_6947,N_6469,N_6507);
or U6948 (N_6948,N_6464,N_6417);
or U6949 (N_6949,N_6615,N_6652);
xnor U6950 (N_6950,N_6697,N_6737);
xnor U6951 (N_6951,N_6758,N_6603);
or U6952 (N_6952,N_6484,N_6410);
nand U6953 (N_6953,N_6664,N_6700);
xnor U6954 (N_6954,N_6649,N_6578);
nand U6955 (N_6955,N_6468,N_6752);
xnor U6956 (N_6956,N_6676,N_6548);
nor U6957 (N_6957,N_6720,N_6708);
or U6958 (N_6958,N_6731,N_6683);
xnor U6959 (N_6959,N_6587,N_6485);
nor U6960 (N_6960,N_6686,N_6436);
or U6961 (N_6961,N_6626,N_6446);
and U6962 (N_6962,N_6555,N_6472);
xnor U6963 (N_6963,N_6719,N_6799);
xnor U6964 (N_6964,N_6463,N_6513);
or U6965 (N_6965,N_6596,N_6514);
and U6966 (N_6966,N_6473,N_6569);
xor U6967 (N_6967,N_6496,N_6554);
nor U6968 (N_6968,N_6563,N_6499);
nand U6969 (N_6969,N_6504,N_6770);
nor U6970 (N_6970,N_6415,N_6684);
nand U6971 (N_6971,N_6769,N_6724);
nor U6972 (N_6972,N_6740,N_6482);
nand U6973 (N_6973,N_6574,N_6636);
and U6974 (N_6974,N_6595,N_6645);
and U6975 (N_6975,N_6409,N_6658);
or U6976 (N_6976,N_6528,N_6477);
xor U6977 (N_6977,N_6564,N_6440);
or U6978 (N_6978,N_6424,N_6531);
nor U6979 (N_6979,N_6723,N_6543);
or U6980 (N_6980,N_6621,N_6701);
nand U6981 (N_6981,N_6535,N_6750);
nand U6982 (N_6982,N_6790,N_6461);
nor U6983 (N_6983,N_6480,N_6588);
xor U6984 (N_6984,N_6465,N_6766);
nand U6985 (N_6985,N_6668,N_6654);
nor U6986 (N_6986,N_6421,N_6733);
xor U6987 (N_6987,N_6631,N_6516);
nor U6988 (N_6988,N_6795,N_6530);
xor U6989 (N_6989,N_6729,N_6624);
xor U6990 (N_6990,N_6663,N_6796);
xnor U6991 (N_6991,N_6653,N_6717);
nand U6992 (N_6992,N_6798,N_6546);
nand U6993 (N_6993,N_6534,N_6604);
and U6994 (N_6994,N_6586,N_6728);
nor U6995 (N_6995,N_6500,N_6678);
xor U6996 (N_6996,N_6434,N_6746);
xor U6997 (N_6997,N_6715,N_6695);
xnor U6998 (N_6998,N_6673,N_6406);
or U6999 (N_6999,N_6512,N_6510);
or U7000 (N_7000,N_6552,N_6487);
and U7001 (N_7001,N_6749,N_6623);
nor U7002 (N_7002,N_6579,N_6593);
nor U7003 (N_7003,N_6662,N_6558);
nand U7004 (N_7004,N_6416,N_6587);
xnor U7005 (N_7005,N_6580,N_6501);
xnor U7006 (N_7006,N_6628,N_6589);
nor U7007 (N_7007,N_6453,N_6795);
or U7008 (N_7008,N_6711,N_6597);
or U7009 (N_7009,N_6709,N_6776);
and U7010 (N_7010,N_6741,N_6403);
nor U7011 (N_7011,N_6776,N_6745);
nor U7012 (N_7012,N_6665,N_6495);
nand U7013 (N_7013,N_6539,N_6636);
and U7014 (N_7014,N_6618,N_6698);
xor U7015 (N_7015,N_6698,N_6423);
nand U7016 (N_7016,N_6564,N_6622);
or U7017 (N_7017,N_6633,N_6651);
xnor U7018 (N_7018,N_6594,N_6704);
xor U7019 (N_7019,N_6698,N_6695);
nor U7020 (N_7020,N_6558,N_6781);
nor U7021 (N_7021,N_6774,N_6414);
nand U7022 (N_7022,N_6658,N_6530);
and U7023 (N_7023,N_6452,N_6657);
and U7024 (N_7024,N_6605,N_6633);
or U7025 (N_7025,N_6517,N_6552);
and U7026 (N_7026,N_6586,N_6776);
or U7027 (N_7027,N_6659,N_6517);
or U7028 (N_7028,N_6673,N_6548);
or U7029 (N_7029,N_6408,N_6619);
nand U7030 (N_7030,N_6447,N_6472);
or U7031 (N_7031,N_6616,N_6682);
nand U7032 (N_7032,N_6553,N_6719);
xor U7033 (N_7033,N_6612,N_6769);
xor U7034 (N_7034,N_6727,N_6511);
xnor U7035 (N_7035,N_6595,N_6694);
nand U7036 (N_7036,N_6776,N_6550);
xnor U7037 (N_7037,N_6656,N_6457);
and U7038 (N_7038,N_6452,N_6470);
nand U7039 (N_7039,N_6590,N_6670);
or U7040 (N_7040,N_6425,N_6467);
or U7041 (N_7041,N_6582,N_6570);
nand U7042 (N_7042,N_6599,N_6538);
or U7043 (N_7043,N_6644,N_6478);
nand U7044 (N_7044,N_6477,N_6670);
or U7045 (N_7045,N_6732,N_6705);
nand U7046 (N_7046,N_6542,N_6548);
xor U7047 (N_7047,N_6623,N_6693);
nand U7048 (N_7048,N_6796,N_6482);
nor U7049 (N_7049,N_6764,N_6600);
or U7050 (N_7050,N_6748,N_6402);
nand U7051 (N_7051,N_6413,N_6523);
or U7052 (N_7052,N_6671,N_6443);
or U7053 (N_7053,N_6683,N_6530);
nand U7054 (N_7054,N_6579,N_6679);
nand U7055 (N_7055,N_6779,N_6634);
nand U7056 (N_7056,N_6656,N_6422);
and U7057 (N_7057,N_6763,N_6709);
xor U7058 (N_7058,N_6774,N_6702);
nand U7059 (N_7059,N_6754,N_6634);
and U7060 (N_7060,N_6752,N_6695);
xor U7061 (N_7061,N_6633,N_6510);
or U7062 (N_7062,N_6450,N_6647);
and U7063 (N_7063,N_6746,N_6571);
xor U7064 (N_7064,N_6689,N_6541);
or U7065 (N_7065,N_6640,N_6715);
nand U7066 (N_7066,N_6721,N_6416);
xor U7067 (N_7067,N_6450,N_6605);
nor U7068 (N_7068,N_6556,N_6737);
nand U7069 (N_7069,N_6636,N_6560);
xor U7070 (N_7070,N_6785,N_6489);
nor U7071 (N_7071,N_6431,N_6512);
or U7072 (N_7072,N_6680,N_6496);
and U7073 (N_7073,N_6559,N_6734);
nand U7074 (N_7074,N_6597,N_6649);
xnor U7075 (N_7075,N_6628,N_6656);
or U7076 (N_7076,N_6509,N_6467);
xor U7077 (N_7077,N_6726,N_6721);
nand U7078 (N_7078,N_6605,N_6554);
or U7079 (N_7079,N_6590,N_6496);
xnor U7080 (N_7080,N_6623,N_6773);
or U7081 (N_7081,N_6425,N_6588);
or U7082 (N_7082,N_6480,N_6571);
or U7083 (N_7083,N_6521,N_6461);
xnor U7084 (N_7084,N_6555,N_6434);
xor U7085 (N_7085,N_6702,N_6534);
nand U7086 (N_7086,N_6759,N_6703);
nand U7087 (N_7087,N_6424,N_6485);
or U7088 (N_7088,N_6698,N_6647);
nor U7089 (N_7089,N_6496,N_6771);
nor U7090 (N_7090,N_6614,N_6480);
nor U7091 (N_7091,N_6428,N_6689);
or U7092 (N_7092,N_6665,N_6404);
or U7093 (N_7093,N_6753,N_6478);
and U7094 (N_7094,N_6592,N_6578);
and U7095 (N_7095,N_6782,N_6539);
nor U7096 (N_7096,N_6484,N_6723);
nand U7097 (N_7097,N_6567,N_6485);
nor U7098 (N_7098,N_6753,N_6744);
nand U7099 (N_7099,N_6675,N_6712);
nand U7100 (N_7100,N_6780,N_6529);
and U7101 (N_7101,N_6575,N_6558);
and U7102 (N_7102,N_6439,N_6403);
and U7103 (N_7103,N_6782,N_6664);
xnor U7104 (N_7104,N_6451,N_6583);
xnor U7105 (N_7105,N_6720,N_6479);
and U7106 (N_7106,N_6657,N_6741);
and U7107 (N_7107,N_6486,N_6773);
xnor U7108 (N_7108,N_6787,N_6456);
and U7109 (N_7109,N_6731,N_6503);
nor U7110 (N_7110,N_6714,N_6708);
or U7111 (N_7111,N_6473,N_6602);
nor U7112 (N_7112,N_6494,N_6730);
and U7113 (N_7113,N_6596,N_6685);
nand U7114 (N_7114,N_6618,N_6515);
nor U7115 (N_7115,N_6545,N_6506);
nor U7116 (N_7116,N_6742,N_6677);
nor U7117 (N_7117,N_6408,N_6502);
or U7118 (N_7118,N_6757,N_6427);
nand U7119 (N_7119,N_6622,N_6714);
nand U7120 (N_7120,N_6634,N_6588);
nand U7121 (N_7121,N_6523,N_6782);
and U7122 (N_7122,N_6638,N_6502);
nand U7123 (N_7123,N_6487,N_6526);
or U7124 (N_7124,N_6634,N_6740);
xor U7125 (N_7125,N_6611,N_6771);
or U7126 (N_7126,N_6685,N_6588);
nor U7127 (N_7127,N_6683,N_6596);
and U7128 (N_7128,N_6676,N_6689);
and U7129 (N_7129,N_6544,N_6782);
nand U7130 (N_7130,N_6540,N_6722);
or U7131 (N_7131,N_6534,N_6643);
xnor U7132 (N_7132,N_6621,N_6608);
and U7133 (N_7133,N_6765,N_6431);
nand U7134 (N_7134,N_6410,N_6482);
nor U7135 (N_7135,N_6537,N_6668);
or U7136 (N_7136,N_6588,N_6608);
xnor U7137 (N_7137,N_6497,N_6670);
nor U7138 (N_7138,N_6468,N_6750);
xnor U7139 (N_7139,N_6400,N_6745);
nand U7140 (N_7140,N_6705,N_6539);
or U7141 (N_7141,N_6512,N_6715);
xor U7142 (N_7142,N_6455,N_6444);
and U7143 (N_7143,N_6478,N_6560);
nand U7144 (N_7144,N_6544,N_6442);
and U7145 (N_7145,N_6639,N_6637);
or U7146 (N_7146,N_6734,N_6477);
or U7147 (N_7147,N_6609,N_6641);
xnor U7148 (N_7148,N_6715,N_6444);
nor U7149 (N_7149,N_6709,N_6732);
and U7150 (N_7150,N_6406,N_6640);
or U7151 (N_7151,N_6433,N_6406);
nand U7152 (N_7152,N_6477,N_6414);
nand U7153 (N_7153,N_6680,N_6598);
or U7154 (N_7154,N_6522,N_6430);
nand U7155 (N_7155,N_6445,N_6487);
and U7156 (N_7156,N_6542,N_6714);
nor U7157 (N_7157,N_6740,N_6596);
xor U7158 (N_7158,N_6552,N_6573);
nand U7159 (N_7159,N_6590,N_6616);
xnor U7160 (N_7160,N_6751,N_6742);
nor U7161 (N_7161,N_6552,N_6472);
or U7162 (N_7162,N_6606,N_6568);
and U7163 (N_7163,N_6556,N_6520);
and U7164 (N_7164,N_6602,N_6618);
and U7165 (N_7165,N_6606,N_6661);
nor U7166 (N_7166,N_6408,N_6717);
or U7167 (N_7167,N_6668,N_6566);
xor U7168 (N_7168,N_6664,N_6720);
nand U7169 (N_7169,N_6574,N_6644);
nand U7170 (N_7170,N_6516,N_6680);
or U7171 (N_7171,N_6497,N_6458);
xnor U7172 (N_7172,N_6593,N_6558);
and U7173 (N_7173,N_6789,N_6662);
nand U7174 (N_7174,N_6724,N_6605);
nor U7175 (N_7175,N_6664,N_6441);
nor U7176 (N_7176,N_6492,N_6673);
and U7177 (N_7177,N_6775,N_6728);
nor U7178 (N_7178,N_6699,N_6707);
nand U7179 (N_7179,N_6700,N_6459);
xor U7180 (N_7180,N_6458,N_6671);
nand U7181 (N_7181,N_6596,N_6592);
nand U7182 (N_7182,N_6687,N_6659);
nand U7183 (N_7183,N_6572,N_6497);
or U7184 (N_7184,N_6751,N_6629);
nand U7185 (N_7185,N_6687,N_6515);
xnor U7186 (N_7186,N_6755,N_6498);
nor U7187 (N_7187,N_6647,N_6611);
or U7188 (N_7188,N_6514,N_6701);
or U7189 (N_7189,N_6642,N_6788);
or U7190 (N_7190,N_6650,N_6401);
or U7191 (N_7191,N_6486,N_6413);
xor U7192 (N_7192,N_6437,N_6486);
nand U7193 (N_7193,N_6550,N_6466);
nand U7194 (N_7194,N_6599,N_6438);
nor U7195 (N_7195,N_6748,N_6761);
xnor U7196 (N_7196,N_6574,N_6678);
nand U7197 (N_7197,N_6608,N_6718);
xor U7198 (N_7198,N_6731,N_6696);
or U7199 (N_7199,N_6662,N_6709);
and U7200 (N_7200,N_6914,N_7110);
nand U7201 (N_7201,N_7177,N_6867);
or U7202 (N_7202,N_6985,N_7064);
nor U7203 (N_7203,N_7100,N_7098);
xor U7204 (N_7204,N_7010,N_6965);
and U7205 (N_7205,N_7070,N_7092);
nand U7206 (N_7206,N_6843,N_6846);
nand U7207 (N_7207,N_7157,N_6803);
or U7208 (N_7208,N_7020,N_7050);
and U7209 (N_7209,N_6928,N_6980);
nor U7210 (N_7210,N_6921,N_7093);
or U7211 (N_7211,N_6924,N_7037);
or U7212 (N_7212,N_7193,N_7131);
or U7213 (N_7213,N_6934,N_7172);
nor U7214 (N_7214,N_7097,N_6839);
nand U7215 (N_7215,N_7057,N_6970);
nor U7216 (N_7216,N_6809,N_6981);
and U7217 (N_7217,N_6957,N_7164);
or U7218 (N_7218,N_6858,N_6910);
or U7219 (N_7219,N_6818,N_7062);
xnor U7220 (N_7220,N_7156,N_7073);
nand U7221 (N_7221,N_6911,N_6856);
or U7222 (N_7222,N_7174,N_6979);
nor U7223 (N_7223,N_6898,N_6935);
nand U7224 (N_7224,N_7138,N_7155);
nand U7225 (N_7225,N_6896,N_7132);
nand U7226 (N_7226,N_7011,N_6923);
and U7227 (N_7227,N_6807,N_6829);
xor U7228 (N_7228,N_6817,N_7001);
or U7229 (N_7229,N_7152,N_7078);
xor U7230 (N_7230,N_6802,N_6853);
nand U7231 (N_7231,N_7016,N_7086);
or U7232 (N_7232,N_7195,N_7180);
nand U7233 (N_7233,N_7075,N_6948);
nor U7234 (N_7234,N_6949,N_7129);
nor U7235 (N_7235,N_6943,N_7041);
and U7236 (N_7236,N_7066,N_6902);
xor U7237 (N_7237,N_7042,N_6929);
and U7238 (N_7238,N_7069,N_7063);
or U7239 (N_7239,N_7154,N_6922);
nand U7240 (N_7240,N_6915,N_7052);
nor U7241 (N_7241,N_7178,N_7198);
xor U7242 (N_7242,N_6897,N_6954);
nand U7243 (N_7243,N_6958,N_7072);
and U7244 (N_7244,N_6968,N_6894);
nor U7245 (N_7245,N_7149,N_7146);
or U7246 (N_7246,N_7007,N_7049);
nor U7247 (N_7247,N_6890,N_6827);
or U7248 (N_7248,N_7189,N_6871);
nor U7249 (N_7249,N_6959,N_6999);
xor U7250 (N_7250,N_6953,N_7036);
xor U7251 (N_7251,N_7060,N_7048);
or U7252 (N_7252,N_7141,N_6878);
nor U7253 (N_7253,N_7142,N_6847);
xor U7254 (N_7254,N_7071,N_7067);
or U7255 (N_7255,N_6904,N_6821);
xor U7256 (N_7256,N_6886,N_7168);
nand U7257 (N_7257,N_6966,N_7051);
nand U7258 (N_7258,N_6905,N_7128);
and U7259 (N_7259,N_7160,N_7044);
nor U7260 (N_7260,N_6945,N_7140);
nand U7261 (N_7261,N_7014,N_7182);
nor U7262 (N_7262,N_7169,N_7135);
or U7263 (N_7263,N_6815,N_6909);
xor U7264 (N_7264,N_6833,N_6864);
xor U7265 (N_7265,N_7088,N_7103);
nand U7266 (N_7266,N_6991,N_7034);
or U7267 (N_7267,N_7023,N_6814);
xor U7268 (N_7268,N_6998,N_7126);
xnor U7269 (N_7269,N_6801,N_7122);
xnor U7270 (N_7270,N_6811,N_6800);
or U7271 (N_7271,N_6891,N_6819);
nand U7272 (N_7272,N_7065,N_7000);
nand U7273 (N_7273,N_6952,N_6820);
xnor U7274 (N_7274,N_6873,N_6836);
or U7275 (N_7275,N_7003,N_7083);
nand U7276 (N_7276,N_7095,N_7194);
nand U7277 (N_7277,N_6863,N_6955);
nand U7278 (N_7278,N_7018,N_6916);
xnor U7279 (N_7279,N_7107,N_6956);
and U7280 (N_7280,N_6984,N_6848);
or U7281 (N_7281,N_6812,N_6927);
nor U7282 (N_7282,N_7101,N_6813);
or U7283 (N_7283,N_6969,N_6860);
or U7284 (N_7284,N_6900,N_6993);
nor U7285 (N_7285,N_6912,N_6887);
or U7286 (N_7286,N_7061,N_7127);
or U7287 (N_7287,N_6964,N_6854);
or U7288 (N_7288,N_7039,N_7183);
or U7289 (N_7289,N_7190,N_7163);
xnor U7290 (N_7290,N_7115,N_6908);
or U7291 (N_7291,N_6889,N_7105);
xnor U7292 (N_7292,N_6825,N_7046);
xnor U7293 (N_7293,N_6987,N_7119);
xnor U7294 (N_7294,N_7108,N_6868);
nand U7295 (N_7295,N_7096,N_7024);
and U7296 (N_7296,N_7147,N_6805);
nand U7297 (N_7297,N_7068,N_7118);
xor U7298 (N_7298,N_6977,N_7079);
xnor U7299 (N_7299,N_7045,N_6884);
and U7300 (N_7300,N_7197,N_7043);
xnor U7301 (N_7301,N_6851,N_6972);
or U7302 (N_7302,N_6947,N_7084);
nand U7303 (N_7303,N_6808,N_7123);
and U7304 (N_7304,N_7176,N_6961);
and U7305 (N_7305,N_6982,N_6804);
or U7306 (N_7306,N_6840,N_6903);
and U7307 (N_7307,N_6842,N_6946);
or U7308 (N_7308,N_6880,N_6992);
or U7309 (N_7309,N_6828,N_6879);
xnor U7310 (N_7310,N_6931,N_6940);
nor U7311 (N_7311,N_7109,N_6865);
xnor U7312 (N_7312,N_7112,N_6845);
xor U7313 (N_7313,N_6855,N_7009);
and U7314 (N_7314,N_7179,N_7031);
and U7315 (N_7315,N_6932,N_7139);
xor U7316 (N_7316,N_6837,N_7058);
or U7317 (N_7317,N_6939,N_6831);
nor U7318 (N_7318,N_7148,N_7161);
and U7319 (N_7319,N_7120,N_6967);
or U7320 (N_7320,N_7038,N_6876);
and U7321 (N_7321,N_6883,N_7099);
or U7322 (N_7322,N_7087,N_6849);
or U7323 (N_7323,N_7158,N_6899);
and U7324 (N_7324,N_7167,N_7106);
nor U7325 (N_7325,N_7114,N_7192);
and U7326 (N_7326,N_6926,N_7030);
nand U7327 (N_7327,N_6941,N_7005);
or U7328 (N_7328,N_6816,N_7173);
nor U7329 (N_7329,N_7027,N_7165);
xor U7330 (N_7330,N_7006,N_6838);
and U7331 (N_7331,N_7134,N_7035);
or U7332 (N_7332,N_6901,N_7002);
or U7333 (N_7333,N_7013,N_7028);
nor U7334 (N_7334,N_7191,N_6933);
nor U7335 (N_7335,N_7125,N_7186);
or U7336 (N_7336,N_6974,N_6989);
nand U7337 (N_7337,N_6823,N_6906);
or U7338 (N_7338,N_7032,N_6937);
xor U7339 (N_7339,N_7159,N_7175);
and U7340 (N_7340,N_6841,N_6810);
nor U7341 (N_7341,N_6874,N_6983);
or U7342 (N_7342,N_6996,N_6895);
nand U7343 (N_7343,N_7077,N_6936);
nor U7344 (N_7344,N_7150,N_6888);
xor U7345 (N_7345,N_6866,N_6962);
xnor U7346 (N_7346,N_6885,N_6986);
xor U7347 (N_7347,N_7082,N_7196);
xor U7348 (N_7348,N_6881,N_7187);
nand U7349 (N_7349,N_6869,N_7145);
or U7350 (N_7350,N_6844,N_7137);
or U7351 (N_7351,N_6951,N_6973);
nor U7352 (N_7352,N_6882,N_6995);
and U7353 (N_7353,N_7124,N_7017);
xor U7354 (N_7354,N_6832,N_6861);
or U7355 (N_7355,N_7091,N_6872);
nand U7356 (N_7356,N_7130,N_7059);
nand U7357 (N_7357,N_6997,N_6990);
nand U7358 (N_7358,N_6930,N_6892);
nand U7359 (N_7359,N_7054,N_7022);
xnor U7360 (N_7360,N_6875,N_6822);
or U7361 (N_7361,N_7021,N_7166);
nand U7362 (N_7362,N_6942,N_7121);
or U7363 (N_7363,N_7144,N_7199);
and U7364 (N_7364,N_7089,N_7184);
or U7365 (N_7365,N_7055,N_7004);
nand U7366 (N_7366,N_7076,N_6920);
nand U7367 (N_7367,N_6830,N_7019);
xnor U7368 (N_7368,N_7029,N_7080);
nor U7369 (N_7369,N_6988,N_6852);
and U7370 (N_7370,N_6960,N_6913);
and U7371 (N_7371,N_6944,N_7026);
and U7372 (N_7372,N_7074,N_7033);
and U7373 (N_7373,N_6938,N_7185);
nand U7374 (N_7374,N_6978,N_7085);
nand U7375 (N_7375,N_6862,N_6963);
and U7376 (N_7376,N_6826,N_6859);
or U7377 (N_7377,N_7053,N_7151);
xor U7378 (N_7378,N_7181,N_7188);
nor U7379 (N_7379,N_6918,N_6950);
nand U7380 (N_7380,N_6806,N_6824);
nand U7381 (N_7381,N_6834,N_7047);
or U7382 (N_7382,N_6850,N_6857);
xor U7383 (N_7383,N_6994,N_6919);
and U7384 (N_7384,N_7117,N_6975);
and U7385 (N_7385,N_7090,N_7133);
xor U7386 (N_7386,N_7012,N_7170);
or U7387 (N_7387,N_7116,N_7015);
or U7388 (N_7388,N_7056,N_7143);
nor U7389 (N_7389,N_6870,N_7111);
or U7390 (N_7390,N_7008,N_7102);
and U7391 (N_7391,N_6971,N_7094);
nand U7392 (N_7392,N_7162,N_7113);
xor U7393 (N_7393,N_7081,N_6976);
xor U7394 (N_7394,N_7040,N_7025);
nand U7395 (N_7395,N_7171,N_7153);
nor U7396 (N_7396,N_6835,N_6877);
nand U7397 (N_7397,N_6907,N_6917);
nor U7398 (N_7398,N_6893,N_6925);
nand U7399 (N_7399,N_7104,N_7136);
and U7400 (N_7400,N_6861,N_6875);
xnor U7401 (N_7401,N_7151,N_7083);
xor U7402 (N_7402,N_6908,N_6911);
xnor U7403 (N_7403,N_6908,N_7029);
nand U7404 (N_7404,N_6938,N_7055);
xor U7405 (N_7405,N_6866,N_6830);
xnor U7406 (N_7406,N_6985,N_7070);
and U7407 (N_7407,N_6868,N_7070);
xor U7408 (N_7408,N_7190,N_7142);
or U7409 (N_7409,N_6850,N_7080);
xor U7410 (N_7410,N_7048,N_7112);
and U7411 (N_7411,N_6908,N_6824);
nor U7412 (N_7412,N_7124,N_7090);
xnor U7413 (N_7413,N_6983,N_7094);
or U7414 (N_7414,N_6967,N_7007);
or U7415 (N_7415,N_7166,N_7124);
and U7416 (N_7416,N_6857,N_7063);
xnor U7417 (N_7417,N_7131,N_7187);
or U7418 (N_7418,N_6935,N_7126);
xor U7419 (N_7419,N_7109,N_6837);
xnor U7420 (N_7420,N_6958,N_7127);
xnor U7421 (N_7421,N_7015,N_7012);
or U7422 (N_7422,N_6929,N_6994);
xnor U7423 (N_7423,N_6933,N_6943);
or U7424 (N_7424,N_6939,N_7110);
xnor U7425 (N_7425,N_6860,N_6885);
nor U7426 (N_7426,N_7122,N_6874);
nor U7427 (N_7427,N_7115,N_7114);
and U7428 (N_7428,N_7075,N_6925);
and U7429 (N_7429,N_7192,N_7103);
nand U7430 (N_7430,N_7143,N_7000);
or U7431 (N_7431,N_7140,N_6901);
or U7432 (N_7432,N_6808,N_7196);
and U7433 (N_7433,N_6929,N_6836);
xnor U7434 (N_7434,N_7123,N_6970);
and U7435 (N_7435,N_6843,N_7104);
xor U7436 (N_7436,N_6997,N_7131);
or U7437 (N_7437,N_7040,N_6840);
nor U7438 (N_7438,N_7129,N_6964);
or U7439 (N_7439,N_6968,N_6993);
nand U7440 (N_7440,N_6922,N_6874);
or U7441 (N_7441,N_7177,N_6948);
xnor U7442 (N_7442,N_7033,N_6979);
xnor U7443 (N_7443,N_6930,N_7068);
nor U7444 (N_7444,N_7137,N_7002);
nor U7445 (N_7445,N_7092,N_7018);
or U7446 (N_7446,N_6954,N_7134);
or U7447 (N_7447,N_6842,N_7080);
nor U7448 (N_7448,N_6869,N_6918);
nor U7449 (N_7449,N_6968,N_7194);
and U7450 (N_7450,N_6953,N_7055);
nor U7451 (N_7451,N_7051,N_7055);
and U7452 (N_7452,N_7043,N_6813);
nor U7453 (N_7453,N_6992,N_7089);
xnor U7454 (N_7454,N_6896,N_6991);
xnor U7455 (N_7455,N_6940,N_6978);
xor U7456 (N_7456,N_6986,N_7173);
or U7457 (N_7457,N_7139,N_7186);
and U7458 (N_7458,N_7067,N_6988);
and U7459 (N_7459,N_6853,N_6953);
or U7460 (N_7460,N_7126,N_7019);
or U7461 (N_7461,N_7132,N_7030);
xor U7462 (N_7462,N_7136,N_6873);
nand U7463 (N_7463,N_6832,N_6988);
or U7464 (N_7464,N_7160,N_7127);
xnor U7465 (N_7465,N_7052,N_7106);
nor U7466 (N_7466,N_7112,N_7186);
and U7467 (N_7467,N_6954,N_6909);
and U7468 (N_7468,N_7148,N_7024);
xor U7469 (N_7469,N_7191,N_6879);
and U7470 (N_7470,N_6882,N_7131);
and U7471 (N_7471,N_6918,N_6879);
or U7472 (N_7472,N_6814,N_6969);
and U7473 (N_7473,N_6902,N_7158);
and U7474 (N_7474,N_6815,N_7095);
nand U7475 (N_7475,N_7173,N_6859);
xnor U7476 (N_7476,N_7186,N_6804);
nor U7477 (N_7477,N_7113,N_7024);
or U7478 (N_7478,N_7156,N_6918);
nor U7479 (N_7479,N_7080,N_6920);
or U7480 (N_7480,N_7073,N_6855);
xor U7481 (N_7481,N_6929,N_7069);
and U7482 (N_7482,N_6976,N_7106);
or U7483 (N_7483,N_7146,N_6843);
nor U7484 (N_7484,N_6985,N_7079);
or U7485 (N_7485,N_7033,N_6808);
or U7486 (N_7486,N_6919,N_7025);
or U7487 (N_7487,N_6933,N_7156);
or U7488 (N_7488,N_6838,N_7108);
or U7489 (N_7489,N_6931,N_7176);
or U7490 (N_7490,N_7053,N_6973);
nand U7491 (N_7491,N_7190,N_6868);
or U7492 (N_7492,N_6869,N_6908);
nor U7493 (N_7493,N_7015,N_6909);
and U7494 (N_7494,N_6927,N_7112);
nand U7495 (N_7495,N_7114,N_6852);
nor U7496 (N_7496,N_6885,N_7057);
or U7497 (N_7497,N_7110,N_7109);
nor U7498 (N_7498,N_6848,N_7101);
xor U7499 (N_7499,N_6965,N_7022);
nor U7500 (N_7500,N_6820,N_7139);
nor U7501 (N_7501,N_6892,N_6885);
nor U7502 (N_7502,N_7166,N_7070);
nor U7503 (N_7503,N_6842,N_7001);
nor U7504 (N_7504,N_6869,N_7014);
nor U7505 (N_7505,N_7072,N_6874);
and U7506 (N_7506,N_7064,N_7170);
nand U7507 (N_7507,N_6900,N_6924);
nand U7508 (N_7508,N_7090,N_6925);
nand U7509 (N_7509,N_7163,N_7009);
nor U7510 (N_7510,N_6880,N_6825);
and U7511 (N_7511,N_7058,N_7016);
and U7512 (N_7512,N_6835,N_7173);
xnor U7513 (N_7513,N_7074,N_6804);
or U7514 (N_7514,N_6967,N_7180);
nor U7515 (N_7515,N_6922,N_6961);
and U7516 (N_7516,N_7115,N_6976);
xnor U7517 (N_7517,N_7168,N_7185);
nor U7518 (N_7518,N_6874,N_6877);
nand U7519 (N_7519,N_6958,N_7007);
nor U7520 (N_7520,N_6814,N_6971);
nor U7521 (N_7521,N_6889,N_6868);
nand U7522 (N_7522,N_7119,N_7170);
xnor U7523 (N_7523,N_7081,N_6933);
nor U7524 (N_7524,N_7033,N_7076);
or U7525 (N_7525,N_7161,N_7133);
and U7526 (N_7526,N_6845,N_6895);
or U7527 (N_7527,N_7062,N_7112);
nand U7528 (N_7528,N_6876,N_6810);
xor U7529 (N_7529,N_7015,N_6808);
and U7530 (N_7530,N_6922,N_7074);
and U7531 (N_7531,N_7146,N_7031);
or U7532 (N_7532,N_6825,N_6953);
or U7533 (N_7533,N_7051,N_6900);
nand U7534 (N_7534,N_7199,N_7096);
nor U7535 (N_7535,N_7057,N_7071);
xnor U7536 (N_7536,N_6935,N_7138);
xnor U7537 (N_7537,N_6813,N_6986);
or U7538 (N_7538,N_6920,N_7153);
or U7539 (N_7539,N_7193,N_6868);
or U7540 (N_7540,N_6965,N_6840);
xnor U7541 (N_7541,N_6893,N_6914);
and U7542 (N_7542,N_6977,N_6892);
and U7543 (N_7543,N_7112,N_7108);
nor U7544 (N_7544,N_7143,N_6970);
and U7545 (N_7545,N_6854,N_6885);
and U7546 (N_7546,N_6920,N_7114);
nand U7547 (N_7547,N_7093,N_6977);
nand U7548 (N_7548,N_7062,N_7131);
nand U7549 (N_7549,N_7041,N_7101);
or U7550 (N_7550,N_7077,N_7089);
xor U7551 (N_7551,N_7000,N_6907);
nor U7552 (N_7552,N_7130,N_6872);
nor U7553 (N_7553,N_7042,N_7097);
nand U7554 (N_7554,N_6930,N_7053);
nor U7555 (N_7555,N_7071,N_6925);
or U7556 (N_7556,N_7169,N_7151);
xnor U7557 (N_7557,N_6912,N_6935);
xnor U7558 (N_7558,N_6963,N_6802);
and U7559 (N_7559,N_6982,N_6999);
xnor U7560 (N_7560,N_7089,N_6955);
and U7561 (N_7561,N_6891,N_7006);
nand U7562 (N_7562,N_6903,N_6895);
nor U7563 (N_7563,N_6889,N_6867);
or U7564 (N_7564,N_6855,N_6895);
and U7565 (N_7565,N_6993,N_6938);
nor U7566 (N_7566,N_6990,N_7034);
and U7567 (N_7567,N_7006,N_7015);
nand U7568 (N_7568,N_6969,N_6851);
or U7569 (N_7569,N_6826,N_6820);
or U7570 (N_7570,N_6955,N_7115);
xor U7571 (N_7571,N_6957,N_6974);
nor U7572 (N_7572,N_7132,N_6880);
nand U7573 (N_7573,N_6841,N_6885);
nor U7574 (N_7574,N_6999,N_7089);
nand U7575 (N_7575,N_6894,N_7107);
xor U7576 (N_7576,N_7058,N_7007);
nor U7577 (N_7577,N_6986,N_6945);
nand U7578 (N_7578,N_6908,N_6885);
xor U7579 (N_7579,N_6969,N_6884);
xor U7580 (N_7580,N_6819,N_6953);
nor U7581 (N_7581,N_7030,N_6959);
and U7582 (N_7582,N_6846,N_6991);
nor U7583 (N_7583,N_6988,N_6965);
nand U7584 (N_7584,N_7054,N_6988);
nand U7585 (N_7585,N_6929,N_7012);
nor U7586 (N_7586,N_7126,N_7151);
nand U7587 (N_7587,N_7106,N_7195);
xnor U7588 (N_7588,N_7109,N_6957);
nand U7589 (N_7589,N_7010,N_6913);
or U7590 (N_7590,N_6958,N_7145);
xnor U7591 (N_7591,N_7155,N_7146);
and U7592 (N_7592,N_7175,N_6872);
xor U7593 (N_7593,N_7064,N_7172);
nand U7594 (N_7594,N_7021,N_6925);
xor U7595 (N_7595,N_7020,N_6811);
nor U7596 (N_7596,N_6823,N_7020);
or U7597 (N_7597,N_6876,N_7029);
xnor U7598 (N_7598,N_7129,N_6808);
nand U7599 (N_7599,N_7156,N_7142);
nor U7600 (N_7600,N_7517,N_7444);
nor U7601 (N_7601,N_7202,N_7293);
nand U7602 (N_7602,N_7290,N_7214);
or U7603 (N_7603,N_7432,N_7337);
nor U7604 (N_7604,N_7429,N_7329);
or U7605 (N_7605,N_7286,N_7566);
nand U7606 (N_7606,N_7474,N_7418);
and U7607 (N_7607,N_7538,N_7531);
nand U7608 (N_7608,N_7525,N_7553);
nand U7609 (N_7609,N_7225,N_7328);
and U7610 (N_7610,N_7381,N_7257);
nor U7611 (N_7611,N_7233,N_7508);
nor U7612 (N_7612,N_7269,N_7273);
nand U7613 (N_7613,N_7407,N_7483);
or U7614 (N_7614,N_7465,N_7281);
xor U7615 (N_7615,N_7468,N_7402);
xor U7616 (N_7616,N_7527,N_7392);
and U7617 (N_7617,N_7368,N_7502);
xnor U7618 (N_7618,N_7327,N_7320);
xnor U7619 (N_7619,N_7416,N_7279);
or U7620 (N_7620,N_7488,N_7388);
nor U7621 (N_7621,N_7394,N_7341);
xor U7622 (N_7622,N_7261,N_7475);
nand U7623 (N_7623,N_7270,N_7535);
or U7624 (N_7624,N_7252,N_7499);
or U7625 (N_7625,N_7289,N_7319);
and U7626 (N_7626,N_7536,N_7588);
or U7627 (N_7627,N_7403,N_7280);
nor U7628 (N_7628,N_7310,N_7396);
and U7629 (N_7629,N_7331,N_7294);
or U7630 (N_7630,N_7464,N_7491);
xor U7631 (N_7631,N_7345,N_7303);
nand U7632 (N_7632,N_7370,N_7282);
and U7633 (N_7633,N_7229,N_7543);
and U7634 (N_7634,N_7262,N_7456);
nand U7635 (N_7635,N_7428,N_7382);
xor U7636 (N_7636,N_7323,N_7458);
and U7637 (N_7637,N_7355,N_7467);
and U7638 (N_7638,N_7235,N_7462);
and U7639 (N_7639,N_7539,N_7529);
or U7640 (N_7640,N_7561,N_7398);
xor U7641 (N_7641,N_7453,N_7524);
and U7642 (N_7642,N_7550,N_7583);
nor U7643 (N_7643,N_7332,N_7520);
nor U7644 (N_7644,N_7503,N_7260);
or U7645 (N_7645,N_7569,N_7457);
nor U7646 (N_7646,N_7292,N_7477);
nand U7647 (N_7647,N_7478,N_7343);
xnor U7648 (N_7648,N_7299,N_7463);
and U7649 (N_7649,N_7454,N_7251);
or U7650 (N_7650,N_7203,N_7208);
and U7651 (N_7651,N_7514,N_7565);
nand U7652 (N_7652,N_7371,N_7461);
and U7653 (N_7653,N_7540,N_7264);
xor U7654 (N_7654,N_7222,N_7228);
nand U7655 (N_7655,N_7515,N_7486);
nand U7656 (N_7656,N_7442,N_7451);
xor U7657 (N_7657,N_7534,N_7557);
xnor U7658 (N_7658,N_7334,N_7239);
nand U7659 (N_7659,N_7356,N_7435);
and U7660 (N_7660,N_7369,N_7563);
or U7661 (N_7661,N_7276,N_7597);
or U7662 (N_7662,N_7577,N_7439);
and U7663 (N_7663,N_7568,N_7227);
nand U7664 (N_7664,N_7390,N_7379);
or U7665 (N_7665,N_7263,N_7243);
xor U7666 (N_7666,N_7570,N_7365);
nor U7667 (N_7667,N_7300,N_7436);
and U7668 (N_7668,N_7242,N_7206);
or U7669 (N_7669,N_7385,N_7267);
nand U7670 (N_7670,N_7250,N_7448);
and U7671 (N_7671,N_7336,N_7359);
or U7672 (N_7672,N_7406,N_7315);
xor U7673 (N_7673,N_7507,N_7265);
nand U7674 (N_7674,N_7528,N_7349);
or U7675 (N_7675,N_7441,N_7312);
and U7676 (N_7676,N_7395,N_7322);
and U7677 (N_7677,N_7351,N_7555);
nand U7678 (N_7678,N_7301,N_7344);
and U7679 (N_7679,N_7339,N_7594);
and U7680 (N_7680,N_7363,N_7479);
and U7681 (N_7681,N_7296,N_7326);
and U7682 (N_7682,N_7496,N_7450);
or U7683 (N_7683,N_7291,N_7231);
xnor U7684 (N_7684,N_7221,N_7505);
nand U7685 (N_7685,N_7518,N_7586);
and U7686 (N_7686,N_7576,N_7284);
nand U7687 (N_7687,N_7596,N_7526);
nor U7688 (N_7688,N_7558,N_7372);
nor U7689 (N_7689,N_7399,N_7590);
or U7690 (N_7690,N_7354,N_7510);
or U7691 (N_7691,N_7480,N_7512);
xor U7692 (N_7692,N_7424,N_7580);
nor U7693 (N_7693,N_7218,N_7256);
nor U7694 (N_7694,N_7469,N_7217);
and U7695 (N_7695,N_7414,N_7546);
nor U7696 (N_7696,N_7367,N_7574);
nand U7697 (N_7697,N_7492,N_7210);
xor U7698 (N_7698,N_7366,N_7241);
nand U7699 (N_7699,N_7500,N_7521);
xor U7700 (N_7700,N_7413,N_7380);
nand U7701 (N_7701,N_7274,N_7417);
and U7702 (N_7702,N_7575,N_7579);
nor U7703 (N_7703,N_7295,N_7446);
or U7704 (N_7704,N_7405,N_7230);
nor U7705 (N_7705,N_7277,N_7308);
xor U7706 (N_7706,N_7266,N_7223);
and U7707 (N_7707,N_7350,N_7393);
nand U7708 (N_7708,N_7591,N_7564);
nand U7709 (N_7709,N_7226,N_7426);
nand U7710 (N_7710,N_7419,N_7324);
xor U7711 (N_7711,N_7335,N_7425);
or U7712 (N_7712,N_7487,N_7578);
and U7713 (N_7713,N_7212,N_7378);
nor U7714 (N_7714,N_7490,N_7430);
or U7715 (N_7715,N_7259,N_7547);
xor U7716 (N_7716,N_7244,N_7346);
xnor U7717 (N_7717,N_7258,N_7421);
nand U7718 (N_7718,N_7585,N_7482);
and U7719 (N_7719,N_7360,N_7330);
or U7720 (N_7720,N_7219,N_7389);
or U7721 (N_7721,N_7495,N_7255);
nand U7722 (N_7722,N_7481,N_7559);
nand U7723 (N_7723,N_7285,N_7216);
nor U7724 (N_7724,N_7240,N_7353);
xnor U7725 (N_7725,N_7422,N_7364);
xor U7726 (N_7726,N_7246,N_7473);
and U7727 (N_7727,N_7560,N_7374);
nand U7728 (N_7728,N_7434,N_7595);
nand U7729 (N_7729,N_7408,N_7567);
nand U7730 (N_7730,N_7213,N_7409);
nor U7731 (N_7731,N_7401,N_7532);
nand U7732 (N_7732,N_7447,N_7599);
and U7733 (N_7733,N_7357,N_7552);
xnor U7734 (N_7734,N_7304,N_7516);
xnor U7735 (N_7735,N_7476,N_7200);
nor U7736 (N_7736,N_7400,N_7236);
xor U7737 (N_7737,N_7541,N_7484);
xor U7738 (N_7738,N_7316,N_7377);
and U7739 (N_7739,N_7438,N_7288);
xor U7740 (N_7740,N_7340,N_7268);
nor U7741 (N_7741,N_7411,N_7506);
nor U7742 (N_7742,N_7373,N_7549);
nor U7743 (N_7743,N_7501,N_7533);
nor U7744 (N_7744,N_7391,N_7497);
xor U7745 (N_7745,N_7249,N_7466);
or U7746 (N_7746,N_7307,N_7358);
xnor U7747 (N_7747,N_7338,N_7211);
or U7748 (N_7748,N_7519,N_7209);
or U7749 (N_7749,N_7207,N_7348);
and U7750 (N_7750,N_7248,N_7412);
nor U7751 (N_7751,N_7498,N_7298);
nand U7752 (N_7752,N_7493,N_7275);
and U7753 (N_7753,N_7237,N_7238);
and U7754 (N_7754,N_7523,N_7537);
or U7755 (N_7755,N_7287,N_7554);
nor U7756 (N_7756,N_7234,N_7573);
nand U7757 (N_7757,N_7224,N_7522);
nand U7758 (N_7758,N_7443,N_7548);
and U7759 (N_7759,N_7271,N_7306);
or U7760 (N_7760,N_7347,N_7309);
xnor U7761 (N_7761,N_7423,N_7592);
or U7762 (N_7762,N_7470,N_7584);
nor U7763 (N_7763,N_7215,N_7551);
nand U7764 (N_7764,N_7587,N_7386);
and U7765 (N_7765,N_7253,N_7556);
xnor U7766 (N_7766,N_7489,N_7232);
and U7767 (N_7767,N_7433,N_7204);
or U7768 (N_7768,N_7283,N_7352);
or U7769 (N_7769,N_7582,N_7245);
xor U7770 (N_7770,N_7437,N_7471);
and U7771 (N_7771,N_7530,N_7297);
and U7772 (N_7772,N_7205,N_7387);
nor U7773 (N_7773,N_7494,N_7220);
nor U7774 (N_7774,N_7254,N_7375);
nor U7775 (N_7775,N_7420,N_7383);
or U7776 (N_7776,N_7427,N_7397);
or U7777 (N_7777,N_7404,N_7460);
nand U7778 (N_7778,N_7321,N_7581);
nand U7779 (N_7779,N_7384,N_7455);
xor U7780 (N_7780,N_7313,N_7589);
xnor U7781 (N_7781,N_7318,N_7305);
xnor U7782 (N_7782,N_7449,N_7593);
or U7783 (N_7783,N_7598,N_7247);
nor U7784 (N_7784,N_7342,N_7415);
nand U7785 (N_7785,N_7376,N_7201);
xor U7786 (N_7786,N_7362,N_7311);
or U7787 (N_7787,N_7562,N_7472);
and U7788 (N_7788,N_7302,N_7542);
nor U7789 (N_7789,N_7572,N_7544);
nor U7790 (N_7790,N_7314,N_7545);
xnor U7791 (N_7791,N_7513,N_7452);
or U7792 (N_7792,N_7504,N_7459);
or U7793 (N_7793,N_7333,N_7440);
nand U7794 (N_7794,N_7445,N_7571);
xor U7795 (N_7795,N_7431,N_7511);
nor U7796 (N_7796,N_7325,N_7410);
or U7797 (N_7797,N_7485,N_7361);
nor U7798 (N_7798,N_7278,N_7272);
nor U7799 (N_7799,N_7509,N_7317);
nand U7800 (N_7800,N_7209,N_7243);
xnor U7801 (N_7801,N_7376,N_7274);
and U7802 (N_7802,N_7437,N_7243);
xor U7803 (N_7803,N_7478,N_7592);
nor U7804 (N_7804,N_7288,N_7566);
nand U7805 (N_7805,N_7515,N_7477);
nor U7806 (N_7806,N_7285,N_7312);
nand U7807 (N_7807,N_7525,N_7382);
or U7808 (N_7808,N_7482,N_7393);
nor U7809 (N_7809,N_7572,N_7476);
nand U7810 (N_7810,N_7351,N_7233);
and U7811 (N_7811,N_7385,N_7229);
or U7812 (N_7812,N_7578,N_7296);
nand U7813 (N_7813,N_7347,N_7267);
xnor U7814 (N_7814,N_7479,N_7279);
nor U7815 (N_7815,N_7500,N_7385);
nand U7816 (N_7816,N_7452,N_7379);
and U7817 (N_7817,N_7445,N_7494);
xor U7818 (N_7818,N_7252,N_7469);
or U7819 (N_7819,N_7439,N_7298);
nand U7820 (N_7820,N_7313,N_7266);
and U7821 (N_7821,N_7565,N_7550);
or U7822 (N_7822,N_7408,N_7493);
nand U7823 (N_7823,N_7442,N_7438);
and U7824 (N_7824,N_7336,N_7395);
xnor U7825 (N_7825,N_7329,N_7220);
nor U7826 (N_7826,N_7334,N_7363);
xnor U7827 (N_7827,N_7419,N_7380);
nand U7828 (N_7828,N_7319,N_7263);
xor U7829 (N_7829,N_7584,N_7563);
or U7830 (N_7830,N_7270,N_7479);
and U7831 (N_7831,N_7475,N_7239);
nor U7832 (N_7832,N_7443,N_7370);
or U7833 (N_7833,N_7420,N_7587);
nand U7834 (N_7834,N_7512,N_7473);
nand U7835 (N_7835,N_7216,N_7369);
nand U7836 (N_7836,N_7359,N_7280);
nand U7837 (N_7837,N_7323,N_7485);
nor U7838 (N_7838,N_7304,N_7577);
xnor U7839 (N_7839,N_7489,N_7314);
nand U7840 (N_7840,N_7487,N_7405);
nand U7841 (N_7841,N_7488,N_7461);
nand U7842 (N_7842,N_7403,N_7364);
nor U7843 (N_7843,N_7449,N_7599);
nor U7844 (N_7844,N_7406,N_7541);
and U7845 (N_7845,N_7267,N_7568);
nor U7846 (N_7846,N_7331,N_7527);
nand U7847 (N_7847,N_7540,N_7387);
or U7848 (N_7848,N_7568,N_7450);
nor U7849 (N_7849,N_7561,N_7566);
or U7850 (N_7850,N_7417,N_7552);
nand U7851 (N_7851,N_7576,N_7538);
nand U7852 (N_7852,N_7495,N_7516);
nor U7853 (N_7853,N_7273,N_7213);
or U7854 (N_7854,N_7461,N_7306);
and U7855 (N_7855,N_7315,N_7359);
or U7856 (N_7856,N_7485,N_7299);
xnor U7857 (N_7857,N_7423,N_7228);
nor U7858 (N_7858,N_7579,N_7331);
nor U7859 (N_7859,N_7548,N_7576);
nor U7860 (N_7860,N_7468,N_7396);
and U7861 (N_7861,N_7233,N_7301);
or U7862 (N_7862,N_7594,N_7253);
or U7863 (N_7863,N_7265,N_7350);
and U7864 (N_7864,N_7383,N_7248);
nor U7865 (N_7865,N_7467,N_7437);
nand U7866 (N_7866,N_7462,N_7483);
and U7867 (N_7867,N_7522,N_7563);
and U7868 (N_7868,N_7491,N_7429);
and U7869 (N_7869,N_7383,N_7567);
and U7870 (N_7870,N_7368,N_7232);
and U7871 (N_7871,N_7387,N_7362);
or U7872 (N_7872,N_7458,N_7524);
xnor U7873 (N_7873,N_7395,N_7213);
and U7874 (N_7874,N_7229,N_7529);
nor U7875 (N_7875,N_7504,N_7379);
nor U7876 (N_7876,N_7553,N_7246);
or U7877 (N_7877,N_7262,N_7401);
nor U7878 (N_7878,N_7593,N_7592);
xnor U7879 (N_7879,N_7566,N_7349);
xor U7880 (N_7880,N_7253,N_7514);
and U7881 (N_7881,N_7479,N_7211);
and U7882 (N_7882,N_7213,N_7279);
and U7883 (N_7883,N_7383,N_7230);
nor U7884 (N_7884,N_7414,N_7516);
xnor U7885 (N_7885,N_7353,N_7253);
nand U7886 (N_7886,N_7311,N_7514);
nor U7887 (N_7887,N_7366,N_7592);
nand U7888 (N_7888,N_7583,N_7201);
xnor U7889 (N_7889,N_7300,N_7350);
nor U7890 (N_7890,N_7549,N_7494);
and U7891 (N_7891,N_7537,N_7516);
nor U7892 (N_7892,N_7561,N_7374);
xnor U7893 (N_7893,N_7290,N_7454);
nor U7894 (N_7894,N_7573,N_7525);
nand U7895 (N_7895,N_7388,N_7253);
nand U7896 (N_7896,N_7293,N_7248);
nor U7897 (N_7897,N_7364,N_7281);
and U7898 (N_7898,N_7598,N_7260);
and U7899 (N_7899,N_7272,N_7341);
or U7900 (N_7900,N_7301,N_7565);
and U7901 (N_7901,N_7380,N_7209);
nand U7902 (N_7902,N_7585,N_7314);
nor U7903 (N_7903,N_7414,N_7208);
or U7904 (N_7904,N_7261,N_7204);
nor U7905 (N_7905,N_7378,N_7488);
xnor U7906 (N_7906,N_7582,N_7400);
nor U7907 (N_7907,N_7475,N_7549);
and U7908 (N_7908,N_7595,N_7272);
nand U7909 (N_7909,N_7276,N_7447);
nor U7910 (N_7910,N_7324,N_7269);
or U7911 (N_7911,N_7450,N_7564);
nor U7912 (N_7912,N_7492,N_7578);
nor U7913 (N_7913,N_7378,N_7407);
nor U7914 (N_7914,N_7597,N_7250);
nand U7915 (N_7915,N_7415,N_7532);
or U7916 (N_7916,N_7241,N_7547);
and U7917 (N_7917,N_7298,N_7267);
nand U7918 (N_7918,N_7305,N_7458);
xnor U7919 (N_7919,N_7357,N_7214);
and U7920 (N_7920,N_7569,N_7336);
nor U7921 (N_7921,N_7519,N_7230);
nor U7922 (N_7922,N_7582,N_7519);
xor U7923 (N_7923,N_7381,N_7457);
nor U7924 (N_7924,N_7541,N_7225);
nor U7925 (N_7925,N_7276,N_7481);
nand U7926 (N_7926,N_7574,N_7345);
and U7927 (N_7927,N_7491,N_7202);
or U7928 (N_7928,N_7563,N_7493);
nor U7929 (N_7929,N_7501,N_7575);
nand U7930 (N_7930,N_7247,N_7547);
nand U7931 (N_7931,N_7205,N_7208);
or U7932 (N_7932,N_7396,N_7248);
or U7933 (N_7933,N_7283,N_7521);
or U7934 (N_7934,N_7229,N_7425);
xor U7935 (N_7935,N_7238,N_7251);
nand U7936 (N_7936,N_7581,N_7305);
xor U7937 (N_7937,N_7246,N_7389);
or U7938 (N_7938,N_7597,N_7380);
nor U7939 (N_7939,N_7529,N_7407);
or U7940 (N_7940,N_7247,N_7408);
or U7941 (N_7941,N_7527,N_7201);
xor U7942 (N_7942,N_7588,N_7441);
nor U7943 (N_7943,N_7506,N_7599);
nor U7944 (N_7944,N_7512,N_7427);
nand U7945 (N_7945,N_7208,N_7202);
xnor U7946 (N_7946,N_7283,N_7322);
and U7947 (N_7947,N_7337,N_7394);
nor U7948 (N_7948,N_7264,N_7404);
xor U7949 (N_7949,N_7357,N_7279);
nand U7950 (N_7950,N_7207,N_7515);
or U7951 (N_7951,N_7484,N_7358);
and U7952 (N_7952,N_7516,N_7290);
and U7953 (N_7953,N_7447,N_7515);
nand U7954 (N_7954,N_7431,N_7595);
nand U7955 (N_7955,N_7285,N_7252);
or U7956 (N_7956,N_7560,N_7591);
or U7957 (N_7957,N_7310,N_7395);
or U7958 (N_7958,N_7221,N_7457);
and U7959 (N_7959,N_7401,N_7251);
xnor U7960 (N_7960,N_7326,N_7541);
nor U7961 (N_7961,N_7461,N_7492);
nand U7962 (N_7962,N_7536,N_7255);
xnor U7963 (N_7963,N_7420,N_7222);
and U7964 (N_7964,N_7392,N_7315);
and U7965 (N_7965,N_7244,N_7268);
nor U7966 (N_7966,N_7212,N_7286);
or U7967 (N_7967,N_7515,N_7469);
or U7968 (N_7968,N_7598,N_7450);
and U7969 (N_7969,N_7410,N_7320);
nand U7970 (N_7970,N_7429,N_7216);
nor U7971 (N_7971,N_7517,N_7237);
nor U7972 (N_7972,N_7212,N_7238);
nor U7973 (N_7973,N_7441,N_7405);
and U7974 (N_7974,N_7577,N_7354);
xor U7975 (N_7975,N_7487,N_7389);
and U7976 (N_7976,N_7273,N_7467);
or U7977 (N_7977,N_7335,N_7551);
or U7978 (N_7978,N_7579,N_7401);
nand U7979 (N_7979,N_7595,N_7395);
or U7980 (N_7980,N_7295,N_7255);
and U7981 (N_7981,N_7380,N_7576);
xnor U7982 (N_7982,N_7323,N_7490);
nor U7983 (N_7983,N_7341,N_7316);
xnor U7984 (N_7984,N_7398,N_7481);
and U7985 (N_7985,N_7563,N_7424);
and U7986 (N_7986,N_7404,N_7552);
or U7987 (N_7987,N_7221,N_7382);
nor U7988 (N_7988,N_7255,N_7346);
xor U7989 (N_7989,N_7259,N_7331);
and U7990 (N_7990,N_7355,N_7421);
and U7991 (N_7991,N_7245,N_7512);
and U7992 (N_7992,N_7478,N_7540);
or U7993 (N_7993,N_7536,N_7350);
and U7994 (N_7994,N_7317,N_7315);
or U7995 (N_7995,N_7373,N_7303);
or U7996 (N_7996,N_7519,N_7382);
or U7997 (N_7997,N_7595,N_7448);
nand U7998 (N_7998,N_7509,N_7591);
nor U7999 (N_7999,N_7493,N_7489);
nand U8000 (N_8000,N_7786,N_7637);
xnor U8001 (N_8001,N_7725,N_7681);
xor U8002 (N_8002,N_7688,N_7694);
xor U8003 (N_8003,N_7923,N_7860);
and U8004 (N_8004,N_7793,N_7812);
nor U8005 (N_8005,N_7900,N_7802);
nor U8006 (N_8006,N_7868,N_7891);
or U8007 (N_8007,N_7924,N_7729);
and U8008 (N_8008,N_7643,N_7787);
xnor U8009 (N_8009,N_7815,N_7999);
or U8010 (N_8010,N_7823,N_7774);
and U8011 (N_8011,N_7761,N_7819);
or U8012 (N_8012,N_7996,N_7913);
nand U8013 (N_8013,N_7888,N_7986);
and U8014 (N_8014,N_7941,N_7696);
xor U8015 (N_8015,N_7775,N_7908);
xor U8016 (N_8016,N_7932,N_7976);
xnor U8017 (N_8017,N_7695,N_7794);
nor U8018 (N_8018,N_7656,N_7658);
nand U8019 (N_8019,N_7828,N_7843);
and U8020 (N_8020,N_7997,N_7871);
nand U8021 (N_8021,N_7726,N_7717);
or U8022 (N_8022,N_7903,N_7773);
nor U8023 (N_8023,N_7865,N_7767);
nand U8024 (N_8024,N_7790,N_7984);
xnor U8025 (N_8025,N_7857,N_7649);
xor U8026 (N_8026,N_7845,N_7937);
or U8027 (N_8027,N_7619,N_7893);
nand U8028 (N_8028,N_7632,N_7780);
nand U8029 (N_8029,N_7973,N_7720);
nand U8030 (N_8030,N_7675,N_7947);
xnor U8031 (N_8031,N_7910,N_7801);
or U8032 (N_8032,N_7712,N_7657);
or U8033 (N_8033,N_7746,N_7853);
or U8034 (N_8034,N_7995,N_7600);
nand U8035 (N_8035,N_7617,N_7735);
nand U8036 (N_8036,N_7918,N_7931);
nor U8037 (N_8037,N_7764,N_7938);
and U8038 (N_8038,N_7710,N_7919);
and U8039 (N_8039,N_7756,N_7651);
nor U8040 (N_8040,N_7623,N_7606);
nor U8041 (N_8041,N_7814,N_7784);
and U8042 (N_8042,N_7856,N_7838);
or U8043 (N_8043,N_7736,N_7977);
nor U8044 (N_8044,N_7788,N_7612);
or U8045 (N_8045,N_7618,N_7895);
nor U8046 (N_8046,N_7816,N_7849);
or U8047 (N_8047,N_7677,N_7882);
xor U8048 (N_8048,N_7806,N_7604);
or U8049 (N_8049,N_7782,N_7754);
nand U8050 (N_8050,N_7669,N_7732);
and U8051 (N_8051,N_7988,N_7930);
xnor U8052 (N_8052,N_7701,N_7832);
and U8053 (N_8053,N_7956,N_7993);
and U8054 (N_8054,N_7664,N_7862);
nand U8055 (N_8055,N_7940,N_7740);
or U8056 (N_8056,N_7797,N_7961);
and U8057 (N_8057,N_7731,N_7934);
nand U8058 (N_8058,N_7834,N_7837);
nor U8059 (N_8059,N_7607,N_7825);
xor U8060 (N_8060,N_7646,N_7647);
nand U8061 (N_8061,N_7808,N_7629);
xor U8062 (N_8062,N_7948,N_7750);
or U8063 (N_8063,N_7749,N_7951);
nand U8064 (N_8064,N_7822,N_7783);
nor U8065 (N_8065,N_7942,N_7943);
nand U8066 (N_8066,N_7693,N_7616);
or U8067 (N_8067,N_7914,N_7689);
nor U8068 (N_8068,N_7737,N_7827);
xnor U8069 (N_8069,N_7809,N_7768);
xnor U8070 (N_8070,N_7707,N_7610);
xnor U8071 (N_8071,N_7818,N_7645);
nand U8072 (N_8072,N_7652,N_7901);
or U8073 (N_8073,N_7846,N_7641);
or U8074 (N_8074,N_7640,N_7660);
or U8075 (N_8075,N_7676,N_7799);
or U8076 (N_8076,N_7962,N_7686);
nand U8077 (N_8077,N_7939,N_7699);
and U8078 (N_8078,N_7602,N_7748);
or U8079 (N_8079,N_7734,N_7906);
nor U8080 (N_8080,N_7839,N_7826);
nor U8081 (N_8081,N_7771,N_7803);
or U8082 (N_8082,N_7776,N_7628);
or U8083 (N_8083,N_7867,N_7935);
nor U8084 (N_8084,N_7911,N_7980);
nor U8085 (N_8085,N_7648,N_7899);
nand U8086 (N_8086,N_7608,N_7795);
nor U8087 (N_8087,N_7892,N_7929);
nor U8088 (N_8088,N_7890,N_7905);
nand U8089 (N_8089,N_7668,N_7998);
xor U8090 (N_8090,N_7915,N_7896);
xnor U8091 (N_8091,N_7703,N_7683);
nand U8092 (N_8092,N_7738,N_7885);
and U8093 (N_8093,N_7863,N_7622);
nand U8094 (N_8094,N_7912,N_7829);
or U8095 (N_8095,N_7954,N_7760);
nand U8096 (N_8096,N_7638,N_7851);
nor U8097 (N_8097,N_7945,N_7855);
or U8098 (N_8098,N_7621,N_7858);
nor U8099 (N_8099,N_7659,N_7848);
nand U8100 (N_8100,N_7953,N_7836);
or U8101 (N_8101,N_7789,N_7679);
or U8102 (N_8102,N_7672,N_7990);
nand U8103 (N_8103,N_7982,N_7747);
xor U8104 (N_8104,N_7922,N_7723);
nor U8105 (N_8105,N_7824,N_7928);
nor U8106 (N_8106,N_7739,N_7876);
or U8107 (N_8107,N_7975,N_7753);
nor U8108 (N_8108,N_7691,N_7921);
or U8109 (N_8109,N_7950,N_7957);
nand U8110 (N_8110,N_7972,N_7633);
nor U8111 (N_8111,N_7847,N_7830);
xnor U8112 (N_8112,N_7878,N_7981);
or U8113 (N_8113,N_7674,N_7969);
nand U8114 (N_8114,N_7682,N_7968);
xnor U8115 (N_8115,N_7898,N_7880);
nand U8116 (N_8116,N_7971,N_7706);
nor U8117 (N_8117,N_7680,N_7964);
xnor U8118 (N_8118,N_7626,N_7779);
or U8119 (N_8119,N_7983,N_7770);
xnor U8120 (N_8120,N_7627,N_7960);
nor U8121 (N_8121,N_7917,N_7639);
or U8122 (N_8122,N_7642,N_7745);
xor U8123 (N_8123,N_7650,N_7897);
nand U8124 (N_8124,N_7869,N_7722);
nand U8125 (N_8125,N_7979,N_7730);
or U8126 (N_8126,N_7821,N_7907);
xor U8127 (N_8127,N_7667,N_7716);
xor U8128 (N_8128,N_7727,N_7886);
or U8129 (N_8129,N_7615,N_7909);
xnor U8130 (N_8130,N_7673,N_7663);
nand U8131 (N_8131,N_7798,N_7835);
and U8132 (N_8132,N_7927,N_7841);
or U8133 (N_8133,N_7958,N_7665);
xnor U8134 (N_8134,N_7967,N_7872);
nor U8135 (N_8135,N_7850,N_7894);
nand U8136 (N_8136,N_7758,N_7970);
nor U8137 (N_8137,N_7772,N_7833);
xnor U8138 (N_8138,N_7933,N_7709);
or U8139 (N_8139,N_7741,N_7743);
and U8140 (N_8140,N_7752,N_7854);
or U8141 (N_8141,N_7733,N_7728);
nor U8142 (N_8142,N_7671,N_7702);
and U8143 (N_8143,N_7714,N_7655);
nor U8144 (N_8144,N_7859,N_7884);
nand U8145 (N_8145,N_7724,N_7611);
or U8146 (N_8146,N_7920,N_7989);
xor U8147 (N_8147,N_7634,N_7994);
xnor U8148 (N_8148,N_7654,N_7791);
nor U8149 (N_8149,N_7718,N_7719);
nor U8150 (N_8150,N_7813,N_7800);
xor U8151 (N_8151,N_7936,N_7966);
or U8152 (N_8152,N_7889,N_7708);
nand U8153 (N_8153,N_7873,N_7778);
and U8154 (N_8154,N_7875,N_7662);
xnor U8155 (N_8155,N_7965,N_7762);
nand U8156 (N_8156,N_7620,N_7631);
nand U8157 (N_8157,N_7944,N_7796);
xor U8158 (N_8158,N_7817,N_7601);
and U8159 (N_8159,N_7624,N_7879);
nand U8160 (N_8160,N_7991,N_7705);
and U8161 (N_8161,N_7811,N_7810);
nor U8162 (N_8162,N_7690,N_7766);
or U8163 (N_8163,N_7613,N_7751);
and U8164 (N_8164,N_7792,N_7804);
xnor U8165 (N_8165,N_7883,N_7763);
or U8166 (N_8166,N_7887,N_7955);
nand U8167 (N_8167,N_7755,N_7757);
and U8168 (N_8168,N_7781,N_7925);
xnor U8169 (N_8169,N_7916,N_7700);
nor U8170 (N_8170,N_7952,N_7877);
xor U8171 (N_8171,N_7713,N_7978);
nor U8172 (N_8172,N_7874,N_7744);
or U8173 (N_8173,N_7864,N_7692);
nor U8174 (N_8174,N_7605,N_7635);
nand U8175 (N_8175,N_7742,N_7870);
nor U8176 (N_8176,N_7670,N_7987);
xor U8177 (N_8177,N_7685,N_7625);
and U8178 (N_8178,N_7926,N_7661);
nand U8179 (N_8179,N_7777,N_7666);
xor U8180 (N_8180,N_7852,N_7636);
and U8181 (N_8181,N_7866,N_7603);
nor U8182 (N_8182,N_7711,N_7721);
and U8183 (N_8183,N_7684,N_7904);
nand U8184 (N_8184,N_7785,N_7678);
xnor U8185 (N_8185,N_7653,N_7609);
xor U8186 (N_8186,N_7614,N_7963);
and U8187 (N_8187,N_7881,N_7630);
and U8188 (N_8188,N_7985,N_7807);
nor U8189 (N_8189,N_7992,N_7974);
and U8190 (N_8190,N_7946,N_7959);
nand U8191 (N_8191,N_7715,N_7759);
xor U8192 (N_8192,N_7805,N_7840);
and U8193 (N_8193,N_7820,N_7769);
and U8194 (N_8194,N_7765,N_7644);
nand U8195 (N_8195,N_7697,N_7949);
nand U8196 (N_8196,N_7704,N_7831);
xor U8197 (N_8197,N_7842,N_7861);
and U8198 (N_8198,N_7844,N_7902);
nand U8199 (N_8199,N_7698,N_7687);
or U8200 (N_8200,N_7768,N_7630);
or U8201 (N_8201,N_7632,N_7932);
nand U8202 (N_8202,N_7732,N_7714);
and U8203 (N_8203,N_7713,N_7732);
nand U8204 (N_8204,N_7721,N_7801);
or U8205 (N_8205,N_7815,N_7624);
nor U8206 (N_8206,N_7739,N_7752);
and U8207 (N_8207,N_7711,N_7986);
xnor U8208 (N_8208,N_7893,N_7938);
nor U8209 (N_8209,N_7621,N_7850);
and U8210 (N_8210,N_7862,N_7808);
and U8211 (N_8211,N_7815,N_7697);
xnor U8212 (N_8212,N_7779,N_7616);
or U8213 (N_8213,N_7763,N_7681);
or U8214 (N_8214,N_7772,N_7710);
and U8215 (N_8215,N_7764,N_7904);
nor U8216 (N_8216,N_7882,N_7641);
xnor U8217 (N_8217,N_7732,N_7976);
nand U8218 (N_8218,N_7852,N_7811);
or U8219 (N_8219,N_7604,N_7652);
nand U8220 (N_8220,N_7711,N_7952);
xnor U8221 (N_8221,N_7826,N_7808);
or U8222 (N_8222,N_7839,N_7857);
and U8223 (N_8223,N_7609,N_7744);
xnor U8224 (N_8224,N_7874,N_7894);
or U8225 (N_8225,N_7940,N_7609);
nor U8226 (N_8226,N_7665,N_7823);
xor U8227 (N_8227,N_7647,N_7775);
nor U8228 (N_8228,N_7613,N_7844);
nor U8229 (N_8229,N_7866,N_7770);
xor U8230 (N_8230,N_7698,N_7701);
xor U8231 (N_8231,N_7751,N_7933);
or U8232 (N_8232,N_7856,N_7975);
nor U8233 (N_8233,N_7601,N_7681);
nor U8234 (N_8234,N_7816,N_7627);
and U8235 (N_8235,N_7965,N_7884);
nand U8236 (N_8236,N_7866,N_7739);
nand U8237 (N_8237,N_7938,N_7996);
and U8238 (N_8238,N_7741,N_7640);
nor U8239 (N_8239,N_7757,N_7878);
nor U8240 (N_8240,N_7720,N_7929);
xnor U8241 (N_8241,N_7706,N_7837);
or U8242 (N_8242,N_7724,N_7965);
nand U8243 (N_8243,N_7850,N_7799);
or U8244 (N_8244,N_7969,N_7904);
xnor U8245 (N_8245,N_7691,N_7786);
and U8246 (N_8246,N_7801,N_7908);
or U8247 (N_8247,N_7727,N_7681);
xor U8248 (N_8248,N_7965,N_7603);
xor U8249 (N_8249,N_7692,N_7776);
or U8250 (N_8250,N_7916,N_7818);
and U8251 (N_8251,N_7757,N_7694);
nand U8252 (N_8252,N_7619,N_7615);
nand U8253 (N_8253,N_7865,N_7841);
or U8254 (N_8254,N_7824,N_7812);
or U8255 (N_8255,N_7807,N_7668);
or U8256 (N_8256,N_7825,N_7742);
and U8257 (N_8257,N_7673,N_7878);
nor U8258 (N_8258,N_7619,N_7973);
nand U8259 (N_8259,N_7911,N_7868);
xor U8260 (N_8260,N_7752,N_7692);
xor U8261 (N_8261,N_7878,N_7974);
xor U8262 (N_8262,N_7843,N_7738);
xor U8263 (N_8263,N_7640,N_7811);
or U8264 (N_8264,N_7792,N_7623);
or U8265 (N_8265,N_7875,N_7813);
nor U8266 (N_8266,N_7675,N_7611);
xnor U8267 (N_8267,N_7955,N_7914);
xnor U8268 (N_8268,N_7868,N_7622);
or U8269 (N_8269,N_7629,N_7735);
or U8270 (N_8270,N_7735,N_7732);
nor U8271 (N_8271,N_7714,N_7965);
or U8272 (N_8272,N_7600,N_7811);
xor U8273 (N_8273,N_7669,N_7854);
nor U8274 (N_8274,N_7782,N_7685);
xor U8275 (N_8275,N_7703,N_7613);
or U8276 (N_8276,N_7892,N_7663);
nand U8277 (N_8277,N_7761,N_7942);
or U8278 (N_8278,N_7768,N_7830);
nand U8279 (N_8279,N_7627,N_7933);
nand U8280 (N_8280,N_7985,N_7906);
xor U8281 (N_8281,N_7979,N_7767);
and U8282 (N_8282,N_7931,N_7928);
or U8283 (N_8283,N_7906,N_7640);
and U8284 (N_8284,N_7829,N_7951);
and U8285 (N_8285,N_7748,N_7738);
nand U8286 (N_8286,N_7866,N_7925);
nor U8287 (N_8287,N_7852,N_7767);
nand U8288 (N_8288,N_7664,N_7888);
and U8289 (N_8289,N_7820,N_7829);
and U8290 (N_8290,N_7875,N_7787);
nor U8291 (N_8291,N_7946,N_7603);
nor U8292 (N_8292,N_7824,N_7745);
xor U8293 (N_8293,N_7807,N_7799);
and U8294 (N_8294,N_7735,N_7869);
nand U8295 (N_8295,N_7685,N_7714);
xnor U8296 (N_8296,N_7648,N_7945);
nor U8297 (N_8297,N_7848,N_7624);
or U8298 (N_8298,N_7749,N_7745);
xor U8299 (N_8299,N_7746,N_7960);
xor U8300 (N_8300,N_7704,N_7702);
nor U8301 (N_8301,N_7772,N_7947);
nand U8302 (N_8302,N_7874,N_7695);
or U8303 (N_8303,N_7884,N_7935);
xor U8304 (N_8304,N_7680,N_7726);
or U8305 (N_8305,N_7791,N_7942);
or U8306 (N_8306,N_7849,N_7863);
nand U8307 (N_8307,N_7852,N_7690);
nand U8308 (N_8308,N_7611,N_7882);
xnor U8309 (N_8309,N_7944,N_7626);
nor U8310 (N_8310,N_7895,N_7931);
or U8311 (N_8311,N_7791,N_7950);
and U8312 (N_8312,N_7848,N_7756);
xor U8313 (N_8313,N_7969,N_7783);
and U8314 (N_8314,N_7897,N_7727);
or U8315 (N_8315,N_7618,N_7745);
nand U8316 (N_8316,N_7644,N_7633);
nor U8317 (N_8317,N_7987,N_7607);
xor U8318 (N_8318,N_7898,N_7815);
or U8319 (N_8319,N_7908,N_7662);
and U8320 (N_8320,N_7737,N_7716);
nor U8321 (N_8321,N_7988,N_7628);
xnor U8322 (N_8322,N_7951,N_7801);
and U8323 (N_8323,N_7823,N_7738);
xor U8324 (N_8324,N_7729,N_7864);
nand U8325 (N_8325,N_7702,N_7755);
and U8326 (N_8326,N_7876,N_7914);
nor U8327 (N_8327,N_7728,N_7627);
xor U8328 (N_8328,N_7629,N_7954);
or U8329 (N_8329,N_7775,N_7734);
and U8330 (N_8330,N_7698,N_7736);
xor U8331 (N_8331,N_7978,N_7773);
xor U8332 (N_8332,N_7781,N_7911);
xor U8333 (N_8333,N_7698,N_7626);
nand U8334 (N_8334,N_7804,N_7667);
nor U8335 (N_8335,N_7713,N_7781);
and U8336 (N_8336,N_7684,N_7845);
or U8337 (N_8337,N_7638,N_7827);
nand U8338 (N_8338,N_7642,N_7743);
or U8339 (N_8339,N_7688,N_7987);
and U8340 (N_8340,N_7670,N_7820);
nor U8341 (N_8341,N_7903,N_7657);
and U8342 (N_8342,N_7825,N_7774);
nor U8343 (N_8343,N_7895,N_7821);
and U8344 (N_8344,N_7831,N_7896);
and U8345 (N_8345,N_7701,N_7977);
nand U8346 (N_8346,N_7998,N_7914);
or U8347 (N_8347,N_7659,N_7968);
nand U8348 (N_8348,N_7912,N_7816);
nand U8349 (N_8349,N_7798,N_7767);
and U8350 (N_8350,N_7812,N_7818);
or U8351 (N_8351,N_7823,N_7959);
xor U8352 (N_8352,N_7995,N_7642);
or U8353 (N_8353,N_7990,N_7681);
or U8354 (N_8354,N_7802,N_7978);
and U8355 (N_8355,N_7790,N_7887);
nand U8356 (N_8356,N_7975,N_7914);
and U8357 (N_8357,N_7780,N_7938);
xnor U8358 (N_8358,N_7739,N_7906);
nand U8359 (N_8359,N_7902,N_7922);
nor U8360 (N_8360,N_7643,N_7756);
nor U8361 (N_8361,N_7776,N_7960);
nand U8362 (N_8362,N_7700,N_7601);
nand U8363 (N_8363,N_7921,N_7957);
and U8364 (N_8364,N_7742,N_7810);
nor U8365 (N_8365,N_7636,N_7734);
xor U8366 (N_8366,N_7786,N_7601);
nand U8367 (N_8367,N_7623,N_7649);
and U8368 (N_8368,N_7977,N_7880);
xnor U8369 (N_8369,N_7855,N_7890);
and U8370 (N_8370,N_7783,N_7801);
and U8371 (N_8371,N_7761,N_7979);
nand U8372 (N_8372,N_7844,N_7609);
or U8373 (N_8373,N_7642,N_7810);
or U8374 (N_8374,N_7637,N_7830);
nor U8375 (N_8375,N_7610,N_7953);
nand U8376 (N_8376,N_7962,N_7951);
nor U8377 (N_8377,N_7755,N_7602);
or U8378 (N_8378,N_7841,N_7844);
or U8379 (N_8379,N_7732,N_7630);
and U8380 (N_8380,N_7644,N_7818);
or U8381 (N_8381,N_7891,N_7841);
xor U8382 (N_8382,N_7933,N_7802);
and U8383 (N_8383,N_7688,N_7862);
nand U8384 (N_8384,N_7799,N_7887);
xnor U8385 (N_8385,N_7757,N_7805);
or U8386 (N_8386,N_7622,N_7843);
nand U8387 (N_8387,N_7983,N_7902);
or U8388 (N_8388,N_7987,N_7831);
and U8389 (N_8389,N_7679,N_7694);
or U8390 (N_8390,N_7980,N_7617);
xor U8391 (N_8391,N_7716,N_7870);
nand U8392 (N_8392,N_7870,N_7660);
nand U8393 (N_8393,N_7602,N_7688);
nor U8394 (N_8394,N_7850,N_7983);
or U8395 (N_8395,N_7934,N_7929);
nand U8396 (N_8396,N_7936,N_7848);
nand U8397 (N_8397,N_7967,N_7762);
nand U8398 (N_8398,N_7926,N_7680);
nand U8399 (N_8399,N_7860,N_7628);
nor U8400 (N_8400,N_8226,N_8095);
nor U8401 (N_8401,N_8307,N_8105);
xor U8402 (N_8402,N_8057,N_8238);
xnor U8403 (N_8403,N_8077,N_8394);
nor U8404 (N_8404,N_8388,N_8175);
xnor U8405 (N_8405,N_8355,N_8348);
xor U8406 (N_8406,N_8242,N_8241);
or U8407 (N_8407,N_8276,N_8194);
nor U8408 (N_8408,N_8038,N_8390);
or U8409 (N_8409,N_8033,N_8032);
or U8410 (N_8410,N_8325,N_8331);
nor U8411 (N_8411,N_8110,N_8120);
or U8412 (N_8412,N_8013,N_8106);
xor U8413 (N_8413,N_8353,N_8220);
nand U8414 (N_8414,N_8107,N_8117);
nand U8415 (N_8415,N_8297,N_8101);
nand U8416 (N_8416,N_8014,N_8396);
and U8417 (N_8417,N_8162,N_8185);
xor U8418 (N_8418,N_8196,N_8158);
nand U8419 (N_8419,N_8367,N_8187);
or U8420 (N_8420,N_8042,N_8317);
or U8421 (N_8421,N_8228,N_8025);
and U8422 (N_8422,N_8052,N_8089);
or U8423 (N_8423,N_8056,N_8362);
or U8424 (N_8424,N_8249,N_8321);
or U8425 (N_8425,N_8364,N_8210);
nor U8426 (N_8426,N_8182,N_8133);
nand U8427 (N_8427,N_8009,N_8229);
nand U8428 (N_8428,N_8280,N_8380);
and U8429 (N_8429,N_8094,N_8285);
nor U8430 (N_8430,N_8327,N_8151);
nor U8431 (N_8431,N_8197,N_8188);
nor U8432 (N_8432,N_8186,N_8000);
and U8433 (N_8433,N_8377,N_8097);
xnor U8434 (N_8434,N_8222,N_8174);
or U8435 (N_8435,N_8273,N_8172);
nor U8436 (N_8436,N_8247,N_8055);
xor U8437 (N_8437,N_8050,N_8116);
xnor U8438 (N_8438,N_8206,N_8250);
nor U8439 (N_8439,N_8119,N_8277);
nand U8440 (N_8440,N_8254,N_8034);
nand U8441 (N_8441,N_8130,N_8230);
or U8442 (N_8442,N_8045,N_8062);
and U8443 (N_8443,N_8223,N_8112);
and U8444 (N_8444,N_8121,N_8350);
nand U8445 (N_8445,N_8272,N_8310);
and U8446 (N_8446,N_8392,N_8290);
nand U8447 (N_8447,N_8203,N_8345);
and U8448 (N_8448,N_8176,N_8083);
nor U8449 (N_8449,N_8265,N_8069);
or U8450 (N_8450,N_8361,N_8385);
nand U8451 (N_8451,N_8293,N_8067);
or U8452 (N_8452,N_8007,N_8227);
nand U8453 (N_8453,N_8259,N_8308);
or U8454 (N_8454,N_8098,N_8044);
nor U8455 (N_8455,N_8163,N_8003);
nor U8456 (N_8456,N_8340,N_8023);
and U8457 (N_8457,N_8011,N_8258);
nor U8458 (N_8458,N_8167,N_8193);
nand U8459 (N_8459,N_8125,N_8204);
nor U8460 (N_8460,N_8066,N_8026);
nand U8461 (N_8461,N_8309,N_8278);
nor U8462 (N_8462,N_8379,N_8306);
xnor U8463 (N_8463,N_8398,N_8156);
nor U8464 (N_8464,N_8288,N_8261);
and U8465 (N_8465,N_8113,N_8147);
or U8466 (N_8466,N_8202,N_8359);
and U8467 (N_8467,N_8161,N_8287);
or U8468 (N_8468,N_8356,N_8240);
nand U8469 (N_8469,N_8036,N_8271);
or U8470 (N_8470,N_8256,N_8096);
nor U8471 (N_8471,N_8257,N_8386);
and U8472 (N_8472,N_8053,N_8005);
nor U8473 (N_8473,N_8059,N_8144);
nand U8474 (N_8474,N_8328,N_8024);
nand U8475 (N_8475,N_8150,N_8270);
xor U8476 (N_8476,N_8252,N_8275);
and U8477 (N_8477,N_8081,N_8199);
nor U8478 (N_8478,N_8114,N_8141);
or U8479 (N_8479,N_8260,N_8195);
nor U8480 (N_8480,N_8311,N_8352);
xnor U8481 (N_8481,N_8375,N_8207);
or U8482 (N_8482,N_8366,N_8086);
or U8483 (N_8483,N_8231,N_8248);
and U8484 (N_8484,N_8164,N_8082);
xor U8485 (N_8485,N_8181,N_8374);
or U8486 (N_8486,N_8190,N_8395);
xor U8487 (N_8487,N_8233,N_8319);
or U8488 (N_8488,N_8103,N_8200);
xnor U8489 (N_8489,N_8216,N_8330);
nand U8490 (N_8490,N_8335,N_8041);
nor U8491 (N_8491,N_8313,N_8262);
xnor U8492 (N_8492,N_8004,N_8111);
and U8493 (N_8493,N_8370,N_8169);
or U8494 (N_8494,N_8138,N_8320);
or U8495 (N_8495,N_8006,N_8279);
or U8496 (N_8496,N_8152,N_8387);
and U8497 (N_8497,N_8391,N_8266);
or U8498 (N_8498,N_8088,N_8142);
and U8499 (N_8499,N_8078,N_8232);
xor U8500 (N_8500,N_8170,N_8047);
or U8501 (N_8501,N_8002,N_8269);
nor U8502 (N_8502,N_8336,N_8393);
or U8503 (N_8503,N_8218,N_8302);
xnor U8504 (N_8504,N_8318,N_8145);
nand U8505 (N_8505,N_8137,N_8104);
nand U8506 (N_8506,N_8108,N_8322);
or U8507 (N_8507,N_8217,N_8018);
or U8508 (N_8508,N_8191,N_8039);
nor U8509 (N_8509,N_8389,N_8369);
xor U8510 (N_8510,N_8068,N_8093);
nor U8511 (N_8511,N_8058,N_8166);
and U8512 (N_8512,N_8008,N_8295);
and U8513 (N_8513,N_8284,N_8315);
or U8514 (N_8514,N_8341,N_8001);
nand U8515 (N_8515,N_8148,N_8236);
xnor U8516 (N_8516,N_8010,N_8134);
nor U8517 (N_8517,N_8209,N_8109);
xor U8518 (N_8518,N_8263,N_8159);
xnor U8519 (N_8519,N_8099,N_8128);
and U8520 (N_8520,N_8212,N_8192);
or U8521 (N_8521,N_8102,N_8079);
nor U8522 (N_8522,N_8296,N_8132);
xnor U8523 (N_8523,N_8333,N_8245);
xor U8524 (N_8524,N_8063,N_8085);
xor U8525 (N_8525,N_8267,N_8211);
or U8526 (N_8526,N_8224,N_8243);
xor U8527 (N_8527,N_8129,N_8179);
nor U8528 (N_8528,N_8100,N_8015);
xnor U8529 (N_8529,N_8251,N_8115);
xor U8530 (N_8530,N_8381,N_8301);
and U8531 (N_8531,N_8118,N_8189);
nor U8532 (N_8532,N_8294,N_8316);
xnor U8533 (N_8533,N_8087,N_8339);
nor U8534 (N_8534,N_8084,N_8289);
nor U8535 (N_8535,N_8153,N_8031);
nor U8536 (N_8536,N_8213,N_8074);
nor U8537 (N_8537,N_8139,N_8040);
nand U8538 (N_8538,N_8171,N_8299);
xnor U8539 (N_8539,N_8030,N_8046);
and U8540 (N_8540,N_8360,N_8126);
nand U8541 (N_8541,N_8165,N_8239);
and U8542 (N_8542,N_8146,N_8051);
or U8543 (N_8543,N_8037,N_8073);
xnor U8544 (N_8544,N_8208,N_8149);
or U8545 (N_8545,N_8016,N_8090);
nand U8546 (N_8546,N_8334,N_8343);
xor U8547 (N_8547,N_8048,N_8358);
and U8548 (N_8548,N_8292,N_8157);
xnor U8549 (N_8549,N_8324,N_8017);
and U8550 (N_8550,N_8180,N_8092);
or U8551 (N_8551,N_8312,N_8168);
or U8552 (N_8552,N_8061,N_8054);
xor U8553 (N_8553,N_8035,N_8219);
nor U8554 (N_8554,N_8291,N_8154);
nor U8555 (N_8555,N_8371,N_8337);
or U8556 (N_8556,N_8215,N_8382);
and U8557 (N_8557,N_8131,N_8205);
xnor U8558 (N_8558,N_8012,N_8298);
xnor U8559 (N_8559,N_8127,N_8143);
xnor U8560 (N_8560,N_8028,N_8368);
or U8561 (N_8561,N_8225,N_8357);
or U8562 (N_8562,N_8303,N_8123);
nor U8563 (N_8563,N_8244,N_8178);
nand U8564 (N_8564,N_8076,N_8383);
nand U8565 (N_8565,N_8160,N_8029);
and U8566 (N_8566,N_8376,N_8019);
nand U8567 (N_8567,N_8027,N_8255);
xor U8568 (N_8568,N_8124,N_8346);
nand U8569 (N_8569,N_8326,N_8198);
xnor U8570 (N_8570,N_8237,N_8060);
xnor U8571 (N_8571,N_8140,N_8020);
or U8572 (N_8572,N_8332,N_8122);
and U8573 (N_8573,N_8323,N_8070);
and U8574 (N_8574,N_8214,N_8378);
nand U8575 (N_8575,N_8268,N_8235);
and U8576 (N_8576,N_8091,N_8234);
nor U8577 (N_8577,N_8064,N_8342);
nor U8578 (N_8578,N_8314,N_8021);
nor U8579 (N_8579,N_8373,N_8264);
xnor U8580 (N_8580,N_8349,N_8305);
or U8581 (N_8581,N_8080,N_8136);
and U8582 (N_8582,N_8363,N_8329);
nand U8583 (N_8583,N_8281,N_8365);
and U8584 (N_8584,N_8177,N_8022);
and U8585 (N_8585,N_8043,N_8384);
nand U8586 (N_8586,N_8300,N_8135);
nand U8587 (N_8587,N_8354,N_8372);
nor U8588 (N_8588,N_8347,N_8155);
xnor U8589 (N_8589,N_8049,N_8283);
xor U8590 (N_8590,N_8184,N_8274);
nand U8591 (N_8591,N_8344,N_8253);
and U8592 (N_8592,N_8065,N_8338);
xnor U8593 (N_8593,N_8201,N_8183);
xnor U8594 (N_8594,N_8173,N_8286);
and U8595 (N_8595,N_8282,N_8071);
and U8596 (N_8596,N_8221,N_8072);
nand U8597 (N_8597,N_8399,N_8304);
nand U8598 (N_8598,N_8351,N_8397);
nand U8599 (N_8599,N_8246,N_8075);
nor U8600 (N_8600,N_8126,N_8036);
and U8601 (N_8601,N_8205,N_8321);
xnor U8602 (N_8602,N_8127,N_8184);
and U8603 (N_8603,N_8168,N_8141);
xnor U8604 (N_8604,N_8384,N_8065);
xor U8605 (N_8605,N_8090,N_8374);
nor U8606 (N_8606,N_8244,N_8173);
xor U8607 (N_8607,N_8137,N_8173);
and U8608 (N_8608,N_8220,N_8213);
or U8609 (N_8609,N_8249,N_8281);
nand U8610 (N_8610,N_8048,N_8159);
xor U8611 (N_8611,N_8289,N_8106);
nor U8612 (N_8612,N_8131,N_8357);
nor U8613 (N_8613,N_8296,N_8069);
nor U8614 (N_8614,N_8125,N_8016);
or U8615 (N_8615,N_8026,N_8205);
xnor U8616 (N_8616,N_8112,N_8100);
and U8617 (N_8617,N_8197,N_8352);
and U8618 (N_8618,N_8347,N_8181);
nand U8619 (N_8619,N_8157,N_8184);
nand U8620 (N_8620,N_8242,N_8123);
xor U8621 (N_8621,N_8374,N_8020);
or U8622 (N_8622,N_8123,N_8192);
and U8623 (N_8623,N_8096,N_8354);
nor U8624 (N_8624,N_8067,N_8210);
and U8625 (N_8625,N_8167,N_8030);
nor U8626 (N_8626,N_8346,N_8147);
xnor U8627 (N_8627,N_8319,N_8155);
and U8628 (N_8628,N_8221,N_8215);
nor U8629 (N_8629,N_8090,N_8152);
nor U8630 (N_8630,N_8044,N_8087);
or U8631 (N_8631,N_8153,N_8276);
xor U8632 (N_8632,N_8391,N_8236);
nand U8633 (N_8633,N_8151,N_8385);
or U8634 (N_8634,N_8153,N_8110);
xnor U8635 (N_8635,N_8007,N_8198);
nor U8636 (N_8636,N_8250,N_8059);
and U8637 (N_8637,N_8031,N_8075);
or U8638 (N_8638,N_8320,N_8216);
or U8639 (N_8639,N_8166,N_8081);
or U8640 (N_8640,N_8340,N_8254);
nand U8641 (N_8641,N_8094,N_8281);
and U8642 (N_8642,N_8056,N_8055);
nand U8643 (N_8643,N_8237,N_8206);
nor U8644 (N_8644,N_8137,N_8398);
or U8645 (N_8645,N_8395,N_8071);
xnor U8646 (N_8646,N_8116,N_8236);
or U8647 (N_8647,N_8169,N_8119);
nor U8648 (N_8648,N_8236,N_8198);
xor U8649 (N_8649,N_8193,N_8159);
and U8650 (N_8650,N_8287,N_8335);
xnor U8651 (N_8651,N_8362,N_8058);
xor U8652 (N_8652,N_8395,N_8127);
nor U8653 (N_8653,N_8078,N_8395);
or U8654 (N_8654,N_8273,N_8166);
or U8655 (N_8655,N_8182,N_8074);
nor U8656 (N_8656,N_8245,N_8213);
or U8657 (N_8657,N_8301,N_8359);
or U8658 (N_8658,N_8168,N_8247);
xnor U8659 (N_8659,N_8309,N_8241);
and U8660 (N_8660,N_8303,N_8252);
or U8661 (N_8661,N_8072,N_8154);
xnor U8662 (N_8662,N_8022,N_8362);
nand U8663 (N_8663,N_8071,N_8294);
or U8664 (N_8664,N_8036,N_8115);
or U8665 (N_8665,N_8150,N_8274);
or U8666 (N_8666,N_8231,N_8001);
and U8667 (N_8667,N_8268,N_8126);
nand U8668 (N_8668,N_8107,N_8360);
xor U8669 (N_8669,N_8067,N_8125);
nand U8670 (N_8670,N_8399,N_8217);
or U8671 (N_8671,N_8101,N_8249);
nand U8672 (N_8672,N_8100,N_8252);
or U8673 (N_8673,N_8023,N_8374);
or U8674 (N_8674,N_8081,N_8310);
and U8675 (N_8675,N_8252,N_8059);
and U8676 (N_8676,N_8201,N_8310);
and U8677 (N_8677,N_8013,N_8224);
nor U8678 (N_8678,N_8163,N_8291);
and U8679 (N_8679,N_8116,N_8364);
and U8680 (N_8680,N_8014,N_8009);
nand U8681 (N_8681,N_8031,N_8357);
and U8682 (N_8682,N_8147,N_8041);
and U8683 (N_8683,N_8218,N_8351);
xor U8684 (N_8684,N_8365,N_8187);
nor U8685 (N_8685,N_8115,N_8254);
nor U8686 (N_8686,N_8195,N_8151);
nand U8687 (N_8687,N_8027,N_8016);
xnor U8688 (N_8688,N_8364,N_8183);
nor U8689 (N_8689,N_8148,N_8289);
and U8690 (N_8690,N_8392,N_8061);
nor U8691 (N_8691,N_8058,N_8109);
nor U8692 (N_8692,N_8261,N_8123);
xnor U8693 (N_8693,N_8277,N_8148);
xor U8694 (N_8694,N_8019,N_8319);
xnor U8695 (N_8695,N_8289,N_8183);
and U8696 (N_8696,N_8316,N_8198);
nand U8697 (N_8697,N_8267,N_8110);
or U8698 (N_8698,N_8187,N_8033);
nand U8699 (N_8699,N_8008,N_8102);
nor U8700 (N_8700,N_8389,N_8304);
xor U8701 (N_8701,N_8338,N_8329);
nand U8702 (N_8702,N_8184,N_8052);
nand U8703 (N_8703,N_8031,N_8252);
nand U8704 (N_8704,N_8062,N_8344);
nor U8705 (N_8705,N_8375,N_8072);
or U8706 (N_8706,N_8198,N_8330);
nand U8707 (N_8707,N_8371,N_8285);
xor U8708 (N_8708,N_8222,N_8271);
or U8709 (N_8709,N_8276,N_8164);
and U8710 (N_8710,N_8066,N_8215);
and U8711 (N_8711,N_8396,N_8377);
or U8712 (N_8712,N_8281,N_8357);
nand U8713 (N_8713,N_8119,N_8393);
xnor U8714 (N_8714,N_8067,N_8050);
and U8715 (N_8715,N_8206,N_8129);
nor U8716 (N_8716,N_8277,N_8006);
or U8717 (N_8717,N_8148,N_8184);
or U8718 (N_8718,N_8345,N_8399);
xnor U8719 (N_8719,N_8025,N_8185);
xor U8720 (N_8720,N_8324,N_8059);
xor U8721 (N_8721,N_8224,N_8003);
and U8722 (N_8722,N_8223,N_8315);
and U8723 (N_8723,N_8150,N_8197);
and U8724 (N_8724,N_8153,N_8313);
nand U8725 (N_8725,N_8015,N_8215);
xnor U8726 (N_8726,N_8042,N_8143);
nor U8727 (N_8727,N_8310,N_8238);
xnor U8728 (N_8728,N_8255,N_8005);
or U8729 (N_8729,N_8248,N_8395);
and U8730 (N_8730,N_8304,N_8018);
or U8731 (N_8731,N_8120,N_8197);
or U8732 (N_8732,N_8381,N_8107);
or U8733 (N_8733,N_8001,N_8165);
nor U8734 (N_8734,N_8044,N_8162);
or U8735 (N_8735,N_8262,N_8110);
nand U8736 (N_8736,N_8138,N_8310);
xnor U8737 (N_8737,N_8097,N_8109);
and U8738 (N_8738,N_8193,N_8208);
or U8739 (N_8739,N_8240,N_8060);
xor U8740 (N_8740,N_8064,N_8263);
nor U8741 (N_8741,N_8002,N_8104);
xor U8742 (N_8742,N_8235,N_8052);
or U8743 (N_8743,N_8349,N_8049);
nor U8744 (N_8744,N_8302,N_8090);
nand U8745 (N_8745,N_8294,N_8087);
nor U8746 (N_8746,N_8294,N_8194);
nand U8747 (N_8747,N_8186,N_8143);
nand U8748 (N_8748,N_8347,N_8033);
and U8749 (N_8749,N_8076,N_8104);
nand U8750 (N_8750,N_8197,N_8161);
and U8751 (N_8751,N_8350,N_8008);
and U8752 (N_8752,N_8207,N_8075);
nor U8753 (N_8753,N_8390,N_8155);
xor U8754 (N_8754,N_8132,N_8250);
nand U8755 (N_8755,N_8389,N_8118);
nor U8756 (N_8756,N_8313,N_8102);
xor U8757 (N_8757,N_8323,N_8047);
xnor U8758 (N_8758,N_8270,N_8346);
and U8759 (N_8759,N_8175,N_8110);
and U8760 (N_8760,N_8017,N_8354);
nor U8761 (N_8761,N_8360,N_8281);
nand U8762 (N_8762,N_8034,N_8332);
or U8763 (N_8763,N_8263,N_8189);
nor U8764 (N_8764,N_8020,N_8158);
nand U8765 (N_8765,N_8305,N_8200);
nand U8766 (N_8766,N_8054,N_8306);
xnor U8767 (N_8767,N_8129,N_8393);
nand U8768 (N_8768,N_8054,N_8272);
xnor U8769 (N_8769,N_8224,N_8316);
nor U8770 (N_8770,N_8352,N_8150);
or U8771 (N_8771,N_8297,N_8204);
or U8772 (N_8772,N_8309,N_8078);
nor U8773 (N_8773,N_8370,N_8202);
or U8774 (N_8774,N_8322,N_8177);
and U8775 (N_8775,N_8387,N_8120);
nand U8776 (N_8776,N_8180,N_8229);
nor U8777 (N_8777,N_8381,N_8114);
nand U8778 (N_8778,N_8143,N_8135);
nor U8779 (N_8779,N_8166,N_8268);
xnor U8780 (N_8780,N_8093,N_8319);
and U8781 (N_8781,N_8307,N_8336);
or U8782 (N_8782,N_8199,N_8035);
nand U8783 (N_8783,N_8161,N_8196);
and U8784 (N_8784,N_8331,N_8146);
nand U8785 (N_8785,N_8034,N_8064);
and U8786 (N_8786,N_8128,N_8055);
nor U8787 (N_8787,N_8366,N_8029);
nand U8788 (N_8788,N_8226,N_8138);
nor U8789 (N_8789,N_8156,N_8334);
nand U8790 (N_8790,N_8026,N_8080);
xor U8791 (N_8791,N_8159,N_8060);
xnor U8792 (N_8792,N_8389,N_8105);
or U8793 (N_8793,N_8167,N_8256);
nor U8794 (N_8794,N_8031,N_8239);
nand U8795 (N_8795,N_8221,N_8087);
xnor U8796 (N_8796,N_8149,N_8391);
xor U8797 (N_8797,N_8063,N_8056);
and U8798 (N_8798,N_8286,N_8222);
and U8799 (N_8799,N_8041,N_8083);
and U8800 (N_8800,N_8487,N_8541);
or U8801 (N_8801,N_8721,N_8714);
xor U8802 (N_8802,N_8430,N_8418);
and U8803 (N_8803,N_8789,N_8411);
xor U8804 (N_8804,N_8703,N_8445);
nor U8805 (N_8805,N_8507,N_8694);
xnor U8806 (N_8806,N_8631,N_8691);
nor U8807 (N_8807,N_8601,N_8655);
nor U8808 (N_8808,N_8427,N_8738);
nand U8809 (N_8809,N_8612,N_8596);
or U8810 (N_8810,N_8491,N_8540);
xor U8811 (N_8811,N_8471,N_8556);
or U8812 (N_8812,N_8737,N_8422);
xor U8813 (N_8813,N_8599,N_8457);
nand U8814 (N_8814,N_8744,N_8643);
nor U8815 (N_8815,N_8695,N_8454);
nand U8816 (N_8816,N_8433,N_8573);
nand U8817 (N_8817,N_8465,N_8787);
nor U8818 (N_8818,N_8494,N_8632);
or U8819 (N_8819,N_8630,N_8505);
nor U8820 (N_8820,N_8482,N_8758);
nand U8821 (N_8821,N_8486,N_8438);
xor U8822 (N_8822,N_8656,N_8460);
nand U8823 (N_8823,N_8652,N_8543);
and U8824 (N_8824,N_8553,N_8773);
nor U8825 (N_8825,N_8751,N_8407);
or U8826 (N_8826,N_8716,N_8653);
nand U8827 (N_8827,N_8511,N_8493);
or U8828 (N_8828,N_8761,N_8475);
nand U8829 (N_8829,N_8429,N_8664);
and U8830 (N_8830,N_8587,N_8712);
xor U8831 (N_8831,N_8565,N_8734);
or U8832 (N_8832,N_8724,N_8709);
nor U8833 (N_8833,N_8776,N_8500);
xnor U8834 (N_8834,N_8674,N_8795);
nor U8835 (N_8835,N_8688,N_8544);
nor U8836 (N_8836,N_8727,N_8686);
xnor U8837 (N_8837,N_8506,N_8641);
and U8838 (N_8838,N_8786,N_8424);
or U8839 (N_8839,N_8697,N_8548);
and U8840 (N_8840,N_8481,N_8654);
or U8841 (N_8841,N_8708,N_8651);
nand U8842 (N_8842,N_8463,N_8749);
and U8843 (N_8843,N_8676,N_8538);
xnor U8844 (N_8844,N_8512,N_8437);
and U8845 (N_8845,N_8770,N_8650);
nor U8846 (N_8846,N_8701,N_8495);
nand U8847 (N_8847,N_8555,N_8683);
and U8848 (N_8848,N_8742,N_8559);
nand U8849 (N_8849,N_8527,N_8530);
nor U8850 (N_8850,N_8696,N_8747);
or U8851 (N_8851,N_8525,N_8726);
xor U8852 (N_8852,N_8444,N_8689);
xnor U8853 (N_8853,N_8693,N_8771);
and U8854 (N_8854,N_8769,N_8488);
nand U8855 (N_8855,N_8649,N_8534);
nand U8856 (N_8856,N_8748,N_8627);
and U8857 (N_8857,N_8637,N_8588);
nand U8858 (N_8858,N_8598,N_8575);
nor U8859 (N_8859,N_8774,N_8797);
xnor U8860 (N_8860,N_8469,N_8467);
xnor U8861 (N_8861,N_8752,N_8662);
xnor U8862 (N_8862,N_8754,N_8432);
xor U8863 (N_8863,N_8459,N_8410);
xor U8864 (N_8864,N_8403,N_8767);
nand U8865 (N_8865,N_8621,N_8515);
nor U8866 (N_8866,N_8570,N_8642);
xor U8867 (N_8867,N_8720,N_8574);
nor U8868 (N_8868,N_8765,N_8585);
xnor U8869 (N_8869,N_8472,N_8740);
and U8870 (N_8870,N_8762,N_8669);
or U8871 (N_8871,N_8455,N_8619);
xor U8872 (N_8872,N_8743,N_8453);
xor U8873 (N_8873,N_8713,N_8434);
nor U8874 (N_8874,N_8690,N_8443);
nor U8875 (N_8875,N_8466,N_8450);
and U8876 (N_8876,N_8673,N_8778);
xor U8877 (N_8877,N_8780,N_8536);
xnor U8878 (N_8878,N_8668,N_8796);
and U8879 (N_8879,N_8603,N_8503);
nand U8880 (N_8880,N_8685,N_8519);
nor U8881 (N_8881,N_8783,N_8745);
and U8882 (N_8882,N_8799,N_8497);
xor U8883 (N_8883,N_8633,N_8647);
and U8884 (N_8884,N_8766,N_8618);
and U8885 (N_8885,N_8564,N_8682);
nor U8886 (N_8886,N_8730,N_8733);
xnor U8887 (N_8887,N_8479,N_8584);
or U8888 (N_8888,N_8666,N_8567);
xnor U8889 (N_8889,N_8547,N_8772);
nand U8890 (N_8890,N_8794,N_8554);
nor U8891 (N_8891,N_8680,N_8725);
nand U8892 (N_8892,N_8423,N_8592);
nor U8893 (N_8893,N_8529,N_8705);
and U8894 (N_8894,N_8657,N_8417);
nor U8895 (N_8895,N_8626,N_8638);
and U8896 (N_8896,N_8611,N_8617);
xnor U8897 (N_8897,N_8792,N_8613);
and U8898 (N_8898,N_8739,N_8604);
or U8899 (N_8899,N_8510,N_8428);
nor U8900 (N_8900,N_8722,N_8615);
and U8901 (N_8901,N_8715,N_8404);
nand U8902 (N_8902,N_8760,N_8671);
or U8903 (N_8903,N_8485,N_8741);
nor U8904 (N_8904,N_8777,N_8661);
nor U8905 (N_8905,N_8711,N_8750);
and U8906 (N_8906,N_8546,N_8706);
nand U8907 (N_8907,N_8470,N_8723);
nor U8908 (N_8908,N_8535,N_8415);
nand U8909 (N_8909,N_8610,N_8436);
and U8910 (N_8910,N_8489,N_8595);
or U8911 (N_8911,N_8421,N_8710);
or U8912 (N_8912,N_8520,N_8717);
and U8913 (N_8913,N_8622,N_8679);
nand U8914 (N_8914,N_8677,N_8458);
nand U8915 (N_8915,N_8502,N_8764);
and U8916 (N_8916,N_8707,N_8522);
nor U8917 (N_8917,N_8498,N_8670);
nor U8918 (N_8918,N_8521,N_8464);
xnor U8919 (N_8919,N_8583,N_8678);
nor U8920 (N_8920,N_8692,N_8524);
xnor U8921 (N_8921,N_8605,N_8478);
nand U8922 (N_8922,N_8542,N_8798);
nor U8923 (N_8923,N_8667,N_8589);
and U8924 (N_8924,N_8514,N_8784);
and U8925 (N_8925,N_8768,N_8609);
nand U8926 (N_8926,N_8518,N_8474);
xor U8927 (N_8927,N_8704,N_8698);
and U8928 (N_8928,N_8572,N_8577);
nand U8929 (N_8929,N_8462,N_8606);
nand U8930 (N_8930,N_8757,N_8639);
or U8931 (N_8931,N_8513,N_8468);
or U8932 (N_8932,N_8408,N_8528);
or U8933 (N_8933,N_8702,N_8425);
and U8934 (N_8934,N_8431,N_8590);
nand U8935 (N_8935,N_8586,N_8456);
nor U8936 (N_8936,N_8480,N_8728);
nand U8937 (N_8937,N_8793,N_8569);
xor U8938 (N_8938,N_8508,N_8791);
or U8939 (N_8939,N_8483,N_8719);
or U8940 (N_8940,N_8620,N_8628);
and U8941 (N_8941,N_8675,N_8729);
xnor U8942 (N_8942,N_8501,N_8517);
xnor U8943 (N_8943,N_8412,N_8687);
nor U8944 (N_8944,N_8681,N_8400);
xnor U8945 (N_8945,N_8645,N_8602);
and U8946 (N_8946,N_8779,N_8623);
or U8947 (N_8947,N_8549,N_8732);
nor U8948 (N_8948,N_8420,N_8452);
nand U8949 (N_8949,N_8477,N_8413);
and U8950 (N_8950,N_8532,N_8447);
or U8951 (N_8951,N_8646,N_8545);
nor U8952 (N_8952,N_8516,N_8579);
or U8953 (N_8953,N_8755,N_8539);
and U8954 (N_8954,N_8523,N_8594);
nand U8955 (N_8955,N_8663,N_8552);
or U8956 (N_8956,N_8785,N_8442);
xor U8957 (N_8957,N_8492,N_8736);
nand U8958 (N_8958,N_8635,N_8566);
nand U8959 (N_8959,N_8665,N_8608);
or U8960 (N_8960,N_8616,N_8557);
and U8961 (N_8961,N_8473,N_8581);
nor U8962 (N_8962,N_8775,N_8526);
nor U8963 (N_8963,N_8568,N_8644);
xor U8964 (N_8964,N_8405,N_8699);
or U8965 (N_8965,N_8561,N_8614);
or U8966 (N_8966,N_8537,N_8781);
and U8967 (N_8967,N_8461,N_8658);
nand U8968 (N_8968,N_8441,N_8648);
nor U8969 (N_8969,N_8640,N_8563);
nand U8970 (N_8970,N_8731,N_8440);
and U8971 (N_8971,N_8735,N_8439);
nand U8972 (N_8972,N_8782,N_8684);
nand U8973 (N_8973,N_8582,N_8788);
nand U8974 (N_8974,N_8660,N_8558);
and U8975 (N_8975,N_8490,N_8448);
and U8976 (N_8976,N_8591,N_8504);
nor U8977 (N_8977,N_8578,N_8629);
and U8978 (N_8978,N_8746,N_8419);
or U8979 (N_8979,N_8634,N_8756);
or U8980 (N_8980,N_8509,N_8401);
xnor U8981 (N_8981,N_8484,N_8659);
nor U8982 (N_8982,N_8550,N_8759);
and U8983 (N_8983,N_8426,N_8718);
nand U8984 (N_8984,N_8672,N_8551);
and U8985 (N_8985,N_8753,N_8790);
nand U8986 (N_8986,N_8763,N_8597);
or U8987 (N_8987,N_8446,N_8449);
and U8988 (N_8988,N_8414,N_8562);
and U8989 (N_8989,N_8451,N_8533);
or U8990 (N_8990,N_8531,N_8593);
and U8991 (N_8991,N_8625,N_8576);
nand U8992 (N_8992,N_8406,N_8624);
or U8993 (N_8993,N_8435,N_8600);
or U8994 (N_8994,N_8409,N_8560);
nand U8995 (N_8995,N_8580,N_8416);
xnor U8996 (N_8996,N_8700,N_8402);
and U8997 (N_8997,N_8607,N_8571);
and U8998 (N_8998,N_8476,N_8496);
and U8999 (N_8999,N_8499,N_8636);
or U9000 (N_9000,N_8541,N_8562);
nand U9001 (N_9001,N_8524,N_8603);
nand U9002 (N_9002,N_8728,N_8635);
nand U9003 (N_9003,N_8491,N_8722);
or U9004 (N_9004,N_8402,N_8546);
nor U9005 (N_9005,N_8686,N_8420);
nand U9006 (N_9006,N_8748,N_8562);
and U9007 (N_9007,N_8483,N_8739);
or U9008 (N_9008,N_8434,N_8406);
and U9009 (N_9009,N_8652,N_8709);
and U9010 (N_9010,N_8634,N_8433);
nand U9011 (N_9011,N_8562,N_8799);
and U9012 (N_9012,N_8402,N_8690);
nor U9013 (N_9013,N_8657,N_8568);
or U9014 (N_9014,N_8787,N_8495);
nor U9015 (N_9015,N_8744,N_8716);
or U9016 (N_9016,N_8559,N_8713);
nor U9017 (N_9017,N_8655,N_8536);
nor U9018 (N_9018,N_8645,N_8573);
xor U9019 (N_9019,N_8502,N_8497);
or U9020 (N_9020,N_8568,N_8546);
nor U9021 (N_9021,N_8471,N_8734);
or U9022 (N_9022,N_8492,N_8488);
or U9023 (N_9023,N_8788,N_8518);
xor U9024 (N_9024,N_8579,N_8475);
or U9025 (N_9025,N_8566,N_8767);
and U9026 (N_9026,N_8541,N_8555);
and U9027 (N_9027,N_8500,N_8629);
nand U9028 (N_9028,N_8640,N_8527);
nor U9029 (N_9029,N_8556,N_8500);
xor U9030 (N_9030,N_8660,N_8533);
xor U9031 (N_9031,N_8688,N_8627);
xor U9032 (N_9032,N_8412,N_8606);
xor U9033 (N_9033,N_8744,N_8519);
xnor U9034 (N_9034,N_8627,N_8484);
or U9035 (N_9035,N_8631,N_8773);
or U9036 (N_9036,N_8731,N_8794);
nor U9037 (N_9037,N_8626,N_8432);
and U9038 (N_9038,N_8721,N_8677);
xnor U9039 (N_9039,N_8521,N_8646);
or U9040 (N_9040,N_8412,N_8796);
and U9041 (N_9041,N_8714,N_8483);
or U9042 (N_9042,N_8707,N_8495);
and U9043 (N_9043,N_8773,N_8723);
and U9044 (N_9044,N_8745,N_8517);
nand U9045 (N_9045,N_8717,N_8672);
xor U9046 (N_9046,N_8512,N_8651);
nand U9047 (N_9047,N_8762,N_8779);
and U9048 (N_9048,N_8494,N_8653);
nor U9049 (N_9049,N_8569,N_8670);
or U9050 (N_9050,N_8779,N_8780);
nand U9051 (N_9051,N_8528,N_8704);
xor U9052 (N_9052,N_8792,N_8438);
xnor U9053 (N_9053,N_8748,N_8504);
and U9054 (N_9054,N_8713,N_8699);
nor U9055 (N_9055,N_8498,N_8468);
or U9056 (N_9056,N_8732,N_8601);
and U9057 (N_9057,N_8585,N_8561);
and U9058 (N_9058,N_8494,N_8658);
and U9059 (N_9059,N_8549,N_8413);
or U9060 (N_9060,N_8680,N_8705);
nor U9061 (N_9061,N_8689,N_8699);
and U9062 (N_9062,N_8404,N_8488);
or U9063 (N_9063,N_8712,N_8678);
xnor U9064 (N_9064,N_8559,N_8577);
nor U9065 (N_9065,N_8744,N_8611);
nand U9066 (N_9066,N_8631,N_8732);
nand U9067 (N_9067,N_8476,N_8536);
xnor U9068 (N_9068,N_8427,N_8701);
and U9069 (N_9069,N_8624,N_8647);
and U9070 (N_9070,N_8584,N_8750);
nand U9071 (N_9071,N_8657,N_8495);
xor U9072 (N_9072,N_8589,N_8742);
nor U9073 (N_9073,N_8753,N_8500);
nand U9074 (N_9074,N_8538,N_8686);
nand U9075 (N_9075,N_8427,N_8545);
nand U9076 (N_9076,N_8584,N_8570);
xor U9077 (N_9077,N_8648,N_8477);
or U9078 (N_9078,N_8618,N_8508);
nor U9079 (N_9079,N_8787,N_8714);
or U9080 (N_9080,N_8483,N_8741);
and U9081 (N_9081,N_8763,N_8682);
nand U9082 (N_9082,N_8710,N_8664);
nand U9083 (N_9083,N_8613,N_8489);
or U9084 (N_9084,N_8595,N_8583);
nand U9085 (N_9085,N_8695,N_8662);
nor U9086 (N_9086,N_8762,N_8443);
nand U9087 (N_9087,N_8646,N_8683);
or U9088 (N_9088,N_8731,N_8721);
and U9089 (N_9089,N_8797,N_8563);
nand U9090 (N_9090,N_8494,N_8624);
or U9091 (N_9091,N_8697,N_8707);
and U9092 (N_9092,N_8411,N_8424);
nor U9093 (N_9093,N_8651,N_8752);
xor U9094 (N_9094,N_8597,N_8404);
nand U9095 (N_9095,N_8564,N_8593);
xor U9096 (N_9096,N_8769,N_8700);
nand U9097 (N_9097,N_8426,N_8703);
nor U9098 (N_9098,N_8645,N_8686);
nand U9099 (N_9099,N_8671,N_8799);
xnor U9100 (N_9100,N_8605,N_8741);
nand U9101 (N_9101,N_8543,N_8720);
nor U9102 (N_9102,N_8692,N_8447);
nor U9103 (N_9103,N_8694,N_8453);
xor U9104 (N_9104,N_8610,N_8600);
xor U9105 (N_9105,N_8736,N_8742);
and U9106 (N_9106,N_8525,N_8596);
and U9107 (N_9107,N_8786,N_8661);
or U9108 (N_9108,N_8500,N_8559);
and U9109 (N_9109,N_8482,N_8743);
nor U9110 (N_9110,N_8790,N_8613);
or U9111 (N_9111,N_8433,N_8540);
and U9112 (N_9112,N_8431,N_8682);
xnor U9113 (N_9113,N_8714,N_8570);
nand U9114 (N_9114,N_8567,N_8737);
or U9115 (N_9115,N_8579,N_8431);
or U9116 (N_9116,N_8539,N_8641);
nand U9117 (N_9117,N_8557,N_8483);
xnor U9118 (N_9118,N_8539,N_8723);
nor U9119 (N_9119,N_8782,N_8586);
xor U9120 (N_9120,N_8759,N_8680);
and U9121 (N_9121,N_8485,N_8555);
xor U9122 (N_9122,N_8745,N_8742);
xnor U9123 (N_9123,N_8500,N_8671);
and U9124 (N_9124,N_8695,N_8573);
xor U9125 (N_9125,N_8722,N_8567);
xnor U9126 (N_9126,N_8783,N_8708);
or U9127 (N_9127,N_8491,N_8588);
and U9128 (N_9128,N_8495,N_8795);
nand U9129 (N_9129,N_8589,N_8455);
nand U9130 (N_9130,N_8400,N_8796);
xnor U9131 (N_9131,N_8560,N_8685);
nand U9132 (N_9132,N_8425,N_8514);
nor U9133 (N_9133,N_8701,N_8577);
nor U9134 (N_9134,N_8528,N_8701);
or U9135 (N_9135,N_8730,N_8644);
nor U9136 (N_9136,N_8796,N_8409);
nand U9137 (N_9137,N_8561,N_8401);
nor U9138 (N_9138,N_8407,N_8588);
xnor U9139 (N_9139,N_8412,N_8584);
nor U9140 (N_9140,N_8748,N_8630);
nor U9141 (N_9141,N_8595,N_8764);
xor U9142 (N_9142,N_8784,N_8777);
xor U9143 (N_9143,N_8711,N_8620);
or U9144 (N_9144,N_8652,N_8573);
or U9145 (N_9145,N_8676,N_8655);
nand U9146 (N_9146,N_8693,N_8630);
nand U9147 (N_9147,N_8574,N_8462);
or U9148 (N_9148,N_8591,N_8697);
nand U9149 (N_9149,N_8573,N_8608);
and U9150 (N_9150,N_8638,N_8546);
and U9151 (N_9151,N_8610,N_8761);
or U9152 (N_9152,N_8543,N_8439);
xnor U9153 (N_9153,N_8583,N_8452);
nor U9154 (N_9154,N_8441,N_8617);
or U9155 (N_9155,N_8530,N_8628);
xnor U9156 (N_9156,N_8441,N_8574);
xnor U9157 (N_9157,N_8593,N_8584);
xor U9158 (N_9158,N_8438,N_8436);
or U9159 (N_9159,N_8522,N_8748);
or U9160 (N_9160,N_8587,N_8505);
xnor U9161 (N_9161,N_8785,N_8416);
and U9162 (N_9162,N_8468,N_8742);
nor U9163 (N_9163,N_8442,N_8497);
nand U9164 (N_9164,N_8510,N_8571);
nor U9165 (N_9165,N_8746,N_8548);
and U9166 (N_9166,N_8759,N_8489);
or U9167 (N_9167,N_8465,N_8558);
nand U9168 (N_9168,N_8680,N_8638);
nor U9169 (N_9169,N_8579,N_8778);
nor U9170 (N_9170,N_8619,N_8425);
xnor U9171 (N_9171,N_8692,N_8740);
nor U9172 (N_9172,N_8489,N_8537);
nor U9173 (N_9173,N_8722,N_8695);
and U9174 (N_9174,N_8587,N_8458);
or U9175 (N_9175,N_8774,N_8715);
and U9176 (N_9176,N_8644,N_8776);
or U9177 (N_9177,N_8626,N_8523);
xnor U9178 (N_9178,N_8701,N_8659);
or U9179 (N_9179,N_8485,N_8758);
or U9180 (N_9180,N_8524,N_8728);
or U9181 (N_9181,N_8713,N_8656);
nand U9182 (N_9182,N_8756,N_8503);
xor U9183 (N_9183,N_8557,N_8506);
and U9184 (N_9184,N_8495,N_8736);
nand U9185 (N_9185,N_8472,N_8465);
and U9186 (N_9186,N_8422,N_8558);
xor U9187 (N_9187,N_8425,N_8438);
nand U9188 (N_9188,N_8766,N_8524);
or U9189 (N_9189,N_8655,N_8618);
xnor U9190 (N_9190,N_8600,N_8573);
nand U9191 (N_9191,N_8522,N_8479);
or U9192 (N_9192,N_8731,N_8468);
xor U9193 (N_9193,N_8671,N_8548);
and U9194 (N_9194,N_8610,N_8680);
nor U9195 (N_9195,N_8504,N_8609);
nand U9196 (N_9196,N_8725,N_8709);
or U9197 (N_9197,N_8483,N_8733);
nand U9198 (N_9198,N_8700,N_8709);
xnor U9199 (N_9199,N_8669,N_8721);
xor U9200 (N_9200,N_8831,N_8855);
xnor U9201 (N_9201,N_8949,N_9105);
or U9202 (N_9202,N_8951,N_9006);
xnor U9203 (N_9203,N_8812,N_8948);
xor U9204 (N_9204,N_9109,N_8870);
and U9205 (N_9205,N_8956,N_9051);
nor U9206 (N_9206,N_8924,N_9155);
nor U9207 (N_9207,N_8844,N_8909);
xor U9208 (N_9208,N_8832,N_8964);
nor U9209 (N_9209,N_9003,N_8874);
nand U9210 (N_9210,N_9094,N_9123);
nand U9211 (N_9211,N_9016,N_9026);
and U9212 (N_9212,N_9045,N_8997);
xnor U9213 (N_9213,N_8973,N_9062);
nand U9214 (N_9214,N_8989,N_8980);
nor U9215 (N_9215,N_9092,N_8972);
nand U9216 (N_9216,N_8925,N_8915);
nand U9217 (N_9217,N_9139,N_8817);
xor U9218 (N_9218,N_9135,N_9112);
nand U9219 (N_9219,N_9015,N_8933);
or U9220 (N_9220,N_8963,N_9127);
nand U9221 (N_9221,N_9028,N_9195);
nor U9222 (N_9222,N_9038,N_8828);
and U9223 (N_9223,N_9115,N_9029);
and U9224 (N_9224,N_9057,N_8861);
or U9225 (N_9225,N_8939,N_8994);
or U9226 (N_9226,N_8877,N_8969);
and U9227 (N_9227,N_8917,N_9149);
or U9228 (N_9228,N_9076,N_8928);
nand U9229 (N_9229,N_9193,N_9021);
xor U9230 (N_9230,N_9128,N_8913);
nor U9231 (N_9231,N_8875,N_8983);
nor U9232 (N_9232,N_8824,N_9072);
nand U9233 (N_9233,N_8955,N_9175);
or U9234 (N_9234,N_9039,N_8970);
nand U9235 (N_9235,N_9025,N_8962);
and U9236 (N_9236,N_9184,N_9060);
nand U9237 (N_9237,N_8981,N_9088);
and U9238 (N_9238,N_9185,N_8846);
xnor U9239 (N_9239,N_9106,N_8911);
nand U9240 (N_9240,N_8823,N_8853);
and U9241 (N_9241,N_8965,N_9120);
xor U9242 (N_9242,N_9170,N_8898);
nand U9243 (N_9243,N_9192,N_9042);
nand U9244 (N_9244,N_8820,N_9138);
nand U9245 (N_9245,N_9001,N_8941);
or U9246 (N_9246,N_9156,N_9098);
or U9247 (N_9247,N_9020,N_9083);
and U9248 (N_9248,N_8868,N_8872);
xnor U9249 (N_9249,N_8991,N_8860);
nor U9250 (N_9250,N_8910,N_8967);
xnor U9251 (N_9251,N_8954,N_9052);
xor U9252 (N_9252,N_8947,N_9125);
and U9253 (N_9253,N_8809,N_8976);
nand U9254 (N_9254,N_8998,N_8923);
and U9255 (N_9255,N_9054,N_8838);
or U9256 (N_9256,N_9085,N_9172);
nand U9257 (N_9257,N_8805,N_8810);
xor U9258 (N_9258,N_8887,N_8827);
nor U9259 (N_9259,N_9103,N_9101);
and U9260 (N_9260,N_9007,N_9143);
nand U9261 (N_9261,N_8834,N_9080);
nor U9262 (N_9262,N_8800,N_8918);
and U9263 (N_9263,N_8878,N_9093);
or U9264 (N_9264,N_8978,N_9087);
nor U9265 (N_9265,N_8806,N_9187);
xnor U9266 (N_9266,N_9102,N_8904);
or U9267 (N_9267,N_9089,N_8808);
and U9268 (N_9268,N_8858,N_8865);
nor U9269 (N_9269,N_9043,N_9009);
and U9270 (N_9270,N_8847,N_9037);
xor U9271 (N_9271,N_9152,N_9142);
and U9272 (N_9272,N_8840,N_9074);
xnor U9273 (N_9273,N_8942,N_8854);
nand U9274 (N_9274,N_9095,N_8891);
nor U9275 (N_9275,N_9111,N_8999);
and U9276 (N_9276,N_8859,N_8835);
and U9277 (N_9277,N_9034,N_8852);
and U9278 (N_9278,N_9131,N_9108);
and U9279 (N_9279,N_8903,N_9058);
nand U9280 (N_9280,N_8818,N_9130);
or U9281 (N_9281,N_9117,N_8975);
nor U9282 (N_9282,N_9032,N_8958);
or U9283 (N_9283,N_8902,N_8934);
nor U9284 (N_9284,N_9159,N_8930);
nor U9285 (N_9285,N_9040,N_8968);
or U9286 (N_9286,N_8936,N_8931);
and U9287 (N_9287,N_9121,N_9066);
and U9288 (N_9288,N_9119,N_8908);
nor U9289 (N_9289,N_8966,N_9000);
or U9290 (N_9290,N_9049,N_9011);
nor U9291 (N_9291,N_8961,N_9146);
or U9292 (N_9292,N_8927,N_8890);
or U9293 (N_9293,N_8893,N_9008);
or U9294 (N_9294,N_8979,N_8984);
xor U9295 (N_9295,N_9036,N_8883);
or U9296 (N_9296,N_9012,N_9134);
and U9297 (N_9297,N_8863,N_9077);
and U9298 (N_9298,N_9166,N_8862);
xnor U9299 (N_9299,N_9019,N_8839);
and U9300 (N_9300,N_9024,N_9099);
and U9301 (N_9301,N_9078,N_9091);
xnor U9302 (N_9302,N_8802,N_9100);
nand U9303 (N_9303,N_8953,N_9071);
nor U9304 (N_9304,N_8914,N_8825);
nor U9305 (N_9305,N_8906,N_8905);
xor U9306 (N_9306,N_9129,N_8900);
and U9307 (N_9307,N_8945,N_9182);
and U9308 (N_9308,N_8952,N_8922);
xor U9309 (N_9309,N_8850,N_9122);
nand U9310 (N_9310,N_9190,N_8921);
and U9311 (N_9311,N_9061,N_9153);
or U9312 (N_9312,N_8841,N_9053);
and U9313 (N_9313,N_8957,N_8990);
and U9314 (N_9314,N_8932,N_9158);
nor U9315 (N_9315,N_9047,N_8851);
or U9316 (N_9316,N_8982,N_9169);
xnor U9317 (N_9317,N_9194,N_8822);
nand U9318 (N_9318,N_9014,N_8833);
xor U9319 (N_9319,N_8896,N_8811);
nand U9320 (N_9320,N_9110,N_8889);
xor U9321 (N_9321,N_8842,N_8880);
and U9322 (N_9322,N_8804,N_8988);
nor U9323 (N_9323,N_9116,N_9018);
nor U9324 (N_9324,N_9147,N_8819);
nand U9325 (N_9325,N_8849,N_8894);
and U9326 (N_9326,N_9073,N_8926);
nand U9327 (N_9327,N_8971,N_8879);
nand U9328 (N_9328,N_8960,N_9160);
nor U9329 (N_9329,N_8814,N_9017);
nand U9330 (N_9330,N_9183,N_9148);
and U9331 (N_9331,N_8946,N_9005);
nand U9332 (N_9332,N_9151,N_8876);
nand U9333 (N_9333,N_8993,N_8867);
and U9334 (N_9334,N_9030,N_9197);
nand U9335 (N_9335,N_8995,N_8856);
xnor U9336 (N_9336,N_9086,N_8829);
and U9337 (N_9337,N_8845,N_8886);
and U9338 (N_9338,N_8974,N_9140);
xor U9339 (N_9339,N_9023,N_8897);
or U9340 (N_9340,N_9199,N_9136);
nand U9341 (N_9341,N_9084,N_9150);
nand U9342 (N_9342,N_9164,N_8821);
xor U9343 (N_9343,N_9163,N_9055);
or U9344 (N_9344,N_8937,N_8884);
nand U9345 (N_9345,N_9165,N_9167);
and U9346 (N_9346,N_9079,N_8848);
xnor U9347 (N_9347,N_8996,N_9180);
xnor U9348 (N_9348,N_9046,N_9145);
nand U9349 (N_9349,N_8885,N_8959);
nand U9350 (N_9350,N_8944,N_8986);
xnor U9351 (N_9351,N_9107,N_9035);
nand U9352 (N_9352,N_9059,N_9104);
nand U9353 (N_9353,N_9067,N_9041);
or U9354 (N_9354,N_8977,N_8943);
or U9355 (N_9355,N_8830,N_9050);
or U9356 (N_9356,N_9022,N_9031);
or U9357 (N_9357,N_9177,N_9141);
nor U9358 (N_9358,N_9056,N_9157);
xor U9359 (N_9359,N_8919,N_9173);
xnor U9360 (N_9360,N_9162,N_9179);
nand U9361 (N_9361,N_9075,N_9081);
nand U9362 (N_9362,N_8907,N_8895);
nor U9363 (N_9363,N_9082,N_8837);
or U9364 (N_9364,N_8929,N_9033);
nand U9365 (N_9365,N_9013,N_9044);
and U9366 (N_9366,N_9070,N_9186);
nand U9367 (N_9367,N_8869,N_9198);
nand U9368 (N_9368,N_9181,N_8985);
xor U9369 (N_9369,N_9133,N_8888);
nand U9370 (N_9370,N_9027,N_9090);
or U9371 (N_9371,N_9063,N_8816);
nand U9372 (N_9372,N_8813,N_8866);
nand U9373 (N_9373,N_8912,N_8873);
nand U9374 (N_9374,N_8857,N_8935);
or U9375 (N_9375,N_8836,N_8843);
or U9376 (N_9376,N_8899,N_8864);
nor U9377 (N_9377,N_9002,N_9069);
nand U9378 (N_9378,N_9144,N_8992);
nor U9379 (N_9379,N_9176,N_9118);
nand U9380 (N_9380,N_9048,N_8950);
nor U9381 (N_9381,N_9137,N_8803);
or U9382 (N_9382,N_8987,N_9171);
xnor U9383 (N_9383,N_9196,N_8807);
and U9384 (N_9384,N_9126,N_8916);
nand U9385 (N_9385,N_8892,N_8826);
nor U9386 (N_9386,N_8940,N_9168);
or U9387 (N_9387,N_9191,N_9174);
xor U9388 (N_9388,N_8815,N_8871);
xor U9389 (N_9389,N_8882,N_8901);
and U9390 (N_9390,N_9132,N_9096);
nor U9391 (N_9391,N_9097,N_8920);
xor U9392 (N_9392,N_9124,N_8881);
and U9393 (N_9393,N_9065,N_8938);
and U9394 (N_9394,N_9064,N_9010);
xor U9395 (N_9395,N_9114,N_9154);
nand U9396 (N_9396,N_9068,N_9004);
and U9397 (N_9397,N_9189,N_8801);
or U9398 (N_9398,N_9161,N_9178);
and U9399 (N_9399,N_9113,N_9188);
or U9400 (N_9400,N_9023,N_8988);
xnor U9401 (N_9401,N_9135,N_9141);
and U9402 (N_9402,N_9045,N_9048);
nand U9403 (N_9403,N_9132,N_9008);
and U9404 (N_9404,N_9055,N_8917);
and U9405 (N_9405,N_8861,N_9194);
nand U9406 (N_9406,N_9033,N_9047);
xnor U9407 (N_9407,N_9164,N_8938);
nand U9408 (N_9408,N_9036,N_9177);
or U9409 (N_9409,N_8982,N_8930);
nor U9410 (N_9410,N_8935,N_9048);
or U9411 (N_9411,N_9021,N_9054);
nor U9412 (N_9412,N_9032,N_8851);
or U9413 (N_9413,N_8818,N_9080);
nand U9414 (N_9414,N_8978,N_9167);
and U9415 (N_9415,N_9056,N_8979);
or U9416 (N_9416,N_9145,N_9156);
or U9417 (N_9417,N_9177,N_8881);
nand U9418 (N_9418,N_8832,N_8881);
nand U9419 (N_9419,N_8912,N_9099);
and U9420 (N_9420,N_8851,N_9153);
or U9421 (N_9421,N_9147,N_8935);
xor U9422 (N_9422,N_8994,N_9154);
nand U9423 (N_9423,N_9137,N_9113);
xor U9424 (N_9424,N_9116,N_8867);
or U9425 (N_9425,N_9064,N_8985);
nor U9426 (N_9426,N_9037,N_8925);
or U9427 (N_9427,N_9041,N_9135);
nand U9428 (N_9428,N_9107,N_8922);
xor U9429 (N_9429,N_8831,N_9174);
or U9430 (N_9430,N_9022,N_8836);
or U9431 (N_9431,N_9030,N_9116);
nand U9432 (N_9432,N_8946,N_8902);
nor U9433 (N_9433,N_8987,N_9134);
and U9434 (N_9434,N_8857,N_8869);
and U9435 (N_9435,N_8879,N_8900);
or U9436 (N_9436,N_9084,N_9195);
xnor U9437 (N_9437,N_9155,N_9048);
or U9438 (N_9438,N_8916,N_9196);
nor U9439 (N_9439,N_8805,N_8970);
xor U9440 (N_9440,N_9155,N_8805);
and U9441 (N_9441,N_8868,N_9061);
or U9442 (N_9442,N_9169,N_9080);
xor U9443 (N_9443,N_9129,N_9173);
xnor U9444 (N_9444,N_9077,N_9041);
nor U9445 (N_9445,N_9082,N_9167);
xor U9446 (N_9446,N_9142,N_8885);
nand U9447 (N_9447,N_8930,N_8800);
nor U9448 (N_9448,N_9142,N_8821);
nand U9449 (N_9449,N_8875,N_9154);
xnor U9450 (N_9450,N_8813,N_8810);
and U9451 (N_9451,N_8949,N_9015);
and U9452 (N_9452,N_8901,N_8961);
xnor U9453 (N_9453,N_8860,N_8974);
and U9454 (N_9454,N_9193,N_8862);
nor U9455 (N_9455,N_9092,N_8890);
xor U9456 (N_9456,N_9180,N_9035);
nand U9457 (N_9457,N_9060,N_8810);
and U9458 (N_9458,N_8936,N_9122);
or U9459 (N_9459,N_9032,N_9124);
nand U9460 (N_9460,N_9188,N_9136);
or U9461 (N_9461,N_9130,N_8945);
and U9462 (N_9462,N_9172,N_8966);
or U9463 (N_9463,N_9139,N_8944);
or U9464 (N_9464,N_9028,N_8880);
and U9465 (N_9465,N_8964,N_9100);
nor U9466 (N_9466,N_9182,N_9187);
and U9467 (N_9467,N_8905,N_9084);
nor U9468 (N_9468,N_9159,N_9060);
nor U9469 (N_9469,N_9005,N_9168);
xor U9470 (N_9470,N_8859,N_8933);
nor U9471 (N_9471,N_8979,N_9050);
or U9472 (N_9472,N_8856,N_9072);
xnor U9473 (N_9473,N_8934,N_9165);
or U9474 (N_9474,N_9186,N_8833);
nand U9475 (N_9475,N_9166,N_8871);
or U9476 (N_9476,N_9021,N_9093);
or U9477 (N_9477,N_8940,N_9151);
and U9478 (N_9478,N_9158,N_9055);
nand U9479 (N_9479,N_8824,N_8904);
or U9480 (N_9480,N_8954,N_9091);
nor U9481 (N_9481,N_8931,N_8861);
and U9482 (N_9482,N_8806,N_9019);
xor U9483 (N_9483,N_8963,N_9117);
and U9484 (N_9484,N_8968,N_8932);
nand U9485 (N_9485,N_8801,N_9161);
xnor U9486 (N_9486,N_8820,N_9029);
nand U9487 (N_9487,N_8825,N_9180);
or U9488 (N_9488,N_8824,N_8866);
nand U9489 (N_9489,N_8928,N_8974);
xor U9490 (N_9490,N_9011,N_8816);
or U9491 (N_9491,N_8942,N_8944);
nor U9492 (N_9492,N_9075,N_9024);
nor U9493 (N_9493,N_9149,N_8845);
and U9494 (N_9494,N_9070,N_9077);
nor U9495 (N_9495,N_8890,N_9091);
nand U9496 (N_9496,N_9079,N_8996);
xor U9497 (N_9497,N_9156,N_9166);
nor U9498 (N_9498,N_9059,N_8895);
nor U9499 (N_9499,N_8885,N_8973);
xnor U9500 (N_9500,N_9023,N_9194);
nor U9501 (N_9501,N_8963,N_8824);
xor U9502 (N_9502,N_9126,N_8966);
xnor U9503 (N_9503,N_9114,N_8935);
or U9504 (N_9504,N_9004,N_9001);
nand U9505 (N_9505,N_9141,N_8934);
xnor U9506 (N_9506,N_8809,N_8884);
xnor U9507 (N_9507,N_8975,N_9009);
xnor U9508 (N_9508,N_8991,N_9084);
and U9509 (N_9509,N_9117,N_8934);
or U9510 (N_9510,N_9034,N_9008);
or U9511 (N_9511,N_8980,N_8893);
nor U9512 (N_9512,N_9093,N_8904);
xnor U9513 (N_9513,N_8840,N_9121);
nand U9514 (N_9514,N_9165,N_8983);
nor U9515 (N_9515,N_8858,N_8857);
and U9516 (N_9516,N_8852,N_8830);
or U9517 (N_9517,N_9141,N_8924);
nor U9518 (N_9518,N_9153,N_8900);
nand U9519 (N_9519,N_9161,N_8915);
or U9520 (N_9520,N_9165,N_8978);
nand U9521 (N_9521,N_9169,N_8986);
and U9522 (N_9522,N_9122,N_9119);
nor U9523 (N_9523,N_9092,N_8804);
nand U9524 (N_9524,N_9177,N_8801);
and U9525 (N_9525,N_9003,N_9032);
or U9526 (N_9526,N_8924,N_8987);
xnor U9527 (N_9527,N_9019,N_9190);
nor U9528 (N_9528,N_8930,N_9058);
nand U9529 (N_9529,N_8953,N_8825);
or U9530 (N_9530,N_9058,N_8932);
xor U9531 (N_9531,N_9157,N_9108);
and U9532 (N_9532,N_9082,N_8828);
nand U9533 (N_9533,N_9192,N_9024);
xor U9534 (N_9534,N_9030,N_9139);
xnor U9535 (N_9535,N_8958,N_9160);
or U9536 (N_9536,N_8990,N_8950);
and U9537 (N_9537,N_9085,N_9114);
nand U9538 (N_9538,N_8925,N_9109);
and U9539 (N_9539,N_9097,N_8969);
nand U9540 (N_9540,N_8966,N_8840);
and U9541 (N_9541,N_9168,N_8895);
xnor U9542 (N_9542,N_9061,N_8950);
and U9543 (N_9543,N_8944,N_8940);
and U9544 (N_9544,N_9182,N_9153);
nand U9545 (N_9545,N_9059,N_8902);
or U9546 (N_9546,N_8887,N_9162);
xnor U9547 (N_9547,N_8889,N_8902);
or U9548 (N_9548,N_9152,N_9101);
xor U9549 (N_9549,N_9087,N_8889);
xnor U9550 (N_9550,N_9095,N_8848);
and U9551 (N_9551,N_8857,N_9071);
and U9552 (N_9552,N_8896,N_9090);
xnor U9553 (N_9553,N_9170,N_9160);
or U9554 (N_9554,N_8966,N_8872);
and U9555 (N_9555,N_9136,N_9167);
nor U9556 (N_9556,N_9104,N_9114);
nor U9557 (N_9557,N_8846,N_9004);
xor U9558 (N_9558,N_9031,N_9070);
and U9559 (N_9559,N_9121,N_8899);
and U9560 (N_9560,N_8922,N_8800);
xor U9561 (N_9561,N_8955,N_8855);
nand U9562 (N_9562,N_8809,N_9038);
nor U9563 (N_9563,N_9083,N_9086);
nand U9564 (N_9564,N_8931,N_8830);
xnor U9565 (N_9565,N_8952,N_9130);
nand U9566 (N_9566,N_9117,N_8929);
or U9567 (N_9567,N_8836,N_8930);
or U9568 (N_9568,N_8846,N_9040);
nand U9569 (N_9569,N_9073,N_8954);
xnor U9570 (N_9570,N_9111,N_9032);
xnor U9571 (N_9571,N_9124,N_9042);
and U9572 (N_9572,N_9185,N_9092);
nand U9573 (N_9573,N_9172,N_8823);
or U9574 (N_9574,N_8888,N_8973);
nor U9575 (N_9575,N_8993,N_8815);
nand U9576 (N_9576,N_8975,N_8917);
and U9577 (N_9577,N_8949,N_9135);
xor U9578 (N_9578,N_9053,N_9065);
nor U9579 (N_9579,N_8892,N_9107);
nand U9580 (N_9580,N_9187,N_9096);
nand U9581 (N_9581,N_9129,N_8933);
nor U9582 (N_9582,N_9157,N_8858);
xnor U9583 (N_9583,N_8929,N_9074);
xor U9584 (N_9584,N_8819,N_9169);
and U9585 (N_9585,N_9150,N_9106);
xnor U9586 (N_9586,N_8825,N_9127);
nand U9587 (N_9587,N_9162,N_8899);
or U9588 (N_9588,N_9051,N_9108);
and U9589 (N_9589,N_9071,N_9179);
nor U9590 (N_9590,N_8980,N_9109);
xnor U9591 (N_9591,N_8952,N_8983);
nor U9592 (N_9592,N_8915,N_9152);
or U9593 (N_9593,N_8879,N_8953);
nor U9594 (N_9594,N_9069,N_8811);
or U9595 (N_9595,N_9194,N_8977);
nor U9596 (N_9596,N_8926,N_8858);
and U9597 (N_9597,N_8856,N_8904);
or U9598 (N_9598,N_8827,N_9120);
or U9599 (N_9599,N_9147,N_8835);
xnor U9600 (N_9600,N_9590,N_9417);
nand U9601 (N_9601,N_9379,N_9233);
or U9602 (N_9602,N_9529,N_9224);
and U9603 (N_9603,N_9201,N_9505);
xnor U9604 (N_9604,N_9205,N_9351);
nor U9605 (N_9605,N_9383,N_9521);
or U9606 (N_9606,N_9561,N_9281);
nor U9607 (N_9607,N_9519,N_9362);
and U9608 (N_9608,N_9592,N_9332);
and U9609 (N_9609,N_9356,N_9585);
nand U9610 (N_9610,N_9532,N_9578);
nand U9611 (N_9611,N_9345,N_9290);
nor U9612 (N_9612,N_9477,N_9352);
or U9613 (N_9613,N_9469,N_9490);
xnor U9614 (N_9614,N_9598,N_9381);
nor U9615 (N_9615,N_9367,N_9230);
nand U9616 (N_9616,N_9577,N_9220);
and U9617 (N_9617,N_9580,N_9441);
or U9618 (N_9618,N_9508,N_9416);
and U9619 (N_9619,N_9338,N_9510);
xor U9620 (N_9620,N_9301,N_9507);
xor U9621 (N_9621,N_9599,N_9213);
xor U9622 (N_9622,N_9438,N_9494);
and U9623 (N_9623,N_9531,N_9273);
or U9624 (N_9624,N_9516,N_9567);
nor U9625 (N_9625,N_9422,N_9455);
nor U9626 (N_9626,N_9323,N_9556);
and U9627 (N_9627,N_9309,N_9265);
xor U9628 (N_9628,N_9513,N_9232);
nand U9629 (N_9629,N_9541,N_9331);
nor U9630 (N_9630,N_9550,N_9304);
or U9631 (N_9631,N_9515,N_9482);
xor U9632 (N_9632,N_9415,N_9387);
and U9633 (N_9633,N_9373,N_9570);
and U9634 (N_9634,N_9405,N_9341);
xnor U9635 (N_9635,N_9231,N_9500);
or U9636 (N_9636,N_9354,N_9461);
nor U9637 (N_9637,N_9202,N_9495);
or U9638 (N_9638,N_9536,N_9451);
xor U9639 (N_9639,N_9374,N_9312);
nor U9640 (N_9640,N_9491,N_9499);
or U9641 (N_9641,N_9384,N_9487);
or U9642 (N_9642,N_9317,N_9294);
nand U9643 (N_9643,N_9307,N_9504);
nor U9644 (N_9644,N_9483,N_9464);
nand U9645 (N_9645,N_9424,N_9446);
nor U9646 (N_9646,N_9474,N_9343);
nand U9647 (N_9647,N_9569,N_9239);
xor U9648 (N_9648,N_9511,N_9584);
and U9649 (N_9649,N_9314,N_9385);
nand U9650 (N_9650,N_9544,N_9412);
nor U9651 (N_9651,N_9501,N_9478);
or U9652 (N_9652,N_9542,N_9223);
xor U9653 (N_9653,N_9523,N_9260);
or U9654 (N_9654,N_9277,N_9439);
nand U9655 (N_9655,N_9392,N_9371);
nand U9656 (N_9656,N_9245,N_9251);
nor U9657 (N_9657,N_9316,N_9472);
xnor U9658 (N_9658,N_9517,N_9503);
or U9659 (N_9659,N_9335,N_9388);
or U9660 (N_9660,N_9574,N_9467);
and U9661 (N_9661,N_9221,N_9305);
xor U9662 (N_9662,N_9407,N_9410);
and U9663 (N_9663,N_9404,N_9207);
nand U9664 (N_9664,N_9400,N_9372);
xor U9665 (N_9665,N_9236,N_9360);
nor U9666 (N_9666,N_9342,N_9428);
nor U9667 (N_9667,N_9576,N_9364);
and U9668 (N_9668,N_9300,N_9234);
and U9669 (N_9669,N_9369,N_9484);
or U9670 (N_9670,N_9526,N_9460);
xor U9671 (N_9671,N_9525,N_9426);
xnor U9672 (N_9672,N_9206,N_9297);
nor U9673 (N_9673,N_9311,N_9434);
and U9674 (N_9674,N_9324,N_9328);
xnor U9675 (N_9675,N_9594,N_9359);
or U9676 (N_9676,N_9571,N_9453);
or U9677 (N_9677,N_9272,N_9226);
nand U9678 (N_9678,N_9255,N_9545);
nor U9679 (N_9679,N_9564,N_9268);
and U9680 (N_9680,N_9361,N_9419);
and U9681 (N_9681,N_9566,N_9572);
xor U9682 (N_9682,N_9411,N_9527);
xor U9683 (N_9683,N_9380,N_9555);
xor U9684 (N_9684,N_9518,N_9241);
nand U9685 (N_9685,N_9459,N_9514);
nand U9686 (N_9686,N_9246,N_9270);
nor U9687 (N_9687,N_9588,N_9480);
nand U9688 (N_9688,N_9222,N_9319);
nand U9689 (N_9689,N_9528,N_9313);
and U9690 (N_9690,N_9449,N_9349);
xor U9691 (N_9691,N_9267,N_9326);
nand U9692 (N_9692,N_9425,N_9302);
nand U9693 (N_9693,N_9211,N_9522);
xor U9694 (N_9694,N_9465,N_9493);
and U9695 (N_9695,N_9492,N_9414);
xor U9696 (N_9696,N_9466,N_9393);
and U9697 (N_9697,N_9225,N_9378);
and U9698 (N_9698,N_9248,N_9558);
and U9699 (N_9699,N_9210,N_9308);
nand U9700 (N_9700,N_9420,N_9554);
and U9701 (N_9701,N_9370,N_9581);
or U9702 (N_9702,N_9448,N_9587);
xnor U9703 (N_9703,N_9442,N_9237);
and U9704 (N_9704,N_9546,N_9204);
nand U9705 (N_9705,N_9346,N_9291);
nor U9706 (N_9706,N_9471,N_9457);
nand U9707 (N_9707,N_9318,N_9427);
nand U9708 (N_9708,N_9247,N_9595);
or U9709 (N_9709,N_9396,N_9252);
or U9710 (N_9710,N_9560,N_9520);
xor U9711 (N_9711,N_9235,N_9573);
nand U9712 (N_9712,N_9200,N_9485);
nor U9713 (N_9713,N_9287,N_9274);
xor U9714 (N_9714,N_9583,N_9450);
and U9715 (N_9715,N_9243,N_9497);
nand U9716 (N_9716,N_9437,N_9533);
nor U9717 (N_9717,N_9279,N_9452);
and U9718 (N_9718,N_9463,N_9445);
xor U9719 (N_9719,N_9266,N_9512);
xnor U9720 (N_9720,N_9489,N_9408);
or U9721 (N_9721,N_9275,N_9218);
and U9722 (N_9722,N_9543,N_9339);
and U9723 (N_9723,N_9292,N_9551);
xnor U9724 (N_9724,N_9325,N_9276);
nor U9725 (N_9725,N_9329,N_9348);
xnor U9726 (N_9726,N_9476,N_9386);
xnor U9727 (N_9727,N_9462,N_9219);
or U9728 (N_9728,N_9436,N_9389);
nand U9729 (N_9729,N_9227,N_9432);
or U9730 (N_9730,N_9303,N_9443);
nor U9731 (N_9731,N_9229,N_9208);
xor U9732 (N_9732,N_9262,N_9336);
nand U9733 (N_9733,N_9582,N_9563);
nand U9734 (N_9734,N_9397,N_9535);
or U9735 (N_9735,N_9358,N_9409);
nor U9736 (N_9736,N_9306,N_9557);
xnor U9737 (N_9737,N_9263,N_9423);
and U9738 (N_9738,N_9586,N_9315);
nand U9739 (N_9739,N_9203,N_9481);
xor U9740 (N_9740,N_9429,N_9575);
or U9741 (N_9741,N_9299,N_9447);
and U9742 (N_9742,N_9261,N_9395);
or U9743 (N_9743,N_9456,N_9548);
nand U9744 (N_9744,N_9391,N_9347);
nor U9745 (N_9745,N_9524,N_9254);
nand U9746 (N_9746,N_9288,N_9547);
xnor U9747 (N_9747,N_9298,N_9209);
or U9748 (N_9748,N_9539,N_9280);
and U9749 (N_9749,N_9394,N_9321);
nand U9750 (N_9750,N_9264,N_9212);
xnor U9751 (N_9751,N_9534,N_9470);
xnor U9752 (N_9752,N_9435,N_9390);
nor U9753 (N_9753,N_9250,N_9402);
xor U9754 (N_9754,N_9431,N_9398);
and U9755 (N_9755,N_9228,N_9216);
nor U9756 (N_9756,N_9355,N_9399);
and U9757 (N_9757,N_9320,N_9363);
nand U9758 (N_9758,N_9552,N_9337);
nand U9759 (N_9759,N_9553,N_9568);
and U9760 (N_9760,N_9350,N_9589);
xnor U9761 (N_9761,N_9256,N_9368);
and U9762 (N_9762,N_9334,N_9295);
or U9763 (N_9763,N_9454,N_9509);
or U9764 (N_9764,N_9418,N_9538);
nand U9765 (N_9765,N_9240,N_9283);
xnor U9766 (N_9766,N_9382,N_9502);
xor U9767 (N_9767,N_9406,N_9488);
xnor U9768 (N_9768,N_9579,N_9440);
xnor U9769 (N_9769,N_9330,N_9282);
and U9770 (N_9770,N_9597,N_9468);
xnor U9771 (N_9771,N_9214,N_9421);
nand U9772 (N_9772,N_9530,N_9498);
xnor U9773 (N_9773,N_9333,N_9296);
nor U9774 (N_9774,N_9249,N_9479);
nor U9775 (N_9775,N_9596,N_9565);
or U9776 (N_9776,N_9413,N_9540);
xor U9777 (N_9777,N_9591,N_9278);
nor U9778 (N_9778,N_9458,N_9549);
xor U9779 (N_9779,N_9475,N_9327);
xor U9780 (N_9780,N_9257,N_9286);
nand U9781 (N_9781,N_9238,N_9537);
or U9782 (N_9782,N_9403,N_9593);
or U9783 (N_9783,N_9215,N_9285);
and U9784 (N_9784,N_9258,N_9293);
or U9785 (N_9785,N_9496,N_9562);
xnor U9786 (N_9786,N_9506,N_9244);
and U9787 (N_9787,N_9433,N_9271);
and U9788 (N_9788,N_9444,N_9217);
xor U9789 (N_9789,N_9357,N_9259);
xnor U9790 (N_9790,N_9344,N_9365);
nor U9791 (N_9791,N_9310,N_9430);
or U9792 (N_9792,N_9377,N_9353);
and U9793 (N_9793,N_9269,N_9486);
or U9794 (N_9794,N_9366,N_9289);
or U9795 (N_9795,N_9340,N_9322);
nor U9796 (N_9796,N_9375,N_9242);
xor U9797 (N_9797,N_9253,N_9376);
or U9798 (N_9798,N_9559,N_9401);
nor U9799 (N_9799,N_9473,N_9284);
nor U9800 (N_9800,N_9200,N_9533);
and U9801 (N_9801,N_9442,N_9348);
or U9802 (N_9802,N_9452,N_9339);
nand U9803 (N_9803,N_9572,N_9585);
xnor U9804 (N_9804,N_9293,N_9538);
or U9805 (N_9805,N_9417,N_9221);
and U9806 (N_9806,N_9320,N_9505);
nor U9807 (N_9807,N_9308,N_9541);
and U9808 (N_9808,N_9421,N_9227);
and U9809 (N_9809,N_9563,N_9479);
nor U9810 (N_9810,N_9202,N_9304);
or U9811 (N_9811,N_9568,N_9547);
or U9812 (N_9812,N_9389,N_9458);
and U9813 (N_9813,N_9413,N_9410);
xor U9814 (N_9814,N_9468,N_9340);
and U9815 (N_9815,N_9341,N_9479);
or U9816 (N_9816,N_9273,N_9235);
nand U9817 (N_9817,N_9596,N_9485);
nand U9818 (N_9818,N_9356,N_9399);
and U9819 (N_9819,N_9548,N_9317);
and U9820 (N_9820,N_9296,N_9594);
and U9821 (N_9821,N_9390,N_9331);
xnor U9822 (N_9822,N_9413,N_9392);
xnor U9823 (N_9823,N_9217,N_9475);
xor U9824 (N_9824,N_9238,N_9243);
nand U9825 (N_9825,N_9540,N_9465);
or U9826 (N_9826,N_9534,N_9396);
nand U9827 (N_9827,N_9443,N_9350);
or U9828 (N_9828,N_9351,N_9397);
or U9829 (N_9829,N_9395,N_9522);
and U9830 (N_9830,N_9359,N_9549);
or U9831 (N_9831,N_9553,N_9508);
nand U9832 (N_9832,N_9457,N_9426);
nand U9833 (N_9833,N_9446,N_9331);
or U9834 (N_9834,N_9540,N_9365);
nand U9835 (N_9835,N_9276,N_9266);
or U9836 (N_9836,N_9476,N_9574);
nor U9837 (N_9837,N_9514,N_9574);
or U9838 (N_9838,N_9426,N_9575);
and U9839 (N_9839,N_9582,N_9235);
nor U9840 (N_9840,N_9301,N_9238);
or U9841 (N_9841,N_9221,N_9210);
or U9842 (N_9842,N_9353,N_9560);
xor U9843 (N_9843,N_9337,N_9526);
xnor U9844 (N_9844,N_9291,N_9441);
nand U9845 (N_9845,N_9392,N_9569);
nand U9846 (N_9846,N_9510,N_9325);
nand U9847 (N_9847,N_9534,N_9293);
and U9848 (N_9848,N_9501,N_9326);
xor U9849 (N_9849,N_9543,N_9294);
nor U9850 (N_9850,N_9582,N_9465);
nand U9851 (N_9851,N_9440,N_9505);
and U9852 (N_9852,N_9413,N_9258);
nand U9853 (N_9853,N_9269,N_9388);
nor U9854 (N_9854,N_9353,N_9216);
and U9855 (N_9855,N_9201,N_9351);
and U9856 (N_9856,N_9492,N_9240);
and U9857 (N_9857,N_9267,N_9508);
nand U9858 (N_9858,N_9375,N_9287);
or U9859 (N_9859,N_9286,N_9542);
or U9860 (N_9860,N_9441,N_9547);
xor U9861 (N_9861,N_9530,N_9309);
nor U9862 (N_9862,N_9211,N_9305);
nand U9863 (N_9863,N_9351,N_9421);
xor U9864 (N_9864,N_9373,N_9380);
xor U9865 (N_9865,N_9410,N_9316);
nand U9866 (N_9866,N_9249,N_9297);
and U9867 (N_9867,N_9579,N_9264);
nand U9868 (N_9868,N_9406,N_9556);
nand U9869 (N_9869,N_9527,N_9477);
nor U9870 (N_9870,N_9452,N_9398);
or U9871 (N_9871,N_9558,N_9480);
xor U9872 (N_9872,N_9407,N_9207);
nand U9873 (N_9873,N_9287,N_9581);
and U9874 (N_9874,N_9387,N_9469);
nand U9875 (N_9875,N_9564,N_9403);
nand U9876 (N_9876,N_9334,N_9441);
nor U9877 (N_9877,N_9392,N_9242);
and U9878 (N_9878,N_9405,N_9534);
nor U9879 (N_9879,N_9418,N_9361);
nand U9880 (N_9880,N_9425,N_9573);
nor U9881 (N_9881,N_9432,N_9503);
or U9882 (N_9882,N_9425,N_9248);
xor U9883 (N_9883,N_9477,N_9582);
and U9884 (N_9884,N_9223,N_9216);
and U9885 (N_9885,N_9512,N_9370);
nor U9886 (N_9886,N_9477,N_9220);
nor U9887 (N_9887,N_9483,N_9577);
nor U9888 (N_9888,N_9389,N_9261);
nand U9889 (N_9889,N_9287,N_9489);
xnor U9890 (N_9890,N_9401,N_9484);
and U9891 (N_9891,N_9486,N_9529);
nand U9892 (N_9892,N_9387,N_9446);
or U9893 (N_9893,N_9526,N_9347);
nor U9894 (N_9894,N_9205,N_9516);
xnor U9895 (N_9895,N_9534,N_9386);
nand U9896 (N_9896,N_9212,N_9513);
nor U9897 (N_9897,N_9408,N_9563);
or U9898 (N_9898,N_9460,N_9489);
and U9899 (N_9899,N_9218,N_9355);
xor U9900 (N_9900,N_9373,N_9514);
nor U9901 (N_9901,N_9365,N_9422);
nor U9902 (N_9902,N_9353,N_9427);
nand U9903 (N_9903,N_9292,N_9399);
nand U9904 (N_9904,N_9597,N_9559);
and U9905 (N_9905,N_9234,N_9351);
or U9906 (N_9906,N_9441,N_9306);
or U9907 (N_9907,N_9404,N_9386);
xor U9908 (N_9908,N_9380,N_9576);
or U9909 (N_9909,N_9344,N_9375);
xnor U9910 (N_9910,N_9419,N_9522);
or U9911 (N_9911,N_9213,N_9568);
and U9912 (N_9912,N_9473,N_9515);
xnor U9913 (N_9913,N_9326,N_9592);
nand U9914 (N_9914,N_9529,N_9474);
and U9915 (N_9915,N_9283,N_9235);
nand U9916 (N_9916,N_9562,N_9218);
nand U9917 (N_9917,N_9387,N_9351);
nor U9918 (N_9918,N_9309,N_9372);
and U9919 (N_9919,N_9502,N_9392);
nand U9920 (N_9920,N_9543,N_9235);
xnor U9921 (N_9921,N_9412,N_9489);
xor U9922 (N_9922,N_9432,N_9548);
or U9923 (N_9923,N_9330,N_9597);
or U9924 (N_9924,N_9241,N_9353);
or U9925 (N_9925,N_9477,N_9427);
and U9926 (N_9926,N_9280,N_9212);
or U9927 (N_9927,N_9235,N_9581);
xor U9928 (N_9928,N_9233,N_9514);
xor U9929 (N_9929,N_9540,N_9220);
and U9930 (N_9930,N_9429,N_9243);
and U9931 (N_9931,N_9371,N_9548);
nand U9932 (N_9932,N_9590,N_9566);
nor U9933 (N_9933,N_9476,N_9216);
or U9934 (N_9934,N_9581,N_9559);
xnor U9935 (N_9935,N_9598,N_9469);
and U9936 (N_9936,N_9278,N_9522);
or U9937 (N_9937,N_9332,N_9564);
nor U9938 (N_9938,N_9311,N_9275);
nor U9939 (N_9939,N_9387,N_9580);
nor U9940 (N_9940,N_9333,N_9424);
nor U9941 (N_9941,N_9276,N_9516);
and U9942 (N_9942,N_9547,N_9597);
or U9943 (N_9943,N_9250,N_9479);
and U9944 (N_9944,N_9372,N_9226);
and U9945 (N_9945,N_9391,N_9504);
or U9946 (N_9946,N_9593,N_9535);
nor U9947 (N_9947,N_9464,N_9243);
xor U9948 (N_9948,N_9253,N_9355);
and U9949 (N_9949,N_9509,N_9586);
and U9950 (N_9950,N_9455,N_9534);
or U9951 (N_9951,N_9228,N_9431);
nand U9952 (N_9952,N_9334,N_9456);
nor U9953 (N_9953,N_9323,N_9461);
and U9954 (N_9954,N_9506,N_9208);
nor U9955 (N_9955,N_9350,N_9541);
and U9956 (N_9956,N_9326,N_9575);
xor U9957 (N_9957,N_9557,N_9591);
or U9958 (N_9958,N_9563,N_9340);
nand U9959 (N_9959,N_9318,N_9391);
xor U9960 (N_9960,N_9248,N_9252);
nor U9961 (N_9961,N_9391,N_9219);
nor U9962 (N_9962,N_9276,N_9474);
or U9963 (N_9963,N_9535,N_9272);
nor U9964 (N_9964,N_9495,N_9244);
nor U9965 (N_9965,N_9249,N_9313);
or U9966 (N_9966,N_9333,N_9569);
nor U9967 (N_9967,N_9499,N_9212);
nor U9968 (N_9968,N_9367,N_9532);
or U9969 (N_9969,N_9550,N_9449);
nand U9970 (N_9970,N_9397,N_9289);
nand U9971 (N_9971,N_9586,N_9495);
and U9972 (N_9972,N_9442,N_9278);
and U9973 (N_9973,N_9358,N_9278);
and U9974 (N_9974,N_9328,N_9376);
and U9975 (N_9975,N_9445,N_9450);
nand U9976 (N_9976,N_9235,N_9560);
or U9977 (N_9977,N_9346,N_9212);
or U9978 (N_9978,N_9283,N_9226);
nand U9979 (N_9979,N_9329,N_9425);
and U9980 (N_9980,N_9356,N_9264);
xor U9981 (N_9981,N_9432,N_9519);
xor U9982 (N_9982,N_9216,N_9536);
nand U9983 (N_9983,N_9288,N_9379);
or U9984 (N_9984,N_9457,N_9395);
nand U9985 (N_9985,N_9505,N_9303);
nand U9986 (N_9986,N_9200,N_9384);
or U9987 (N_9987,N_9355,N_9523);
nand U9988 (N_9988,N_9419,N_9347);
xnor U9989 (N_9989,N_9470,N_9591);
xor U9990 (N_9990,N_9372,N_9249);
xnor U9991 (N_9991,N_9556,N_9234);
nor U9992 (N_9992,N_9255,N_9248);
xor U9993 (N_9993,N_9260,N_9532);
nand U9994 (N_9994,N_9518,N_9583);
nor U9995 (N_9995,N_9226,N_9421);
xor U9996 (N_9996,N_9535,N_9373);
xor U9997 (N_9997,N_9206,N_9363);
and U9998 (N_9998,N_9353,N_9458);
and U9999 (N_9999,N_9371,N_9430);
or U10000 (N_10000,N_9607,N_9878);
or U10001 (N_10001,N_9813,N_9941);
or U10002 (N_10002,N_9685,N_9912);
or U10003 (N_10003,N_9815,N_9672);
nor U10004 (N_10004,N_9677,N_9872);
xnor U10005 (N_10005,N_9879,N_9737);
nand U10006 (N_10006,N_9951,N_9786);
xnor U10007 (N_10007,N_9663,N_9850);
xnor U10008 (N_10008,N_9741,N_9969);
nand U10009 (N_10009,N_9642,N_9958);
xor U10010 (N_10010,N_9604,N_9844);
nand U10011 (N_10011,N_9706,N_9954);
and U10012 (N_10012,N_9933,N_9673);
or U10013 (N_10013,N_9890,N_9876);
xnor U10014 (N_10014,N_9978,N_9659);
and U10015 (N_10015,N_9873,N_9687);
or U10016 (N_10016,N_9603,N_9913);
nand U10017 (N_10017,N_9667,N_9789);
nand U10018 (N_10018,N_9788,N_9654);
or U10019 (N_10019,N_9960,N_9992);
xnor U10020 (N_10020,N_9961,N_9932);
and U10021 (N_10021,N_9860,N_9718);
and U10022 (N_10022,N_9605,N_9657);
nor U10023 (N_10023,N_9660,N_9797);
nand U10024 (N_10024,N_9675,N_9758);
xor U10025 (N_10025,N_9802,N_9602);
nand U10026 (N_10026,N_9778,N_9921);
and U10027 (N_10027,N_9926,N_9753);
nand U10028 (N_10028,N_9980,N_9828);
and U10029 (N_10029,N_9865,N_9875);
nand U10030 (N_10030,N_9708,N_9738);
nor U10031 (N_10031,N_9819,N_9909);
xor U10032 (N_10032,N_9982,N_9920);
nor U10033 (N_10033,N_9855,N_9769);
xor U10034 (N_10034,N_9952,N_9714);
nor U10035 (N_10035,N_9653,N_9794);
nor U10036 (N_10036,N_9745,N_9742);
or U10037 (N_10037,N_9820,N_9720);
nor U10038 (N_10038,N_9825,N_9793);
nand U10039 (N_10039,N_9867,N_9905);
and U10040 (N_10040,N_9956,N_9883);
and U10041 (N_10041,N_9732,N_9785);
and U10042 (N_10042,N_9767,N_9988);
and U10043 (N_10043,N_9827,N_9638);
and U10044 (N_10044,N_9822,N_9947);
xnor U10045 (N_10045,N_9811,N_9935);
and U10046 (N_10046,N_9632,N_9945);
and U10047 (N_10047,N_9981,N_9974);
xor U10048 (N_10048,N_9645,N_9678);
nor U10049 (N_10049,N_9998,N_9948);
xor U10050 (N_10050,N_9782,N_9842);
or U10051 (N_10051,N_9666,N_9936);
xor U10052 (N_10052,N_9818,N_9962);
and U10053 (N_10053,N_9757,N_9845);
and U10054 (N_10054,N_9702,N_9655);
xor U10055 (N_10055,N_9907,N_9885);
nand U10056 (N_10056,N_9836,N_9634);
and U10057 (N_10057,N_9967,N_9834);
nand U10058 (N_10058,N_9959,N_9930);
or U10059 (N_10059,N_9996,N_9650);
and U10060 (N_10060,N_9643,N_9616);
nor U10061 (N_10061,N_9692,N_9977);
nor U10062 (N_10062,N_9739,N_9862);
and U10063 (N_10063,N_9887,N_9929);
or U10064 (N_10064,N_9937,N_9826);
nand U10065 (N_10065,N_9814,N_9976);
nand U10066 (N_10066,N_9630,N_9622);
nand U10067 (N_10067,N_9970,N_9640);
nand U10068 (N_10068,N_9777,N_9779);
and U10069 (N_10069,N_9669,N_9809);
xor U10070 (N_10070,N_9609,N_9759);
and U10071 (N_10071,N_9829,N_9953);
and U10072 (N_10072,N_9755,N_9805);
xnor U10073 (N_10073,N_9899,N_9696);
or U10074 (N_10074,N_9621,N_9983);
nor U10075 (N_10075,N_9727,N_9715);
xnor U10076 (N_10076,N_9808,N_9812);
or U10077 (N_10077,N_9939,N_9735);
and U10078 (N_10078,N_9631,N_9641);
and U10079 (N_10079,N_9656,N_9651);
xor U10080 (N_10080,N_9636,N_9683);
nand U10081 (N_10081,N_9858,N_9944);
nand U10082 (N_10082,N_9816,N_9923);
or U10083 (N_10083,N_9810,N_9756);
nand U10084 (N_10084,N_9821,N_9750);
xor U10085 (N_10085,N_9796,N_9963);
and U10086 (N_10086,N_9868,N_9997);
and U10087 (N_10087,N_9721,N_9830);
nand U10088 (N_10088,N_9852,N_9924);
nand U10089 (N_10089,N_9851,N_9861);
or U10090 (N_10090,N_9902,N_9774);
and U10091 (N_10091,N_9882,N_9938);
xnor U10092 (N_10092,N_9646,N_9712);
nand U10093 (N_10093,N_9940,N_9679);
and U10094 (N_10094,N_9984,N_9760);
or U10095 (N_10095,N_9994,N_9698);
or U10096 (N_10096,N_9689,N_9693);
or U10097 (N_10097,N_9849,N_9620);
nand U10098 (N_10098,N_9991,N_9705);
or U10099 (N_10099,N_9823,N_9990);
xor U10100 (N_10100,N_9623,N_9649);
or U10101 (N_10101,N_9743,N_9763);
nand U10102 (N_10102,N_9859,N_9608);
nor U10103 (N_10103,N_9931,N_9754);
and U10104 (N_10104,N_9837,N_9627);
or U10105 (N_10105,N_9892,N_9880);
xor U10106 (N_10106,N_9889,N_9787);
xnor U10107 (N_10107,N_9717,N_9729);
xor U10108 (N_10108,N_9606,N_9847);
or U10109 (N_10109,N_9668,N_9765);
nand U10110 (N_10110,N_9671,N_9662);
xnor U10111 (N_10111,N_9695,N_9874);
and U10112 (N_10112,N_9615,N_9619);
and U10113 (N_10113,N_9824,N_9895);
xnor U10114 (N_10114,N_9985,N_9888);
and U10115 (N_10115,N_9870,N_9807);
nand U10116 (N_10116,N_9803,N_9910);
nand U10117 (N_10117,N_9833,N_9674);
nor U10118 (N_10118,N_9770,N_9731);
nor U10119 (N_10119,N_9904,N_9886);
nand U10120 (N_10120,N_9676,N_9804);
xnor U10121 (N_10121,N_9658,N_9934);
or U10122 (N_10122,N_9749,N_9800);
or U10123 (N_10123,N_9681,N_9841);
nand U10124 (N_10124,N_9764,N_9617);
and U10125 (N_10125,N_9752,N_9791);
nand U10126 (N_10126,N_9831,N_9748);
nand U10127 (N_10127,N_9848,N_9968);
xor U10128 (N_10128,N_9915,N_9894);
nand U10129 (N_10129,N_9801,N_9942);
or U10130 (N_10130,N_9661,N_9680);
and U10131 (N_10131,N_9792,N_9795);
nand U10132 (N_10132,N_9776,N_9629);
nor U10133 (N_10133,N_9798,N_9625);
nor U10134 (N_10134,N_9916,N_9857);
or U10135 (N_10135,N_9744,N_9635);
nor U10136 (N_10136,N_9928,N_9688);
or U10137 (N_10137,N_9704,N_9711);
or U10138 (N_10138,N_9647,N_9747);
xnor U10139 (N_10139,N_9896,N_9613);
xor U10140 (N_10140,N_9866,N_9652);
nand U10141 (N_10141,N_9740,N_9703);
and U10142 (N_10142,N_9987,N_9806);
xnor U10143 (N_10143,N_9768,N_9919);
nor U10144 (N_10144,N_9908,N_9835);
or U10145 (N_10145,N_9843,N_9697);
xor U10146 (N_10146,N_9900,N_9897);
xor U10147 (N_10147,N_9684,N_9611);
nand U10148 (N_10148,N_9736,N_9964);
or U10149 (N_10149,N_9781,N_9869);
nor U10150 (N_10150,N_9863,N_9832);
xnor U10151 (N_10151,N_9709,N_9690);
or U10152 (N_10152,N_9898,N_9881);
xor U10153 (N_10153,N_9871,N_9734);
or U10154 (N_10154,N_9975,N_9965);
xor U10155 (N_10155,N_9775,N_9946);
and U10156 (N_10156,N_9628,N_9922);
xor U10157 (N_10157,N_9639,N_9906);
nor U10158 (N_10158,N_9618,N_9817);
nor U10159 (N_10159,N_9893,N_9884);
nand U10160 (N_10160,N_9700,N_9903);
and U10161 (N_10161,N_9986,N_9644);
nor U10162 (N_10162,N_9726,N_9971);
or U10163 (N_10163,N_9624,N_9979);
xnor U10164 (N_10164,N_9725,N_9966);
xnor U10165 (N_10165,N_9957,N_9633);
nand U10166 (N_10166,N_9600,N_9917);
nor U10167 (N_10167,N_9989,N_9761);
nor U10168 (N_10168,N_9790,N_9648);
nor U10169 (N_10169,N_9772,N_9840);
and U10170 (N_10170,N_9601,N_9995);
and U10171 (N_10171,N_9927,N_9846);
or U10172 (N_10172,N_9722,N_9955);
or U10173 (N_10173,N_9780,N_9854);
xor U10174 (N_10174,N_9877,N_9723);
or U10175 (N_10175,N_9838,N_9713);
xor U10176 (N_10176,N_9670,N_9864);
or U10177 (N_10177,N_9783,N_9891);
or U10178 (N_10178,N_9691,N_9724);
nor U10179 (N_10179,N_9943,N_9694);
or U10180 (N_10180,N_9733,N_9925);
xnor U10181 (N_10181,N_9637,N_9773);
nor U10182 (N_10182,N_9853,N_9614);
and U10183 (N_10183,N_9746,N_9973);
nor U10184 (N_10184,N_9999,N_9707);
nand U10185 (N_10185,N_9972,N_9839);
nor U10186 (N_10186,N_9710,N_9766);
and U10187 (N_10187,N_9784,N_9699);
and U10188 (N_10188,N_9856,N_9612);
xor U10189 (N_10189,N_9918,N_9664);
and U10190 (N_10190,N_9771,N_9799);
nor U10191 (N_10191,N_9762,N_9911);
or U10192 (N_10192,N_9949,N_9682);
and U10193 (N_10193,N_9626,N_9716);
nor U10194 (N_10194,N_9751,N_9730);
nor U10195 (N_10195,N_9686,N_9901);
and U10196 (N_10196,N_9701,N_9728);
or U10197 (N_10197,N_9719,N_9610);
and U10198 (N_10198,N_9914,N_9665);
and U10199 (N_10199,N_9950,N_9993);
nor U10200 (N_10200,N_9849,N_9954);
and U10201 (N_10201,N_9732,N_9931);
or U10202 (N_10202,N_9900,N_9911);
and U10203 (N_10203,N_9993,N_9854);
nor U10204 (N_10204,N_9841,N_9859);
nor U10205 (N_10205,N_9961,N_9937);
nor U10206 (N_10206,N_9868,N_9879);
xor U10207 (N_10207,N_9674,N_9735);
xor U10208 (N_10208,N_9862,N_9613);
and U10209 (N_10209,N_9973,N_9841);
nand U10210 (N_10210,N_9744,N_9607);
or U10211 (N_10211,N_9736,N_9870);
or U10212 (N_10212,N_9814,N_9805);
or U10213 (N_10213,N_9727,N_9742);
nand U10214 (N_10214,N_9674,N_9744);
and U10215 (N_10215,N_9849,N_9889);
and U10216 (N_10216,N_9740,N_9672);
or U10217 (N_10217,N_9799,N_9944);
nor U10218 (N_10218,N_9651,N_9699);
nand U10219 (N_10219,N_9824,N_9716);
nand U10220 (N_10220,N_9677,N_9728);
xnor U10221 (N_10221,N_9616,N_9817);
and U10222 (N_10222,N_9863,N_9943);
nor U10223 (N_10223,N_9878,N_9756);
nor U10224 (N_10224,N_9617,N_9672);
or U10225 (N_10225,N_9904,N_9771);
and U10226 (N_10226,N_9969,N_9636);
xor U10227 (N_10227,N_9893,N_9967);
or U10228 (N_10228,N_9806,N_9619);
xnor U10229 (N_10229,N_9700,N_9945);
xnor U10230 (N_10230,N_9713,N_9965);
nand U10231 (N_10231,N_9647,N_9820);
and U10232 (N_10232,N_9601,N_9973);
and U10233 (N_10233,N_9781,N_9632);
and U10234 (N_10234,N_9611,N_9979);
or U10235 (N_10235,N_9861,N_9836);
nor U10236 (N_10236,N_9751,N_9946);
xor U10237 (N_10237,N_9755,N_9743);
or U10238 (N_10238,N_9763,N_9703);
nor U10239 (N_10239,N_9879,N_9894);
nor U10240 (N_10240,N_9614,N_9732);
or U10241 (N_10241,N_9911,N_9971);
and U10242 (N_10242,N_9879,N_9985);
nor U10243 (N_10243,N_9750,N_9690);
nand U10244 (N_10244,N_9720,N_9961);
nor U10245 (N_10245,N_9947,N_9996);
and U10246 (N_10246,N_9956,N_9858);
nor U10247 (N_10247,N_9738,N_9876);
or U10248 (N_10248,N_9836,N_9721);
or U10249 (N_10249,N_9900,N_9753);
nand U10250 (N_10250,N_9785,N_9907);
and U10251 (N_10251,N_9943,N_9636);
or U10252 (N_10252,N_9649,N_9828);
xnor U10253 (N_10253,N_9918,N_9838);
xnor U10254 (N_10254,N_9878,N_9995);
and U10255 (N_10255,N_9916,N_9989);
nor U10256 (N_10256,N_9935,N_9896);
nand U10257 (N_10257,N_9707,N_9737);
and U10258 (N_10258,N_9801,N_9991);
xor U10259 (N_10259,N_9769,N_9602);
or U10260 (N_10260,N_9748,N_9823);
xnor U10261 (N_10261,N_9920,N_9756);
xor U10262 (N_10262,N_9615,N_9659);
xor U10263 (N_10263,N_9769,N_9863);
nor U10264 (N_10264,N_9636,N_9611);
nand U10265 (N_10265,N_9857,N_9684);
nor U10266 (N_10266,N_9745,N_9980);
or U10267 (N_10267,N_9782,N_9857);
and U10268 (N_10268,N_9649,N_9969);
xor U10269 (N_10269,N_9713,N_9745);
xor U10270 (N_10270,N_9890,N_9714);
xor U10271 (N_10271,N_9601,N_9869);
xor U10272 (N_10272,N_9891,N_9999);
nand U10273 (N_10273,N_9669,N_9814);
or U10274 (N_10274,N_9893,N_9965);
xnor U10275 (N_10275,N_9977,N_9741);
or U10276 (N_10276,N_9984,N_9751);
nand U10277 (N_10277,N_9628,N_9653);
and U10278 (N_10278,N_9632,N_9690);
and U10279 (N_10279,N_9802,N_9878);
or U10280 (N_10280,N_9863,N_9873);
or U10281 (N_10281,N_9705,N_9605);
nor U10282 (N_10282,N_9821,N_9627);
xor U10283 (N_10283,N_9787,N_9847);
nor U10284 (N_10284,N_9892,N_9983);
xnor U10285 (N_10285,N_9778,N_9684);
and U10286 (N_10286,N_9765,N_9738);
nand U10287 (N_10287,N_9948,N_9888);
nor U10288 (N_10288,N_9729,N_9892);
nand U10289 (N_10289,N_9978,N_9884);
or U10290 (N_10290,N_9627,N_9775);
nand U10291 (N_10291,N_9622,N_9602);
nand U10292 (N_10292,N_9674,N_9855);
xor U10293 (N_10293,N_9649,N_9848);
and U10294 (N_10294,N_9835,N_9603);
and U10295 (N_10295,N_9813,N_9765);
nand U10296 (N_10296,N_9829,N_9818);
xor U10297 (N_10297,N_9901,N_9894);
nand U10298 (N_10298,N_9626,N_9784);
nand U10299 (N_10299,N_9697,N_9823);
or U10300 (N_10300,N_9618,N_9695);
and U10301 (N_10301,N_9771,N_9726);
or U10302 (N_10302,N_9732,N_9627);
or U10303 (N_10303,N_9917,N_9780);
nor U10304 (N_10304,N_9658,N_9670);
and U10305 (N_10305,N_9858,N_9625);
or U10306 (N_10306,N_9840,N_9953);
nor U10307 (N_10307,N_9731,N_9846);
or U10308 (N_10308,N_9849,N_9616);
or U10309 (N_10309,N_9823,N_9760);
xor U10310 (N_10310,N_9931,N_9831);
or U10311 (N_10311,N_9716,N_9870);
or U10312 (N_10312,N_9803,N_9652);
nand U10313 (N_10313,N_9718,N_9654);
nor U10314 (N_10314,N_9966,N_9672);
and U10315 (N_10315,N_9843,N_9876);
nor U10316 (N_10316,N_9631,N_9824);
nand U10317 (N_10317,N_9982,N_9722);
or U10318 (N_10318,N_9921,N_9604);
or U10319 (N_10319,N_9861,N_9866);
xnor U10320 (N_10320,N_9787,N_9744);
or U10321 (N_10321,N_9970,N_9746);
and U10322 (N_10322,N_9709,N_9708);
and U10323 (N_10323,N_9829,N_9678);
or U10324 (N_10324,N_9662,N_9727);
nor U10325 (N_10325,N_9921,N_9687);
nand U10326 (N_10326,N_9646,N_9855);
and U10327 (N_10327,N_9945,N_9955);
nor U10328 (N_10328,N_9743,N_9975);
xnor U10329 (N_10329,N_9685,N_9644);
xor U10330 (N_10330,N_9622,N_9650);
nor U10331 (N_10331,N_9976,N_9929);
nand U10332 (N_10332,N_9755,N_9904);
nor U10333 (N_10333,N_9895,N_9902);
or U10334 (N_10334,N_9983,N_9894);
and U10335 (N_10335,N_9964,N_9785);
and U10336 (N_10336,N_9865,N_9778);
nand U10337 (N_10337,N_9624,N_9700);
or U10338 (N_10338,N_9747,N_9969);
xnor U10339 (N_10339,N_9779,N_9949);
nand U10340 (N_10340,N_9649,N_9799);
xor U10341 (N_10341,N_9754,N_9941);
or U10342 (N_10342,N_9850,N_9655);
nor U10343 (N_10343,N_9653,N_9926);
nor U10344 (N_10344,N_9735,N_9794);
nand U10345 (N_10345,N_9944,N_9667);
nor U10346 (N_10346,N_9609,N_9768);
nand U10347 (N_10347,N_9824,N_9652);
nor U10348 (N_10348,N_9662,N_9665);
or U10349 (N_10349,N_9843,N_9630);
or U10350 (N_10350,N_9871,N_9657);
xnor U10351 (N_10351,N_9683,N_9702);
and U10352 (N_10352,N_9652,N_9675);
nor U10353 (N_10353,N_9697,N_9628);
nand U10354 (N_10354,N_9845,N_9920);
nand U10355 (N_10355,N_9852,N_9731);
and U10356 (N_10356,N_9604,N_9654);
or U10357 (N_10357,N_9855,N_9789);
and U10358 (N_10358,N_9795,N_9850);
nor U10359 (N_10359,N_9706,N_9699);
xnor U10360 (N_10360,N_9880,N_9794);
xor U10361 (N_10361,N_9600,N_9812);
nand U10362 (N_10362,N_9780,N_9768);
or U10363 (N_10363,N_9675,N_9888);
nor U10364 (N_10364,N_9705,N_9609);
xor U10365 (N_10365,N_9683,N_9757);
and U10366 (N_10366,N_9867,N_9711);
nor U10367 (N_10367,N_9964,N_9632);
and U10368 (N_10368,N_9689,N_9697);
or U10369 (N_10369,N_9997,N_9822);
nand U10370 (N_10370,N_9605,N_9715);
and U10371 (N_10371,N_9708,N_9935);
nand U10372 (N_10372,N_9880,N_9906);
nand U10373 (N_10373,N_9875,N_9911);
nor U10374 (N_10374,N_9799,N_9783);
nor U10375 (N_10375,N_9845,N_9769);
xor U10376 (N_10376,N_9835,N_9992);
nand U10377 (N_10377,N_9676,N_9793);
xor U10378 (N_10378,N_9865,N_9677);
nor U10379 (N_10379,N_9986,N_9931);
or U10380 (N_10380,N_9819,N_9669);
xor U10381 (N_10381,N_9776,N_9613);
nand U10382 (N_10382,N_9791,N_9918);
xor U10383 (N_10383,N_9653,N_9899);
and U10384 (N_10384,N_9813,N_9686);
nor U10385 (N_10385,N_9854,N_9899);
and U10386 (N_10386,N_9684,N_9780);
nand U10387 (N_10387,N_9713,N_9651);
nor U10388 (N_10388,N_9935,N_9919);
nor U10389 (N_10389,N_9789,N_9864);
nor U10390 (N_10390,N_9632,N_9775);
or U10391 (N_10391,N_9834,N_9844);
and U10392 (N_10392,N_9876,N_9722);
and U10393 (N_10393,N_9696,N_9884);
xor U10394 (N_10394,N_9706,N_9691);
or U10395 (N_10395,N_9766,N_9872);
and U10396 (N_10396,N_9623,N_9651);
xnor U10397 (N_10397,N_9666,N_9854);
and U10398 (N_10398,N_9644,N_9915);
and U10399 (N_10399,N_9773,N_9774);
xor U10400 (N_10400,N_10337,N_10158);
or U10401 (N_10401,N_10372,N_10336);
or U10402 (N_10402,N_10246,N_10174);
nand U10403 (N_10403,N_10308,N_10284);
or U10404 (N_10404,N_10026,N_10213);
nand U10405 (N_10405,N_10115,N_10369);
nand U10406 (N_10406,N_10389,N_10041);
nand U10407 (N_10407,N_10097,N_10101);
or U10408 (N_10408,N_10128,N_10143);
nand U10409 (N_10409,N_10069,N_10286);
or U10410 (N_10410,N_10098,N_10083);
xnor U10411 (N_10411,N_10334,N_10192);
nand U10412 (N_10412,N_10347,N_10253);
nor U10413 (N_10413,N_10385,N_10200);
nand U10414 (N_10414,N_10323,N_10298);
xnor U10415 (N_10415,N_10395,N_10359);
nor U10416 (N_10416,N_10289,N_10208);
or U10417 (N_10417,N_10032,N_10022);
xnor U10418 (N_10418,N_10079,N_10147);
nor U10419 (N_10419,N_10312,N_10166);
or U10420 (N_10420,N_10126,N_10081);
nand U10421 (N_10421,N_10309,N_10038);
nor U10422 (N_10422,N_10316,N_10145);
and U10423 (N_10423,N_10295,N_10074);
or U10424 (N_10424,N_10018,N_10182);
xor U10425 (N_10425,N_10155,N_10057);
xor U10426 (N_10426,N_10184,N_10288);
nand U10427 (N_10427,N_10193,N_10102);
and U10428 (N_10428,N_10090,N_10072);
and U10429 (N_10429,N_10037,N_10362);
nor U10430 (N_10430,N_10168,N_10133);
nand U10431 (N_10431,N_10394,N_10346);
nor U10432 (N_10432,N_10159,N_10358);
nand U10433 (N_10433,N_10297,N_10196);
nor U10434 (N_10434,N_10290,N_10396);
or U10435 (N_10435,N_10172,N_10361);
nor U10436 (N_10436,N_10356,N_10380);
nand U10437 (N_10437,N_10390,N_10229);
and U10438 (N_10438,N_10164,N_10398);
or U10439 (N_10439,N_10215,N_10244);
xnor U10440 (N_10440,N_10017,N_10034);
nor U10441 (N_10441,N_10315,N_10342);
nand U10442 (N_10442,N_10139,N_10241);
nand U10443 (N_10443,N_10082,N_10216);
nor U10444 (N_10444,N_10392,N_10219);
or U10445 (N_10445,N_10066,N_10170);
or U10446 (N_10446,N_10043,N_10094);
or U10447 (N_10447,N_10360,N_10189);
xnor U10448 (N_10448,N_10169,N_10258);
nand U10449 (N_10449,N_10077,N_10096);
nor U10450 (N_10450,N_10171,N_10131);
and U10451 (N_10451,N_10203,N_10059);
or U10452 (N_10452,N_10020,N_10012);
nor U10453 (N_10453,N_10248,N_10245);
and U10454 (N_10454,N_10270,N_10095);
xnor U10455 (N_10455,N_10089,N_10302);
xor U10456 (N_10456,N_10156,N_10365);
nand U10457 (N_10457,N_10324,N_10035);
xor U10458 (N_10458,N_10052,N_10354);
or U10459 (N_10459,N_10019,N_10209);
or U10460 (N_10460,N_10186,N_10294);
and U10461 (N_10461,N_10195,N_10344);
nand U10462 (N_10462,N_10242,N_10153);
nand U10463 (N_10463,N_10254,N_10296);
nand U10464 (N_10464,N_10125,N_10163);
and U10465 (N_10465,N_10278,N_10367);
nor U10466 (N_10466,N_10050,N_10279);
nor U10467 (N_10467,N_10224,N_10055);
nor U10468 (N_10468,N_10188,N_10007);
or U10469 (N_10469,N_10107,N_10104);
and U10470 (N_10470,N_10024,N_10013);
and U10471 (N_10471,N_10060,N_10363);
nor U10472 (N_10472,N_10048,N_10259);
nand U10473 (N_10473,N_10078,N_10280);
nor U10474 (N_10474,N_10162,N_10165);
or U10475 (N_10475,N_10393,N_10322);
or U10476 (N_10476,N_10268,N_10185);
nand U10477 (N_10477,N_10267,N_10181);
xnor U10478 (N_10478,N_10148,N_10004);
and U10479 (N_10479,N_10223,N_10033);
nand U10480 (N_10480,N_10202,N_10029);
or U10481 (N_10481,N_10087,N_10343);
and U10482 (N_10482,N_10122,N_10300);
xor U10483 (N_10483,N_10371,N_10157);
or U10484 (N_10484,N_10311,N_10199);
and U10485 (N_10485,N_10063,N_10333);
nand U10486 (N_10486,N_10282,N_10243);
nor U10487 (N_10487,N_10330,N_10210);
nand U10488 (N_10488,N_10136,N_10387);
xor U10489 (N_10489,N_10044,N_10218);
xor U10490 (N_10490,N_10002,N_10046);
xor U10491 (N_10491,N_10092,N_10221);
nand U10492 (N_10492,N_10368,N_10146);
or U10493 (N_10493,N_10255,N_10240);
and U10494 (N_10494,N_10379,N_10320);
nand U10495 (N_10495,N_10226,N_10138);
and U10496 (N_10496,N_10269,N_10287);
and U10497 (N_10497,N_10349,N_10008);
nand U10498 (N_10498,N_10326,N_10071);
nor U10499 (N_10499,N_10051,N_10124);
xor U10500 (N_10500,N_10023,N_10027);
nand U10501 (N_10501,N_10307,N_10137);
nor U10502 (N_10502,N_10317,N_10160);
nor U10503 (N_10503,N_10374,N_10187);
xor U10504 (N_10504,N_10212,N_10227);
nand U10505 (N_10505,N_10238,N_10119);
xnor U10506 (N_10506,N_10306,N_10266);
xnor U10507 (N_10507,N_10109,N_10014);
xnor U10508 (N_10508,N_10351,N_10388);
xor U10509 (N_10509,N_10257,N_10377);
xor U10510 (N_10510,N_10305,N_10304);
xor U10511 (N_10511,N_10299,N_10262);
or U10512 (N_10512,N_10353,N_10339);
and U10513 (N_10513,N_10025,N_10154);
nor U10514 (N_10514,N_10141,N_10001);
xor U10515 (N_10515,N_10039,N_10085);
and U10516 (N_10516,N_10194,N_10335);
nand U10517 (N_10517,N_10142,N_10263);
nand U10518 (N_10518,N_10237,N_10180);
or U10519 (N_10519,N_10381,N_10364);
and U10520 (N_10520,N_10178,N_10277);
nor U10521 (N_10521,N_10045,N_10283);
and U10522 (N_10522,N_10250,N_10161);
xnor U10523 (N_10523,N_10325,N_10175);
xor U10524 (N_10524,N_10274,N_10345);
or U10525 (N_10525,N_10061,N_10047);
xor U10526 (N_10526,N_10327,N_10129);
or U10527 (N_10527,N_10231,N_10005);
xor U10528 (N_10528,N_10127,N_10239);
or U10529 (N_10529,N_10016,N_10247);
nor U10530 (N_10530,N_10106,N_10073);
or U10531 (N_10531,N_10230,N_10121);
nor U10532 (N_10532,N_10350,N_10285);
and U10533 (N_10533,N_10273,N_10015);
xor U10534 (N_10534,N_10197,N_10201);
and U10535 (N_10535,N_10319,N_10233);
xnor U10536 (N_10536,N_10214,N_10293);
xnor U10537 (N_10537,N_10383,N_10217);
xnor U10538 (N_10538,N_10149,N_10384);
nand U10539 (N_10539,N_10318,N_10291);
nor U10540 (N_10540,N_10144,N_10204);
xor U10541 (N_10541,N_10112,N_10252);
and U10542 (N_10542,N_10100,N_10338);
nand U10543 (N_10543,N_10067,N_10151);
or U10544 (N_10544,N_10340,N_10190);
nor U10545 (N_10545,N_10140,N_10135);
and U10546 (N_10546,N_10275,N_10206);
nor U10547 (N_10547,N_10068,N_10150);
and U10548 (N_10548,N_10292,N_10232);
or U10549 (N_10549,N_10056,N_10006);
xor U10550 (N_10550,N_10321,N_10220);
nor U10551 (N_10551,N_10062,N_10028);
nor U10552 (N_10552,N_10234,N_10328);
xor U10553 (N_10553,N_10132,N_10003);
or U10554 (N_10554,N_10040,N_10103);
nor U10555 (N_10555,N_10386,N_10198);
and U10556 (N_10556,N_10167,N_10281);
nand U10557 (N_10557,N_10251,N_10370);
or U10558 (N_10558,N_10049,N_10348);
and U10559 (N_10559,N_10108,N_10355);
xnor U10560 (N_10560,N_10314,N_10009);
or U10561 (N_10561,N_10134,N_10260);
nand U10562 (N_10562,N_10352,N_10177);
and U10563 (N_10563,N_10152,N_10235);
nand U10564 (N_10564,N_10310,N_10375);
xor U10565 (N_10565,N_10091,N_10391);
and U10566 (N_10566,N_10021,N_10113);
and U10567 (N_10567,N_10114,N_10276);
and U10568 (N_10568,N_10225,N_10265);
nor U10569 (N_10569,N_10064,N_10123);
and U10570 (N_10570,N_10053,N_10130);
or U10571 (N_10571,N_10010,N_10031);
nand U10572 (N_10572,N_10211,N_10173);
or U10573 (N_10573,N_10331,N_10256);
or U10574 (N_10574,N_10093,N_10301);
nor U10575 (N_10575,N_10222,N_10341);
nand U10576 (N_10576,N_10249,N_10030);
nand U10577 (N_10577,N_10000,N_10118);
nand U10578 (N_10578,N_10272,N_10110);
nand U10579 (N_10579,N_10111,N_10176);
or U10580 (N_10580,N_10399,N_10382);
and U10581 (N_10581,N_10236,N_10084);
nor U10582 (N_10582,N_10373,N_10183);
nand U10583 (N_10583,N_10117,N_10088);
nand U10584 (N_10584,N_10076,N_10054);
nor U10585 (N_10585,N_10332,N_10329);
nand U10586 (N_10586,N_10080,N_10205);
nand U10587 (N_10587,N_10011,N_10036);
and U10588 (N_10588,N_10075,N_10366);
and U10589 (N_10589,N_10313,N_10116);
or U10590 (N_10590,N_10099,N_10179);
nor U10591 (N_10591,N_10042,N_10065);
nand U10592 (N_10592,N_10261,N_10058);
xor U10593 (N_10593,N_10105,N_10207);
or U10594 (N_10594,N_10303,N_10357);
and U10595 (N_10595,N_10120,N_10378);
or U10596 (N_10596,N_10397,N_10070);
or U10597 (N_10597,N_10376,N_10086);
and U10598 (N_10598,N_10191,N_10271);
nand U10599 (N_10599,N_10264,N_10228);
nand U10600 (N_10600,N_10118,N_10033);
and U10601 (N_10601,N_10225,N_10068);
nor U10602 (N_10602,N_10000,N_10262);
nor U10603 (N_10603,N_10053,N_10087);
or U10604 (N_10604,N_10100,N_10217);
or U10605 (N_10605,N_10337,N_10270);
nor U10606 (N_10606,N_10218,N_10382);
or U10607 (N_10607,N_10057,N_10253);
or U10608 (N_10608,N_10277,N_10371);
nor U10609 (N_10609,N_10115,N_10140);
and U10610 (N_10610,N_10007,N_10120);
xor U10611 (N_10611,N_10171,N_10382);
nand U10612 (N_10612,N_10272,N_10049);
nor U10613 (N_10613,N_10070,N_10097);
nor U10614 (N_10614,N_10239,N_10365);
nand U10615 (N_10615,N_10229,N_10358);
nor U10616 (N_10616,N_10277,N_10157);
and U10617 (N_10617,N_10384,N_10076);
nor U10618 (N_10618,N_10239,N_10186);
xor U10619 (N_10619,N_10242,N_10077);
nor U10620 (N_10620,N_10121,N_10340);
or U10621 (N_10621,N_10332,N_10086);
nor U10622 (N_10622,N_10180,N_10118);
nand U10623 (N_10623,N_10019,N_10052);
and U10624 (N_10624,N_10009,N_10082);
or U10625 (N_10625,N_10308,N_10162);
xor U10626 (N_10626,N_10304,N_10336);
and U10627 (N_10627,N_10272,N_10289);
xor U10628 (N_10628,N_10032,N_10177);
and U10629 (N_10629,N_10386,N_10121);
xor U10630 (N_10630,N_10034,N_10014);
nand U10631 (N_10631,N_10288,N_10085);
nand U10632 (N_10632,N_10312,N_10117);
xor U10633 (N_10633,N_10061,N_10121);
xor U10634 (N_10634,N_10272,N_10324);
or U10635 (N_10635,N_10145,N_10055);
or U10636 (N_10636,N_10018,N_10212);
nor U10637 (N_10637,N_10207,N_10095);
xnor U10638 (N_10638,N_10188,N_10041);
nor U10639 (N_10639,N_10294,N_10236);
xor U10640 (N_10640,N_10397,N_10148);
and U10641 (N_10641,N_10364,N_10185);
nor U10642 (N_10642,N_10061,N_10019);
and U10643 (N_10643,N_10334,N_10361);
nand U10644 (N_10644,N_10207,N_10318);
and U10645 (N_10645,N_10152,N_10356);
or U10646 (N_10646,N_10096,N_10314);
xor U10647 (N_10647,N_10273,N_10000);
nand U10648 (N_10648,N_10166,N_10274);
or U10649 (N_10649,N_10114,N_10135);
or U10650 (N_10650,N_10384,N_10394);
nor U10651 (N_10651,N_10026,N_10268);
nand U10652 (N_10652,N_10321,N_10117);
xnor U10653 (N_10653,N_10120,N_10322);
nor U10654 (N_10654,N_10148,N_10262);
nor U10655 (N_10655,N_10094,N_10297);
or U10656 (N_10656,N_10301,N_10221);
or U10657 (N_10657,N_10048,N_10072);
and U10658 (N_10658,N_10017,N_10201);
and U10659 (N_10659,N_10129,N_10259);
xnor U10660 (N_10660,N_10270,N_10286);
nor U10661 (N_10661,N_10145,N_10092);
nor U10662 (N_10662,N_10287,N_10068);
nor U10663 (N_10663,N_10032,N_10107);
xor U10664 (N_10664,N_10121,N_10077);
xor U10665 (N_10665,N_10276,N_10149);
or U10666 (N_10666,N_10233,N_10006);
nor U10667 (N_10667,N_10376,N_10036);
nor U10668 (N_10668,N_10162,N_10386);
nand U10669 (N_10669,N_10046,N_10028);
and U10670 (N_10670,N_10103,N_10136);
xor U10671 (N_10671,N_10122,N_10101);
and U10672 (N_10672,N_10385,N_10030);
nand U10673 (N_10673,N_10166,N_10344);
nand U10674 (N_10674,N_10028,N_10191);
nand U10675 (N_10675,N_10043,N_10183);
and U10676 (N_10676,N_10075,N_10209);
and U10677 (N_10677,N_10123,N_10237);
and U10678 (N_10678,N_10183,N_10329);
and U10679 (N_10679,N_10238,N_10236);
nor U10680 (N_10680,N_10297,N_10247);
nand U10681 (N_10681,N_10391,N_10247);
and U10682 (N_10682,N_10061,N_10298);
nor U10683 (N_10683,N_10183,N_10021);
nand U10684 (N_10684,N_10041,N_10390);
and U10685 (N_10685,N_10087,N_10044);
and U10686 (N_10686,N_10250,N_10007);
xnor U10687 (N_10687,N_10347,N_10074);
xnor U10688 (N_10688,N_10365,N_10314);
nor U10689 (N_10689,N_10218,N_10094);
nand U10690 (N_10690,N_10095,N_10268);
or U10691 (N_10691,N_10269,N_10179);
xnor U10692 (N_10692,N_10159,N_10041);
and U10693 (N_10693,N_10034,N_10095);
nand U10694 (N_10694,N_10187,N_10159);
nor U10695 (N_10695,N_10155,N_10243);
or U10696 (N_10696,N_10000,N_10396);
xnor U10697 (N_10697,N_10377,N_10222);
nor U10698 (N_10698,N_10014,N_10278);
or U10699 (N_10699,N_10381,N_10186);
or U10700 (N_10700,N_10236,N_10132);
nor U10701 (N_10701,N_10279,N_10268);
nor U10702 (N_10702,N_10286,N_10131);
xor U10703 (N_10703,N_10104,N_10287);
and U10704 (N_10704,N_10296,N_10001);
or U10705 (N_10705,N_10376,N_10135);
and U10706 (N_10706,N_10025,N_10394);
or U10707 (N_10707,N_10390,N_10110);
nor U10708 (N_10708,N_10123,N_10272);
nand U10709 (N_10709,N_10151,N_10128);
and U10710 (N_10710,N_10071,N_10177);
and U10711 (N_10711,N_10254,N_10078);
nor U10712 (N_10712,N_10327,N_10309);
xor U10713 (N_10713,N_10064,N_10220);
xor U10714 (N_10714,N_10369,N_10109);
nor U10715 (N_10715,N_10229,N_10257);
nor U10716 (N_10716,N_10232,N_10115);
and U10717 (N_10717,N_10034,N_10080);
nor U10718 (N_10718,N_10380,N_10136);
xnor U10719 (N_10719,N_10281,N_10264);
xnor U10720 (N_10720,N_10010,N_10127);
nand U10721 (N_10721,N_10177,N_10096);
or U10722 (N_10722,N_10089,N_10059);
xnor U10723 (N_10723,N_10234,N_10189);
nand U10724 (N_10724,N_10240,N_10168);
xor U10725 (N_10725,N_10310,N_10373);
xnor U10726 (N_10726,N_10233,N_10257);
nor U10727 (N_10727,N_10315,N_10387);
nand U10728 (N_10728,N_10388,N_10143);
nor U10729 (N_10729,N_10334,N_10024);
or U10730 (N_10730,N_10316,N_10291);
nor U10731 (N_10731,N_10036,N_10332);
or U10732 (N_10732,N_10242,N_10304);
and U10733 (N_10733,N_10291,N_10383);
nand U10734 (N_10734,N_10123,N_10285);
or U10735 (N_10735,N_10373,N_10079);
and U10736 (N_10736,N_10230,N_10124);
or U10737 (N_10737,N_10196,N_10232);
or U10738 (N_10738,N_10012,N_10177);
or U10739 (N_10739,N_10042,N_10020);
or U10740 (N_10740,N_10293,N_10308);
and U10741 (N_10741,N_10318,N_10351);
or U10742 (N_10742,N_10233,N_10377);
nand U10743 (N_10743,N_10160,N_10299);
nor U10744 (N_10744,N_10081,N_10003);
nor U10745 (N_10745,N_10079,N_10214);
xnor U10746 (N_10746,N_10361,N_10376);
or U10747 (N_10747,N_10129,N_10054);
xnor U10748 (N_10748,N_10027,N_10297);
nand U10749 (N_10749,N_10264,N_10040);
or U10750 (N_10750,N_10293,N_10376);
xnor U10751 (N_10751,N_10066,N_10065);
xnor U10752 (N_10752,N_10276,N_10009);
nor U10753 (N_10753,N_10117,N_10191);
and U10754 (N_10754,N_10223,N_10277);
nor U10755 (N_10755,N_10042,N_10054);
or U10756 (N_10756,N_10307,N_10302);
or U10757 (N_10757,N_10119,N_10011);
or U10758 (N_10758,N_10088,N_10048);
nor U10759 (N_10759,N_10377,N_10019);
xnor U10760 (N_10760,N_10158,N_10194);
nand U10761 (N_10761,N_10205,N_10311);
nor U10762 (N_10762,N_10237,N_10044);
nand U10763 (N_10763,N_10032,N_10096);
nor U10764 (N_10764,N_10103,N_10375);
and U10765 (N_10765,N_10003,N_10376);
nand U10766 (N_10766,N_10289,N_10298);
or U10767 (N_10767,N_10047,N_10260);
nor U10768 (N_10768,N_10244,N_10324);
xnor U10769 (N_10769,N_10161,N_10099);
and U10770 (N_10770,N_10132,N_10335);
nor U10771 (N_10771,N_10199,N_10152);
nand U10772 (N_10772,N_10181,N_10011);
nand U10773 (N_10773,N_10215,N_10206);
nor U10774 (N_10774,N_10348,N_10083);
or U10775 (N_10775,N_10228,N_10184);
or U10776 (N_10776,N_10375,N_10104);
and U10777 (N_10777,N_10289,N_10040);
and U10778 (N_10778,N_10230,N_10182);
and U10779 (N_10779,N_10049,N_10394);
xnor U10780 (N_10780,N_10138,N_10140);
or U10781 (N_10781,N_10010,N_10216);
xnor U10782 (N_10782,N_10021,N_10003);
and U10783 (N_10783,N_10329,N_10260);
nor U10784 (N_10784,N_10108,N_10089);
and U10785 (N_10785,N_10183,N_10155);
or U10786 (N_10786,N_10344,N_10280);
xnor U10787 (N_10787,N_10330,N_10033);
xnor U10788 (N_10788,N_10264,N_10033);
nor U10789 (N_10789,N_10276,N_10029);
nor U10790 (N_10790,N_10270,N_10223);
and U10791 (N_10791,N_10173,N_10106);
or U10792 (N_10792,N_10068,N_10394);
nor U10793 (N_10793,N_10146,N_10192);
nor U10794 (N_10794,N_10363,N_10177);
nand U10795 (N_10795,N_10367,N_10104);
nand U10796 (N_10796,N_10011,N_10009);
nand U10797 (N_10797,N_10029,N_10003);
or U10798 (N_10798,N_10094,N_10319);
nor U10799 (N_10799,N_10019,N_10016);
or U10800 (N_10800,N_10466,N_10665);
nor U10801 (N_10801,N_10799,N_10548);
or U10802 (N_10802,N_10745,N_10472);
or U10803 (N_10803,N_10423,N_10620);
nor U10804 (N_10804,N_10737,N_10404);
nor U10805 (N_10805,N_10497,N_10516);
and U10806 (N_10806,N_10743,N_10792);
and U10807 (N_10807,N_10483,N_10447);
xnor U10808 (N_10808,N_10781,N_10616);
nand U10809 (N_10809,N_10568,N_10793);
xnor U10810 (N_10810,N_10601,N_10409);
nand U10811 (N_10811,N_10473,N_10580);
nand U10812 (N_10812,N_10612,N_10509);
xor U10813 (N_10813,N_10740,N_10408);
or U10814 (N_10814,N_10564,N_10689);
nor U10815 (N_10815,N_10632,N_10557);
and U10816 (N_10816,N_10419,N_10566);
nor U10817 (N_10817,N_10546,N_10436);
xor U10818 (N_10818,N_10674,N_10687);
nor U10819 (N_10819,N_10695,N_10673);
or U10820 (N_10820,N_10592,N_10782);
xor U10821 (N_10821,N_10463,N_10403);
and U10822 (N_10822,N_10505,N_10727);
xnor U10823 (N_10823,N_10449,N_10575);
or U10824 (N_10824,N_10607,N_10427);
nor U10825 (N_10825,N_10615,N_10595);
or U10826 (N_10826,N_10424,N_10726);
and U10827 (N_10827,N_10597,N_10747);
xnor U10828 (N_10828,N_10414,N_10433);
and U10829 (N_10829,N_10650,N_10780);
or U10830 (N_10830,N_10406,N_10678);
xnor U10831 (N_10831,N_10554,N_10664);
or U10832 (N_10832,N_10738,N_10559);
xor U10833 (N_10833,N_10587,N_10659);
or U10834 (N_10834,N_10759,N_10776);
or U10835 (N_10835,N_10670,N_10426);
and U10836 (N_10836,N_10733,N_10448);
nor U10837 (N_10837,N_10774,N_10555);
nand U10838 (N_10838,N_10490,N_10688);
nand U10839 (N_10839,N_10736,N_10489);
and U10840 (N_10840,N_10734,N_10491);
nor U10841 (N_10841,N_10567,N_10437);
nor U10842 (N_10842,N_10703,N_10715);
or U10843 (N_10843,N_10502,N_10639);
or U10844 (N_10844,N_10493,N_10467);
nand U10845 (N_10845,N_10712,N_10479);
nor U10846 (N_10846,N_10698,N_10750);
and U10847 (N_10847,N_10637,N_10589);
nand U10848 (N_10848,N_10649,N_10513);
and U10849 (N_10849,N_10422,N_10662);
and U10850 (N_10850,N_10600,N_10768);
nor U10851 (N_10851,N_10481,N_10432);
and U10852 (N_10852,N_10465,N_10443);
and U10853 (N_10853,N_10638,N_10631);
nand U10854 (N_10854,N_10605,N_10458);
or U10855 (N_10855,N_10484,N_10746);
nand U10856 (N_10856,N_10748,N_10783);
nor U10857 (N_10857,N_10681,N_10648);
xnor U10858 (N_10858,N_10462,N_10453);
xor U10859 (N_10859,N_10586,N_10635);
nand U10860 (N_10860,N_10794,N_10428);
nor U10861 (N_10861,N_10769,N_10573);
nor U10862 (N_10862,N_10593,N_10732);
nor U10863 (N_10863,N_10524,N_10450);
and U10864 (N_10864,N_10477,N_10588);
or U10865 (N_10865,N_10417,N_10470);
nand U10866 (N_10866,N_10692,N_10496);
or U10867 (N_10867,N_10617,N_10739);
and U10868 (N_10868,N_10621,N_10603);
xor U10869 (N_10869,N_10552,N_10645);
nor U10870 (N_10870,N_10412,N_10511);
and U10871 (N_10871,N_10656,N_10787);
nor U10872 (N_10872,N_10435,N_10576);
or U10873 (N_10873,N_10789,N_10682);
and U10874 (N_10874,N_10723,N_10476);
or U10875 (N_10875,N_10651,N_10475);
or U10876 (N_10876,N_10558,N_10766);
nand U10877 (N_10877,N_10722,N_10400);
xor U10878 (N_10878,N_10791,N_10492);
nand U10879 (N_10879,N_10411,N_10684);
xor U10880 (N_10880,N_10760,N_10533);
xor U10881 (N_10881,N_10425,N_10613);
and U10882 (N_10882,N_10752,N_10440);
nand U10883 (N_10883,N_10728,N_10551);
nor U10884 (N_10884,N_10764,N_10667);
xor U10885 (N_10885,N_10630,N_10691);
nand U10886 (N_10886,N_10507,N_10503);
xor U10887 (N_10887,N_10754,N_10522);
and U10888 (N_10888,N_10619,N_10498);
xor U10889 (N_10889,N_10699,N_10536);
and U10890 (N_10890,N_10686,N_10707);
and U10891 (N_10891,N_10625,N_10478);
nand U10892 (N_10892,N_10622,N_10790);
nor U10893 (N_10893,N_10401,N_10755);
nor U10894 (N_10894,N_10626,N_10742);
and U10895 (N_10895,N_10532,N_10501);
nor U10896 (N_10896,N_10685,N_10461);
nand U10897 (N_10897,N_10429,N_10714);
or U10898 (N_10898,N_10506,N_10430);
and U10899 (N_10899,N_10758,N_10713);
xor U10900 (N_10900,N_10494,N_10556);
nand U10901 (N_10901,N_10640,N_10633);
and U10902 (N_10902,N_10526,N_10629);
xor U10903 (N_10903,N_10721,N_10679);
nand U10904 (N_10904,N_10534,N_10569);
or U10905 (N_10905,N_10416,N_10460);
nand U10906 (N_10906,N_10661,N_10608);
or U10907 (N_10907,N_10761,N_10598);
nand U10908 (N_10908,N_10653,N_10624);
and U10909 (N_10909,N_10451,N_10610);
and U10910 (N_10910,N_10459,N_10495);
or U10911 (N_10911,N_10562,N_10700);
xor U10912 (N_10912,N_10599,N_10675);
xor U10913 (N_10913,N_10521,N_10413);
and U10914 (N_10914,N_10464,N_10751);
and U10915 (N_10915,N_10690,N_10488);
nor U10916 (N_10916,N_10770,N_10796);
or U10917 (N_10917,N_10410,N_10441);
or U10918 (N_10918,N_10765,N_10518);
nand U10919 (N_10919,N_10545,N_10654);
nand U10920 (N_10920,N_10560,N_10510);
or U10921 (N_10921,N_10402,N_10535);
xor U10922 (N_10922,N_10655,N_10749);
and U10923 (N_10923,N_10701,N_10515);
xor U10924 (N_10924,N_10676,N_10704);
and U10925 (N_10925,N_10549,N_10596);
xnor U10926 (N_10926,N_10731,N_10779);
nor U10927 (N_10927,N_10643,N_10778);
and U10928 (N_10928,N_10657,N_10572);
and U10929 (N_10929,N_10717,N_10594);
or U10930 (N_10930,N_10585,N_10531);
or U10931 (N_10931,N_10504,N_10438);
and U10932 (N_10932,N_10777,N_10672);
nand U10933 (N_10933,N_10445,N_10762);
and U10934 (N_10934,N_10487,N_10718);
nor U10935 (N_10935,N_10540,N_10647);
xor U10936 (N_10936,N_10538,N_10454);
or U10937 (N_10937,N_10604,N_10628);
or U10938 (N_10938,N_10456,N_10602);
xor U10939 (N_10939,N_10544,N_10431);
nor U10940 (N_10940,N_10702,N_10668);
nand U10941 (N_10941,N_10452,N_10627);
nor U10942 (N_10942,N_10652,N_10486);
nor U10943 (N_10943,N_10710,N_10418);
nor U10944 (N_10944,N_10663,N_10442);
nor U10945 (N_10945,N_10694,N_10658);
xor U10946 (N_10946,N_10517,N_10756);
nand U10947 (N_10947,N_10553,N_10798);
or U10948 (N_10948,N_10581,N_10720);
or U10949 (N_10949,N_10611,N_10542);
or U10950 (N_10950,N_10623,N_10767);
nand U10951 (N_10951,N_10706,N_10405);
nor U10952 (N_10952,N_10669,N_10499);
nand U10953 (N_10953,N_10457,N_10529);
or U10954 (N_10954,N_10579,N_10530);
and U10955 (N_10955,N_10570,N_10512);
nor U10956 (N_10956,N_10471,N_10527);
nor U10957 (N_10957,N_10729,N_10583);
or U10958 (N_10958,N_10520,N_10683);
and U10959 (N_10959,N_10671,N_10480);
and U10960 (N_10960,N_10709,N_10716);
xor U10961 (N_10961,N_10636,N_10420);
and U10962 (N_10962,N_10724,N_10577);
or U10963 (N_10963,N_10757,N_10641);
nor U10964 (N_10964,N_10693,N_10725);
or U10965 (N_10965,N_10609,N_10474);
and U10966 (N_10966,N_10711,N_10618);
nor U10967 (N_10967,N_10574,N_10439);
and U10968 (N_10968,N_10696,N_10784);
nor U10969 (N_10969,N_10508,N_10571);
xor U10970 (N_10970,N_10705,N_10642);
xnor U10971 (N_10971,N_10500,N_10519);
or U10972 (N_10972,N_10775,N_10550);
or U10973 (N_10973,N_10415,N_10614);
nand U10974 (N_10974,N_10735,N_10646);
or U10975 (N_10975,N_10785,N_10590);
or U10976 (N_10976,N_10773,N_10525);
nor U10977 (N_10977,N_10578,N_10455);
or U10978 (N_10978,N_10547,N_10719);
xor U10979 (N_10979,N_10772,N_10528);
xor U10980 (N_10980,N_10680,N_10565);
nand U10981 (N_10981,N_10537,N_10666);
and U10982 (N_10982,N_10543,N_10514);
nor U10983 (N_10983,N_10591,N_10797);
and U10984 (N_10984,N_10697,N_10744);
xor U10985 (N_10985,N_10582,N_10771);
nor U10986 (N_10986,N_10730,N_10753);
nor U10987 (N_10987,N_10660,N_10421);
nand U10988 (N_10988,N_10606,N_10485);
and U10989 (N_10989,N_10561,N_10468);
xor U10990 (N_10990,N_10469,N_10763);
xor U10991 (N_10991,N_10708,N_10584);
xnor U10992 (N_10992,N_10407,N_10644);
nor U10993 (N_10993,N_10741,N_10786);
nor U10994 (N_10994,N_10539,N_10563);
xor U10995 (N_10995,N_10788,N_10446);
xnor U10996 (N_10996,N_10795,N_10523);
xnor U10997 (N_10997,N_10677,N_10541);
nor U10998 (N_10998,N_10634,N_10482);
xnor U10999 (N_10999,N_10444,N_10434);
and U11000 (N_11000,N_10670,N_10518);
nor U11001 (N_11001,N_10713,N_10442);
nor U11002 (N_11002,N_10625,N_10744);
nand U11003 (N_11003,N_10732,N_10799);
or U11004 (N_11004,N_10762,N_10469);
nand U11005 (N_11005,N_10637,N_10639);
xnor U11006 (N_11006,N_10543,N_10689);
nor U11007 (N_11007,N_10401,N_10708);
xor U11008 (N_11008,N_10674,N_10738);
or U11009 (N_11009,N_10780,N_10693);
nor U11010 (N_11010,N_10674,N_10494);
or U11011 (N_11011,N_10612,N_10610);
and U11012 (N_11012,N_10671,N_10763);
or U11013 (N_11013,N_10794,N_10546);
nand U11014 (N_11014,N_10485,N_10400);
or U11015 (N_11015,N_10554,N_10403);
or U11016 (N_11016,N_10511,N_10755);
or U11017 (N_11017,N_10787,N_10680);
or U11018 (N_11018,N_10735,N_10473);
nor U11019 (N_11019,N_10705,N_10635);
and U11020 (N_11020,N_10776,N_10697);
xnor U11021 (N_11021,N_10552,N_10453);
nand U11022 (N_11022,N_10758,N_10608);
and U11023 (N_11023,N_10753,N_10638);
nand U11024 (N_11024,N_10714,N_10762);
xor U11025 (N_11025,N_10784,N_10583);
and U11026 (N_11026,N_10791,N_10639);
nand U11027 (N_11027,N_10472,N_10443);
or U11028 (N_11028,N_10731,N_10532);
xor U11029 (N_11029,N_10490,N_10752);
nand U11030 (N_11030,N_10753,N_10430);
nor U11031 (N_11031,N_10522,N_10684);
or U11032 (N_11032,N_10554,N_10542);
and U11033 (N_11033,N_10406,N_10745);
nor U11034 (N_11034,N_10628,N_10445);
and U11035 (N_11035,N_10556,N_10466);
or U11036 (N_11036,N_10411,N_10714);
nand U11037 (N_11037,N_10502,N_10524);
nor U11038 (N_11038,N_10479,N_10741);
nor U11039 (N_11039,N_10487,N_10401);
or U11040 (N_11040,N_10479,N_10562);
xnor U11041 (N_11041,N_10594,N_10543);
nand U11042 (N_11042,N_10780,N_10441);
nand U11043 (N_11043,N_10449,N_10599);
or U11044 (N_11044,N_10793,N_10629);
or U11045 (N_11045,N_10777,N_10402);
nand U11046 (N_11046,N_10622,N_10471);
xor U11047 (N_11047,N_10425,N_10701);
xor U11048 (N_11048,N_10527,N_10445);
nand U11049 (N_11049,N_10539,N_10567);
nand U11050 (N_11050,N_10774,N_10711);
and U11051 (N_11051,N_10438,N_10446);
xnor U11052 (N_11052,N_10745,N_10711);
xor U11053 (N_11053,N_10754,N_10752);
nand U11054 (N_11054,N_10627,N_10523);
and U11055 (N_11055,N_10758,N_10442);
xnor U11056 (N_11056,N_10722,N_10635);
nand U11057 (N_11057,N_10614,N_10501);
nand U11058 (N_11058,N_10449,N_10701);
xor U11059 (N_11059,N_10497,N_10465);
or U11060 (N_11060,N_10602,N_10585);
nand U11061 (N_11061,N_10746,N_10598);
and U11062 (N_11062,N_10738,N_10730);
and U11063 (N_11063,N_10560,N_10413);
xor U11064 (N_11064,N_10714,N_10651);
nand U11065 (N_11065,N_10649,N_10505);
nor U11066 (N_11066,N_10696,N_10594);
or U11067 (N_11067,N_10500,N_10627);
nor U11068 (N_11068,N_10710,N_10632);
xnor U11069 (N_11069,N_10786,N_10419);
or U11070 (N_11070,N_10430,N_10709);
nor U11071 (N_11071,N_10459,N_10527);
xor U11072 (N_11072,N_10411,N_10671);
or U11073 (N_11073,N_10458,N_10685);
nor U11074 (N_11074,N_10686,N_10505);
nor U11075 (N_11075,N_10575,N_10440);
or U11076 (N_11076,N_10493,N_10445);
or U11077 (N_11077,N_10727,N_10473);
xnor U11078 (N_11078,N_10412,N_10748);
nand U11079 (N_11079,N_10793,N_10547);
and U11080 (N_11080,N_10726,N_10427);
xor U11081 (N_11081,N_10613,N_10523);
nand U11082 (N_11082,N_10675,N_10534);
or U11083 (N_11083,N_10681,N_10646);
and U11084 (N_11084,N_10676,N_10736);
or U11085 (N_11085,N_10763,N_10492);
or U11086 (N_11086,N_10791,N_10431);
and U11087 (N_11087,N_10709,N_10446);
nor U11088 (N_11088,N_10590,N_10573);
and U11089 (N_11089,N_10477,N_10616);
nand U11090 (N_11090,N_10536,N_10515);
nand U11091 (N_11091,N_10589,N_10442);
and U11092 (N_11092,N_10606,N_10448);
and U11093 (N_11093,N_10673,N_10655);
nand U11094 (N_11094,N_10626,N_10770);
or U11095 (N_11095,N_10431,N_10479);
nand U11096 (N_11096,N_10431,N_10480);
nand U11097 (N_11097,N_10412,N_10478);
xor U11098 (N_11098,N_10555,N_10717);
and U11099 (N_11099,N_10576,N_10752);
nand U11100 (N_11100,N_10445,N_10566);
nor U11101 (N_11101,N_10724,N_10414);
nor U11102 (N_11102,N_10493,N_10521);
nand U11103 (N_11103,N_10722,N_10589);
or U11104 (N_11104,N_10475,N_10499);
xor U11105 (N_11105,N_10529,N_10638);
or U11106 (N_11106,N_10530,N_10768);
and U11107 (N_11107,N_10441,N_10419);
and U11108 (N_11108,N_10600,N_10734);
nor U11109 (N_11109,N_10564,N_10451);
and U11110 (N_11110,N_10568,N_10681);
and U11111 (N_11111,N_10707,N_10790);
or U11112 (N_11112,N_10623,N_10739);
and U11113 (N_11113,N_10672,N_10421);
or U11114 (N_11114,N_10656,N_10633);
nand U11115 (N_11115,N_10667,N_10531);
and U11116 (N_11116,N_10691,N_10468);
or U11117 (N_11117,N_10590,N_10560);
xor U11118 (N_11118,N_10653,N_10673);
or U11119 (N_11119,N_10780,N_10601);
and U11120 (N_11120,N_10578,N_10698);
and U11121 (N_11121,N_10567,N_10729);
xor U11122 (N_11122,N_10641,N_10440);
or U11123 (N_11123,N_10776,N_10430);
or U11124 (N_11124,N_10574,N_10580);
or U11125 (N_11125,N_10438,N_10674);
xnor U11126 (N_11126,N_10673,N_10685);
or U11127 (N_11127,N_10416,N_10535);
and U11128 (N_11128,N_10543,N_10617);
nand U11129 (N_11129,N_10633,N_10755);
or U11130 (N_11130,N_10590,N_10622);
xnor U11131 (N_11131,N_10769,N_10477);
nor U11132 (N_11132,N_10695,N_10679);
nand U11133 (N_11133,N_10437,N_10733);
or U11134 (N_11134,N_10480,N_10694);
and U11135 (N_11135,N_10783,N_10502);
xor U11136 (N_11136,N_10542,N_10606);
and U11137 (N_11137,N_10516,N_10440);
xnor U11138 (N_11138,N_10422,N_10776);
nor U11139 (N_11139,N_10732,N_10638);
and U11140 (N_11140,N_10666,N_10727);
xor U11141 (N_11141,N_10713,N_10696);
xor U11142 (N_11142,N_10518,N_10663);
xnor U11143 (N_11143,N_10763,N_10478);
xnor U11144 (N_11144,N_10590,N_10519);
or U11145 (N_11145,N_10752,N_10775);
xor U11146 (N_11146,N_10526,N_10592);
and U11147 (N_11147,N_10432,N_10420);
xor U11148 (N_11148,N_10691,N_10724);
or U11149 (N_11149,N_10776,N_10431);
and U11150 (N_11150,N_10549,N_10681);
or U11151 (N_11151,N_10615,N_10673);
nand U11152 (N_11152,N_10581,N_10445);
or U11153 (N_11153,N_10690,N_10481);
nor U11154 (N_11154,N_10527,N_10669);
nand U11155 (N_11155,N_10418,N_10409);
xnor U11156 (N_11156,N_10500,N_10451);
nand U11157 (N_11157,N_10573,N_10705);
or U11158 (N_11158,N_10430,N_10792);
nor U11159 (N_11159,N_10489,N_10563);
nor U11160 (N_11160,N_10772,N_10755);
xor U11161 (N_11161,N_10409,N_10583);
or U11162 (N_11162,N_10662,N_10515);
or U11163 (N_11163,N_10642,N_10755);
or U11164 (N_11164,N_10744,N_10598);
nor U11165 (N_11165,N_10517,N_10664);
xnor U11166 (N_11166,N_10572,N_10626);
nand U11167 (N_11167,N_10787,N_10675);
nand U11168 (N_11168,N_10611,N_10756);
nand U11169 (N_11169,N_10777,N_10553);
xnor U11170 (N_11170,N_10728,N_10463);
and U11171 (N_11171,N_10708,N_10647);
nand U11172 (N_11172,N_10569,N_10768);
or U11173 (N_11173,N_10570,N_10629);
xor U11174 (N_11174,N_10459,N_10713);
nand U11175 (N_11175,N_10707,N_10699);
or U11176 (N_11176,N_10633,N_10657);
nor U11177 (N_11177,N_10540,N_10576);
or U11178 (N_11178,N_10665,N_10425);
xor U11179 (N_11179,N_10762,N_10656);
xor U11180 (N_11180,N_10464,N_10536);
xor U11181 (N_11181,N_10597,N_10406);
nor U11182 (N_11182,N_10788,N_10577);
and U11183 (N_11183,N_10498,N_10657);
xnor U11184 (N_11184,N_10535,N_10658);
nor U11185 (N_11185,N_10541,N_10737);
or U11186 (N_11186,N_10505,N_10638);
nand U11187 (N_11187,N_10515,N_10499);
nand U11188 (N_11188,N_10672,N_10417);
xor U11189 (N_11189,N_10796,N_10518);
nand U11190 (N_11190,N_10544,N_10542);
or U11191 (N_11191,N_10654,N_10565);
and U11192 (N_11192,N_10775,N_10477);
or U11193 (N_11193,N_10464,N_10720);
xnor U11194 (N_11194,N_10609,N_10705);
nor U11195 (N_11195,N_10596,N_10765);
nor U11196 (N_11196,N_10755,N_10590);
nand U11197 (N_11197,N_10635,N_10664);
and U11198 (N_11198,N_10497,N_10788);
nor U11199 (N_11199,N_10740,N_10715);
and U11200 (N_11200,N_10952,N_11089);
or U11201 (N_11201,N_11096,N_10923);
or U11202 (N_11202,N_11189,N_10858);
xor U11203 (N_11203,N_11047,N_11155);
and U11204 (N_11204,N_11146,N_10967);
and U11205 (N_11205,N_10913,N_10899);
nor U11206 (N_11206,N_10903,N_10963);
and U11207 (N_11207,N_10974,N_10922);
nor U11208 (N_11208,N_11012,N_11185);
nand U11209 (N_11209,N_11053,N_11070);
or U11210 (N_11210,N_11084,N_10984);
or U11211 (N_11211,N_11137,N_10805);
nand U11212 (N_11212,N_11027,N_11003);
nand U11213 (N_11213,N_11190,N_11001);
nor U11214 (N_11214,N_11095,N_10990);
or U11215 (N_11215,N_11107,N_11090);
or U11216 (N_11216,N_11011,N_10890);
or U11217 (N_11217,N_10883,N_10991);
and U11218 (N_11218,N_11044,N_11031);
nand U11219 (N_11219,N_10848,N_10989);
or U11220 (N_11220,N_11197,N_11111);
xor U11221 (N_11221,N_11079,N_11145);
or U11222 (N_11222,N_11166,N_11103);
xnor U11223 (N_11223,N_10813,N_11061);
xor U11224 (N_11224,N_11159,N_10821);
nand U11225 (N_11225,N_11083,N_10933);
nor U11226 (N_11226,N_10867,N_10915);
xor U11227 (N_11227,N_10983,N_10981);
and U11228 (N_11228,N_11177,N_11151);
or U11229 (N_11229,N_10947,N_10893);
and U11230 (N_11230,N_10875,N_11033);
xor U11231 (N_11231,N_11040,N_10908);
nor U11232 (N_11232,N_11086,N_10855);
nor U11233 (N_11233,N_10907,N_11029);
or U11234 (N_11234,N_10801,N_11057);
nor U11235 (N_11235,N_11100,N_10942);
and U11236 (N_11236,N_10824,N_11091);
xor U11237 (N_11237,N_10844,N_11039);
and U11238 (N_11238,N_11056,N_11052);
or U11239 (N_11239,N_10940,N_10959);
and U11240 (N_11240,N_10862,N_11023);
xor U11241 (N_11241,N_10819,N_10803);
nor U11242 (N_11242,N_10955,N_11182);
xnor U11243 (N_11243,N_11188,N_11119);
xor U11244 (N_11244,N_10982,N_10970);
xor U11245 (N_11245,N_11180,N_10904);
nand U11246 (N_11246,N_11055,N_11051);
and U11247 (N_11247,N_11148,N_10887);
or U11248 (N_11248,N_11198,N_11002);
nand U11249 (N_11249,N_10934,N_10889);
nand U11250 (N_11250,N_11192,N_11058);
and U11251 (N_11251,N_10835,N_11021);
or U11252 (N_11252,N_11004,N_11127);
nor U11253 (N_11253,N_10920,N_10895);
and U11254 (N_11254,N_11115,N_11042);
nand U11255 (N_11255,N_11160,N_10857);
and U11256 (N_11256,N_10918,N_11175);
nor U11257 (N_11257,N_11035,N_10914);
nand U11258 (N_11258,N_11026,N_10976);
nand U11259 (N_11259,N_11196,N_10971);
xor U11260 (N_11260,N_10810,N_10945);
or U11261 (N_11261,N_11123,N_10850);
or U11262 (N_11262,N_11135,N_11105);
and U11263 (N_11263,N_10825,N_10870);
and U11264 (N_11264,N_11109,N_11036);
and U11265 (N_11265,N_11114,N_11032);
xor U11266 (N_11266,N_11049,N_10832);
nor U11267 (N_11267,N_11161,N_11162);
xnor U11268 (N_11268,N_11149,N_11007);
nand U11269 (N_11269,N_10897,N_10972);
or U11270 (N_11270,N_10996,N_11138);
or U11271 (N_11271,N_10938,N_10891);
and U11272 (N_11272,N_10849,N_10854);
or U11273 (N_11273,N_10878,N_10941);
and U11274 (N_11274,N_10969,N_11064);
or U11275 (N_11275,N_10826,N_11076);
or U11276 (N_11276,N_11018,N_11173);
nand U11277 (N_11277,N_11099,N_10912);
or U11278 (N_11278,N_10900,N_11092);
or U11279 (N_11279,N_11120,N_10980);
and U11280 (N_11280,N_11010,N_11179);
and U11281 (N_11281,N_10806,N_11122);
and U11282 (N_11282,N_10874,N_11030);
xor U11283 (N_11283,N_11067,N_10808);
nor U11284 (N_11284,N_10979,N_10929);
xnor U11285 (N_11285,N_10815,N_11020);
xor U11286 (N_11286,N_11153,N_11069);
xor U11287 (N_11287,N_11174,N_10919);
nand U11288 (N_11288,N_11104,N_10954);
nand U11289 (N_11289,N_11106,N_11037);
nand U11290 (N_11290,N_11006,N_11134);
xnor U11291 (N_11291,N_11050,N_11184);
xor U11292 (N_11292,N_10968,N_11195);
and U11293 (N_11293,N_10881,N_11028);
xor U11294 (N_11294,N_11139,N_10909);
nand U11295 (N_11295,N_10966,N_11169);
and U11296 (N_11296,N_11087,N_10902);
nor U11297 (N_11297,N_11140,N_10856);
or U11298 (N_11298,N_10987,N_11063);
nor U11299 (N_11299,N_10859,N_10910);
nor U11300 (N_11300,N_11014,N_10841);
nor U11301 (N_11301,N_10949,N_11022);
nor U11302 (N_11302,N_10994,N_10992);
nor U11303 (N_11303,N_10939,N_11136);
nor U11304 (N_11304,N_10818,N_11019);
and U11305 (N_11305,N_10911,N_11009);
or U11306 (N_11306,N_11129,N_11116);
nand U11307 (N_11307,N_10937,N_10995);
nand U11308 (N_11308,N_11117,N_10827);
nand U11309 (N_11309,N_10960,N_10864);
or U11310 (N_11310,N_11034,N_11025);
and U11311 (N_11311,N_10879,N_11194);
xnor U11312 (N_11312,N_10814,N_10965);
nand U11313 (N_11313,N_11038,N_10873);
and U11314 (N_11314,N_10950,N_11152);
nor U11315 (N_11315,N_10868,N_10901);
nor U11316 (N_11316,N_11059,N_10928);
xnor U11317 (N_11317,N_11163,N_11143);
and U11318 (N_11318,N_11000,N_11072);
nor U11319 (N_11319,N_10834,N_11112);
or U11320 (N_11320,N_11172,N_11156);
or U11321 (N_11321,N_10964,N_11132);
xnor U11322 (N_11322,N_10880,N_10829);
or U11323 (N_11323,N_11073,N_11071);
or U11324 (N_11324,N_11158,N_11082);
xor U11325 (N_11325,N_11126,N_10894);
or U11326 (N_11326,N_10885,N_10946);
nand U11327 (N_11327,N_10988,N_11017);
or U11328 (N_11328,N_10986,N_11150);
xnor U11329 (N_11329,N_10816,N_10927);
xnor U11330 (N_11330,N_11154,N_10957);
xor U11331 (N_11331,N_10936,N_11142);
nor U11332 (N_11332,N_11013,N_11077);
xnor U11333 (N_11333,N_11125,N_10905);
and U11334 (N_11334,N_10842,N_10943);
or U11335 (N_11335,N_11054,N_10853);
and U11336 (N_11336,N_10930,N_11081);
nor U11337 (N_11337,N_11165,N_11102);
nand U11338 (N_11338,N_11098,N_11066);
nand U11339 (N_11339,N_10944,N_10993);
nand U11340 (N_11340,N_10863,N_11178);
nor U11341 (N_11341,N_10807,N_10998);
and U11342 (N_11342,N_11130,N_10869);
xnor U11343 (N_11343,N_10932,N_10876);
nand U11344 (N_11344,N_10871,N_11168);
xor U11345 (N_11345,N_11016,N_10877);
nor U11346 (N_11346,N_10837,N_11124);
or U11347 (N_11347,N_11097,N_11147);
or U11348 (N_11348,N_10811,N_11110);
xnor U11349 (N_11349,N_10861,N_10843);
xnor U11350 (N_11350,N_10962,N_10925);
xor U11351 (N_11351,N_10898,N_10978);
and U11352 (N_11352,N_11118,N_10906);
xnor U11353 (N_11353,N_11108,N_10948);
nor U11354 (N_11354,N_11170,N_10833);
and U11355 (N_11355,N_11068,N_11121);
nor U11356 (N_11356,N_11133,N_11176);
xnor U11357 (N_11357,N_11060,N_10958);
nor U11358 (N_11358,N_11141,N_11074);
nand U11359 (N_11359,N_11113,N_10823);
xor U11360 (N_11360,N_11183,N_10884);
xnor U11361 (N_11361,N_11088,N_10830);
and U11362 (N_11362,N_11065,N_10896);
xnor U11363 (N_11363,N_10985,N_10997);
xor U11364 (N_11364,N_10851,N_10838);
and U11365 (N_11365,N_11167,N_10866);
or U11366 (N_11366,N_11101,N_10804);
xnor U11367 (N_11367,N_11085,N_10951);
xor U11368 (N_11368,N_11024,N_11181);
and U11369 (N_11369,N_10809,N_11093);
nand U11370 (N_11370,N_11075,N_11144);
or U11371 (N_11371,N_11078,N_11080);
and U11372 (N_11372,N_11046,N_11171);
nand U11373 (N_11373,N_10935,N_11131);
xnor U11374 (N_11374,N_10973,N_11062);
xnor U11375 (N_11375,N_10931,N_10845);
xor U11376 (N_11376,N_11015,N_11005);
and U11377 (N_11377,N_10800,N_10892);
xor U11378 (N_11378,N_10860,N_10846);
and U11379 (N_11379,N_11193,N_10812);
nand U11380 (N_11380,N_10999,N_11186);
nor U11381 (N_11381,N_10977,N_11045);
nor U11382 (N_11382,N_10802,N_10924);
nor U11383 (N_11383,N_11041,N_11199);
nand U11384 (N_11384,N_10921,N_10847);
and U11385 (N_11385,N_10852,N_10926);
nand U11386 (N_11386,N_10882,N_10840);
nor U11387 (N_11387,N_10839,N_10831);
and U11388 (N_11388,N_11164,N_10820);
or U11389 (N_11389,N_10817,N_10888);
nand U11390 (N_11390,N_10975,N_10836);
nand U11391 (N_11391,N_10886,N_11157);
nand U11392 (N_11392,N_10956,N_11187);
and U11393 (N_11393,N_10916,N_11094);
nor U11394 (N_11394,N_11043,N_10828);
and U11395 (N_11395,N_11008,N_10953);
xnor U11396 (N_11396,N_10822,N_10961);
nand U11397 (N_11397,N_11048,N_10865);
or U11398 (N_11398,N_11128,N_11191);
or U11399 (N_11399,N_10872,N_10917);
or U11400 (N_11400,N_11169,N_10948);
nor U11401 (N_11401,N_10884,N_10814);
nand U11402 (N_11402,N_10946,N_11164);
xnor U11403 (N_11403,N_10971,N_10975);
nor U11404 (N_11404,N_10854,N_11177);
nor U11405 (N_11405,N_10819,N_11042);
nor U11406 (N_11406,N_11090,N_11190);
nand U11407 (N_11407,N_10909,N_11084);
nor U11408 (N_11408,N_10923,N_10926);
nor U11409 (N_11409,N_11120,N_11153);
xor U11410 (N_11410,N_11077,N_11192);
xnor U11411 (N_11411,N_11145,N_11121);
xnor U11412 (N_11412,N_11160,N_10821);
and U11413 (N_11413,N_10817,N_11078);
and U11414 (N_11414,N_11118,N_11087);
or U11415 (N_11415,N_11031,N_10947);
nor U11416 (N_11416,N_10809,N_11011);
and U11417 (N_11417,N_11183,N_11156);
and U11418 (N_11418,N_11078,N_10915);
or U11419 (N_11419,N_10831,N_10859);
nand U11420 (N_11420,N_11043,N_10948);
nor U11421 (N_11421,N_11085,N_10945);
nand U11422 (N_11422,N_11086,N_11071);
nand U11423 (N_11423,N_11112,N_11029);
nand U11424 (N_11424,N_10906,N_10889);
nand U11425 (N_11425,N_10865,N_10920);
or U11426 (N_11426,N_10884,N_11113);
or U11427 (N_11427,N_11061,N_11106);
nor U11428 (N_11428,N_11085,N_10833);
or U11429 (N_11429,N_10898,N_10818);
xnor U11430 (N_11430,N_10812,N_11174);
or U11431 (N_11431,N_10888,N_11197);
or U11432 (N_11432,N_10897,N_10864);
and U11433 (N_11433,N_11043,N_10921);
nand U11434 (N_11434,N_11146,N_10940);
nor U11435 (N_11435,N_11034,N_10925);
or U11436 (N_11436,N_10954,N_11025);
nor U11437 (N_11437,N_10938,N_11123);
and U11438 (N_11438,N_11052,N_10923);
or U11439 (N_11439,N_11001,N_11015);
xnor U11440 (N_11440,N_10951,N_10822);
or U11441 (N_11441,N_11073,N_11191);
and U11442 (N_11442,N_11176,N_11081);
and U11443 (N_11443,N_10841,N_11077);
and U11444 (N_11444,N_11014,N_10881);
xor U11445 (N_11445,N_10817,N_11027);
xor U11446 (N_11446,N_11127,N_11028);
and U11447 (N_11447,N_10854,N_10995);
or U11448 (N_11448,N_10843,N_10807);
nand U11449 (N_11449,N_11140,N_11038);
and U11450 (N_11450,N_10991,N_11178);
nor U11451 (N_11451,N_11198,N_10835);
nand U11452 (N_11452,N_11092,N_10971);
xor U11453 (N_11453,N_11025,N_11063);
xnor U11454 (N_11454,N_10927,N_11114);
and U11455 (N_11455,N_11184,N_10912);
nand U11456 (N_11456,N_10918,N_10895);
and U11457 (N_11457,N_10976,N_11041);
nor U11458 (N_11458,N_11145,N_11055);
xnor U11459 (N_11459,N_11108,N_11015);
and U11460 (N_11460,N_11062,N_10990);
xor U11461 (N_11461,N_11074,N_10838);
nand U11462 (N_11462,N_10874,N_11032);
or U11463 (N_11463,N_11092,N_10855);
nor U11464 (N_11464,N_11002,N_11132);
nand U11465 (N_11465,N_11098,N_10871);
and U11466 (N_11466,N_11046,N_10943);
nor U11467 (N_11467,N_11121,N_10907);
or U11468 (N_11468,N_10898,N_10948);
nand U11469 (N_11469,N_10814,N_11146);
xnor U11470 (N_11470,N_11132,N_10897);
nor U11471 (N_11471,N_11152,N_11077);
or U11472 (N_11472,N_10940,N_11112);
or U11473 (N_11473,N_10986,N_11199);
or U11474 (N_11474,N_10865,N_10968);
and U11475 (N_11475,N_11139,N_11011);
nor U11476 (N_11476,N_10837,N_10813);
nor U11477 (N_11477,N_10822,N_11062);
or U11478 (N_11478,N_11173,N_11081);
nor U11479 (N_11479,N_10835,N_10938);
or U11480 (N_11480,N_11027,N_11094);
or U11481 (N_11481,N_10880,N_10926);
and U11482 (N_11482,N_10841,N_11098);
and U11483 (N_11483,N_11005,N_10812);
or U11484 (N_11484,N_11166,N_11177);
nor U11485 (N_11485,N_11117,N_11041);
or U11486 (N_11486,N_10923,N_10932);
xor U11487 (N_11487,N_10828,N_11148);
nor U11488 (N_11488,N_11065,N_10927);
nor U11489 (N_11489,N_10970,N_11042);
nor U11490 (N_11490,N_10922,N_11076);
and U11491 (N_11491,N_11198,N_10996);
and U11492 (N_11492,N_11059,N_10976);
nand U11493 (N_11493,N_11022,N_10887);
or U11494 (N_11494,N_11051,N_11087);
and U11495 (N_11495,N_10976,N_11089);
nor U11496 (N_11496,N_10978,N_10860);
nand U11497 (N_11497,N_11030,N_10905);
nand U11498 (N_11498,N_10817,N_11051);
nand U11499 (N_11499,N_11184,N_11189);
nor U11500 (N_11500,N_11124,N_11169);
nand U11501 (N_11501,N_11000,N_11029);
xnor U11502 (N_11502,N_10855,N_10820);
or U11503 (N_11503,N_11129,N_11119);
xor U11504 (N_11504,N_10964,N_11063);
xnor U11505 (N_11505,N_11027,N_10926);
and U11506 (N_11506,N_10869,N_11078);
xnor U11507 (N_11507,N_11109,N_11130);
nor U11508 (N_11508,N_10874,N_11138);
nand U11509 (N_11509,N_11138,N_11136);
xnor U11510 (N_11510,N_11083,N_10914);
and U11511 (N_11511,N_11179,N_11095);
xnor U11512 (N_11512,N_10894,N_11049);
nand U11513 (N_11513,N_10860,N_10863);
nor U11514 (N_11514,N_10800,N_11002);
xnor U11515 (N_11515,N_10891,N_10968);
nand U11516 (N_11516,N_11053,N_10819);
or U11517 (N_11517,N_10844,N_10939);
nor U11518 (N_11518,N_11017,N_11010);
and U11519 (N_11519,N_11060,N_11133);
and U11520 (N_11520,N_10893,N_10812);
nor U11521 (N_11521,N_11175,N_10800);
xor U11522 (N_11522,N_11180,N_11052);
nor U11523 (N_11523,N_10845,N_11039);
nand U11524 (N_11524,N_11061,N_11056);
nor U11525 (N_11525,N_10995,N_11131);
nor U11526 (N_11526,N_10920,N_11098);
nor U11527 (N_11527,N_11038,N_11177);
nor U11528 (N_11528,N_11177,N_10856);
and U11529 (N_11529,N_11025,N_10819);
nand U11530 (N_11530,N_10904,N_10947);
nor U11531 (N_11531,N_11195,N_10957);
nand U11532 (N_11532,N_11011,N_10888);
nor U11533 (N_11533,N_10843,N_10986);
nand U11534 (N_11534,N_11128,N_10866);
and U11535 (N_11535,N_11096,N_11092);
nand U11536 (N_11536,N_11059,N_10978);
or U11537 (N_11537,N_10938,N_10874);
or U11538 (N_11538,N_10948,N_10830);
nor U11539 (N_11539,N_11022,N_10900);
xor U11540 (N_11540,N_10841,N_11031);
nand U11541 (N_11541,N_11020,N_10807);
xor U11542 (N_11542,N_11078,N_11001);
and U11543 (N_11543,N_10928,N_11053);
nor U11544 (N_11544,N_11092,N_10977);
and U11545 (N_11545,N_11124,N_10875);
nand U11546 (N_11546,N_10957,N_11090);
and U11547 (N_11547,N_11106,N_10922);
nand U11548 (N_11548,N_10808,N_11111);
and U11549 (N_11549,N_11180,N_10960);
xnor U11550 (N_11550,N_10944,N_10898);
nand U11551 (N_11551,N_10950,N_11100);
and U11552 (N_11552,N_10906,N_10876);
or U11553 (N_11553,N_11111,N_11149);
and U11554 (N_11554,N_11017,N_11023);
nand U11555 (N_11555,N_11030,N_10809);
or U11556 (N_11556,N_11198,N_10927);
and U11557 (N_11557,N_10816,N_10969);
xor U11558 (N_11558,N_10880,N_11103);
or U11559 (N_11559,N_10942,N_11148);
nor U11560 (N_11560,N_10960,N_10812);
xor U11561 (N_11561,N_10984,N_11066);
and U11562 (N_11562,N_10914,N_11070);
xnor U11563 (N_11563,N_11063,N_11045);
and U11564 (N_11564,N_10807,N_10917);
nand U11565 (N_11565,N_11137,N_11121);
nor U11566 (N_11566,N_11023,N_11071);
or U11567 (N_11567,N_11162,N_11038);
nand U11568 (N_11568,N_11048,N_10899);
xnor U11569 (N_11569,N_10940,N_10868);
and U11570 (N_11570,N_10984,N_10977);
and U11571 (N_11571,N_11150,N_11155);
nor U11572 (N_11572,N_10824,N_11113);
and U11573 (N_11573,N_10886,N_11126);
nor U11574 (N_11574,N_10981,N_10975);
xor U11575 (N_11575,N_11109,N_10918);
nor U11576 (N_11576,N_10930,N_10868);
nand U11577 (N_11577,N_10924,N_11159);
nor U11578 (N_11578,N_10869,N_10942);
xor U11579 (N_11579,N_10981,N_11001);
nor U11580 (N_11580,N_10926,N_11091);
xnor U11581 (N_11581,N_10996,N_10977);
nand U11582 (N_11582,N_10947,N_11119);
xnor U11583 (N_11583,N_11192,N_11089);
nand U11584 (N_11584,N_10813,N_10998);
nor U11585 (N_11585,N_10804,N_10909);
nand U11586 (N_11586,N_11120,N_10982);
or U11587 (N_11587,N_10826,N_11100);
and U11588 (N_11588,N_11049,N_10960);
nand U11589 (N_11589,N_11133,N_10882);
xor U11590 (N_11590,N_10919,N_10929);
or U11591 (N_11591,N_11177,N_11088);
and U11592 (N_11592,N_10900,N_10950);
nor U11593 (N_11593,N_11193,N_11100);
or U11594 (N_11594,N_10935,N_11158);
and U11595 (N_11595,N_10975,N_10926);
xor U11596 (N_11596,N_11078,N_11014);
and U11597 (N_11597,N_10835,N_11003);
or U11598 (N_11598,N_11112,N_10950);
and U11599 (N_11599,N_11132,N_10845);
and U11600 (N_11600,N_11387,N_11507);
or U11601 (N_11601,N_11218,N_11456);
or U11602 (N_11602,N_11212,N_11516);
nor U11603 (N_11603,N_11541,N_11531);
or U11604 (N_11604,N_11463,N_11572);
nor U11605 (N_11605,N_11328,N_11564);
xor U11606 (N_11606,N_11331,N_11332);
and U11607 (N_11607,N_11539,N_11496);
xnor U11608 (N_11608,N_11549,N_11380);
xor U11609 (N_11609,N_11390,N_11426);
or U11610 (N_11610,N_11499,N_11268);
nand U11611 (N_11611,N_11545,N_11478);
nand U11612 (N_11612,N_11480,N_11430);
xor U11613 (N_11613,N_11391,N_11299);
and U11614 (N_11614,N_11568,N_11479);
or U11615 (N_11615,N_11360,N_11276);
xnor U11616 (N_11616,N_11442,N_11384);
xor U11617 (N_11617,N_11469,N_11425);
xor U11618 (N_11618,N_11403,N_11528);
or U11619 (N_11619,N_11309,N_11215);
or U11620 (N_11620,N_11301,N_11586);
nor U11621 (N_11621,N_11407,N_11295);
or U11622 (N_11622,N_11352,N_11418);
xnor U11623 (N_11623,N_11548,N_11251);
nor U11624 (N_11624,N_11433,N_11252);
or U11625 (N_11625,N_11269,N_11560);
or U11626 (N_11626,N_11209,N_11312);
nor U11627 (N_11627,N_11376,N_11386);
or U11628 (N_11628,N_11534,N_11382);
nand U11629 (N_11629,N_11226,N_11282);
or U11630 (N_11630,N_11562,N_11489);
or U11631 (N_11631,N_11434,N_11570);
xor U11632 (N_11632,N_11363,N_11513);
nand U11633 (N_11633,N_11359,N_11241);
and U11634 (N_11634,N_11378,N_11428);
and U11635 (N_11635,N_11599,N_11298);
or U11636 (N_11636,N_11581,N_11579);
or U11637 (N_11637,N_11449,N_11592);
and U11638 (N_11638,N_11294,N_11419);
and U11639 (N_11639,N_11244,N_11341);
or U11640 (N_11640,N_11435,N_11556);
xor U11641 (N_11641,N_11321,N_11367);
and U11642 (N_11642,N_11221,N_11240);
xnor U11643 (N_11643,N_11527,N_11211);
nor U11644 (N_11644,N_11559,N_11490);
nor U11645 (N_11645,N_11389,N_11373);
nand U11646 (N_11646,N_11492,N_11342);
xnor U11647 (N_11647,N_11291,N_11219);
or U11648 (N_11648,N_11439,N_11566);
or U11649 (N_11649,N_11246,N_11208);
xnor U11650 (N_11650,N_11544,N_11473);
or U11651 (N_11651,N_11420,N_11506);
or U11652 (N_11652,N_11510,N_11257);
nand U11653 (N_11653,N_11200,N_11595);
nor U11654 (N_11654,N_11394,N_11271);
and U11655 (N_11655,N_11227,N_11228);
nand U11656 (N_11656,N_11577,N_11340);
and U11657 (N_11657,N_11333,N_11455);
and U11658 (N_11658,N_11265,N_11270);
and U11659 (N_11659,N_11542,N_11488);
or U11660 (N_11660,N_11225,N_11578);
or U11661 (N_11661,N_11329,N_11565);
xor U11662 (N_11662,N_11432,N_11302);
nand U11663 (N_11663,N_11520,N_11346);
xor U11664 (N_11664,N_11279,N_11445);
or U11665 (N_11665,N_11247,N_11524);
nand U11666 (N_11666,N_11512,N_11344);
xnor U11667 (N_11667,N_11514,N_11235);
and U11668 (N_11668,N_11258,N_11347);
nor U11669 (N_11669,N_11417,N_11261);
nand U11670 (N_11670,N_11438,N_11300);
nand U11671 (N_11671,N_11594,N_11323);
xor U11672 (N_11672,N_11451,N_11374);
and U11673 (N_11673,N_11508,N_11343);
or U11674 (N_11674,N_11204,N_11547);
or U11675 (N_11675,N_11305,N_11237);
nand U11676 (N_11676,N_11307,N_11290);
nand U11677 (N_11677,N_11248,N_11551);
and U11678 (N_11678,N_11379,N_11518);
nor U11679 (N_11679,N_11362,N_11475);
xor U11680 (N_11680,N_11303,N_11459);
and U11681 (N_11681,N_11392,N_11327);
nor U11682 (N_11682,N_11519,N_11447);
nand U11683 (N_11683,N_11535,N_11530);
nand U11684 (N_11684,N_11325,N_11210);
nand U11685 (N_11685,N_11231,N_11207);
nor U11686 (N_11686,N_11414,N_11203);
and U11687 (N_11687,N_11423,N_11311);
or U11688 (N_11688,N_11486,N_11259);
and U11689 (N_11689,N_11267,N_11297);
and U11690 (N_11690,N_11366,N_11404);
xnor U11691 (N_11691,N_11324,N_11316);
or U11692 (N_11692,N_11584,N_11401);
and U11693 (N_11693,N_11277,N_11427);
or U11694 (N_11694,N_11571,N_11422);
nand U11695 (N_11695,N_11353,N_11448);
or U11696 (N_11696,N_11233,N_11381);
nor U11697 (N_11697,N_11457,N_11483);
or U11698 (N_11698,N_11306,N_11273);
xor U11699 (N_11699,N_11375,N_11262);
and U11700 (N_11700,N_11266,N_11310);
or U11701 (N_11701,N_11576,N_11393);
xor U11702 (N_11702,N_11356,N_11440);
or U11703 (N_11703,N_11256,N_11536);
xnor U11704 (N_11704,N_11216,N_11320);
and U11705 (N_11705,N_11365,N_11245);
nand U11706 (N_11706,N_11337,N_11253);
nand U11707 (N_11707,N_11283,N_11238);
nand U11708 (N_11708,N_11398,N_11357);
xor U11709 (N_11709,N_11526,N_11355);
and U11710 (N_11710,N_11591,N_11339);
nor U11711 (N_11711,N_11400,N_11315);
and U11712 (N_11712,N_11491,N_11288);
nor U11713 (N_11713,N_11285,N_11250);
or U11714 (N_11714,N_11412,N_11354);
and U11715 (N_11715,N_11350,N_11361);
xnor U11716 (N_11716,N_11487,N_11505);
xnor U11717 (N_11717,N_11550,N_11567);
nor U11718 (N_11718,N_11585,N_11351);
xnor U11719 (N_11719,N_11263,N_11569);
nor U11720 (N_11720,N_11255,N_11460);
xnor U11721 (N_11721,N_11415,N_11485);
nand U11722 (N_11722,N_11590,N_11254);
nand U11723 (N_11723,N_11436,N_11540);
nor U11724 (N_11724,N_11217,N_11429);
or U11725 (N_11725,N_11532,N_11575);
xor U11726 (N_11726,N_11249,N_11336);
or U11727 (N_11727,N_11424,N_11206);
or U11728 (N_11728,N_11474,N_11214);
nand U11729 (N_11729,N_11476,N_11509);
and U11730 (N_11730,N_11421,N_11552);
xor U11731 (N_11731,N_11533,N_11236);
nand U11732 (N_11732,N_11468,N_11561);
xnor U11733 (N_11733,N_11296,N_11588);
xnor U11734 (N_11734,N_11322,N_11213);
xor U11735 (N_11735,N_11477,N_11289);
or U11736 (N_11736,N_11287,N_11593);
and U11737 (N_11737,N_11345,N_11493);
nand U11738 (N_11738,N_11280,N_11314);
xor U11739 (N_11739,N_11563,N_11454);
nand U11740 (N_11740,N_11453,N_11371);
xnor U11741 (N_11741,N_11443,N_11502);
xor U11742 (N_11742,N_11281,N_11441);
or U11743 (N_11743,N_11555,N_11348);
xnor U11744 (N_11744,N_11402,N_11222);
xor U11745 (N_11745,N_11272,N_11239);
nand U11746 (N_11746,N_11501,N_11597);
nand U11747 (N_11747,N_11464,N_11525);
or U11748 (N_11748,N_11446,N_11395);
nand U11749 (N_11749,N_11465,N_11368);
xor U11750 (N_11750,N_11462,N_11529);
xor U11751 (N_11751,N_11399,N_11292);
or U11752 (N_11752,N_11554,N_11405);
and U11753 (N_11753,N_11264,N_11515);
and U11754 (N_11754,N_11330,N_11408);
xor U11755 (N_11755,N_11369,N_11484);
nor U11756 (N_11756,N_11243,N_11431);
and U11757 (N_11757,N_11286,N_11284);
and U11758 (N_11758,N_11503,N_11543);
or U11759 (N_11759,N_11495,N_11504);
xor U11760 (N_11760,N_11260,N_11500);
xnor U11761 (N_11761,N_11582,N_11466);
nor U11762 (N_11762,N_11358,N_11293);
or U11763 (N_11763,N_11319,N_11234);
or U11764 (N_11764,N_11523,N_11229);
nand U11765 (N_11765,N_11553,N_11494);
and U11766 (N_11766,N_11372,N_11377);
nand U11767 (N_11767,N_11497,N_11230);
xor U11768 (N_11768,N_11558,N_11589);
or U11769 (N_11769,N_11383,N_11223);
and U11770 (N_11770,N_11202,N_11467);
nor U11771 (N_11771,N_11538,N_11482);
and U11772 (N_11772,N_11517,N_11557);
or U11773 (N_11773,N_11370,N_11587);
nand U11774 (N_11774,N_11452,N_11317);
nand U11775 (N_11775,N_11522,N_11470);
xor U11776 (N_11776,N_11413,N_11521);
and U11777 (N_11777,N_11511,N_11498);
or U11778 (N_11778,N_11349,N_11278);
nand U11779 (N_11779,N_11409,N_11334);
and U11780 (N_11780,N_11574,N_11232);
nor U11781 (N_11781,N_11308,N_11326);
xnor U11782 (N_11782,N_11437,N_11410);
xor U11783 (N_11783,N_11406,N_11546);
nand U11784 (N_11784,N_11205,N_11596);
nor U11785 (N_11785,N_11388,N_11313);
nor U11786 (N_11786,N_11338,N_11242);
nor U11787 (N_11787,N_11274,N_11583);
nand U11788 (N_11788,N_11364,N_11580);
and U11789 (N_11789,N_11275,N_11450);
nor U11790 (N_11790,N_11472,N_11411);
nor U11791 (N_11791,N_11537,N_11385);
and U11792 (N_11792,N_11220,N_11481);
nand U11793 (N_11793,N_11318,N_11471);
xor U11794 (N_11794,N_11458,N_11444);
nor U11795 (N_11795,N_11598,N_11201);
xor U11796 (N_11796,N_11416,N_11396);
nand U11797 (N_11797,N_11304,N_11397);
xor U11798 (N_11798,N_11573,N_11224);
xnor U11799 (N_11799,N_11335,N_11461);
nand U11800 (N_11800,N_11249,N_11397);
and U11801 (N_11801,N_11561,N_11438);
and U11802 (N_11802,N_11418,N_11498);
xnor U11803 (N_11803,N_11517,N_11414);
nand U11804 (N_11804,N_11517,N_11528);
nand U11805 (N_11805,N_11384,N_11471);
xnor U11806 (N_11806,N_11201,N_11255);
or U11807 (N_11807,N_11387,N_11392);
nand U11808 (N_11808,N_11465,N_11514);
or U11809 (N_11809,N_11412,N_11304);
nor U11810 (N_11810,N_11467,N_11469);
xnor U11811 (N_11811,N_11541,N_11564);
and U11812 (N_11812,N_11373,N_11203);
nand U11813 (N_11813,N_11222,N_11526);
nor U11814 (N_11814,N_11481,N_11215);
and U11815 (N_11815,N_11431,N_11562);
nand U11816 (N_11816,N_11321,N_11533);
nand U11817 (N_11817,N_11450,N_11469);
xnor U11818 (N_11818,N_11261,N_11446);
xor U11819 (N_11819,N_11288,N_11348);
xnor U11820 (N_11820,N_11473,N_11361);
nand U11821 (N_11821,N_11325,N_11233);
or U11822 (N_11822,N_11274,N_11251);
nand U11823 (N_11823,N_11239,N_11286);
xnor U11824 (N_11824,N_11545,N_11442);
or U11825 (N_11825,N_11208,N_11408);
nand U11826 (N_11826,N_11489,N_11414);
or U11827 (N_11827,N_11266,N_11398);
nand U11828 (N_11828,N_11429,N_11281);
and U11829 (N_11829,N_11310,N_11202);
xor U11830 (N_11830,N_11431,N_11484);
or U11831 (N_11831,N_11459,N_11274);
or U11832 (N_11832,N_11585,N_11208);
xor U11833 (N_11833,N_11230,N_11289);
and U11834 (N_11834,N_11543,N_11211);
and U11835 (N_11835,N_11515,N_11297);
nor U11836 (N_11836,N_11534,N_11451);
nand U11837 (N_11837,N_11415,N_11580);
xnor U11838 (N_11838,N_11356,N_11484);
xnor U11839 (N_11839,N_11542,N_11517);
xor U11840 (N_11840,N_11592,N_11415);
nor U11841 (N_11841,N_11417,N_11414);
nand U11842 (N_11842,N_11408,N_11215);
and U11843 (N_11843,N_11402,N_11581);
and U11844 (N_11844,N_11524,N_11460);
nand U11845 (N_11845,N_11575,N_11352);
nand U11846 (N_11846,N_11202,N_11332);
nor U11847 (N_11847,N_11516,N_11566);
nor U11848 (N_11848,N_11449,N_11203);
nor U11849 (N_11849,N_11255,N_11400);
or U11850 (N_11850,N_11539,N_11471);
nand U11851 (N_11851,N_11444,N_11244);
nand U11852 (N_11852,N_11453,N_11436);
nand U11853 (N_11853,N_11346,N_11483);
xor U11854 (N_11854,N_11436,N_11503);
xor U11855 (N_11855,N_11575,N_11300);
xor U11856 (N_11856,N_11519,N_11229);
and U11857 (N_11857,N_11430,N_11335);
and U11858 (N_11858,N_11499,N_11421);
nor U11859 (N_11859,N_11592,N_11377);
nor U11860 (N_11860,N_11524,N_11397);
or U11861 (N_11861,N_11439,N_11408);
or U11862 (N_11862,N_11258,N_11335);
xor U11863 (N_11863,N_11521,N_11327);
or U11864 (N_11864,N_11248,N_11453);
nand U11865 (N_11865,N_11541,N_11481);
nor U11866 (N_11866,N_11473,N_11536);
nand U11867 (N_11867,N_11357,N_11401);
nor U11868 (N_11868,N_11539,N_11387);
xor U11869 (N_11869,N_11509,N_11598);
nor U11870 (N_11870,N_11558,N_11240);
and U11871 (N_11871,N_11577,N_11472);
and U11872 (N_11872,N_11579,N_11491);
or U11873 (N_11873,N_11517,N_11430);
and U11874 (N_11874,N_11534,N_11256);
xor U11875 (N_11875,N_11242,N_11414);
xnor U11876 (N_11876,N_11475,N_11326);
xnor U11877 (N_11877,N_11599,N_11389);
nor U11878 (N_11878,N_11493,N_11221);
nand U11879 (N_11879,N_11206,N_11543);
xor U11880 (N_11880,N_11424,N_11224);
xnor U11881 (N_11881,N_11551,N_11258);
and U11882 (N_11882,N_11290,N_11446);
and U11883 (N_11883,N_11270,N_11528);
nand U11884 (N_11884,N_11231,N_11215);
nor U11885 (N_11885,N_11329,N_11561);
xor U11886 (N_11886,N_11552,N_11401);
or U11887 (N_11887,N_11290,N_11339);
and U11888 (N_11888,N_11528,N_11578);
nor U11889 (N_11889,N_11537,N_11353);
xnor U11890 (N_11890,N_11435,N_11216);
or U11891 (N_11891,N_11381,N_11363);
xor U11892 (N_11892,N_11369,N_11422);
xor U11893 (N_11893,N_11455,N_11331);
nand U11894 (N_11894,N_11214,N_11483);
nor U11895 (N_11895,N_11239,N_11294);
and U11896 (N_11896,N_11220,N_11251);
nor U11897 (N_11897,N_11568,N_11492);
or U11898 (N_11898,N_11409,N_11517);
or U11899 (N_11899,N_11441,N_11481);
nor U11900 (N_11900,N_11287,N_11404);
nand U11901 (N_11901,N_11538,N_11239);
nand U11902 (N_11902,N_11285,N_11497);
and U11903 (N_11903,N_11315,N_11254);
nor U11904 (N_11904,N_11392,N_11302);
nand U11905 (N_11905,N_11205,N_11224);
nor U11906 (N_11906,N_11477,N_11561);
nand U11907 (N_11907,N_11210,N_11460);
nor U11908 (N_11908,N_11225,N_11324);
and U11909 (N_11909,N_11296,N_11293);
and U11910 (N_11910,N_11301,N_11254);
and U11911 (N_11911,N_11509,N_11354);
or U11912 (N_11912,N_11540,N_11342);
and U11913 (N_11913,N_11447,N_11419);
nand U11914 (N_11914,N_11392,N_11226);
nor U11915 (N_11915,N_11490,N_11402);
xnor U11916 (N_11916,N_11283,N_11243);
nand U11917 (N_11917,N_11533,N_11245);
and U11918 (N_11918,N_11591,N_11267);
nand U11919 (N_11919,N_11495,N_11337);
or U11920 (N_11920,N_11258,N_11336);
nor U11921 (N_11921,N_11463,N_11295);
and U11922 (N_11922,N_11462,N_11503);
nand U11923 (N_11923,N_11395,N_11295);
nor U11924 (N_11924,N_11409,N_11258);
nand U11925 (N_11925,N_11502,N_11500);
xnor U11926 (N_11926,N_11586,N_11352);
or U11927 (N_11927,N_11519,N_11204);
or U11928 (N_11928,N_11221,N_11598);
or U11929 (N_11929,N_11294,N_11364);
and U11930 (N_11930,N_11354,N_11335);
xor U11931 (N_11931,N_11374,N_11237);
xnor U11932 (N_11932,N_11499,N_11478);
xor U11933 (N_11933,N_11256,N_11214);
nor U11934 (N_11934,N_11348,N_11589);
nor U11935 (N_11935,N_11200,N_11241);
nand U11936 (N_11936,N_11538,N_11245);
xnor U11937 (N_11937,N_11226,N_11296);
nor U11938 (N_11938,N_11513,N_11319);
or U11939 (N_11939,N_11312,N_11569);
or U11940 (N_11940,N_11442,N_11399);
or U11941 (N_11941,N_11451,N_11531);
and U11942 (N_11942,N_11342,N_11310);
or U11943 (N_11943,N_11453,N_11349);
nor U11944 (N_11944,N_11419,N_11261);
nor U11945 (N_11945,N_11247,N_11551);
nand U11946 (N_11946,N_11342,N_11559);
or U11947 (N_11947,N_11553,N_11359);
or U11948 (N_11948,N_11459,N_11585);
nand U11949 (N_11949,N_11572,N_11492);
xnor U11950 (N_11950,N_11586,N_11407);
nand U11951 (N_11951,N_11243,N_11492);
or U11952 (N_11952,N_11215,N_11579);
and U11953 (N_11953,N_11310,N_11374);
and U11954 (N_11954,N_11252,N_11265);
or U11955 (N_11955,N_11248,N_11524);
xor U11956 (N_11956,N_11431,N_11400);
xnor U11957 (N_11957,N_11248,N_11330);
nor U11958 (N_11958,N_11470,N_11383);
or U11959 (N_11959,N_11507,N_11267);
nor U11960 (N_11960,N_11285,N_11505);
nor U11961 (N_11961,N_11444,N_11495);
or U11962 (N_11962,N_11520,N_11356);
nor U11963 (N_11963,N_11546,N_11403);
nand U11964 (N_11964,N_11599,N_11464);
nand U11965 (N_11965,N_11460,N_11484);
and U11966 (N_11966,N_11503,N_11318);
xor U11967 (N_11967,N_11210,N_11292);
xnor U11968 (N_11968,N_11526,N_11358);
nor U11969 (N_11969,N_11509,N_11266);
and U11970 (N_11970,N_11404,N_11369);
nor U11971 (N_11971,N_11301,N_11588);
and U11972 (N_11972,N_11438,N_11249);
nand U11973 (N_11973,N_11206,N_11212);
and U11974 (N_11974,N_11265,N_11522);
nand U11975 (N_11975,N_11308,N_11418);
nor U11976 (N_11976,N_11206,N_11409);
xnor U11977 (N_11977,N_11458,N_11334);
and U11978 (N_11978,N_11546,N_11272);
or U11979 (N_11979,N_11463,N_11577);
and U11980 (N_11980,N_11374,N_11539);
nand U11981 (N_11981,N_11345,N_11219);
xnor U11982 (N_11982,N_11285,N_11516);
nor U11983 (N_11983,N_11542,N_11350);
or U11984 (N_11984,N_11327,N_11297);
and U11985 (N_11985,N_11531,N_11512);
nand U11986 (N_11986,N_11450,N_11506);
nor U11987 (N_11987,N_11549,N_11553);
and U11988 (N_11988,N_11583,N_11261);
nor U11989 (N_11989,N_11432,N_11308);
and U11990 (N_11990,N_11428,N_11460);
nor U11991 (N_11991,N_11400,N_11257);
or U11992 (N_11992,N_11453,N_11442);
or U11993 (N_11993,N_11242,N_11545);
xnor U11994 (N_11994,N_11598,N_11447);
nor U11995 (N_11995,N_11302,N_11344);
xnor U11996 (N_11996,N_11403,N_11208);
and U11997 (N_11997,N_11262,N_11231);
or U11998 (N_11998,N_11293,N_11514);
xnor U11999 (N_11999,N_11565,N_11569);
or U12000 (N_12000,N_11850,N_11724);
nor U12001 (N_12001,N_11754,N_11795);
and U12002 (N_12002,N_11786,N_11934);
nor U12003 (N_12003,N_11875,N_11717);
and U12004 (N_12004,N_11680,N_11682);
or U12005 (N_12005,N_11723,N_11778);
and U12006 (N_12006,N_11700,N_11887);
nor U12007 (N_12007,N_11952,N_11982);
xor U12008 (N_12008,N_11613,N_11731);
nand U12009 (N_12009,N_11602,N_11898);
nand U12010 (N_12010,N_11752,N_11812);
nand U12011 (N_12011,N_11943,N_11806);
nand U12012 (N_12012,N_11766,N_11758);
and U12013 (N_12013,N_11616,N_11954);
and U12014 (N_12014,N_11902,N_11990);
nor U12015 (N_12015,N_11819,N_11994);
xor U12016 (N_12016,N_11715,N_11671);
nand U12017 (N_12017,N_11894,N_11980);
xnor U12018 (N_12018,N_11647,N_11824);
nand U12019 (N_12019,N_11790,N_11788);
and U12020 (N_12020,N_11820,N_11776);
nor U12021 (N_12021,N_11794,N_11876);
xnor U12022 (N_12022,N_11753,N_11730);
nor U12023 (N_12023,N_11770,N_11608);
and U12024 (N_12024,N_11698,N_11912);
and U12025 (N_12025,N_11746,N_11796);
nand U12026 (N_12026,N_11967,N_11621);
and U12027 (N_12027,N_11683,N_11692);
xor U12028 (N_12028,N_11989,N_11813);
nand U12029 (N_12029,N_11638,N_11888);
or U12030 (N_12030,N_11914,N_11609);
nor U12031 (N_12031,N_11726,N_11665);
nor U12032 (N_12032,N_11631,N_11699);
nand U12033 (N_12033,N_11827,N_11991);
xor U12034 (N_12034,N_11856,N_11840);
nand U12035 (N_12035,N_11646,N_11889);
or U12036 (N_12036,N_11949,N_11689);
nand U12037 (N_12037,N_11624,N_11627);
or U12038 (N_12038,N_11670,N_11904);
xor U12039 (N_12039,N_11821,N_11641);
nand U12040 (N_12040,N_11880,N_11755);
and U12041 (N_12041,N_11639,N_11760);
nand U12042 (N_12042,N_11618,N_11725);
xnor U12043 (N_12043,N_11668,N_11635);
or U12044 (N_12044,N_11958,N_11906);
nor U12045 (N_12045,N_11779,N_11977);
nand U12046 (N_12046,N_11964,N_11745);
xor U12047 (N_12047,N_11716,N_11910);
nor U12048 (N_12048,N_11860,N_11858);
or U12049 (N_12049,N_11893,N_11793);
nor U12050 (N_12050,N_11749,N_11721);
nor U12051 (N_12051,N_11686,N_11973);
xor U12052 (N_12052,N_11604,N_11871);
nand U12053 (N_12053,N_11764,N_11787);
nor U12054 (N_12054,N_11763,N_11789);
and U12055 (N_12055,N_11942,N_11679);
xnor U12056 (N_12056,N_11714,N_11999);
nand U12057 (N_12057,N_11853,N_11828);
and U12058 (N_12058,N_11917,N_11862);
xnor U12059 (N_12059,N_11945,N_11899);
xor U12060 (N_12060,N_11685,N_11773);
and U12061 (N_12061,N_11817,N_11831);
xnor U12062 (N_12062,N_11959,N_11815);
nor U12063 (N_12063,N_11722,N_11644);
nor U12064 (N_12064,N_11935,N_11688);
nand U12065 (N_12065,N_11802,N_11907);
nor U12066 (N_12066,N_11791,N_11709);
xor U12067 (N_12067,N_11883,N_11941);
nor U12068 (N_12068,N_11933,N_11744);
nand U12069 (N_12069,N_11829,N_11854);
nand U12070 (N_12070,N_11866,N_11610);
or U12071 (N_12071,N_11948,N_11693);
and U12072 (N_12072,N_11834,N_11861);
xor U12073 (N_12073,N_11878,N_11735);
xor U12074 (N_12074,N_11600,N_11605);
xor U12075 (N_12075,N_11658,N_11841);
and U12076 (N_12076,N_11626,N_11676);
xnor U12077 (N_12077,N_11909,N_11783);
and U12078 (N_12078,N_11785,N_11847);
or U12079 (N_12079,N_11923,N_11897);
or U12080 (N_12080,N_11983,N_11984);
and U12081 (N_12081,N_11988,N_11678);
or U12082 (N_12082,N_11781,N_11937);
xnor U12083 (N_12083,N_11739,N_11975);
xnor U12084 (N_12084,N_11891,N_11661);
nor U12085 (N_12085,N_11657,N_11884);
nor U12086 (N_12086,N_11921,N_11712);
xor U12087 (N_12087,N_11896,N_11986);
nand U12088 (N_12088,N_11979,N_11911);
and U12089 (N_12089,N_11908,N_11625);
nor U12090 (N_12090,N_11656,N_11895);
nor U12091 (N_12091,N_11792,N_11701);
nor U12092 (N_12092,N_11675,N_11614);
or U12093 (N_12093,N_11966,N_11633);
nand U12094 (N_12094,N_11762,N_11777);
and U12095 (N_12095,N_11747,N_11929);
nor U12096 (N_12096,N_11940,N_11603);
or U12097 (N_12097,N_11711,N_11851);
and U12098 (N_12098,N_11843,N_11863);
nand U12099 (N_12099,N_11873,N_11920);
and U12100 (N_12100,N_11913,N_11767);
xnor U12101 (N_12101,N_11833,N_11844);
or U12102 (N_12102,N_11947,N_11901);
and U12103 (N_12103,N_11642,N_11607);
or U12104 (N_12104,N_11771,N_11710);
xnor U12105 (N_12105,N_11927,N_11832);
nor U12106 (N_12106,N_11669,N_11737);
nand U12107 (N_12107,N_11892,N_11836);
xor U12108 (N_12108,N_11719,N_11772);
or U12109 (N_12109,N_11932,N_11830);
nor U12110 (N_12110,N_11885,N_11846);
nand U12111 (N_12111,N_11981,N_11759);
nor U12112 (N_12112,N_11780,N_11992);
or U12113 (N_12113,N_11708,N_11867);
and U12114 (N_12114,N_11713,N_11944);
or U12115 (N_12115,N_11743,N_11696);
nor U12116 (N_12116,N_11769,N_11838);
xor U12117 (N_12117,N_11740,N_11842);
and U12118 (N_12118,N_11852,N_11922);
or U12119 (N_12119,N_11868,N_11687);
nand U12120 (N_12120,N_11742,N_11651);
or U12121 (N_12121,N_11877,N_11957);
and U12122 (N_12122,N_11918,N_11667);
xnor U12123 (N_12123,N_11629,N_11648);
xnor U12124 (N_12124,N_11799,N_11775);
xnor U12125 (N_12125,N_11652,N_11619);
nand U12126 (N_12126,N_11951,N_11872);
or U12127 (N_12127,N_11707,N_11808);
and U12128 (N_12128,N_11645,N_11919);
nor U12129 (N_12129,N_11765,N_11653);
xnor U12130 (N_12130,N_11774,N_11650);
nand U12131 (N_12131,N_11695,N_11797);
nand U12132 (N_12132,N_11968,N_11729);
nor U12133 (N_12133,N_11677,N_11601);
nand U12134 (N_12134,N_11800,N_11950);
xor U12135 (N_12135,N_11874,N_11637);
nor U12136 (N_12136,N_11620,N_11643);
and U12137 (N_12137,N_11750,N_11663);
nand U12138 (N_12138,N_11628,N_11636);
nor U12139 (N_12139,N_11998,N_11963);
or U12140 (N_12140,N_11926,N_11818);
and U12141 (N_12141,N_11936,N_11703);
or U12142 (N_12142,N_11816,N_11946);
nand U12143 (N_12143,N_11810,N_11811);
xor U12144 (N_12144,N_11809,N_11659);
nor U12145 (N_12145,N_11974,N_11886);
nor U12146 (N_12146,N_11865,N_11741);
or U12147 (N_12147,N_11751,N_11634);
and U12148 (N_12148,N_11969,N_11997);
nor U12149 (N_12149,N_11807,N_11674);
or U12150 (N_12150,N_11837,N_11903);
or U12151 (N_12151,N_11953,N_11697);
nor U12152 (N_12152,N_11732,N_11915);
or U12153 (N_12153,N_11761,N_11839);
nor U12154 (N_12154,N_11718,N_11870);
or U12155 (N_12155,N_11823,N_11814);
nor U12156 (N_12156,N_11690,N_11938);
xor U12157 (N_12157,N_11782,N_11655);
or U12158 (N_12158,N_11632,N_11673);
and U12159 (N_12159,N_11640,N_11855);
or U12160 (N_12160,N_11976,N_11857);
nor U12161 (N_12161,N_11623,N_11704);
xnor U12162 (N_12162,N_11955,N_11924);
nand U12163 (N_12163,N_11826,N_11881);
nor U12164 (N_12164,N_11672,N_11930);
nor U12165 (N_12165,N_11734,N_11939);
and U12166 (N_12166,N_11803,N_11664);
or U12167 (N_12167,N_11702,N_11606);
nor U12168 (N_12168,N_11728,N_11845);
or U12169 (N_12169,N_11705,N_11798);
xnor U12170 (N_12170,N_11617,N_11733);
nor U12171 (N_12171,N_11622,N_11993);
xor U12172 (N_12172,N_11978,N_11848);
nor U12173 (N_12173,N_11971,N_11987);
nand U12174 (N_12174,N_11649,N_11801);
nor U12175 (N_12175,N_11849,N_11931);
nor U12176 (N_12176,N_11864,N_11666);
and U12177 (N_12177,N_11961,N_11905);
or U12178 (N_12178,N_11900,N_11748);
xnor U12179 (N_12179,N_11706,N_11615);
xor U12180 (N_12180,N_11660,N_11962);
or U12181 (N_12181,N_11995,N_11694);
and U12182 (N_12182,N_11879,N_11681);
or U12183 (N_12183,N_11960,N_11859);
nor U12184 (N_12184,N_11965,N_11928);
nor U12185 (N_12185,N_11611,N_11835);
or U12186 (N_12186,N_11925,N_11720);
xnor U12187 (N_12187,N_11869,N_11662);
nand U12188 (N_12188,N_11916,N_11985);
nor U12189 (N_12189,N_11727,N_11972);
xor U12190 (N_12190,N_11882,N_11691);
nor U12191 (N_12191,N_11822,N_11805);
nor U12192 (N_12192,N_11756,N_11654);
and U12193 (N_12193,N_11684,N_11757);
and U12194 (N_12194,N_11612,N_11890);
or U12195 (N_12195,N_11996,N_11630);
nor U12196 (N_12196,N_11804,N_11970);
and U12197 (N_12197,N_11825,N_11784);
nor U12198 (N_12198,N_11736,N_11956);
and U12199 (N_12199,N_11738,N_11768);
and U12200 (N_12200,N_11684,N_11904);
nand U12201 (N_12201,N_11797,N_11811);
nor U12202 (N_12202,N_11643,N_11826);
and U12203 (N_12203,N_11675,N_11747);
nand U12204 (N_12204,N_11681,N_11799);
and U12205 (N_12205,N_11722,N_11991);
or U12206 (N_12206,N_11906,N_11921);
or U12207 (N_12207,N_11642,N_11653);
or U12208 (N_12208,N_11917,N_11975);
and U12209 (N_12209,N_11800,N_11663);
nor U12210 (N_12210,N_11754,N_11895);
nor U12211 (N_12211,N_11698,N_11997);
xnor U12212 (N_12212,N_11859,N_11903);
xnor U12213 (N_12213,N_11861,N_11758);
nor U12214 (N_12214,N_11967,N_11898);
nor U12215 (N_12215,N_11719,N_11786);
or U12216 (N_12216,N_11832,N_11825);
or U12217 (N_12217,N_11736,N_11685);
xnor U12218 (N_12218,N_11617,N_11905);
and U12219 (N_12219,N_11961,N_11783);
xor U12220 (N_12220,N_11698,N_11999);
nor U12221 (N_12221,N_11913,N_11854);
and U12222 (N_12222,N_11840,N_11630);
xor U12223 (N_12223,N_11765,N_11929);
xor U12224 (N_12224,N_11667,N_11675);
or U12225 (N_12225,N_11801,N_11776);
nor U12226 (N_12226,N_11823,N_11972);
xor U12227 (N_12227,N_11655,N_11753);
and U12228 (N_12228,N_11953,N_11956);
and U12229 (N_12229,N_11958,N_11618);
nor U12230 (N_12230,N_11654,N_11851);
or U12231 (N_12231,N_11916,N_11810);
nand U12232 (N_12232,N_11713,N_11776);
nor U12233 (N_12233,N_11633,N_11659);
and U12234 (N_12234,N_11888,N_11883);
and U12235 (N_12235,N_11988,N_11685);
nor U12236 (N_12236,N_11785,N_11620);
nand U12237 (N_12237,N_11818,N_11900);
and U12238 (N_12238,N_11739,N_11772);
or U12239 (N_12239,N_11657,N_11961);
nand U12240 (N_12240,N_11879,N_11603);
nor U12241 (N_12241,N_11964,N_11777);
xnor U12242 (N_12242,N_11601,N_11742);
nor U12243 (N_12243,N_11664,N_11951);
nand U12244 (N_12244,N_11871,N_11744);
xnor U12245 (N_12245,N_11920,N_11862);
xnor U12246 (N_12246,N_11930,N_11760);
xor U12247 (N_12247,N_11622,N_11627);
and U12248 (N_12248,N_11716,N_11851);
nor U12249 (N_12249,N_11973,N_11788);
nor U12250 (N_12250,N_11851,N_11690);
and U12251 (N_12251,N_11907,N_11657);
xor U12252 (N_12252,N_11878,N_11830);
xnor U12253 (N_12253,N_11980,N_11906);
xor U12254 (N_12254,N_11636,N_11917);
or U12255 (N_12255,N_11632,N_11843);
xor U12256 (N_12256,N_11701,N_11717);
xor U12257 (N_12257,N_11862,N_11679);
xor U12258 (N_12258,N_11664,N_11781);
nand U12259 (N_12259,N_11814,N_11940);
nand U12260 (N_12260,N_11606,N_11958);
and U12261 (N_12261,N_11751,N_11631);
and U12262 (N_12262,N_11730,N_11980);
nand U12263 (N_12263,N_11731,N_11810);
nor U12264 (N_12264,N_11900,N_11689);
nand U12265 (N_12265,N_11819,N_11942);
nor U12266 (N_12266,N_11636,N_11785);
nand U12267 (N_12267,N_11926,N_11696);
nand U12268 (N_12268,N_11790,N_11735);
xor U12269 (N_12269,N_11800,N_11868);
nor U12270 (N_12270,N_11993,N_11929);
xor U12271 (N_12271,N_11701,N_11889);
nor U12272 (N_12272,N_11606,N_11956);
xnor U12273 (N_12273,N_11864,N_11894);
nand U12274 (N_12274,N_11772,N_11609);
nor U12275 (N_12275,N_11768,N_11721);
and U12276 (N_12276,N_11992,N_11850);
nor U12277 (N_12277,N_11962,N_11782);
or U12278 (N_12278,N_11661,N_11755);
nand U12279 (N_12279,N_11668,N_11967);
nor U12280 (N_12280,N_11983,N_11772);
or U12281 (N_12281,N_11652,N_11807);
nor U12282 (N_12282,N_11957,N_11831);
xnor U12283 (N_12283,N_11823,N_11902);
nor U12284 (N_12284,N_11832,N_11848);
nor U12285 (N_12285,N_11702,N_11670);
and U12286 (N_12286,N_11661,N_11939);
nor U12287 (N_12287,N_11896,N_11958);
nor U12288 (N_12288,N_11794,N_11743);
nor U12289 (N_12289,N_11934,N_11849);
nor U12290 (N_12290,N_11787,N_11886);
nor U12291 (N_12291,N_11868,N_11905);
or U12292 (N_12292,N_11895,N_11783);
nor U12293 (N_12293,N_11629,N_11635);
and U12294 (N_12294,N_11854,N_11936);
or U12295 (N_12295,N_11761,N_11873);
xor U12296 (N_12296,N_11945,N_11908);
or U12297 (N_12297,N_11677,N_11742);
and U12298 (N_12298,N_11729,N_11689);
xnor U12299 (N_12299,N_11689,N_11992);
nand U12300 (N_12300,N_11947,N_11676);
or U12301 (N_12301,N_11604,N_11970);
nand U12302 (N_12302,N_11898,N_11880);
or U12303 (N_12303,N_11611,N_11608);
xor U12304 (N_12304,N_11949,N_11825);
nor U12305 (N_12305,N_11944,N_11707);
nor U12306 (N_12306,N_11631,N_11887);
nor U12307 (N_12307,N_11767,N_11642);
nand U12308 (N_12308,N_11995,N_11863);
and U12309 (N_12309,N_11921,N_11803);
nand U12310 (N_12310,N_11863,N_11918);
and U12311 (N_12311,N_11819,N_11878);
nor U12312 (N_12312,N_11723,N_11748);
nor U12313 (N_12313,N_11672,N_11635);
or U12314 (N_12314,N_11846,N_11988);
or U12315 (N_12315,N_11756,N_11678);
xor U12316 (N_12316,N_11787,N_11797);
nor U12317 (N_12317,N_11935,N_11784);
xnor U12318 (N_12318,N_11928,N_11899);
or U12319 (N_12319,N_11646,N_11743);
nand U12320 (N_12320,N_11783,N_11715);
xnor U12321 (N_12321,N_11742,N_11824);
and U12322 (N_12322,N_11618,N_11716);
and U12323 (N_12323,N_11797,N_11934);
xnor U12324 (N_12324,N_11730,N_11786);
nor U12325 (N_12325,N_11825,N_11641);
or U12326 (N_12326,N_11729,N_11809);
xnor U12327 (N_12327,N_11622,N_11965);
or U12328 (N_12328,N_11655,N_11895);
nor U12329 (N_12329,N_11687,N_11807);
and U12330 (N_12330,N_11776,N_11646);
xnor U12331 (N_12331,N_11891,N_11901);
xnor U12332 (N_12332,N_11795,N_11964);
xor U12333 (N_12333,N_11745,N_11629);
xnor U12334 (N_12334,N_11857,N_11916);
xor U12335 (N_12335,N_11614,N_11653);
xor U12336 (N_12336,N_11951,N_11785);
nor U12337 (N_12337,N_11933,N_11669);
and U12338 (N_12338,N_11690,N_11625);
nand U12339 (N_12339,N_11875,N_11751);
nor U12340 (N_12340,N_11790,N_11845);
and U12341 (N_12341,N_11719,N_11935);
or U12342 (N_12342,N_11604,N_11961);
or U12343 (N_12343,N_11989,N_11836);
xnor U12344 (N_12344,N_11751,N_11749);
nand U12345 (N_12345,N_11983,N_11987);
and U12346 (N_12346,N_11672,N_11923);
xor U12347 (N_12347,N_11875,N_11946);
and U12348 (N_12348,N_11958,N_11672);
or U12349 (N_12349,N_11873,N_11896);
nor U12350 (N_12350,N_11801,N_11673);
nand U12351 (N_12351,N_11720,N_11909);
xor U12352 (N_12352,N_11722,N_11634);
nor U12353 (N_12353,N_11701,N_11939);
and U12354 (N_12354,N_11811,N_11892);
nand U12355 (N_12355,N_11863,N_11884);
and U12356 (N_12356,N_11918,N_11689);
or U12357 (N_12357,N_11787,N_11963);
or U12358 (N_12358,N_11993,N_11891);
nor U12359 (N_12359,N_11696,N_11765);
xnor U12360 (N_12360,N_11881,N_11959);
nand U12361 (N_12361,N_11809,N_11798);
nor U12362 (N_12362,N_11886,N_11881);
nand U12363 (N_12363,N_11887,N_11677);
xnor U12364 (N_12364,N_11783,N_11813);
or U12365 (N_12365,N_11714,N_11954);
and U12366 (N_12366,N_11693,N_11898);
nor U12367 (N_12367,N_11702,N_11793);
and U12368 (N_12368,N_11793,N_11898);
or U12369 (N_12369,N_11805,N_11656);
xnor U12370 (N_12370,N_11883,N_11906);
or U12371 (N_12371,N_11911,N_11787);
and U12372 (N_12372,N_11835,N_11633);
and U12373 (N_12373,N_11601,N_11744);
or U12374 (N_12374,N_11875,N_11919);
or U12375 (N_12375,N_11617,N_11971);
xor U12376 (N_12376,N_11700,N_11757);
or U12377 (N_12377,N_11787,N_11808);
and U12378 (N_12378,N_11630,N_11649);
nor U12379 (N_12379,N_11754,N_11794);
and U12380 (N_12380,N_11681,N_11892);
nor U12381 (N_12381,N_11680,N_11944);
or U12382 (N_12382,N_11628,N_11614);
and U12383 (N_12383,N_11642,N_11695);
xnor U12384 (N_12384,N_11798,N_11773);
or U12385 (N_12385,N_11884,N_11868);
and U12386 (N_12386,N_11837,N_11641);
xor U12387 (N_12387,N_11655,N_11775);
nor U12388 (N_12388,N_11647,N_11839);
nand U12389 (N_12389,N_11946,N_11672);
xor U12390 (N_12390,N_11642,N_11661);
nor U12391 (N_12391,N_11969,N_11830);
and U12392 (N_12392,N_11801,N_11717);
and U12393 (N_12393,N_11936,N_11875);
nor U12394 (N_12394,N_11976,N_11790);
and U12395 (N_12395,N_11675,N_11732);
and U12396 (N_12396,N_11768,N_11613);
nor U12397 (N_12397,N_11689,N_11697);
nand U12398 (N_12398,N_11723,N_11638);
or U12399 (N_12399,N_11772,N_11826);
or U12400 (N_12400,N_12297,N_12215);
or U12401 (N_12401,N_12340,N_12094);
nand U12402 (N_12402,N_12351,N_12132);
nor U12403 (N_12403,N_12211,N_12219);
or U12404 (N_12404,N_12346,N_12320);
nand U12405 (N_12405,N_12333,N_12205);
nor U12406 (N_12406,N_12078,N_12111);
xor U12407 (N_12407,N_12118,N_12249);
nand U12408 (N_12408,N_12122,N_12031);
nor U12409 (N_12409,N_12197,N_12265);
nor U12410 (N_12410,N_12278,N_12238);
and U12411 (N_12411,N_12166,N_12364);
nor U12412 (N_12412,N_12355,N_12201);
and U12413 (N_12413,N_12144,N_12315);
nor U12414 (N_12414,N_12001,N_12058);
nand U12415 (N_12415,N_12353,N_12038);
xnor U12416 (N_12416,N_12223,N_12218);
nand U12417 (N_12417,N_12212,N_12011);
or U12418 (N_12418,N_12076,N_12334);
xor U12419 (N_12419,N_12075,N_12077);
nor U12420 (N_12420,N_12039,N_12323);
or U12421 (N_12421,N_12348,N_12108);
xnor U12422 (N_12422,N_12307,N_12309);
or U12423 (N_12423,N_12386,N_12004);
nor U12424 (N_12424,N_12327,N_12109);
or U12425 (N_12425,N_12347,N_12274);
nand U12426 (N_12426,N_12081,N_12266);
nor U12427 (N_12427,N_12016,N_12252);
xor U12428 (N_12428,N_12222,N_12377);
and U12429 (N_12429,N_12200,N_12380);
nand U12430 (N_12430,N_12032,N_12234);
xnor U12431 (N_12431,N_12220,N_12376);
nand U12432 (N_12432,N_12088,N_12126);
nand U12433 (N_12433,N_12229,N_12100);
xor U12434 (N_12434,N_12378,N_12103);
and U12435 (N_12435,N_12285,N_12368);
nor U12436 (N_12436,N_12165,N_12383);
nand U12437 (N_12437,N_12370,N_12231);
and U12438 (N_12438,N_12124,N_12034);
nand U12439 (N_12439,N_12180,N_12008);
or U12440 (N_12440,N_12208,N_12299);
or U12441 (N_12441,N_12157,N_12134);
nand U12442 (N_12442,N_12254,N_12375);
or U12443 (N_12443,N_12324,N_12046);
or U12444 (N_12444,N_12236,N_12350);
xnor U12445 (N_12445,N_12233,N_12015);
and U12446 (N_12446,N_12174,N_12171);
xnor U12447 (N_12447,N_12105,N_12248);
xnor U12448 (N_12448,N_12083,N_12151);
xnor U12449 (N_12449,N_12337,N_12176);
or U12450 (N_12450,N_12025,N_12204);
nand U12451 (N_12451,N_12009,N_12255);
nand U12452 (N_12452,N_12059,N_12012);
and U12453 (N_12453,N_12360,N_12147);
or U12454 (N_12454,N_12245,N_12028);
nor U12455 (N_12455,N_12087,N_12116);
or U12456 (N_12456,N_12128,N_12125);
nand U12457 (N_12457,N_12371,N_12095);
or U12458 (N_12458,N_12247,N_12318);
nand U12459 (N_12459,N_12206,N_12057);
xor U12460 (N_12460,N_12013,N_12336);
or U12461 (N_12461,N_12101,N_12106);
nand U12462 (N_12462,N_12258,N_12048);
nand U12463 (N_12463,N_12143,N_12372);
nor U12464 (N_12464,N_12352,N_12262);
or U12465 (N_12465,N_12163,N_12399);
and U12466 (N_12466,N_12369,N_12096);
or U12467 (N_12467,N_12127,N_12068);
xnor U12468 (N_12468,N_12186,N_12043);
xnor U12469 (N_12469,N_12185,N_12005);
xnor U12470 (N_12470,N_12183,N_12207);
and U12471 (N_12471,N_12289,N_12036);
xnor U12472 (N_12472,N_12045,N_12021);
or U12473 (N_12473,N_12269,N_12029);
nand U12474 (N_12474,N_12339,N_12209);
nand U12475 (N_12475,N_12317,N_12395);
xor U12476 (N_12476,N_12062,N_12253);
and U12477 (N_12477,N_12026,N_12193);
xnor U12478 (N_12478,N_12225,N_12121);
nand U12479 (N_12479,N_12194,N_12330);
xor U12480 (N_12480,N_12308,N_12052);
nand U12481 (N_12481,N_12051,N_12343);
nor U12482 (N_12482,N_12304,N_12305);
or U12483 (N_12483,N_12182,N_12136);
nor U12484 (N_12484,N_12164,N_12130);
and U12485 (N_12485,N_12049,N_12177);
xor U12486 (N_12486,N_12161,N_12356);
nor U12487 (N_12487,N_12006,N_12374);
and U12488 (N_12488,N_12316,N_12153);
xor U12489 (N_12489,N_12089,N_12159);
nor U12490 (N_12490,N_12060,N_12002);
nor U12491 (N_12491,N_12091,N_12071);
and U12492 (N_12492,N_12251,N_12181);
xor U12493 (N_12493,N_12342,N_12148);
nand U12494 (N_12494,N_12150,N_12063);
and U12495 (N_12495,N_12198,N_12079);
and U12496 (N_12496,N_12240,N_12366);
or U12497 (N_12497,N_12267,N_12263);
nand U12498 (N_12498,N_12155,N_12199);
nor U12499 (N_12499,N_12170,N_12385);
xor U12500 (N_12500,N_12064,N_12196);
nor U12501 (N_12501,N_12397,N_12053);
nand U12502 (N_12502,N_12033,N_12168);
nand U12503 (N_12503,N_12080,N_12129);
or U12504 (N_12504,N_12050,N_12288);
or U12505 (N_12505,N_12373,N_12329);
xnor U12506 (N_12506,N_12141,N_12092);
or U12507 (N_12507,N_12287,N_12393);
nand U12508 (N_12508,N_12362,N_12396);
nor U12509 (N_12509,N_12345,N_12056);
or U12510 (N_12510,N_12135,N_12314);
xnor U12511 (N_12511,N_12110,N_12149);
nor U12512 (N_12512,N_12246,N_12169);
and U12513 (N_12513,N_12392,N_12226);
xor U12514 (N_12514,N_12260,N_12067);
and U12515 (N_12515,N_12044,N_12082);
or U12516 (N_12516,N_12104,N_12300);
or U12517 (N_12517,N_12384,N_12298);
nand U12518 (N_12518,N_12295,N_12379);
xnor U12519 (N_12519,N_12030,N_12283);
nand U12520 (N_12520,N_12107,N_12224);
or U12521 (N_12521,N_12213,N_12018);
nand U12522 (N_12522,N_12023,N_12230);
or U12523 (N_12523,N_12243,N_12172);
nor U12524 (N_12524,N_12332,N_12156);
or U12525 (N_12525,N_12037,N_12321);
xor U12526 (N_12526,N_12162,N_12202);
nor U12527 (N_12527,N_12261,N_12047);
nor U12528 (N_12528,N_12041,N_12024);
or U12529 (N_12529,N_12235,N_12311);
xnor U12530 (N_12530,N_12173,N_12301);
xnor U12531 (N_12531,N_12146,N_12228);
xnor U12532 (N_12532,N_12072,N_12007);
nand U12533 (N_12533,N_12123,N_12066);
or U12534 (N_12534,N_12354,N_12296);
xnor U12535 (N_12535,N_12195,N_12270);
and U12536 (N_12536,N_12137,N_12341);
nor U12537 (N_12537,N_12085,N_12000);
and U12538 (N_12538,N_12112,N_12221);
and U12539 (N_12539,N_12139,N_12099);
xnor U12540 (N_12540,N_12187,N_12133);
xor U12541 (N_12541,N_12294,N_12256);
nand U12542 (N_12542,N_12264,N_12325);
nor U12543 (N_12543,N_12097,N_12398);
nor U12544 (N_12544,N_12335,N_12084);
or U12545 (N_12545,N_12098,N_12313);
nand U12546 (N_12546,N_12070,N_12019);
and U12547 (N_12547,N_12331,N_12138);
or U12548 (N_12548,N_12268,N_12189);
xnor U12549 (N_12549,N_12061,N_12250);
nand U12550 (N_12550,N_12237,N_12387);
xor U12551 (N_12551,N_12291,N_12145);
nand U12552 (N_12552,N_12178,N_12086);
nand U12553 (N_12553,N_12271,N_12282);
xnor U12554 (N_12554,N_12382,N_12120);
or U12555 (N_12555,N_12119,N_12010);
nand U12556 (N_12556,N_12027,N_12303);
and U12557 (N_12557,N_12179,N_12167);
and U12558 (N_12558,N_12276,N_12306);
xor U12559 (N_12559,N_12114,N_12326);
nand U12560 (N_12560,N_12093,N_12394);
or U12561 (N_12561,N_12003,N_12055);
or U12562 (N_12562,N_12319,N_12239);
nor U12563 (N_12563,N_12281,N_12090);
xor U12564 (N_12564,N_12054,N_12328);
and U12565 (N_12565,N_12279,N_12277);
and U12566 (N_12566,N_12359,N_12131);
nor U12567 (N_12567,N_12020,N_12257);
and U12568 (N_12568,N_12293,N_12184);
xnor U12569 (N_12569,N_12217,N_12290);
nand U12570 (N_12570,N_12160,N_12188);
nor U12571 (N_12571,N_12175,N_12286);
nand U12572 (N_12572,N_12065,N_12273);
xnor U12573 (N_12573,N_12272,N_12192);
and U12574 (N_12574,N_12338,N_12312);
xnor U12575 (N_12575,N_12391,N_12073);
and U12576 (N_12576,N_12280,N_12115);
nand U12577 (N_12577,N_12284,N_12113);
xnor U12578 (N_12578,N_12361,N_12381);
and U12579 (N_12579,N_12154,N_12022);
nor U12580 (N_12580,N_12242,N_12322);
nor U12581 (N_12581,N_12140,N_12358);
or U12582 (N_12582,N_12214,N_12365);
and U12583 (N_12583,N_12158,N_12142);
nor U12584 (N_12584,N_12203,N_12244);
or U12585 (N_12585,N_12102,N_12040);
nand U12586 (N_12586,N_12069,N_12259);
and U12587 (N_12587,N_12302,N_12388);
xnor U12588 (N_12588,N_12117,N_12191);
xor U12589 (N_12589,N_12017,N_12363);
nor U12590 (N_12590,N_12389,N_12241);
nand U12591 (N_12591,N_12275,N_12310);
xnor U12592 (N_12592,N_12390,N_12042);
xnor U12593 (N_12593,N_12190,N_12035);
or U12594 (N_12594,N_12074,N_12216);
nor U12595 (N_12595,N_12349,N_12344);
or U12596 (N_12596,N_12210,N_12232);
nand U12597 (N_12597,N_12357,N_12014);
and U12598 (N_12598,N_12367,N_12152);
nand U12599 (N_12599,N_12292,N_12227);
nor U12600 (N_12600,N_12279,N_12299);
nand U12601 (N_12601,N_12360,N_12189);
or U12602 (N_12602,N_12102,N_12264);
xnor U12603 (N_12603,N_12381,N_12176);
nand U12604 (N_12604,N_12286,N_12274);
xnor U12605 (N_12605,N_12281,N_12339);
nor U12606 (N_12606,N_12196,N_12387);
nor U12607 (N_12607,N_12204,N_12030);
and U12608 (N_12608,N_12277,N_12065);
and U12609 (N_12609,N_12300,N_12031);
or U12610 (N_12610,N_12014,N_12131);
or U12611 (N_12611,N_12077,N_12355);
nor U12612 (N_12612,N_12005,N_12310);
nand U12613 (N_12613,N_12393,N_12066);
nor U12614 (N_12614,N_12011,N_12358);
and U12615 (N_12615,N_12254,N_12064);
nor U12616 (N_12616,N_12048,N_12205);
xor U12617 (N_12617,N_12395,N_12375);
or U12618 (N_12618,N_12123,N_12230);
or U12619 (N_12619,N_12332,N_12043);
nor U12620 (N_12620,N_12207,N_12178);
xor U12621 (N_12621,N_12006,N_12382);
and U12622 (N_12622,N_12229,N_12155);
or U12623 (N_12623,N_12296,N_12073);
xor U12624 (N_12624,N_12040,N_12265);
or U12625 (N_12625,N_12339,N_12116);
xnor U12626 (N_12626,N_12084,N_12113);
or U12627 (N_12627,N_12178,N_12169);
and U12628 (N_12628,N_12121,N_12224);
or U12629 (N_12629,N_12120,N_12218);
nor U12630 (N_12630,N_12241,N_12233);
nand U12631 (N_12631,N_12200,N_12015);
xnor U12632 (N_12632,N_12071,N_12081);
nand U12633 (N_12633,N_12347,N_12393);
nand U12634 (N_12634,N_12382,N_12067);
xnor U12635 (N_12635,N_12041,N_12330);
and U12636 (N_12636,N_12304,N_12361);
nor U12637 (N_12637,N_12376,N_12049);
nand U12638 (N_12638,N_12266,N_12330);
nor U12639 (N_12639,N_12268,N_12126);
nand U12640 (N_12640,N_12232,N_12208);
or U12641 (N_12641,N_12047,N_12140);
xnor U12642 (N_12642,N_12398,N_12190);
nand U12643 (N_12643,N_12179,N_12124);
nand U12644 (N_12644,N_12161,N_12206);
nor U12645 (N_12645,N_12162,N_12009);
and U12646 (N_12646,N_12392,N_12287);
nand U12647 (N_12647,N_12032,N_12111);
and U12648 (N_12648,N_12030,N_12274);
or U12649 (N_12649,N_12251,N_12303);
and U12650 (N_12650,N_12382,N_12361);
nor U12651 (N_12651,N_12036,N_12171);
nor U12652 (N_12652,N_12156,N_12365);
and U12653 (N_12653,N_12007,N_12015);
and U12654 (N_12654,N_12128,N_12384);
xnor U12655 (N_12655,N_12160,N_12154);
or U12656 (N_12656,N_12265,N_12276);
nand U12657 (N_12657,N_12165,N_12348);
nor U12658 (N_12658,N_12382,N_12004);
xor U12659 (N_12659,N_12038,N_12363);
nand U12660 (N_12660,N_12338,N_12198);
xnor U12661 (N_12661,N_12226,N_12317);
nand U12662 (N_12662,N_12330,N_12360);
and U12663 (N_12663,N_12059,N_12247);
nand U12664 (N_12664,N_12188,N_12029);
and U12665 (N_12665,N_12319,N_12043);
xnor U12666 (N_12666,N_12351,N_12228);
nand U12667 (N_12667,N_12229,N_12058);
xor U12668 (N_12668,N_12323,N_12082);
xnor U12669 (N_12669,N_12021,N_12067);
or U12670 (N_12670,N_12318,N_12031);
or U12671 (N_12671,N_12123,N_12383);
nor U12672 (N_12672,N_12337,N_12061);
and U12673 (N_12673,N_12270,N_12289);
nand U12674 (N_12674,N_12189,N_12198);
nand U12675 (N_12675,N_12253,N_12012);
xor U12676 (N_12676,N_12343,N_12095);
nand U12677 (N_12677,N_12150,N_12049);
or U12678 (N_12678,N_12352,N_12062);
or U12679 (N_12679,N_12325,N_12136);
nand U12680 (N_12680,N_12341,N_12129);
nor U12681 (N_12681,N_12296,N_12134);
nand U12682 (N_12682,N_12107,N_12040);
or U12683 (N_12683,N_12230,N_12100);
nor U12684 (N_12684,N_12173,N_12207);
or U12685 (N_12685,N_12032,N_12108);
or U12686 (N_12686,N_12285,N_12091);
xnor U12687 (N_12687,N_12130,N_12232);
nor U12688 (N_12688,N_12356,N_12293);
nor U12689 (N_12689,N_12103,N_12213);
nor U12690 (N_12690,N_12326,N_12309);
nand U12691 (N_12691,N_12193,N_12136);
nor U12692 (N_12692,N_12135,N_12259);
xor U12693 (N_12693,N_12107,N_12172);
or U12694 (N_12694,N_12286,N_12184);
xor U12695 (N_12695,N_12212,N_12251);
or U12696 (N_12696,N_12074,N_12293);
nand U12697 (N_12697,N_12268,N_12178);
nand U12698 (N_12698,N_12341,N_12313);
nand U12699 (N_12699,N_12137,N_12315);
or U12700 (N_12700,N_12086,N_12379);
nor U12701 (N_12701,N_12117,N_12009);
nand U12702 (N_12702,N_12366,N_12345);
or U12703 (N_12703,N_12183,N_12190);
and U12704 (N_12704,N_12129,N_12335);
nor U12705 (N_12705,N_12104,N_12315);
nor U12706 (N_12706,N_12211,N_12124);
and U12707 (N_12707,N_12237,N_12314);
nand U12708 (N_12708,N_12261,N_12247);
nand U12709 (N_12709,N_12370,N_12189);
nor U12710 (N_12710,N_12286,N_12331);
nor U12711 (N_12711,N_12158,N_12123);
xor U12712 (N_12712,N_12012,N_12366);
nor U12713 (N_12713,N_12099,N_12284);
or U12714 (N_12714,N_12272,N_12119);
and U12715 (N_12715,N_12312,N_12390);
nand U12716 (N_12716,N_12192,N_12151);
or U12717 (N_12717,N_12003,N_12196);
xnor U12718 (N_12718,N_12086,N_12126);
nor U12719 (N_12719,N_12396,N_12269);
nand U12720 (N_12720,N_12107,N_12328);
xor U12721 (N_12721,N_12236,N_12130);
nor U12722 (N_12722,N_12378,N_12052);
and U12723 (N_12723,N_12031,N_12022);
nor U12724 (N_12724,N_12089,N_12132);
xnor U12725 (N_12725,N_12266,N_12006);
xor U12726 (N_12726,N_12070,N_12274);
xor U12727 (N_12727,N_12030,N_12314);
and U12728 (N_12728,N_12364,N_12141);
nand U12729 (N_12729,N_12311,N_12221);
nand U12730 (N_12730,N_12313,N_12008);
xor U12731 (N_12731,N_12160,N_12039);
or U12732 (N_12732,N_12382,N_12069);
or U12733 (N_12733,N_12237,N_12246);
nand U12734 (N_12734,N_12060,N_12254);
or U12735 (N_12735,N_12013,N_12231);
or U12736 (N_12736,N_12307,N_12177);
or U12737 (N_12737,N_12112,N_12262);
or U12738 (N_12738,N_12239,N_12056);
nand U12739 (N_12739,N_12394,N_12290);
xnor U12740 (N_12740,N_12121,N_12105);
or U12741 (N_12741,N_12206,N_12393);
xor U12742 (N_12742,N_12354,N_12179);
and U12743 (N_12743,N_12200,N_12078);
and U12744 (N_12744,N_12130,N_12169);
and U12745 (N_12745,N_12186,N_12281);
nand U12746 (N_12746,N_12098,N_12118);
nand U12747 (N_12747,N_12110,N_12022);
and U12748 (N_12748,N_12254,N_12389);
or U12749 (N_12749,N_12329,N_12138);
nor U12750 (N_12750,N_12161,N_12307);
and U12751 (N_12751,N_12331,N_12018);
nor U12752 (N_12752,N_12162,N_12350);
xnor U12753 (N_12753,N_12268,N_12351);
or U12754 (N_12754,N_12028,N_12107);
nor U12755 (N_12755,N_12071,N_12148);
or U12756 (N_12756,N_12149,N_12389);
nor U12757 (N_12757,N_12353,N_12143);
nor U12758 (N_12758,N_12046,N_12107);
or U12759 (N_12759,N_12108,N_12119);
xnor U12760 (N_12760,N_12286,N_12091);
and U12761 (N_12761,N_12375,N_12080);
and U12762 (N_12762,N_12292,N_12147);
nor U12763 (N_12763,N_12053,N_12066);
and U12764 (N_12764,N_12142,N_12225);
or U12765 (N_12765,N_12376,N_12321);
and U12766 (N_12766,N_12121,N_12285);
xor U12767 (N_12767,N_12134,N_12387);
and U12768 (N_12768,N_12194,N_12357);
xor U12769 (N_12769,N_12144,N_12375);
nand U12770 (N_12770,N_12019,N_12270);
nand U12771 (N_12771,N_12028,N_12141);
or U12772 (N_12772,N_12114,N_12061);
or U12773 (N_12773,N_12395,N_12075);
and U12774 (N_12774,N_12213,N_12109);
nor U12775 (N_12775,N_12357,N_12185);
or U12776 (N_12776,N_12352,N_12375);
and U12777 (N_12777,N_12268,N_12258);
nand U12778 (N_12778,N_12303,N_12388);
and U12779 (N_12779,N_12233,N_12363);
and U12780 (N_12780,N_12072,N_12329);
or U12781 (N_12781,N_12106,N_12144);
xor U12782 (N_12782,N_12185,N_12386);
nand U12783 (N_12783,N_12333,N_12340);
nor U12784 (N_12784,N_12207,N_12269);
nor U12785 (N_12785,N_12154,N_12272);
xnor U12786 (N_12786,N_12343,N_12205);
or U12787 (N_12787,N_12193,N_12188);
nor U12788 (N_12788,N_12351,N_12050);
or U12789 (N_12789,N_12062,N_12086);
or U12790 (N_12790,N_12080,N_12163);
and U12791 (N_12791,N_12171,N_12210);
or U12792 (N_12792,N_12195,N_12271);
or U12793 (N_12793,N_12254,N_12036);
xor U12794 (N_12794,N_12231,N_12278);
and U12795 (N_12795,N_12081,N_12023);
xnor U12796 (N_12796,N_12102,N_12014);
nor U12797 (N_12797,N_12286,N_12066);
nand U12798 (N_12798,N_12395,N_12267);
nor U12799 (N_12799,N_12276,N_12288);
or U12800 (N_12800,N_12768,N_12566);
and U12801 (N_12801,N_12619,N_12775);
and U12802 (N_12802,N_12488,N_12578);
or U12803 (N_12803,N_12766,N_12626);
xnor U12804 (N_12804,N_12494,N_12581);
xor U12805 (N_12805,N_12618,N_12753);
and U12806 (N_12806,N_12634,N_12749);
and U12807 (N_12807,N_12602,N_12695);
or U12808 (N_12808,N_12497,N_12798);
nand U12809 (N_12809,N_12704,N_12452);
and U12810 (N_12810,N_12457,N_12662);
and U12811 (N_12811,N_12633,N_12759);
nand U12812 (N_12812,N_12622,N_12489);
xor U12813 (N_12813,N_12527,N_12482);
nor U12814 (N_12814,N_12792,N_12454);
xor U12815 (N_12815,N_12438,N_12614);
and U12816 (N_12816,N_12673,N_12598);
nand U12817 (N_12817,N_12711,N_12441);
xor U12818 (N_12818,N_12716,N_12642);
nor U12819 (N_12819,N_12537,N_12606);
xor U12820 (N_12820,N_12552,N_12620);
xnor U12821 (N_12821,N_12461,N_12684);
nor U12822 (N_12822,N_12443,N_12594);
nand U12823 (N_12823,N_12465,N_12474);
and U12824 (N_12824,N_12558,N_12706);
nand U12825 (N_12825,N_12669,N_12691);
nand U12826 (N_12826,N_12750,N_12694);
or U12827 (N_12827,N_12425,N_12720);
nor U12828 (N_12828,N_12591,N_12421);
xor U12829 (N_12829,N_12464,N_12540);
and U12830 (N_12830,N_12504,N_12472);
and U12831 (N_12831,N_12685,N_12420);
nor U12832 (N_12832,N_12569,N_12455);
or U12833 (N_12833,N_12616,N_12439);
nand U12834 (N_12834,N_12791,N_12650);
nand U12835 (N_12835,N_12526,N_12430);
and U12836 (N_12836,N_12734,N_12415);
or U12837 (N_12837,N_12479,N_12700);
nor U12838 (N_12838,N_12723,N_12740);
nor U12839 (N_12839,N_12608,N_12646);
nor U12840 (N_12840,N_12764,N_12492);
xor U12841 (N_12841,N_12607,N_12469);
nand U12842 (N_12842,N_12730,N_12551);
or U12843 (N_12843,N_12466,N_12409);
or U12844 (N_12844,N_12681,N_12543);
or U12845 (N_12845,N_12567,N_12468);
xor U12846 (N_12846,N_12408,N_12604);
nand U12847 (N_12847,N_12617,N_12568);
nand U12848 (N_12848,N_12649,N_12529);
nand U12849 (N_12849,N_12476,N_12635);
and U12850 (N_12850,N_12582,N_12583);
nand U12851 (N_12851,N_12776,N_12678);
nand U12852 (N_12852,N_12536,N_12784);
xor U12853 (N_12853,N_12667,N_12697);
or U12854 (N_12854,N_12771,N_12689);
or U12855 (N_12855,N_12419,N_12495);
and U12856 (N_12856,N_12613,N_12609);
nor U12857 (N_12857,N_12571,N_12687);
nand U12858 (N_12858,N_12570,N_12629);
nand U12859 (N_12859,N_12541,N_12718);
and U12860 (N_12860,N_12799,N_12450);
xnor U12861 (N_12861,N_12444,N_12757);
nand U12862 (N_12862,N_12714,N_12755);
nor U12863 (N_12863,N_12721,N_12564);
nand U12864 (N_12864,N_12493,N_12535);
or U12865 (N_12865,N_12590,N_12789);
nand U12866 (N_12866,N_12478,N_12502);
nand U12867 (N_12867,N_12625,N_12402);
xnor U12868 (N_12868,N_12675,N_12555);
nand U12869 (N_12869,N_12440,N_12525);
or U12870 (N_12870,N_12656,N_12507);
and U12871 (N_12871,N_12505,N_12756);
or U12872 (N_12872,N_12696,N_12434);
and U12873 (N_12873,N_12795,N_12702);
nor U12874 (N_12874,N_12418,N_12615);
nor U12875 (N_12875,N_12778,N_12719);
nand U12876 (N_12876,N_12772,N_12705);
nor U12877 (N_12877,N_12773,N_12530);
xor U12878 (N_12878,N_12788,N_12751);
and U12879 (N_12879,N_12400,N_12793);
xnor U12880 (N_12880,N_12477,N_12761);
nor U12881 (N_12881,N_12576,N_12542);
and U12882 (N_12882,N_12524,N_12729);
nor U12883 (N_12883,N_12636,N_12501);
nand U12884 (N_12884,N_12644,N_12545);
nor U12885 (N_12885,N_12484,N_12514);
nand U12886 (N_12886,N_12538,N_12404);
xnor U12887 (N_12887,N_12796,N_12426);
xor U12888 (N_12888,N_12442,N_12413);
nor U12889 (N_12889,N_12496,N_12630);
or U12890 (N_12890,N_12447,N_12786);
nor U12891 (N_12891,N_12417,N_12645);
and U12892 (N_12892,N_12648,N_12470);
xor U12893 (N_12893,N_12412,N_12676);
or U12894 (N_12894,N_12429,N_12544);
or U12895 (N_12895,N_12592,N_12547);
or U12896 (N_12896,N_12411,N_12448);
nor U12897 (N_12897,N_12491,N_12782);
and U12898 (N_12898,N_12549,N_12522);
or U12899 (N_12899,N_12638,N_12783);
and U12900 (N_12900,N_12774,N_12679);
nor U12901 (N_12901,N_12785,N_12473);
or U12902 (N_12902,N_12588,N_12428);
nand U12903 (N_12903,N_12713,N_12692);
nor U12904 (N_12904,N_12610,N_12556);
nor U12905 (N_12905,N_12456,N_12666);
or U12906 (N_12906,N_12769,N_12672);
and U12907 (N_12907,N_12765,N_12518);
nand U12908 (N_12908,N_12603,N_12739);
and U12909 (N_12909,N_12690,N_12657);
or U12910 (N_12910,N_12715,N_12532);
nand U12911 (N_12911,N_12490,N_12637);
or U12912 (N_12912,N_12708,N_12698);
nor U12913 (N_12913,N_12741,N_12480);
or U12914 (N_12914,N_12560,N_12737);
xnor U12915 (N_12915,N_12674,N_12742);
or U12916 (N_12916,N_12520,N_12762);
or U12917 (N_12917,N_12611,N_12748);
nor U12918 (N_12918,N_12665,N_12758);
nand U12919 (N_12919,N_12760,N_12410);
and U12920 (N_12920,N_12462,N_12595);
nor U12921 (N_12921,N_12565,N_12521);
or U12922 (N_12922,N_12458,N_12597);
nand U12923 (N_12923,N_12660,N_12601);
nor U12924 (N_12924,N_12643,N_12780);
and U12925 (N_12925,N_12531,N_12652);
nor U12926 (N_12926,N_12509,N_12627);
and U12927 (N_12927,N_12746,N_12677);
and U12928 (N_12928,N_12471,N_12767);
or U12929 (N_12929,N_12743,N_12516);
nor U12930 (N_12930,N_12580,N_12640);
and U12931 (N_12931,N_12572,N_12671);
or U12932 (N_12932,N_12453,N_12574);
or U12933 (N_12933,N_12423,N_12724);
xor U12934 (N_12934,N_12550,N_12658);
nor U12935 (N_12935,N_12513,N_12651);
or U12936 (N_12936,N_12585,N_12770);
xnor U12937 (N_12937,N_12639,N_12414);
xor U12938 (N_12938,N_12699,N_12432);
and U12939 (N_12939,N_12463,N_12703);
and U12940 (N_12940,N_12794,N_12779);
nor U12941 (N_12941,N_12406,N_12736);
nor U12942 (N_12942,N_12459,N_12435);
nand U12943 (N_12943,N_12486,N_12733);
or U12944 (N_12944,N_12573,N_12722);
and U12945 (N_12945,N_12424,N_12562);
or U12946 (N_12946,N_12707,N_12559);
and U12947 (N_12947,N_12523,N_12460);
nand U12948 (N_12948,N_12500,N_12483);
or U12949 (N_12949,N_12589,N_12534);
and U12950 (N_12950,N_12731,N_12744);
nor U12951 (N_12951,N_12709,N_12519);
nand U12952 (N_12952,N_12451,N_12510);
xnor U12953 (N_12953,N_12754,N_12427);
nand U12954 (N_12954,N_12431,N_12624);
nand U12955 (N_12955,N_12664,N_12403);
or U12956 (N_12956,N_12499,N_12686);
xor U12957 (N_12957,N_12584,N_12683);
nor U12958 (N_12958,N_12632,N_12732);
nand U12959 (N_12959,N_12512,N_12670);
and U12960 (N_12960,N_12710,N_12745);
nand U12961 (N_12961,N_12481,N_12485);
or U12962 (N_12962,N_12680,N_12747);
or U12963 (N_12963,N_12668,N_12623);
xnor U12964 (N_12964,N_12449,N_12790);
xor U12965 (N_12965,N_12659,N_12561);
nor U12966 (N_12966,N_12548,N_12475);
nor U12967 (N_12967,N_12612,N_12647);
xnor U12968 (N_12968,N_12599,N_12554);
or U12969 (N_12969,N_12787,N_12605);
nand U12970 (N_12970,N_12577,N_12416);
or U12971 (N_12971,N_12628,N_12655);
nor U12972 (N_12972,N_12553,N_12436);
or U12973 (N_12973,N_12506,N_12641);
nor U12974 (N_12974,N_12797,N_12735);
or U12975 (N_12975,N_12433,N_12517);
nor U12976 (N_12976,N_12487,N_12407);
xnor U12977 (N_12977,N_12728,N_12717);
nor U12978 (N_12978,N_12701,N_12563);
nor U12979 (N_12979,N_12533,N_12586);
nand U12980 (N_12980,N_12725,N_12682);
nand U12981 (N_12981,N_12726,N_12546);
xor U12982 (N_12982,N_12727,N_12781);
xnor U12983 (N_12983,N_12498,N_12693);
nand U12984 (N_12984,N_12653,N_12446);
or U12985 (N_12985,N_12437,N_12405);
nor U12986 (N_12986,N_12752,N_12528);
or U12987 (N_12987,N_12663,N_12593);
or U12988 (N_12988,N_12596,N_12738);
xnor U12989 (N_12989,N_12445,N_12712);
nand U12990 (N_12990,N_12557,N_12688);
nor U12991 (N_12991,N_12763,N_12401);
or U12992 (N_12992,N_12579,N_12515);
and U12993 (N_12993,N_12631,N_12661);
xnor U12994 (N_12994,N_12621,N_12575);
and U12995 (N_12995,N_12654,N_12511);
nand U12996 (N_12996,N_12539,N_12467);
nor U12997 (N_12997,N_12587,N_12600);
or U12998 (N_12998,N_12422,N_12503);
nor U12999 (N_12999,N_12508,N_12777);
or U13000 (N_13000,N_12691,N_12794);
nand U13001 (N_13001,N_12411,N_12413);
nor U13002 (N_13002,N_12532,N_12595);
nor U13003 (N_13003,N_12431,N_12646);
or U13004 (N_13004,N_12470,N_12678);
nand U13005 (N_13005,N_12772,N_12515);
nor U13006 (N_13006,N_12774,N_12586);
nor U13007 (N_13007,N_12669,N_12689);
nand U13008 (N_13008,N_12448,N_12798);
and U13009 (N_13009,N_12501,N_12417);
xnor U13010 (N_13010,N_12571,N_12489);
nand U13011 (N_13011,N_12703,N_12433);
or U13012 (N_13012,N_12457,N_12732);
xor U13013 (N_13013,N_12470,N_12659);
xnor U13014 (N_13014,N_12538,N_12470);
nor U13015 (N_13015,N_12774,N_12491);
or U13016 (N_13016,N_12497,N_12476);
or U13017 (N_13017,N_12752,N_12641);
or U13018 (N_13018,N_12561,N_12679);
or U13019 (N_13019,N_12707,N_12494);
and U13020 (N_13020,N_12687,N_12445);
nor U13021 (N_13021,N_12469,N_12571);
nand U13022 (N_13022,N_12577,N_12653);
or U13023 (N_13023,N_12587,N_12690);
and U13024 (N_13024,N_12792,N_12749);
xnor U13025 (N_13025,N_12664,N_12419);
or U13026 (N_13026,N_12754,N_12419);
and U13027 (N_13027,N_12462,N_12533);
or U13028 (N_13028,N_12774,N_12705);
and U13029 (N_13029,N_12421,N_12621);
nor U13030 (N_13030,N_12518,N_12691);
or U13031 (N_13031,N_12631,N_12573);
nand U13032 (N_13032,N_12793,N_12564);
and U13033 (N_13033,N_12502,N_12788);
and U13034 (N_13034,N_12413,N_12727);
or U13035 (N_13035,N_12662,N_12444);
xnor U13036 (N_13036,N_12466,N_12508);
nor U13037 (N_13037,N_12681,N_12775);
nand U13038 (N_13038,N_12593,N_12436);
nand U13039 (N_13039,N_12679,N_12769);
nand U13040 (N_13040,N_12597,N_12769);
nand U13041 (N_13041,N_12686,N_12497);
nand U13042 (N_13042,N_12797,N_12769);
xor U13043 (N_13043,N_12770,N_12724);
and U13044 (N_13044,N_12792,N_12579);
nand U13045 (N_13045,N_12553,N_12539);
or U13046 (N_13046,N_12636,N_12498);
and U13047 (N_13047,N_12605,N_12511);
xnor U13048 (N_13048,N_12523,N_12731);
nand U13049 (N_13049,N_12513,N_12643);
nor U13050 (N_13050,N_12626,N_12754);
nor U13051 (N_13051,N_12750,N_12459);
and U13052 (N_13052,N_12552,N_12761);
or U13053 (N_13053,N_12425,N_12691);
and U13054 (N_13054,N_12556,N_12449);
or U13055 (N_13055,N_12612,N_12796);
nor U13056 (N_13056,N_12688,N_12489);
or U13057 (N_13057,N_12611,N_12436);
xnor U13058 (N_13058,N_12518,N_12419);
xor U13059 (N_13059,N_12405,N_12550);
or U13060 (N_13060,N_12739,N_12775);
or U13061 (N_13061,N_12489,N_12591);
nand U13062 (N_13062,N_12536,N_12679);
nand U13063 (N_13063,N_12725,N_12795);
xnor U13064 (N_13064,N_12640,N_12562);
and U13065 (N_13065,N_12712,N_12489);
xnor U13066 (N_13066,N_12515,N_12767);
nor U13067 (N_13067,N_12614,N_12622);
nor U13068 (N_13068,N_12473,N_12650);
nand U13069 (N_13069,N_12746,N_12476);
xnor U13070 (N_13070,N_12706,N_12673);
nand U13071 (N_13071,N_12432,N_12497);
nand U13072 (N_13072,N_12404,N_12602);
nand U13073 (N_13073,N_12443,N_12424);
and U13074 (N_13074,N_12548,N_12595);
or U13075 (N_13075,N_12757,N_12503);
xor U13076 (N_13076,N_12429,N_12622);
or U13077 (N_13077,N_12699,N_12725);
or U13078 (N_13078,N_12724,N_12718);
or U13079 (N_13079,N_12618,N_12527);
nor U13080 (N_13080,N_12450,N_12611);
and U13081 (N_13081,N_12694,N_12769);
nor U13082 (N_13082,N_12763,N_12400);
nand U13083 (N_13083,N_12762,N_12723);
nand U13084 (N_13084,N_12413,N_12685);
xor U13085 (N_13085,N_12600,N_12512);
xor U13086 (N_13086,N_12481,N_12559);
xnor U13087 (N_13087,N_12433,N_12601);
and U13088 (N_13088,N_12786,N_12622);
nand U13089 (N_13089,N_12440,N_12686);
xnor U13090 (N_13090,N_12692,N_12510);
nand U13091 (N_13091,N_12617,N_12642);
and U13092 (N_13092,N_12524,N_12786);
and U13093 (N_13093,N_12408,N_12665);
or U13094 (N_13094,N_12622,N_12658);
xnor U13095 (N_13095,N_12579,N_12430);
nand U13096 (N_13096,N_12489,N_12402);
nand U13097 (N_13097,N_12706,N_12552);
nand U13098 (N_13098,N_12516,N_12448);
nor U13099 (N_13099,N_12561,N_12609);
or U13100 (N_13100,N_12721,N_12703);
nand U13101 (N_13101,N_12599,N_12428);
nand U13102 (N_13102,N_12704,N_12483);
xnor U13103 (N_13103,N_12554,N_12721);
or U13104 (N_13104,N_12728,N_12473);
nor U13105 (N_13105,N_12516,N_12624);
nand U13106 (N_13106,N_12739,N_12522);
and U13107 (N_13107,N_12651,N_12622);
and U13108 (N_13108,N_12594,N_12751);
and U13109 (N_13109,N_12500,N_12417);
or U13110 (N_13110,N_12765,N_12579);
and U13111 (N_13111,N_12780,N_12543);
nand U13112 (N_13112,N_12764,N_12585);
and U13113 (N_13113,N_12477,N_12745);
nand U13114 (N_13114,N_12595,N_12416);
nor U13115 (N_13115,N_12510,N_12425);
xnor U13116 (N_13116,N_12644,N_12739);
nor U13117 (N_13117,N_12405,N_12487);
nor U13118 (N_13118,N_12639,N_12710);
nand U13119 (N_13119,N_12677,N_12414);
and U13120 (N_13120,N_12560,N_12606);
or U13121 (N_13121,N_12627,N_12587);
xor U13122 (N_13122,N_12714,N_12428);
and U13123 (N_13123,N_12471,N_12644);
or U13124 (N_13124,N_12479,N_12435);
and U13125 (N_13125,N_12431,N_12539);
and U13126 (N_13126,N_12616,N_12717);
and U13127 (N_13127,N_12549,N_12423);
nor U13128 (N_13128,N_12484,N_12536);
nor U13129 (N_13129,N_12528,N_12666);
and U13130 (N_13130,N_12666,N_12736);
nor U13131 (N_13131,N_12754,N_12596);
nor U13132 (N_13132,N_12738,N_12409);
or U13133 (N_13133,N_12662,N_12756);
nor U13134 (N_13134,N_12546,N_12760);
nor U13135 (N_13135,N_12404,N_12596);
xnor U13136 (N_13136,N_12489,N_12452);
or U13137 (N_13137,N_12506,N_12630);
or U13138 (N_13138,N_12638,N_12511);
xnor U13139 (N_13139,N_12757,N_12746);
nand U13140 (N_13140,N_12555,N_12463);
xor U13141 (N_13141,N_12453,N_12694);
nor U13142 (N_13142,N_12624,N_12567);
nor U13143 (N_13143,N_12706,N_12456);
nor U13144 (N_13144,N_12667,N_12778);
nor U13145 (N_13145,N_12587,N_12685);
xor U13146 (N_13146,N_12594,N_12742);
or U13147 (N_13147,N_12667,N_12740);
xnor U13148 (N_13148,N_12429,N_12734);
or U13149 (N_13149,N_12452,N_12517);
nand U13150 (N_13150,N_12581,N_12648);
nor U13151 (N_13151,N_12426,N_12477);
or U13152 (N_13152,N_12524,N_12503);
nand U13153 (N_13153,N_12783,N_12672);
nand U13154 (N_13154,N_12735,N_12601);
and U13155 (N_13155,N_12660,N_12753);
nand U13156 (N_13156,N_12798,N_12485);
nor U13157 (N_13157,N_12731,N_12556);
or U13158 (N_13158,N_12466,N_12568);
xor U13159 (N_13159,N_12595,N_12673);
and U13160 (N_13160,N_12517,N_12451);
xor U13161 (N_13161,N_12798,N_12665);
nor U13162 (N_13162,N_12563,N_12508);
or U13163 (N_13163,N_12755,N_12561);
and U13164 (N_13164,N_12775,N_12655);
xnor U13165 (N_13165,N_12404,N_12787);
and U13166 (N_13166,N_12589,N_12451);
or U13167 (N_13167,N_12488,N_12718);
nor U13168 (N_13168,N_12731,N_12481);
or U13169 (N_13169,N_12513,N_12430);
nor U13170 (N_13170,N_12578,N_12442);
or U13171 (N_13171,N_12584,N_12746);
nand U13172 (N_13172,N_12658,N_12648);
and U13173 (N_13173,N_12607,N_12648);
xnor U13174 (N_13174,N_12736,N_12537);
nand U13175 (N_13175,N_12690,N_12681);
xor U13176 (N_13176,N_12563,N_12728);
nor U13177 (N_13177,N_12400,N_12765);
xor U13178 (N_13178,N_12762,N_12508);
and U13179 (N_13179,N_12538,N_12534);
nand U13180 (N_13180,N_12778,N_12551);
nand U13181 (N_13181,N_12697,N_12775);
nand U13182 (N_13182,N_12683,N_12719);
nand U13183 (N_13183,N_12522,N_12734);
nor U13184 (N_13184,N_12441,N_12741);
nor U13185 (N_13185,N_12461,N_12588);
or U13186 (N_13186,N_12602,N_12656);
xor U13187 (N_13187,N_12784,N_12679);
xor U13188 (N_13188,N_12435,N_12710);
xor U13189 (N_13189,N_12698,N_12554);
xnor U13190 (N_13190,N_12570,N_12498);
xor U13191 (N_13191,N_12525,N_12513);
and U13192 (N_13192,N_12650,N_12469);
or U13193 (N_13193,N_12412,N_12702);
or U13194 (N_13194,N_12583,N_12608);
xor U13195 (N_13195,N_12629,N_12463);
and U13196 (N_13196,N_12481,N_12473);
and U13197 (N_13197,N_12640,N_12445);
and U13198 (N_13198,N_12702,N_12469);
nor U13199 (N_13199,N_12407,N_12446);
nand U13200 (N_13200,N_12927,N_13198);
or U13201 (N_13201,N_12916,N_13031);
xor U13202 (N_13202,N_13125,N_13005);
xor U13203 (N_13203,N_12826,N_13008);
or U13204 (N_13204,N_12896,N_13123);
or U13205 (N_13205,N_13121,N_12821);
nor U13206 (N_13206,N_13174,N_12893);
or U13207 (N_13207,N_12935,N_12862);
or U13208 (N_13208,N_13185,N_13016);
and U13209 (N_13209,N_13180,N_12960);
xor U13210 (N_13210,N_12998,N_13143);
xor U13211 (N_13211,N_13086,N_13095);
or U13212 (N_13212,N_13151,N_13149);
or U13213 (N_13213,N_13052,N_13085);
or U13214 (N_13214,N_13136,N_12802);
and U13215 (N_13215,N_12973,N_12990);
xnor U13216 (N_13216,N_12995,N_13043);
nor U13217 (N_13217,N_13128,N_13000);
or U13218 (N_13218,N_12808,N_12909);
xnor U13219 (N_13219,N_12817,N_12866);
nand U13220 (N_13220,N_13059,N_12987);
nor U13221 (N_13221,N_12875,N_13058);
and U13222 (N_13222,N_12843,N_12848);
or U13223 (N_13223,N_13036,N_13178);
nand U13224 (N_13224,N_12977,N_13044);
nand U13225 (N_13225,N_13153,N_13120);
and U13226 (N_13226,N_13080,N_13155);
nor U13227 (N_13227,N_13173,N_13161);
or U13228 (N_13228,N_13041,N_13199);
or U13229 (N_13229,N_13145,N_12822);
nor U13230 (N_13230,N_13187,N_13147);
nand U13231 (N_13231,N_12984,N_12865);
nand U13232 (N_13232,N_13159,N_13137);
xnor U13233 (N_13233,N_13148,N_12912);
and U13234 (N_13234,N_13109,N_13091);
nand U13235 (N_13235,N_12938,N_12873);
and U13236 (N_13236,N_12810,N_13133);
nand U13237 (N_13237,N_12887,N_13119);
nand U13238 (N_13238,N_12807,N_13167);
nor U13239 (N_13239,N_13077,N_12829);
xnor U13240 (N_13240,N_12971,N_12853);
xnor U13241 (N_13241,N_12936,N_12823);
or U13242 (N_13242,N_13009,N_13152);
and U13243 (N_13243,N_12950,N_13154);
or U13244 (N_13244,N_13027,N_13038);
or U13245 (N_13245,N_13090,N_12918);
and U13246 (N_13246,N_12937,N_13045);
nor U13247 (N_13247,N_13103,N_12898);
nand U13248 (N_13248,N_12851,N_13061);
and U13249 (N_13249,N_13017,N_12943);
nor U13250 (N_13250,N_12888,N_12827);
nor U13251 (N_13251,N_12922,N_12884);
xor U13252 (N_13252,N_12994,N_13189);
nand U13253 (N_13253,N_13093,N_12815);
xor U13254 (N_13254,N_13078,N_13081);
nor U13255 (N_13255,N_13050,N_12871);
and U13256 (N_13256,N_13066,N_13165);
and U13257 (N_13257,N_12881,N_12805);
xor U13258 (N_13258,N_12889,N_12835);
or U13259 (N_13259,N_12902,N_12814);
and U13260 (N_13260,N_12868,N_13113);
nor U13261 (N_13261,N_12955,N_12944);
or U13262 (N_13262,N_13042,N_13089);
or U13263 (N_13263,N_13131,N_13194);
xnor U13264 (N_13264,N_12852,N_12906);
nand U13265 (N_13265,N_12818,N_13169);
or U13266 (N_13266,N_13019,N_12953);
xnor U13267 (N_13267,N_12919,N_13073);
and U13268 (N_13268,N_12804,N_12886);
and U13269 (N_13269,N_12964,N_12904);
and U13270 (N_13270,N_13141,N_12933);
xnor U13271 (N_13271,N_13063,N_13029);
nand U13272 (N_13272,N_12882,N_13030);
or U13273 (N_13273,N_13138,N_13060);
nor U13274 (N_13274,N_12983,N_13157);
nand U13275 (N_13275,N_13182,N_13076);
nor U13276 (N_13276,N_13162,N_12966);
nor U13277 (N_13277,N_12980,N_13082);
or U13278 (N_13278,N_12917,N_13134);
or U13279 (N_13279,N_12908,N_13057);
or U13280 (N_13280,N_13135,N_13156);
nand U13281 (N_13281,N_13075,N_13101);
and U13282 (N_13282,N_13014,N_13195);
nor U13283 (N_13283,N_12856,N_12969);
xor U13284 (N_13284,N_13018,N_12877);
or U13285 (N_13285,N_13188,N_12883);
nand U13286 (N_13286,N_12861,N_13102);
nand U13287 (N_13287,N_12842,N_13107);
nand U13288 (N_13288,N_12874,N_12974);
xor U13289 (N_13289,N_12924,N_13183);
xnor U13290 (N_13290,N_12981,N_13003);
nor U13291 (N_13291,N_12858,N_12905);
and U13292 (N_13292,N_12870,N_13158);
nand U13293 (N_13293,N_12867,N_13186);
nand U13294 (N_13294,N_13055,N_13142);
or U13295 (N_13295,N_13111,N_13022);
and U13296 (N_13296,N_12907,N_12920);
or U13297 (N_13297,N_13065,N_12869);
nand U13298 (N_13298,N_13098,N_12812);
xor U13299 (N_13299,N_13124,N_12986);
nand U13300 (N_13300,N_12876,N_13172);
nand U13301 (N_13301,N_12976,N_13049);
and U13302 (N_13302,N_12985,N_12885);
xnor U13303 (N_13303,N_13072,N_12975);
or U13304 (N_13304,N_12849,N_13079);
or U13305 (N_13305,N_12838,N_12962);
and U13306 (N_13306,N_13074,N_12982);
and U13307 (N_13307,N_13023,N_13177);
nand U13308 (N_13308,N_13071,N_13032);
nor U13309 (N_13309,N_12941,N_12844);
and U13310 (N_13310,N_12967,N_12839);
or U13311 (N_13311,N_12999,N_12993);
or U13312 (N_13312,N_13037,N_13164);
xnor U13313 (N_13313,N_13114,N_13004);
nor U13314 (N_13314,N_13013,N_12897);
nand U13315 (N_13315,N_13006,N_13115);
nor U13316 (N_13316,N_12928,N_12951);
xnor U13317 (N_13317,N_13092,N_13070);
and U13318 (N_13318,N_12949,N_13139);
or U13319 (N_13319,N_12830,N_13051);
and U13320 (N_13320,N_12952,N_12940);
or U13321 (N_13321,N_13034,N_13068);
or U13322 (N_13322,N_12854,N_12946);
nor U13323 (N_13323,N_13021,N_12819);
xnor U13324 (N_13324,N_12824,N_13160);
and U13325 (N_13325,N_13025,N_13190);
and U13326 (N_13326,N_13012,N_13094);
xor U13327 (N_13327,N_13083,N_13104);
xnor U13328 (N_13328,N_12925,N_13140);
xnor U13329 (N_13329,N_12978,N_12846);
xor U13330 (N_13330,N_13196,N_12947);
xnor U13331 (N_13331,N_12880,N_12892);
or U13332 (N_13332,N_12934,N_12872);
xnor U13333 (N_13333,N_13179,N_12948);
and U13334 (N_13334,N_12942,N_12864);
or U13335 (N_13335,N_13106,N_12970);
nor U13336 (N_13336,N_12837,N_13110);
nand U13337 (N_13337,N_12855,N_13002);
and U13338 (N_13338,N_13181,N_13132);
and U13339 (N_13339,N_13117,N_13105);
nor U13340 (N_13340,N_12988,N_13112);
xnor U13341 (N_13341,N_12836,N_13171);
or U13342 (N_13342,N_13062,N_12956);
xnor U13343 (N_13343,N_12991,N_13011);
and U13344 (N_13344,N_13166,N_12800);
nor U13345 (N_13345,N_12923,N_13067);
nor U13346 (N_13346,N_12930,N_13064);
and U13347 (N_13347,N_13020,N_12914);
nand U13348 (N_13348,N_12813,N_12857);
xnor U13349 (N_13349,N_12894,N_12911);
or U13350 (N_13350,N_13087,N_13024);
and U13351 (N_13351,N_13168,N_12891);
or U13352 (N_13352,N_12828,N_12965);
and U13353 (N_13353,N_12820,N_13069);
nand U13354 (N_13354,N_12895,N_12913);
nor U13355 (N_13355,N_13039,N_12859);
and U13356 (N_13356,N_13193,N_13197);
or U13357 (N_13357,N_12929,N_12841);
xnor U13358 (N_13358,N_13053,N_13126);
or U13359 (N_13359,N_12958,N_13088);
nand U13360 (N_13360,N_12879,N_12921);
or U13361 (N_13361,N_12963,N_12900);
xnor U13362 (N_13362,N_12860,N_13116);
nor U13363 (N_13363,N_13129,N_13118);
and U13364 (N_13364,N_12878,N_13127);
nand U13365 (N_13365,N_13084,N_12903);
xor U13366 (N_13366,N_12945,N_12992);
nor U13367 (N_13367,N_12850,N_12845);
nor U13368 (N_13368,N_12831,N_12915);
xnor U13369 (N_13369,N_12954,N_13175);
nor U13370 (N_13370,N_13047,N_13046);
nand U13371 (N_13371,N_13028,N_12834);
xor U13372 (N_13372,N_12809,N_13097);
or U13373 (N_13373,N_12863,N_13146);
nor U13374 (N_13374,N_12811,N_12847);
and U13375 (N_13375,N_13056,N_13144);
and U13376 (N_13376,N_13150,N_13176);
xnor U13377 (N_13377,N_12931,N_12901);
or U13378 (N_13378,N_13191,N_13001);
and U13379 (N_13379,N_13040,N_12806);
and U13380 (N_13380,N_13099,N_12816);
nor U13381 (N_13381,N_13163,N_12832);
nor U13382 (N_13382,N_13170,N_12996);
or U13383 (N_13383,N_12825,N_13108);
nor U13384 (N_13384,N_12961,N_13048);
xnor U13385 (N_13385,N_13192,N_13130);
or U13386 (N_13386,N_12972,N_12890);
nor U13387 (N_13387,N_13007,N_12968);
nand U13388 (N_13388,N_12989,N_13035);
nor U13389 (N_13389,N_13184,N_12997);
nor U13390 (N_13390,N_12910,N_13015);
or U13391 (N_13391,N_13096,N_13122);
nor U13392 (N_13392,N_13033,N_12959);
or U13393 (N_13393,N_12932,N_13054);
and U13394 (N_13394,N_12899,N_12939);
and U13395 (N_13395,N_12979,N_12803);
nand U13396 (N_13396,N_13100,N_12833);
nor U13397 (N_13397,N_13010,N_12957);
or U13398 (N_13398,N_13026,N_12801);
nand U13399 (N_13399,N_12840,N_12926);
and U13400 (N_13400,N_12988,N_13109);
or U13401 (N_13401,N_13111,N_13049);
nand U13402 (N_13402,N_12838,N_13040);
and U13403 (N_13403,N_12981,N_13147);
xnor U13404 (N_13404,N_12934,N_12845);
and U13405 (N_13405,N_12902,N_12816);
or U13406 (N_13406,N_12928,N_12967);
or U13407 (N_13407,N_13080,N_12877);
nor U13408 (N_13408,N_13035,N_13121);
nand U13409 (N_13409,N_13053,N_12909);
or U13410 (N_13410,N_12956,N_13154);
nand U13411 (N_13411,N_13185,N_12862);
or U13412 (N_13412,N_13134,N_12928);
nand U13413 (N_13413,N_13078,N_13116);
nor U13414 (N_13414,N_12876,N_12939);
nand U13415 (N_13415,N_12879,N_12997);
and U13416 (N_13416,N_13164,N_12801);
nor U13417 (N_13417,N_13102,N_13139);
or U13418 (N_13418,N_12814,N_13086);
nor U13419 (N_13419,N_12807,N_13053);
and U13420 (N_13420,N_12984,N_12879);
nor U13421 (N_13421,N_12810,N_13155);
nand U13422 (N_13422,N_13154,N_12818);
nand U13423 (N_13423,N_12825,N_13048);
xor U13424 (N_13424,N_13078,N_12899);
xor U13425 (N_13425,N_13172,N_13158);
xnor U13426 (N_13426,N_13010,N_13126);
nand U13427 (N_13427,N_12962,N_12923);
nand U13428 (N_13428,N_12877,N_13123);
and U13429 (N_13429,N_13194,N_13195);
xor U13430 (N_13430,N_13050,N_13007);
nand U13431 (N_13431,N_12941,N_13137);
nand U13432 (N_13432,N_12871,N_12832);
and U13433 (N_13433,N_13069,N_12804);
xor U13434 (N_13434,N_12867,N_13062);
nor U13435 (N_13435,N_13144,N_12931);
nand U13436 (N_13436,N_12836,N_12844);
xnor U13437 (N_13437,N_13105,N_12857);
and U13438 (N_13438,N_12801,N_12940);
and U13439 (N_13439,N_13076,N_13106);
and U13440 (N_13440,N_12848,N_12993);
or U13441 (N_13441,N_13094,N_13042);
xnor U13442 (N_13442,N_13043,N_12890);
nand U13443 (N_13443,N_12901,N_13000);
xnor U13444 (N_13444,N_13039,N_12880);
xor U13445 (N_13445,N_13160,N_12954);
nand U13446 (N_13446,N_12805,N_13124);
and U13447 (N_13447,N_13161,N_13164);
nand U13448 (N_13448,N_13076,N_13048);
and U13449 (N_13449,N_12953,N_13087);
nand U13450 (N_13450,N_13026,N_12837);
nand U13451 (N_13451,N_13097,N_13107);
and U13452 (N_13452,N_12858,N_13075);
or U13453 (N_13453,N_12898,N_13051);
and U13454 (N_13454,N_12955,N_13186);
nor U13455 (N_13455,N_12985,N_13058);
nand U13456 (N_13456,N_13075,N_13198);
nor U13457 (N_13457,N_13192,N_13079);
nor U13458 (N_13458,N_12854,N_12921);
or U13459 (N_13459,N_12930,N_12990);
xor U13460 (N_13460,N_13177,N_12940);
xnor U13461 (N_13461,N_12821,N_13041);
xnor U13462 (N_13462,N_13133,N_13148);
and U13463 (N_13463,N_12829,N_12903);
or U13464 (N_13464,N_12966,N_13156);
nand U13465 (N_13465,N_12924,N_12928);
and U13466 (N_13466,N_12862,N_12849);
nor U13467 (N_13467,N_12835,N_13018);
xor U13468 (N_13468,N_12885,N_13046);
xnor U13469 (N_13469,N_12967,N_12977);
or U13470 (N_13470,N_12823,N_12949);
nor U13471 (N_13471,N_12840,N_12969);
xor U13472 (N_13472,N_12921,N_13061);
nor U13473 (N_13473,N_12812,N_13010);
xnor U13474 (N_13474,N_12953,N_13067);
or U13475 (N_13475,N_12966,N_12968);
xnor U13476 (N_13476,N_12899,N_13058);
and U13477 (N_13477,N_13012,N_12950);
xnor U13478 (N_13478,N_13168,N_13105);
and U13479 (N_13479,N_12910,N_13169);
xnor U13480 (N_13480,N_12859,N_13042);
or U13481 (N_13481,N_12905,N_13015);
nand U13482 (N_13482,N_13027,N_12967);
nand U13483 (N_13483,N_12941,N_13039);
nand U13484 (N_13484,N_13103,N_13177);
or U13485 (N_13485,N_13172,N_13067);
xor U13486 (N_13486,N_12868,N_13095);
nor U13487 (N_13487,N_12992,N_12831);
and U13488 (N_13488,N_13121,N_13070);
or U13489 (N_13489,N_12961,N_13146);
nor U13490 (N_13490,N_12910,N_12967);
or U13491 (N_13491,N_13088,N_12828);
and U13492 (N_13492,N_12984,N_13048);
nand U13493 (N_13493,N_12909,N_12924);
and U13494 (N_13494,N_13196,N_13169);
nor U13495 (N_13495,N_12815,N_13157);
xnor U13496 (N_13496,N_13023,N_13089);
nand U13497 (N_13497,N_13012,N_13193);
or U13498 (N_13498,N_12942,N_12803);
nor U13499 (N_13499,N_12910,N_13069);
or U13500 (N_13500,N_13193,N_13036);
nor U13501 (N_13501,N_13024,N_13112);
xor U13502 (N_13502,N_13013,N_13002);
nand U13503 (N_13503,N_12957,N_12816);
nand U13504 (N_13504,N_12837,N_13105);
xnor U13505 (N_13505,N_13032,N_13004);
nand U13506 (N_13506,N_12873,N_13007);
nand U13507 (N_13507,N_13111,N_12898);
nand U13508 (N_13508,N_13123,N_13022);
and U13509 (N_13509,N_13060,N_12953);
nor U13510 (N_13510,N_12817,N_12823);
or U13511 (N_13511,N_12933,N_13092);
nor U13512 (N_13512,N_13026,N_12826);
nand U13513 (N_13513,N_13155,N_12926);
xnor U13514 (N_13514,N_13083,N_12809);
nand U13515 (N_13515,N_13080,N_13168);
xnor U13516 (N_13516,N_12837,N_13048);
nor U13517 (N_13517,N_12934,N_12933);
nand U13518 (N_13518,N_13042,N_13151);
and U13519 (N_13519,N_13142,N_13109);
nand U13520 (N_13520,N_12892,N_13049);
and U13521 (N_13521,N_12931,N_13078);
nand U13522 (N_13522,N_13158,N_12818);
nor U13523 (N_13523,N_12870,N_13192);
nor U13524 (N_13524,N_13116,N_12980);
and U13525 (N_13525,N_12965,N_13186);
nor U13526 (N_13526,N_12851,N_13108);
or U13527 (N_13527,N_13076,N_12902);
and U13528 (N_13528,N_13045,N_12830);
and U13529 (N_13529,N_13194,N_12816);
or U13530 (N_13530,N_12981,N_12814);
nor U13531 (N_13531,N_12869,N_12873);
nor U13532 (N_13532,N_12840,N_13159);
nand U13533 (N_13533,N_13142,N_12924);
xnor U13534 (N_13534,N_12960,N_13045);
nor U13535 (N_13535,N_12801,N_13034);
or U13536 (N_13536,N_12852,N_13068);
nand U13537 (N_13537,N_13077,N_12851);
and U13538 (N_13538,N_13188,N_12960);
nor U13539 (N_13539,N_12897,N_13146);
or U13540 (N_13540,N_13083,N_13069);
nor U13541 (N_13541,N_12831,N_12957);
xor U13542 (N_13542,N_13199,N_12958);
nand U13543 (N_13543,N_13073,N_12878);
nand U13544 (N_13544,N_13009,N_12857);
xor U13545 (N_13545,N_13088,N_13103);
or U13546 (N_13546,N_13097,N_12949);
or U13547 (N_13547,N_12890,N_13035);
nor U13548 (N_13548,N_12940,N_13009);
and U13549 (N_13549,N_12948,N_12913);
and U13550 (N_13550,N_12871,N_13151);
or U13551 (N_13551,N_12864,N_13199);
and U13552 (N_13552,N_13049,N_13010);
nor U13553 (N_13553,N_12958,N_13081);
and U13554 (N_13554,N_13049,N_13112);
and U13555 (N_13555,N_13143,N_13059);
nand U13556 (N_13556,N_12952,N_13193);
and U13557 (N_13557,N_12960,N_13021);
xnor U13558 (N_13558,N_13164,N_12944);
or U13559 (N_13559,N_12980,N_13167);
or U13560 (N_13560,N_12902,N_13054);
nand U13561 (N_13561,N_12849,N_13104);
nand U13562 (N_13562,N_12895,N_13011);
xnor U13563 (N_13563,N_13162,N_12924);
or U13564 (N_13564,N_13176,N_13040);
nand U13565 (N_13565,N_12954,N_13177);
nand U13566 (N_13566,N_12829,N_12888);
and U13567 (N_13567,N_13187,N_12820);
and U13568 (N_13568,N_13013,N_12952);
xnor U13569 (N_13569,N_13015,N_13067);
xnor U13570 (N_13570,N_12812,N_12893);
or U13571 (N_13571,N_13163,N_12954);
xor U13572 (N_13572,N_13052,N_13125);
nor U13573 (N_13573,N_12975,N_13102);
or U13574 (N_13574,N_13027,N_12850);
nand U13575 (N_13575,N_12963,N_13147);
or U13576 (N_13576,N_13023,N_12889);
and U13577 (N_13577,N_12923,N_12871);
xnor U13578 (N_13578,N_12983,N_13119);
nor U13579 (N_13579,N_12965,N_13004);
xor U13580 (N_13580,N_13152,N_13116);
nand U13581 (N_13581,N_13070,N_13024);
or U13582 (N_13582,N_12972,N_13126);
nand U13583 (N_13583,N_12948,N_13159);
or U13584 (N_13584,N_12800,N_13104);
or U13585 (N_13585,N_13102,N_12931);
nor U13586 (N_13586,N_12850,N_13136);
and U13587 (N_13587,N_12906,N_12950);
or U13588 (N_13588,N_13133,N_13019);
nand U13589 (N_13589,N_13158,N_13109);
nand U13590 (N_13590,N_13013,N_13044);
nand U13591 (N_13591,N_12998,N_13138);
nor U13592 (N_13592,N_12873,N_13180);
or U13593 (N_13593,N_13155,N_13063);
or U13594 (N_13594,N_12981,N_13192);
or U13595 (N_13595,N_12865,N_12854);
or U13596 (N_13596,N_12899,N_13129);
nor U13597 (N_13597,N_13084,N_13106);
xnor U13598 (N_13598,N_12985,N_13074);
nor U13599 (N_13599,N_13090,N_13069);
and U13600 (N_13600,N_13462,N_13567);
xor U13601 (N_13601,N_13565,N_13375);
nand U13602 (N_13602,N_13449,N_13555);
nand U13603 (N_13603,N_13478,N_13350);
nor U13604 (N_13604,N_13303,N_13274);
and U13605 (N_13605,N_13558,N_13212);
nor U13606 (N_13606,N_13517,N_13559);
nor U13607 (N_13607,N_13439,N_13522);
nand U13608 (N_13608,N_13442,N_13473);
xnor U13609 (N_13609,N_13214,N_13236);
nor U13610 (N_13610,N_13286,N_13532);
and U13611 (N_13611,N_13505,N_13344);
or U13612 (N_13612,N_13431,N_13351);
or U13613 (N_13613,N_13382,N_13346);
or U13614 (N_13614,N_13409,N_13363);
and U13615 (N_13615,N_13432,N_13593);
or U13616 (N_13616,N_13483,N_13299);
or U13617 (N_13617,N_13407,N_13334);
nand U13618 (N_13618,N_13383,N_13541);
nand U13619 (N_13619,N_13571,N_13368);
and U13620 (N_13620,N_13598,N_13211);
xor U13621 (N_13621,N_13531,N_13373);
and U13622 (N_13622,N_13279,N_13437);
or U13623 (N_13623,N_13465,N_13513);
nand U13624 (N_13624,N_13496,N_13448);
nor U13625 (N_13625,N_13525,N_13592);
nor U13626 (N_13626,N_13302,N_13335);
xnor U13627 (N_13627,N_13219,N_13262);
nor U13628 (N_13628,N_13464,N_13200);
nand U13629 (N_13629,N_13440,N_13342);
or U13630 (N_13630,N_13239,N_13340);
and U13631 (N_13631,N_13562,N_13281);
and U13632 (N_13632,N_13206,N_13284);
or U13633 (N_13633,N_13394,N_13282);
nand U13634 (N_13634,N_13570,N_13597);
and U13635 (N_13635,N_13402,N_13378);
nor U13636 (N_13636,N_13248,N_13201);
or U13637 (N_13637,N_13307,N_13450);
or U13638 (N_13638,N_13263,N_13313);
nand U13639 (N_13639,N_13452,N_13495);
nor U13640 (N_13640,N_13438,N_13546);
nand U13641 (N_13641,N_13332,N_13535);
xnor U13642 (N_13642,N_13228,N_13243);
xor U13643 (N_13643,N_13494,N_13434);
nand U13644 (N_13644,N_13456,N_13360);
and U13645 (N_13645,N_13331,N_13226);
xnor U13646 (N_13646,N_13466,N_13249);
nand U13647 (N_13647,N_13428,N_13581);
xor U13648 (N_13648,N_13575,N_13547);
or U13649 (N_13649,N_13359,N_13485);
xnor U13650 (N_13650,N_13347,N_13328);
and U13651 (N_13651,N_13451,N_13543);
and U13652 (N_13652,N_13361,N_13572);
xor U13653 (N_13653,N_13512,N_13493);
nor U13654 (N_13654,N_13396,N_13523);
nor U13655 (N_13655,N_13553,N_13395);
nand U13656 (N_13656,N_13362,N_13519);
and U13657 (N_13657,N_13476,N_13413);
xnor U13658 (N_13658,N_13242,N_13253);
xnor U13659 (N_13659,N_13492,N_13227);
and U13660 (N_13660,N_13251,N_13549);
nor U13661 (N_13661,N_13424,N_13540);
and U13662 (N_13662,N_13579,N_13345);
xnor U13663 (N_13663,N_13468,N_13422);
and U13664 (N_13664,N_13416,N_13502);
nand U13665 (N_13665,N_13415,N_13392);
nand U13666 (N_13666,N_13386,N_13270);
xnor U13667 (N_13667,N_13480,N_13235);
nor U13668 (N_13668,N_13315,N_13290);
nor U13669 (N_13669,N_13229,N_13365);
or U13670 (N_13670,N_13305,N_13268);
and U13671 (N_13671,N_13204,N_13588);
xor U13672 (N_13672,N_13246,N_13323);
nor U13673 (N_13673,N_13387,N_13410);
or U13674 (N_13674,N_13300,N_13427);
or U13675 (N_13675,N_13591,N_13234);
or U13676 (N_13676,N_13528,N_13520);
nand U13677 (N_13677,N_13599,N_13319);
or U13678 (N_13678,N_13459,N_13534);
nand U13679 (N_13679,N_13475,N_13258);
or U13680 (N_13680,N_13418,N_13423);
nand U13681 (N_13681,N_13306,N_13288);
and U13682 (N_13682,N_13544,N_13318);
nand U13683 (N_13683,N_13557,N_13232);
or U13684 (N_13684,N_13230,N_13587);
nand U13685 (N_13685,N_13568,N_13467);
nor U13686 (N_13686,N_13436,N_13533);
nor U13687 (N_13687,N_13421,N_13419);
and U13688 (N_13688,N_13316,N_13356);
or U13689 (N_13689,N_13329,N_13218);
or U13690 (N_13690,N_13393,N_13381);
nand U13691 (N_13691,N_13370,N_13577);
or U13692 (N_13692,N_13404,N_13384);
or U13693 (N_13693,N_13231,N_13510);
nor U13694 (N_13694,N_13330,N_13297);
and U13695 (N_13695,N_13414,N_13515);
and U13696 (N_13696,N_13397,N_13489);
or U13697 (N_13697,N_13576,N_13398);
xor U13698 (N_13698,N_13560,N_13526);
xnor U13699 (N_13699,N_13324,N_13596);
xnor U13700 (N_13700,N_13245,N_13585);
nand U13701 (N_13701,N_13474,N_13429);
xnor U13702 (N_13702,N_13304,N_13321);
nand U13703 (N_13703,N_13376,N_13314);
xor U13704 (N_13704,N_13203,N_13275);
nand U13705 (N_13705,N_13590,N_13222);
or U13706 (N_13706,N_13269,N_13417);
and U13707 (N_13707,N_13457,N_13582);
nor U13708 (N_13708,N_13453,N_13385);
or U13709 (N_13709,N_13529,N_13287);
and U13710 (N_13710,N_13339,N_13564);
nand U13711 (N_13711,N_13390,N_13511);
and U13712 (N_13712,N_13447,N_13482);
or U13713 (N_13713,N_13471,N_13430);
or U13714 (N_13714,N_13488,N_13561);
nor U13715 (N_13715,N_13556,N_13355);
nand U13716 (N_13716,N_13366,N_13477);
and U13717 (N_13717,N_13272,N_13291);
nor U13718 (N_13718,N_13244,N_13213);
and U13719 (N_13719,N_13372,N_13551);
and U13720 (N_13720,N_13259,N_13285);
and U13721 (N_13721,N_13516,N_13354);
nor U13722 (N_13722,N_13518,N_13472);
or U13723 (N_13723,N_13377,N_13460);
xnor U13724 (N_13724,N_13357,N_13504);
or U13725 (N_13725,N_13371,N_13374);
nor U13726 (N_13726,N_13389,N_13276);
and U13727 (N_13727,N_13349,N_13224);
xnor U13728 (N_13728,N_13257,N_13348);
xnor U13729 (N_13729,N_13469,N_13539);
nand U13730 (N_13730,N_13310,N_13209);
or U13731 (N_13731,N_13484,N_13364);
and U13732 (N_13732,N_13580,N_13479);
or U13733 (N_13733,N_13283,N_13278);
xor U13734 (N_13734,N_13341,N_13406);
nor U13735 (N_13735,N_13503,N_13205);
nand U13736 (N_13736,N_13490,N_13216);
or U13737 (N_13737,N_13481,N_13501);
and U13738 (N_13738,N_13552,N_13458);
nand U13739 (N_13739,N_13260,N_13352);
and U13740 (N_13740,N_13554,N_13238);
or U13741 (N_13741,N_13542,N_13207);
nor U13742 (N_13742,N_13507,N_13426);
and U13743 (N_13743,N_13367,N_13536);
or U13744 (N_13744,N_13595,N_13233);
or U13745 (N_13745,N_13548,N_13566);
nor U13746 (N_13746,N_13264,N_13309);
xnor U13747 (N_13747,N_13240,N_13358);
nor U13748 (N_13748,N_13261,N_13210);
xor U13749 (N_13749,N_13301,N_13399);
xnor U13750 (N_13750,N_13320,N_13538);
nor U13751 (N_13751,N_13594,N_13308);
nand U13752 (N_13752,N_13509,N_13454);
nand U13753 (N_13753,N_13225,N_13223);
xnor U13754 (N_13754,N_13435,N_13250);
nand U13755 (N_13755,N_13208,N_13470);
or U13756 (N_13756,N_13545,N_13217);
or U13757 (N_13757,N_13338,N_13498);
xor U13758 (N_13758,N_13506,N_13569);
xor U13759 (N_13759,N_13312,N_13521);
xnor U13760 (N_13760,N_13491,N_13343);
nand U13761 (N_13761,N_13292,N_13563);
nor U13762 (N_13762,N_13527,N_13322);
nand U13763 (N_13763,N_13369,N_13586);
nand U13764 (N_13764,N_13441,N_13550);
xor U13765 (N_13765,N_13220,N_13271);
xnor U13766 (N_13766,N_13241,N_13405);
xor U13767 (N_13767,N_13277,N_13508);
or U13768 (N_13768,N_13411,N_13336);
nand U13769 (N_13769,N_13514,N_13353);
nand U13770 (N_13770,N_13295,N_13379);
and U13771 (N_13771,N_13412,N_13486);
nand U13772 (N_13772,N_13433,N_13497);
nand U13773 (N_13773,N_13443,N_13391);
nor U13774 (N_13774,N_13267,N_13455);
nor U13775 (N_13775,N_13326,N_13254);
or U13776 (N_13776,N_13294,N_13237);
xnor U13777 (N_13777,N_13325,N_13289);
xor U13778 (N_13778,N_13524,N_13589);
nor U13779 (N_13779,N_13298,N_13425);
and U13780 (N_13780,N_13247,N_13583);
xnor U13781 (N_13781,N_13296,N_13293);
nor U13782 (N_13782,N_13420,N_13273);
or U13783 (N_13783,N_13499,N_13445);
xor U13784 (N_13784,N_13333,N_13380);
xor U13785 (N_13785,N_13317,N_13401);
and U13786 (N_13786,N_13574,N_13400);
nand U13787 (N_13787,N_13255,N_13202);
nor U13788 (N_13788,N_13463,N_13578);
or U13789 (N_13789,N_13403,N_13584);
nand U13790 (N_13790,N_13215,N_13537);
or U13791 (N_13791,N_13265,N_13388);
nand U13792 (N_13792,N_13408,N_13221);
nand U13793 (N_13793,N_13530,N_13500);
nand U13794 (N_13794,N_13280,N_13444);
xnor U13795 (N_13795,N_13252,N_13266);
nor U13796 (N_13796,N_13256,N_13461);
and U13797 (N_13797,N_13327,N_13311);
nand U13798 (N_13798,N_13337,N_13487);
xor U13799 (N_13799,N_13446,N_13573);
xnor U13800 (N_13800,N_13333,N_13547);
and U13801 (N_13801,N_13426,N_13347);
or U13802 (N_13802,N_13523,N_13510);
or U13803 (N_13803,N_13247,N_13375);
nand U13804 (N_13804,N_13461,N_13310);
nor U13805 (N_13805,N_13376,N_13307);
or U13806 (N_13806,N_13578,N_13272);
nand U13807 (N_13807,N_13467,N_13266);
or U13808 (N_13808,N_13377,N_13489);
nor U13809 (N_13809,N_13520,N_13312);
or U13810 (N_13810,N_13524,N_13596);
nor U13811 (N_13811,N_13225,N_13407);
nand U13812 (N_13812,N_13526,N_13554);
xnor U13813 (N_13813,N_13230,N_13424);
xnor U13814 (N_13814,N_13491,N_13312);
or U13815 (N_13815,N_13431,N_13347);
and U13816 (N_13816,N_13371,N_13466);
xnor U13817 (N_13817,N_13272,N_13533);
and U13818 (N_13818,N_13282,N_13510);
nor U13819 (N_13819,N_13379,N_13233);
and U13820 (N_13820,N_13483,N_13215);
and U13821 (N_13821,N_13352,N_13336);
nor U13822 (N_13822,N_13253,N_13334);
or U13823 (N_13823,N_13522,N_13536);
and U13824 (N_13824,N_13428,N_13297);
or U13825 (N_13825,N_13408,N_13528);
nand U13826 (N_13826,N_13276,N_13472);
or U13827 (N_13827,N_13356,N_13299);
xor U13828 (N_13828,N_13253,N_13341);
and U13829 (N_13829,N_13224,N_13597);
or U13830 (N_13830,N_13335,N_13398);
nor U13831 (N_13831,N_13587,N_13413);
and U13832 (N_13832,N_13587,N_13519);
xnor U13833 (N_13833,N_13432,N_13450);
or U13834 (N_13834,N_13568,N_13525);
nor U13835 (N_13835,N_13276,N_13227);
xnor U13836 (N_13836,N_13593,N_13468);
or U13837 (N_13837,N_13454,N_13287);
nor U13838 (N_13838,N_13524,N_13474);
or U13839 (N_13839,N_13313,N_13581);
xnor U13840 (N_13840,N_13228,N_13233);
xnor U13841 (N_13841,N_13226,N_13531);
or U13842 (N_13842,N_13371,N_13363);
and U13843 (N_13843,N_13376,N_13377);
and U13844 (N_13844,N_13392,N_13568);
nor U13845 (N_13845,N_13297,N_13383);
and U13846 (N_13846,N_13559,N_13525);
xnor U13847 (N_13847,N_13295,N_13582);
nor U13848 (N_13848,N_13324,N_13582);
nor U13849 (N_13849,N_13352,N_13299);
xnor U13850 (N_13850,N_13288,N_13562);
nand U13851 (N_13851,N_13358,N_13540);
and U13852 (N_13852,N_13596,N_13390);
nor U13853 (N_13853,N_13461,N_13436);
nand U13854 (N_13854,N_13292,N_13519);
nor U13855 (N_13855,N_13209,N_13555);
and U13856 (N_13856,N_13370,N_13349);
xor U13857 (N_13857,N_13398,N_13548);
xnor U13858 (N_13858,N_13513,N_13358);
nand U13859 (N_13859,N_13461,N_13393);
nor U13860 (N_13860,N_13408,N_13527);
nand U13861 (N_13861,N_13508,N_13530);
nand U13862 (N_13862,N_13365,N_13302);
nor U13863 (N_13863,N_13518,N_13443);
xnor U13864 (N_13864,N_13438,N_13354);
and U13865 (N_13865,N_13527,N_13582);
nor U13866 (N_13866,N_13318,N_13534);
nand U13867 (N_13867,N_13202,N_13305);
and U13868 (N_13868,N_13455,N_13217);
and U13869 (N_13869,N_13271,N_13391);
or U13870 (N_13870,N_13492,N_13472);
or U13871 (N_13871,N_13472,N_13330);
nor U13872 (N_13872,N_13341,N_13598);
nand U13873 (N_13873,N_13221,N_13307);
and U13874 (N_13874,N_13344,N_13298);
and U13875 (N_13875,N_13595,N_13458);
xor U13876 (N_13876,N_13576,N_13545);
nor U13877 (N_13877,N_13209,N_13358);
xor U13878 (N_13878,N_13494,N_13543);
nand U13879 (N_13879,N_13230,N_13273);
nor U13880 (N_13880,N_13450,N_13541);
or U13881 (N_13881,N_13377,N_13352);
nand U13882 (N_13882,N_13336,N_13229);
nor U13883 (N_13883,N_13220,N_13259);
nand U13884 (N_13884,N_13271,N_13200);
and U13885 (N_13885,N_13599,N_13325);
nor U13886 (N_13886,N_13325,N_13421);
nor U13887 (N_13887,N_13203,N_13519);
nand U13888 (N_13888,N_13255,N_13343);
nand U13889 (N_13889,N_13550,N_13365);
or U13890 (N_13890,N_13474,N_13203);
nor U13891 (N_13891,N_13321,N_13527);
and U13892 (N_13892,N_13284,N_13247);
or U13893 (N_13893,N_13403,N_13477);
or U13894 (N_13894,N_13445,N_13436);
nand U13895 (N_13895,N_13266,N_13530);
xnor U13896 (N_13896,N_13574,N_13295);
nand U13897 (N_13897,N_13424,N_13244);
or U13898 (N_13898,N_13260,N_13244);
or U13899 (N_13899,N_13236,N_13255);
nor U13900 (N_13900,N_13576,N_13378);
and U13901 (N_13901,N_13588,N_13451);
nor U13902 (N_13902,N_13550,N_13487);
nor U13903 (N_13903,N_13274,N_13234);
xor U13904 (N_13904,N_13367,N_13339);
or U13905 (N_13905,N_13244,N_13265);
and U13906 (N_13906,N_13419,N_13467);
nand U13907 (N_13907,N_13540,N_13535);
and U13908 (N_13908,N_13479,N_13263);
or U13909 (N_13909,N_13295,N_13487);
or U13910 (N_13910,N_13269,N_13446);
and U13911 (N_13911,N_13493,N_13255);
nand U13912 (N_13912,N_13525,N_13505);
and U13913 (N_13913,N_13348,N_13279);
nand U13914 (N_13914,N_13521,N_13425);
nand U13915 (N_13915,N_13348,N_13410);
nor U13916 (N_13916,N_13541,N_13322);
nand U13917 (N_13917,N_13348,N_13304);
nand U13918 (N_13918,N_13417,N_13500);
nor U13919 (N_13919,N_13424,N_13576);
and U13920 (N_13920,N_13409,N_13432);
xor U13921 (N_13921,N_13398,N_13491);
xor U13922 (N_13922,N_13207,N_13358);
xnor U13923 (N_13923,N_13243,N_13527);
nand U13924 (N_13924,N_13303,N_13427);
and U13925 (N_13925,N_13477,N_13537);
or U13926 (N_13926,N_13583,N_13369);
nor U13927 (N_13927,N_13208,N_13415);
and U13928 (N_13928,N_13225,N_13313);
nand U13929 (N_13929,N_13213,N_13250);
or U13930 (N_13930,N_13227,N_13597);
xnor U13931 (N_13931,N_13491,N_13300);
nor U13932 (N_13932,N_13257,N_13513);
xor U13933 (N_13933,N_13392,N_13208);
and U13934 (N_13934,N_13346,N_13208);
and U13935 (N_13935,N_13318,N_13240);
nor U13936 (N_13936,N_13517,N_13573);
nand U13937 (N_13937,N_13428,N_13555);
xnor U13938 (N_13938,N_13538,N_13476);
nand U13939 (N_13939,N_13591,N_13307);
or U13940 (N_13940,N_13271,N_13414);
or U13941 (N_13941,N_13444,N_13572);
nor U13942 (N_13942,N_13464,N_13342);
and U13943 (N_13943,N_13339,N_13389);
nand U13944 (N_13944,N_13474,N_13355);
nand U13945 (N_13945,N_13392,N_13517);
or U13946 (N_13946,N_13311,N_13540);
nand U13947 (N_13947,N_13224,N_13356);
xor U13948 (N_13948,N_13319,N_13211);
nand U13949 (N_13949,N_13515,N_13398);
nor U13950 (N_13950,N_13549,N_13314);
xor U13951 (N_13951,N_13245,N_13227);
xor U13952 (N_13952,N_13592,N_13200);
or U13953 (N_13953,N_13428,N_13479);
xnor U13954 (N_13954,N_13430,N_13456);
nor U13955 (N_13955,N_13517,N_13566);
and U13956 (N_13956,N_13359,N_13501);
nand U13957 (N_13957,N_13597,N_13384);
xor U13958 (N_13958,N_13241,N_13438);
nand U13959 (N_13959,N_13597,N_13254);
nor U13960 (N_13960,N_13251,N_13499);
or U13961 (N_13961,N_13345,N_13550);
and U13962 (N_13962,N_13512,N_13254);
nand U13963 (N_13963,N_13457,N_13320);
xnor U13964 (N_13964,N_13401,N_13212);
and U13965 (N_13965,N_13570,N_13508);
and U13966 (N_13966,N_13473,N_13335);
nand U13967 (N_13967,N_13459,N_13350);
xnor U13968 (N_13968,N_13290,N_13566);
xor U13969 (N_13969,N_13439,N_13313);
and U13970 (N_13970,N_13526,N_13420);
nand U13971 (N_13971,N_13372,N_13378);
or U13972 (N_13972,N_13205,N_13341);
nor U13973 (N_13973,N_13207,N_13516);
nand U13974 (N_13974,N_13477,N_13516);
nand U13975 (N_13975,N_13526,N_13446);
nand U13976 (N_13976,N_13416,N_13533);
nor U13977 (N_13977,N_13236,N_13478);
nor U13978 (N_13978,N_13225,N_13446);
nand U13979 (N_13979,N_13516,N_13339);
or U13980 (N_13980,N_13433,N_13569);
xnor U13981 (N_13981,N_13232,N_13210);
or U13982 (N_13982,N_13319,N_13517);
xor U13983 (N_13983,N_13391,N_13287);
xnor U13984 (N_13984,N_13498,N_13434);
nor U13985 (N_13985,N_13529,N_13598);
and U13986 (N_13986,N_13303,N_13405);
nand U13987 (N_13987,N_13383,N_13395);
or U13988 (N_13988,N_13238,N_13431);
or U13989 (N_13989,N_13525,N_13323);
nor U13990 (N_13990,N_13449,N_13387);
xor U13991 (N_13991,N_13491,N_13378);
and U13992 (N_13992,N_13415,N_13386);
xor U13993 (N_13993,N_13554,N_13411);
xor U13994 (N_13994,N_13453,N_13498);
or U13995 (N_13995,N_13435,N_13212);
nor U13996 (N_13996,N_13265,N_13262);
xor U13997 (N_13997,N_13573,N_13451);
xnor U13998 (N_13998,N_13351,N_13570);
and U13999 (N_13999,N_13480,N_13465);
and U14000 (N_14000,N_13977,N_13703);
nand U14001 (N_14001,N_13695,N_13995);
xor U14002 (N_14002,N_13798,N_13710);
nor U14003 (N_14003,N_13910,N_13832);
and U14004 (N_14004,N_13766,N_13824);
or U14005 (N_14005,N_13749,N_13634);
nor U14006 (N_14006,N_13854,N_13905);
xnor U14007 (N_14007,N_13946,N_13731);
xor U14008 (N_14008,N_13717,N_13663);
nor U14009 (N_14009,N_13902,N_13688);
or U14010 (N_14010,N_13778,N_13967);
xnor U14011 (N_14011,N_13779,N_13654);
nand U14012 (N_14012,N_13785,N_13775);
nand U14013 (N_14013,N_13940,N_13857);
nand U14014 (N_14014,N_13895,N_13974);
and U14015 (N_14015,N_13860,N_13852);
nand U14016 (N_14016,N_13845,N_13755);
xnor U14017 (N_14017,N_13738,N_13791);
nor U14018 (N_14018,N_13614,N_13605);
nand U14019 (N_14019,N_13632,N_13835);
nand U14020 (N_14020,N_13891,N_13963);
nor U14021 (N_14021,N_13828,N_13748);
and U14022 (N_14022,N_13647,N_13660);
nand U14023 (N_14023,N_13990,N_13999);
xor U14024 (N_14024,N_13689,N_13783);
or U14025 (N_14025,N_13867,N_13697);
or U14026 (N_14026,N_13822,N_13800);
and U14027 (N_14027,N_13741,N_13880);
nand U14028 (N_14028,N_13737,N_13613);
nand U14029 (N_14029,N_13997,N_13769);
and U14030 (N_14030,N_13865,N_13996);
and U14031 (N_14031,N_13933,N_13991);
or U14032 (N_14032,N_13674,N_13621);
and U14033 (N_14033,N_13984,N_13883);
nand U14034 (N_14034,N_13774,N_13941);
nor U14035 (N_14035,N_13809,N_13793);
xor U14036 (N_14036,N_13978,N_13842);
or U14037 (N_14037,N_13698,N_13623);
and U14038 (N_14038,N_13758,N_13707);
nand U14039 (N_14039,N_13627,N_13912);
and U14040 (N_14040,N_13616,N_13976);
nand U14041 (N_14041,N_13722,N_13730);
xor U14042 (N_14042,N_13924,N_13615);
and U14043 (N_14043,N_13879,N_13643);
nand U14044 (N_14044,N_13840,N_13992);
nor U14045 (N_14045,N_13848,N_13813);
and U14046 (N_14046,N_13770,N_13786);
or U14047 (N_14047,N_13931,N_13952);
xnor U14048 (N_14048,N_13752,N_13728);
nor U14049 (N_14049,N_13885,N_13921);
nor U14050 (N_14050,N_13636,N_13890);
and U14051 (N_14051,N_13907,N_13768);
nor U14052 (N_14052,N_13911,N_13641);
xnor U14053 (N_14053,N_13829,N_13837);
and U14054 (N_14054,N_13670,N_13713);
nor U14055 (N_14055,N_13987,N_13882);
xnor U14056 (N_14056,N_13716,N_13754);
or U14057 (N_14057,N_13724,N_13900);
nand U14058 (N_14058,N_13757,N_13954);
and U14059 (N_14059,N_13934,N_13745);
nor U14060 (N_14060,N_13711,N_13795);
and U14061 (N_14061,N_13998,N_13781);
nand U14062 (N_14062,N_13847,N_13734);
or U14063 (N_14063,N_13985,N_13986);
or U14064 (N_14064,N_13676,N_13659);
and U14065 (N_14065,N_13973,N_13846);
xnor U14066 (N_14066,N_13815,N_13638);
and U14067 (N_14067,N_13886,N_13953);
nand U14068 (N_14068,N_13942,N_13756);
and U14069 (N_14069,N_13718,N_13988);
nor U14070 (N_14070,N_13858,N_13762);
or U14071 (N_14071,N_13893,N_13979);
nand U14072 (N_14072,N_13826,N_13620);
and U14073 (N_14073,N_13935,N_13746);
or U14074 (N_14074,N_13888,N_13792);
and U14075 (N_14075,N_13794,N_13936);
and U14076 (N_14076,N_13819,N_13980);
and U14077 (N_14077,N_13628,N_13773);
nand U14078 (N_14078,N_13830,N_13971);
nor U14079 (N_14079,N_13972,N_13807);
or U14080 (N_14080,N_13721,N_13646);
xor U14081 (N_14081,N_13831,N_13870);
nor U14082 (N_14082,N_13603,N_13960);
and U14083 (N_14083,N_13926,N_13648);
or U14084 (N_14084,N_13868,N_13771);
and U14085 (N_14085,N_13827,N_13784);
or U14086 (N_14086,N_13622,N_13694);
and U14087 (N_14087,N_13918,N_13661);
or U14088 (N_14088,N_13751,N_13612);
or U14089 (N_14089,N_13704,N_13675);
nor U14090 (N_14090,N_13619,N_13683);
xor U14091 (N_14091,N_13958,N_13602);
and U14092 (N_14092,N_13764,N_13642);
and U14093 (N_14093,N_13962,N_13925);
nand U14094 (N_14094,N_13719,N_13964);
xor U14095 (N_14095,N_13851,N_13617);
xnor U14096 (N_14096,N_13733,N_13650);
or U14097 (N_14097,N_13903,N_13959);
nor U14098 (N_14098,N_13966,N_13631);
nand U14099 (N_14099,N_13677,N_13812);
nand U14100 (N_14100,N_13850,N_13790);
xnor U14101 (N_14101,N_13869,N_13825);
nand U14102 (N_14102,N_13693,N_13801);
and U14103 (N_14103,N_13994,N_13708);
xnor U14104 (N_14104,N_13901,N_13797);
nor U14105 (N_14105,N_13906,N_13706);
or U14106 (N_14106,N_13920,N_13929);
and U14107 (N_14107,N_13908,N_13821);
nand U14108 (N_14108,N_13899,N_13943);
nor U14109 (N_14109,N_13843,N_13653);
and U14110 (N_14110,N_13725,N_13853);
nand U14111 (N_14111,N_13637,N_13604);
xnor U14112 (N_14112,N_13866,N_13889);
and U14113 (N_14113,N_13923,N_13624);
nand U14114 (N_14114,N_13715,N_13665);
xnor U14115 (N_14115,N_13639,N_13606);
xnor U14116 (N_14116,N_13804,N_13836);
and U14117 (N_14117,N_13873,N_13626);
xnor U14118 (N_14118,N_13607,N_13789);
and U14119 (N_14119,N_13818,N_13989);
nand U14120 (N_14120,N_13742,N_13983);
and U14121 (N_14121,N_13914,N_13656);
xnor U14122 (N_14122,N_13814,N_13699);
xnor U14123 (N_14123,N_13823,N_13981);
nand U14124 (N_14124,N_13743,N_13690);
nor U14125 (N_14125,N_13782,N_13961);
or U14126 (N_14126,N_13787,N_13796);
xor U14127 (N_14127,N_13856,N_13610);
nand U14128 (N_14128,N_13937,N_13720);
nor U14129 (N_14129,N_13927,N_13919);
nor U14130 (N_14130,N_13727,N_13965);
nor U14131 (N_14131,N_13601,N_13732);
xor U14132 (N_14132,N_13817,N_13803);
xor U14133 (N_14133,N_13834,N_13687);
or U14134 (N_14134,N_13735,N_13750);
or U14135 (N_14135,N_13916,N_13896);
and U14136 (N_14136,N_13679,N_13609);
or U14137 (N_14137,N_13651,N_13859);
xor U14138 (N_14138,N_13863,N_13714);
xor U14139 (N_14139,N_13608,N_13645);
nand U14140 (N_14140,N_13881,N_13664);
or U14141 (N_14141,N_13633,N_13649);
nor U14142 (N_14142,N_13776,N_13658);
or U14143 (N_14143,N_13874,N_13671);
and U14144 (N_14144,N_13810,N_13662);
xnor U14145 (N_14145,N_13672,N_13682);
xnor U14146 (N_14146,N_13767,N_13898);
nand U14147 (N_14147,N_13932,N_13820);
xor U14148 (N_14148,N_13744,N_13740);
or U14149 (N_14149,N_13894,N_13928);
or U14150 (N_14150,N_13917,N_13666);
or U14151 (N_14151,N_13841,N_13897);
or U14152 (N_14152,N_13669,N_13849);
and U14153 (N_14153,N_13780,N_13944);
nor U14154 (N_14154,N_13839,N_13833);
nand U14155 (N_14155,N_13844,N_13955);
and U14156 (N_14156,N_13957,N_13709);
and U14157 (N_14157,N_13982,N_13763);
and U14158 (N_14158,N_13765,N_13761);
and U14159 (N_14159,N_13805,N_13806);
and U14160 (N_14160,N_13686,N_13700);
and U14161 (N_14161,N_13705,N_13655);
or U14162 (N_14162,N_13951,N_13993);
nor U14163 (N_14163,N_13673,N_13600);
and U14164 (N_14164,N_13876,N_13930);
or U14165 (N_14165,N_13777,N_13652);
xnor U14166 (N_14166,N_13726,N_13945);
nand U14167 (N_14167,N_13802,N_13629);
or U14168 (N_14168,N_13861,N_13939);
and U14169 (N_14169,N_13970,N_13947);
and U14170 (N_14170,N_13838,N_13739);
nand U14171 (N_14171,N_13772,N_13913);
xnor U14172 (N_14172,N_13701,N_13799);
nand U14173 (N_14173,N_13904,N_13681);
xnor U14174 (N_14174,N_13887,N_13692);
nand U14175 (N_14175,N_13788,N_13948);
or U14176 (N_14176,N_13892,N_13667);
and U14177 (N_14177,N_13884,N_13949);
nand U14178 (N_14178,N_13611,N_13685);
nor U14179 (N_14179,N_13968,N_13915);
or U14180 (N_14180,N_13877,N_13691);
nand U14181 (N_14181,N_13875,N_13635);
and U14182 (N_14182,N_13922,N_13640);
nor U14183 (N_14183,N_13680,N_13702);
nor U14184 (N_14184,N_13760,N_13956);
xnor U14185 (N_14185,N_13630,N_13811);
and U14186 (N_14186,N_13736,N_13871);
or U14187 (N_14187,N_13938,N_13684);
nand U14188 (N_14188,N_13950,N_13678);
nor U14189 (N_14189,N_13696,N_13878);
and U14190 (N_14190,N_13729,N_13723);
nand U14191 (N_14191,N_13657,N_13618);
nor U14192 (N_14192,N_13644,N_13909);
and U14193 (N_14193,N_13747,N_13855);
or U14194 (N_14194,N_13969,N_13808);
nor U14195 (N_14195,N_13668,N_13864);
or U14196 (N_14196,N_13975,N_13816);
or U14197 (N_14197,N_13872,N_13759);
and U14198 (N_14198,N_13712,N_13625);
or U14199 (N_14199,N_13753,N_13862);
nor U14200 (N_14200,N_13912,N_13676);
xnor U14201 (N_14201,N_13736,N_13604);
xor U14202 (N_14202,N_13735,N_13892);
or U14203 (N_14203,N_13609,N_13722);
nor U14204 (N_14204,N_13672,N_13649);
xor U14205 (N_14205,N_13907,N_13688);
xnor U14206 (N_14206,N_13656,N_13962);
xor U14207 (N_14207,N_13963,N_13998);
nor U14208 (N_14208,N_13717,N_13669);
nor U14209 (N_14209,N_13680,N_13810);
nand U14210 (N_14210,N_13959,N_13954);
or U14211 (N_14211,N_13895,N_13907);
xnor U14212 (N_14212,N_13612,N_13615);
xor U14213 (N_14213,N_13844,N_13736);
and U14214 (N_14214,N_13668,N_13680);
nor U14215 (N_14215,N_13949,N_13714);
and U14216 (N_14216,N_13725,N_13820);
and U14217 (N_14217,N_13979,N_13675);
or U14218 (N_14218,N_13717,N_13752);
xor U14219 (N_14219,N_13770,N_13789);
or U14220 (N_14220,N_13846,N_13761);
or U14221 (N_14221,N_13700,N_13795);
xor U14222 (N_14222,N_13804,N_13918);
or U14223 (N_14223,N_13687,N_13894);
xnor U14224 (N_14224,N_13798,N_13872);
nor U14225 (N_14225,N_13780,N_13759);
xnor U14226 (N_14226,N_13708,N_13638);
nor U14227 (N_14227,N_13954,N_13627);
and U14228 (N_14228,N_13738,N_13781);
xnor U14229 (N_14229,N_13783,N_13971);
nor U14230 (N_14230,N_13682,N_13958);
nor U14231 (N_14231,N_13832,N_13749);
xor U14232 (N_14232,N_13856,N_13847);
nor U14233 (N_14233,N_13858,N_13866);
xor U14234 (N_14234,N_13615,N_13935);
xnor U14235 (N_14235,N_13802,N_13861);
nand U14236 (N_14236,N_13920,N_13648);
xor U14237 (N_14237,N_13905,N_13998);
and U14238 (N_14238,N_13608,N_13853);
or U14239 (N_14239,N_13996,N_13775);
nand U14240 (N_14240,N_13891,N_13894);
nand U14241 (N_14241,N_13884,N_13769);
or U14242 (N_14242,N_13796,N_13965);
xnor U14243 (N_14243,N_13712,N_13746);
nor U14244 (N_14244,N_13706,N_13984);
nor U14245 (N_14245,N_13874,N_13808);
nand U14246 (N_14246,N_13619,N_13785);
or U14247 (N_14247,N_13700,N_13894);
xor U14248 (N_14248,N_13604,N_13900);
nand U14249 (N_14249,N_13939,N_13849);
nand U14250 (N_14250,N_13734,N_13908);
or U14251 (N_14251,N_13690,N_13763);
xor U14252 (N_14252,N_13686,N_13638);
or U14253 (N_14253,N_13729,N_13604);
and U14254 (N_14254,N_13841,N_13779);
nor U14255 (N_14255,N_13950,N_13815);
and U14256 (N_14256,N_13819,N_13701);
or U14257 (N_14257,N_13688,N_13940);
nor U14258 (N_14258,N_13631,N_13904);
xnor U14259 (N_14259,N_13674,N_13701);
nand U14260 (N_14260,N_13943,N_13733);
or U14261 (N_14261,N_13952,N_13735);
nor U14262 (N_14262,N_13861,N_13947);
nand U14263 (N_14263,N_13624,N_13892);
and U14264 (N_14264,N_13965,N_13687);
nand U14265 (N_14265,N_13988,N_13998);
nand U14266 (N_14266,N_13936,N_13937);
or U14267 (N_14267,N_13878,N_13987);
or U14268 (N_14268,N_13982,N_13770);
nand U14269 (N_14269,N_13841,N_13794);
or U14270 (N_14270,N_13821,N_13865);
xnor U14271 (N_14271,N_13787,N_13730);
or U14272 (N_14272,N_13997,N_13702);
xor U14273 (N_14273,N_13659,N_13807);
xnor U14274 (N_14274,N_13900,N_13631);
and U14275 (N_14275,N_13831,N_13998);
and U14276 (N_14276,N_13856,N_13914);
and U14277 (N_14277,N_13767,N_13813);
or U14278 (N_14278,N_13720,N_13985);
or U14279 (N_14279,N_13941,N_13841);
nor U14280 (N_14280,N_13648,N_13895);
nand U14281 (N_14281,N_13853,N_13994);
nor U14282 (N_14282,N_13806,N_13950);
nand U14283 (N_14283,N_13978,N_13636);
xor U14284 (N_14284,N_13769,N_13726);
or U14285 (N_14285,N_13805,N_13604);
xor U14286 (N_14286,N_13887,N_13953);
or U14287 (N_14287,N_13833,N_13768);
or U14288 (N_14288,N_13756,N_13701);
and U14289 (N_14289,N_13901,N_13699);
and U14290 (N_14290,N_13770,N_13917);
nor U14291 (N_14291,N_13621,N_13650);
and U14292 (N_14292,N_13871,N_13996);
nand U14293 (N_14293,N_13698,N_13717);
or U14294 (N_14294,N_13878,N_13921);
or U14295 (N_14295,N_13944,N_13795);
nand U14296 (N_14296,N_13890,N_13994);
and U14297 (N_14297,N_13696,N_13613);
xor U14298 (N_14298,N_13725,N_13689);
nand U14299 (N_14299,N_13675,N_13877);
or U14300 (N_14300,N_13784,N_13963);
nor U14301 (N_14301,N_13690,N_13760);
nor U14302 (N_14302,N_13665,N_13904);
xor U14303 (N_14303,N_13806,N_13611);
xnor U14304 (N_14304,N_13637,N_13911);
nand U14305 (N_14305,N_13812,N_13994);
xnor U14306 (N_14306,N_13747,N_13655);
and U14307 (N_14307,N_13810,N_13843);
nor U14308 (N_14308,N_13764,N_13682);
xor U14309 (N_14309,N_13777,N_13942);
nand U14310 (N_14310,N_13706,N_13832);
or U14311 (N_14311,N_13619,N_13742);
and U14312 (N_14312,N_13778,N_13873);
nand U14313 (N_14313,N_13712,N_13682);
and U14314 (N_14314,N_13792,N_13806);
nand U14315 (N_14315,N_13691,N_13616);
or U14316 (N_14316,N_13657,N_13611);
xnor U14317 (N_14317,N_13859,N_13836);
and U14318 (N_14318,N_13851,N_13686);
nor U14319 (N_14319,N_13762,N_13730);
or U14320 (N_14320,N_13943,N_13711);
and U14321 (N_14321,N_13600,N_13674);
and U14322 (N_14322,N_13971,N_13677);
xor U14323 (N_14323,N_13829,N_13877);
nor U14324 (N_14324,N_13883,N_13743);
xor U14325 (N_14325,N_13628,N_13977);
nor U14326 (N_14326,N_13713,N_13778);
xnor U14327 (N_14327,N_13869,N_13854);
xor U14328 (N_14328,N_13979,N_13718);
nor U14329 (N_14329,N_13760,N_13959);
nor U14330 (N_14330,N_13886,N_13605);
xnor U14331 (N_14331,N_13724,N_13883);
nand U14332 (N_14332,N_13670,N_13663);
nor U14333 (N_14333,N_13990,N_13900);
and U14334 (N_14334,N_13688,N_13973);
or U14335 (N_14335,N_13629,N_13634);
and U14336 (N_14336,N_13839,N_13841);
nand U14337 (N_14337,N_13936,N_13720);
nor U14338 (N_14338,N_13836,N_13856);
and U14339 (N_14339,N_13939,N_13605);
nor U14340 (N_14340,N_13855,N_13940);
nor U14341 (N_14341,N_13624,N_13994);
nand U14342 (N_14342,N_13864,N_13803);
nor U14343 (N_14343,N_13640,N_13673);
and U14344 (N_14344,N_13877,N_13896);
nor U14345 (N_14345,N_13980,N_13829);
nor U14346 (N_14346,N_13794,N_13986);
nor U14347 (N_14347,N_13659,N_13933);
nand U14348 (N_14348,N_13730,N_13770);
nand U14349 (N_14349,N_13843,N_13687);
or U14350 (N_14350,N_13944,N_13800);
nand U14351 (N_14351,N_13928,N_13738);
nand U14352 (N_14352,N_13867,N_13744);
nor U14353 (N_14353,N_13899,N_13868);
nand U14354 (N_14354,N_13952,N_13719);
nor U14355 (N_14355,N_13758,N_13830);
and U14356 (N_14356,N_13768,N_13772);
and U14357 (N_14357,N_13694,N_13875);
and U14358 (N_14358,N_13793,N_13967);
nor U14359 (N_14359,N_13616,N_13610);
or U14360 (N_14360,N_13954,N_13813);
or U14361 (N_14361,N_13780,N_13891);
or U14362 (N_14362,N_13728,N_13958);
xnor U14363 (N_14363,N_13713,N_13678);
nor U14364 (N_14364,N_13922,N_13968);
and U14365 (N_14365,N_13946,N_13779);
or U14366 (N_14366,N_13809,N_13949);
and U14367 (N_14367,N_13802,N_13913);
nand U14368 (N_14368,N_13731,N_13657);
and U14369 (N_14369,N_13957,N_13775);
xor U14370 (N_14370,N_13772,N_13931);
nand U14371 (N_14371,N_13945,N_13650);
or U14372 (N_14372,N_13997,N_13642);
nand U14373 (N_14373,N_13709,N_13908);
nor U14374 (N_14374,N_13625,N_13788);
or U14375 (N_14375,N_13982,N_13701);
nor U14376 (N_14376,N_13746,N_13675);
and U14377 (N_14377,N_13723,N_13895);
or U14378 (N_14378,N_13913,N_13616);
and U14379 (N_14379,N_13982,N_13790);
or U14380 (N_14380,N_13895,N_13643);
nor U14381 (N_14381,N_13934,N_13809);
nand U14382 (N_14382,N_13635,N_13871);
nor U14383 (N_14383,N_13795,N_13625);
and U14384 (N_14384,N_13817,N_13637);
nand U14385 (N_14385,N_13806,N_13998);
nand U14386 (N_14386,N_13856,N_13788);
nand U14387 (N_14387,N_13642,N_13819);
and U14388 (N_14388,N_13646,N_13732);
xnor U14389 (N_14389,N_13992,N_13651);
nand U14390 (N_14390,N_13908,N_13998);
xnor U14391 (N_14391,N_13876,N_13911);
and U14392 (N_14392,N_13832,N_13956);
nor U14393 (N_14393,N_13711,N_13908);
nand U14394 (N_14394,N_13651,N_13631);
nand U14395 (N_14395,N_13955,N_13843);
nor U14396 (N_14396,N_13802,N_13640);
nor U14397 (N_14397,N_13998,N_13982);
and U14398 (N_14398,N_13742,N_13653);
and U14399 (N_14399,N_13867,N_13650);
or U14400 (N_14400,N_14001,N_14011);
xnor U14401 (N_14401,N_14226,N_14049);
and U14402 (N_14402,N_14197,N_14233);
nand U14403 (N_14403,N_14002,N_14339);
nor U14404 (N_14404,N_14219,N_14315);
nand U14405 (N_14405,N_14034,N_14269);
nand U14406 (N_14406,N_14014,N_14057);
xor U14407 (N_14407,N_14274,N_14341);
nand U14408 (N_14408,N_14060,N_14294);
xor U14409 (N_14409,N_14130,N_14027);
nand U14410 (N_14410,N_14096,N_14129);
and U14411 (N_14411,N_14046,N_14218);
and U14412 (N_14412,N_14352,N_14280);
nand U14413 (N_14413,N_14263,N_14298);
nor U14414 (N_14414,N_14392,N_14330);
or U14415 (N_14415,N_14119,N_14088);
or U14416 (N_14416,N_14191,N_14351);
and U14417 (N_14417,N_14248,N_14094);
and U14418 (N_14418,N_14070,N_14177);
nand U14419 (N_14419,N_14246,N_14319);
xor U14420 (N_14420,N_14005,N_14376);
nor U14421 (N_14421,N_14105,N_14328);
xnor U14422 (N_14422,N_14097,N_14286);
and U14423 (N_14423,N_14116,N_14213);
nand U14424 (N_14424,N_14064,N_14379);
xnor U14425 (N_14425,N_14321,N_14384);
nor U14426 (N_14426,N_14399,N_14290);
nand U14427 (N_14427,N_14056,N_14017);
and U14428 (N_14428,N_14222,N_14388);
nand U14429 (N_14429,N_14131,N_14079);
or U14430 (N_14430,N_14077,N_14291);
nand U14431 (N_14431,N_14053,N_14302);
nor U14432 (N_14432,N_14145,N_14113);
nor U14433 (N_14433,N_14344,N_14036);
and U14434 (N_14434,N_14110,N_14215);
xnor U14435 (N_14435,N_14121,N_14369);
and U14436 (N_14436,N_14041,N_14147);
nand U14437 (N_14437,N_14182,N_14255);
or U14438 (N_14438,N_14163,N_14062);
nand U14439 (N_14439,N_14391,N_14135);
and U14440 (N_14440,N_14155,N_14366);
nor U14441 (N_14441,N_14132,N_14074);
or U14442 (N_14442,N_14223,N_14152);
nand U14443 (N_14443,N_14178,N_14254);
and U14444 (N_14444,N_14196,N_14313);
or U14445 (N_14445,N_14109,N_14349);
xnor U14446 (N_14446,N_14217,N_14043);
or U14447 (N_14447,N_14220,N_14148);
xor U14448 (N_14448,N_14314,N_14000);
nand U14449 (N_14449,N_14111,N_14098);
or U14450 (N_14450,N_14203,N_14021);
xor U14451 (N_14451,N_14040,N_14168);
nor U14452 (N_14452,N_14186,N_14106);
or U14453 (N_14453,N_14125,N_14316);
or U14454 (N_14454,N_14176,N_14342);
nor U14455 (N_14455,N_14347,N_14227);
nand U14456 (N_14456,N_14063,N_14212);
nor U14457 (N_14457,N_14209,N_14237);
or U14458 (N_14458,N_14076,N_14231);
and U14459 (N_14459,N_14066,N_14257);
or U14460 (N_14460,N_14085,N_14229);
xor U14461 (N_14461,N_14193,N_14086);
nand U14462 (N_14462,N_14282,N_14309);
nor U14463 (N_14463,N_14337,N_14236);
nor U14464 (N_14464,N_14181,N_14183);
and U14465 (N_14465,N_14234,N_14007);
and U14466 (N_14466,N_14354,N_14323);
and U14467 (N_14467,N_14245,N_14200);
xnor U14468 (N_14468,N_14170,N_14325);
nor U14469 (N_14469,N_14242,N_14118);
or U14470 (N_14470,N_14382,N_14311);
nor U14471 (N_14471,N_14375,N_14289);
and U14472 (N_14472,N_14358,N_14367);
or U14473 (N_14473,N_14093,N_14346);
or U14474 (N_14474,N_14292,N_14268);
xor U14475 (N_14475,N_14138,N_14159);
or U14476 (N_14476,N_14397,N_14164);
nand U14477 (N_14477,N_14322,N_14338);
nand U14478 (N_14478,N_14238,N_14276);
or U14479 (N_14479,N_14260,N_14241);
nand U14480 (N_14480,N_14089,N_14386);
nor U14481 (N_14481,N_14026,N_14195);
nor U14482 (N_14482,N_14123,N_14146);
nor U14483 (N_14483,N_14144,N_14272);
nor U14484 (N_14484,N_14104,N_14273);
and U14485 (N_14485,N_14004,N_14187);
and U14486 (N_14486,N_14305,N_14381);
and U14487 (N_14487,N_14161,N_14327);
nor U14488 (N_14488,N_14264,N_14301);
xnor U14489 (N_14489,N_14059,N_14265);
or U14490 (N_14490,N_14051,N_14370);
xnor U14491 (N_14491,N_14012,N_14359);
or U14492 (N_14492,N_14133,N_14010);
xnor U14493 (N_14493,N_14283,N_14030);
nand U14494 (N_14494,N_14120,N_14281);
nand U14495 (N_14495,N_14023,N_14253);
nand U14496 (N_14496,N_14162,N_14006);
nand U14497 (N_14497,N_14232,N_14211);
and U14498 (N_14498,N_14340,N_14050);
and U14499 (N_14499,N_14015,N_14297);
or U14500 (N_14500,N_14204,N_14158);
nor U14501 (N_14501,N_14039,N_14154);
nand U14502 (N_14502,N_14172,N_14078);
nand U14503 (N_14503,N_14019,N_14372);
nor U14504 (N_14504,N_14277,N_14320);
or U14505 (N_14505,N_14267,N_14099);
nor U14506 (N_14506,N_14160,N_14380);
nand U14507 (N_14507,N_14084,N_14042);
xor U14508 (N_14508,N_14013,N_14368);
nand U14509 (N_14509,N_14044,N_14312);
xor U14510 (N_14510,N_14115,N_14166);
or U14511 (N_14511,N_14174,N_14091);
nor U14512 (N_14512,N_14167,N_14171);
xor U14513 (N_14513,N_14261,N_14103);
nor U14514 (N_14514,N_14235,N_14072);
xor U14515 (N_14515,N_14045,N_14396);
or U14516 (N_14516,N_14071,N_14208);
xnor U14517 (N_14517,N_14175,N_14390);
xor U14518 (N_14518,N_14357,N_14387);
and U14519 (N_14519,N_14240,N_14033);
nand U14520 (N_14520,N_14134,N_14127);
nor U14521 (N_14521,N_14285,N_14150);
or U14522 (N_14522,N_14249,N_14201);
nor U14523 (N_14523,N_14139,N_14259);
and U14524 (N_14524,N_14081,N_14279);
nand U14525 (N_14525,N_14100,N_14102);
nand U14526 (N_14526,N_14061,N_14136);
xor U14527 (N_14527,N_14028,N_14336);
xnor U14528 (N_14528,N_14124,N_14117);
or U14529 (N_14529,N_14278,N_14024);
nand U14530 (N_14530,N_14216,N_14065);
or U14531 (N_14531,N_14262,N_14304);
and U14532 (N_14532,N_14087,N_14295);
or U14533 (N_14533,N_14225,N_14080);
and U14534 (N_14534,N_14029,N_14244);
and U14535 (N_14535,N_14250,N_14389);
nand U14536 (N_14536,N_14362,N_14032);
xor U14537 (N_14537,N_14108,N_14090);
xnor U14538 (N_14538,N_14334,N_14239);
and U14539 (N_14539,N_14114,N_14035);
or U14540 (N_14540,N_14037,N_14092);
nand U14541 (N_14541,N_14266,N_14069);
nor U14542 (N_14542,N_14317,N_14303);
or U14543 (N_14543,N_14306,N_14149);
nor U14544 (N_14544,N_14271,N_14126);
and U14545 (N_14545,N_14300,N_14307);
nor U14546 (N_14546,N_14350,N_14107);
nor U14547 (N_14547,N_14385,N_14188);
xor U14548 (N_14548,N_14251,N_14202);
and U14549 (N_14549,N_14140,N_14252);
nor U14550 (N_14550,N_14009,N_14169);
xnor U14551 (N_14551,N_14016,N_14355);
xor U14552 (N_14552,N_14363,N_14371);
nor U14553 (N_14553,N_14308,N_14332);
or U14554 (N_14554,N_14398,N_14048);
nand U14555 (N_14555,N_14329,N_14361);
nor U14556 (N_14556,N_14377,N_14345);
and U14557 (N_14557,N_14192,N_14142);
xor U14558 (N_14558,N_14373,N_14270);
and U14559 (N_14559,N_14194,N_14343);
or U14560 (N_14560,N_14364,N_14067);
nor U14561 (N_14561,N_14185,N_14365);
or U14562 (N_14562,N_14189,N_14256);
xnor U14563 (N_14563,N_14157,N_14083);
nor U14564 (N_14564,N_14020,N_14247);
nor U14565 (N_14565,N_14173,N_14331);
nor U14566 (N_14566,N_14275,N_14378);
or U14567 (N_14567,N_14112,N_14333);
xor U14568 (N_14568,N_14224,N_14258);
xor U14569 (N_14569,N_14075,N_14198);
or U14570 (N_14570,N_14205,N_14383);
xnor U14571 (N_14571,N_14151,N_14095);
nor U14572 (N_14572,N_14052,N_14210);
xor U14573 (N_14573,N_14288,N_14393);
and U14574 (N_14574,N_14395,N_14228);
nor U14575 (N_14575,N_14353,N_14287);
nand U14576 (N_14576,N_14141,N_14214);
xor U14577 (N_14577,N_14073,N_14128);
and U14578 (N_14578,N_14068,N_14122);
or U14579 (N_14579,N_14394,N_14047);
nand U14580 (N_14580,N_14082,N_14143);
and U14581 (N_14581,N_14230,N_14324);
xor U14582 (N_14582,N_14101,N_14360);
nand U14583 (N_14583,N_14335,N_14284);
or U14584 (N_14584,N_14031,N_14003);
nor U14585 (N_14585,N_14054,N_14310);
nor U14586 (N_14586,N_14326,N_14180);
nand U14587 (N_14587,N_14207,N_14199);
nor U14588 (N_14588,N_14184,N_14165);
and U14589 (N_14589,N_14221,N_14022);
nor U14590 (N_14590,N_14318,N_14348);
nor U14591 (N_14591,N_14018,N_14299);
nor U14592 (N_14592,N_14243,N_14293);
and U14593 (N_14593,N_14206,N_14058);
nor U14594 (N_14594,N_14008,N_14153);
xor U14595 (N_14595,N_14025,N_14055);
and U14596 (N_14596,N_14190,N_14356);
xnor U14597 (N_14597,N_14137,N_14296);
xor U14598 (N_14598,N_14038,N_14374);
nand U14599 (N_14599,N_14156,N_14179);
nand U14600 (N_14600,N_14311,N_14250);
or U14601 (N_14601,N_14028,N_14224);
nor U14602 (N_14602,N_14321,N_14101);
nor U14603 (N_14603,N_14390,N_14253);
or U14604 (N_14604,N_14059,N_14028);
nor U14605 (N_14605,N_14146,N_14147);
nand U14606 (N_14606,N_14028,N_14073);
xnor U14607 (N_14607,N_14315,N_14323);
xor U14608 (N_14608,N_14298,N_14367);
xnor U14609 (N_14609,N_14351,N_14082);
nor U14610 (N_14610,N_14120,N_14110);
nor U14611 (N_14611,N_14098,N_14049);
nor U14612 (N_14612,N_14158,N_14333);
xnor U14613 (N_14613,N_14314,N_14215);
xnor U14614 (N_14614,N_14258,N_14091);
or U14615 (N_14615,N_14256,N_14080);
nor U14616 (N_14616,N_14319,N_14356);
and U14617 (N_14617,N_14219,N_14011);
or U14618 (N_14618,N_14014,N_14196);
or U14619 (N_14619,N_14187,N_14068);
nand U14620 (N_14620,N_14186,N_14136);
xnor U14621 (N_14621,N_14008,N_14098);
and U14622 (N_14622,N_14292,N_14010);
nor U14623 (N_14623,N_14315,N_14298);
xnor U14624 (N_14624,N_14194,N_14072);
nor U14625 (N_14625,N_14396,N_14037);
nand U14626 (N_14626,N_14133,N_14207);
xor U14627 (N_14627,N_14272,N_14294);
nor U14628 (N_14628,N_14363,N_14072);
nand U14629 (N_14629,N_14303,N_14371);
xnor U14630 (N_14630,N_14193,N_14019);
xnor U14631 (N_14631,N_14156,N_14067);
xnor U14632 (N_14632,N_14254,N_14271);
nand U14633 (N_14633,N_14055,N_14315);
nor U14634 (N_14634,N_14144,N_14032);
nor U14635 (N_14635,N_14351,N_14091);
and U14636 (N_14636,N_14015,N_14236);
nor U14637 (N_14637,N_14296,N_14226);
and U14638 (N_14638,N_14378,N_14331);
xnor U14639 (N_14639,N_14143,N_14301);
nand U14640 (N_14640,N_14374,N_14287);
or U14641 (N_14641,N_14260,N_14056);
nand U14642 (N_14642,N_14337,N_14008);
nor U14643 (N_14643,N_14043,N_14308);
nand U14644 (N_14644,N_14376,N_14370);
nand U14645 (N_14645,N_14399,N_14144);
nor U14646 (N_14646,N_14018,N_14249);
or U14647 (N_14647,N_14273,N_14259);
nor U14648 (N_14648,N_14356,N_14205);
or U14649 (N_14649,N_14302,N_14145);
nor U14650 (N_14650,N_14138,N_14087);
nor U14651 (N_14651,N_14029,N_14376);
and U14652 (N_14652,N_14397,N_14024);
and U14653 (N_14653,N_14077,N_14074);
nor U14654 (N_14654,N_14357,N_14259);
or U14655 (N_14655,N_14025,N_14254);
and U14656 (N_14656,N_14260,N_14214);
nand U14657 (N_14657,N_14057,N_14013);
nand U14658 (N_14658,N_14071,N_14181);
and U14659 (N_14659,N_14030,N_14163);
or U14660 (N_14660,N_14244,N_14053);
or U14661 (N_14661,N_14349,N_14372);
nand U14662 (N_14662,N_14081,N_14271);
or U14663 (N_14663,N_14269,N_14025);
xor U14664 (N_14664,N_14356,N_14176);
or U14665 (N_14665,N_14049,N_14385);
nor U14666 (N_14666,N_14328,N_14155);
xnor U14667 (N_14667,N_14145,N_14337);
nor U14668 (N_14668,N_14075,N_14229);
nor U14669 (N_14669,N_14152,N_14065);
nand U14670 (N_14670,N_14213,N_14128);
and U14671 (N_14671,N_14305,N_14040);
or U14672 (N_14672,N_14133,N_14364);
or U14673 (N_14673,N_14123,N_14250);
nor U14674 (N_14674,N_14249,N_14144);
xnor U14675 (N_14675,N_14024,N_14009);
nand U14676 (N_14676,N_14004,N_14061);
xnor U14677 (N_14677,N_14168,N_14116);
or U14678 (N_14678,N_14146,N_14003);
xor U14679 (N_14679,N_14075,N_14122);
or U14680 (N_14680,N_14128,N_14226);
or U14681 (N_14681,N_14240,N_14383);
or U14682 (N_14682,N_14050,N_14149);
or U14683 (N_14683,N_14249,N_14314);
xor U14684 (N_14684,N_14016,N_14173);
and U14685 (N_14685,N_14149,N_14253);
nand U14686 (N_14686,N_14351,N_14096);
and U14687 (N_14687,N_14268,N_14368);
nor U14688 (N_14688,N_14109,N_14098);
or U14689 (N_14689,N_14274,N_14312);
xnor U14690 (N_14690,N_14050,N_14140);
and U14691 (N_14691,N_14095,N_14079);
nor U14692 (N_14692,N_14276,N_14222);
or U14693 (N_14693,N_14082,N_14276);
nor U14694 (N_14694,N_14083,N_14359);
nand U14695 (N_14695,N_14134,N_14008);
or U14696 (N_14696,N_14395,N_14129);
nor U14697 (N_14697,N_14371,N_14048);
or U14698 (N_14698,N_14040,N_14297);
nand U14699 (N_14699,N_14053,N_14399);
and U14700 (N_14700,N_14046,N_14368);
nand U14701 (N_14701,N_14030,N_14005);
nor U14702 (N_14702,N_14066,N_14221);
or U14703 (N_14703,N_14171,N_14092);
nand U14704 (N_14704,N_14329,N_14009);
xor U14705 (N_14705,N_14152,N_14164);
or U14706 (N_14706,N_14339,N_14336);
xor U14707 (N_14707,N_14342,N_14048);
xnor U14708 (N_14708,N_14344,N_14064);
or U14709 (N_14709,N_14009,N_14281);
or U14710 (N_14710,N_14197,N_14121);
or U14711 (N_14711,N_14257,N_14316);
or U14712 (N_14712,N_14100,N_14087);
nand U14713 (N_14713,N_14031,N_14235);
and U14714 (N_14714,N_14053,N_14212);
and U14715 (N_14715,N_14069,N_14175);
nand U14716 (N_14716,N_14188,N_14096);
or U14717 (N_14717,N_14210,N_14247);
nor U14718 (N_14718,N_14156,N_14377);
nor U14719 (N_14719,N_14152,N_14110);
xor U14720 (N_14720,N_14303,N_14190);
nor U14721 (N_14721,N_14381,N_14015);
or U14722 (N_14722,N_14196,N_14104);
xnor U14723 (N_14723,N_14151,N_14277);
or U14724 (N_14724,N_14015,N_14377);
and U14725 (N_14725,N_14371,N_14201);
and U14726 (N_14726,N_14050,N_14254);
nor U14727 (N_14727,N_14269,N_14115);
nand U14728 (N_14728,N_14342,N_14219);
or U14729 (N_14729,N_14267,N_14061);
and U14730 (N_14730,N_14102,N_14013);
nand U14731 (N_14731,N_14155,N_14078);
xnor U14732 (N_14732,N_14184,N_14190);
xor U14733 (N_14733,N_14164,N_14186);
nor U14734 (N_14734,N_14201,N_14009);
or U14735 (N_14735,N_14068,N_14180);
or U14736 (N_14736,N_14139,N_14154);
or U14737 (N_14737,N_14373,N_14228);
or U14738 (N_14738,N_14160,N_14243);
xnor U14739 (N_14739,N_14274,N_14246);
or U14740 (N_14740,N_14057,N_14047);
nand U14741 (N_14741,N_14305,N_14066);
xnor U14742 (N_14742,N_14293,N_14177);
and U14743 (N_14743,N_14352,N_14218);
nand U14744 (N_14744,N_14336,N_14246);
nor U14745 (N_14745,N_14273,N_14204);
xor U14746 (N_14746,N_14107,N_14062);
nor U14747 (N_14747,N_14206,N_14287);
nand U14748 (N_14748,N_14106,N_14021);
and U14749 (N_14749,N_14101,N_14381);
xnor U14750 (N_14750,N_14054,N_14125);
xor U14751 (N_14751,N_14248,N_14235);
xor U14752 (N_14752,N_14224,N_14211);
xor U14753 (N_14753,N_14083,N_14310);
nor U14754 (N_14754,N_14200,N_14333);
xnor U14755 (N_14755,N_14356,N_14027);
nor U14756 (N_14756,N_14050,N_14141);
nand U14757 (N_14757,N_14054,N_14269);
nor U14758 (N_14758,N_14108,N_14273);
nor U14759 (N_14759,N_14057,N_14258);
or U14760 (N_14760,N_14027,N_14324);
or U14761 (N_14761,N_14041,N_14279);
nor U14762 (N_14762,N_14358,N_14288);
nand U14763 (N_14763,N_14251,N_14342);
nand U14764 (N_14764,N_14024,N_14246);
nor U14765 (N_14765,N_14142,N_14026);
or U14766 (N_14766,N_14051,N_14212);
and U14767 (N_14767,N_14293,N_14252);
nor U14768 (N_14768,N_14059,N_14276);
and U14769 (N_14769,N_14178,N_14245);
or U14770 (N_14770,N_14304,N_14350);
nand U14771 (N_14771,N_14101,N_14158);
nand U14772 (N_14772,N_14399,N_14291);
or U14773 (N_14773,N_14208,N_14206);
nor U14774 (N_14774,N_14264,N_14199);
and U14775 (N_14775,N_14275,N_14294);
xnor U14776 (N_14776,N_14313,N_14125);
or U14777 (N_14777,N_14153,N_14178);
and U14778 (N_14778,N_14360,N_14073);
and U14779 (N_14779,N_14357,N_14075);
nand U14780 (N_14780,N_14023,N_14172);
or U14781 (N_14781,N_14068,N_14207);
and U14782 (N_14782,N_14312,N_14382);
or U14783 (N_14783,N_14091,N_14358);
nor U14784 (N_14784,N_14229,N_14126);
nor U14785 (N_14785,N_14137,N_14088);
nand U14786 (N_14786,N_14040,N_14101);
or U14787 (N_14787,N_14013,N_14157);
or U14788 (N_14788,N_14039,N_14347);
nor U14789 (N_14789,N_14161,N_14054);
and U14790 (N_14790,N_14008,N_14133);
or U14791 (N_14791,N_14099,N_14161);
xor U14792 (N_14792,N_14297,N_14294);
xor U14793 (N_14793,N_14387,N_14197);
xnor U14794 (N_14794,N_14274,N_14120);
nand U14795 (N_14795,N_14312,N_14057);
xor U14796 (N_14796,N_14328,N_14008);
and U14797 (N_14797,N_14148,N_14348);
xnor U14798 (N_14798,N_14017,N_14396);
or U14799 (N_14799,N_14231,N_14336);
xnor U14800 (N_14800,N_14439,N_14726);
nand U14801 (N_14801,N_14590,N_14548);
nor U14802 (N_14802,N_14767,N_14443);
or U14803 (N_14803,N_14445,N_14556);
xor U14804 (N_14804,N_14588,N_14469);
nor U14805 (N_14805,N_14668,N_14665);
nor U14806 (N_14806,N_14483,N_14456);
and U14807 (N_14807,N_14576,N_14538);
xnor U14808 (N_14808,N_14671,N_14698);
or U14809 (N_14809,N_14741,N_14579);
xnor U14810 (N_14810,N_14670,N_14693);
xor U14811 (N_14811,N_14429,N_14787);
nor U14812 (N_14812,N_14617,N_14653);
xor U14813 (N_14813,N_14416,N_14684);
or U14814 (N_14814,N_14449,N_14441);
nand U14815 (N_14815,N_14446,N_14614);
xnor U14816 (N_14816,N_14746,N_14605);
xnor U14817 (N_14817,N_14646,N_14494);
xor U14818 (N_14818,N_14629,N_14453);
xor U14819 (N_14819,N_14474,N_14794);
nor U14820 (N_14820,N_14473,N_14496);
and U14821 (N_14821,N_14448,N_14475);
nand U14822 (N_14822,N_14708,N_14573);
nor U14823 (N_14823,N_14550,N_14751);
nor U14824 (N_14824,N_14768,N_14481);
and U14825 (N_14825,N_14484,N_14509);
or U14826 (N_14826,N_14781,N_14765);
nor U14827 (N_14827,N_14712,N_14485);
xnor U14828 (N_14828,N_14597,N_14709);
or U14829 (N_14829,N_14454,N_14498);
or U14830 (N_14830,N_14707,N_14601);
nand U14831 (N_14831,N_14417,N_14592);
and U14832 (N_14832,N_14557,N_14603);
and U14833 (N_14833,N_14566,N_14716);
and U14834 (N_14834,N_14784,N_14740);
or U14835 (N_14835,N_14559,N_14526);
nor U14836 (N_14836,N_14562,N_14694);
or U14837 (N_14837,N_14774,N_14761);
nand U14838 (N_14838,N_14404,N_14622);
or U14839 (N_14839,N_14535,N_14493);
nor U14840 (N_14840,N_14611,N_14524);
and U14841 (N_14841,N_14422,N_14640);
and U14842 (N_14842,N_14609,N_14489);
nand U14843 (N_14843,N_14459,N_14735);
xnor U14844 (N_14844,N_14683,N_14487);
and U14845 (N_14845,N_14642,N_14599);
and U14846 (N_14846,N_14407,N_14775);
xor U14847 (N_14847,N_14773,N_14516);
nand U14848 (N_14848,N_14447,N_14703);
or U14849 (N_14849,N_14503,N_14744);
nor U14850 (N_14850,N_14674,N_14728);
xor U14851 (N_14851,N_14754,N_14421);
xor U14852 (N_14852,N_14560,N_14772);
nand U14853 (N_14853,N_14687,N_14546);
xor U14854 (N_14854,N_14659,N_14541);
nand U14855 (N_14855,N_14434,N_14507);
or U14856 (N_14856,N_14565,N_14680);
or U14857 (N_14857,N_14467,N_14705);
nor U14858 (N_14858,N_14654,N_14673);
and U14859 (N_14859,N_14762,N_14490);
xor U14860 (N_14860,N_14607,N_14491);
or U14861 (N_14861,N_14410,N_14587);
xor U14862 (N_14862,N_14702,N_14630);
nor U14863 (N_14863,N_14488,N_14661);
and U14864 (N_14864,N_14770,N_14461);
nand U14865 (N_14865,N_14613,N_14499);
and U14866 (N_14866,N_14504,N_14505);
or U14867 (N_14867,N_14413,N_14512);
nand U14868 (N_14868,N_14479,N_14675);
or U14869 (N_14869,N_14433,N_14634);
xnor U14870 (N_14870,N_14732,N_14482);
nor U14871 (N_14871,N_14627,N_14650);
nor U14872 (N_14872,N_14756,N_14570);
xnor U14873 (N_14873,N_14688,N_14706);
or U14874 (N_14874,N_14409,N_14700);
xor U14875 (N_14875,N_14628,N_14760);
xor U14876 (N_14876,N_14666,N_14460);
or U14877 (N_14877,N_14594,N_14604);
and U14878 (N_14878,N_14697,N_14455);
nor U14879 (N_14879,N_14658,N_14518);
xor U14880 (N_14880,N_14465,N_14695);
nand U14881 (N_14881,N_14737,N_14637);
or U14882 (N_14882,N_14739,N_14419);
nor U14883 (N_14883,N_14572,N_14759);
nand U14884 (N_14884,N_14478,N_14633);
xor U14885 (N_14885,N_14452,N_14574);
and U14886 (N_14886,N_14591,N_14791);
nand U14887 (N_14887,N_14644,N_14648);
nor U14888 (N_14888,N_14427,N_14782);
xnor U14889 (N_14889,N_14729,N_14779);
or U14890 (N_14890,N_14625,N_14677);
nor U14891 (N_14891,N_14651,N_14515);
and U14892 (N_14892,N_14508,N_14406);
nand U14893 (N_14893,N_14582,N_14730);
nor U14894 (N_14894,N_14602,N_14797);
xor U14895 (N_14895,N_14401,N_14785);
nand U14896 (N_14896,N_14486,N_14776);
xnor U14897 (N_14897,N_14533,N_14616);
and U14898 (N_14898,N_14529,N_14757);
or U14899 (N_14899,N_14621,N_14636);
or U14900 (N_14900,N_14647,N_14585);
nand U14901 (N_14901,N_14711,N_14721);
xnor U14902 (N_14902,N_14542,N_14436);
xor U14903 (N_14903,N_14631,N_14710);
nor U14904 (N_14904,N_14685,N_14725);
nand U14905 (N_14905,N_14743,N_14718);
or U14906 (N_14906,N_14714,N_14497);
or U14907 (N_14907,N_14742,N_14411);
or U14908 (N_14908,N_14788,N_14750);
xnor U14909 (N_14909,N_14639,N_14662);
xnor U14910 (N_14910,N_14563,N_14495);
nand U14911 (N_14911,N_14564,N_14476);
nor U14912 (N_14912,N_14780,N_14593);
xnor U14913 (N_14913,N_14571,N_14790);
xnor U14914 (N_14914,N_14552,N_14778);
or U14915 (N_14915,N_14462,N_14681);
xnor U14916 (N_14916,N_14736,N_14606);
and U14917 (N_14917,N_14747,N_14466);
or U14918 (N_14918,N_14511,N_14589);
xnor U14919 (N_14919,N_14480,N_14502);
or U14920 (N_14920,N_14428,N_14470);
nand U14921 (N_14921,N_14764,N_14769);
and U14922 (N_14922,N_14715,N_14492);
nor U14923 (N_14923,N_14414,N_14442);
and U14924 (N_14924,N_14690,N_14438);
and U14925 (N_14925,N_14624,N_14405);
xor U14926 (N_14926,N_14667,N_14510);
xnor U14927 (N_14927,N_14412,N_14575);
or U14928 (N_14928,N_14686,N_14522);
and U14929 (N_14929,N_14523,N_14514);
nor U14930 (N_14930,N_14635,N_14766);
nand U14931 (N_14931,N_14596,N_14777);
nand U14932 (N_14932,N_14724,N_14701);
nand U14933 (N_14933,N_14457,N_14420);
or U14934 (N_14934,N_14558,N_14451);
nor U14935 (N_14935,N_14799,N_14643);
and U14936 (N_14936,N_14540,N_14792);
nand U14937 (N_14937,N_14699,N_14795);
and U14938 (N_14938,N_14402,N_14423);
nor U14939 (N_14939,N_14623,N_14672);
and U14940 (N_14940,N_14752,N_14689);
nor U14941 (N_14941,N_14471,N_14657);
and U14942 (N_14942,N_14458,N_14415);
or U14943 (N_14943,N_14444,N_14620);
xnor U14944 (N_14944,N_14612,N_14734);
nand U14945 (N_14945,N_14568,N_14626);
nor U14946 (N_14946,N_14722,N_14638);
or U14947 (N_14947,N_14525,N_14749);
and U14948 (N_14948,N_14440,N_14619);
xnor U14949 (N_14949,N_14437,N_14534);
and U14950 (N_14950,N_14696,N_14472);
nor U14951 (N_14951,N_14679,N_14656);
and U14952 (N_14952,N_14663,N_14745);
or U14953 (N_14953,N_14418,N_14408);
and U14954 (N_14954,N_14727,N_14468);
or U14955 (N_14955,N_14748,N_14555);
nor U14956 (N_14956,N_14581,N_14615);
nand U14957 (N_14957,N_14608,N_14551);
nand U14958 (N_14958,N_14763,N_14669);
or U14959 (N_14959,N_14506,N_14723);
and U14960 (N_14960,N_14691,N_14731);
nor U14961 (N_14961,N_14600,N_14664);
and U14962 (N_14962,N_14513,N_14755);
nand U14963 (N_14963,N_14610,N_14431);
nand U14964 (N_14964,N_14561,N_14539);
xnor U14965 (N_14965,N_14598,N_14719);
or U14966 (N_14966,N_14425,N_14530);
nand U14967 (N_14967,N_14632,N_14584);
and U14968 (N_14968,N_14517,N_14704);
and U14969 (N_14969,N_14583,N_14738);
or U14970 (N_14970,N_14798,N_14578);
nor U14971 (N_14971,N_14586,N_14547);
nor U14972 (N_14972,N_14520,N_14536);
nand U14973 (N_14973,N_14783,N_14676);
nor U14974 (N_14974,N_14758,N_14531);
or U14975 (N_14975,N_14595,N_14521);
and U14976 (N_14976,N_14435,N_14753);
nand U14977 (N_14977,N_14652,N_14464);
nor U14978 (N_14978,N_14477,N_14682);
nor U14979 (N_14979,N_14789,N_14655);
and U14980 (N_14980,N_14426,N_14660);
xor U14981 (N_14981,N_14545,N_14463);
nand U14982 (N_14982,N_14793,N_14430);
nor U14983 (N_14983,N_14527,N_14400);
or U14984 (N_14984,N_14528,N_14553);
nor U14985 (N_14985,N_14649,N_14645);
and U14986 (N_14986,N_14580,N_14537);
or U14987 (N_14987,N_14532,N_14500);
xnor U14988 (N_14988,N_14424,N_14554);
nor U14989 (N_14989,N_14567,N_14403);
and U14990 (N_14990,N_14771,N_14692);
nor U14991 (N_14991,N_14519,N_14733);
xnor U14992 (N_14992,N_14549,N_14450);
or U14993 (N_14993,N_14569,N_14501);
and U14994 (N_14994,N_14717,N_14678);
nor U14995 (N_14995,N_14618,N_14796);
and U14996 (N_14996,N_14713,N_14543);
nand U14997 (N_14997,N_14577,N_14786);
nand U14998 (N_14998,N_14432,N_14641);
nor U14999 (N_14999,N_14544,N_14720);
nor U15000 (N_15000,N_14697,N_14418);
nor U15001 (N_15001,N_14478,N_14795);
nor U15002 (N_15002,N_14490,N_14777);
and U15003 (N_15003,N_14488,N_14659);
and U15004 (N_15004,N_14450,N_14725);
nand U15005 (N_15005,N_14622,N_14576);
xnor U15006 (N_15006,N_14767,N_14691);
nor U15007 (N_15007,N_14621,N_14477);
nor U15008 (N_15008,N_14647,N_14616);
or U15009 (N_15009,N_14669,N_14647);
and U15010 (N_15010,N_14457,N_14587);
xnor U15011 (N_15011,N_14529,N_14760);
and U15012 (N_15012,N_14561,N_14767);
nor U15013 (N_15013,N_14462,N_14563);
or U15014 (N_15014,N_14486,N_14670);
nand U15015 (N_15015,N_14479,N_14671);
nor U15016 (N_15016,N_14666,N_14431);
or U15017 (N_15017,N_14716,N_14627);
and U15018 (N_15018,N_14410,N_14596);
or U15019 (N_15019,N_14528,N_14431);
nor U15020 (N_15020,N_14745,N_14630);
nand U15021 (N_15021,N_14774,N_14677);
nand U15022 (N_15022,N_14709,N_14572);
or U15023 (N_15023,N_14761,N_14460);
and U15024 (N_15024,N_14613,N_14497);
xnor U15025 (N_15025,N_14490,N_14688);
nand U15026 (N_15026,N_14626,N_14689);
nor U15027 (N_15027,N_14751,N_14535);
nand U15028 (N_15028,N_14430,N_14559);
or U15029 (N_15029,N_14712,N_14726);
or U15030 (N_15030,N_14691,N_14554);
or U15031 (N_15031,N_14755,N_14566);
or U15032 (N_15032,N_14507,N_14501);
nor U15033 (N_15033,N_14664,N_14648);
nand U15034 (N_15034,N_14450,N_14608);
xnor U15035 (N_15035,N_14456,N_14730);
xnor U15036 (N_15036,N_14695,N_14626);
and U15037 (N_15037,N_14543,N_14657);
nor U15038 (N_15038,N_14664,N_14446);
nand U15039 (N_15039,N_14686,N_14790);
nor U15040 (N_15040,N_14510,N_14679);
nor U15041 (N_15041,N_14462,N_14688);
xor U15042 (N_15042,N_14484,N_14634);
nor U15043 (N_15043,N_14784,N_14492);
and U15044 (N_15044,N_14717,N_14536);
xor U15045 (N_15045,N_14500,N_14503);
nor U15046 (N_15046,N_14773,N_14482);
and U15047 (N_15047,N_14619,N_14770);
nor U15048 (N_15048,N_14641,N_14492);
nor U15049 (N_15049,N_14504,N_14500);
and U15050 (N_15050,N_14637,N_14665);
nor U15051 (N_15051,N_14698,N_14498);
nand U15052 (N_15052,N_14609,N_14564);
nand U15053 (N_15053,N_14665,N_14590);
and U15054 (N_15054,N_14571,N_14484);
and U15055 (N_15055,N_14576,N_14468);
and U15056 (N_15056,N_14791,N_14519);
nor U15057 (N_15057,N_14617,N_14510);
and U15058 (N_15058,N_14533,N_14535);
or U15059 (N_15059,N_14469,N_14508);
and U15060 (N_15060,N_14795,N_14671);
and U15061 (N_15061,N_14410,N_14401);
or U15062 (N_15062,N_14672,N_14676);
or U15063 (N_15063,N_14540,N_14667);
nor U15064 (N_15064,N_14607,N_14634);
nand U15065 (N_15065,N_14726,N_14430);
nor U15066 (N_15066,N_14583,N_14750);
or U15067 (N_15067,N_14633,N_14616);
and U15068 (N_15068,N_14739,N_14530);
nand U15069 (N_15069,N_14691,N_14444);
nand U15070 (N_15070,N_14500,N_14606);
nor U15071 (N_15071,N_14729,N_14766);
nor U15072 (N_15072,N_14525,N_14686);
nor U15073 (N_15073,N_14710,N_14754);
and U15074 (N_15074,N_14410,N_14771);
nor U15075 (N_15075,N_14540,N_14788);
nor U15076 (N_15076,N_14496,N_14798);
xor U15077 (N_15077,N_14402,N_14672);
nor U15078 (N_15078,N_14660,N_14482);
xnor U15079 (N_15079,N_14758,N_14581);
nand U15080 (N_15080,N_14443,N_14590);
or U15081 (N_15081,N_14414,N_14629);
nor U15082 (N_15082,N_14649,N_14476);
and U15083 (N_15083,N_14474,N_14713);
nor U15084 (N_15084,N_14669,N_14412);
and U15085 (N_15085,N_14796,N_14603);
nand U15086 (N_15086,N_14546,N_14486);
xor U15087 (N_15087,N_14622,N_14658);
nand U15088 (N_15088,N_14682,N_14741);
and U15089 (N_15089,N_14452,N_14584);
or U15090 (N_15090,N_14563,N_14637);
or U15091 (N_15091,N_14645,N_14679);
nand U15092 (N_15092,N_14539,N_14456);
or U15093 (N_15093,N_14645,N_14638);
xnor U15094 (N_15094,N_14526,N_14705);
nor U15095 (N_15095,N_14742,N_14575);
xnor U15096 (N_15096,N_14484,N_14794);
xnor U15097 (N_15097,N_14624,N_14796);
nor U15098 (N_15098,N_14593,N_14755);
xor U15099 (N_15099,N_14709,N_14553);
nand U15100 (N_15100,N_14604,N_14557);
and U15101 (N_15101,N_14457,N_14477);
or U15102 (N_15102,N_14469,N_14551);
and U15103 (N_15103,N_14514,N_14521);
and U15104 (N_15104,N_14570,N_14512);
nor U15105 (N_15105,N_14743,N_14663);
and U15106 (N_15106,N_14770,N_14718);
and U15107 (N_15107,N_14555,N_14790);
and U15108 (N_15108,N_14714,N_14783);
and U15109 (N_15109,N_14645,N_14676);
or U15110 (N_15110,N_14727,N_14568);
or U15111 (N_15111,N_14534,N_14776);
or U15112 (N_15112,N_14542,N_14445);
or U15113 (N_15113,N_14460,N_14627);
or U15114 (N_15114,N_14479,N_14526);
xor U15115 (N_15115,N_14455,N_14788);
and U15116 (N_15116,N_14409,N_14439);
nand U15117 (N_15117,N_14405,N_14540);
and U15118 (N_15118,N_14497,N_14659);
xnor U15119 (N_15119,N_14589,N_14607);
or U15120 (N_15120,N_14602,N_14460);
nor U15121 (N_15121,N_14429,N_14425);
or U15122 (N_15122,N_14515,N_14539);
nand U15123 (N_15123,N_14726,N_14461);
and U15124 (N_15124,N_14429,N_14515);
or U15125 (N_15125,N_14566,N_14414);
and U15126 (N_15126,N_14574,N_14651);
xor U15127 (N_15127,N_14425,N_14412);
and U15128 (N_15128,N_14696,N_14662);
nand U15129 (N_15129,N_14449,N_14773);
xnor U15130 (N_15130,N_14529,N_14773);
and U15131 (N_15131,N_14478,N_14772);
or U15132 (N_15132,N_14427,N_14731);
or U15133 (N_15133,N_14485,N_14465);
nand U15134 (N_15134,N_14686,N_14786);
and U15135 (N_15135,N_14411,N_14650);
xnor U15136 (N_15136,N_14618,N_14456);
nand U15137 (N_15137,N_14599,N_14648);
or U15138 (N_15138,N_14740,N_14761);
or U15139 (N_15139,N_14650,N_14603);
nand U15140 (N_15140,N_14620,N_14760);
nor U15141 (N_15141,N_14534,N_14596);
or U15142 (N_15142,N_14593,N_14742);
xnor U15143 (N_15143,N_14583,N_14693);
nand U15144 (N_15144,N_14427,N_14734);
nand U15145 (N_15145,N_14707,N_14706);
and U15146 (N_15146,N_14588,N_14473);
or U15147 (N_15147,N_14769,N_14558);
nand U15148 (N_15148,N_14606,N_14523);
nand U15149 (N_15149,N_14641,N_14758);
nand U15150 (N_15150,N_14621,N_14610);
nand U15151 (N_15151,N_14669,N_14782);
nor U15152 (N_15152,N_14447,N_14739);
nor U15153 (N_15153,N_14555,N_14739);
nand U15154 (N_15154,N_14439,N_14579);
and U15155 (N_15155,N_14754,N_14457);
or U15156 (N_15156,N_14483,N_14582);
xnor U15157 (N_15157,N_14787,N_14537);
and U15158 (N_15158,N_14460,N_14568);
xor U15159 (N_15159,N_14636,N_14708);
and U15160 (N_15160,N_14478,N_14734);
nor U15161 (N_15161,N_14464,N_14693);
nor U15162 (N_15162,N_14489,N_14433);
nand U15163 (N_15163,N_14425,N_14641);
xnor U15164 (N_15164,N_14687,N_14547);
xor U15165 (N_15165,N_14520,N_14745);
and U15166 (N_15166,N_14576,N_14440);
xor U15167 (N_15167,N_14753,N_14720);
nand U15168 (N_15168,N_14596,N_14608);
nor U15169 (N_15169,N_14604,N_14539);
nor U15170 (N_15170,N_14564,N_14487);
and U15171 (N_15171,N_14560,N_14405);
xor U15172 (N_15172,N_14767,N_14452);
and U15173 (N_15173,N_14797,N_14418);
and U15174 (N_15174,N_14605,N_14429);
xor U15175 (N_15175,N_14490,N_14619);
or U15176 (N_15176,N_14658,N_14640);
nand U15177 (N_15177,N_14641,N_14698);
xnor U15178 (N_15178,N_14426,N_14631);
xor U15179 (N_15179,N_14567,N_14423);
and U15180 (N_15180,N_14640,N_14458);
and U15181 (N_15181,N_14743,N_14480);
or U15182 (N_15182,N_14505,N_14630);
xnor U15183 (N_15183,N_14598,N_14648);
nor U15184 (N_15184,N_14625,N_14572);
xnor U15185 (N_15185,N_14510,N_14722);
or U15186 (N_15186,N_14630,N_14615);
and U15187 (N_15187,N_14608,N_14656);
nor U15188 (N_15188,N_14620,N_14716);
xnor U15189 (N_15189,N_14506,N_14553);
or U15190 (N_15190,N_14515,N_14427);
and U15191 (N_15191,N_14526,N_14694);
nor U15192 (N_15192,N_14648,N_14406);
and U15193 (N_15193,N_14505,N_14748);
xnor U15194 (N_15194,N_14504,N_14525);
or U15195 (N_15195,N_14545,N_14797);
nand U15196 (N_15196,N_14608,N_14421);
nor U15197 (N_15197,N_14626,N_14684);
nand U15198 (N_15198,N_14786,N_14677);
xor U15199 (N_15199,N_14522,N_14460);
and U15200 (N_15200,N_14917,N_15085);
nor U15201 (N_15201,N_15080,N_14922);
xor U15202 (N_15202,N_14816,N_14851);
nor U15203 (N_15203,N_14959,N_14827);
nand U15204 (N_15204,N_15088,N_14898);
and U15205 (N_15205,N_15052,N_14872);
nor U15206 (N_15206,N_15054,N_15047);
nor U15207 (N_15207,N_15147,N_15187);
or U15208 (N_15208,N_15102,N_14954);
nand U15209 (N_15209,N_15117,N_15049);
xnor U15210 (N_15210,N_14863,N_14808);
and U15211 (N_15211,N_14975,N_14810);
nor U15212 (N_15212,N_15002,N_15060);
xor U15213 (N_15213,N_15029,N_14853);
and U15214 (N_15214,N_15083,N_14821);
and U15215 (N_15215,N_14901,N_14847);
or U15216 (N_15216,N_15086,N_14987);
or U15217 (N_15217,N_15158,N_15172);
nand U15218 (N_15218,N_15070,N_14981);
and U15219 (N_15219,N_15061,N_15048);
and U15220 (N_15220,N_14891,N_14836);
and U15221 (N_15221,N_14871,N_15171);
and U15222 (N_15222,N_14913,N_15067);
nor U15223 (N_15223,N_15149,N_14904);
and U15224 (N_15224,N_14920,N_15125);
nor U15225 (N_15225,N_15160,N_15089);
nand U15226 (N_15226,N_15079,N_14854);
or U15227 (N_15227,N_14865,N_15011);
nor U15228 (N_15228,N_15164,N_15022);
and U15229 (N_15229,N_15134,N_15126);
nor U15230 (N_15230,N_14970,N_14958);
nor U15231 (N_15231,N_15182,N_15152);
or U15232 (N_15232,N_15065,N_14817);
and U15233 (N_15233,N_14979,N_14903);
nor U15234 (N_15234,N_14824,N_15076);
nor U15235 (N_15235,N_15123,N_15021);
or U15236 (N_15236,N_14826,N_15169);
and U15237 (N_15237,N_15075,N_14960);
and U15238 (N_15238,N_14848,N_14866);
xnor U15239 (N_15239,N_14962,N_15000);
nor U15240 (N_15240,N_15057,N_15176);
nand U15241 (N_15241,N_14837,N_15135);
nor U15242 (N_15242,N_15013,N_14804);
xnor U15243 (N_15243,N_15017,N_15096);
nand U15244 (N_15244,N_14961,N_14845);
xnor U15245 (N_15245,N_14870,N_15133);
nor U15246 (N_15246,N_14932,N_14947);
and U15247 (N_15247,N_14820,N_14976);
and U15248 (N_15248,N_15090,N_14807);
nor U15249 (N_15249,N_14839,N_14941);
xor U15250 (N_15250,N_14998,N_14923);
xnor U15251 (N_15251,N_15181,N_15092);
nor U15252 (N_15252,N_15094,N_14800);
and U15253 (N_15253,N_15183,N_14914);
and U15254 (N_15254,N_15168,N_14900);
xnor U15255 (N_15255,N_14929,N_14840);
and U15256 (N_15256,N_14972,N_14936);
and U15257 (N_15257,N_15018,N_15120);
or U15258 (N_15258,N_14966,N_15151);
nand U15259 (N_15259,N_14812,N_14968);
or U15260 (N_15260,N_15110,N_15154);
or U15261 (N_15261,N_15106,N_15156);
nor U15262 (N_15262,N_15107,N_14874);
nor U15263 (N_15263,N_14855,N_14973);
nand U15264 (N_15264,N_15051,N_14942);
nor U15265 (N_15265,N_15167,N_15097);
xor U15266 (N_15266,N_15004,N_14902);
or U15267 (N_15267,N_15100,N_14894);
or U15268 (N_15268,N_15050,N_14869);
xnor U15269 (N_15269,N_14825,N_15024);
nor U15270 (N_15270,N_14938,N_15184);
or U15271 (N_15271,N_14974,N_14802);
nor U15272 (N_15272,N_15109,N_15069);
and U15273 (N_15273,N_14830,N_14993);
xor U15274 (N_15274,N_14828,N_14896);
nand U15275 (N_15275,N_14842,N_14887);
xnor U15276 (N_15276,N_14818,N_15148);
and U15277 (N_15277,N_14911,N_14809);
nand U15278 (N_15278,N_15045,N_15030);
and U15279 (N_15279,N_15119,N_15073);
nor U15280 (N_15280,N_15179,N_15115);
nand U15281 (N_15281,N_15023,N_15032);
nor U15282 (N_15282,N_15019,N_15192);
xnor U15283 (N_15283,N_15136,N_15180);
nand U15284 (N_15284,N_15016,N_15108);
xnor U15285 (N_15285,N_15140,N_15153);
nor U15286 (N_15286,N_15145,N_14864);
nor U15287 (N_15287,N_14886,N_14875);
xor U15288 (N_15288,N_15071,N_15084);
or U15289 (N_15289,N_15101,N_15193);
xor U15290 (N_15290,N_14967,N_15034);
and U15291 (N_15291,N_14969,N_15078);
nand U15292 (N_15292,N_14832,N_15173);
xor U15293 (N_15293,N_14949,N_14850);
or U15294 (N_15294,N_14943,N_14990);
nor U15295 (N_15295,N_15035,N_15129);
nor U15296 (N_15296,N_15178,N_14957);
and U15297 (N_15297,N_15118,N_15068);
xor U15298 (N_15298,N_15170,N_14950);
xor U15299 (N_15299,N_15143,N_14986);
nor U15300 (N_15300,N_14814,N_15053);
xor U15301 (N_15301,N_14956,N_14978);
xnor U15302 (N_15302,N_14838,N_14984);
nand U15303 (N_15303,N_15026,N_14843);
nand U15304 (N_15304,N_14857,N_14926);
xor U15305 (N_15305,N_15194,N_14835);
or U15306 (N_15306,N_15038,N_14822);
xnor U15307 (N_15307,N_14861,N_15103);
or U15308 (N_15308,N_15175,N_14852);
or U15309 (N_15309,N_15020,N_15037);
nor U15310 (N_15310,N_14803,N_14940);
nor U15311 (N_15311,N_15091,N_15114);
or U15312 (N_15312,N_14805,N_15138);
xor U15313 (N_15313,N_14884,N_15044);
nand U15314 (N_15314,N_15198,N_14908);
xor U15315 (N_15315,N_14819,N_14948);
nor U15316 (N_15316,N_15093,N_14895);
and U15317 (N_15317,N_14888,N_14955);
nor U15318 (N_15318,N_15095,N_14909);
xor U15319 (N_15319,N_14897,N_14893);
xnor U15320 (N_15320,N_15064,N_14879);
nor U15321 (N_15321,N_15112,N_15042);
nand U15322 (N_15322,N_14833,N_15121);
xnor U15323 (N_15323,N_15185,N_15196);
nor U15324 (N_15324,N_14907,N_14905);
or U15325 (N_15325,N_14930,N_15144);
nand U15326 (N_15326,N_14935,N_15014);
xor U15327 (N_15327,N_15190,N_14931);
nand U15328 (N_15328,N_14933,N_15197);
nand U15329 (N_15329,N_14877,N_15141);
xnor U15330 (N_15330,N_15074,N_15028);
xor U15331 (N_15331,N_14939,N_15174);
or U15332 (N_15332,N_15003,N_15157);
nand U15333 (N_15333,N_14921,N_14867);
or U15334 (N_15334,N_15191,N_14995);
xnor U15335 (N_15335,N_14937,N_14996);
xnor U15336 (N_15336,N_14878,N_15188);
nand U15337 (N_15337,N_14983,N_14859);
nand U15338 (N_15338,N_15039,N_15056);
and U15339 (N_15339,N_15146,N_15033);
xnor U15340 (N_15340,N_14811,N_15010);
and U15341 (N_15341,N_14841,N_15124);
nor U15342 (N_15342,N_14882,N_14846);
nand U15343 (N_15343,N_14934,N_14889);
and U15344 (N_15344,N_15177,N_14952);
nand U15345 (N_15345,N_14801,N_14806);
xor U15346 (N_15346,N_14999,N_14989);
nor U15347 (N_15347,N_15186,N_15062);
and U15348 (N_15348,N_15155,N_14858);
nand U15349 (N_15349,N_14951,N_15162);
nor U15350 (N_15350,N_14997,N_14965);
or U15351 (N_15351,N_14985,N_14919);
nand U15352 (N_15352,N_14971,N_14924);
xnor U15353 (N_15353,N_15015,N_15199);
nand U15354 (N_15354,N_15063,N_14868);
nand U15355 (N_15355,N_14944,N_15066);
nand U15356 (N_15356,N_14906,N_14890);
nand U15357 (N_15357,N_15006,N_14925);
nand U15358 (N_15358,N_14946,N_14823);
nand U15359 (N_15359,N_14964,N_15009);
and U15360 (N_15360,N_15036,N_15165);
xor U15361 (N_15361,N_15132,N_15001);
nand U15362 (N_15362,N_14953,N_15113);
and U15363 (N_15363,N_15087,N_14988);
xor U15364 (N_15364,N_15128,N_14918);
and U15365 (N_15365,N_15127,N_14856);
and U15366 (N_15366,N_14831,N_14982);
nor U15367 (N_15367,N_15025,N_15031);
and U15368 (N_15368,N_14991,N_15159);
or U15369 (N_15369,N_14860,N_15161);
and U15370 (N_15370,N_14916,N_14899);
or U15371 (N_15371,N_15055,N_15142);
or U15372 (N_15372,N_14873,N_15098);
nand U15373 (N_15373,N_15059,N_14862);
nand U15374 (N_15374,N_15008,N_15137);
nand U15375 (N_15375,N_15105,N_15027);
nand U15376 (N_15376,N_15111,N_14813);
nor U15377 (N_15377,N_15139,N_15130);
xnor U15378 (N_15378,N_15005,N_14915);
or U15379 (N_15379,N_15099,N_15043);
nand U15380 (N_15380,N_15116,N_15150);
and U15381 (N_15381,N_15166,N_15163);
xor U15382 (N_15382,N_15007,N_14881);
and U15383 (N_15383,N_14945,N_14849);
xor U15384 (N_15384,N_14992,N_14892);
nor U15385 (N_15385,N_14928,N_15077);
nor U15386 (N_15386,N_15040,N_15041);
xor U15387 (N_15387,N_14980,N_14963);
xor U15388 (N_15388,N_15046,N_14912);
xor U15389 (N_15389,N_14927,N_14910);
nor U15390 (N_15390,N_14994,N_15082);
xor U15391 (N_15391,N_15081,N_14883);
nor U15392 (N_15392,N_15012,N_15104);
nand U15393 (N_15393,N_15189,N_14876);
or U15394 (N_15394,N_14885,N_14880);
and U15395 (N_15395,N_15122,N_14815);
or U15396 (N_15396,N_15058,N_14844);
xor U15397 (N_15397,N_15131,N_15195);
nor U15398 (N_15398,N_14834,N_14829);
xor U15399 (N_15399,N_15072,N_14977);
and U15400 (N_15400,N_15076,N_15121);
or U15401 (N_15401,N_15049,N_14890);
xnor U15402 (N_15402,N_14964,N_15173);
and U15403 (N_15403,N_14910,N_14885);
or U15404 (N_15404,N_15056,N_14903);
nor U15405 (N_15405,N_14998,N_14861);
or U15406 (N_15406,N_14951,N_15121);
xor U15407 (N_15407,N_15186,N_15126);
and U15408 (N_15408,N_15098,N_14856);
and U15409 (N_15409,N_14806,N_15013);
xnor U15410 (N_15410,N_14936,N_15161);
nor U15411 (N_15411,N_14813,N_15052);
or U15412 (N_15412,N_14902,N_15107);
and U15413 (N_15413,N_14808,N_15162);
nor U15414 (N_15414,N_14923,N_15031);
xnor U15415 (N_15415,N_14956,N_14983);
and U15416 (N_15416,N_15180,N_14940);
xnor U15417 (N_15417,N_14938,N_14886);
and U15418 (N_15418,N_15146,N_14874);
nor U15419 (N_15419,N_15049,N_15170);
nor U15420 (N_15420,N_15131,N_14868);
or U15421 (N_15421,N_15002,N_14985);
and U15422 (N_15422,N_14932,N_15083);
or U15423 (N_15423,N_15188,N_14904);
nor U15424 (N_15424,N_14815,N_14943);
xnor U15425 (N_15425,N_14860,N_15145);
nand U15426 (N_15426,N_15007,N_14914);
or U15427 (N_15427,N_15162,N_14831);
xnor U15428 (N_15428,N_15047,N_14957);
or U15429 (N_15429,N_15188,N_15157);
nand U15430 (N_15430,N_14891,N_14972);
xnor U15431 (N_15431,N_15120,N_15144);
xor U15432 (N_15432,N_15076,N_15190);
nand U15433 (N_15433,N_15032,N_14805);
or U15434 (N_15434,N_14850,N_15158);
nor U15435 (N_15435,N_15098,N_14842);
or U15436 (N_15436,N_14974,N_15166);
and U15437 (N_15437,N_15020,N_15092);
nor U15438 (N_15438,N_14954,N_14914);
nor U15439 (N_15439,N_14887,N_14899);
or U15440 (N_15440,N_15078,N_14981);
and U15441 (N_15441,N_14993,N_15055);
and U15442 (N_15442,N_15125,N_14914);
xor U15443 (N_15443,N_15171,N_15174);
nand U15444 (N_15444,N_14952,N_14903);
and U15445 (N_15445,N_15089,N_15142);
nand U15446 (N_15446,N_14941,N_14887);
nand U15447 (N_15447,N_14968,N_14814);
or U15448 (N_15448,N_15065,N_14865);
and U15449 (N_15449,N_15091,N_14818);
or U15450 (N_15450,N_14823,N_15092);
and U15451 (N_15451,N_14903,N_15144);
xnor U15452 (N_15452,N_14956,N_14969);
nor U15453 (N_15453,N_14842,N_15126);
nand U15454 (N_15454,N_14829,N_14806);
and U15455 (N_15455,N_14828,N_15133);
xor U15456 (N_15456,N_14829,N_15057);
nor U15457 (N_15457,N_15073,N_14819);
nor U15458 (N_15458,N_15132,N_15041);
nor U15459 (N_15459,N_14964,N_15146);
nand U15460 (N_15460,N_15189,N_15157);
or U15461 (N_15461,N_15156,N_14950);
or U15462 (N_15462,N_15145,N_14849);
and U15463 (N_15463,N_15143,N_14890);
nand U15464 (N_15464,N_14804,N_15134);
nor U15465 (N_15465,N_14842,N_14920);
and U15466 (N_15466,N_14876,N_14943);
nor U15467 (N_15467,N_15017,N_14965);
and U15468 (N_15468,N_14949,N_15054);
nand U15469 (N_15469,N_14860,N_14802);
nor U15470 (N_15470,N_14867,N_14997);
or U15471 (N_15471,N_14971,N_14816);
nand U15472 (N_15472,N_15195,N_14904);
nor U15473 (N_15473,N_15175,N_14891);
and U15474 (N_15474,N_15068,N_15164);
and U15475 (N_15475,N_14886,N_14990);
nor U15476 (N_15476,N_14811,N_14814);
and U15477 (N_15477,N_14858,N_15158);
and U15478 (N_15478,N_14858,N_14853);
nor U15479 (N_15479,N_14853,N_15118);
nand U15480 (N_15480,N_14800,N_14971);
nand U15481 (N_15481,N_14980,N_15094);
or U15482 (N_15482,N_14853,N_15047);
or U15483 (N_15483,N_14806,N_15170);
xor U15484 (N_15484,N_15065,N_14892);
or U15485 (N_15485,N_15016,N_15032);
xor U15486 (N_15486,N_14844,N_14845);
nor U15487 (N_15487,N_15101,N_15003);
or U15488 (N_15488,N_15018,N_15037);
xnor U15489 (N_15489,N_15167,N_14879);
xnor U15490 (N_15490,N_14848,N_15024);
nand U15491 (N_15491,N_14805,N_15134);
nand U15492 (N_15492,N_14993,N_15182);
and U15493 (N_15493,N_14834,N_14988);
or U15494 (N_15494,N_15172,N_15161);
and U15495 (N_15495,N_15027,N_14906);
or U15496 (N_15496,N_14818,N_14959);
and U15497 (N_15497,N_15008,N_14967);
nor U15498 (N_15498,N_14913,N_15089);
nand U15499 (N_15499,N_14849,N_14809);
and U15500 (N_15500,N_15162,N_15124);
nor U15501 (N_15501,N_15149,N_14974);
xnor U15502 (N_15502,N_14976,N_14997);
nor U15503 (N_15503,N_15191,N_14825);
xnor U15504 (N_15504,N_14909,N_15107);
xnor U15505 (N_15505,N_14844,N_15005);
xnor U15506 (N_15506,N_15193,N_14934);
xor U15507 (N_15507,N_15167,N_14892);
xnor U15508 (N_15508,N_15005,N_15177);
nor U15509 (N_15509,N_15151,N_15187);
or U15510 (N_15510,N_14921,N_15013);
or U15511 (N_15511,N_15159,N_15133);
and U15512 (N_15512,N_14855,N_14817);
nand U15513 (N_15513,N_15060,N_15068);
and U15514 (N_15514,N_14899,N_15005);
xnor U15515 (N_15515,N_14903,N_15143);
xnor U15516 (N_15516,N_15120,N_15177);
or U15517 (N_15517,N_15158,N_15046);
or U15518 (N_15518,N_15048,N_15157);
or U15519 (N_15519,N_14934,N_14920);
and U15520 (N_15520,N_15072,N_15062);
nor U15521 (N_15521,N_15003,N_14809);
nor U15522 (N_15522,N_15083,N_15120);
xor U15523 (N_15523,N_15084,N_15067);
xor U15524 (N_15524,N_15121,N_15118);
or U15525 (N_15525,N_14865,N_15093);
nor U15526 (N_15526,N_14891,N_15026);
xor U15527 (N_15527,N_15037,N_14889);
nor U15528 (N_15528,N_15192,N_14991);
nand U15529 (N_15529,N_14874,N_15007);
and U15530 (N_15530,N_15045,N_14910);
and U15531 (N_15531,N_15148,N_15138);
or U15532 (N_15532,N_14853,N_14957);
xor U15533 (N_15533,N_15193,N_15059);
and U15534 (N_15534,N_14871,N_14825);
and U15535 (N_15535,N_14982,N_14925);
nor U15536 (N_15536,N_15016,N_14997);
xor U15537 (N_15537,N_15125,N_15009);
nand U15538 (N_15538,N_15151,N_14936);
nor U15539 (N_15539,N_14910,N_15182);
and U15540 (N_15540,N_15149,N_14986);
nand U15541 (N_15541,N_14853,N_14993);
or U15542 (N_15542,N_15036,N_15005);
nand U15543 (N_15543,N_14871,N_15177);
nand U15544 (N_15544,N_15182,N_15062);
nor U15545 (N_15545,N_15172,N_14967);
nand U15546 (N_15546,N_14915,N_15020);
xor U15547 (N_15547,N_14999,N_14892);
nand U15548 (N_15548,N_15064,N_15088);
xor U15549 (N_15549,N_14971,N_14950);
xnor U15550 (N_15550,N_15086,N_14883);
nor U15551 (N_15551,N_15001,N_15008);
nand U15552 (N_15552,N_14966,N_15163);
nand U15553 (N_15553,N_15142,N_15014);
xnor U15554 (N_15554,N_15077,N_15058);
or U15555 (N_15555,N_15057,N_15038);
or U15556 (N_15556,N_15032,N_14950);
or U15557 (N_15557,N_14807,N_15062);
nor U15558 (N_15558,N_15003,N_14984);
nand U15559 (N_15559,N_14954,N_14881);
and U15560 (N_15560,N_15023,N_15198);
xnor U15561 (N_15561,N_15102,N_15140);
or U15562 (N_15562,N_14980,N_14886);
and U15563 (N_15563,N_15113,N_14870);
or U15564 (N_15564,N_15097,N_15119);
xnor U15565 (N_15565,N_15124,N_14894);
xor U15566 (N_15566,N_14898,N_14820);
xnor U15567 (N_15567,N_15183,N_14823);
and U15568 (N_15568,N_14916,N_14869);
xnor U15569 (N_15569,N_15033,N_15002);
and U15570 (N_15570,N_15021,N_14966);
nand U15571 (N_15571,N_15129,N_14930);
and U15572 (N_15572,N_15139,N_14994);
nand U15573 (N_15573,N_15195,N_15176);
nand U15574 (N_15574,N_15002,N_14939);
nand U15575 (N_15575,N_14860,N_14836);
xnor U15576 (N_15576,N_14865,N_15120);
or U15577 (N_15577,N_14944,N_15046);
nand U15578 (N_15578,N_15129,N_14939);
nor U15579 (N_15579,N_14942,N_14986);
nand U15580 (N_15580,N_14869,N_14816);
nand U15581 (N_15581,N_15189,N_14954);
nand U15582 (N_15582,N_15092,N_14869);
nand U15583 (N_15583,N_14833,N_14825);
and U15584 (N_15584,N_14830,N_14846);
nand U15585 (N_15585,N_15149,N_15005);
nor U15586 (N_15586,N_14857,N_15087);
xor U15587 (N_15587,N_15186,N_15022);
and U15588 (N_15588,N_14908,N_14891);
and U15589 (N_15589,N_15031,N_15133);
or U15590 (N_15590,N_14886,N_15159);
and U15591 (N_15591,N_15153,N_15054);
or U15592 (N_15592,N_14859,N_15040);
nand U15593 (N_15593,N_15007,N_15073);
and U15594 (N_15594,N_14988,N_14889);
nand U15595 (N_15595,N_15007,N_15189);
and U15596 (N_15596,N_15198,N_14943);
or U15597 (N_15597,N_14965,N_14847);
xnor U15598 (N_15598,N_15060,N_15176);
and U15599 (N_15599,N_14805,N_15097);
or U15600 (N_15600,N_15405,N_15377);
xor U15601 (N_15601,N_15489,N_15424);
or U15602 (N_15602,N_15378,N_15292);
xnor U15603 (N_15603,N_15535,N_15294);
xor U15604 (N_15604,N_15420,N_15313);
or U15605 (N_15605,N_15317,N_15464);
nand U15606 (N_15606,N_15568,N_15500);
nor U15607 (N_15607,N_15279,N_15347);
or U15608 (N_15608,N_15573,N_15213);
or U15609 (N_15609,N_15280,N_15579);
and U15610 (N_15610,N_15277,N_15283);
nand U15611 (N_15611,N_15487,N_15570);
and U15612 (N_15612,N_15444,N_15381);
or U15613 (N_15613,N_15565,N_15215);
xnor U15614 (N_15614,N_15597,N_15338);
and U15615 (N_15615,N_15567,N_15574);
nor U15616 (N_15616,N_15484,N_15514);
and U15617 (N_15617,N_15512,N_15376);
or U15618 (N_15618,N_15441,N_15527);
and U15619 (N_15619,N_15486,N_15380);
and U15620 (N_15620,N_15284,N_15558);
or U15621 (N_15621,N_15418,N_15416);
xor U15622 (N_15622,N_15547,N_15504);
or U15623 (N_15623,N_15218,N_15415);
nand U15624 (N_15624,N_15373,N_15581);
nor U15625 (N_15625,N_15458,N_15289);
xor U15626 (N_15626,N_15261,N_15511);
nand U15627 (N_15627,N_15226,N_15485);
xor U15628 (N_15628,N_15201,N_15503);
nor U15629 (N_15629,N_15519,N_15236);
nand U15630 (N_15630,N_15440,N_15245);
and U15631 (N_15631,N_15260,N_15293);
nand U15632 (N_15632,N_15372,N_15240);
nor U15633 (N_15633,N_15276,N_15454);
xor U15634 (N_15634,N_15355,N_15305);
xor U15635 (N_15635,N_15216,N_15554);
xor U15636 (N_15636,N_15219,N_15266);
nand U15637 (N_15637,N_15346,N_15259);
and U15638 (N_15638,N_15571,N_15231);
and U15639 (N_15639,N_15361,N_15368);
and U15640 (N_15640,N_15587,N_15457);
nor U15641 (N_15641,N_15479,N_15359);
xor U15642 (N_15642,N_15350,N_15434);
nand U15643 (N_15643,N_15401,N_15330);
nand U15644 (N_15644,N_15497,N_15447);
and U15645 (N_15645,N_15495,N_15501);
nor U15646 (N_15646,N_15370,N_15446);
nor U15647 (N_15647,N_15431,N_15311);
xnor U15648 (N_15648,N_15507,N_15445);
nor U15649 (N_15649,N_15423,N_15584);
nand U15650 (N_15650,N_15212,N_15349);
xnor U15651 (N_15651,N_15598,N_15302);
nand U15652 (N_15652,N_15451,N_15220);
or U15653 (N_15653,N_15273,N_15256);
xnor U15654 (N_15654,N_15417,N_15477);
and U15655 (N_15655,N_15426,N_15510);
and U15656 (N_15656,N_15335,N_15551);
or U15657 (N_15657,N_15360,N_15327);
nor U15658 (N_15658,N_15304,N_15433);
xnor U15659 (N_15659,N_15421,N_15287);
and U15660 (N_15660,N_15351,N_15463);
or U15661 (N_15661,N_15333,N_15233);
or U15662 (N_15662,N_15369,N_15400);
nand U15663 (N_15663,N_15515,N_15436);
or U15664 (N_15664,N_15412,N_15337);
xor U15665 (N_15665,N_15270,N_15462);
or U15666 (N_15666,N_15599,N_15564);
or U15667 (N_15667,N_15448,N_15460);
nand U15668 (N_15668,N_15248,N_15344);
or U15669 (N_15669,N_15468,N_15288);
nor U15670 (N_15670,N_15403,N_15592);
xnor U15671 (N_15671,N_15528,N_15529);
or U15672 (N_15672,N_15353,N_15221);
or U15673 (N_15673,N_15275,N_15472);
nand U15674 (N_15674,N_15365,N_15588);
xor U15675 (N_15675,N_15395,N_15589);
or U15676 (N_15676,N_15237,N_15427);
nor U15677 (N_15677,N_15550,N_15322);
xor U15678 (N_15678,N_15591,N_15538);
or U15679 (N_15679,N_15202,N_15223);
and U15680 (N_15680,N_15580,N_15315);
and U15681 (N_15681,N_15517,N_15384);
and U15682 (N_15682,N_15291,N_15482);
or U15683 (N_15683,N_15374,N_15402);
nor U15684 (N_15684,N_15257,N_15522);
and U15685 (N_15685,N_15227,N_15228);
or U15686 (N_15686,N_15300,N_15306);
and U15687 (N_15687,N_15453,N_15467);
and U15688 (N_15688,N_15540,N_15536);
nand U15689 (N_15689,N_15366,N_15407);
nand U15690 (N_15690,N_15391,N_15326);
and U15691 (N_15691,N_15543,N_15548);
and U15692 (N_15692,N_15576,N_15207);
or U15693 (N_15693,N_15471,N_15362);
and U15694 (N_15694,N_15569,N_15585);
xnor U15695 (N_15695,N_15537,N_15388);
nand U15696 (N_15696,N_15475,N_15235);
or U15697 (N_15697,N_15480,N_15438);
or U15698 (N_15698,N_15532,N_15252);
xnor U15699 (N_15699,N_15549,N_15367);
nand U15700 (N_15700,N_15269,N_15559);
and U15701 (N_15701,N_15524,N_15296);
or U15702 (N_15702,N_15465,N_15325);
nand U15703 (N_15703,N_15483,N_15394);
and U15704 (N_15704,N_15340,N_15319);
nor U15705 (N_15705,N_15469,N_15490);
or U15706 (N_15706,N_15267,N_15443);
or U15707 (N_15707,N_15309,N_15345);
nand U15708 (N_15708,N_15336,N_15506);
nand U15709 (N_15709,N_15307,N_15274);
and U15710 (N_15710,N_15520,N_15525);
xnor U15711 (N_15711,N_15290,N_15281);
and U15712 (N_15712,N_15531,N_15238);
nor U15713 (N_15713,N_15390,N_15250);
xor U15714 (N_15714,N_15314,N_15398);
or U15715 (N_15715,N_15208,N_15234);
nor U15716 (N_15716,N_15502,N_15328);
xor U15717 (N_15717,N_15232,N_15386);
nor U15718 (N_15718,N_15357,N_15393);
nand U15719 (N_15719,N_15432,N_15348);
and U15720 (N_15720,N_15324,N_15387);
nor U15721 (N_15721,N_15541,N_15254);
and U15722 (N_15722,N_15255,N_15299);
nor U15723 (N_15723,N_15200,N_15382);
or U15724 (N_15724,N_15316,N_15264);
nor U15725 (N_15725,N_15542,N_15523);
nor U15726 (N_15726,N_15561,N_15498);
and U15727 (N_15727,N_15509,N_15556);
nor U15728 (N_15728,N_15329,N_15363);
or U15729 (N_15729,N_15318,N_15310);
or U15730 (N_15730,N_15578,N_15545);
or U15731 (N_15731,N_15225,N_15411);
xnor U15732 (N_15732,N_15452,N_15566);
nand U15733 (N_15733,N_15358,N_15271);
nand U15734 (N_15734,N_15364,N_15332);
or U15735 (N_15735,N_15526,N_15456);
and U15736 (N_15736,N_15513,N_15303);
nor U15737 (N_15737,N_15244,N_15214);
and U15738 (N_15738,N_15383,N_15222);
and U15739 (N_15739,N_15435,N_15505);
nor U15740 (N_15740,N_15552,N_15521);
nand U15741 (N_15741,N_15466,N_15494);
nand U15742 (N_15742,N_15210,N_15389);
and U15743 (N_15743,N_15473,N_15243);
xnor U15744 (N_15744,N_15575,N_15408);
nand U15745 (N_15745,N_15413,N_15242);
or U15746 (N_15746,N_15204,N_15251);
or U15747 (N_15747,N_15459,N_15499);
or U15748 (N_15748,N_15409,N_15553);
or U15749 (N_15749,N_15491,N_15428);
nand U15750 (N_15750,N_15206,N_15385);
nor U15751 (N_15751,N_15334,N_15392);
or U15752 (N_15752,N_15582,N_15481);
and U15753 (N_15753,N_15422,N_15331);
nor U15754 (N_15754,N_15211,N_15341);
and U15755 (N_15755,N_15375,N_15590);
or U15756 (N_15756,N_15285,N_15419);
xor U15757 (N_15757,N_15474,N_15282);
and U15758 (N_15758,N_15450,N_15354);
or U15759 (N_15759,N_15308,N_15298);
or U15760 (N_15760,N_15476,N_15301);
nand U15761 (N_15761,N_15246,N_15268);
or U15762 (N_15762,N_15449,N_15356);
xor U15763 (N_15763,N_15249,N_15278);
nor U15764 (N_15764,N_15247,N_15461);
and U15765 (N_15765,N_15496,N_15312);
nand U15766 (N_15766,N_15262,N_15533);
xnor U15767 (N_15767,N_15203,N_15410);
xnor U15768 (N_15768,N_15230,N_15492);
xor U15769 (N_15769,N_15263,N_15253);
or U15770 (N_15770,N_15518,N_15544);
and U15771 (N_15771,N_15286,N_15572);
nand U15772 (N_15772,N_15379,N_15258);
nand U15773 (N_15773,N_15586,N_15209);
nor U15774 (N_15774,N_15439,N_15594);
nor U15775 (N_15775,N_15470,N_15371);
xor U15776 (N_15776,N_15399,N_15339);
or U15777 (N_15777,N_15562,N_15404);
and U15778 (N_15778,N_15297,N_15425);
xor U15779 (N_15779,N_15352,N_15321);
or U15780 (N_15780,N_15534,N_15530);
and U15781 (N_15781,N_15595,N_15320);
xor U15782 (N_15782,N_15323,N_15343);
and U15783 (N_15783,N_15539,N_15241);
nand U15784 (N_15784,N_15593,N_15437);
and U15785 (N_15785,N_15205,N_15406);
and U15786 (N_15786,N_15396,N_15596);
and U15787 (N_15787,N_15397,N_15442);
nand U15788 (N_15788,N_15508,N_15493);
nand U15789 (N_15789,N_15229,N_15546);
or U15790 (N_15790,N_15295,N_15429);
and U15791 (N_15791,N_15488,N_15342);
and U15792 (N_15792,N_15455,N_15555);
xor U15793 (N_15793,N_15516,N_15557);
and U15794 (N_15794,N_15239,N_15265);
nor U15795 (N_15795,N_15430,N_15563);
xor U15796 (N_15796,N_15478,N_15583);
nor U15797 (N_15797,N_15577,N_15224);
nand U15798 (N_15798,N_15414,N_15272);
or U15799 (N_15799,N_15217,N_15560);
xnor U15800 (N_15800,N_15244,N_15540);
nor U15801 (N_15801,N_15337,N_15571);
nor U15802 (N_15802,N_15271,N_15269);
and U15803 (N_15803,N_15570,N_15426);
xor U15804 (N_15804,N_15463,N_15348);
xnor U15805 (N_15805,N_15543,N_15210);
nor U15806 (N_15806,N_15321,N_15375);
nand U15807 (N_15807,N_15347,N_15341);
and U15808 (N_15808,N_15470,N_15315);
and U15809 (N_15809,N_15571,N_15424);
or U15810 (N_15810,N_15480,N_15338);
xor U15811 (N_15811,N_15530,N_15206);
nor U15812 (N_15812,N_15485,N_15471);
nor U15813 (N_15813,N_15465,N_15539);
or U15814 (N_15814,N_15342,N_15585);
or U15815 (N_15815,N_15445,N_15515);
xor U15816 (N_15816,N_15263,N_15379);
nor U15817 (N_15817,N_15380,N_15566);
xnor U15818 (N_15818,N_15408,N_15250);
nand U15819 (N_15819,N_15394,N_15298);
or U15820 (N_15820,N_15584,N_15449);
and U15821 (N_15821,N_15531,N_15390);
nor U15822 (N_15822,N_15424,N_15578);
or U15823 (N_15823,N_15326,N_15222);
nor U15824 (N_15824,N_15484,N_15367);
and U15825 (N_15825,N_15295,N_15547);
xnor U15826 (N_15826,N_15340,N_15435);
or U15827 (N_15827,N_15217,N_15563);
or U15828 (N_15828,N_15351,N_15459);
xor U15829 (N_15829,N_15323,N_15473);
nor U15830 (N_15830,N_15205,N_15329);
nand U15831 (N_15831,N_15539,N_15327);
xnor U15832 (N_15832,N_15231,N_15282);
nor U15833 (N_15833,N_15594,N_15472);
and U15834 (N_15834,N_15216,N_15341);
nand U15835 (N_15835,N_15406,N_15328);
nand U15836 (N_15836,N_15493,N_15495);
nor U15837 (N_15837,N_15338,N_15364);
nor U15838 (N_15838,N_15326,N_15236);
or U15839 (N_15839,N_15334,N_15225);
nand U15840 (N_15840,N_15201,N_15483);
and U15841 (N_15841,N_15330,N_15568);
and U15842 (N_15842,N_15342,N_15493);
and U15843 (N_15843,N_15471,N_15543);
nor U15844 (N_15844,N_15573,N_15261);
xnor U15845 (N_15845,N_15502,N_15479);
or U15846 (N_15846,N_15560,N_15272);
xor U15847 (N_15847,N_15443,N_15588);
and U15848 (N_15848,N_15504,N_15325);
nor U15849 (N_15849,N_15214,N_15341);
or U15850 (N_15850,N_15206,N_15456);
and U15851 (N_15851,N_15540,N_15265);
xor U15852 (N_15852,N_15325,N_15573);
xnor U15853 (N_15853,N_15342,N_15247);
and U15854 (N_15854,N_15312,N_15479);
nand U15855 (N_15855,N_15241,N_15218);
nand U15856 (N_15856,N_15471,N_15520);
nand U15857 (N_15857,N_15400,N_15414);
nor U15858 (N_15858,N_15552,N_15274);
nor U15859 (N_15859,N_15572,N_15421);
and U15860 (N_15860,N_15344,N_15431);
nand U15861 (N_15861,N_15456,N_15538);
or U15862 (N_15862,N_15511,N_15361);
and U15863 (N_15863,N_15273,N_15269);
nand U15864 (N_15864,N_15209,N_15208);
nor U15865 (N_15865,N_15471,N_15536);
nor U15866 (N_15866,N_15234,N_15464);
nand U15867 (N_15867,N_15231,N_15484);
xor U15868 (N_15868,N_15372,N_15491);
and U15869 (N_15869,N_15239,N_15508);
nand U15870 (N_15870,N_15487,N_15339);
xor U15871 (N_15871,N_15425,N_15427);
nand U15872 (N_15872,N_15587,N_15522);
nor U15873 (N_15873,N_15426,N_15235);
xor U15874 (N_15874,N_15582,N_15313);
nand U15875 (N_15875,N_15486,N_15278);
xor U15876 (N_15876,N_15483,N_15282);
or U15877 (N_15877,N_15586,N_15462);
nor U15878 (N_15878,N_15454,N_15556);
xnor U15879 (N_15879,N_15310,N_15456);
xor U15880 (N_15880,N_15355,N_15530);
or U15881 (N_15881,N_15401,N_15475);
xor U15882 (N_15882,N_15238,N_15565);
nor U15883 (N_15883,N_15547,N_15452);
nand U15884 (N_15884,N_15506,N_15411);
nor U15885 (N_15885,N_15309,N_15266);
and U15886 (N_15886,N_15392,N_15416);
xor U15887 (N_15887,N_15414,N_15474);
nor U15888 (N_15888,N_15534,N_15207);
nand U15889 (N_15889,N_15400,N_15280);
nand U15890 (N_15890,N_15595,N_15324);
nor U15891 (N_15891,N_15504,N_15259);
nand U15892 (N_15892,N_15467,N_15478);
nand U15893 (N_15893,N_15376,N_15214);
xor U15894 (N_15894,N_15422,N_15224);
or U15895 (N_15895,N_15512,N_15304);
xor U15896 (N_15896,N_15476,N_15460);
or U15897 (N_15897,N_15222,N_15536);
nor U15898 (N_15898,N_15291,N_15406);
nand U15899 (N_15899,N_15422,N_15440);
and U15900 (N_15900,N_15298,N_15260);
or U15901 (N_15901,N_15415,N_15493);
nand U15902 (N_15902,N_15250,N_15493);
and U15903 (N_15903,N_15432,N_15550);
xnor U15904 (N_15904,N_15210,N_15492);
or U15905 (N_15905,N_15546,N_15377);
nor U15906 (N_15906,N_15470,N_15414);
or U15907 (N_15907,N_15513,N_15202);
and U15908 (N_15908,N_15334,N_15391);
nor U15909 (N_15909,N_15451,N_15484);
xor U15910 (N_15910,N_15403,N_15320);
nand U15911 (N_15911,N_15389,N_15203);
nand U15912 (N_15912,N_15257,N_15220);
or U15913 (N_15913,N_15258,N_15540);
or U15914 (N_15914,N_15244,N_15423);
nor U15915 (N_15915,N_15421,N_15223);
or U15916 (N_15916,N_15408,N_15500);
nor U15917 (N_15917,N_15311,N_15404);
and U15918 (N_15918,N_15400,N_15223);
nand U15919 (N_15919,N_15379,N_15281);
or U15920 (N_15920,N_15245,N_15531);
nand U15921 (N_15921,N_15378,N_15287);
or U15922 (N_15922,N_15581,N_15528);
or U15923 (N_15923,N_15458,N_15269);
or U15924 (N_15924,N_15348,N_15305);
nor U15925 (N_15925,N_15292,N_15592);
xor U15926 (N_15926,N_15278,N_15415);
nand U15927 (N_15927,N_15399,N_15303);
xor U15928 (N_15928,N_15281,N_15250);
and U15929 (N_15929,N_15459,N_15415);
xnor U15930 (N_15930,N_15441,N_15451);
or U15931 (N_15931,N_15332,N_15428);
nor U15932 (N_15932,N_15331,N_15347);
and U15933 (N_15933,N_15204,N_15425);
nor U15934 (N_15934,N_15314,N_15239);
nand U15935 (N_15935,N_15352,N_15413);
nand U15936 (N_15936,N_15523,N_15279);
nor U15937 (N_15937,N_15344,N_15594);
and U15938 (N_15938,N_15415,N_15353);
nor U15939 (N_15939,N_15552,N_15303);
or U15940 (N_15940,N_15287,N_15571);
and U15941 (N_15941,N_15440,N_15351);
nand U15942 (N_15942,N_15371,N_15341);
or U15943 (N_15943,N_15293,N_15431);
or U15944 (N_15944,N_15218,N_15401);
nor U15945 (N_15945,N_15202,N_15544);
nand U15946 (N_15946,N_15427,N_15509);
or U15947 (N_15947,N_15385,N_15359);
xor U15948 (N_15948,N_15446,N_15578);
and U15949 (N_15949,N_15577,N_15435);
xor U15950 (N_15950,N_15479,N_15410);
or U15951 (N_15951,N_15303,N_15498);
nand U15952 (N_15952,N_15539,N_15412);
nor U15953 (N_15953,N_15391,N_15593);
nor U15954 (N_15954,N_15293,N_15415);
nor U15955 (N_15955,N_15280,N_15318);
nor U15956 (N_15956,N_15485,N_15396);
nor U15957 (N_15957,N_15383,N_15323);
xnor U15958 (N_15958,N_15252,N_15290);
nand U15959 (N_15959,N_15215,N_15572);
xor U15960 (N_15960,N_15451,N_15529);
and U15961 (N_15961,N_15526,N_15390);
xor U15962 (N_15962,N_15226,N_15569);
and U15963 (N_15963,N_15247,N_15331);
nor U15964 (N_15964,N_15453,N_15278);
nor U15965 (N_15965,N_15404,N_15287);
nor U15966 (N_15966,N_15348,N_15354);
xor U15967 (N_15967,N_15213,N_15347);
xor U15968 (N_15968,N_15553,N_15212);
and U15969 (N_15969,N_15247,N_15401);
nand U15970 (N_15970,N_15299,N_15261);
nand U15971 (N_15971,N_15438,N_15219);
and U15972 (N_15972,N_15281,N_15261);
nand U15973 (N_15973,N_15332,N_15217);
or U15974 (N_15974,N_15533,N_15545);
nor U15975 (N_15975,N_15582,N_15228);
or U15976 (N_15976,N_15345,N_15213);
and U15977 (N_15977,N_15311,N_15452);
xnor U15978 (N_15978,N_15595,N_15537);
nand U15979 (N_15979,N_15540,N_15495);
nand U15980 (N_15980,N_15346,N_15265);
and U15981 (N_15981,N_15429,N_15250);
xnor U15982 (N_15982,N_15467,N_15496);
nand U15983 (N_15983,N_15535,N_15396);
xor U15984 (N_15984,N_15477,N_15595);
and U15985 (N_15985,N_15481,N_15324);
or U15986 (N_15986,N_15328,N_15527);
or U15987 (N_15987,N_15516,N_15414);
xnor U15988 (N_15988,N_15543,N_15493);
or U15989 (N_15989,N_15560,N_15359);
or U15990 (N_15990,N_15238,N_15208);
and U15991 (N_15991,N_15365,N_15485);
nor U15992 (N_15992,N_15512,N_15232);
and U15993 (N_15993,N_15308,N_15393);
nor U15994 (N_15994,N_15319,N_15391);
xor U15995 (N_15995,N_15290,N_15578);
and U15996 (N_15996,N_15438,N_15489);
xor U15997 (N_15997,N_15321,N_15269);
nor U15998 (N_15998,N_15414,N_15210);
nor U15999 (N_15999,N_15492,N_15413);
nor U16000 (N_16000,N_15730,N_15717);
nand U16001 (N_16001,N_15826,N_15877);
xnor U16002 (N_16002,N_15851,N_15956);
or U16003 (N_16003,N_15873,N_15806);
and U16004 (N_16004,N_15880,N_15749);
nand U16005 (N_16005,N_15901,N_15807);
or U16006 (N_16006,N_15817,N_15603);
and U16007 (N_16007,N_15846,N_15794);
nand U16008 (N_16008,N_15709,N_15978);
xor U16009 (N_16009,N_15699,N_15975);
xor U16010 (N_16010,N_15763,N_15947);
xor U16011 (N_16011,N_15795,N_15819);
nand U16012 (N_16012,N_15813,N_15649);
or U16013 (N_16013,N_15816,N_15606);
nand U16014 (N_16014,N_15604,N_15923);
and U16015 (N_16015,N_15886,N_15928);
nand U16016 (N_16016,N_15658,N_15666);
nand U16017 (N_16017,N_15944,N_15919);
nand U16018 (N_16018,N_15702,N_15836);
nand U16019 (N_16019,N_15905,N_15645);
and U16020 (N_16020,N_15661,N_15866);
or U16021 (N_16021,N_15825,N_15933);
and U16022 (N_16022,N_15850,N_15861);
xnor U16023 (N_16023,N_15954,N_15829);
xnor U16024 (N_16024,N_15963,N_15692);
xnor U16025 (N_16025,N_15831,N_15881);
nand U16026 (N_16026,N_15788,N_15799);
nand U16027 (N_16027,N_15811,N_15776);
or U16028 (N_16028,N_15862,N_15700);
nand U16029 (N_16029,N_15659,N_15821);
and U16030 (N_16030,N_15753,N_15674);
nand U16031 (N_16031,N_15999,N_15609);
and U16032 (N_16032,N_15723,N_15654);
or U16033 (N_16033,N_15728,N_15926);
nor U16034 (N_16034,N_15874,N_15959);
and U16035 (N_16035,N_15958,N_15859);
nor U16036 (N_16036,N_15962,N_15839);
nand U16037 (N_16037,N_15968,N_15631);
xor U16038 (N_16038,N_15619,N_15929);
nor U16039 (N_16039,N_15745,N_15747);
nand U16040 (N_16040,N_15814,N_15852);
xnor U16041 (N_16041,N_15685,N_15868);
nand U16042 (N_16042,N_15610,N_15760);
nand U16043 (N_16043,N_15894,N_15650);
xor U16044 (N_16044,N_15774,N_15693);
nor U16045 (N_16045,N_15718,N_15639);
nor U16046 (N_16046,N_15884,N_15720);
nor U16047 (N_16047,N_15969,N_15696);
xnor U16048 (N_16048,N_15653,N_15707);
nor U16049 (N_16049,N_15917,N_15634);
and U16050 (N_16050,N_15855,N_15823);
or U16051 (N_16051,N_15660,N_15784);
and U16052 (N_16052,N_15725,N_15988);
nor U16053 (N_16053,N_15927,N_15907);
xor U16054 (N_16054,N_15620,N_15986);
or U16055 (N_16055,N_15783,N_15942);
or U16056 (N_16056,N_15759,N_15902);
xnor U16057 (N_16057,N_15970,N_15845);
and U16058 (N_16058,N_15936,N_15945);
xnor U16059 (N_16059,N_15980,N_15990);
nand U16060 (N_16060,N_15695,N_15883);
nand U16061 (N_16061,N_15792,N_15913);
or U16062 (N_16062,N_15912,N_15617);
nand U16063 (N_16063,N_15853,N_15683);
and U16064 (N_16064,N_15726,N_15681);
nor U16065 (N_16065,N_15847,N_15734);
and U16066 (N_16066,N_15885,N_15729);
or U16067 (N_16067,N_15614,N_15932);
xor U16068 (N_16068,N_15808,N_15744);
nand U16069 (N_16069,N_15967,N_15899);
and U16070 (N_16070,N_15870,N_15757);
nand U16071 (N_16071,N_15641,N_15764);
nand U16072 (N_16072,N_15882,N_15798);
or U16073 (N_16073,N_15727,N_15930);
nor U16074 (N_16074,N_15860,N_15979);
xor U16075 (N_16075,N_15671,N_15876);
nor U16076 (N_16076,N_15837,N_15964);
nor U16077 (N_16077,N_15697,N_15626);
xor U16078 (N_16078,N_15663,N_15676);
nor U16079 (N_16079,N_15624,N_15678);
nor U16080 (N_16080,N_15736,N_15731);
nand U16081 (N_16081,N_15655,N_15898);
and U16082 (N_16082,N_15843,N_15890);
nor U16083 (N_16083,N_15849,N_15906);
nor U16084 (N_16084,N_15686,N_15949);
xor U16085 (N_16085,N_15802,N_15743);
nand U16086 (N_16086,N_15935,N_15690);
nor U16087 (N_16087,N_15698,N_15952);
nor U16088 (N_16088,N_15780,N_15710);
nor U16089 (N_16089,N_15721,N_15995);
xor U16090 (N_16090,N_15937,N_15976);
and U16091 (N_16091,N_15679,N_15801);
or U16092 (N_16092,N_15623,N_15786);
and U16093 (N_16093,N_15787,N_15818);
and U16094 (N_16094,N_15955,N_15946);
nand U16095 (N_16095,N_15869,N_15835);
xnor U16096 (N_16096,N_15943,N_15785);
nor U16097 (N_16097,N_15633,N_15684);
nor U16098 (N_16098,N_15605,N_15887);
and U16099 (N_16099,N_15939,N_15992);
or U16100 (N_16100,N_15878,N_15998);
nand U16101 (N_16101,N_15694,N_15983);
nor U16102 (N_16102,N_15652,N_15800);
xnor U16103 (N_16103,N_15618,N_15613);
nand U16104 (N_16104,N_15796,N_15803);
nand U16105 (N_16105,N_15770,N_15600);
xnor U16106 (N_16106,N_15879,N_15948);
nor U16107 (N_16107,N_15965,N_15724);
or U16108 (N_16108,N_15656,N_15682);
or U16109 (N_16109,N_15782,N_15896);
or U16110 (N_16110,N_15601,N_15889);
or U16111 (N_16111,N_15841,N_15820);
nor U16112 (N_16112,N_15621,N_15767);
xnor U16113 (N_16113,N_15891,N_15822);
nor U16114 (N_16114,N_15922,N_15857);
nand U16115 (N_16115,N_15925,N_15677);
and U16116 (N_16116,N_15627,N_15810);
and U16117 (N_16117,N_15758,N_15672);
xor U16118 (N_16118,N_15625,N_15914);
nor U16119 (N_16119,N_15765,N_15966);
xnor U16120 (N_16120,N_15797,N_15670);
and U16121 (N_16121,N_15704,N_15608);
nand U16122 (N_16122,N_15971,N_15643);
and U16123 (N_16123,N_15669,N_15637);
or U16124 (N_16124,N_15804,N_15775);
nor U16125 (N_16125,N_15675,N_15646);
nor U16126 (N_16126,N_15773,N_15602);
and U16127 (N_16127,N_15838,N_15994);
and U16128 (N_16128,N_15708,N_15630);
nand U16129 (N_16129,N_15858,N_15715);
nand U16130 (N_16130,N_15746,N_15742);
or U16131 (N_16131,N_15647,N_15974);
xor U16132 (N_16132,N_15812,N_15716);
nor U16133 (N_16133,N_15739,N_15738);
xnor U16134 (N_16134,N_15931,N_15805);
and U16135 (N_16135,N_15636,N_15916);
and U16136 (N_16136,N_15635,N_15934);
and U16137 (N_16137,N_15832,N_15993);
xnor U16138 (N_16138,N_15960,N_15793);
nor U16139 (N_16139,N_15893,N_15701);
or U16140 (N_16140,N_15789,N_15953);
nand U16141 (N_16141,N_15688,N_15856);
or U16142 (N_16142,N_15622,N_15985);
nor U16143 (N_16143,N_15973,N_15827);
and U16144 (N_16144,N_15834,N_15915);
or U16145 (N_16145,N_15703,N_15778);
nor U16146 (N_16146,N_15651,N_15909);
xor U16147 (N_16147,N_15900,N_15673);
nor U16148 (N_16148,N_15872,N_15779);
and U16149 (N_16149,N_15712,N_15769);
and U16150 (N_16150,N_15781,N_15908);
or U16151 (N_16151,N_15719,N_15830);
nand U16152 (N_16152,N_15828,N_15733);
xnor U16153 (N_16153,N_15997,N_15640);
xor U16154 (N_16154,N_15981,N_15903);
xor U16155 (N_16155,N_15748,N_15918);
xnor U16156 (N_16156,N_15689,N_15977);
xnor U16157 (N_16157,N_15750,N_15754);
xnor U16158 (N_16158,N_15612,N_15895);
xor U16159 (N_16159,N_15951,N_15991);
xor U16160 (N_16160,N_15972,N_15809);
nor U16161 (N_16161,N_15768,N_15833);
and U16162 (N_16162,N_15615,N_15888);
xor U16163 (N_16163,N_15941,N_15665);
nor U16164 (N_16164,N_15735,N_15867);
or U16165 (N_16165,N_15705,N_15611);
nor U16166 (N_16166,N_15629,N_15854);
xnor U16167 (N_16167,N_15755,N_15940);
and U16168 (N_16168,N_15989,N_15824);
or U16169 (N_16169,N_15657,N_15911);
or U16170 (N_16170,N_15687,N_15722);
nor U16171 (N_16171,N_15844,N_15987);
nor U16172 (N_16172,N_15741,N_15642);
nor U16173 (N_16173,N_15713,N_15751);
and U16174 (N_16174,N_15732,N_15737);
xor U16175 (N_16175,N_15950,N_15772);
xor U16176 (N_16176,N_15644,N_15662);
and U16177 (N_16177,N_15815,N_15897);
xor U16178 (N_16178,N_15777,N_15982);
nor U16179 (N_16179,N_15910,N_15924);
and U16180 (N_16180,N_15961,N_15766);
and U16181 (N_16181,N_15628,N_15752);
or U16182 (N_16182,N_15864,N_15842);
and U16183 (N_16183,N_15848,N_15711);
nand U16184 (N_16184,N_15791,N_15865);
nor U16185 (N_16185,N_15840,N_15771);
nor U16186 (N_16186,N_15667,N_15680);
and U16187 (N_16187,N_15648,N_15714);
or U16188 (N_16188,N_15638,N_15875);
nand U16189 (N_16189,N_15668,N_15957);
or U16190 (N_16190,N_15921,N_15616);
and U16191 (N_16191,N_15984,N_15904);
and U16192 (N_16192,N_15761,N_15756);
or U16193 (N_16193,N_15762,N_15691);
or U16194 (N_16194,N_15632,N_15938);
nand U16195 (N_16195,N_15790,N_15664);
nand U16196 (N_16196,N_15871,N_15892);
xnor U16197 (N_16197,N_15740,N_15706);
xnor U16198 (N_16198,N_15607,N_15996);
xor U16199 (N_16199,N_15920,N_15863);
nand U16200 (N_16200,N_15663,N_15776);
xor U16201 (N_16201,N_15848,N_15824);
or U16202 (N_16202,N_15770,N_15967);
xnor U16203 (N_16203,N_15984,N_15945);
nor U16204 (N_16204,N_15937,N_15842);
nor U16205 (N_16205,N_15633,N_15852);
nand U16206 (N_16206,N_15807,N_15962);
nor U16207 (N_16207,N_15613,N_15765);
nand U16208 (N_16208,N_15964,N_15779);
and U16209 (N_16209,N_15920,N_15663);
nand U16210 (N_16210,N_15832,N_15867);
nor U16211 (N_16211,N_15847,N_15756);
nand U16212 (N_16212,N_15820,N_15697);
nand U16213 (N_16213,N_15914,N_15902);
xor U16214 (N_16214,N_15676,N_15951);
or U16215 (N_16215,N_15623,N_15614);
nand U16216 (N_16216,N_15712,N_15706);
or U16217 (N_16217,N_15800,N_15620);
or U16218 (N_16218,N_15914,N_15794);
or U16219 (N_16219,N_15785,N_15946);
and U16220 (N_16220,N_15809,N_15964);
or U16221 (N_16221,N_15636,N_15965);
nor U16222 (N_16222,N_15802,N_15936);
nand U16223 (N_16223,N_15635,N_15909);
or U16224 (N_16224,N_15937,N_15741);
and U16225 (N_16225,N_15668,N_15942);
xnor U16226 (N_16226,N_15938,N_15830);
xnor U16227 (N_16227,N_15680,N_15938);
nand U16228 (N_16228,N_15700,N_15717);
and U16229 (N_16229,N_15841,N_15842);
and U16230 (N_16230,N_15709,N_15725);
and U16231 (N_16231,N_15735,N_15659);
xor U16232 (N_16232,N_15719,N_15952);
or U16233 (N_16233,N_15864,N_15887);
and U16234 (N_16234,N_15739,N_15788);
xor U16235 (N_16235,N_15938,N_15693);
or U16236 (N_16236,N_15766,N_15638);
nand U16237 (N_16237,N_15934,N_15913);
or U16238 (N_16238,N_15789,N_15816);
nand U16239 (N_16239,N_15869,N_15998);
or U16240 (N_16240,N_15654,N_15963);
nor U16241 (N_16241,N_15800,N_15632);
and U16242 (N_16242,N_15684,N_15801);
or U16243 (N_16243,N_15987,N_15688);
nor U16244 (N_16244,N_15970,N_15957);
nand U16245 (N_16245,N_15828,N_15989);
and U16246 (N_16246,N_15687,N_15819);
nand U16247 (N_16247,N_15845,N_15954);
and U16248 (N_16248,N_15973,N_15762);
and U16249 (N_16249,N_15903,N_15902);
and U16250 (N_16250,N_15768,N_15619);
or U16251 (N_16251,N_15860,N_15997);
and U16252 (N_16252,N_15676,N_15693);
or U16253 (N_16253,N_15756,N_15867);
nand U16254 (N_16254,N_15753,N_15762);
or U16255 (N_16255,N_15902,N_15623);
nand U16256 (N_16256,N_15886,N_15604);
xnor U16257 (N_16257,N_15790,N_15768);
and U16258 (N_16258,N_15748,N_15684);
xor U16259 (N_16259,N_15769,N_15725);
and U16260 (N_16260,N_15931,N_15946);
or U16261 (N_16261,N_15742,N_15860);
or U16262 (N_16262,N_15616,N_15951);
nand U16263 (N_16263,N_15991,N_15603);
xor U16264 (N_16264,N_15756,N_15943);
nand U16265 (N_16265,N_15957,N_15848);
nor U16266 (N_16266,N_15695,N_15767);
xor U16267 (N_16267,N_15850,N_15977);
nor U16268 (N_16268,N_15644,N_15947);
nor U16269 (N_16269,N_15739,N_15850);
or U16270 (N_16270,N_15692,N_15754);
and U16271 (N_16271,N_15919,N_15914);
xnor U16272 (N_16272,N_15726,N_15896);
and U16273 (N_16273,N_15771,N_15959);
nor U16274 (N_16274,N_15812,N_15658);
xnor U16275 (N_16275,N_15819,N_15959);
xor U16276 (N_16276,N_15818,N_15635);
nand U16277 (N_16277,N_15796,N_15930);
nand U16278 (N_16278,N_15830,N_15732);
xor U16279 (N_16279,N_15950,N_15761);
xor U16280 (N_16280,N_15858,N_15882);
or U16281 (N_16281,N_15872,N_15806);
and U16282 (N_16282,N_15871,N_15760);
nor U16283 (N_16283,N_15971,N_15821);
xnor U16284 (N_16284,N_15928,N_15915);
and U16285 (N_16285,N_15939,N_15798);
or U16286 (N_16286,N_15900,N_15647);
nor U16287 (N_16287,N_15923,N_15848);
nor U16288 (N_16288,N_15720,N_15863);
and U16289 (N_16289,N_15939,N_15854);
nor U16290 (N_16290,N_15678,N_15847);
xnor U16291 (N_16291,N_15625,N_15963);
xor U16292 (N_16292,N_15679,N_15968);
and U16293 (N_16293,N_15692,N_15676);
xnor U16294 (N_16294,N_15970,N_15889);
xnor U16295 (N_16295,N_15667,N_15641);
xnor U16296 (N_16296,N_15881,N_15732);
and U16297 (N_16297,N_15700,N_15803);
or U16298 (N_16298,N_15741,N_15748);
nand U16299 (N_16299,N_15642,N_15668);
nand U16300 (N_16300,N_15628,N_15936);
nand U16301 (N_16301,N_15908,N_15680);
nand U16302 (N_16302,N_15710,N_15901);
nor U16303 (N_16303,N_15609,N_15752);
xor U16304 (N_16304,N_15918,N_15740);
and U16305 (N_16305,N_15934,N_15943);
nand U16306 (N_16306,N_15760,N_15969);
or U16307 (N_16307,N_15683,N_15831);
or U16308 (N_16308,N_15999,N_15819);
or U16309 (N_16309,N_15822,N_15858);
or U16310 (N_16310,N_15694,N_15776);
nor U16311 (N_16311,N_15968,N_15694);
xor U16312 (N_16312,N_15625,N_15835);
nor U16313 (N_16313,N_15603,N_15955);
nand U16314 (N_16314,N_15719,N_15757);
or U16315 (N_16315,N_15741,N_15885);
nor U16316 (N_16316,N_15942,N_15817);
nand U16317 (N_16317,N_15860,N_15727);
nand U16318 (N_16318,N_15697,N_15843);
and U16319 (N_16319,N_15734,N_15812);
and U16320 (N_16320,N_15638,N_15753);
nor U16321 (N_16321,N_15988,N_15924);
nand U16322 (N_16322,N_15649,N_15976);
and U16323 (N_16323,N_15753,N_15678);
nor U16324 (N_16324,N_15627,N_15863);
or U16325 (N_16325,N_15779,N_15613);
and U16326 (N_16326,N_15833,N_15955);
and U16327 (N_16327,N_15664,N_15793);
nor U16328 (N_16328,N_15725,N_15637);
nand U16329 (N_16329,N_15912,N_15768);
and U16330 (N_16330,N_15866,N_15711);
nand U16331 (N_16331,N_15840,N_15960);
or U16332 (N_16332,N_15890,N_15728);
xnor U16333 (N_16333,N_15751,N_15877);
nor U16334 (N_16334,N_15857,N_15630);
xnor U16335 (N_16335,N_15756,N_15775);
and U16336 (N_16336,N_15723,N_15637);
nand U16337 (N_16337,N_15966,N_15956);
nand U16338 (N_16338,N_15767,N_15660);
nor U16339 (N_16339,N_15953,N_15685);
xor U16340 (N_16340,N_15946,N_15659);
and U16341 (N_16341,N_15814,N_15710);
and U16342 (N_16342,N_15956,N_15603);
nor U16343 (N_16343,N_15602,N_15671);
xor U16344 (N_16344,N_15834,N_15953);
nor U16345 (N_16345,N_15805,N_15927);
xor U16346 (N_16346,N_15672,N_15643);
xor U16347 (N_16347,N_15617,N_15910);
nand U16348 (N_16348,N_15930,N_15876);
nand U16349 (N_16349,N_15796,N_15736);
xor U16350 (N_16350,N_15798,N_15896);
or U16351 (N_16351,N_15961,N_15804);
nor U16352 (N_16352,N_15870,N_15639);
and U16353 (N_16353,N_15816,N_15956);
or U16354 (N_16354,N_15976,N_15671);
nor U16355 (N_16355,N_15816,N_15685);
nand U16356 (N_16356,N_15995,N_15623);
nor U16357 (N_16357,N_15683,N_15935);
nor U16358 (N_16358,N_15667,N_15737);
nor U16359 (N_16359,N_15807,N_15974);
nor U16360 (N_16360,N_15899,N_15932);
and U16361 (N_16361,N_15669,N_15893);
xnor U16362 (N_16362,N_15825,N_15787);
xnor U16363 (N_16363,N_15854,N_15791);
nand U16364 (N_16364,N_15966,N_15680);
and U16365 (N_16365,N_15649,N_15934);
nand U16366 (N_16366,N_15717,N_15963);
and U16367 (N_16367,N_15996,N_15962);
or U16368 (N_16368,N_15855,N_15804);
xnor U16369 (N_16369,N_15896,N_15792);
or U16370 (N_16370,N_15734,N_15836);
xor U16371 (N_16371,N_15988,N_15769);
or U16372 (N_16372,N_15690,N_15926);
and U16373 (N_16373,N_15831,N_15781);
or U16374 (N_16374,N_15630,N_15836);
or U16375 (N_16375,N_15892,N_15678);
xnor U16376 (N_16376,N_15730,N_15701);
or U16377 (N_16377,N_15820,N_15927);
nand U16378 (N_16378,N_15678,N_15831);
and U16379 (N_16379,N_15820,N_15868);
nand U16380 (N_16380,N_15772,N_15728);
or U16381 (N_16381,N_15722,N_15655);
nand U16382 (N_16382,N_15709,N_15688);
and U16383 (N_16383,N_15603,N_15994);
and U16384 (N_16384,N_15673,N_15920);
xor U16385 (N_16385,N_15802,N_15884);
xnor U16386 (N_16386,N_15739,N_15863);
xnor U16387 (N_16387,N_15982,N_15730);
nand U16388 (N_16388,N_15993,N_15890);
nor U16389 (N_16389,N_15744,N_15889);
or U16390 (N_16390,N_15916,N_15754);
and U16391 (N_16391,N_15609,N_15705);
xor U16392 (N_16392,N_15695,N_15759);
and U16393 (N_16393,N_15625,N_15855);
nor U16394 (N_16394,N_15670,N_15925);
nand U16395 (N_16395,N_15638,N_15779);
and U16396 (N_16396,N_15901,N_15737);
nand U16397 (N_16397,N_15920,N_15661);
and U16398 (N_16398,N_15733,N_15692);
or U16399 (N_16399,N_15842,N_15633);
xnor U16400 (N_16400,N_16058,N_16292);
nand U16401 (N_16401,N_16187,N_16396);
nand U16402 (N_16402,N_16256,N_16259);
xnor U16403 (N_16403,N_16080,N_16209);
or U16404 (N_16404,N_16244,N_16345);
nor U16405 (N_16405,N_16068,N_16231);
or U16406 (N_16406,N_16309,N_16019);
nor U16407 (N_16407,N_16316,N_16239);
nor U16408 (N_16408,N_16198,N_16172);
and U16409 (N_16409,N_16332,N_16321);
and U16410 (N_16410,N_16092,N_16386);
or U16411 (N_16411,N_16000,N_16300);
nand U16412 (N_16412,N_16188,N_16039);
xnor U16413 (N_16413,N_16212,N_16295);
xnor U16414 (N_16414,N_16016,N_16328);
or U16415 (N_16415,N_16148,N_16296);
nand U16416 (N_16416,N_16192,N_16166);
or U16417 (N_16417,N_16369,N_16367);
or U16418 (N_16418,N_16299,N_16226);
xnor U16419 (N_16419,N_16103,N_16069);
and U16420 (N_16420,N_16252,N_16027);
nor U16421 (N_16421,N_16145,N_16325);
nand U16422 (N_16422,N_16276,N_16306);
nor U16423 (N_16423,N_16077,N_16267);
xor U16424 (N_16424,N_16125,N_16211);
and U16425 (N_16425,N_16379,N_16380);
or U16426 (N_16426,N_16186,N_16032);
or U16427 (N_16427,N_16385,N_16283);
or U16428 (N_16428,N_16261,N_16157);
xor U16429 (N_16429,N_16035,N_16288);
nand U16430 (N_16430,N_16324,N_16112);
nand U16431 (N_16431,N_16051,N_16050);
and U16432 (N_16432,N_16302,N_16353);
nor U16433 (N_16433,N_16093,N_16114);
or U16434 (N_16434,N_16098,N_16207);
nor U16435 (N_16435,N_16291,N_16201);
nand U16436 (N_16436,N_16257,N_16001);
or U16437 (N_16437,N_16010,N_16245);
and U16438 (N_16438,N_16355,N_16116);
nor U16439 (N_16439,N_16161,N_16219);
and U16440 (N_16440,N_16394,N_16247);
nor U16441 (N_16441,N_16173,N_16225);
and U16442 (N_16442,N_16313,N_16360);
xor U16443 (N_16443,N_16197,N_16237);
xor U16444 (N_16444,N_16224,N_16007);
nand U16445 (N_16445,N_16356,N_16134);
xnor U16446 (N_16446,N_16154,N_16274);
and U16447 (N_16447,N_16323,N_16193);
nand U16448 (N_16448,N_16085,N_16130);
or U16449 (N_16449,N_16253,N_16030);
or U16450 (N_16450,N_16170,N_16012);
nand U16451 (N_16451,N_16352,N_16133);
nand U16452 (N_16452,N_16311,N_16117);
and U16453 (N_16453,N_16370,N_16329);
nand U16454 (N_16454,N_16376,N_16229);
xor U16455 (N_16455,N_16189,N_16087);
or U16456 (N_16456,N_16047,N_16158);
xor U16457 (N_16457,N_16041,N_16395);
nor U16458 (N_16458,N_16287,N_16241);
nand U16459 (N_16459,N_16242,N_16095);
nor U16460 (N_16460,N_16118,N_16089);
xnor U16461 (N_16461,N_16342,N_16137);
xnor U16462 (N_16462,N_16235,N_16371);
nor U16463 (N_16463,N_16143,N_16307);
and U16464 (N_16464,N_16293,N_16390);
nand U16465 (N_16465,N_16090,N_16046);
and U16466 (N_16466,N_16375,N_16185);
xnor U16467 (N_16467,N_16020,N_16216);
nor U16468 (N_16468,N_16270,N_16009);
nor U16469 (N_16469,N_16150,N_16255);
nor U16470 (N_16470,N_16026,N_16331);
and U16471 (N_16471,N_16183,N_16123);
xor U16472 (N_16472,N_16398,N_16251);
and U16473 (N_16473,N_16358,N_16072);
nor U16474 (N_16474,N_16205,N_16322);
and U16475 (N_16475,N_16228,N_16160);
nor U16476 (N_16476,N_16124,N_16003);
nor U16477 (N_16477,N_16347,N_16122);
or U16478 (N_16478,N_16094,N_16220);
and U16479 (N_16479,N_16289,N_16024);
nand U16480 (N_16480,N_16042,N_16275);
xor U16481 (N_16481,N_16036,N_16061);
nor U16482 (N_16482,N_16344,N_16002);
nand U16483 (N_16483,N_16233,N_16073);
xnor U16484 (N_16484,N_16281,N_16031);
and U16485 (N_16485,N_16250,N_16301);
xor U16486 (N_16486,N_16303,N_16317);
nand U16487 (N_16487,N_16100,N_16204);
nor U16488 (N_16488,N_16128,N_16013);
or U16489 (N_16489,N_16146,N_16203);
nor U16490 (N_16490,N_16081,N_16343);
nand U16491 (N_16491,N_16179,N_16222);
nand U16492 (N_16492,N_16097,N_16131);
xor U16493 (N_16493,N_16254,N_16140);
and U16494 (N_16494,N_16159,N_16333);
and U16495 (N_16495,N_16071,N_16164);
nor U16496 (N_16496,N_16298,N_16004);
xnor U16497 (N_16497,N_16372,N_16113);
or U16498 (N_16498,N_16389,N_16162);
xor U16499 (N_16499,N_16149,N_16091);
nor U16500 (N_16500,N_16282,N_16266);
nand U16501 (N_16501,N_16327,N_16104);
nor U16502 (N_16502,N_16215,N_16320);
xor U16503 (N_16503,N_16199,N_16297);
xnor U16504 (N_16504,N_16284,N_16147);
nand U16505 (N_16505,N_16070,N_16022);
or U16506 (N_16506,N_16017,N_16008);
xor U16507 (N_16507,N_16191,N_16121);
and U16508 (N_16508,N_16045,N_16221);
or U16509 (N_16509,N_16110,N_16078);
nand U16510 (N_16510,N_16277,N_16060);
nand U16511 (N_16511,N_16101,N_16037);
nand U16512 (N_16512,N_16139,N_16065);
or U16513 (N_16513,N_16377,N_16048);
and U16514 (N_16514,N_16136,N_16054);
and U16515 (N_16515,N_16373,N_16105);
nand U16516 (N_16516,N_16057,N_16388);
or U16517 (N_16517,N_16273,N_16319);
and U16518 (N_16518,N_16168,N_16314);
nand U16519 (N_16519,N_16264,N_16176);
and U16520 (N_16520,N_16337,N_16208);
or U16521 (N_16521,N_16269,N_16310);
or U16522 (N_16522,N_16141,N_16397);
and U16523 (N_16523,N_16082,N_16290);
nand U16524 (N_16524,N_16387,N_16362);
or U16525 (N_16525,N_16243,N_16006);
or U16526 (N_16526,N_16234,N_16218);
and U16527 (N_16527,N_16294,N_16318);
xor U16528 (N_16528,N_16153,N_16248);
xor U16529 (N_16529,N_16126,N_16106);
or U16530 (N_16530,N_16062,N_16079);
xor U16531 (N_16531,N_16383,N_16088);
and U16532 (N_16532,N_16053,N_16015);
and U16533 (N_16533,N_16262,N_16336);
and U16534 (N_16534,N_16338,N_16005);
nor U16535 (N_16535,N_16393,N_16346);
nor U16536 (N_16536,N_16305,N_16210);
and U16537 (N_16537,N_16206,N_16272);
nand U16538 (N_16538,N_16349,N_16392);
nand U16539 (N_16539,N_16308,N_16359);
nand U16540 (N_16540,N_16232,N_16044);
or U16541 (N_16541,N_16240,N_16304);
xnor U16542 (N_16542,N_16155,N_16363);
xor U16543 (N_16543,N_16357,N_16075);
and U16544 (N_16544,N_16107,N_16011);
nor U16545 (N_16545,N_16135,N_16217);
or U16546 (N_16546,N_16230,N_16102);
and U16547 (N_16547,N_16055,N_16200);
or U16548 (N_16548,N_16194,N_16351);
and U16549 (N_16549,N_16144,N_16120);
xnor U16550 (N_16550,N_16064,N_16014);
nor U16551 (N_16551,N_16182,N_16067);
or U16552 (N_16552,N_16214,N_16056);
and U16553 (N_16553,N_16127,N_16119);
nand U16554 (N_16554,N_16021,N_16043);
or U16555 (N_16555,N_16341,N_16029);
xor U16556 (N_16556,N_16086,N_16028);
xnor U16557 (N_16557,N_16315,N_16018);
nor U16558 (N_16558,N_16171,N_16227);
xnor U16559 (N_16559,N_16178,N_16181);
xnor U16560 (N_16560,N_16034,N_16278);
nor U16561 (N_16561,N_16350,N_16268);
xnor U16562 (N_16562,N_16165,N_16142);
and U16563 (N_16563,N_16156,N_16196);
nand U16564 (N_16564,N_16354,N_16132);
xnor U16565 (N_16565,N_16258,N_16213);
and U16566 (N_16566,N_16190,N_16083);
and U16567 (N_16567,N_16151,N_16382);
nand U16568 (N_16568,N_16052,N_16152);
or U16569 (N_16569,N_16368,N_16374);
xnor U16570 (N_16570,N_16169,N_16384);
or U16571 (N_16571,N_16175,N_16339);
and U16572 (N_16572,N_16285,N_16040);
or U16573 (N_16573,N_16108,N_16115);
and U16574 (N_16574,N_16334,N_16038);
xnor U16575 (N_16575,N_16059,N_16049);
xnor U16576 (N_16576,N_16111,N_16280);
or U16577 (N_16577,N_16260,N_16138);
and U16578 (N_16578,N_16279,N_16109);
xor U16579 (N_16579,N_16174,N_16249);
and U16580 (N_16580,N_16366,N_16364);
or U16581 (N_16581,N_16025,N_16084);
nand U16582 (N_16582,N_16236,N_16180);
and U16583 (N_16583,N_16381,N_16023);
xnor U16584 (N_16584,N_16033,N_16361);
nor U16585 (N_16585,N_16391,N_16184);
nor U16586 (N_16586,N_16238,N_16163);
nor U16587 (N_16587,N_16312,N_16202);
xnor U16588 (N_16588,N_16223,N_16365);
xnor U16589 (N_16589,N_16263,N_16066);
nor U16590 (N_16590,N_16246,N_16195);
and U16591 (N_16591,N_16326,N_16378);
nor U16592 (N_16592,N_16099,N_16340);
or U16593 (N_16593,N_16286,N_16063);
nand U16594 (N_16594,N_16076,N_16167);
or U16595 (N_16595,N_16265,N_16096);
and U16596 (N_16596,N_16271,N_16177);
and U16597 (N_16597,N_16330,N_16335);
and U16598 (N_16598,N_16348,N_16129);
and U16599 (N_16599,N_16074,N_16399);
xor U16600 (N_16600,N_16110,N_16094);
nor U16601 (N_16601,N_16250,N_16333);
nand U16602 (N_16602,N_16088,N_16318);
or U16603 (N_16603,N_16054,N_16195);
xnor U16604 (N_16604,N_16166,N_16354);
and U16605 (N_16605,N_16269,N_16350);
nand U16606 (N_16606,N_16037,N_16273);
or U16607 (N_16607,N_16321,N_16059);
xnor U16608 (N_16608,N_16257,N_16272);
or U16609 (N_16609,N_16123,N_16180);
or U16610 (N_16610,N_16075,N_16017);
xnor U16611 (N_16611,N_16161,N_16224);
nor U16612 (N_16612,N_16006,N_16388);
or U16613 (N_16613,N_16180,N_16284);
nor U16614 (N_16614,N_16030,N_16231);
nand U16615 (N_16615,N_16052,N_16245);
nand U16616 (N_16616,N_16352,N_16129);
nor U16617 (N_16617,N_16008,N_16162);
nand U16618 (N_16618,N_16134,N_16378);
xnor U16619 (N_16619,N_16283,N_16117);
nor U16620 (N_16620,N_16307,N_16062);
or U16621 (N_16621,N_16364,N_16029);
nand U16622 (N_16622,N_16173,N_16123);
nor U16623 (N_16623,N_16044,N_16125);
and U16624 (N_16624,N_16190,N_16208);
or U16625 (N_16625,N_16374,N_16390);
xnor U16626 (N_16626,N_16283,N_16319);
nand U16627 (N_16627,N_16047,N_16138);
xnor U16628 (N_16628,N_16318,N_16013);
nor U16629 (N_16629,N_16320,N_16336);
and U16630 (N_16630,N_16105,N_16039);
nor U16631 (N_16631,N_16167,N_16056);
and U16632 (N_16632,N_16007,N_16119);
or U16633 (N_16633,N_16305,N_16369);
nand U16634 (N_16634,N_16324,N_16301);
xor U16635 (N_16635,N_16003,N_16170);
xnor U16636 (N_16636,N_16223,N_16315);
nand U16637 (N_16637,N_16388,N_16239);
nor U16638 (N_16638,N_16080,N_16075);
nor U16639 (N_16639,N_16237,N_16019);
or U16640 (N_16640,N_16147,N_16057);
and U16641 (N_16641,N_16109,N_16139);
nand U16642 (N_16642,N_16346,N_16024);
nand U16643 (N_16643,N_16133,N_16383);
xnor U16644 (N_16644,N_16056,N_16121);
nor U16645 (N_16645,N_16306,N_16388);
nor U16646 (N_16646,N_16319,N_16235);
nand U16647 (N_16647,N_16149,N_16009);
nor U16648 (N_16648,N_16006,N_16012);
and U16649 (N_16649,N_16066,N_16372);
xnor U16650 (N_16650,N_16272,N_16320);
xor U16651 (N_16651,N_16316,N_16019);
nor U16652 (N_16652,N_16146,N_16184);
xnor U16653 (N_16653,N_16004,N_16354);
and U16654 (N_16654,N_16172,N_16330);
xor U16655 (N_16655,N_16031,N_16236);
nor U16656 (N_16656,N_16067,N_16346);
and U16657 (N_16657,N_16359,N_16197);
nor U16658 (N_16658,N_16169,N_16237);
nor U16659 (N_16659,N_16176,N_16025);
xor U16660 (N_16660,N_16243,N_16027);
xor U16661 (N_16661,N_16224,N_16397);
or U16662 (N_16662,N_16054,N_16368);
xor U16663 (N_16663,N_16142,N_16333);
nor U16664 (N_16664,N_16277,N_16154);
nor U16665 (N_16665,N_16215,N_16024);
nor U16666 (N_16666,N_16391,N_16019);
nor U16667 (N_16667,N_16168,N_16118);
xnor U16668 (N_16668,N_16029,N_16287);
xor U16669 (N_16669,N_16052,N_16129);
nor U16670 (N_16670,N_16094,N_16172);
or U16671 (N_16671,N_16248,N_16117);
and U16672 (N_16672,N_16066,N_16031);
and U16673 (N_16673,N_16100,N_16127);
nor U16674 (N_16674,N_16166,N_16082);
nand U16675 (N_16675,N_16230,N_16307);
nor U16676 (N_16676,N_16323,N_16119);
nand U16677 (N_16677,N_16306,N_16045);
or U16678 (N_16678,N_16099,N_16161);
xor U16679 (N_16679,N_16019,N_16208);
xor U16680 (N_16680,N_16085,N_16183);
nor U16681 (N_16681,N_16076,N_16026);
nor U16682 (N_16682,N_16075,N_16074);
nand U16683 (N_16683,N_16172,N_16261);
and U16684 (N_16684,N_16098,N_16368);
xor U16685 (N_16685,N_16221,N_16236);
nor U16686 (N_16686,N_16291,N_16070);
xnor U16687 (N_16687,N_16110,N_16238);
nor U16688 (N_16688,N_16318,N_16378);
nor U16689 (N_16689,N_16371,N_16364);
nor U16690 (N_16690,N_16399,N_16351);
nand U16691 (N_16691,N_16016,N_16092);
or U16692 (N_16692,N_16073,N_16080);
xnor U16693 (N_16693,N_16092,N_16221);
nand U16694 (N_16694,N_16262,N_16270);
or U16695 (N_16695,N_16304,N_16014);
and U16696 (N_16696,N_16198,N_16065);
nor U16697 (N_16697,N_16270,N_16036);
xnor U16698 (N_16698,N_16389,N_16396);
xnor U16699 (N_16699,N_16327,N_16315);
and U16700 (N_16700,N_16339,N_16162);
nor U16701 (N_16701,N_16317,N_16287);
or U16702 (N_16702,N_16173,N_16020);
and U16703 (N_16703,N_16079,N_16140);
and U16704 (N_16704,N_16001,N_16193);
and U16705 (N_16705,N_16323,N_16366);
nor U16706 (N_16706,N_16288,N_16253);
xor U16707 (N_16707,N_16098,N_16023);
xor U16708 (N_16708,N_16208,N_16304);
or U16709 (N_16709,N_16266,N_16071);
xor U16710 (N_16710,N_16240,N_16341);
xnor U16711 (N_16711,N_16270,N_16213);
nor U16712 (N_16712,N_16344,N_16243);
nand U16713 (N_16713,N_16350,N_16155);
and U16714 (N_16714,N_16188,N_16000);
nand U16715 (N_16715,N_16124,N_16192);
nand U16716 (N_16716,N_16162,N_16102);
or U16717 (N_16717,N_16061,N_16157);
nor U16718 (N_16718,N_16255,N_16021);
nor U16719 (N_16719,N_16228,N_16060);
xor U16720 (N_16720,N_16130,N_16003);
and U16721 (N_16721,N_16278,N_16221);
and U16722 (N_16722,N_16092,N_16170);
or U16723 (N_16723,N_16005,N_16390);
and U16724 (N_16724,N_16039,N_16357);
nand U16725 (N_16725,N_16222,N_16206);
or U16726 (N_16726,N_16039,N_16374);
or U16727 (N_16727,N_16231,N_16017);
and U16728 (N_16728,N_16267,N_16140);
or U16729 (N_16729,N_16002,N_16015);
nand U16730 (N_16730,N_16102,N_16304);
nand U16731 (N_16731,N_16264,N_16247);
and U16732 (N_16732,N_16387,N_16263);
nor U16733 (N_16733,N_16032,N_16288);
or U16734 (N_16734,N_16223,N_16375);
xnor U16735 (N_16735,N_16113,N_16115);
and U16736 (N_16736,N_16160,N_16318);
nor U16737 (N_16737,N_16305,N_16259);
xor U16738 (N_16738,N_16209,N_16225);
nor U16739 (N_16739,N_16111,N_16126);
nand U16740 (N_16740,N_16162,N_16174);
nor U16741 (N_16741,N_16218,N_16060);
nor U16742 (N_16742,N_16073,N_16349);
nor U16743 (N_16743,N_16088,N_16301);
xnor U16744 (N_16744,N_16013,N_16119);
xor U16745 (N_16745,N_16366,N_16091);
and U16746 (N_16746,N_16378,N_16014);
nand U16747 (N_16747,N_16213,N_16044);
and U16748 (N_16748,N_16278,N_16395);
xor U16749 (N_16749,N_16103,N_16019);
and U16750 (N_16750,N_16270,N_16071);
nand U16751 (N_16751,N_16058,N_16368);
or U16752 (N_16752,N_16097,N_16115);
nor U16753 (N_16753,N_16018,N_16340);
nor U16754 (N_16754,N_16372,N_16029);
and U16755 (N_16755,N_16024,N_16371);
nand U16756 (N_16756,N_16281,N_16246);
nand U16757 (N_16757,N_16375,N_16363);
or U16758 (N_16758,N_16182,N_16277);
or U16759 (N_16759,N_16141,N_16148);
xor U16760 (N_16760,N_16199,N_16322);
nor U16761 (N_16761,N_16105,N_16007);
nor U16762 (N_16762,N_16121,N_16054);
xor U16763 (N_16763,N_16023,N_16165);
nor U16764 (N_16764,N_16383,N_16326);
nor U16765 (N_16765,N_16050,N_16321);
nor U16766 (N_16766,N_16039,N_16021);
or U16767 (N_16767,N_16235,N_16389);
or U16768 (N_16768,N_16347,N_16133);
xnor U16769 (N_16769,N_16060,N_16002);
nor U16770 (N_16770,N_16024,N_16373);
and U16771 (N_16771,N_16094,N_16282);
nor U16772 (N_16772,N_16305,N_16108);
nand U16773 (N_16773,N_16098,N_16129);
and U16774 (N_16774,N_16327,N_16383);
and U16775 (N_16775,N_16114,N_16116);
xor U16776 (N_16776,N_16274,N_16322);
or U16777 (N_16777,N_16305,N_16134);
xnor U16778 (N_16778,N_16166,N_16216);
or U16779 (N_16779,N_16230,N_16114);
nor U16780 (N_16780,N_16132,N_16393);
xnor U16781 (N_16781,N_16117,N_16127);
nor U16782 (N_16782,N_16058,N_16032);
nand U16783 (N_16783,N_16300,N_16034);
and U16784 (N_16784,N_16223,N_16366);
and U16785 (N_16785,N_16288,N_16258);
nand U16786 (N_16786,N_16098,N_16385);
and U16787 (N_16787,N_16143,N_16395);
nand U16788 (N_16788,N_16208,N_16261);
nor U16789 (N_16789,N_16387,N_16299);
xnor U16790 (N_16790,N_16192,N_16104);
nand U16791 (N_16791,N_16190,N_16146);
or U16792 (N_16792,N_16094,N_16359);
nand U16793 (N_16793,N_16372,N_16086);
and U16794 (N_16794,N_16124,N_16069);
xnor U16795 (N_16795,N_16038,N_16296);
or U16796 (N_16796,N_16175,N_16135);
nand U16797 (N_16797,N_16050,N_16302);
nor U16798 (N_16798,N_16278,N_16242);
and U16799 (N_16799,N_16051,N_16225);
nand U16800 (N_16800,N_16418,N_16650);
or U16801 (N_16801,N_16474,N_16628);
and U16802 (N_16802,N_16477,N_16454);
nand U16803 (N_16803,N_16589,N_16508);
and U16804 (N_16804,N_16700,N_16750);
and U16805 (N_16805,N_16408,N_16681);
nor U16806 (N_16806,N_16780,N_16459);
or U16807 (N_16807,N_16555,N_16666);
and U16808 (N_16808,N_16724,N_16582);
and U16809 (N_16809,N_16580,N_16514);
xnor U16810 (N_16810,N_16435,N_16601);
and U16811 (N_16811,N_16787,N_16438);
xnor U16812 (N_16812,N_16558,N_16665);
xnor U16813 (N_16813,N_16563,N_16789);
nor U16814 (N_16814,N_16494,N_16691);
and U16815 (N_16815,N_16626,N_16584);
or U16816 (N_16816,N_16554,N_16766);
xnor U16817 (N_16817,N_16637,N_16442);
nand U16818 (N_16818,N_16686,N_16460);
xor U16819 (N_16819,N_16746,N_16506);
or U16820 (N_16820,N_16448,N_16549);
or U16821 (N_16821,N_16415,N_16706);
nor U16822 (N_16822,N_16577,N_16515);
or U16823 (N_16823,N_16463,N_16575);
nor U16824 (N_16824,N_16550,N_16649);
and U16825 (N_16825,N_16720,N_16597);
xor U16826 (N_16826,N_16511,N_16775);
or U16827 (N_16827,N_16736,N_16436);
or U16828 (N_16828,N_16756,N_16687);
nor U16829 (N_16829,N_16528,N_16581);
nor U16830 (N_16830,N_16531,N_16461);
xnor U16831 (N_16831,N_16598,N_16529);
or U16832 (N_16832,N_16604,N_16782);
xor U16833 (N_16833,N_16699,N_16743);
nand U16834 (N_16834,N_16496,N_16499);
or U16835 (N_16835,N_16507,N_16772);
or U16836 (N_16836,N_16771,N_16532);
nand U16837 (N_16837,N_16457,N_16505);
and U16838 (N_16838,N_16497,N_16420);
and U16839 (N_16839,N_16786,N_16530);
nor U16840 (N_16840,N_16556,N_16672);
and U16841 (N_16841,N_16472,N_16535);
xnor U16842 (N_16842,N_16546,N_16462);
nor U16843 (N_16843,N_16609,N_16657);
or U16844 (N_16844,N_16483,N_16548);
or U16845 (N_16845,N_16605,N_16762);
and U16846 (N_16846,N_16465,N_16547);
and U16847 (N_16847,N_16551,N_16446);
nand U16848 (N_16848,N_16576,N_16519);
and U16849 (N_16849,N_16553,N_16527);
and U16850 (N_16850,N_16467,N_16674);
and U16851 (N_16851,N_16659,N_16417);
or U16852 (N_16852,N_16414,N_16578);
and U16853 (N_16853,N_16748,N_16760);
xnor U16854 (N_16854,N_16450,N_16757);
nand U16855 (N_16855,N_16413,N_16595);
nand U16856 (N_16856,N_16725,N_16486);
nand U16857 (N_16857,N_16693,N_16723);
nor U16858 (N_16858,N_16492,N_16793);
and U16859 (N_16859,N_16466,N_16770);
and U16860 (N_16860,N_16468,N_16737);
nand U16861 (N_16861,N_16751,N_16721);
or U16862 (N_16862,N_16475,N_16726);
nor U16863 (N_16863,N_16685,N_16574);
nor U16864 (N_16864,N_16630,N_16664);
and U16865 (N_16865,N_16579,N_16753);
nand U16866 (N_16866,N_16570,N_16640);
and U16867 (N_16867,N_16729,N_16440);
nand U16868 (N_16868,N_16799,N_16710);
nand U16869 (N_16869,N_16641,N_16635);
or U16870 (N_16870,N_16485,N_16490);
nand U16871 (N_16871,N_16545,N_16647);
nor U16872 (N_16872,N_16404,N_16732);
and U16873 (N_16873,N_16792,N_16429);
xor U16874 (N_16874,N_16402,N_16749);
nand U16875 (N_16875,N_16670,N_16731);
nor U16876 (N_16876,N_16480,N_16716);
nor U16877 (N_16877,N_16752,N_16433);
nor U16878 (N_16878,N_16648,N_16758);
xor U16879 (N_16879,N_16608,N_16774);
nor U16880 (N_16880,N_16606,N_16719);
and U16881 (N_16881,N_16453,N_16484);
xor U16882 (N_16882,N_16524,N_16638);
or U16883 (N_16883,N_16777,N_16423);
and U16884 (N_16884,N_16416,N_16741);
and U16885 (N_16885,N_16702,N_16464);
xnor U16886 (N_16886,N_16500,N_16562);
nor U16887 (N_16887,N_16526,N_16498);
xor U16888 (N_16888,N_16487,N_16671);
nor U16889 (N_16889,N_16730,N_16619);
nand U16890 (N_16890,N_16747,N_16596);
nor U16891 (N_16891,N_16714,N_16654);
nor U16892 (N_16892,N_16411,N_16407);
nand U16893 (N_16893,N_16458,N_16540);
and U16894 (N_16894,N_16697,N_16593);
nor U16895 (N_16895,N_16481,N_16400);
or U16896 (N_16896,N_16668,N_16734);
xnor U16897 (N_16897,N_16785,N_16509);
xor U16898 (N_16898,N_16642,N_16445);
and U16899 (N_16899,N_16471,N_16684);
nand U16900 (N_16900,N_16663,N_16624);
and U16901 (N_16901,N_16425,N_16620);
and U16902 (N_16902,N_16444,N_16443);
or U16903 (N_16903,N_16561,N_16566);
nand U16904 (N_16904,N_16735,N_16560);
and U16905 (N_16905,N_16586,N_16763);
and U16906 (N_16906,N_16406,N_16738);
nand U16907 (N_16907,N_16779,N_16470);
nand U16908 (N_16908,N_16572,N_16541);
nor U16909 (N_16909,N_16431,N_16667);
and U16910 (N_16910,N_16634,N_16449);
or U16911 (N_16911,N_16502,N_16517);
nand U16912 (N_16912,N_16631,N_16653);
or U16913 (N_16913,N_16790,N_16701);
or U16914 (N_16914,N_16501,N_16590);
and U16915 (N_16915,N_16405,N_16759);
nand U16916 (N_16916,N_16569,N_16543);
nand U16917 (N_16917,N_16652,N_16504);
nor U16918 (N_16918,N_16727,N_16711);
nand U16919 (N_16919,N_16646,N_16503);
nor U16920 (N_16920,N_16669,N_16643);
or U16921 (N_16921,N_16675,N_16683);
and U16922 (N_16922,N_16542,N_16767);
nand U16923 (N_16923,N_16567,N_16441);
nor U16924 (N_16924,N_16520,N_16603);
xnor U16925 (N_16925,N_16692,N_16718);
or U16926 (N_16926,N_16455,N_16655);
or U16927 (N_16927,N_16587,N_16403);
or U16928 (N_16928,N_16476,N_16594);
nor U16929 (N_16929,N_16565,N_16493);
nor U16930 (N_16930,N_16784,N_16591);
or U16931 (N_16931,N_16522,N_16518);
xnor U16932 (N_16932,N_16409,N_16533);
nor U16933 (N_16933,N_16614,N_16645);
or U16934 (N_16934,N_16615,N_16568);
xnor U16935 (N_16935,N_16695,N_16682);
nor U16936 (N_16936,N_16797,N_16611);
nand U16937 (N_16937,N_16778,N_16717);
or U16938 (N_16938,N_16796,N_16573);
nor U16939 (N_16939,N_16539,N_16709);
nand U16940 (N_16940,N_16712,N_16610);
nor U16941 (N_16941,N_16678,N_16689);
nand U16942 (N_16942,N_16469,N_16421);
and U16943 (N_16943,N_16636,N_16708);
nor U16944 (N_16944,N_16742,N_16783);
or U16945 (N_16945,N_16625,N_16516);
xor U16946 (N_16946,N_16456,N_16617);
or U16947 (N_16947,N_16588,N_16537);
xor U16948 (N_16948,N_16536,N_16552);
or U16949 (N_16949,N_16680,N_16629);
and U16950 (N_16950,N_16739,N_16607);
xor U16951 (N_16951,N_16733,N_16510);
nor U16952 (N_16952,N_16713,N_16583);
nor U16953 (N_16953,N_16571,N_16679);
nand U16954 (N_16954,N_16776,N_16616);
or U16955 (N_16955,N_16744,N_16621);
or U16956 (N_16956,N_16622,N_16432);
nand U16957 (N_16957,N_16677,N_16754);
nor U16958 (N_16958,N_16764,N_16612);
nor U16959 (N_16959,N_16644,N_16479);
and U16960 (N_16960,N_16495,N_16427);
xnor U16961 (N_16961,N_16559,N_16639);
or U16962 (N_16962,N_16437,N_16781);
nand U16963 (N_16963,N_16534,N_16410);
xnor U16964 (N_16964,N_16694,N_16434);
nor U16965 (N_16965,N_16696,N_16632);
nor U16966 (N_16966,N_16791,N_16794);
or U16967 (N_16967,N_16525,N_16544);
nor U16968 (N_16968,N_16765,N_16656);
nor U16969 (N_16969,N_16447,N_16478);
and U16970 (N_16970,N_16660,N_16491);
nand U16971 (N_16971,N_16673,N_16651);
or U16972 (N_16972,N_16428,N_16773);
nand U16973 (N_16973,N_16745,N_16722);
xnor U16974 (N_16974,N_16488,N_16564);
nor U16975 (N_16975,N_16513,N_16419);
nor U16976 (N_16976,N_16627,N_16676);
xnor U16977 (N_16977,N_16698,N_16439);
xor U16978 (N_16978,N_16755,N_16633);
nor U16979 (N_16979,N_16512,N_16538);
or U16980 (N_16980,N_16705,N_16426);
nor U16981 (N_16981,N_16661,N_16703);
nor U16982 (N_16982,N_16422,N_16602);
or U16983 (N_16983,N_16482,N_16473);
nor U16984 (N_16984,N_16613,N_16451);
and U16985 (N_16985,N_16728,N_16430);
xnor U16986 (N_16986,N_16523,N_16769);
nor U16987 (N_16987,N_16690,N_16401);
nand U16988 (N_16988,N_16795,N_16599);
xor U16989 (N_16989,N_16704,N_16662);
xor U16990 (N_16990,N_16452,N_16707);
nor U16991 (N_16991,N_16740,N_16688);
xnor U16992 (N_16992,N_16412,N_16623);
and U16993 (N_16993,N_16600,N_16761);
and U16994 (N_16994,N_16521,N_16618);
or U16995 (N_16995,N_16489,N_16768);
xor U16996 (N_16996,N_16658,N_16557);
xnor U16997 (N_16997,N_16788,N_16585);
or U16998 (N_16998,N_16798,N_16592);
and U16999 (N_16999,N_16715,N_16424);
or U17000 (N_17000,N_16584,N_16518);
or U17001 (N_17001,N_16718,N_16578);
nor U17002 (N_17002,N_16548,N_16606);
nand U17003 (N_17003,N_16507,N_16587);
nor U17004 (N_17004,N_16589,N_16473);
and U17005 (N_17005,N_16698,N_16774);
or U17006 (N_17006,N_16459,N_16688);
or U17007 (N_17007,N_16716,N_16526);
nor U17008 (N_17008,N_16680,N_16450);
nor U17009 (N_17009,N_16547,N_16546);
or U17010 (N_17010,N_16627,N_16458);
nor U17011 (N_17011,N_16726,N_16508);
nand U17012 (N_17012,N_16686,N_16487);
xnor U17013 (N_17013,N_16493,N_16700);
nand U17014 (N_17014,N_16777,N_16630);
nor U17015 (N_17015,N_16689,N_16688);
or U17016 (N_17016,N_16424,N_16734);
or U17017 (N_17017,N_16500,N_16738);
nand U17018 (N_17018,N_16463,N_16735);
xnor U17019 (N_17019,N_16422,N_16556);
nand U17020 (N_17020,N_16587,N_16736);
nand U17021 (N_17021,N_16598,N_16474);
and U17022 (N_17022,N_16640,N_16591);
and U17023 (N_17023,N_16559,N_16444);
nand U17024 (N_17024,N_16672,N_16761);
or U17025 (N_17025,N_16470,N_16563);
nand U17026 (N_17026,N_16755,N_16754);
and U17027 (N_17027,N_16701,N_16575);
or U17028 (N_17028,N_16458,N_16429);
or U17029 (N_17029,N_16550,N_16700);
or U17030 (N_17030,N_16499,N_16509);
nor U17031 (N_17031,N_16704,N_16652);
or U17032 (N_17032,N_16545,N_16507);
nor U17033 (N_17033,N_16750,N_16680);
nor U17034 (N_17034,N_16633,N_16680);
nand U17035 (N_17035,N_16536,N_16663);
or U17036 (N_17036,N_16748,N_16771);
or U17037 (N_17037,N_16641,N_16475);
or U17038 (N_17038,N_16691,N_16671);
xor U17039 (N_17039,N_16424,N_16510);
nor U17040 (N_17040,N_16722,N_16776);
and U17041 (N_17041,N_16528,N_16702);
and U17042 (N_17042,N_16672,N_16545);
nand U17043 (N_17043,N_16594,N_16796);
or U17044 (N_17044,N_16561,N_16514);
nor U17045 (N_17045,N_16493,N_16766);
and U17046 (N_17046,N_16437,N_16491);
or U17047 (N_17047,N_16706,N_16544);
or U17048 (N_17048,N_16505,N_16484);
or U17049 (N_17049,N_16476,N_16707);
and U17050 (N_17050,N_16722,N_16504);
nor U17051 (N_17051,N_16402,N_16663);
and U17052 (N_17052,N_16635,N_16438);
xor U17053 (N_17053,N_16500,N_16430);
xor U17054 (N_17054,N_16551,N_16481);
nor U17055 (N_17055,N_16757,N_16613);
nor U17056 (N_17056,N_16653,N_16427);
or U17057 (N_17057,N_16629,N_16765);
nor U17058 (N_17058,N_16761,N_16568);
nor U17059 (N_17059,N_16584,N_16564);
and U17060 (N_17060,N_16761,N_16641);
nor U17061 (N_17061,N_16431,N_16711);
or U17062 (N_17062,N_16717,N_16699);
nor U17063 (N_17063,N_16504,N_16459);
nand U17064 (N_17064,N_16782,N_16611);
and U17065 (N_17065,N_16470,N_16493);
nor U17066 (N_17066,N_16562,N_16797);
or U17067 (N_17067,N_16426,N_16499);
and U17068 (N_17068,N_16581,N_16661);
xor U17069 (N_17069,N_16514,N_16434);
nand U17070 (N_17070,N_16554,N_16477);
or U17071 (N_17071,N_16683,N_16690);
xnor U17072 (N_17072,N_16594,N_16434);
nor U17073 (N_17073,N_16622,N_16708);
and U17074 (N_17074,N_16445,N_16544);
or U17075 (N_17075,N_16656,N_16427);
nor U17076 (N_17076,N_16680,N_16674);
nor U17077 (N_17077,N_16791,N_16490);
or U17078 (N_17078,N_16780,N_16774);
or U17079 (N_17079,N_16552,N_16682);
nand U17080 (N_17080,N_16737,N_16606);
xor U17081 (N_17081,N_16667,N_16757);
nand U17082 (N_17082,N_16751,N_16518);
or U17083 (N_17083,N_16509,N_16551);
and U17084 (N_17084,N_16438,N_16466);
or U17085 (N_17085,N_16578,N_16443);
and U17086 (N_17086,N_16657,N_16670);
and U17087 (N_17087,N_16480,N_16775);
xor U17088 (N_17088,N_16506,N_16779);
and U17089 (N_17089,N_16792,N_16727);
nor U17090 (N_17090,N_16630,N_16521);
nor U17091 (N_17091,N_16494,N_16444);
xor U17092 (N_17092,N_16797,N_16485);
and U17093 (N_17093,N_16561,N_16443);
nand U17094 (N_17094,N_16662,N_16561);
nor U17095 (N_17095,N_16462,N_16516);
nand U17096 (N_17096,N_16667,N_16547);
nor U17097 (N_17097,N_16755,N_16485);
nand U17098 (N_17098,N_16528,N_16496);
nor U17099 (N_17099,N_16650,N_16668);
xor U17100 (N_17100,N_16524,N_16633);
nand U17101 (N_17101,N_16702,N_16668);
or U17102 (N_17102,N_16551,N_16489);
nor U17103 (N_17103,N_16423,N_16692);
nor U17104 (N_17104,N_16592,N_16453);
nand U17105 (N_17105,N_16686,N_16468);
nand U17106 (N_17106,N_16474,N_16777);
nand U17107 (N_17107,N_16438,N_16514);
and U17108 (N_17108,N_16713,N_16411);
nor U17109 (N_17109,N_16689,N_16777);
and U17110 (N_17110,N_16423,N_16724);
nand U17111 (N_17111,N_16773,N_16751);
nor U17112 (N_17112,N_16485,N_16691);
nor U17113 (N_17113,N_16790,N_16466);
xor U17114 (N_17114,N_16612,N_16403);
nor U17115 (N_17115,N_16622,N_16794);
nor U17116 (N_17116,N_16677,N_16570);
xor U17117 (N_17117,N_16756,N_16686);
nand U17118 (N_17118,N_16447,N_16721);
or U17119 (N_17119,N_16579,N_16794);
or U17120 (N_17120,N_16717,N_16462);
nand U17121 (N_17121,N_16485,N_16455);
xnor U17122 (N_17122,N_16760,N_16638);
and U17123 (N_17123,N_16664,N_16636);
xor U17124 (N_17124,N_16698,N_16705);
nand U17125 (N_17125,N_16502,N_16521);
nand U17126 (N_17126,N_16638,N_16619);
and U17127 (N_17127,N_16652,N_16539);
or U17128 (N_17128,N_16669,N_16602);
and U17129 (N_17129,N_16676,N_16528);
or U17130 (N_17130,N_16684,N_16424);
nand U17131 (N_17131,N_16770,N_16429);
xnor U17132 (N_17132,N_16767,N_16550);
nand U17133 (N_17133,N_16610,N_16519);
and U17134 (N_17134,N_16525,N_16670);
xor U17135 (N_17135,N_16756,N_16434);
xnor U17136 (N_17136,N_16621,N_16465);
and U17137 (N_17137,N_16684,N_16488);
and U17138 (N_17138,N_16544,N_16651);
nor U17139 (N_17139,N_16588,N_16546);
xnor U17140 (N_17140,N_16735,N_16631);
or U17141 (N_17141,N_16626,N_16534);
nor U17142 (N_17142,N_16667,N_16666);
and U17143 (N_17143,N_16786,N_16572);
xnor U17144 (N_17144,N_16415,N_16684);
nor U17145 (N_17145,N_16684,N_16588);
and U17146 (N_17146,N_16667,N_16429);
xor U17147 (N_17147,N_16725,N_16422);
nand U17148 (N_17148,N_16778,N_16651);
xor U17149 (N_17149,N_16479,N_16783);
or U17150 (N_17150,N_16699,N_16443);
nor U17151 (N_17151,N_16425,N_16700);
nand U17152 (N_17152,N_16573,N_16576);
or U17153 (N_17153,N_16769,N_16410);
and U17154 (N_17154,N_16788,N_16648);
nand U17155 (N_17155,N_16653,N_16551);
and U17156 (N_17156,N_16465,N_16535);
nand U17157 (N_17157,N_16534,N_16540);
nor U17158 (N_17158,N_16770,N_16430);
xor U17159 (N_17159,N_16754,N_16611);
nor U17160 (N_17160,N_16738,N_16695);
xnor U17161 (N_17161,N_16590,N_16476);
nor U17162 (N_17162,N_16438,N_16716);
xor U17163 (N_17163,N_16583,N_16550);
or U17164 (N_17164,N_16760,N_16515);
or U17165 (N_17165,N_16786,N_16495);
or U17166 (N_17166,N_16673,N_16689);
nand U17167 (N_17167,N_16748,N_16505);
nor U17168 (N_17168,N_16674,N_16408);
or U17169 (N_17169,N_16683,N_16461);
xor U17170 (N_17170,N_16423,N_16527);
or U17171 (N_17171,N_16783,N_16511);
nor U17172 (N_17172,N_16773,N_16679);
and U17173 (N_17173,N_16430,N_16449);
or U17174 (N_17174,N_16738,N_16524);
or U17175 (N_17175,N_16407,N_16419);
and U17176 (N_17176,N_16533,N_16655);
nor U17177 (N_17177,N_16703,N_16662);
nor U17178 (N_17178,N_16415,N_16544);
nor U17179 (N_17179,N_16480,N_16485);
and U17180 (N_17180,N_16495,N_16504);
xnor U17181 (N_17181,N_16606,N_16550);
xor U17182 (N_17182,N_16624,N_16598);
nor U17183 (N_17183,N_16455,N_16484);
or U17184 (N_17184,N_16572,N_16466);
xnor U17185 (N_17185,N_16721,N_16782);
nor U17186 (N_17186,N_16797,N_16546);
or U17187 (N_17187,N_16479,N_16454);
xor U17188 (N_17188,N_16790,N_16586);
or U17189 (N_17189,N_16787,N_16430);
or U17190 (N_17190,N_16525,N_16545);
nor U17191 (N_17191,N_16739,N_16501);
nand U17192 (N_17192,N_16606,N_16598);
nor U17193 (N_17193,N_16756,N_16456);
nor U17194 (N_17194,N_16495,N_16733);
or U17195 (N_17195,N_16519,N_16798);
xor U17196 (N_17196,N_16741,N_16464);
and U17197 (N_17197,N_16447,N_16622);
nor U17198 (N_17198,N_16506,N_16504);
or U17199 (N_17199,N_16759,N_16456);
or U17200 (N_17200,N_17161,N_17128);
and U17201 (N_17201,N_16820,N_17007);
xor U17202 (N_17202,N_16806,N_16929);
nand U17203 (N_17203,N_17137,N_17092);
or U17204 (N_17204,N_16944,N_16976);
nor U17205 (N_17205,N_17018,N_17168);
nor U17206 (N_17206,N_16932,N_17165);
xor U17207 (N_17207,N_16936,N_16913);
nor U17208 (N_17208,N_17117,N_16873);
xnor U17209 (N_17209,N_16895,N_17043);
xnor U17210 (N_17210,N_16979,N_17016);
xnor U17211 (N_17211,N_16974,N_16961);
nand U17212 (N_17212,N_17170,N_17179);
or U17213 (N_17213,N_17021,N_17014);
nand U17214 (N_17214,N_16856,N_16993);
and U17215 (N_17215,N_17143,N_16811);
or U17216 (N_17216,N_16845,N_17035);
or U17217 (N_17217,N_17140,N_16835);
and U17218 (N_17218,N_17011,N_17139);
xnor U17219 (N_17219,N_17039,N_17191);
nor U17220 (N_17220,N_17041,N_16824);
or U17221 (N_17221,N_17006,N_16855);
or U17222 (N_17222,N_17138,N_17122);
or U17223 (N_17223,N_17188,N_16848);
and U17224 (N_17224,N_17129,N_16916);
xor U17225 (N_17225,N_17163,N_17031);
and U17226 (N_17226,N_17113,N_16902);
and U17227 (N_17227,N_17005,N_16962);
nor U17228 (N_17228,N_16963,N_16868);
nor U17229 (N_17229,N_16886,N_16928);
nand U17230 (N_17230,N_17083,N_17156);
and U17231 (N_17231,N_16870,N_17193);
and U17232 (N_17232,N_17030,N_17104);
or U17233 (N_17233,N_17105,N_17114);
and U17234 (N_17234,N_16947,N_17171);
xor U17235 (N_17235,N_17094,N_17025);
and U17236 (N_17236,N_17065,N_16818);
or U17237 (N_17237,N_17093,N_17123);
or U17238 (N_17238,N_17084,N_16851);
and U17239 (N_17239,N_16866,N_16849);
and U17240 (N_17240,N_17075,N_17009);
nand U17241 (N_17241,N_17125,N_16987);
xor U17242 (N_17242,N_17149,N_17101);
nor U17243 (N_17243,N_17108,N_16900);
and U17244 (N_17244,N_17133,N_16903);
nand U17245 (N_17245,N_17056,N_16893);
xnor U17246 (N_17246,N_17106,N_16803);
xor U17247 (N_17247,N_17098,N_16949);
nor U17248 (N_17248,N_16834,N_17173);
nor U17249 (N_17249,N_16800,N_17130);
xor U17250 (N_17250,N_17053,N_16844);
or U17251 (N_17251,N_17144,N_17012);
xor U17252 (N_17252,N_16983,N_16846);
xor U17253 (N_17253,N_17126,N_16807);
and U17254 (N_17254,N_16920,N_16842);
xnor U17255 (N_17255,N_17028,N_16897);
or U17256 (N_17256,N_16970,N_17184);
xnor U17257 (N_17257,N_16841,N_16812);
and U17258 (N_17258,N_16881,N_17196);
and U17259 (N_17259,N_17090,N_17008);
or U17260 (N_17260,N_17095,N_16859);
nor U17261 (N_17261,N_16911,N_16805);
and U17262 (N_17262,N_16830,N_17097);
or U17263 (N_17263,N_16864,N_17153);
or U17264 (N_17264,N_16925,N_17112);
nor U17265 (N_17265,N_16819,N_16907);
nand U17266 (N_17266,N_16892,N_16843);
nand U17267 (N_17267,N_17077,N_16879);
or U17268 (N_17268,N_17058,N_16998);
xor U17269 (N_17269,N_17116,N_16831);
nor U17270 (N_17270,N_16852,N_17109);
xnor U17271 (N_17271,N_16858,N_17175);
xnor U17272 (N_17272,N_17051,N_16999);
and U17273 (N_17273,N_17004,N_16923);
and U17274 (N_17274,N_16939,N_17029);
or U17275 (N_17275,N_16853,N_17087);
and U17276 (N_17276,N_16874,N_17054);
or U17277 (N_17277,N_16869,N_16991);
xnor U17278 (N_17278,N_17189,N_16816);
and U17279 (N_17279,N_17042,N_16954);
nor U17280 (N_17280,N_16885,N_16808);
xor U17281 (N_17281,N_17024,N_16880);
and U17282 (N_17282,N_17060,N_17038);
nor U17283 (N_17283,N_17145,N_17180);
nor U17284 (N_17284,N_16933,N_17048);
nor U17285 (N_17285,N_16942,N_16978);
and U17286 (N_17286,N_16876,N_16964);
nor U17287 (N_17287,N_17176,N_17010);
nor U17288 (N_17288,N_16931,N_16956);
or U17289 (N_17289,N_16965,N_17096);
nand U17290 (N_17290,N_16995,N_16969);
and U17291 (N_17291,N_17119,N_17071);
nor U17292 (N_17292,N_16989,N_17107);
nand U17293 (N_17293,N_16912,N_17082);
nor U17294 (N_17294,N_17121,N_16814);
nand U17295 (N_17295,N_17019,N_17147);
or U17296 (N_17296,N_16982,N_16822);
nand U17297 (N_17297,N_16810,N_17000);
xnor U17298 (N_17298,N_17072,N_16952);
xnor U17299 (N_17299,N_17037,N_17169);
nand U17300 (N_17300,N_16914,N_16966);
nand U17301 (N_17301,N_16972,N_17111);
and U17302 (N_17302,N_16959,N_16943);
nor U17303 (N_17303,N_17044,N_17124);
nand U17304 (N_17304,N_16909,N_17194);
and U17305 (N_17305,N_16825,N_17167);
nor U17306 (N_17306,N_16817,N_16935);
xor U17307 (N_17307,N_17036,N_17131);
or U17308 (N_17308,N_17059,N_17057);
nand U17309 (N_17309,N_17192,N_16891);
nor U17310 (N_17310,N_16804,N_17183);
nor U17311 (N_17311,N_17164,N_17066);
nand U17312 (N_17312,N_17034,N_17063);
nor U17313 (N_17313,N_17148,N_17089);
and U17314 (N_17314,N_16945,N_17052);
nand U17315 (N_17315,N_16847,N_16850);
and U17316 (N_17316,N_16941,N_17085);
nor U17317 (N_17317,N_16973,N_17067);
or U17318 (N_17318,N_17182,N_16986);
or U17319 (N_17319,N_16996,N_16890);
nand U17320 (N_17320,N_17046,N_17103);
and U17321 (N_17321,N_17199,N_16938);
or U17322 (N_17322,N_16946,N_16829);
nor U17323 (N_17323,N_17154,N_16927);
and U17324 (N_17324,N_17178,N_16905);
nor U17325 (N_17325,N_16930,N_16968);
or U17326 (N_17326,N_16827,N_17190);
xor U17327 (N_17327,N_16865,N_17186);
nor U17328 (N_17328,N_16839,N_17015);
nand U17329 (N_17329,N_17002,N_16937);
or U17330 (N_17330,N_16984,N_17146);
xnor U17331 (N_17331,N_17166,N_17068);
and U17332 (N_17332,N_17088,N_16823);
xor U17333 (N_17333,N_16918,N_17079);
or U17334 (N_17334,N_16860,N_16826);
or U17335 (N_17335,N_16813,N_16828);
nor U17336 (N_17336,N_16884,N_17078);
or U17337 (N_17337,N_17158,N_16971);
or U17338 (N_17338,N_17141,N_16904);
nand U17339 (N_17339,N_17181,N_17074);
xor U17340 (N_17340,N_17073,N_16955);
and U17341 (N_17341,N_16940,N_17135);
nor U17342 (N_17342,N_16901,N_17050);
xor U17343 (N_17343,N_16926,N_16980);
xor U17344 (N_17344,N_16888,N_17160);
and U17345 (N_17345,N_16836,N_17003);
or U17346 (N_17346,N_17159,N_17155);
and U17347 (N_17347,N_17120,N_16896);
nand U17348 (N_17348,N_17150,N_16882);
nand U17349 (N_17349,N_17127,N_17080);
xnor U17350 (N_17350,N_17152,N_16833);
or U17351 (N_17351,N_17023,N_16840);
xor U17352 (N_17352,N_17157,N_17064);
nand U17353 (N_17353,N_16917,N_17061);
nor U17354 (N_17354,N_16953,N_16908);
nor U17355 (N_17355,N_16915,N_16867);
and U17356 (N_17356,N_16988,N_17055);
nand U17357 (N_17357,N_17047,N_16994);
nor U17358 (N_17358,N_16877,N_17091);
xnor U17359 (N_17359,N_17017,N_16815);
xor U17360 (N_17360,N_16906,N_16861);
and U17361 (N_17361,N_16821,N_16863);
nand U17362 (N_17362,N_16957,N_16894);
nand U17363 (N_17363,N_17197,N_16922);
and U17364 (N_17364,N_17045,N_17177);
nand U17365 (N_17365,N_17100,N_17026);
xor U17366 (N_17366,N_16958,N_16883);
nor U17367 (N_17367,N_16948,N_17110);
or U17368 (N_17368,N_17198,N_16977);
nor U17369 (N_17369,N_16862,N_17086);
xnor U17370 (N_17370,N_17102,N_16898);
and U17371 (N_17371,N_17032,N_16838);
or U17372 (N_17372,N_16924,N_17001);
nand U17373 (N_17373,N_17027,N_17081);
xor U17374 (N_17374,N_16878,N_16919);
and U17375 (N_17375,N_16802,N_17195);
and U17376 (N_17376,N_17136,N_16910);
xor U17377 (N_17377,N_17115,N_17033);
and U17378 (N_17378,N_16967,N_17076);
nor U17379 (N_17379,N_17099,N_16997);
nand U17380 (N_17380,N_16875,N_17022);
or U17381 (N_17381,N_16857,N_17132);
nor U17382 (N_17382,N_16951,N_16934);
xnor U17383 (N_17383,N_16981,N_16899);
nor U17384 (N_17384,N_16801,N_17185);
or U17385 (N_17385,N_17062,N_16990);
nand U17386 (N_17386,N_17013,N_16832);
or U17387 (N_17387,N_17172,N_16985);
or U17388 (N_17388,N_16992,N_16854);
or U17389 (N_17389,N_17049,N_17134);
nor U17390 (N_17390,N_17187,N_16872);
xor U17391 (N_17391,N_16887,N_16921);
and U17392 (N_17392,N_17069,N_16837);
and U17393 (N_17393,N_17151,N_17040);
nand U17394 (N_17394,N_17162,N_16809);
xor U17395 (N_17395,N_16889,N_16960);
or U17396 (N_17396,N_17118,N_17174);
xor U17397 (N_17397,N_17070,N_16871);
or U17398 (N_17398,N_16950,N_17142);
nand U17399 (N_17399,N_17020,N_16975);
nor U17400 (N_17400,N_17023,N_17031);
nand U17401 (N_17401,N_17049,N_17011);
nor U17402 (N_17402,N_16875,N_17124);
nand U17403 (N_17403,N_17079,N_16851);
nand U17404 (N_17404,N_16903,N_17022);
and U17405 (N_17405,N_17023,N_17005);
and U17406 (N_17406,N_16974,N_16831);
nor U17407 (N_17407,N_17015,N_17168);
nor U17408 (N_17408,N_16849,N_17148);
and U17409 (N_17409,N_16959,N_17082);
or U17410 (N_17410,N_17022,N_16906);
or U17411 (N_17411,N_16854,N_17176);
xnor U17412 (N_17412,N_16971,N_17157);
and U17413 (N_17413,N_17182,N_17051);
nor U17414 (N_17414,N_16833,N_17003);
xnor U17415 (N_17415,N_16866,N_16969);
and U17416 (N_17416,N_17073,N_17050);
nand U17417 (N_17417,N_16944,N_16883);
xor U17418 (N_17418,N_16864,N_16888);
and U17419 (N_17419,N_17129,N_17065);
nor U17420 (N_17420,N_17040,N_16989);
and U17421 (N_17421,N_17023,N_17166);
nand U17422 (N_17422,N_17165,N_16815);
xor U17423 (N_17423,N_16932,N_16940);
or U17424 (N_17424,N_17146,N_16947);
xor U17425 (N_17425,N_16952,N_16849);
or U17426 (N_17426,N_17197,N_17196);
nand U17427 (N_17427,N_16837,N_17189);
and U17428 (N_17428,N_16911,N_17083);
nor U17429 (N_17429,N_16834,N_16869);
nand U17430 (N_17430,N_16934,N_16851);
xor U17431 (N_17431,N_16919,N_16938);
xor U17432 (N_17432,N_16975,N_17149);
xnor U17433 (N_17433,N_17153,N_17118);
or U17434 (N_17434,N_17081,N_17163);
or U17435 (N_17435,N_17107,N_17070);
nand U17436 (N_17436,N_16813,N_17179);
xor U17437 (N_17437,N_16805,N_16900);
xnor U17438 (N_17438,N_16809,N_16930);
nor U17439 (N_17439,N_16806,N_17042);
and U17440 (N_17440,N_16934,N_16917);
and U17441 (N_17441,N_17085,N_16943);
xnor U17442 (N_17442,N_16928,N_16812);
nand U17443 (N_17443,N_16958,N_16964);
and U17444 (N_17444,N_17124,N_17198);
and U17445 (N_17445,N_16911,N_16900);
xor U17446 (N_17446,N_17096,N_16941);
nor U17447 (N_17447,N_17036,N_16885);
nor U17448 (N_17448,N_17033,N_16800);
or U17449 (N_17449,N_16886,N_17092);
nor U17450 (N_17450,N_16872,N_16842);
nand U17451 (N_17451,N_16835,N_17180);
xor U17452 (N_17452,N_17192,N_17058);
xor U17453 (N_17453,N_16930,N_16995);
nand U17454 (N_17454,N_16935,N_16973);
xnor U17455 (N_17455,N_17039,N_16898);
and U17456 (N_17456,N_17162,N_17169);
or U17457 (N_17457,N_17167,N_17012);
xnor U17458 (N_17458,N_16814,N_17100);
or U17459 (N_17459,N_16959,N_17047);
xnor U17460 (N_17460,N_16988,N_16804);
nand U17461 (N_17461,N_17085,N_16881);
and U17462 (N_17462,N_16976,N_16801);
xor U17463 (N_17463,N_16833,N_17110);
and U17464 (N_17464,N_16848,N_16974);
nand U17465 (N_17465,N_17092,N_17120);
nand U17466 (N_17466,N_16976,N_17188);
and U17467 (N_17467,N_17036,N_16956);
xnor U17468 (N_17468,N_17104,N_16888);
nor U17469 (N_17469,N_16816,N_16930);
nor U17470 (N_17470,N_16926,N_16858);
or U17471 (N_17471,N_16936,N_17103);
xor U17472 (N_17472,N_17138,N_17019);
nand U17473 (N_17473,N_16918,N_17006);
and U17474 (N_17474,N_17041,N_17070);
nor U17475 (N_17475,N_16881,N_17027);
nor U17476 (N_17476,N_17161,N_17069);
or U17477 (N_17477,N_16985,N_17161);
nor U17478 (N_17478,N_16832,N_16838);
or U17479 (N_17479,N_17103,N_17165);
xor U17480 (N_17480,N_17049,N_16930);
and U17481 (N_17481,N_16966,N_16834);
and U17482 (N_17482,N_16918,N_17139);
xnor U17483 (N_17483,N_16911,N_16893);
nor U17484 (N_17484,N_17090,N_16822);
and U17485 (N_17485,N_17126,N_17085);
xnor U17486 (N_17486,N_17041,N_16917);
and U17487 (N_17487,N_16964,N_16869);
nand U17488 (N_17488,N_17122,N_17195);
and U17489 (N_17489,N_17013,N_16993);
or U17490 (N_17490,N_17100,N_16908);
or U17491 (N_17491,N_17042,N_16868);
nand U17492 (N_17492,N_16995,N_17058);
xnor U17493 (N_17493,N_16939,N_16948);
nand U17494 (N_17494,N_16812,N_16879);
or U17495 (N_17495,N_17147,N_16809);
nand U17496 (N_17496,N_16824,N_17031);
and U17497 (N_17497,N_16808,N_17081);
or U17498 (N_17498,N_17094,N_16928);
or U17499 (N_17499,N_16916,N_17018);
xnor U17500 (N_17500,N_16864,N_16869);
nand U17501 (N_17501,N_16887,N_17118);
or U17502 (N_17502,N_16868,N_16978);
nor U17503 (N_17503,N_17163,N_17065);
xnor U17504 (N_17504,N_16836,N_16908);
xor U17505 (N_17505,N_16891,N_17013);
nor U17506 (N_17506,N_16972,N_17139);
xnor U17507 (N_17507,N_16907,N_17105);
or U17508 (N_17508,N_16909,N_17017);
xor U17509 (N_17509,N_16924,N_16846);
xor U17510 (N_17510,N_16872,N_17084);
nand U17511 (N_17511,N_17099,N_17089);
and U17512 (N_17512,N_16959,N_16992);
xor U17513 (N_17513,N_16970,N_16904);
nand U17514 (N_17514,N_16846,N_16814);
xnor U17515 (N_17515,N_16835,N_16844);
and U17516 (N_17516,N_16932,N_17162);
nor U17517 (N_17517,N_17102,N_17077);
nand U17518 (N_17518,N_16992,N_16906);
nor U17519 (N_17519,N_16808,N_17075);
and U17520 (N_17520,N_17178,N_16945);
or U17521 (N_17521,N_16916,N_16971);
nand U17522 (N_17522,N_17194,N_17062);
nor U17523 (N_17523,N_16965,N_16976);
xnor U17524 (N_17524,N_17164,N_17173);
nand U17525 (N_17525,N_17177,N_17144);
or U17526 (N_17526,N_17177,N_17150);
or U17527 (N_17527,N_16972,N_16876);
and U17528 (N_17528,N_16840,N_16843);
or U17529 (N_17529,N_17057,N_16902);
or U17530 (N_17530,N_17174,N_17108);
nand U17531 (N_17531,N_17004,N_16849);
nor U17532 (N_17532,N_16911,N_16941);
xnor U17533 (N_17533,N_16897,N_16899);
nor U17534 (N_17534,N_16908,N_16839);
or U17535 (N_17535,N_17088,N_17059);
and U17536 (N_17536,N_17186,N_17035);
nor U17537 (N_17537,N_16826,N_17067);
and U17538 (N_17538,N_16822,N_16867);
xor U17539 (N_17539,N_17192,N_16900);
nor U17540 (N_17540,N_17050,N_16976);
or U17541 (N_17541,N_17149,N_16930);
nor U17542 (N_17542,N_16965,N_17122);
nor U17543 (N_17543,N_17047,N_17095);
nor U17544 (N_17544,N_17142,N_17116);
and U17545 (N_17545,N_16996,N_16926);
nand U17546 (N_17546,N_17180,N_17130);
xnor U17547 (N_17547,N_16976,N_16839);
nor U17548 (N_17548,N_16879,N_16889);
nor U17549 (N_17549,N_16853,N_16802);
and U17550 (N_17550,N_16886,N_16941);
xor U17551 (N_17551,N_16911,N_16955);
nand U17552 (N_17552,N_17020,N_17170);
and U17553 (N_17553,N_16805,N_16872);
nand U17554 (N_17554,N_16829,N_17063);
or U17555 (N_17555,N_16944,N_16826);
or U17556 (N_17556,N_16958,N_16909);
xnor U17557 (N_17557,N_16974,N_16937);
and U17558 (N_17558,N_17136,N_16940);
xnor U17559 (N_17559,N_17005,N_16822);
or U17560 (N_17560,N_17041,N_16946);
and U17561 (N_17561,N_17089,N_17075);
and U17562 (N_17562,N_17049,N_16984);
and U17563 (N_17563,N_17047,N_17024);
nand U17564 (N_17564,N_17065,N_16910);
xnor U17565 (N_17565,N_16813,N_17149);
nand U17566 (N_17566,N_16819,N_16805);
nor U17567 (N_17567,N_16978,N_17051);
nor U17568 (N_17568,N_16895,N_16840);
or U17569 (N_17569,N_16963,N_17032);
and U17570 (N_17570,N_16824,N_17007);
xor U17571 (N_17571,N_16907,N_17176);
and U17572 (N_17572,N_17016,N_16859);
and U17573 (N_17573,N_17161,N_17045);
nor U17574 (N_17574,N_16961,N_16999);
nor U17575 (N_17575,N_16886,N_16852);
nand U17576 (N_17576,N_16881,N_17187);
nand U17577 (N_17577,N_16920,N_16868);
or U17578 (N_17578,N_16851,N_17081);
nor U17579 (N_17579,N_17005,N_17060);
and U17580 (N_17580,N_16911,N_17166);
or U17581 (N_17581,N_17035,N_16914);
nor U17582 (N_17582,N_17112,N_16934);
nor U17583 (N_17583,N_16840,N_17055);
and U17584 (N_17584,N_17024,N_16801);
nand U17585 (N_17585,N_16810,N_17107);
and U17586 (N_17586,N_16931,N_16970);
and U17587 (N_17587,N_17102,N_16985);
xnor U17588 (N_17588,N_17146,N_17017);
xnor U17589 (N_17589,N_17186,N_16807);
and U17590 (N_17590,N_17169,N_16923);
xnor U17591 (N_17591,N_16940,N_17172);
or U17592 (N_17592,N_16911,N_17175);
nand U17593 (N_17593,N_16884,N_16824);
xor U17594 (N_17594,N_16871,N_16975);
and U17595 (N_17595,N_16888,N_17050);
and U17596 (N_17596,N_17079,N_17008);
or U17597 (N_17597,N_17009,N_17177);
nand U17598 (N_17598,N_17068,N_17167);
or U17599 (N_17599,N_16971,N_16872);
and U17600 (N_17600,N_17525,N_17258);
nor U17601 (N_17601,N_17243,N_17387);
xor U17602 (N_17602,N_17323,N_17331);
xor U17603 (N_17603,N_17244,N_17463);
nand U17604 (N_17604,N_17529,N_17499);
and U17605 (N_17605,N_17375,N_17496);
xnor U17606 (N_17606,N_17272,N_17543);
nor U17607 (N_17607,N_17384,N_17536);
xor U17608 (N_17608,N_17478,N_17549);
nand U17609 (N_17609,N_17462,N_17203);
nand U17610 (N_17610,N_17268,N_17237);
xnor U17611 (N_17611,N_17240,N_17520);
or U17612 (N_17612,N_17297,N_17298);
nand U17613 (N_17613,N_17363,N_17382);
nand U17614 (N_17614,N_17381,N_17226);
nor U17615 (N_17615,N_17311,N_17353);
nor U17616 (N_17616,N_17335,N_17236);
or U17617 (N_17617,N_17424,N_17595);
xor U17618 (N_17618,N_17523,N_17285);
nand U17619 (N_17619,N_17430,N_17339);
xnor U17620 (N_17620,N_17429,N_17326);
xor U17621 (N_17621,N_17581,N_17325);
xor U17622 (N_17622,N_17474,N_17421);
and U17623 (N_17623,N_17577,N_17359);
and U17624 (N_17624,N_17368,N_17344);
and U17625 (N_17625,N_17567,N_17234);
nand U17626 (N_17626,N_17396,N_17253);
nand U17627 (N_17627,N_17211,N_17231);
nor U17628 (N_17628,N_17510,N_17437);
xnor U17629 (N_17629,N_17400,N_17535);
nand U17630 (N_17630,N_17470,N_17342);
nand U17631 (N_17631,N_17449,N_17241);
and U17632 (N_17632,N_17334,N_17455);
xor U17633 (N_17633,N_17447,N_17544);
or U17634 (N_17634,N_17362,N_17355);
xor U17635 (N_17635,N_17386,N_17218);
and U17636 (N_17636,N_17318,N_17440);
or U17637 (N_17637,N_17521,N_17419);
xor U17638 (N_17638,N_17372,N_17300);
nor U17639 (N_17639,N_17327,N_17371);
nor U17640 (N_17640,N_17502,N_17225);
xnor U17641 (N_17641,N_17286,N_17201);
nor U17642 (N_17642,N_17385,N_17330);
xnor U17643 (N_17643,N_17484,N_17338);
nand U17644 (N_17644,N_17566,N_17279);
and U17645 (N_17645,N_17505,N_17433);
or U17646 (N_17646,N_17369,N_17441);
or U17647 (N_17647,N_17235,N_17345);
nand U17648 (N_17648,N_17533,N_17217);
or U17649 (N_17649,N_17545,N_17263);
and U17650 (N_17650,N_17580,N_17299);
nand U17651 (N_17651,N_17402,N_17585);
xor U17652 (N_17652,N_17420,N_17598);
nor U17653 (N_17653,N_17374,N_17264);
and U17654 (N_17654,N_17360,N_17219);
xnor U17655 (N_17655,N_17357,N_17262);
nor U17656 (N_17656,N_17404,N_17464);
or U17657 (N_17657,N_17426,N_17354);
nand U17658 (N_17658,N_17341,N_17316);
nor U17659 (N_17659,N_17251,N_17548);
xor U17660 (N_17660,N_17207,N_17451);
nand U17661 (N_17661,N_17432,N_17352);
xor U17662 (N_17662,N_17442,N_17295);
and U17663 (N_17663,N_17301,N_17278);
nor U17664 (N_17664,N_17337,N_17412);
or U17665 (N_17665,N_17434,N_17305);
nor U17666 (N_17666,N_17541,N_17356);
nor U17667 (N_17667,N_17489,N_17568);
xnor U17668 (N_17668,N_17348,N_17347);
xor U17669 (N_17669,N_17200,N_17438);
xor U17670 (N_17670,N_17229,N_17423);
nor U17671 (N_17671,N_17560,N_17389);
xnor U17672 (N_17672,N_17376,N_17303);
or U17673 (N_17673,N_17287,N_17469);
nor U17674 (N_17674,N_17427,N_17254);
nor U17675 (N_17675,N_17212,N_17572);
nor U17676 (N_17676,N_17488,N_17480);
nand U17677 (N_17677,N_17365,N_17422);
nor U17678 (N_17678,N_17216,N_17313);
nor U17679 (N_17679,N_17343,N_17448);
nor U17680 (N_17680,N_17494,N_17340);
nand U17681 (N_17681,N_17519,N_17565);
nand U17682 (N_17682,N_17271,N_17500);
nand U17683 (N_17683,N_17370,N_17594);
nor U17684 (N_17684,N_17332,N_17582);
or U17685 (N_17685,N_17573,N_17406);
nand U17686 (N_17686,N_17399,N_17576);
xor U17687 (N_17687,N_17288,N_17466);
xnor U17688 (N_17688,N_17329,N_17485);
nor U17689 (N_17689,N_17592,N_17537);
or U17690 (N_17690,N_17373,N_17579);
or U17691 (N_17691,N_17491,N_17249);
or U17692 (N_17692,N_17558,N_17516);
xor U17693 (N_17693,N_17569,N_17208);
nand U17694 (N_17694,N_17364,N_17407);
and U17695 (N_17695,N_17564,N_17250);
nor U17696 (N_17696,N_17597,N_17482);
nand U17697 (N_17697,N_17479,N_17380);
nand U17698 (N_17698,N_17508,N_17498);
xor U17699 (N_17699,N_17350,N_17293);
nor U17700 (N_17700,N_17450,N_17290);
xor U17701 (N_17701,N_17457,N_17459);
or U17702 (N_17702,N_17314,N_17409);
xnor U17703 (N_17703,N_17307,N_17501);
xor U17704 (N_17704,N_17490,N_17524);
and U17705 (N_17705,N_17248,N_17439);
or U17706 (N_17706,N_17443,N_17528);
nand U17707 (N_17707,N_17532,N_17550);
nor U17708 (N_17708,N_17454,N_17283);
nand U17709 (N_17709,N_17214,N_17487);
nand U17710 (N_17710,N_17559,N_17265);
and U17711 (N_17711,N_17242,N_17260);
or U17712 (N_17712,N_17276,N_17238);
or U17713 (N_17713,N_17435,N_17493);
or U17714 (N_17714,N_17289,N_17274);
or U17715 (N_17715,N_17509,N_17252);
xor U17716 (N_17716,N_17492,N_17591);
xor U17717 (N_17717,N_17257,N_17551);
nand U17718 (N_17718,N_17408,N_17280);
or U17719 (N_17719,N_17539,N_17391);
and U17720 (N_17720,N_17306,N_17518);
xor U17721 (N_17721,N_17220,N_17570);
xnor U17722 (N_17722,N_17465,N_17224);
and U17723 (N_17723,N_17270,N_17593);
nand U17724 (N_17724,N_17379,N_17590);
nand U17725 (N_17725,N_17294,N_17552);
and U17726 (N_17726,N_17351,N_17273);
nor U17727 (N_17727,N_17296,N_17246);
xor U17728 (N_17728,N_17497,N_17481);
and U17729 (N_17729,N_17383,N_17452);
xnor U17730 (N_17730,N_17205,N_17349);
nand U17731 (N_17731,N_17336,N_17247);
and U17732 (N_17732,N_17284,N_17410);
or U17733 (N_17733,N_17308,N_17575);
or U17734 (N_17734,N_17392,N_17514);
nand U17735 (N_17735,N_17227,N_17504);
nor U17736 (N_17736,N_17534,N_17328);
xnor U17737 (N_17737,N_17589,N_17390);
or U17738 (N_17738,N_17553,N_17411);
and U17739 (N_17739,N_17259,N_17425);
xor U17740 (N_17740,N_17586,N_17315);
nand U17741 (N_17741,N_17292,N_17506);
nand U17742 (N_17742,N_17267,N_17394);
nor U17743 (N_17743,N_17239,N_17403);
or U17744 (N_17744,N_17233,N_17277);
or U17745 (N_17745,N_17495,N_17511);
or U17746 (N_17746,N_17230,N_17310);
or U17747 (N_17747,N_17414,N_17358);
nor U17748 (N_17748,N_17255,N_17312);
xor U17749 (N_17749,N_17599,N_17486);
or U17750 (N_17750,N_17526,N_17460);
and U17751 (N_17751,N_17324,N_17269);
and U17752 (N_17752,N_17477,N_17527);
nor U17753 (N_17753,N_17282,N_17538);
and U17754 (N_17754,N_17317,N_17587);
nand U17755 (N_17755,N_17291,N_17503);
or U17756 (N_17756,N_17461,N_17377);
xor U17757 (N_17757,N_17322,N_17221);
xor U17758 (N_17758,N_17563,N_17446);
or U17759 (N_17759,N_17388,N_17513);
or U17760 (N_17760,N_17418,N_17584);
or U17761 (N_17761,N_17522,N_17395);
nor U17762 (N_17762,N_17431,N_17204);
and U17763 (N_17763,N_17578,N_17215);
or U17764 (N_17764,N_17476,N_17417);
nand U17765 (N_17765,N_17393,N_17401);
or U17766 (N_17766,N_17574,N_17596);
or U17767 (N_17767,N_17547,N_17398);
or U17768 (N_17768,N_17228,N_17453);
or U17769 (N_17769,N_17542,N_17320);
nor U17770 (N_17770,N_17266,N_17361);
or U17771 (N_17771,N_17472,N_17309);
and U17772 (N_17772,N_17571,N_17468);
nand U17773 (N_17773,N_17213,N_17232);
or U17774 (N_17774,N_17531,N_17475);
xor U17775 (N_17775,N_17557,N_17554);
nor U17776 (N_17776,N_17588,N_17405);
nor U17777 (N_17777,N_17321,N_17378);
nand U17778 (N_17778,N_17397,N_17556);
nor U17779 (N_17779,N_17562,N_17415);
xnor U17780 (N_17780,N_17333,N_17467);
nor U17781 (N_17781,N_17206,N_17456);
or U17782 (N_17782,N_17540,N_17275);
nor U17783 (N_17783,N_17202,N_17281);
nor U17784 (N_17784,N_17210,N_17223);
or U17785 (N_17785,N_17302,N_17483);
nor U17786 (N_17786,N_17471,N_17445);
nand U17787 (N_17787,N_17367,N_17583);
xor U17788 (N_17788,N_17245,N_17346);
xnor U17789 (N_17789,N_17444,N_17517);
xor U17790 (N_17790,N_17256,N_17413);
xor U17791 (N_17791,N_17304,N_17458);
nand U17792 (N_17792,N_17546,N_17209);
and U17793 (N_17793,N_17473,N_17366);
or U17794 (N_17794,N_17515,N_17561);
nand U17795 (N_17795,N_17319,N_17555);
nor U17796 (N_17796,N_17507,N_17512);
or U17797 (N_17797,N_17436,N_17428);
nor U17798 (N_17798,N_17416,N_17222);
nand U17799 (N_17799,N_17261,N_17530);
nand U17800 (N_17800,N_17297,N_17287);
nand U17801 (N_17801,N_17279,N_17556);
nor U17802 (N_17802,N_17543,N_17573);
xor U17803 (N_17803,N_17296,N_17207);
xor U17804 (N_17804,N_17278,N_17422);
and U17805 (N_17805,N_17413,N_17261);
or U17806 (N_17806,N_17538,N_17532);
nor U17807 (N_17807,N_17278,N_17264);
nor U17808 (N_17808,N_17367,N_17239);
nand U17809 (N_17809,N_17379,N_17499);
nor U17810 (N_17810,N_17299,N_17555);
xnor U17811 (N_17811,N_17458,N_17403);
xnor U17812 (N_17812,N_17349,N_17486);
xnor U17813 (N_17813,N_17566,N_17554);
nand U17814 (N_17814,N_17533,N_17447);
nor U17815 (N_17815,N_17401,N_17267);
and U17816 (N_17816,N_17571,N_17560);
xnor U17817 (N_17817,N_17486,N_17543);
nor U17818 (N_17818,N_17297,N_17508);
or U17819 (N_17819,N_17212,N_17502);
or U17820 (N_17820,N_17367,N_17439);
nand U17821 (N_17821,N_17457,N_17388);
nor U17822 (N_17822,N_17577,N_17208);
nor U17823 (N_17823,N_17247,N_17571);
xnor U17824 (N_17824,N_17526,N_17510);
or U17825 (N_17825,N_17317,N_17275);
and U17826 (N_17826,N_17478,N_17479);
nor U17827 (N_17827,N_17226,N_17457);
nor U17828 (N_17828,N_17424,N_17316);
or U17829 (N_17829,N_17559,N_17512);
and U17830 (N_17830,N_17307,N_17352);
or U17831 (N_17831,N_17343,N_17570);
or U17832 (N_17832,N_17436,N_17569);
nor U17833 (N_17833,N_17258,N_17329);
and U17834 (N_17834,N_17238,N_17509);
nor U17835 (N_17835,N_17302,N_17356);
nand U17836 (N_17836,N_17463,N_17410);
and U17837 (N_17837,N_17223,N_17415);
xnor U17838 (N_17838,N_17471,N_17409);
or U17839 (N_17839,N_17428,N_17346);
xnor U17840 (N_17840,N_17228,N_17517);
or U17841 (N_17841,N_17524,N_17343);
and U17842 (N_17842,N_17348,N_17380);
nor U17843 (N_17843,N_17524,N_17339);
xor U17844 (N_17844,N_17210,N_17435);
xor U17845 (N_17845,N_17502,N_17486);
and U17846 (N_17846,N_17320,N_17451);
nand U17847 (N_17847,N_17262,N_17211);
xnor U17848 (N_17848,N_17201,N_17493);
or U17849 (N_17849,N_17535,N_17599);
or U17850 (N_17850,N_17534,N_17593);
or U17851 (N_17851,N_17234,N_17335);
and U17852 (N_17852,N_17426,N_17556);
nand U17853 (N_17853,N_17241,N_17290);
or U17854 (N_17854,N_17336,N_17483);
xnor U17855 (N_17855,N_17379,N_17473);
and U17856 (N_17856,N_17496,N_17270);
nor U17857 (N_17857,N_17227,N_17465);
nand U17858 (N_17858,N_17488,N_17561);
nor U17859 (N_17859,N_17575,N_17249);
nand U17860 (N_17860,N_17431,N_17521);
nand U17861 (N_17861,N_17473,N_17485);
or U17862 (N_17862,N_17515,N_17288);
nor U17863 (N_17863,N_17548,N_17259);
nand U17864 (N_17864,N_17328,N_17268);
or U17865 (N_17865,N_17598,N_17337);
and U17866 (N_17866,N_17349,N_17214);
xnor U17867 (N_17867,N_17295,N_17578);
or U17868 (N_17868,N_17419,N_17423);
and U17869 (N_17869,N_17271,N_17349);
nand U17870 (N_17870,N_17513,N_17392);
and U17871 (N_17871,N_17425,N_17354);
nand U17872 (N_17872,N_17582,N_17587);
nor U17873 (N_17873,N_17534,N_17365);
nand U17874 (N_17874,N_17352,N_17472);
xor U17875 (N_17875,N_17496,N_17290);
xnor U17876 (N_17876,N_17279,N_17248);
nor U17877 (N_17877,N_17579,N_17293);
nand U17878 (N_17878,N_17335,N_17287);
xor U17879 (N_17879,N_17355,N_17369);
or U17880 (N_17880,N_17339,N_17452);
nand U17881 (N_17881,N_17566,N_17407);
nor U17882 (N_17882,N_17243,N_17247);
nor U17883 (N_17883,N_17309,N_17336);
nor U17884 (N_17884,N_17442,N_17206);
and U17885 (N_17885,N_17214,N_17395);
nand U17886 (N_17886,N_17317,N_17272);
and U17887 (N_17887,N_17460,N_17375);
xnor U17888 (N_17888,N_17441,N_17546);
nor U17889 (N_17889,N_17506,N_17306);
nand U17890 (N_17890,N_17544,N_17372);
and U17891 (N_17891,N_17577,N_17335);
nor U17892 (N_17892,N_17235,N_17290);
nand U17893 (N_17893,N_17364,N_17567);
xor U17894 (N_17894,N_17438,N_17465);
nand U17895 (N_17895,N_17450,N_17460);
or U17896 (N_17896,N_17247,N_17260);
or U17897 (N_17897,N_17429,N_17346);
and U17898 (N_17898,N_17586,N_17509);
xnor U17899 (N_17899,N_17525,N_17578);
nand U17900 (N_17900,N_17504,N_17226);
nor U17901 (N_17901,N_17333,N_17253);
nand U17902 (N_17902,N_17239,N_17410);
or U17903 (N_17903,N_17481,N_17207);
or U17904 (N_17904,N_17591,N_17310);
nor U17905 (N_17905,N_17205,N_17418);
or U17906 (N_17906,N_17336,N_17487);
or U17907 (N_17907,N_17421,N_17340);
nand U17908 (N_17908,N_17333,N_17268);
and U17909 (N_17909,N_17503,N_17584);
nor U17910 (N_17910,N_17515,N_17351);
or U17911 (N_17911,N_17434,N_17449);
or U17912 (N_17912,N_17419,N_17511);
and U17913 (N_17913,N_17427,N_17373);
and U17914 (N_17914,N_17300,N_17438);
or U17915 (N_17915,N_17425,N_17486);
nand U17916 (N_17916,N_17418,N_17276);
xnor U17917 (N_17917,N_17408,N_17483);
and U17918 (N_17918,N_17443,N_17464);
nor U17919 (N_17919,N_17281,N_17559);
xor U17920 (N_17920,N_17394,N_17406);
nor U17921 (N_17921,N_17459,N_17471);
or U17922 (N_17922,N_17354,N_17398);
or U17923 (N_17923,N_17225,N_17372);
xor U17924 (N_17924,N_17287,N_17580);
and U17925 (N_17925,N_17342,N_17491);
nand U17926 (N_17926,N_17391,N_17540);
nor U17927 (N_17927,N_17565,N_17323);
nor U17928 (N_17928,N_17538,N_17512);
nor U17929 (N_17929,N_17439,N_17539);
nand U17930 (N_17930,N_17582,N_17355);
nand U17931 (N_17931,N_17264,N_17551);
xnor U17932 (N_17932,N_17483,N_17280);
nand U17933 (N_17933,N_17459,N_17240);
nand U17934 (N_17934,N_17486,N_17548);
xnor U17935 (N_17935,N_17379,N_17422);
nand U17936 (N_17936,N_17282,N_17588);
nand U17937 (N_17937,N_17460,N_17259);
or U17938 (N_17938,N_17385,N_17220);
nand U17939 (N_17939,N_17307,N_17545);
and U17940 (N_17940,N_17449,N_17371);
and U17941 (N_17941,N_17241,N_17379);
nor U17942 (N_17942,N_17250,N_17419);
nor U17943 (N_17943,N_17394,N_17422);
or U17944 (N_17944,N_17371,N_17301);
xor U17945 (N_17945,N_17418,N_17402);
or U17946 (N_17946,N_17383,N_17406);
nand U17947 (N_17947,N_17379,N_17335);
and U17948 (N_17948,N_17483,N_17273);
and U17949 (N_17949,N_17279,N_17369);
nor U17950 (N_17950,N_17325,N_17319);
and U17951 (N_17951,N_17395,N_17246);
xnor U17952 (N_17952,N_17551,N_17364);
nand U17953 (N_17953,N_17433,N_17372);
nor U17954 (N_17954,N_17210,N_17313);
or U17955 (N_17955,N_17412,N_17462);
or U17956 (N_17956,N_17443,N_17320);
nor U17957 (N_17957,N_17413,N_17339);
and U17958 (N_17958,N_17453,N_17227);
nor U17959 (N_17959,N_17321,N_17457);
or U17960 (N_17960,N_17398,N_17242);
xnor U17961 (N_17961,N_17255,N_17396);
and U17962 (N_17962,N_17590,N_17499);
or U17963 (N_17963,N_17478,N_17313);
xor U17964 (N_17964,N_17507,N_17572);
nor U17965 (N_17965,N_17375,N_17424);
nand U17966 (N_17966,N_17591,N_17232);
nor U17967 (N_17967,N_17280,N_17490);
or U17968 (N_17968,N_17228,N_17462);
or U17969 (N_17969,N_17490,N_17555);
xor U17970 (N_17970,N_17224,N_17547);
xnor U17971 (N_17971,N_17448,N_17307);
xor U17972 (N_17972,N_17560,N_17311);
or U17973 (N_17973,N_17579,N_17557);
and U17974 (N_17974,N_17262,N_17319);
nor U17975 (N_17975,N_17223,N_17205);
nand U17976 (N_17976,N_17271,N_17223);
nand U17977 (N_17977,N_17219,N_17434);
or U17978 (N_17978,N_17552,N_17291);
nor U17979 (N_17979,N_17443,N_17408);
or U17980 (N_17980,N_17596,N_17338);
xor U17981 (N_17981,N_17444,N_17287);
and U17982 (N_17982,N_17371,N_17304);
or U17983 (N_17983,N_17532,N_17497);
or U17984 (N_17984,N_17505,N_17313);
nor U17985 (N_17985,N_17567,N_17590);
nor U17986 (N_17986,N_17264,N_17449);
xor U17987 (N_17987,N_17304,N_17494);
xnor U17988 (N_17988,N_17439,N_17382);
xor U17989 (N_17989,N_17583,N_17402);
xor U17990 (N_17990,N_17215,N_17534);
and U17991 (N_17991,N_17356,N_17305);
nor U17992 (N_17992,N_17409,N_17371);
nor U17993 (N_17993,N_17257,N_17575);
nor U17994 (N_17994,N_17567,N_17298);
nand U17995 (N_17995,N_17336,N_17359);
xor U17996 (N_17996,N_17592,N_17542);
nor U17997 (N_17997,N_17510,N_17562);
or U17998 (N_17998,N_17493,N_17208);
and U17999 (N_17999,N_17321,N_17303);
xor U18000 (N_18000,N_17776,N_17991);
xnor U18001 (N_18001,N_17648,N_17888);
nand U18002 (N_18002,N_17979,N_17716);
and U18003 (N_18003,N_17929,N_17905);
nor U18004 (N_18004,N_17824,N_17729);
nor U18005 (N_18005,N_17677,N_17971);
nand U18006 (N_18006,N_17753,N_17615);
nor U18007 (N_18007,N_17742,N_17918);
xor U18008 (N_18008,N_17965,N_17827);
nand U18009 (N_18009,N_17993,N_17895);
xor U18010 (N_18010,N_17869,N_17883);
xnor U18011 (N_18011,N_17631,N_17690);
and U18012 (N_18012,N_17823,N_17967);
nor U18013 (N_18013,N_17604,N_17860);
or U18014 (N_18014,N_17975,N_17841);
or U18015 (N_18015,N_17725,N_17878);
nand U18016 (N_18016,N_17645,N_17897);
nand U18017 (N_18017,N_17923,N_17899);
or U18018 (N_18018,N_17763,N_17986);
xor U18019 (N_18019,N_17813,N_17704);
nand U18020 (N_18020,N_17987,N_17658);
and U18021 (N_18021,N_17737,N_17885);
xor U18022 (N_18022,N_17675,N_17711);
xnor U18023 (N_18023,N_17830,N_17727);
nor U18024 (N_18024,N_17890,N_17811);
or U18025 (N_18025,N_17849,N_17721);
and U18026 (N_18026,N_17747,N_17728);
and U18027 (N_18027,N_17958,N_17980);
nor U18028 (N_18028,N_17892,N_17735);
nand U18029 (N_18029,N_17682,N_17843);
and U18030 (N_18030,N_17619,N_17853);
nor U18031 (N_18031,N_17802,N_17751);
xor U18032 (N_18032,N_17624,N_17653);
nor U18033 (N_18033,N_17616,N_17801);
xnor U18034 (N_18034,N_17950,N_17748);
nand U18035 (N_18035,N_17870,N_17997);
xnor U18036 (N_18036,N_17931,N_17695);
or U18037 (N_18037,N_17663,N_17673);
or U18038 (N_18038,N_17693,N_17768);
xnor U18039 (N_18039,N_17731,N_17854);
or U18040 (N_18040,N_17994,N_17646);
or U18041 (N_18041,N_17654,N_17844);
or U18042 (N_18042,N_17617,N_17627);
nand U18043 (N_18043,N_17710,N_17852);
xor U18044 (N_18044,N_17644,N_17746);
and U18045 (N_18045,N_17964,N_17911);
xor U18046 (N_18046,N_17800,N_17809);
nor U18047 (N_18047,N_17708,N_17679);
nand U18048 (N_18048,N_17933,N_17612);
nand U18049 (N_18049,N_17879,N_17819);
xnor U18050 (N_18050,N_17607,N_17797);
nor U18051 (N_18051,N_17699,N_17600);
and U18052 (N_18052,N_17915,N_17973);
xnor U18053 (N_18053,N_17769,N_17842);
nand U18054 (N_18054,N_17903,N_17688);
and U18055 (N_18055,N_17835,N_17686);
xor U18056 (N_18056,N_17629,N_17639);
xnor U18057 (N_18057,N_17957,N_17807);
nor U18058 (N_18058,N_17920,N_17651);
xor U18059 (N_18059,N_17745,N_17775);
or U18060 (N_18060,N_17910,N_17655);
nand U18061 (N_18061,N_17744,N_17766);
xnor U18062 (N_18062,N_17926,N_17674);
or U18063 (N_18063,N_17839,N_17714);
xnor U18064 (N_18064,N_17630,N_17762);
nor U18065 (N_18065,N_17656,N_17937);
nor U18066 (N_18066,N_17804,N_17755);
or U18067 (N_18067,N_17966,N_17738);
or U18068 (N_18068,N_17712,N_17850);
and U18069 (N_18069,N_17720,N_17988);
or U18070 (N_18070,N_17855,N_17603);
xnor U18071 (N_18071,N_17730,N_17758);
xnor U18072 (N_18072,N_17664,N_17652);
nor U18073 (N_18073,N_17628,N_17779);
or U18074 (N_18074,N_17941,N_17691);
nand U18075 (N_18075,N_17756,N_17622);
nand U18076 (N_18076,N_17798,N_17906);
and U18077 (N_18077,N_17613,N_17626);
nor U18078 (N_18078,N_17799,N_17680);
nand U18079 (N_18079,N_17930,N_17828);
nor U18080 (N_18080,N_17689,N_17947);
nor U18081 (N_18081,N_17970,N_17785);
nor U18082 (N_18082,N_17977,N_17794);
and U18083 (N_18083,N_17927,N_17700);
nor U18084 (N_18084,N_17882,N_17916);
and U18085 (N_18085,N_17900,N_17896);
xnor U18086 (N_18086,N_17732,N_17759);
and U18087 (N_18087,N_17635,N_17694);
and U18088 (N_18088,N_17998,N_17940);
and U18089 (N_18089,N_17873,N_17810);
nand U18090 (N_18090,N_17862,N_17670);
nor U18091 (N_18091,N_17938,N_17898);
or U18092 (N_18092,N_17698,N_17995);
xnor U18093 (N_18093,N_17985,N_17917);
or U18094 (N_18094,N_17960,N_17925);
nor U18095 (N_18095,N_17783,N_17601);
nor U18096 (N_18096,N_17959,N_17932);
xor U18097 (N_18097,N_17914,N_17936);
and U18098 (N_18098,N_17788,N_17750);
xor U18099 (N_18099,N_17934,N_17761);
or U18100 (N_18100,N_17924,N_17724);
xor U18101 (N_18101,N_17846,N_17790);
nor U18102 (N_18102,N_17889,N_17871);
and U18103 (N_18103,N_17868,N_17864);
and U18104 (N_18104,N_17726,N_17837);
and U18105 (N_18105,N_17713,N_17697);
or U18106 (N_18106,N_17902,N_17657);
nand U18107 (N_18107,N_17719,N_17989);
xnor U18108 (N_18108,N_17901,N_17672);
nand U18109 (N_18109,N_17954,N_17981);
nand U18110 (N_18110,N_17808,N_17687);
and U18111 (N_18111,N_17784,N_17952);
and U18112 (N_18112,N_17787,N_17661);
nor U18113 (N_18113,N_17770,N_17949);
or U18114 (N_18114,N_17962,N_17963);
or U18115 (N_18115,N_17821,N_17618);
nand U18116 (N_18116,N_17848,N_17647);
and U18117 (N_18117,N_17637,N_17845);
nand U18118 (N_18118,N_17669,N_17928);
xnor U18119 (N_18119,N_17822,N_17831);
nor U18120 (N_18120,N_17610,N_17935);
xnor U18121 (N_18121,N_17772,N_17847);
xnor U18122 (N_18122,N_17771,N_17707);
nor U18123 (N_18123,N_17706,N_17786);
nand U18124 (N_18124,N_17678,N_17741);
and U18125 (N_18125,N_17829,N_17765);
nor U18126 (N_18126,N_17815,N_17764);
xnor U18127 (N_18127,N_17715,N_17832);
nand U18128 (N_18128,N_17736,N_17881);
or U18129 (N_18129,N_17956,N_17773);
xor U18130 (N_18130,N_17705,N_17781);
and U18131 (N_18131,N_17836,N_17752);
nor U18132 (N_18132,N_17662,N_17921);
nor U18133 (N_18133,N_17817,N_17820);
or U18134 (N_18134,N_17876,N_17996);
nor U18135 (N_18135,N_17609,N_17792);
nor U18136 (N_18136,N_17945,N_17880);
nand U18137 (N_18137,N_17884,N_17733);
and U18138 (N_18138,N_17668,N_17623);
or U18139 (N_18139,N_17886,N_17757);
and U18140 (N_18140,N_17739,N_17782);
nor U18141 (N_18141,N_17702,N_17649);
nor U18142 (N_18142,N_17974,N_17803);
nand U18143 (N_18143,N_17833,N_17942);
and U18144 (N_18144,N_17907,N_17774);
xnor U18145 (N_18145,N_17806,N_17908);
xor U18146 (N_18146,N_17760,N_17717);
nor U18147 (N_18147,N_17778,N_17922);
nor U18148 (N_18148,N_17633,N_17972);
or U18149 (N_18149,N_17969,N_17812);
nand U18150 (N_18150,N_17780,N_17777);
and U18151 (N_18151,N_17632,N_17826);
xnor U18152 (N_18152,N_17789,N_17861);
xnor U18153 (N_18153,N_17961,N_17805);
and U18154 (N_18154,N_17904,N_17754);
and U18155 (N_18155,N_17866,N_17685);
xor U18156 (N_18156,N_17894,N_17865);
nor U18157 (N_18157,N_17667,N_17968);
or U18158 (N_18158,N_17703,N_17857);
and U18159 (N_18159,N_17621,N_17749);
xor U18160 (N_18160,N_17709,N_17681);
nand U18161 (N_18161,N_17978,N_17608);
nor U18162 (N_18162,N_17666,N_17740);
nor U18163 (N_18163,N_17796,N_17641);
nand U18164 (N_18164,N_17696,N_17640);
or U18165 (N_18165,N_17951,N_17891);
and U18166 (N_18166,N_17814,N_17913);
and U18167 (N_18167,N_17877,N_17909);
nor U18168 (N_18168,N_17636,N_17851);
or U18169 (N_18169,N_17944,N_17953);
and U18170 (N_18170,N_17722,N_17834);
and U18171 (N_18171,N_17943,N_17818);
and U18172 (N_18172,N_17718,N_17791);
xnor U18173 (N_18173,N_17692,N_17955);
or U18174 (N_18174,N_17665,N_17867);
and U18175 (N_18175,N_17684,N_17838);
nand U18176 (N_18176,N_17983,N_17912);
or U18177 (N_18177,N_17874,N_17606);
or U18178 (N_18178,N_17650,N_17984);
nand U18179 (N_18179,N_17659,N_17825);
nand U18180 (N_18180,N_17863,N_17614);
nor U18181 (N_18181,N_17946,N_17723);
xor U18182 (N_18182,N_17743,N_17634);
and U18183 (N_18183,N_17872,N_17893);
nor U18184 (N_18184,N_17793,N_17816);
xor U18185 (N_18185,N_17671,N_17875);
or U18186 (N_18186,N_17795,N_17643);
nor U18187 (N_18187,N_17602,N_17999);
nand U18188 (N_18188,N_17767,N_17982);
nand U18189 (N_18189,N_17859,N_17948);
or U18190 (N_18190,N_17858,N_17611);
nand U18191 (N_18191,N_17620,N_17676);
or U18192 (N_18192,N_17701,N_17976);
or U18193 (N_18193,N_17734,N_17840);
nand U18194 (N_18194,N_17605,N_17919);
xnor U18195 (N_18195,N_17939,N_17638);
and U18196 (N_18196,N_17990,N_17856);
nand U18197 (N_18197,N_17887,N_17683);
nor U18198 (N_18198,N_17660,N_17992);
nand U18199 (N_18199,N_17625,N_17642);
and U18200 (N_18200,N_17947,N_17973);
or U18201 (N_18201,N_17902,N_17722);
nand U18202 (N_18202,N_17601,N_17680);
xor U18203 (N_18203,N_17734,N_17793);
and U18204 (N_18204,N_17940,N_17801);
xor U18205 (N_18205,N_17724,N_17846);
xnor U18206 (N_18206,N_17974,N_17947);
or U18207 (N_18207,N_17696,N_17812);
xnor U18208 (N_18208,N_17664,N_17797);
xnor U18209 (N_18209,N_17869,N_17606);
and U18210 (N_18210,N_17611,N_17800);
nand U18211 (N_18211,N_17857,N_17679);
nand U18212 (N_18212,N_17769,N_17968);
xnor U18213 (N_18213,N_17936,N_17782);
xor U18214 (N_18214,N_17998,N_17765);
or U18215 (N_18215,N_17686,N_17675);
xor U18216 (N_18216,N_17849,N_17855);
or U18217 (N_18217,N_17916,N_17723);
or U18218 (N_18218,N_17953,N_17984);
xnor U18219 (N_18219,N_17758,N_17798);
or U18220 (N_18220,N_17808,N_17910);
and U18221 (N_18221,N_17955,N_17973);
and U18222 (N_18222,N_17924,N_17848);
nor U18223 (N_18223,N_17881,N_17762);
nor U18224 (N_18224,N_17794,N_17996);
or U18225 (N_18225,N_17888,N_17695);
and U18226 (N_18226,N_17892,N_17814);
or U18227 (N_18227,N_17960,N_17852);
or U18228 (N_18228,N_17916,N_17708);
or U18229 (N_18229,N_17656,N_17754);
xnor U18230 (N_18230,N_17848,N_17861);
and U18231 (N_18231,N_17642,N_17710);
nand U18232 (N_18232,N_17740,N_17954);
nor U18233 (N_18233,N_17635,N_17817);
nand U18234 (N_18234,N_17944,N_17701);
nand U18235 (N_18235,N_17927,N_17693);
nand U18236 (N_18236,N_17892,N_17977);
or U18237 (N_18237,N_17879,N_17939);
and U18238 (N_18238,N_17816,N_17706);
and U18239 (N_18239,N_17954,N_17719);
xor U18240 (N_18240,N_17793,N_17840);
nand U18241 (N_18241,N_17894,N_17784);
nor U18242 (N_18242,N_17667,N_17735);
and U18243 (N_18243,N_17898,N_17734);
or U18244 (N_18244,N_17770,N_17623);
xor U18245 (N_18245,N_17871,N_17616);
xor U18246 (N_18246,N_17883,N_17604);
xor U18247 (N_18247,N_17737,N_17757);
xnor U18248 (N_18248,N_17742,N_17628);
nor U18249 (N_18249,N_17990,N_17796);
nor U18250 (N_18250,N_17936,N_17746);
nor U18251 (N_18251,N_17824,N_17608);
and U18252 (N_18252,N_17910,N_17665);
xor U18253 (N_18253,N_17691,N_17677);
xnor U18254 (N_18254,N_17886,N_17798);
or U18255 (N_18255,N_17696,N_17660);
nand U18256 (N_18256,N_17892,N_17850);
and U18257 (N_18257,N_17722,N_17964);
nand U18258 (N_18258,N_17679,N_17941);
or U18259 (N_18259,N_17697,N_17609);
nor U18260 (N_18260,N_17706,N_17758);
or U18261 (N_18261,N_17928,N_17621);
nor U18262 (N_18262,N_17952,N_17914);
nand U18263 (N_18263,N_17710,N_17919);
nand U18264 (N_18264,N_17753,N_17640);
or U18265 (N_18265,N_17892,N_17890);
nor U18266 (N_18266,N_17825,N_17776);
nor U18267 (N_18267,N_17973,N_17688);
or U18268 (N_18268,N_17861,N_17726);
or U18269 (N_18269,N_17940,N_17925);
xor U18270 (N_18270,N_17824,N_17724);
xor U18271 (N_18271,N_17939,N_17647);
or U18272 (N_18272,N_17999,N_17825);
nand U18273 (N_18273,N_17853,N_17800);
or U18274 (N_18274,N_17660,N_17654);
and U18275 (N_18275,N_17864,N_17847);
nand U18276 (N_18276,N_17919,N_17826);
xnor U18277 (N_18277,N_17997,N_17796);
nor U18278 (N_18278,N_17910,N_17915);
nand U18279 (N_18279,N_17928,N_17874);
or U18280 (N_18280,N_17696,N_17789);
xor U18281 (N_18281,N_17851,N_17729);
and U18282 (N_18282,N_17858,N_17794);
and U18283 (N_18283,N_17600,N_17666);
and U18284 (N_18284,N_17780,N_17879);
or U18285 (N_18285,N_17992,N_17672);
nor U18286 (N_18286,N_17818,N_17927);
xnor U18287 (N_18287,N_17785,N_17876);
nand U18288 (N_18288,N_17675,N_17833);
nand U18289 (N_18289,N_17840,N_17937);
nand U18290 (N_18290,N_17805,N_17854);
and U18291 (N_18291,N_17875,N_17737);
and U18292 (N_18292,N_17955,N_17717);
and U18293 (N_18293,N_17946,N_17803);
or U18294 (N_18294,N_17985,N_17833);
nor U18295 (N_18295,N_17780,N_17899);
or U18296 (N_18296,N_17921,N_17838);
nor U18297 (N_18297,N_17813,N_17628);
nand U18298 (N_18298,N_17665,N_17857);
xor U18299 (N_18299,N_17698,N_17942);
and U18300 (N_18300,N_17734,N_17765);
or U18301 (N_18301,N_17810,N_17742);
xor U18302 (N_18302,N_17915,N_17722);
nor U18303 (N_18303,N_17771,N_17782);
and U18304 (N_18304,N_17705,N_17735);
or U18305 (N_18305,N_17947,N_17852);
and U18306 (N_18306,N_17996,N_17715);
nor U18307 (N_18307,N_17900,N_17779);
nand U18308 (N_18308,N_17932,N_17633);
or U18309 (N_18309,N_17903,N_17788);
and U18310 (N_18310,N_17996,N_17734);
nor U18311 (N_18311,N_17986,N_17809);
and U18312 (N_18312,N_17699,N_17974);
or U18313 (N_18313,N_17900,N_17693);
or U18314 (N_18314,N_17608,N_17851);
nand U18315 (N_18315,N_17962,N_17796);
or U18316 (N_18316,N_17648,N_17777);
and U18317 (N_18317,N_17761,N_17744);
and U18318 (N_18318,N_17657,N_17722);
nor U18319 (N_18319,N_17659,N_17873);
or U18320 (N_18320,N_17796,N_17889);
nor U18321 (N_18321,N_17976,N_17725);
xnor U18322 (N_18322,N_17719,N_17756);
nand U18323 (N_18323,N_17859,N_17855);
or U18324 (N_18324,N_17840,N_17611);
and U18325 (N_18325,N_17902,N_17725);
and U18326 (N_18326,N_17909,N_17853);
nand U18327 (N_18327,N_17970,N_17705);
nand U18328 (N_18328,N_17683,N_17662);
and U18329 (N_18329,N_17677,N_17866);
nand U18330 (N_18330,N_17711,N_17910);
xnor U18331 (N_18331,N_17616,N_17845);
nor U18332 (N_18332,N_17939,N_17906);
xnor U18333 (N_18333,N_17781,N_17989);
xnor U18334 (N_18334,N_17819,N_17853);
xnor U18335 (N_18335,N_17951,N_17708);
or U18336 (N_18336,N_17836,N_17929);
xnor U18337 (N_18337,N_17915,N_17941);
nand U18338 (N_18338,N_17982,N_17708);
nor U18339 (N_18339,N_17987,N_17650);
nor U18340 (N_18340,N_17987,N_17874);
or U18341 (N_18341,N_17888,N_17828);
or U18342 (N_18342,N_17910,N_17901);
nor U18343 (N_18343,N_17921,N_17753);
or U18344 (N_18344,N_17987,N_17938);
nand U18345 (N_18345,N_17896,N_17851);
nand U18346 (N_18346,N_17726,N_17813);
nor U18347 (N_18347,N_17958,N_17796);
nand U18348 (N_18348,N_17941,N_17665);
or U18349 (N_18349,N_17741,N_17640);
nor U18350 (N_18350,N_17943,N_17860);
nand U18351 (N_18351,N_17601,N_17895);
or U18352 (N_18352,N_17795,N_17922);
xor U18353 (N_18353,N_17901,N_17791);
and U18354 (N_18354,N_17806,N_17749);
nor U18355 (N_18355,N_17831,N_17803);
xor U18356 (N_18356,N_17888,N_17653);
nand U18357 (N_18357,N_17909,N_17770);
or U18358 (N_18358,N_17923,N_17600);
xnor U18359 (N_18359,N_17638,N_17605);
nor U18360 (N_18360,N_17725,N_17614);
or U18361 (N_18361,N_17869,N_17811);
xor U18362 (N_18362,N_17675,N_17844);
and U18363 (N_18363,N_17844,N_17910);
nor U18364 (N_18364,N_17675,N_17949);
and U18365 (N_18365,N_17638,N_17867);
nor U18366 (N_18366,N_17830,N_17780);
and U18367 (N_18367,N_17750,N_17847);
or U18368 (N_18368,N_17616,N_17964);
xor U18369 (N_18369,N_17981,N_17986);
and U18370 (N_18370,N_17950,N_17651);
or U18371 (N_18371,N_17957,N_17997);
xnor U18372 (N_18372,N_17827,N_17639);
nor U18373 (N_18373,N_17955,N_17677);
and U18374 (N_18374,N_17885,N_17692);
xnor U18375 (N_18375,N_17613,N_17853);
xor U18376 (N_18376,N_17824,N_17725);
xor U18377 (N_18377,N_17671,N_17753);
or U18378 (N_18378,N_17798,N_17945);
xnor U18379 (N_18379,N_17691,N_17783);
nand U18380 (N_18380,N_17840,N_17843);
or U18381 (N_18381,N_17981,N_17710);
nand U18382 (N_18382,N_17771,N_17703);
nand U18383 (N_18383,N_17856,N_17883);
nand U18384 (N_18384,N_17738,N_17799);
and U18385 (N_18385,N_17955,N_17835);
nor U18386 (N_18386,N_17830,N_17801);
nor U18387 (N_18387,N_17699,N_17706);
xnor U18388 (N_18388,N_17852,N_17707);
or U18389 (N_18389,N_17957,N_17634);
and U18390 (N_18390,N_17758,N_17866);
nand U18391 (N_18391,N_17860,N_17625);
or U18392 (N_18392,N_17910,N_17751);
xnor U18393 (N_18393,N_17959,N_17952);
nand U18394 (N_18394,N_17870,N_17648);
nor U18395 (N_18395,N_17958,N_17783);
xor U18396 (N_18396,N_17770,N_17884);
xnor U18397 (N_18397,N_17700,N_17748);
and U18398 (N_18398,N_17867,N_17816);
xnor U18399 (N_18399,N_17759,N_17913);
nand U18400 (N_18400,N_18032,N_18152);
and U18401 (N_18401,N_18165,N_18214);
nor U18402 (N_18402,N_18205,N_18069);
nor U18403 (N_18403,N_18235,N_18372);
or U18404 (N_18404,N_18121,N_18182);
nand U18405 (N_18405,N_18241,N_18019);
or U18406 (N_18406,N_18000,N_18197);
nor U18407 (N_18407,N_18074,N_18359);
and U18408 (N_18408,N_18288,N_18078);
nor U18409 (N_18409,N_18128,N_18090);
nand U18410 (N_18410,N_18124,N_18357);
nor U18411 (N_18411,N_18106,N_18271);
and U18412 (N_18412,N_18306,N_18260);
xnor U18413 (N_18413,N_18058,N_18111);
nand U18414 (N_18414,N_18355,N_18342);
xor U18415 (N_18415,N_18335,N_18356);
and U18416 (N_18416,N_18139,N_18274);
or U18417 (N_18417,N_18167,N_18251);
xnor U18418 (N_18418,N_18303,N_18300);
nand U18419 (N_18419,N_18277,N_18224);
nor U18420 (N_18420,N_18118,N_18311);
xnor U18421 (N_18421,N_18201,N_18374);
or U18422 (N_18422,N_18172,N_18313);
xor U18423 (N_18423,N_18004,N_18093);
nand U18424 (N_18424,N_18168,N_18364);
xor U18425 (N_18425,N_18006,N_18315);
nand U18426 (N_18426,N_18248,N_18089);
and U18427 (N_18427,N_18247,N_18350);
nor U18428 (N_18428,N_18353,N_18378);
nand U18429 (N_18429,N_18179,N_18320);
xor U18430 (N_18430,N_18102,N_18107);
and U18431 (N_18431,N_18367,N_18203);
xnor U18432 (N_18432,N_18098,N_18200);
nand U18433 (N_18433,N_18029,N_18162);
xor U18434 (N_18434,N_18227,N_18123);
or U18435 (N_18435,N_18264,N_18043);
nand U18436 (N_18436,N_18084,N_18243);
or U18437 (N_18437,N_18094,N_18016);
xor U18438 (N_18438,N_18075,N_18083);
nor U18439 (N_18439,N_18164,N_18337);
and U18440 (N_18440,N_18012,N_18304);
nor U18441 (N_18441,N_18081,N_18163);
or U18442 (N_18442,N_18092,N_18021);
nand U18443 (N_18443,N_18289,N_18238);
and U18444 (N_18444,N_18343,N_18041);
nor U18445 (N_18445,N_18381,N_18030);
nand U18446 (N_18446,N_18129,N_18368);
nor U18447 (N_18447,N_18250,N_18190);
or U18448 (N_18448,N_18044,N_18209);
xnor U18449 (N_18449,N_18064,N_18176);
or U18450 (N_18450,N_18284,N_18377);
and U18451 (N_18451,N_18317,N_18026);
or U18452 (N_18452,N_18354,N_18252);
and U18453 (N_18453,N_18134,N_18397);
or U18454 (N_18454,N_18031,N_18216);
and U18455 (N_18455,N_18067,N_18398);
and U18456 (N_18456,N_18314,N_18148);
nand U18457 (N_18457,N_18301,N_18399);
nor U18458 (N_18458,N_18346,N_18358);
xor U18459 (N_18459,N_18322,N_18285);
nand U18460 (N_18460,N_18215,N_18033);
xnor U18461 (N_18461,N_18345,N_18228);
nor U18462 (N_18462,N_18347,N_18151);
nor U18463 (N_18463,N_18157,N_18333);
xnor U18464 (N_18464,N_18115,N_18234);
or U18465 (N_18465,N_18109,N_18059);
or U18466 (N_18466,N_18376,N_18174);
xor U18467 (N_18467,N_18253,N_18045);
or U18468 (N_18468,N_18291,N_18237);
nor U18469 (N_18469,N_18334,N_18126);
or U18470 (N_18470,N_18037,N_18052);
or U18471 (N_18471,N_18395,N_18036);
and U18472 (N_18472,N_18338,N_18208);
xor U18473 (N_18473,N_18013,N_18087);
and U18474 (N_18474,N_18020,N_18137);
nand U18475 (N_18475,N_18387,N_18386);
xor U18476 (N_18476,N_18096,N_18221);
nand U18477 (N_18477,N_18014,N_18257);
nand U18478 (N_18478,N_18155,N_18170);
xnor U18479 (N_18479,N_18336,N_18103);
nor U18480 (N_18480,N_18144,N_18082);
or U18481 (N_18481,N_18344,N_18242);
or U18482 (N_18482,N_18175,N_18024);
nand U18483 (N_18483,N_18255,N_18113);
xnor U18484 (N_18484,N_18140,N_18049);
nor U18485 (N_18485,N_18352,N_18389);
nor U18486 (N_18486,N_18097,N_18181);
nand U18487 (N_18487,N_18196,N_18373);
or U18488 (N_18488,N_18068,N_18239);
xor U18489 (N_18489,N_18070,N_18204);
nor U18490 (N_18490,N_18233,N_18263);
nand U18491 (N_18491,N_18307,N_18022);
and U18492 (N_18492,N_18138,N_18363);
and U18493 (N_18493,N_18323,N_18171);
xnor U18494 (N_18494,N_18072,N_18226);
or U18495 (N_18495,N_18153,N_18293);
xnor U18496 (N_18496,N_18266,N_18051);
or U18497 (N_18497,N_18169,N_18076);
nor U18498 (N_18498,N_18254,N_18360);
xnor U18499 (N_18499,N_18276,N_18133);
and U18500 (N_18500,N_18127,N_18244);
nor U18501 (N_18501,N_18340,N_18003);
nand U18502 (N_18502,N_18027,N_18268);
nor U18503 (N_18503,N_18213,N_18310);
xnor U18504 (N_18504,N_18281,N_18091);
nand U18505 (N_18505,N_18206,N_18286);
and U18506 (N_18506,N_18001,N_18391);
nor U18507 (N_18507,N_18073,N_18015);
xor U18508 (N_18508,N_18278,N_18189);
or U18509 (N_18509,N_18010,N_18222);
xnor U18510 (N_18510,N_18161,N_18256);
xor U18511 (N_18511,N_18086,N_18230);
xnor U18512 (N_18512,N_18055,N_18393);
nor U18513 (N_18513,N_18180,N_18194);
nand U18514 (N_18514,N_18132,N_18283);
or U18515 (N_18515,N_18063,N_18223);
xnor U18516 (N_18516,N_18120,N_18394);
nor U18517 (N_18517,N_18219,N_18187);
nor U18518 (N_18518,N_18341,N_18100);
xnor U18519 (N_18519,N_18231,N_18195);
nand U18520 (N_18520,N_18108,N_18142);
or U18521 (N_18521,N_18249,N_18380);
nor U18522 (N_18522,N_18366,N_18327);
and U18523 (N_18523,N_18296,N_18185);
nor U18524 (N_18524,N_18125,N_18156);
nor U18525 (N_18525,N_18028,N_18057);
or U18526 (N_18526,N_18330,N_18265);
nor U18527 (N_18527,N_18130,N_18023);
xor U18528 (N_18528,N_18385,N_18259);
or U18529 (N_18529,N_18302,N_18066);
xnor U18530 (N_18530,N_18245,N_18305);
or U18531 (N_18531,N_18105,N_18038);
or U18532 (N_18532,N_18297,N_18048);
and U18533 (N_18533,N_18316,N_18034);
and U18534 (N_18534,N_18351,N_18217);
and U18535 (N_18535,N_18388,N_18077);
nand U18536 (N_18536,N_18396,N_18309);
nand U18537 (N_18537,N_18065,N_18240);
and U18538 (N_18538,N_18047,N_18273);
or U18539 (N_18539,N_18225,N_18390);
nor U18540 (N_18540,N_18246,N_18101);
xor U18541 (N_18541,N_18158,N_18112);
or U18542 (N_18542,N_18079,N_18099);
nor U18543 (N_18543,N_18329,N_18236);
nor U18544 (N_18544,N_18318,N_18116);
nand U18545 (N_18545,N_18184,N_18198);
or U18546 (N_18546,N_18375,N_18060);
nand U18547 (N_18547,N_18150,N_18299);
nand U18548 (N_18548,N_18362,N_18009);
or U18549 (N_18549,N_18280,N_18370);
nand U18550 (N_18550,N_18007,N_18183);
and U18551 (N_18551,N_18326,N_18365);
and U18552 (N_18552,N_18218,N_18011);
or U18553 (N_18553,N_18191,N_18328);
and U18554 (N_18554,N_18080,N_18122);
and U18555 (N_18555,N_18002,N_18319);
and U18556 (N_18556,N_18202,N_18017);
and U18557 (N_18557,N_18262,N_18384);
nand U18558 (N_18558,N_18261,N_18258);
or U18559 (N_18559,N_18348,N_18383);
xnor U18560 (N_18560,N_18095,N_18008);
and U18561 (N_18561,N_18324,N_18178);
xnor U18562 (N_18562,N_18061,N_18292);
and U18563 (N_18563,N_18220,N_18325);
nand U18564 (N_18564,N_18207,N_18177);
or U18565 (N_18565,N_18193,N_18272);
nand U18566 (N_18566,N_18339,N_18210);
nand U18567 (N_18567,N_18298,N_18149);
or U18568 (N_18568,N_18104,N_18166);
nand U18569 (N_18569,N_18173,N_18025);
nand U18570 (N_18570,N_18275,N_18135);
and U18571 (N_18571,N_18211,N_18308);
and U18572 (N_18572,N_18119,N_18294);
xor U18573 (N_18573,N_18186,N_18143);
nand U18574 (N_18574,N_18332,N_18062);
and U18575 (N_18575,N_18279,N_18270);
nor U18576 (N_18576,N_18229,N_18136);
nand U18577 (N_18577,N_18146,N_18361);
xnor U18578 (N_18578,N_18312,N_18040);
and U18579 (N_18579,N_18039,N_18141);
nor U18580 (N_18580,N_18232,N_18088);
or U18581 (N_18581,N_18295,N_18159);
and U18582 (N_18582,N_18188,N_18054);
nand U18583 (N_18583,N_18382,N_18071);
nand U18584 (N_18584,N_18056,N_18053);
xnor U18585 (N_18585,N_18267,N_18212);
or U18586 (N_18586,N_18371,N_18199);
or U18587 (N_18587,N_18145,N_18349);
xor U18588 (N_18588,N_18160,N_18321);
nor U18589 (N_18589,N_18269,N_18042);
nor U18590 (N_18590,N_18290,N_18282);
nand U18591 (N_18591,N_18085,N_18331);
nand U18592 (N_18592,N_18154,N_18147);
and U18593 (N_18593,N_18035,N_18050);
nor U18594 (N_18594,N_18110,N_18287);
or U18595 (N_18595,N_18046,N_18192);
nor U18596 (N_18596,N_18114,N_18369);
or U18597 (N_18597,N_18005,N_18131);
or U18598 (N_18598,N_18379,N_18117);
nor U18599 (N_18599,N_18018,N_18392);
and U18600 (N_18600,N_18022,N_18351);
xnor U18601 (N_18601,N_18030,N_18088);
nor U18602 (N_18602,N_18324,N_18311);
and U18603 (N_18603,N_18024,N_18086);
xnor U18604 (N_18604,N_18038,N_18369);
nor U18605 (N_18605,N_18282,N_18031);
and U18606 (N_18606,N_18126,N_18098);
nand U18607 (N_18607,N_18237,N_18019);
xnor U18608 (N_18608,N_18244,N_18058);
or U18609 (N_18609,N_18272,N_18323);
or U18610 (N_18610,N_18267,N_18280);
nor U18611 (N_18611,N_18260,N_18011);
and U18612 (N_18612,N_18266,N_18195);
nand U18613 (N_18613,N_18286,N_18299);
nand U18614 (N_18614,N_18331,N_18336);
and U18615 (N_18615,N_18127,N_18155);
xnor U18616 (N_18616,N_18161,N_18327);
xnor U18617 (N_18617,N_18258,N_18140);
nor U18618 (N_18618,N_18271,N_18347);
nand U18619 (N_18619,N_18098,N_18387);
nand U18620 (N_18620,N_18306,N_18139);
and U18621 (N_18621,N_18303,N_18261);
xor U18622 (N_18622,N_18205,N_18145);
xnor U18623 (N_18623,N_18031,N_18309);
xnor U18624 (N_18624,N_18319,N_18109);
xor U18625 (N_18625,N_18099,N_18313);
nor U18626 (N_18626,N_18128,N_18197);
nor U18627 (N_18627,N_18105,N_18270);
or U18628 (N_18628,N_18285,N_18193);
nand U18629 (N_18629,N_18026,N_18043);
nand U18630 (N_18630,N_18316,N_18337);
xor U18631 (N_18631,N_18233,N_18074);
nand U18632 (N_18632,N_18033,N_18243);
nand U18633 (N_18633,N_18392,N_18329);
or U18634 (N_18634,N_18311,N_18005);
xnor U18635 (N_18635,N_18134,N_18275);
nand U18636 (N_18636,N_18077,N_18013);
nor U18637 (N_18637,N_18364,N_18291);
nand U18638 (N_18638,N_18308,N_18040);
xor U18639 (N_18639,N_18390,N_18030);
or U18640 (N_18640,N_18367,N_18071);
nor U18641 (N_18641,N_18142,N_18199);
and U18642 (N_18642,N_18393,N_18025);
and U18643 (N_18643,N_18096,N_18374);
and U18644 (N_18644,N_18033,N_18232);
or U18645 (N_18645,N_18017,N_18027);
or U18646 (N_18646,N_18139,N_18332);
and U18647 (N_18647,N_18300,N_18099);
and U18648 (N_18648,N_18204,N_18017);
nand U18649 (N_18649,N_18185,N_18141);
xor U18650 (N_18650,N_18156,N_18272);
and U18651 (N_18651,N_18292,N_18274);
nand U18652 (N_18652,N_18319,N_18396);
nor U18653 (N_18653,N_18247,N_18198);
nand U18654 (N_18654,N_18367,N_18157);
and U18655 (N_18655,N_18098,N_18341);
or U18656 (N_18656,N_18327,N_18296);
nand U18657 (N_18657,N_18294,N_18385);
or U18658 (N_18658,N_18242,N_18254);
xor U18659 (N_18659,N_18216,N_18095);
nand U18660 (N_18660,N_18360,N_18094);
nand U18661 (N_18661,N_18364,N_18094);
nor U18662 (N_18662,N_18143,N_18161);
xnor U18663 (N_18663,N_18180,N_18317);
nand U18664 (N_18664,N_18065,N_18279);
xnor U18665 (N_18665,N_18032,N_18072);
or U18666 (N_18666,N_18022,N_18314);
and U18667 (N_18667,N_18344,N_18188);
nor U18668 (N_18668,N_18147,N_18369);
xor U18669 (N_18669,N_18075,N_18142);
or U18670 (N_18670,N_18098,N_18133);
nand U18671 (N_18671,N_18221,N_18262);
or U18672 (N_18672,N_18146,N_18112);
and U18673 (N_18673,N_18103,N_18276);
nor U18674 (N_18674,N_18223,N_18356);
xnor U18675 (N_18675,N_18011,N_18312);
nand U18676 (N_18676,N_18391,N_18078);
xnor U18677 (N_18677,N_18149,N_18289);
xor U18678 (N_18678,N_18119,N_18277);
and U18679 (N_18679,N_18204,N_18374);
nand U18680 (N_18680,N_18187,N_18013);
or U18681 (N_18681,N_18315,N_18147);
and U18682 (N_18682,N_18141,N_18145);
nand U18683 (N_18683,N_18367,N_18364);
and U18684 (N_18684,N_18294,N_18276);
and U18685 (N_18685,N_18057,N_18047);
or U18686 (N_18686,N_18372,N_18166);
xnor U18687 (N_18687,N_18210,N_18326);
or U18688 (N_18688,N_18102,N_18197);
xor U18689 (N_18689,N_18320,N_18310);
nand U18690 (N_18690,N_18029,N_18270);
nand U18691 (N_18691,N_18218,N_18381);
and U18692 (N_18692,N_18181,N_18150);
and U18693 (N_18693,N_18001,N_18371);
xnor U18694 (N_18694,N_18275,N_18350);
nor U18695 (N_18695,N_18213,N_18212);
and U18696 (N_18696,N_18212,N_18164);
xor U18697 (N_18697,N_18255,N_18207);
and U18698 (N_18698,N_18234,N_18356);
and U18699 (N_18699,N_18075,N_18199);
nand U18700 (N_18700,N_18391,N_18316);
and U18701 (N_18701,N_18317,N_18292);
xor U18702 (N_18702,N_18338,N_18216);
or U18703 (N_18703,N_18339,N_18245);
and U18704 (N_18704,N_18008,N_18028);
nand U18705 (N_18705,N_18141,N_18274);
nand U18706 (N_18706,N_18023,N_18166);
and U18707 (N_18707,N_18099,N_18169);
xnor U18708 (N_18708,N_18254,N_18144);
nor U18709 (N_18709,N_18384,N_18248);
and U18710 (N_18710,N_18120,N_18386);
or U18711 (N_18711,N_18336,N_18074);
xor U18712 (N_18712,N_18263,N_18393);
xnor U18713 (N_18713,N_18011,N_18042);
and U18714 (N_18714,N_18169,N_18350);
nor U18715 (N_18715,N_18385,N_18048);
nand U18716 (N_18716,N_18187,N_18080);
nor U18717 (N_18717,N_18066,N_18356);
and U18718 (N_18718,N_18150,N_18384);
nand U18719 (N_18719,N_18050,N_18207);
and U18720 (N_18720,N_18287,N_18093);
and U18721 (N_18721,N_18287,N_18297);
nor U18722 (N_18722,N_18390,N_18044);
xnor U18723 (N_18723,N_18075,N_18061);
and U18724 (N_18724,N_18338,N_18186);
or U18725 (N_18725,N_18048,N_18333);
nand U18726 (N_18726,N_18258,N_18153);
or U18727 (N_18727,N_18222,N_18274);
nor U18728 (N_18728,N_18372,N_18317);
nor U18729 (N_18729,N_18043,N_18289);
and U18730 (N_18730,N_18318,N_18275);
nand U18731 (N_18731,N_18240,N_18133);
or U18732 (N_18732,N_18207,N_18223);
nor U18733 (N_18733,N_18325,N_18344);
nor U18734 (N_18734,N_18109,N_18310);
nor U18735 (N_18735,N_18332,N_18038);
nand U18736 (N_18736,N_18272,N_18159);
xor U18737 (N_18737,N_18336,N_18381);
and U18738 (N_18738,N_18202,N_18184);
nor U18739 (N_18739,N_18135,N_18144);
nor U18740 (N_18740,N_18007,N_18203);
xnor U18741 (N_18741,N_18071,N_18256);
nor U18742 (N_18742,N_18252,N_18050);
and U18743 (N_18743,N_18189,N_18285);
or U18744 (N_18744,N_18345,N_18191);
xnor U18745 (N_18745,N_18278,N_18260);
nor U18746 (N_18746,N_18065,N_18141);
nor U18747 (N_18747,N_18123,N_18230);
nand U18748 (N_18748,N_18030,N_18396);
and U18749 (N_18749,N_18092,N_18024);
xor U18750 (N_18750,N_18137,N_18242);
xnor U18751 (N_18751,N_18045,N_18149);
or U18752 (N_18752,N_18038,N_18157);
xnor U18753 (N_18753,N_18121,N_18248);
and U18754 (N_18754,N_18108,N_18236);
or U18755 (N_18755,N_18057,N_18310);
or U18756 (N_18756,N_18298,N_18257);
or U18757 (N_18757,N_18304,N_18224);
and U18758 (N_18758,N_18254,N_18108);
nor U18759 (N_18759,N_18022,N_18397);
or U18760 (N_18760,N_18004,N_18210);
or U18761 (N_18761,N_18058,N_18335);
nor U18762 (N_18762,N_18210,N_18370);
nand U18763 (N_18763,N_18122,N_18133);
xor U18764 (N_18764,N_18380,N_18280);
xnor U18765 (N_18765,N_18144,N_18194);
nand U18766 (N_18766,N_18037,N_18241);
and U18767 (N_18767,N_18093,N_18273);
or U18768 (N_18768,N_18269,N_18390);
nor U18769 (N_18769,N_18331,N_18340);
xor U18770 (N_18770,N_18198,N_18114);
or U18771 (N_18771,N_18037,N_18248);
and U18772 (N_18772,N_18387,N_18291);
nand U18773 (N_18773,N_18227,N_18163);
nand U18774 (N_18774,N_18297,N_18347);
nor U18775 (N_18775,N_18037,N_18296);
nor U18776 (N_18776,N_18393,N_18297);
nor U18777 (N_18777,N_18156,N_18295);
and U18778 (N_18778,N_18362,N_18203);
and U18779 (N_18779,N_18282,N_18198);
nand U18780 (N_18780,N_18105,N_18174);
nor U18781 (N_18781,N_18372,N_18229);
or U18782 (N_18782,N_18043,N_18188);
and U18783 (N_18783,N_18350,N_18386);
xnor U18784 (N_18784,N_18235,N_18128);
and U18785 (N_18785,N_18309,N_18248);
and U18786 (N_18786,N_18165,N_18115);
xnor U18787 (N_18787,N_18172,N_18036);
nor U18788 (N_18788,N_18087,N_18132);
or U18789 (N_18789,N_18361,N_18215);
xnor U18790 (N_18790,N_18265,N_18324);
nor U18791 (N_18791,N_18265,N_18098);
xor U18792 (N_18792,N_18285,N_18119);
and U18793 (N_18793,N_18313,N_18325);
nor U18794 (N_18794,N_18273,N_18248);
and U18795 (N_18795,N_18113,N_18316);
nor U18796 (N_18796,N_18081,N_18288);
or U18797 (N_18797,N_18350,N_18013);
nor U18798 (N_18798,N_18399,N_18063);
xnor U18799 (N_18799,N_18308,N_18314);
xnor U18800 (N_18800,N_18580,N_18572);
or U18801 (N_18801,N_18615,N_18622);
and U18802 (N_18802,N_18701,N_18737);
nand U18803 (N_18803,N_18550,N_18487);
nand U18804 (N_18804,N_18512,N_18457);
and U18805 (N_18805,N_18412,N_18650);
or U18806 (N_18806,N_18534,N_18728);
nor U18807 (N_18807,N_18593,N_18418);
xnor U18808 (N_18808,N_18716,N_18536);
xor U18809 (N_18809,N_18627,N_18634);
nor U18810 (N_18810,N_18604,N_18796);
xor U18811 (N_18811,N_18744,N_18416);
xnor U18812 (N_18812,N_18519,N_18433);
nand U18813 (N_18813,N_18422,N_18426);
and U18814 (N_18814,N_18733,N_18724);
and U18815 (N_18815,N_18540,N_18405);
and U18816 (N_18816,N_18669,N_18791);
and U18817 (N_18817,N_18727,N_18612);
and U18818 (N_18818,N_18779,N_18662);
nand U18819 (N_18819,N_18432,N_18456);
nor U18820 (N_18820,N_18569,N_18657);
xnor U18821 (N_18821,N_18786,N_18640);
xor U18822 (N_18822,N_18764,N_18408);
or U18823 (N_18823,N_18795,N_18503);
and U18824 (N_18824,N_18517,N_18450);
nand U18825 (N_18825,N_18467,N_18749);
and U18826 (N_18826,N_18476,N_18792);
xnor U18827 (N_18827,N_18601,N_18680);
and U18828 (N_18828,N_18451,N_18788);
and U18829 (N_18829,N_18410,N_18472);
nor U18830 (N_18830,N_18531,N_18409);
nand U18831 (N_18831,N_18676,N_18685);
nor U18832 (N_18832,N_18417,N_18637);
and U18833 (N_18833,N_18736,N_18571);
nor U18834 (N_18834,N_18780,N_18789);
nand U18835 (N_18835,N_18548,N_18730);
xnor U18836 (N_18836,N_18756,N_18643);
xor U18837 (N_18837,N_18523,N_18694);
nor U18838 (N_18838,N_18673,N_18753);
xnor U18839 (N_18839,N_18696,N_18771);
and U18840 (N_18840,N_18507,N_18579);
and U18841 (N_18841,N_18630,N_18504);
nor U18842 (N_18842,N_18443,N_18436);
and U18843 (N_18843,N_18570,N_18718);
nor U18844 (N_18844,N_18755,N_18751);
xor U18845 (N_18845,N_18427,N_18715);
nor U18846 (N_18846,N_18794,N_18679);
nand U18847 (N_18847,N_18624,N_18797);
or U18848 (N_18848,N_18793,N_18494);
nand U18849 (N_18849,N_18459,N_18402);
nand U18850 (N_18850,N_18545,N_18552);
or U18851 (N_18851,N_18524,N_18629);
nand U18852 (N_18852,N_18614,N_18485);
and U18853 (N_18853,N_18777,N_18430);
or U18854 (N_18854,N_18605,N_18463);
nor U18855 (N_18855,N_18522,N_18717);
xnor U18856 (N_18856,N_18513,N_18576);
nand U18857 (N_18857,N_18760,N_18675);
nor U18858 (N_18858,N_18404,N_18510);
nor U18859 (N_18859,N_18681,N_18722);
or U18860 (N_18860,N_18619,N_18496);
and U18861 (N_18861,N_18471,N_18709);
nor U18862 (N_18862,N_18411,N_18773);
nor U18863 (N_18863,N_18732,N_18420);
and U18864 (N_18864,N_18678,N_18769);
nand U18865 (N_18865,N_18484,N_18491);
and U18866 (N_18866,N_18700,N_18582);
nor U18867 (N_18867,N_18719,N_18564);
and U18868 (N_18868,N_18474,N_18714);
nor U18869 (N_18869,N_18492,N_18557);
xnor U18870 (N_18870,N_18466,N_18697);
nand U18871 (N_18871,N_18489,N_18446);
and U18872 (N_18872,N_18584,N_18514);
and U18873 (N_18873,N_18508,N_18734);
nor U18874 (N_18874,N_18691,N_18664);
or U18875 (N_18875,N_18578,N_18588);
and U18876 (N_18876,N_18704,N_18563);
xor U18877 (N_18877,N_18558,N_18415);
or U18878 (N_18878,N_18782,N_18677);
nor U18879 (N_18879,N_18766,N_18767);
nor U18880 (N_18880,N_18652,N_18441);
and U18881 (N_18881,N_18470,N_18549);
and U18882 (N_18882,N_18428,N_18535);
nand U18883 (N_18883,N_18455,N_18538);
and U18884 (N_18884,N_18618,N_18687);
nor U18885 (N_18885,N_18639,N_18596);
or U18886 (N_18886,N_18444,N_18628);
xor U18887 (N_18887,N_18661,N_18401);
and U18888 (N_18888,N_18665,N_18663);
and U18889 (N_18889,N_18790,N_18620);
nor U18890 (N_18890,N_18617,N_18725);
nand U18891 (N_18891,N_18595,N_18465);
nor U18892 (N_18892,N_18464,N_18787);
and U18893 (N_18893,N_18561,N_18559);
nand U18894 (N_18894,N_18473,N_18439);
and U18895 (N_18895,N_18742,N_18554);
or U18896 (N_18896,N_18530,N_18560);
xnor U18897 (N_18897,N_18688,N_18525);
and U18898 (N_18898,N_18635,N_18425);
and U18899 (N_18899,N_18692,N_18509);
xor U18900 (N_18900,N_18798,N_18672);
or U18901 (N_18901,N_18602,N_18458);
and U18902 (N_18902,N_18479,N_18775);
and U18903 (N_18903,N_18651,N_18641);
and U18904 (N_18904,N_18452,N_18448);
or U18905 (N_18905,N_18495,N_18453);
nor U18906 (N_18906,N_18565,N_18750);
nor U18907 (N_18907,N_18625,N_18532);
and U18908 (N_18908,N_18726,N_18480);
and U18909 (N_18909,N_18445,N_18746);
and U18910 (N_18910,N_18702,N_18407);
xnor U18911 (N_18911,N_18553,N_18539);
and U18912 (N_18912,N_18449,N_18747);
or U18913 (N_18913,N_18555,N_18486);
or U18914 (N_18914,N_18655,N_18528);
xnor U18915 (N_18915,N_18761,N_18429);
xor U18916 (N_18916,N_18613,N_18499);
xor U18917 (N_18917,N_18784,N_18493);
xnor U18918 (N_18918,N_18656,N_18590);
or U18919 (N_18919,N_18518,N_18666);
and U18920 (N_18920,N_18757,N_18583);
nor U18921 (N_18921,N_18638,N_18686);
or U18922 (N_18922,N_18556,N_18671);
nand U18923 (N_18923,N_18482,N_18670);
nand U18924 (N_18924,N_18646,N_18573);
and U18925 (N_18925,N_18785,N_18469);
and U18926 (N_18926,N_18424,N_18501);
nor U18927 (N_18927,N_18438,N_18581);
or U18928 (N_18928,N_18649,N_18607);
and U18929 (N_18929,N_18698,N_18546);
nor U18930 (N_18930,N_18644,N_18413);
nor U18931 (N_18931,N_18772,N_18440);
nor U18932 (N_18932,N_18575,N_18659);
and U18933 (N_18933,N_18597,N_18707);
nor U18934 (N_18934,N_18414,N_18543);
xor U18935 (N_18935,N_18460,N_18592);
and U18936 (N_18936,N_18711,N_18654);
and U18937 (N_18937,N_18738,N_18591);
or U18938 (N_18938,N_18699,N_18632);
nand U18939 (N_18939,N_18674,N_18689);
and U18940 (N_18940,N_18713,N_18435);
nor U18941 (N_18941,N_18647,N_18481);
nand U18942 (N_18942,N_18748,N_18488);
nand U18943 (N_18943,N_18537,N_18626);
and U18944 (N_18944,N_18434,N_18475);
nor U18945 (N_18945,N_18631,N_18693);
nor U18946 (N_18946,N_18527,N_18500);
and U18947 (N_18947,N_18447,N_18403);
nand U18948 (N_18948,N_18498,N_18653);
nand U18949 (N_18949,N_18419,N_18759);
xnor U18950 (N_18950,N_18778,N_18754);
nor U18951 (N_18951,N_18533,N_18682);
or U18952 (N_18952,N_18490,N_18623);
nand U18953 (N_18953,N_18603,N_18589);
or U18954 (N_18954,N_18743,N_18526);
nand U18955 (N_18955,N_18710,N_18502);
xnor U18956 (N_18956,N_18609,N_18723);
nand U18957 (N_18957,N_18648,N_18568);
xor U18958 (N_18958,N_18721,N_18421);
and U18959 (N_18959,N_18542,N_18768);
nor U18960 (N_18960,N_18454,N_18520);
xor U18961 (N_18961,N_18642,N_18529);
or U18962 (N_18962,N_18712,N_18478);
and U18963 (N_18963,N_18598,N_18762);
and U18964 (N_18964,N_18729,N_18765);
xnor U18965 (N_18965,N_18683,N_18621);
or U18966 (N_18966,N_18741,N_18468);
nor U18967 (N_18967,N_18551,N_18660);
and U18968 (N_18968,N_18431,N_18585);
nand U18969 (N_18969,N_18477,N_18586);
and U18970 (N_18970,N_18406,N_18776);
nand U18971 (N_18971,N_18781,N_18783);
nand U18972 (N_18972,N_18544,N_18774);
xnor U18973 (N_18973,N_18516,N_18608);
nand U18974 (N_18974,N_18600,N_18442);
nor U18975 (N_18975,N_18423,N_18610);
nor U18976 (N_18976,N_18645,N_18599);
nand U18977 (N_18977,N_18611,N_18770);
nand U18978 (N_18978,N_18511,N_18752);
nor U18979 (N_18979,N_18483,N_18739);
and U18980 (N_18980,N_18735,N_18577);
or U18981 (N_18981,N_18758,N_18461);
nor U18982 (N_18982,N_18462,N_18799);
or U18983 (N_18983,N_18515,N_18731);
or U18984 (N_18984,N_18740,N_18705);
nor U18985 (N_18985,N_18668,N_18636);
or U18986 (N_18986,N_18521,N_18566);
nor U18987 (N_18987,N_18633,N_18400);
xnor U18988 (N_18988,N_18562,N_18567);
and U18989 (N_18989,N_18506,N_18667);
nor U18990 (N_18990,N_18690,N_18497);
or U18991 (N_18991,N_18505,N_18541);
nand U18992 (N_18992,N_18574,N_18547);
or U18993 (N_18993,N_18616,N_18708);
nor U18994 (N_18994,N_18594,N_18587);
or U18995 (N_18995,N_18703,N_18763);
nand U18996 (N_18996,N_18706,N_18695);
nand U18997 (N_18997,N_18720,N_18745);
or U18998 (N_18998,N_18606,N_18658);
nand U18999 (N_18999,N_18684,N_18437);
xor U19000 (N_19000,N_18664,N_18441);
nand U19001 (N_19001,N_18706,N_18478);
nor U19002 (N_19002,N_18594,N_18419);
xor U19003 (N_19003,N_18718,N_18575);
nor U19004 (N_19004,N_18769,N_18677);
nand U19005 (N_19005,N_18729,N_18622);
or U19006 (N_19006,N_18633,N_18721);
nand U19007 (N_19007,N_18530,N_18540);
nand U19008 (N_19008,N_18716,N_18796);
nor U19009 (N_19009,N_18449,N_18610);
or U19010 (N_19010,N_18410,N_18484);
xor U19011 (N_19011,N_18671,N_18715);
nor U19012 (N_19012,N_18466,N_18726);
nor U19013 (N_19013,N_18448,N_18608);
nor U19014 (N_19014,N_18536,N_18432);
nor U19015 (N_19015,N_18529,N_18672);
and U19016 (N_19016,N_18460,N_18614);
xnor U19017 (N_19017,N_18459,N_18471);
or U19018 (N_19018,N_18464,N_18652);
nand U19019 (N_19019,N_18479,N_18494);
nand U19020 (N_19020,N_18649,N_18435);
and U19021 (N_19021,N_18776,N_18763);
nand U19022 (N_19022,N_18729,N_18714);
and U19023 (N_19023,N_18781,N_18694);
nor U19024 (N_19024,N_18631,N_18505);
nand U19025 (N_19025,N_18569,N_18680);
or U19026 (N_19026,N_18619,N_18548);
nor U19027 (N_19027,N_18432,N_18635);
xnor U19028 (N_19028,N_18680,N_18424);
and U19029 (N_19029,N_18711,N_18708);
and U19030 (N_19030,N_18604,N_18524);
nand U19031 (N_19031,N_18551,N_18643);
nand U19032 (N_19032,N_18739,N_18616);
nor U19033 (N_19033,N_18768,N_18537);
nand U19034 (N_19034,N_18401,N_18781);
xor U19035 (N_19035,N_18578,N_18628);
xor U19036 (N_19036,N_18492,N_18453);
and U19037 (N_19037,N_18490,N_18667);
xnor U19038 (N_19038,N_18592,N_18652);
xor U19039 (N_19039,N_18646,N_18534);
nor U19040 (N_19040,N_18657,N_18702);
and U19041 (N_19041,N_18657,N_18685);
nand U19042 (N_19042,N_18561,N_18730);
nand U19043 (N_19043,N_18562,N_18424);
nor U19044 (N_19044,N_18429,N_18510);
or U19045 (N_19045,N_18459,N_18662);
nand U19046 (N_19046,N_18573,N_18659);
nor U19047 (N_19047,N_18498,N_18664);
nand U19048 (N_19048,N_18610,N_18648);
or U19049 (N_19049,N_18742,N_18707);
nor U19050 (N_19050,N_18674,N_18652);
or U19051 (N_19051,N_18671,N_18764);
nand U19052 (N_19052,N_18430,N_18589);
xnor U19053 (N_19053,N_18617,N_18737);
and U19054 (N_19054,N_18726,N_18475);
and U19055 (N_19055,N_18442,N_18591);
and U19056 (N_19056,N_18500,N_18781);
xnor U19057 (N_19057,N_18782,N_18757);
nand U19058 (N_19058,N_18605,N_18724);
xnor U19059 (N_19059,N_18686,N_18563);
xnor U19060 (N_19060,N_18611,N_18771);
nand U19061 (N_19061,N_18440,N_18419);
and U19062 (N_19062,N_18751,N_18638);
nor U19063 (N_19063,N_18673,N_18512);
nand U19064 (N_19064,N_18751,N_18582);
and U19065 (N_19065,N_18789,N_18412);
or U19066 (N_19066,N_18789,N_18488);
nor U19067 (N_19067,N_18704,N_18553);
nor U19068 (N_19068,N_18624,N_18418);
xnor U19069 (N_19069,N_18711,N_18409);
or U19070 (N_19070,N_18518,N_18650);
xor U19071 (N_19071,N_18422,N_18652);
or U19072 (N_19072,N_18504,N_18561);
or U19073 (N_19073,N_18410,N_18457);
nand U19074 (N_19074,N_18524,N_18679);
or U19075 (N_19075,N_18757,N_18588);
nand U19076 (N_19076,N_18774,N_18468);
and U19077 (N_19077,N_18793,N_18596);
or U19078 (N_19078,N_18510,N_18416);
or U19079 (N_19079,N_18769,N_18483);
nor U19080 (N_19080,N_18471,N_18607);
and U19081 (N_19081,N_18453,N_18440);
xor U19082 (N_19082,N_18671,N_18588);
and U19083 (N_19083,N_18797,N_18608);
nor U19084 (N_19084,N_18602,N_18570);
and U19085 (N_19085,N_18684,N_18766);
and U19086 (N_19086,N_18736,N_18653);
or U19087 (N_19087,N_18403,N_18777);
and U19088 (N_19088,N_18457,N_18771);
nor U19089 (N_19089,N_18608,N_18597);
nor U19090 (N_19090,N_18581,N_18457);
xor U19091 (N_19091,N_18707,N_18519);
nor U19092 (N_19092,N_18673,N_18421);
or U19093 (N_19093,N_18429,N_18557);
or U19094 (N_19094,N_18694,N_18735);
xnor U19095 (N_19095,N_18522,N_18498);
nand U19096 (N_19096,N_18428,N_18769);
nor U19097 (N_19097,N_18723,N_18626);
and U19098 (N_19098,N_18448,N_18688);
xnor U19099 (N_19099,N_18563,N_18491);
and U19100 (N_19100,N_18624,N_18404);
nand U19101 (N_19101,N_18562,N_18577);
and U19102 (N_19102,N_18536,N_18754);
xnor U19103 (N_19103,N_18460,N_18751);
xnor U19104 (N_19104,N_18465,N_18557);
nor U19105 (N_19105,N_18616,N_18799);
and U19106 (N_19106,N_18449,N_18591);
xor U19107 (N_19107,N_18630,N_18521);
or U19108 (N_19108,N_18510,N_18463);
nand U19109 (N_19109,N_18654,N_18451);
and U19110 (N_19110,N_18407,N_18683);
xor U19111 (N_19111,N_18683,N_18535);
nor U19112 (N_19112,N_18667,N_18512);
nand U19113 (N_19113,N_18563,N_18775);
or U19114 (N_19114,N_18605,N_18526);
or U19115 (N_19115,N_18755,N_18559);
nand U19116 (N_19116,N_18608,N_18415);
xnor U19117 (N_19117,N_18465,N_18716);
or U19118 (N_19118,N_18768,N_18548);
nand U19119 (N_19119,N_18628,N_18622);
and U19120 (N_19120,N_18593,N_18515);
nand U19121 (N_19121,N_18479,N_18509);
nand U19122 (N_19122,N_18439,N_18462);
and U19123 (N_19123,N_18706,N_18666);
nor U19124 (N_19124,N_18554,N_18765);
nor U19125 (N_19125,N_18755,N_18507);
xnor U19126 (N_19126,N_18435,N_18568);
or U19127 (N_19127,N_18402,N_18420);
or U19128 (N_19128,N_18548,N_18704);
nand U19129 (N_19129,N_18402,N_18687);
xnor U19130 (N_19130,N_18426,N_18662);
nand U19131 (N_19131,N_18661,N_18670);
nand U19132 (N_19132,N_18660,N_18405);
and U19133 (N_19133,N_18457,N_18568);
nor U19134 (N_19134,N_18580,N_18677);
or U19135 (N_19135,N_18572,N_18672);
nor U19136 (N_19136,N_18682,N_18686);
xnor U19137 (N_19137,N_18757,N_18492);
xor U19138 (N_19138,N_18691,N_18537);
and U19139 (N_19139,N_18767,N_18748);
nand U19140 (N_19140,N_18790,N_18462);
or U19141 (N_19141,N_18789,N_18669);
nor U19142 (N_19142,N_18685,N_18454);
and U19143 (N_19143,N_18510,N_18498);
xnor U19144 (N_19144,N_18729,N_18439);
xnor U19145 (N_19145,N_18498,N_18482);
xor U19146 (N_19146,N_18581,N_18566);
or U19147 (N_19147,N_18442,N_18400);
nand U19148 (N_19148,N_18621,N_18655);
nor U19149 (N_19149,N_18748,N_18684);
or U19150 (N_19150,N_18609,N_18744);
nor U19151 (N_19151,N_18453,N_18712);
nor U19152 (N_19152,N_18646,N_18588);
nor U19153 (N_19153,N_18789,N_18506);
nor U19154 (N_19154,N_18707,N_18533);
xnor U19155 (N_19155,N_18555,N_18472);
xor U19156 (N_19156,N_18797,N_18657);
nand U19157 (N_19157,N_18544,N_18630);
or U19158 (N_19158,N_18410,N_18548);
or U19159 (N_19159,N_18736,N_18646);
xor U19160 (N_19160,N_18434,N_18698);
xor U19161 (N_19161,N_18483,N_18551);
xnor U19162 (N_19162,N_18592,N_18424);
and U19163 (N_19163,N_18540,N_18650);
and U19164 (N_19164,N_18684,N_18586);
xnor U19165 (N_19165,N_18439,N_18671);
nand U19166 (N_19166,N_18689,N_18544);
or U19167 (N_19167,N_18639,N_18551);
nand U19168 (N_19168,N_18538,N_18777);
and U19169 (N_19169,N_18693,N_18574);
and U19170 (N_19170,N_18728,N_18643);
or U19171 (N_19171,N_18435,N_18747);
and U19172 (N_19172,N_18587,N_18590);
or U19173 (N_19173,N_18759,N_18709);
nand U19174 (N_19174,N_18670,N_18471);
nor U19175 (N_19175,N_18610,N_18471);
and U19176 (N_19176,N_18400,N_18471);
xor U19177 (N_19177,N_18484,N_18736);
or U19178 (N_19178,N_18644,N_18761);
and U19179 (N_19179,N_18408,N_18512);
nor U19180 (N_19180,N_18698,N_18752);
nor U19181 (N_19181,N_18635,N_18679);
nand U19182 (N_19182,N_18489,N_18755);
nand U19183 (N_19183,N_18598,N_18726);
or U19184 (N_19184,N_18621,N_18726);
nor U19185 (N_19185,N_18533,N_18798);
or U19186 (N_19186,N_18470,N_18717);
xor U19187 (N_19187,N_18791,N_18478);
and U19188 (N_19188,N_18628,N_18433);
xnor U19189 (N_19189,N_18725,N_18615);
nor U19190 (N_19190,N_18427,N_18568);
nand U19191 (N_19191,N_18667,N_18559);
xnor U19192 (N_19192,N_18781,N_18476);
nand U19193 (N_19193,N_18632,N_18576);
nand U19194 (N_19194,N_18584,N_18613);
or U19195 (N_19195,N_18572,N_18462);
nor U19196 (N_19196,N_18790,N_18544);
or U19197 (N_19197,N_18772,N_18745);
or U19198 (N_19198,N_18648,N_18481);
and U19199 (N_19199,N_18649,N_18727);
nand U19200 (N_19200,N_18977,N_18911);
nand U19201 (N_19201,N_19126,N_19104);
and U19202 (N_19202,N_19078,N_19062);
xnor U19203 (N_19203,N_19100,N_18978);
and U19204 (N_19204,N_19158,N_18938);
xnor U19205 (N_19205,N_19005,N_19068);
or U19206 (N_19206,N_18960,N_18934);
xor U19207 (N_19207,N_18948,N_18820);
nand U19208 (N_19208,N_19165,N_18915);
xor U19209 (N_19209,N_19169,N_18933);
xnor U19210 (N_19210,N_18965,N_18821);
nand U19211 (N_19211,N_19040,N_19018);
and U19212 (N_19212,N_18957,N_18877);
nand U19213 (N_19213,N_18861,N_19108);
nand U19214 (N_19214,N_18856,N_19039);
nand U19215 (N_19215,N_19167,N_19138);
nand U19216 (N_19216,N_19008,N_19171);
xnor U19217 (N_19217,N_18912,N_18890);
or U19218 (N_19218,N_19073,N_19007);
and U19219 (N_19219,N_18905,N_19177);
or U19220 (N_19220,N_19127,N_19174);
and U19221 (N_19221,N_19155,N_19082);
or U19222 (N_19222,N_18909,N_19188);
nand U19223 (N_19223,N_18805,N_18967);
or U19224 (N_19224,N_18896,N_19044);
and U19225 (N_19225,N_18963,N_19020);
nand U19226 (N_19226,N_18956,N_19032);
and U19227 (N_19227,N_18832,N_18835);
nand U19228 (N_19228,N_19069,N_19098);
nor U19229 (N_19229,N_18970,N_19016);
xor U19230 (N_19230,N_18989,N_19178);
and U19231 (N_19231,N_19019,N_19148);
nand U19232 (N_19232,N_18959,N_18941);
nand U19233 (N_19233,N_19195,N_19114);
nand U19234 (N_19234,N_18922,N_18863);
or U19235 (N_19235,N_19183,N_18964);
xor U19236 (N_19236,N_18972,N_18897);
xnor U19237 (N_19237,N_18924,N_18853);
nor U19238 (N_19238,N_19197,N_19058);
nand U19239 (N_19239,N_19063,N_19053);
nand U19240 (N_19240,N_19103,N_19000);
nor U19241 (N_19241,N_18873,N_18914);
and U19242 (N_19242,N_19124,N_18810);
and U19243 (N_19243,N_18893,N_19064);
and U19244 (N_19244,N_19006,N_19043);
xor U19245 (N_19245,N_19077,N_18973);
xor U19246 (N_19246,N_19041,N_19050);
nor U19247 (N_19247,N_19164,N_18874);
xor U19248 (N_19248,N_18900,N_18994);
nand U19249 (N_19249,N_19060,N_18871);
xor U19250 (N_19250,N_19031,N_18981);
nand U19251 (N_19251,N_18860,N_19010);
xnor U19252 (N_19252,N_18879,N_19110);
or U19253 (N_19253,N_19087,N_18818);
nand U19254 (N_19254,N_18817,N_19046);
and U19255 (N_19255,N_19091,N_18845);
xor U19256 (N_19256,N_19187,N_19025);
nand U19257 (N_19257,N_18951,N_18840);
nor U19258 (N_19258,N_18991,N_19162);
xnor U19259 (N_19259,N_18867,N_18891);
xor U19260 (N_19260,N_18855,N_19049);
nand U19261 (N_19261,N_19083,N_18906);
and U19262 (N_19262,N_19052,N_19160);
or U19263 (N_19263,N_19115,N_18859);
or U19264 (N_19264,N_19106,N_18878);
nor U19265 (N_19265,N_19189,N_18995);
and U19266 (N_19266,N_19139,N_19185);
and U19267 (N_19267,N_19092,N_19030);
nand U19268 (N_19268,N_18892,N_18904);
or U19269 (N_19269,N_19065,N_18940);
nor U19270 (N_19270,N_18986,N_18823);
xnor U19271 (N_19271,N_18936,N_19140);
nor U19272 (N_19272,N_19094,N_18926);
xor U19273 (N_19273,N_18869,N_19099);
or U19274 (N_19274,N_19081,N_19107);
xnor U19275 (N_19275,N_18819,N_18919);
nand U19276 (N_19276,N_18885,N_18917);
or U19277 (N_19277,N_18827,N_18945);
nand U19278 (N_19278,N_19113,N_19133);
or U19279 (N_19279,N_18982,N_18990);
nand U19280 (N_19280,N_19157,N_18803);
and U19281 (N_19281,N_19128,N_18908);
nor U19282 (N_19282,N_18841,N_19059);
nor U19283 (N_19283,N_19004,N_18851);
and U19284 (N_19284,N_19153,N_19074);
nor U19285 (N_19285,N_18907,N_19036);
and U19286 (N_19286,N_18898,N_18983);
or U19287 (N_19287,N_18999,N_19066);
xnor U19288 (N_19288,N_18932,N_18998);
xnor U19289 (N_19289,N_19003,N_19193);
or U19290 (N_19290,N_18969,N_19037);
nor U19291 (N_19291,N_18954,N_19051);
or U19292 (N_19292,N_18825,N_19180);
nand U19293 (N_19293,N_18889,N_19079);
xor U19294 (N_19294,N_18808,N_19116);
or U19295 (N_19295,N_18918,N_18836);
and U19296 (N_19296,N_18868,N_18833);
nor U19297 (N_19297,N_18947,N_19028);
nand U19298 (N_19298,N_19084,N_18834);
nand U19299 (N_19299,N_19117,N_18946);
nor U19300 (N_19300,N_18801,N_19149);
or U19301 (N_19301,N_19154,N_19194);
nand U19302 (N_19302,N_18826,N_19009);
and U19303 (N_19303,N_19159,N_19191);
or U19304 (N_19304,N_19181,N_19123);
nor U19305 (N_19305,N_18910,N_19150);
nand U19306 (N_19306,N_18958,N_18854);
nand U19307 (N_19307,N_18976,N_18935);
xnor U19308 (N_19308,N_19070,N_18992);
nor U19309 (N_19309,N_19024,N_19146);
and U19310 (N_19310,N_18850,N_18939);
nand U19311 (N_19311,N_19170,N_18997);
nand U19312 (N_19312,N_19125,N_19075);
nor U19313 (N_19313,N_19067,N_19135);
nand U19314 (N_19314,N_18942,N_18987);
or U19315 (N_19315,N_18930,N_18804);
nand U19316 (N_19316,N_18852,N_19002);
or U19317 (N_19317,N_18929,N_19076);
or U19318 (N_19318,N_18949,N_18952);
or U19319 (N_19319,N_18884,N_18846);
nand U19320 (N_19320,N_19111,N_19045);
xnor U19321 (N_19321,N_18802,N_19142);
nor U19322 (N_19322,N_19122,N_19144);
nand U19323 (N_19323,N_19042,N_18858);
nand U19324 (N_19324,N_18928,N_18815);
xor U19325 (N_19325,N_19130,N_18937);
nand U19326 (N_19326,N_18923,N_19119);
xnor U19327 (N_19327,N_19109,N_19012);
and U19328 (N_19328,N_19120,N_18822);
xnor U19329 (N_19329,N_18882,N_18876);
nand U19330 (N_19330,N_19055,N_18872);
nand U19331 (N_19331,N_19179,N_19121);
or U19332 (N_19332,N_19054,N_19132);
and U19333 (N_19333,N_19001,N_19141);
nor U19334 (N_19334,N_19145,N_18988);
xor U19335 (N_19335,N_19021,N_18881);
nor U19336 (N_19336,N_18807,N_19080);
nor U19337 (N_19337,N_18980,N_18849);
nand U19338 (N_19338,N_19026,N_18979);
nor U19339 (N_19339,N_19061,N_19101);
nor U19340 (N_19340,N_18866,N_19112);
xnor U19341 (N_19341,N_18864,N_18894);
or U19342 (N_19342,N_19072,N_19151);
nand U19343 (N_19343,N_19027,N_19152);
and U19344 (N_19344,N_18962,N_18811);
or U19345 (N_19345,N_19017,N_18828);
and U19346 (N_19346,N_18943,N_19192);
nor U19347 (N_19347,N_19047,N_19071);
or U19348 (N_19348,N_19038,N_18812);
and U19349 (N_19349,N_18955,N_18927);
xor U19350 (N_19350,N_19096,N_19168);
nand U19351 (N_19351,N_19057,N_19198);
or U19352 (N_19352,N_19176,N_19090);
nand U19353 (N_19353,N_19011,N_18862);
or U19354 (N_19354,N_19173,N_19190);
or U19355 (N_19355,N_18880,N_18903);
xor U19356 (N_19356,N_18996,N_18839);
xor U19357 (N_19357,N_19035,N_19033);
xnor U19358 (N_19358,N_18824,N_19129);
and U19359 (N_19359,N_19136,N_19097);
and U19360 (N_19360,N_19014,N_19175);
or U19361 (N_19361,N_18895,N_19143);
and U19362 (N_19362,N_18950,N_19134);
nor U19363 (N_19363,N_19093,N_18848);
or U19364 (N_19364,N_18971,N_19199);
nor U19365 (N_19365,N_18842,N_18931);
and U19366 (N_19366,N_18953,N_18993);
nor U19367 (N_19367,N_18844,N_19147);
xor U19368 (N_19368,N_18966,N_18916);
and U19369 (N_19369,N_18975,N_19029);
and U19370 (N_19370,N_18816,N_18837);
nand U19371 (N_19371,N_18857,N_18865);
and U19372 (N_19372,N_19166,N_18875);
or U19373 (N_19373,N_19184,N_19172);
nor U19374 (N_19374,N_19015,N_19089);
or U19375 (N_19375,N_19161,N_18901);
nand U19376 (N_19376,N_18974,N_19186);
xnor U19377 (N_19377,N_18961,N_19182);
nand U19378 (N_19378,N_18829,N_18944);
xnor U19379 (N_19379,N_18984,N_19085);
xor U19380 (N_19380,N_19048,N_18913);
or U19381 (N_19381,N_19086,N_18870);
or U19382 (N_19382,N_19034,N_19013);
and U19383 (N_19383,N_18920,N_19118);
and U19384 (N_19384,N_19137,N_18831);
or U19385 (N_19385,N_18809,N_18888);
xnor U19386 (N_19386,N_18838,N_19023);
nor U19387 (N_19387,N_19056,N_19095);
nand U19388 (N_19388,N_19102,N_18800);
or U19389 (N_19389,N_19131,N_18985);
nor U19390 (N_19390,N_18847,N_18886);
or U19391 (N_19391,N_19156,N_19105);
xnor U19392 (N_19392,N_18921,N_18813);
nand U19393 (N_19393,N_18883,N_19163);
nor U19394 (N_19394,N_18968,N_18887);
nand U19395 (N_19395,N_18843,N_18806);
xor U19396 (N_19396,N_19088,N_18814);
or U19397 (N_19397,N_18830,N_18925);
and U19398 (N_19398,N_18899,N_19196);
nor U19399 (N_19399,N_19022,N_18902);
and U19400 (N_19400,N_18945,N_19019);
xnor U19401 (N_19401,N_18942,N_19015);
and U19402 (N_19402,N_19072,N_18890);
xnor U19403 (N_19403,N_18840,N_18868);
and U19404 (N_19404,N_19154,N_19067);
nand U19405 (N_19405,N_19176,N_18861);
nand U19406 (N_19406,N_19076,N_19103);
and U19407 (N_19407,N_19196,N_18900);
xnor U19408 (N_19408,N_18822,N_19000);
nand U19409 (N_19409,N_18906,N_18881);
and U19410 (N_19410,N_19037,N_19084);
and U19411 (N_19411,N_18922,N_18823);
xor U19412 (N_19412,N_19178,N_18992);
xnor U19413 (N_19413,N_18907,N_19055);
xnor U19414 (N_19414,N_19146,N_18832);
nand U19415 (N_19415,N_19199,N_19186);
and U19416 (N_19416,N_18904,N_18875);
nor U19417 (N_19417,N_18878,N_19035);
nand U19418 (N_19418,N_18895,N_18916);
nand U19419 (N_19419,N_19088,N_18999);
or U19420 (N_19420,N_19003,N_18843);
xor U19421 (N_19421,N_18811,N_19038);
xor U19422 (N_19422,N_19095,N_18975);
and U19423 (N_19423,N_18952,N_18872);
nand U19424 (N_19424,N_18922,N_18841);
nand U19425 (N_19425,N_19085,N_19152);
and U19426 (N_19426,N_19040,N_19071);
nor U19427 (N_19427,N_18850,N_19121);
nor U19428 (N_19428,N_19008,N_18934);
or U19429 (N_19429,N_18935,N_19076);
nor U19430 (N_19430,N_18813,N_18970);
xnor U19431 (N_19431,N_19033,N_19145);
nor U19432 (N_19432,N_18941,N_19005);
xnor U19433 (N_19433,N_19114,N_19199);
or U19434 (N_19434,N_19195,N_18907);
nor U19435 (N_19435,N_18930,N_19175);
or U19436 (N_19436,N_18990,N_19149);
nand U19437 (N_19437,N_18838,N_18902);
and U19438 (N_19438,N_19185,N_19003);
or U19439 (N_19439,N_19119,N_18901);
or U19440 (N_19440,N_18912,N_19095);
nor U19441 (N_19441,N_18864,N_18982);
nor U19442 (N_19442,N_19195,N_19147);
nand U19443 (N_19443,N_18896,N_19168);
nor U19444 (N_19444,N_18841,N_19120);
or U19445 (N_19445,N_18981,N_18937);
nand U19446 (N_19446,N_19164,N_19130);
or U19447 (N_19447,N_18956,N_18951);
nand U19448 (N_19448,N_19156,N_18952);
and U19449 (N_19449,N_19116,N_19026);
nand U19450 (N_19450,N_19125,N_19152);
xnor U19451 (N_19451,N_19092,N_18949);
nand U19452 (N_19452,N_18852,N_19060);
or U19453 (N_19453,N_19070,N_18892);
xor U19454 (N_19454,N_18958,N_19133);
or U19455 (N_19455,N_19106,N_18867);
or U19456 (N_19456,N_19090,N_19041);
nor U19457 (N_19457,N_18812,N_19034);
or U19458 (N_19458,N_19110,N_18876);
or U19459 (N_19459,N_18862,N_18836);
nor U19460 (N_19460,N_18925,N_19105);
xor U19461 (N_19461,N_18848,N_19184);
nor U19462 (N_19462,N_19191,N_18881);
nor U19463 (N_19463,N_18953,N_18845);
or U19464 (N_19464,N_18865,N_19133);
xor U19465 (N_19465,N_19032,N_19170);
nand U19466 (N_19466,N_18883,N_19131);
xnor U19467 (N_19467,N_18890,N_19104);
nor U19468 (N_19468,N_19141,N_18838);
xnor U19469 (N_19469,N_19126,N_19147);
and U19470 (N_19470,N_19195,N_18811);
and U19471 (N_19471,N_18951,N_18929);
nor U19472 (N_19472,N_19010,N_18970);
nand U19473 (N_19473,N_18899,N_18806);
nand U19474 (N_19474,N_19111,N_19081);
nor U19475 (N_19475,N_18855,N_19059);
nand U19476 (N_19476,N_18891,N_18976);
xor U19477 (N_19477,N_19170,N_18981);
or U19478 (N_19478,N_19063,N_18838);
or U19479 (N_19479,N_18934,N_18927);
and U19480 (N_19480,N_19125,N_19002);
xnor U19481 (N_19481,N_18904,N_19150);
or U19482 (N_19482,N_18803,N_18849);
or U19483 (N_19483,N_18800,N_19018);
xor U19484 (N_19484,N_19019,N_18845);
and U19485 (N_19485,N_19187,N_19193);
nor U19486 (N_19486,N_18891,N_18991);
xor U19487 (N_19487,N_19116,N_18843);
nand U19488 (N_19488,N_19160,N_19033);
or U19489 (N_19489,N_19127,N_18814);
and U19490 (N_19490,N_18853,N_19132);
nand U19491 (N_19491,N_18989,N_19115);
nand U19492 (N_19492,N_19070,N_19009);
or U19493 (N_19493,N_18813,N_19095);
xnor U19494 (N_19494,N_18981,N_19128);
xor U19495 (N_19495,N_19047,N_18944);
and U19496 (N_19496,N_18822,N_19153);
or U19497 (N_19497,N_19195,N_19023);
nand U19498 (N_19498,N_19179,N_19161);
or U19499 (N_19499,N_18910,N_19126);
and U19500 (N_19500,N_19144,N_18841);
and U19501 (N_19501,N_19098,N_18896);
and U19502 (N_19502,N_18887,N_18915);
nor U19503 (N_19503,N_18847,N_19059);
nand U19504 (N_19504,N_19152,N_19187);
or U19505 (N_19505,N_19136,N_19028);
or U19506 (N_19506,N_18824,N_19138);
nor U19507 (N_19507,N_18848,N_18816);
and U19508 (N_19508,N_18863,N_18969);
or U19509 (N_19509,N_19082,N_18878);
nor U19510 (N_19510,N_19041,N_19016);
and U19511 (N_19511,N_19027,N_18975);
nand U19512 (N_19512,N_19143,N_19048);
nand U19513 (N_19513,N_19169,N_19195);
nor U19514 (N_19514,N_18920,N_18871);
nand U19515 (N_19515,N_19045,N_18885);
nor U19516 (N_19516,N_18866,N_19063);
xnor U19517 (N_19517,N_19050,N_18975);
nor U19518 (N_19518,N_18985,N_19113);
nand U19519 (N_19519,N_18958,N_18826);
and U19520 (N_19520,N_18948,N_18909);
nand U19521 (N_19521,N_18971,N_18960);
and U19522 (N_19522,N_19064,N_18989);
nand U19523 (N_19523,N_19089,N_18812);
nand U19524 (N_19524,N_19079,N_18993);
xnor U19525 (N_19525,N_19169,N_19051);
and U19526 (N_19526,N_19134,N_19113);
xnor U19527 (N_19527,N_19168,N_19037);
xor U19528 (N_19528,N_18961,N_19004);
xor U19529 (N_19529,N_19079,N_19197);
or U19530 (N_19530,N_19070,N_19043);
xnor U19531 (N_19531,N_19049,N_19041);
nor U19532 (N_19532,N_19076,N_19033);
nand U19533 (N_19533,N_19191,N_19172);
nor U19534 (N_19534,N_18924,N_19145);
xnor U19535 (N_19535,N_18803,N_19087);
or U19536 (N_19536,N_18809,N_18934);
nand U19537 (N_19537,N_19079,N_19146);
nand U19538 (N_19538,N_19011,N_19115);
xor U19539 (N_19539,N_19093,N_18984);
and U19540 (N_19540,N_19083,N_19109);
nand U19541 (N_19541,N_18891,N_19143);
and U19542 (N_19542,N_18934,N_19064);
xnor U19543 (N_19543,N_19150,N_19062);
or U19544 (N_19544,N_19060,N_19165);
and U19545 (N_19545,N_18957,N_19188);
xor U19546 (N_19546,N_19137,N_19033);
or U19547 (N_19547,N_19075,N_18958);
nor U19548 (N_19548,N_18903,N_19084);
nor U19549 (N_19549,N_19058,N_19002);
xor U19550 (N_19550,N_19062,N_18876);
or U19551 (N_19551,N_18998,N_18818);
or U19552 (N_19552,N_18896,N_18884);
or U19553 (N_19553,N_18944,N_19159);
nand U19554 (N_19554,N_19120,N_19127);
and U19555 (N_19555,N_19077,N_19139);
xor U19556 (N_19556,N_18986,N_19019);
and U19557 (N_19557,N_18831,N_18899);
or U19558 (N_19558,N_19083,N_19003);
nor U19559 (N_19559,N_19144,N_18969);
and U19560 (N_19560,N_19186,N_18897);
or U19561 (N_19561,N_19030,N_19021);
nand U19562 (N_19562,N_18807,N_18970);
and U19563 (N_19563,N_18888,N_18913);
nand U19564 (N_19564,N_19142,N_19078);
nor U19565 (N_19565,N_18994,N_19062);
and U19566 (N_19566,N_19051,N_18815);
nor U19567 (N_19567,N_18867,N_18870);
nor U19568 (N_19568,N_18932,N_18978);
xnor U19569 (N_19569,N_19167,N_19112);
nor U19570 (N_19570,N_19195,N_18991);
nor U19571 (N_19571,N_18885,N_18925);
xor U19572 (N_19572,N_19058,N_19116);
and U19573 (N_19573,N_19134,N_19175);
or U19574 (N_19574,N_19133,N_19057);
and U19575 (N_19575,N_19156,N_18821);
or U19576 (N_19576,N_19151,N_18846);
nand U19577 (N_19577,N_18925,N_19162);
nand U19578 (N_19578,N_19095,N_18992);
xnor U19579 (N_19579,N_19193,N_19179);
xor U19580 (N_19580,N_18873,N_18939);
and U19581 (N_19581,N_18802,N_18980);
xor U19582 (N_19582,N_19134,N_19121);
xnor U19583 (N_19583,N_19021,N_19061);
or U19584 (N_19584,N_18910,N_18990);
xnor U19585 (N_19585,N_18910,N_18804);
xnor U19586 (N_19586,N_19038,N_18825);
nand U19587 (N_19587,N_18931,N_19024);
nor U19588 (N_19588,N_19154,N_19050);
or U19589 (N_19589,N_19005,N_18818);
nand U19590 (N_19590,N_19111,N_19085);
nor U19591 (N_19591,N_19139,N_19189);
or U19592 (N_19592,N_19113,N_19067);
xnor U19593 (N_19593,N_18855,N_19075);
xnor U19594 (N_19594,N_19100,N_18876);
xnor U19595 (N_19595,N_18810,N_19114);
nor U19596 (N_19596,N_19035,N_18876);
xnor U19597 (N_19597,N_18933,N_18875);
and U19598 (N_19598,N_18854,N_19190);
xor U19599 (N_19599,N_19014,N_18877);
or U19600 (N_19600,N_19411,N_19386);
and U19601 (N_19601,N_19494,N_19356);
nand U19602 (N_19602,N_19544,N_19400);
xor U19603 (N_19603,N_19585,N_19481);
and U19604 (N_19604,N_19398,N_19428);
nor U19605 (N_19605,N_19422,N_19420);
xor U19606 (N_19606,N_19203,N_19553);
nand U19607 (N_19607,N_19249,N_19449);
nor U19608 (N_19608,N_19247,N_19275);
nand U19609 (N_19609,N_19404,N_19427);
xnor U19610 (N_19610,N_19507,N_19451);
nand U19611 (N_19611,N_19522,N_19321);
nor U19612 (N_19612,N_19573,N_19378);
or U19613 (N_19613,N_19556,N_19220);
or U19614 (N_19614,N_19260,N_19520);
nor U19615 (N_19615,N_19397,N_19468);
or U19616 (N_19616,N_19314,N_19264);
nor U19617 (N_19617,N_19515,N_19228);
and U19618 (N_19618,N_19240,N_19273);
nor U19619 (N_19619,N_19326,N_19571);
nand U19620 (N_19620,N_19509,N_19483);
nand U19621 (N_19621,N_19535,N_19232);
nand U19622 (N_19622,N_19288,N_19435);
nand U19623 (N_19623,N_19452,N_19538);
and U19624 (N_19624,N_19224,N_19338);
and U19625 (N_19625,N_19320,N_19590);
nand U19626 (N_19626,N_19343,N_19396);
xor U19627 (N_19627,N_19230,N_19564);
nand U19628 (N_19628,N_19349,N_19513);
xnor U19629 (N_19629,N_19236,N_19512);
nor U19630 (N_19630,N_19462,N_19209);
nor U19631 (N_19631,N_19225,N_19303);
nand U19632 (N_19632,N_19256,N_19545);
or U19633 (N_19633,N_19293,N_19310);
nand U19634 (N_19634,N_19329,N_19467);
nand U19635 (N_19635,N_19202,N_19279);
or U19636 (N_19636,N_19269,N_19437);
nor U19637 (N_19637,N_19215,N_19252);
nand U19638 (N_19638,N_19237,N_19315);
nor U19639 (N_19639,N_19563,N_19548);
nor U19640 (N_19640,N_19583,N_19339);
and U19641 (N_19641,N_19245,N_19527);
or U19642 (N_19642,N_19489,N_19487);
nor U19643 (N_19643,N_19214,N_19325);
or U19644 (N_19644,N_19376,N_19547);
or U19645 (N_19645,N_19501,N_19204);
or U19646 (N_19646,N_19473,N_19519);
nand U19647 (N_19647,N_19283,N_19503);
nor U19648 (N_19648,N_19351,N_19357);
or U19649 (N_19649,N_19340,N_19381);
and U19650 (N_19650,N_19323,N_19432);
nor U19651 (N_19651,N_19518,N_19348);
xnor U19652 (N_19652,N_19254,N_19524);
and U19653 (N_19653,N_19271,N_19425);
nand U19654 (N_19654,N_19387,N_19354);
and U19655 (N_19655,N_19221,N_19307);
nand U19656 (N_19656,N_19447,N_19346);
nor U19657 (N_19657,N_19484,N_19574);
or U19658 (N_19658,N_19289,N_19317);
and U19659 (N_19659,N_19436,N_19372);
nand U19660 (N_19660,N_19470,N_19559);
nand U19661 (N_19661,N_19294,N_19341);
xor U19662 (N_19662,N_19366,N_19213);
nand U19663 (N_19663,N_19443,N_19312);
and U19664 (N_19664,N_19486,N_19291);
and U19665 (N_19665,N_19448,N_19597);
xor U19666 (N_19666,N_19485,N_19560);
nand U19667 (N_19667,N_19296,N_19408);
or U19668 (N_19668,N_19498,N_19458);
xor U19669 (N_19669,N_19304,N_19227);
or U19670 (N_19670,N_19334,N_19217);
nand U19671 (N_19671,N_19566,N_19586);
nand U19672 (N_19672,N_19385,N_19546);
and U19673 (N_19673,N_19570,N_19444);
nor U19674 (N_19674,N_19445,N_19457);
nor U19675 (N_19675,N_19479,N_19588);
xor U19676 (N_19676,N_19337,N_19375);
nand U19677 (N_19677,N_19584,N_19596);
nor U19678 (N_19678,N_19565,N_19426);
xor U19679 (N_19679,N_19345,N_19270);
nand U19680 (N_19680,N_19592,N_19241);
and U19681 (N_19681,N_19532,N_19305);
xor U19682 (N_19682,N_19402,N_19414);
xor U19683 (N_19683,N_19201,N_19261);
and U19684 (N_19684,N_19322,N_19555);
nand U19685 (N_19685,N_19401,N_19374);
xor U19686 (N_19686,N_19332,N_19405);
nand U19687 (N_19687,N_19311,N_19461);
or U19688 (N_19688,N_19211,N_19355);
and U19689 (N_19689,N_19530,N_19309);
xor U19690 (N_19690,N_19395,N_19529);
or U19691 (N_19691,N_19502,N_19430);
or U19692 (N_19692,N_19222,N_19251);
xnor U19693 (N_19693,N_19336,N_19272);
xnor U19694 (N_19694,N_19300,N_19536);
xnor U19695 (N_19695,N_19281,N_19490);
and U19696 (N_19696,N_19394,N_19301);
xnor U19697 (N_19697,N_19393,N_19233);
xnor U19698 (N_19698,N_19347,N_19576);
or U19699 (N_19699,N_19480,N_19413);
nor U19700 (N_19700,N_19379,N_19558);
or U19701 (N_19701,N_19495,N_19582);
and U19702 (N_19702,N_19516,N_19313);
nand U19703 (N_19703,N_19499,N_19331);
nand U19704 (N_19704,N_19297,N_19239);
xor U19705 (N_19705,N_19364,N_19265);
or U19706 (N_19706,N_19416,N_19223);
and U19707 (N_19707,N_19390,N_19561);
nor U19708 (N_19708,N_19433,N_19243);
or U19709 (N_19709,N_19287,N_19205);
xnor U19710 (N_19710,N_19464,N_19212);
nand U19711 (N_19711,N_19568,N_19333);
xor U19712 (N_19712,N_19500,N_19327);
xnor U19713 (N_19713,N_19308,N_19382);
nor U19714 (N_19714,N_19284,N_19295);
and U19715 (N_19715,N_19302,N_19244);
and U19716 (N_19716,N_19593,N_19504);
xnor U19717 (N_19717,N_19533,N_19362);
nor U19718 (N_19718,N_19591,N_19492);
or U19719 (N_19719,N_19474,N_19580);
or U19720 (N_19720,N_19219,N_19207);
or U19721 (N_19721,N_19440,N_19478);
xnor U19722 (N_19722,N_19497,N_19299);
nor U19723 (N_19723,N_19388,N_19482);
nor U19724 (N_19724,N_19539,N_19350);
nor U19725 (N_19725,N_19517,N_19406);
xnor U19726 (N_19726,N_19208,N_19423);
nand U19727 (N_19727,N_19369,N_19569);
nand U19728 (N_19728,N_19218,N_19292);
nand U19729 (N_19729,N_19344,N_19368);
or U19730 (N_19730,N_19267,N_19463);
xor U19731 (N_19731,N_19456,N_19521);
nand U19732 (N_19732,N_19363,N_19472);
or U19733 (N_19733,N_19598,N_19259);
and U19734 (N_19734,N_19324,N_19419);
xnor U19735 (N_19735,N_19358,N_19442);
xnor U19736 (N_19736,N_19206,N_19216);
nor U19737 (N_19737,N_19526,N_19562);
xor U19738 (N_19738,N_19282,N_19391);
nor U19739 (N_19739,N_19450,N_19231);
nor U19740 (N_19740,N_19431,N_19525);
and U19741 (N_19741,N_19255,N_19438);
nand U19742 (N_19742,N_19274,N_19465);
nor U19743 (N_19743,N_19567,N_19542);
and U19744 (N_19744,N_19412,N_19528);
nor U19745 (N_19745,N_19316,N_19266);
nor U19746 (N_19746,N_19454,N_19534);
or U19747 (N_19747,N_19599,N_19543);
nand U19748 (N_19748,N_19359,N_19429);
xnor U19749 (N_19749,N_19392,N_19410);
and U19750 (N_19750,N_19551,N_19238);
and U19751 (N_19751,N_19491,N_19263);
nor U19752 (N_19752,N_19373,N_19550);
nor U19753 (N_19753,N_19407,N_19549);
and U19754 (N_19754,N_19572,N_19276);
or U19755 (N_19755,N_19441,N_19403);
xor U19756 (N_19756,N_19257,N_19514);
nor U19757 (N_19757,N_19258,N_19421);
nor U19758 (N_19758,N_19476,N_19371);
xor U19759 (N_19759,N_19285,N_19268);
nand U19760 (N_19760,N_19510,N_19577);
xor U19761 (N_19761,N_19234,N_19328);
nor U19762 (N_19762,N_19506,N_19552);
xnor U19763 (N_19763,N_19434,N_19537);
nor U19764 (N_19764,N_19523,N_19242);
xor U19765 (N_19765,N_19466,N_19581);
and U19766 (N_19766,N_19469,N_19511);
nor U19767 (N_19767,N_19280,N_19318);
xnor U19768 (N_19768,N_19578,N_19319);
and U19769 (N_19769,N_19508,N_19541);
nand U19770 (N_19770,N_19384,N_19235);
nand U19771 (N_19771,N_19383,N_19342);
nand U19772 (N_19772,N_19370,N_19594);
or U19773 (N_19773,N_19475,N_19360);
or U19774 (N_19774,N_19496,N_19290);
xnor U19775 (N_19775,N_19587,N_19557);
nor U19776 (N_19776,N_19262,N_19455);
xnor U19777 (N_19777,N_19446,N_19389);
nor U19778 (N_19778,N_19453,N_19417);
or U19779 (N_19779,N_19286,N_19531);
or U19780 (N_19780,N_19253,N_19540);
nand U19781 (N_19781,N_19471,N_19418);
or U19782 (N_19782,N_19459,N_19306);
nand U19783 (N_19783,N_19399,N_19505);
xor U19784 (N_19784,N_19415,N_19298);
xor U19785 (N_19785,N_19589,N_19367);
nor U19786 (N_19786,N_19575,N_19439);
nor U19787 (N_19787,N_19226,N_19352);
xor U19788 (N_19788,N_19409,N_19488);
or U19789 (N_19789,N_19460,N_19377);
nor U19790 (N_19790,N_19579,N_19210);
xnor U19791 (N_19791,N_19250,N_19200);
xor U19792 (N_19792,N_19353,N_19365);
nor U19793 (N_19793,N_19361,N_19477);
xnor U19794 (N_19794,N_19595,N_19277);
and U19795 (N_19795,N_19248,N_19278);
nand U19796 (N_19796,N_19330,N_19380);
xnor U19797 (N_19797,N_19493,N_19554);
nor U19798 (N_19798,N_19229,N_19246);
or U19799 (N_19799,N_19424,N_19335);
or U19800 (N_19800,N_19283,N_19236);
and U19801 (N_19801,N_19208,N_19579);
nor U19802 (N_19802,N_19297,N_19259);
xnor U19803 (N_19803,N_19341,N_19305);
or U19804 (N_19804,N_19427,N_19389);
xnor U19805 (N_19805,N_19502,N_19297);
nand U19806 (N_19806,N_19345,N_19595);
and U19807 (N_19807,N_19377,N_19340);
xnor U19808 (N_19808,N_19233,N_19245);
and U19809 (N_19809,N_19531,N_19420);
and U19810 (N_19810,N_19581,N_19273);
nand U19811 (N_19811,N_19490,N_19565);
and U19812 (N_19812,N_19339,N_19361);
xnor U19813 (N_19813,N_19572,N_19576);
or U19814 (N_19814,N_19575,N_19507);
nor U19815 (N_19815,N_19247,N_19486);
or U19816 (N_19816,N_19381,N_19382);
and U19817 (N_19817,N_19398,N_19207);
and U19818 (N_19818,N_19373,N_19213);
nand U19819 (N_19819,N_19581,N_19479);
or U19820 (N_19820,N_19283,N_19474);
nor U19821 (N_19821,N_19379,N_19362);
nor U19822 (N_19822,N_19566,N_19402);
nand U19823 (N_19823,N_19405,N_19298);
or U19824 (N_19824,N_19486,N_19287);
or U19825 (N_19825,N_19313,N_19565);
and U19826 (N_19826,N_19353,N_19384);
or U19827 (N_19827,N_19436,N_19513);
nand U19828 (N_19828,N_19428,N_19430);
or U19829 (N_19829,N_19490,N_19454);
or U19830 (N_19830,N_19396,N_19389);
nand U19831 (N_19831,N_19471,N_19330);
or U19832 (N_19832,N_19486,N_19592);
nor U19833 (N_19833,N_19567,N_19583);
or U19834 (N_19834,N_19203,N_19520);
nand U19835 (N_19835,N_19320,N_19345);
nor U19836 (N_19836,N_19414,N_19283);
xnor U19837 (N_19837,N_19428,N_19578);
xnor U19838 (N_19838,N_19416,N_19527);
nor U19839 (N_19839,N_19580,N_19297);
nand U19840 (N_19840,N_19543,N_19569);
xnor U19841 (N_19841,N_19220,N_19303);
xnor U19842 (N_19842,N_19260,N_19213);
xnor U19843 (N_19843,N_19261,N_19408);
nor U19844 (N_19844,N_19241,N_19569);
xor U19845 (N_19845,N_19487,N_19431);
xnor U19846 (N_19846,N_19599,N_19472);
nor U19847 (N_19847,N_19508,N_19269);
or U19848 (N_19848,N_19356,N_19238);
or U19849 (N_19849,N_19492,N_19262);
xor U19850 (N_19850,N_19559,N_19442);
or U19851 (N_19851,N_19353,N_19203);
xor U19852 (N_19852,N_19533,N_19491);
nand U19853 (N_19853,N_19545,N_19499);
or U19854 (N_19854,N_19252,N_19517);
xor U19855 (N_19855,N_19545,N_19380);
nand U19856 (N_19856,N_19368,N_19573);
or U19857 (N_19857,N_19260,N_19478);
xnor U19858 (N_19858,N_19382,N_19203);
xnor U19859 (N_19859,N_19204,N_19219);
or U19860 (N_19860,N_19344,N_19534);
nand U19861 (N_19861,N_19503,N_19308);
and U19862 (N_19862,N_19401,N_19311);
or U19863 (N_19863,N_19309,N_19364);
or U19864 (N_19864,N_19276,N_19496);
or U19865 (N_19865,N_19369,N_19531);
nand U19866 (N_19866,N_19414,N_19451);
and U19867 (N_19867,N_19286,N_19550);
nand U19868 (N_19868,N_19557,N_19323);
nor U19869 (N_19869,N_19539,N_19514);
or U19870 (N_19870,N_19327,N_19202);
and U19871 (N_19871,N_19362,N_19339);
or U19872 (N_19872,N_19539,N_19526);
nand U19873 (N_19873,N_19482,N_19533);
nand U19874 (N_19874,N_19451,N_19268);
xnor U19875 (N_19875,N_19392,N_19384);
and U19876 (N_19876,N_19436,N_19540);
nand U19877 (N_19877,N_19337,N_19211);
nand U19878 (N_19878,N_19575,N_19416);
nor U19879 (N_19879,N_19316,N_19557);
xor U19880 (N_19880,N_19267,N_19217);
and U19881 (N_19881,N_19335,N_19238);
or U19882 (N_19882,N_19410,N_19333);
and U19883 (N_19883,N_19537,N_19532);
nor U19884 (N_19884,N_19494,N_19484);
or U19885 (N_19885,N_19590,N_19296);
nor U19886 (N_19886,N_19276,N_19232);
xor U19887 (N_19887,N_19564,N_19344);
nor U19888 (N_19888,N_19301,N_19586);
nand U19889 (N_19889,N_19402,N_19515);
nor U19890 (N_19890,N_19354,N_19514);
nor U19891 (N_19891,N_19523,N_19454);
and U19892 (N_19892,N_19221,N_19596);
nor U19893 (N_19893,N_19570,N_19201);
and U19894 (N_19894,N_19498,N_19345);
and U19895 (N_19895,N_19594,N_19298);
and U19896 (N_19896,N_19312,N_19264);
or U19897 (N_19897,N_19489,N_19269);
and U19898 (N_19898,N_19466,N_19479);
xor U19899 (N_19899,N_19426,N_19227);
and U19900 (N_19900,N_19332,N_19269);
xnor U19901 (N_19901,N_19277,N_19311);
and U19902 (N_19902,N_19412,N_19595);
nand U19903 (N_19903,N_19516,N_19382);
and U19904 (N_19904,N_19247,N_19439);
nand U19905 (N_19905,N_19414,N_19326);
xnor U19906 (N_19906,N_19278,N_19531);
xor U19907 (N_19907,N_19595,N_19419);
or U19908 (N_19908,N_19474,N_19482);
or U19909 (N_19909,N_19304,N_19585);
nor U19910 (N_19910,N_19514,N_19223);
and U19911 (N_19911,N_19592,N_19320);
nand U19912 (N_19912,N_19544,N_19387);
nand U19913 (N_19913,N_19239,N_19375);
and U19914 (N_19914,N_19496,N_19503);
nor U19915 (N_19915,N_19529,N_19212);
and U19916 (N_19916,N_19485,N_19463);
nand U19917 (N_19917,N_19227,N_19332);
xor U19918 (N_19918,N_19387,N_19589);
nor U19919 (N_19919,N_19358,N_19360);
or U19920 (N_19920,N_19297,N_19493);
xnor U19921 (N_19921,N_19537,N_19349);
nor U19922 (N_19922,N_19378,N_19287);
xor U19923 (N_19923,N_19564,N_19513);
nand U19924 (N_19924,N_19212,N_19368);
or U19925 (N_19925,N_19227,N_19298);
nand U19926 (N_19926,N_19370,N_19520);
or U19927 (N_19927,N_19461,N_19309);
or U19928 (N_19928,N_19542,N_19400);
xnor U19929 (N_19929,N_19477,N_19412);
nand U19930 (N_19930,N_19327,N_19501);
nand U19931 (N_19931,N_19301,N_19592);
xnor U19932 (N_19932,N_19353,N_19579);
nand U19933 (N_19933,N_19469,N_19328);
nor U19934 (N_19934,N_19356,N_19410);
or U19935 (N_19935,N_19328,N_19323);
or U19936 (N_19936,N_19205,N_19360);
nor U19937 (N_19937,N_19589,N_19507);
xor U19938 (N_19938,N_19396,N_19230);
nand U19939 (N_19939,N_19247,N_19341);
nand U19940 (N_19940,N_19211,N_19231);
nor U19941 (N_19941,N_19375,N_19302);
and U19942 (N_19942,N_19344,N_19269);
nand U19943 (N_19943,N_19541,N_19564);
and U19944 (N_19944,N_19392,N_19553);
nor U19945 (N_19945,N_19583,N_19563);
xor U19946 (N_19946,N_19342,N_19244);
or U19947 (N_19947,N_19370,N_19200);
and U19948 (N_19948,N_19425,N_19383);
nor U19949 (N_19949,N_19534,N_19499);
or U19950 (N_19950,N_19272,N_19405);
nor U19951 (N_19951,N_19309,N_19418);
or U19952 (N_19952,N_19524,N_19563);
nor U19953 (N_19953,N_19594,N_19486);
nor U19954 (N_19954,N_19344,N_19509);
xnor U19955 (N_19955,N_19598,N_19468);
xor U19956 (N_19956,N_19558,N_19551);
or U19957 (N_19957,N_19430,N_19269);
and U19958 (N_19958,N_19264,N_19233);
nand U19959 (N_19959,N_19207,N_19419);
or U19960 (N_19960,N_19306,N_19494);
or U19961 (N_19961,N_19425,N_19468);
and U19962 (N_19962,N_19554,N_19367);
nand U19963 (N_19963,N_19221,N_19594);
and U19964 (N_19964,N_19205,N_19535);
nor U19965 (N_19965,N_19459,N_19218);
nor U19966 (N_19966,N_19292,N_19421);
nand U19967 (N_19967,N_19379,N_19270);
xor U19968 (N_19968,N_19459,N_19437);
or U19969 (N_19969,N_19550,N_19442);
nor U19970 (N_19970,N_19535,N_19362);
or U19971 (N_19971,N_19466,N_19307);
nand U19972 (N_19972,N_19230,N_19546);
xnor U19973 (N_19973,N_19277,N_19280);
and U19974 (N_19974,N_19241,N_19577);
nor U19975 (N_19975,N_19282,N_19525);
and U19976 (N_19976,N_19577,N_19225);
or U19977 (N_19977,N_19302,N_19397);
xnor U19978 (N_19978,N_19296,N_19270);
nand U19979 (N_19979,N_19480,N_19367);
and U19980 (N_19980,N_19556,N_19512);
nor U19981 (N_19981,N_19391,N_19477);
xnor U19982 (N_19982,N_19381,N_19542);
nand U19983 (N_19983,N_19376,N_19425);
and U19984 (N_19984,N_19303,N_19488);
and U19985 (N_19985,N_19510,N_19459);
or U19986 (N_19986,N_19548,N_19333);
xor U19987 (N_19987,N_19470,N_19448);
nand U19988 (N_19988,N_19202,N_19490);
xor U19989 (N_19989,N_19311,N_19534);
xor U19990 (N_19990,N_19531,N_19347);
nand U19991 (N_19991,N_19372,N_19458);
and U19992 (N_19992,N_19466,N_19287);
nand U19993 (N_19993,N_19456,N_19225);
or U19994 (N_19994,N_19421,N_19270);
nand U19995 (N_19995,N_19490,N_19343);
and U19996 (N_19996,N_19332,N_19316);
or U19997 (N_19997,N_19527,N_19270);
nand U19998 (N_19998,N_19347,N_19234);
or U19999 (N_19999,N_19534,N_19238);
xnor UO_0 (O_0,N_19977,N_19932);
xnor UO_1 (O_1,N_19879,N_19781);
nor UO_2 (O_2,N_19975,N_19695);
or UO_3 (O_3,N_19682,N_19804);
nor UO_4 (O_4,N_19883,N_19807);
nor UO_5 (O_5,N_19637,N_19618);
and UO_6 (O_6,N_19736,N_19826);
or UO_7 (O_7,N_19706,N_19945);
and UO_8 (O_8,N_19741,N_19727);
nor UO_9 (O_9,N_19800,N_19904);
nand UO_10 (O_10,N_19663,N_19942);
nand UO_11 (O_11,N_19978,N_19992);
nand UO_12 (O_12,N_19656,N_19608);
nand UO_13 (O_13,N_19995,N_19858);
or UO_14 (O_14,N_19615,N_19888);
nand UO_15 (O_15,N_19642,N_19960);
nor UO_16 (O_16,N_19782,N_19653);
and UO_17 (O_17,N_19770,N_19696);
nand UO_18 (O_18,N_19668,N_19863);
or UO_19 (O_19,N_19751,N_19735);
or UO_20 (O_20,N_19830,N_19646);
xor UO_21 (O_21,N_19929,N_19843);
and UO_22 (O_22,N_19723,N_19624);
nand UO_23 (O_23,N_19725,N_19604);
or UO_24 (O_24,N_19925,N_19897);
nand UO_25 (O_25,N_19930,N_19916);
xor UO_26 (O_26,N_19705,N_19625);
nor UO_27 (O_27,N_19760,N_19822);
xor UO_28 (O_28,N_19794,N_19733);
and UO_29 (O_29,N_19892,N_19693);
nor UO_30 (O_30,N_19600,N_19640);
xor UO_31 (O_31,N_19886,N_19674);
nand UO_32 (O_32,N_19748,N_19805);
and UO_33 (O_33,N_19610,N_19685);
or UO_34 (O_34,N_19710,N_19711);
nand UO_35 (O_35,N_19671,N_19780);
or UO_36 (O_36,N_19766,N_19660);
or UO_37 (O_37,N_19670,N_19881);
xor UO_38 (O_38,N_19820,N_19810);
nand UO_39 (O_39,N_19729,N_19678);
or UO_40 (O_40,N_19988,N_19935);
nor UO_41 (O_41,N_19687,N_19971);
nor UO_42 (O_42,N_19914,N_19801);
or UO_43 (O_43,N_19823,N_19737);
xor UO_44 (O_44,N_19908,N_19722);
xnor UO_45 (O_45,N_19901,N_19745);
nor UO_46 (O_46,N_19959,N_19601);
nand UO_47 (O_47,N_19899,N_19814);
and UO_48 (O_48,N_19979,N_19708);
nor UO_49 (O_49,N_19652,N_19633);
nand UO_50 (O_50,N_19967,N_19755);
xor UO_51 (O_51,N_19949,N_19752);
nand UO_52 (O_52,N_19815,N_19709);
nand UO_53 (O_53,N_19628,N_19836);
nand UO_54 (O_54,N_19641,N_19769);
xor UO_55 (O_55,N_19746,N_19956);
and UO_56 (O_56,N_19655,N_19811);
or UO_57 (O_57,N_19664,N_19626);
nor UO_58 (O_58,N_19789,N_19889);
xnor UO_59 (O_59,N_19684,N_19764);
nor UO_60 (O_60,N_19784,N_19884);
nor UO_61 (O_61,N_19944,N_19720);
and UO_62 (O_62,N_19985,N_19790);
xnor UO_63 (O_63,N_19661,N_19919);
xor UO_64 (O_64,N_19703,N_19953);
nor UO_65 (O_65,N_19767,N_19990);
and UO_66 (O_66,N_19976,N_19906);
or UO_67 (O_67,N_19856,N_19861);
nor UO_68 (O_68,N_19832,N_19970);
and UO_69 (O_69,N_19827,N_19749);
or UO_70 (O_70,N_19650,N_19845);
and UO_71 (O_71,N_19799,N_19756);
nor UO_72 (O_72,N_19852,N_19905);
xnor UO_73 (O_73,N_19715,N_19707);
or UO_74 (O_74,N_19818,N_19853);
and UO_75 (O_75,N_19817,N_19923);
nand UO_76 (O_76,N_19623,N_19659);
nand UO_77 (O_77,N_19651,N_19885);
and UO_78 (O_78,N_19982,N_19997);
xnor UO_79 (O_79,N_19986,N_19834);
and UO_80 (O_80,N_19855,N_19948);
or UO_81 (O_81,N_19957,N_19658);
xor UO_82 (O_82,N_19833,N_19849);
xor UO_83 (O_83,N_19964,N_19648);
or UO_84 (O_84,N_19851,N_19808);
or UO_85 (O_85,N_19828,N_19943);
xor UO_86 (O_86,N_19732,N_19819);
nand UO_87 (O_87,N_19803,N_19854);
xor UO_88 (O_88,N_19873,N_19621);
and UO_89 (O_89,N_19968,N_19972);
or UO_90 (O_90,N_19680,N_19759);
and UO_91 (O_91,N_19643,N_19765);
nor UO_92 (O_92,N_19872,N_19974);
and UO_93 (O_93,N_19900,N_19644);
nor UO_94 (O_94,N_19719,N_19910);
nor UO_95 (O_95,N_19848,N_19862);
nand UO_96 (O_96,N_19816,N_19902);
nor UO_97 (O_97,N_19688,N_19950);
or UO_98 (O_98,N_19981,N_19859);
and UO_99 (O_99,N_19645,N_19860);
nand UO_100 (O_100,N_19934,N_19742);
xor UO_101 (O_101,N_19697,N_19619);
nand UO_102 (O_102,N_19809,N_19931);
nor UO_103 (O_103,N_19679,N_19913);
nor UO_104 (O_104,N_19896,N_19840);
and UO_105 (O_105,N_19673,N_19864);
and UO_106 (O_106,N_19771,N_19839);
nand UO_107 (O_107,N_19890,N_19993);
or UO_108 (O_108,N_19724,N_19714);
nor UO_109 (O_109,N_19795,N_19717);
xor UO_110 (O_110,N_19947,N_19675);
xnor UO_111 (O_111,N_19639,N_19969);
xnor UO_112 (O_112,N_19785,N_19987);
and UO_113 (O_113,N_19605,N_19607);
nand UO_114 (O_114,N_19991,N_19824);
or UO_115 (O_115,N_19692,N_19683);
and UO_116 (O_116,N_19937,N_19716);
and UO_117 (O_117,N_19747,N_19734);
and UO_118 (O_118,N_19691,N_19617);
nor UO_119 (O_119,N_19676,N_19880);
xnor UO_120 (O_120,N_19891,N_19689);
or UO_121 (O_121,N_19787,N_19939);
or UO_122 (O_122,N_19926,N_19783);
nand UO_123 (O_123,N_19632,N_19850);
or UO_124 (O_124,N_19893,N_19806);
nor UO_125 (O_125,N_19768,N_19966);
nand UO_126 (O_126,N_19775,N_19793);
or UO_127 (O_127,N_19999,N_19686);
or UO_128 (O_128,N_19779,N_19989);
nand UO_129 (O_129,N_19772,N_19665);
nand UO_130 (O_130,N_19928,N_19667);
nor UO_131 (O_131,N_19718,N_19763);
xor UO_132 (O_132,N_19699,N_19857);
or UO_133 (O_133,N_19761,N_19955);
nor UO_134 (O_134,N_19704,N_19980);
nor UO_135 (O_135,N_19915,N_19941);
or UO_136 (O_136,N_19662,N_19887);
or UO_137 (O_137,N_19954,N_19630);
nand UO_138 (O_138,N_19868,N_19831);
or UO_139 (O_139,N_19962,N_19698);
and UO_140 (O_140,N_19757,N_19702);
nor UO_141 (O_141,N_19796,N_19701);
nand UO_142 (O_142,N_19998,N_19754);
nor UO_143 (O_143,N_19921,N_19825);
or UO_144 (O_144,N_19917,N_19774);
xnor UO_145 (O_145,N_19627,N_19614);
and UO_146 (O_146,N_19963,N_19791);
nand UO_147 (O_147,N_19842,N_19813);
or UO_148 (O_148,N_19762,N_19984);
nor UO_149 (O_149,N_19797,N_19920);
or UO_150 (O_150,N_19635,N_19638);
and UO_151 (O_151,N_19933,N_19983);
and UO_152 (O_152,N_19753,N_19609);
or UO_153 (O_153,N_19778,N_19835);
and UO_154 (O_154,N_19750,N_19788);
or UO_155 (O_155,N_19631,N_19792);
xor UO_156 (O_156,N_19867,N_19922);
or UO_157 (O_157,N_19713,N_19620);
or UO_158 (O_158,N_19629,N_19654);
nand UO_159 (O_159,N_19712,N_19829);
or UO_160 (O_160,N_19647,N_19669);
nor UO_161 (O_161,N_19951,N_19878);
nor UO_162 (O_162,N_19602,N_19838);
nor UO_163 (O_163,N_19903,N_19773);
nand UO_164 (O_164,N_19907,N_19690);
nand UO_165 (O_165,N_19847,N_19649);
xor UO_166 (O_166,N_19739,N_19961);
or UO_167 (O_167,N_19865,N_19681);
nand UO_168 (O_168,N_19877,N_19996);
nor UO_169 (O_169,N_19924,N_19728);
nor UO_170 (O_170,N_19634,N_19870);
xnor UO_171 (O_171,N_19731,N_19694);
nand UO_172 (O_172,N_19958,N_19613);
nor UO_173 (O_173,N_19776,N_19821);
and UO_174 (O_174,N_19918,N_19612);
and UO_175 (O_175,N_19895,N_19940);
xnor UO_176 (O_176,N_19841,N_19927);
nor UO_177 (O_177,N_19666,N_19952);
xor UO_178 (O_178,N_19812,N_19657);
nand UO_179 (O_179,N_19874,N_19758);
nor UO_180 (O_180,N_19622,N_19911);
nand UO_181 (O_181,N_19837,N_19938);
xnor UO_182 (O_182,N_19973,N_19740);
nand UO_183 (O_183,N_19677,N_19898);
xnor UO_184 (O_184,N_19871,N_19616);
nor UO_185 (O_185,N_19700,N_19606);
and UO_186 (O_186,N_19744,N_19994);
nand UO_187 (O_187,N_19721,N_19802);
and UO_188 (O_188,N_19786,N_19603);
xnor UO_189 (O_189,N_19946,N_19798);
or UO_190 (O_190,N_19875,N_19912);
nand UO_191 (O_191,N_19866,N_19730);
and UO_192 (O_192,N_19738,N_19726);
or UO_193 (O_193,N_19876,N_19611);
and UO_194 (O_194,N_19672,N_19846);
xor UO_195 (O_195,N_19965,N_19743);
nand UO_196 (O_196,N_19909,N_19869);
xor UO_197 (O_197,N_19777,N_19882);
xor UO_198 (O_198,N_19636,N_19894);
or UO_199 (O_199,N_19844,N_19936);
nand UO_200 (O_200,N_19945,N_19815);
nor UO_201 (O_201,N_19628,N_19665);
or UO_202 (O_202,N_19941,N_19604);
xnor UO_203 (O_203,N_19912,N_19893);
or UO_204 (O_204,N_19872,N_19887);
xor UO_205 (O_205,N_19772,N_19675);
and UO_206 (O_206,N_19912,N_19622);
xor UO_207 (O_207,N_19926,N_19706);
nor UO_208 (O_208,N_19823,N_19837);
and UO_209 (O_209,N_19730,N_19616);
nand UO_210 (O_210,N_19648,N_19697);
nor UO_211 (O_211,N_19976,N_19885);
xor UO_212 (O_212,N_19742,N_19608);
or UO_213 (O_213,N_19667,N_19802);
and UO_214 (O_214,N_19984,N_19684);
and UO_215 (O_215,N_19894,N_19929);
nand UO_216 (O_216,N_19742,N_19785);
xor UO_217 (O_217,N_19796,N_19782);
and UO_218 (O_218,N_19791,N_19685);
xor UO_219 (O_219,N_19784,N_19822);
or UO_220 (O_220,N_19876,N_19999);
nand UO_221 (O_221,N_19754,N_19926);
nor UO_222 (O_222,N_19737,N_19871);
xor UO_223 (O_223,N_19624,N_19812);
or UO_224 (O_224,N_19746,N_19738);
nand UO_225 (O_225,N_19990,N_19696);
and UO_226 (O_226,N_19913,N_19699);
or UO_227 (O_227,N_19829,N_19961);
nand UO_228 (O_228,N_19734,N_19832);
or UO_229 (O_229,N_19973,N_19753);
and UO_230 (O_230,N_19764,N_19674);
or UO_231 (O_231,N_19779,N_19637);
xnor UO_232 (O_232,N_19894,N_19957);
or UO_233 (O_233,N_19878,N_19766);
nand UO_234 (O_234,N_19631,N_19808);
or UO_235 (O_235,N_19884,N_19690);
or UO_236 (O_236,N_19851,N_19883);
and UO_237 (O_237,N_19952,N_19932);
nor UO_238 (O_238,N_19806,N_19957);
nor UO_239 (O_239,N_19828,N_19991);
xnor UO_240 (O_240,N_19918,N_19702);
xnor UO_241 (O_241,N_19804,N_19866);
nand UO_242 (O_242,N_19718,N_19924);
xor UO_243 (O_243,N_19801,N_19887);
and UO_244 (O_244,N_19943,N_19623);
nor UO_245 (O_245,N_19843,N_19739);
and UO_246 (O_246,N_19786,N_19667);
and UO_247 (O_247,N_19939,N_19727);
and UO_248 (O_248,N_19788,N_19863);
or UO_249 (O_249,N_19622,N_19767);
or UO_250 (O_250,N_19771,N_19952);
or UO_251 (O_251,N_19606,N_19722);
and UO_252 (O_252,N_19921,N_19624);
xnor UO_253 (O_253,N_19985,N_19891);
xnor UO_254 (O_254,N_19613,N_19803);
and UO_255 (O_255,N_19932,N_19785);
nor UO_256 (O_256,N_19737,N_19757);
nand UO_257 (O_257,N_19721,N_19853);
nand UO_258 (O_258,N_19927,N_19975);
nor UO_259 (O_259,N_19990,N_19956);
xnor UO_260 (O_260,N_19656,N_19753);
nor UO_261 (O_261,N_19638,N_19787);
or UO_262 (O_262,N_19961,N_19864);
and UO_263 (O_263,N_19724,N_19705);
nor UO_264 (O_264,N_19883,N_19872);
and UO_265 (O_265,N_19912,N_19923);
xor UO_266 (O_266,N_19733,N_19717);
xnor UO_267 (O_267,N_19874,N_19848);
nand UO_268 (O_268,N_19963,N_19945);
and UO_269 (O_269,N_19712,N_19701);
xnor UO_270 (O_270,N_19714,N_19972);
and UO_271 (O_271,N_19679,N_19701);
xnor UO_272 (O_272,N_19901,N_19752);
xnor UO_273 (O_273,N_19926,N_19998);
xnor UO_274 (O_274,N_19698,N_19785);
xor UO_275 (O_275,N_19993,N_19702);
or UO_276 (O_276,N_19883,N_19712);
and UO_277 (O_277,N_19847,N_19850);
or UO_278 (O_278,N_19684,N_19986);
nand UO_279 (O_279,N_19720,N_19876);
and UO_280 (O_280,N_19740,N_19772);
nand UO_281 (O_281,N_19917,N_19648);
and UO_282 (O_282,N_19953,N_19968);
and UO_283 (O_283,N_19974,N_19859);
nor UO_284 (O_284,N_19948,N_19814);
xor UO_285 (O_285,N_19908,N_19775);
xor UO_286 (O_286,N_19790,N_19762);
xnor UO_287 (O_287,N_19753,N_19635);
nand UO_288 (O_288,N_19737,N_19842);
xor UO_289 (O_289,N_19755,N_19650);
or UO_290 (O_290,N_19843,N_19663);
and UO_291 (O_291,N_19823,N_19754);
nor UO_292 (O_292,N_19823,N_19995);
nor UO_293 (O_293,N_19793,N_19988);
nor UO_294 (O_294,N_19621,N_19712);
nor UO_295 (O_295,N_19645,N_19965);
and UO_296 (O_296,N_19983,N_19858);
and UO_297 (O_297,N_19908,N_19988);
or UO_298 (O_298,N_19807,N_19610);
or UO_299 (O_299,N_19959,N_19685);
and UO_300 (O_300,N_19735,N_19848);
xor UO_301 (O_301,N_19915,N_19923);
xnor UO_302 (O_302,N_19878,N_19707);
or UO_303 (O_303,N_19930,N_19850);
nand UO_304 (O_304,N_19969,N_19954);
xor UO_305 (O_305,N_19806,N_19775);
xor UO_306 (O_306,N_19617,N_19651);
nand UO_307 (O_307,N_19875,N_19782);
nand UO_308 (O_308,N_19760,N_19640);
or UO_309 (O_309,N_19658,N_19683);
xnor UO_310 (O_310,N_19803,N_19797);
nor UO_311 (O_311,N_19798,N_19792);
xnor UO_312 (O_312,N_19877,N_19739);
or UO_313 (O_313,N_19939,N_19854);
xnor UO_314 (O_314,N_19818,N_19806);
xor UO_315 (O_315,N_19650,N_19617);
xnor UO_316 (O_316,N_19622,N_19999);
nor UO_317 (O_317,N_19744,N_19627);
or UO_318 (O_318,N_19721,N_19914);
nand UO_319 (O_319,N_19739,N_19829);
and UO_320 (O_320,N_19912,N_19840);
nand UO_321 (O_321,N_19781,N_19888);
nor UO_322 (O_322,N_19802,N_19770);
xor UO_323 (O_323,N_19935,N_19784);
or UO_324 (O_324,N_19953,N_19990);
nand UO_325 (O_325,N_19658,N_19920);
or UO_326 (O_326,N_19655,N_19601);
nor UO_327 (O_327,N_19676,N_19767);
xnor UO_328 (O_328,N_19748,N_19759);
and UO_329 (O_329,N_19788,N_19847);
nand UO_330 (O_330,N_19963,N_19770);
and UO_331 (O_331,N_19780,N_19934);
and UO_332 (O_332,N_19686,N_19933);
xor UO_333 (O_333,N_19783,N_19827);
xor UO_334 (O_334,N_19913,N_19773);
nor UO_335 (O_335,N_19920,N_19861);
or UO_336 (O_336,N_19867,N_19713);
nor UO_337 (O_337,N_19984,N_19894);
xnor UO_338 (O_338,N_19916,N_19857);
nor UO_339 (O_339,N_19684,N_19921);
xnor UO_340 (O_340,N_19652,N_19816);
nor UO_341 (O_341,N_19740,N_19709);
or UO_342 (O_342,N_19812,N_19794);
and UO_343 (O_343,N_19684,N_19928);
or UO_344 (O_344,N_19750,N_19945);
or UO_345 (O_345,N_19690,N_19867);
or UO_346 (O_346,N_19621,N_19791);
or UO_347 (O_347,N_19629,N_19847);
xnor UO_348 (O_348,N_19614,N_19761);
and UO_349 (O_349,N_19700,N_19737);
nor UO_350 (O_350,N_19705,N_19846);
and UO_351 (O_351,N_19671,N_19675);
and UO_352 (O_352,N_19735,N_19736);
xor UO_353 (O_353,N_19990,N_19949);
and UO_354 (O_354,N_19966,N_19824);
xor UO_355 (O_355,N_19769,N_19778);
or UO_356 (O_356,N_19941,N_19614);
nand UO_357 (O_357,N_19646,N_19846);
nand UO_358 (O_358,N_19667,N_19902);
and UO_359 (O_359,N_19878,N_19998);
nor UO_360 (O_360,N_19998,N_19741);
or UO_361 (O_361,N_19665,N_19982);
xor UO_362 (O_362,N_19999,N_19767);
or UO_363 (O_363,N_19931,N_19912);
and UO_364 (O_364,N_19829,N_19727);
xnor UO_365 (O_365,N_19635,N_19734);
or UO_366 (O_366,N_19845,N_19963);
nand UO_367 (O_367,N_19727,N_19811);
xnor UO_368 (O_368,N_19802,N_19856);
nor UO_369 (O_369,N_19696,N_19700);
nand UO_370 (O_370,N_19816,N_19683);
nor UO_371 (O_371,N_19884,N_19911);
xnor UO_372 (O_372,N_19672,N_19870);
xnor UO_373 (O_373,N_19831,N_19900);
xor UO_374 (O_374,N_19717,N_19649);
nor UO_375 (O_375,N_19886,N_19885);
xnor UO_376 (O_376,N_19955,N_19964);
or UO_377 (O_377,N_19932,N_19766);
xor UO_378 (O_378,N_19950,N_19762);
or UO_379 (O_379,N_19964,N_19920);
nand UO_380 (O_380,N_19939,N_19658);
xnor UO_381 (O_381,N_19947,N_19873);
nand UO_382 (O_382,N_19997,N_19900);
and UO_383 (O_383,N_19666,N_19619);
and UO_384 (O_384,N_19818,N_19956);
and UO_385 (O_385,N_19693,N_19880);
nand UO_386 (O_386,N_19683,N_19906);
xor UO_387 (O_387,N_19851,N_19944);
nand UO_388 (O_388,N_19881,N_19672);
nor UO_389 (O_389,N_19770,N_19726);
nor UO_390 (O_390,N_19659,N_19942);
nor UO_391 (O_391,N_19928,N_19975);
and UO_392 (O_392,N_19674,N_19852);
or UO_393 (O_393,N_19840,N_19699);
nand UO_394 (O_394,N_19687,N_19676);
nand UO_395 (O_395,N_19867,N_19824);
xnor UO_396 (O_396,N_19726,N_19640);
and UO_397 (O_397,N_19790,N_19992);
or UO_398 (O_398,N_19732,N_19963);
or UO_399 (O_399,N_19842,N_19613);
and UO_400 (O_400,N_19764,N_19819);
xor UO_401 (O_401,N_19974,N_19790);
or UO_402 (O_402,N_19963,N_19985);
or UO_403 (O_403,N_19901,N_19668);
nor UO_404 (O_404,N_19858,N_19963);
or UO_405 (O_405,N_19818,N_19994);
and UO_406 (O_406,N_19662,N_19894);
nand UO_407 (O_407,N_19844,N_19627);
nand UO_408 (O_408,N_19856,N_19913);
or UO_409 (O_409,N_19751,N_19765);
xor UO_410 (O_410,N_19963,N_19673);
and UO_411 (O_411,N_19945,N_19755);
xnor UO_412 (O_412,N_19797,N_19716);
xor UO_413 (O_413,N_19643,N_19959);
xnor UO_414 (O_414,N_19987,N_19702);
nor UO_415 (O_415,N_19908,N_19842);
nor UO_416 (O_416,N_19611,N_19702);
or UO_417 (O_417,N_19608,N_19848);
and UO_418 (O_418,N_19909,N_19809);
nand UO_419 (O_419,N_19661,N_19778);
and UO_420 (O_420,N_19845,N_19677);
nor UO_421 (O_421,N_19690,N_19650);
or UO_422 (O_422,N_19809,N_19609);
and UO_423 (O_423,N_19869,N_19937);
or UO_424 (O_424,N_19626,N_19923);
or UO_425 (O_425,N_19834,N_19750);
nand UO_426 (O_426,N_19735,N_19613);
or UO_427 (O_427,N_19853,N_19653);
or UO_428 (O_428,N_19761,N_19838);
and UO_429 (O_429,N_19969,N_19617);
nand UO_430 (O_430,N_19822,N_19743);
xor UO_431 (O_431,N_19680,N_19834);
xnor UO_432 (O_432,N_19885,N_19945);
or UO_433 (O_433,N_19776,N_19708);
nor UO_434 (O_434,N_19819,N_19946);
nor UO_435 (O_435,N_19877,N_19967);
xor UO_436 (O_436,N_19973,N_19806);
nand UO_437 (O_437,N_19630,N_19711);
or UO_438 (O_438,N_19812,N_19910);
or UO_439 (O_439,N_19876,N_19624);
xor UO_440 (O_440,N_19707,N_19772);
and UO_441 (O_441,N_19699,N_19858);
or UO_442 (O_442,N_19732,N_19949);
nor UO_443 (O_443,N_19885,N_19967);
nor UO_444 (O_444,N_19797,N_19766);
nand UO_445 (O_445,N_19835,N_19704);
xor UO_446 (O_446,N_19934,N_19957);
nor UO_447 (O_447,N_19738,N_19962);
or UO_448 (O_448,N_19647,N_19999);
nand UO_449 (O_449,N_19819,N_19990);
or UO_450 (O_450,N_19873,N_19695);
and UO_451 (O_451,N_19600,N_19842);
xnor UO_452 (O_452,N_19867,N_19714);
or UO_453 (O_453,N_19658,N_19695);
nand UO_454 (O_454,N_19750,N_19773);
xor UO_455 (O_455,N_19736,N_19697);
nor UO_456 (O_456,N_19828,N_19958);
or UO_457 (O_457,N_19777,N_19839);
xor UO_458 (O_458,N_19959,N_19716);
and UO_459 (O_459,N_19706,N_19988);
or UO_460 (O_460,N_19882,N_19719);
or UO_461 (O_461,N_19605,N_19610);
and UO_462 (O_462,N_19603,N_19831);
xnor UO_463 (O_463,N_19867,N_19709);
nand UO_464 (O_464,N_19675,N_19836);
nor UO_465 (O_465,N_19690,N_19828);
nor UO_466 (O_466,N_19862,N_19895);
nand UO_467 (O_467,N_19738,N_19870);
or UO_468 (O_468,N_19933,N_19733);
and UO_469 (O_469,N_19965,N_19922);
xnor UO_470 (O_470,N_19820,N_19610);
or UO_471 (O_471,N_19824,N_19931);
nor UO_472 (O_472,N_19647,N_19730);
xor UO_473 (O_473,N_19735,N_19894);
or UO_474 (O_474,N_19847,N_19961);
and UO_475 (O_475,N_19761,N_19731);
or UO_476 (O_476,N_19781,N_19640);
and UO_477 (O_477,N_19719,N_19869);
nor UO_478 (O_478,N_19899,N_19801);
and UO_479 (O_479,N_19763,N_19900);
and UO_480 (O_480,N_19831,N_19608);
or UO_481 (O_481,N_19896,N_19709);
and UO_482 (O_482,N_19755,N_19705);
or UO_483 (O_483,N_19697,N_19975);
nor UO_484 (O_484,N_19855,N_19812);
nor UO_485 (O_485,N_19811,N_19972);
nor UO_486 (O_486,N_19670,N_19961);
nand UO_487 (O_487,N_19943,N_19741);
nor UO_488 (O_488,N_19720,N_19866);
nor UO_489 (O_489,N_19823,N_19930);
xor UO_490 (O_490,N_19765,N_19968);
nor UO_491 (O_491,N_19741,N_19918);
xnor UO_492 (O_492,N_19865,N_19848);
xor UO_493 (O_493,N_19978,N_19636);
xnor UO_494 (O_494,N_19702,N_19671);
nor UO_495 (O_495,N_19733,N_19807);
nor UO_496 (O_496,N_19753,N_19811);
and UO_497 (O_497,N_19993,N_19755);
and UO_498 (O_498,N_19751,N_19811);
nand UO_499 (O_499,N_19747,N_19643);
and UO_500 (O_500,N_19914,N_19955);
and UO_501 (O_501,N_19780,N_19864);
xor UO_502 (O_502,N_19920,N_19610);
or UO_503 (O_503,N_19893,N_19791);
or UO_504 (O_504,N_19669,N_19877);
nor UO_505 (O_505,N_19607,N_19611);
or UO_506 (O_506,N_19626,N_19685);
nand UO_507 (O_507,N_19684,N_19880);
xor UO_508 (O_508,N_19729,N_19805);
and UO_509 (O_509,N_19918,N_19692);
xor UO_510 (O_510,N_19861,N_19988);
or UO_511 (O_511,N_19625,N_19977);
and UO_512 (O_512,N_19814,N_19627);
nor UO_513 (O_513,N_19847,N_19907);
nor UO_514 (O_514,N_19921,N_19970);
or UO_515 (O_515,N_19953,N_19829);
or UO_516 (O_516,N_19639,N_19866);
or UO_517 (O_517,N_19661,N_19909);
and UO_518 (O_518,N_19730,N_19668);
xor UO_519 (O_519,N_19958,N_19834);
xor UO_520 (O_520,N_19900,N_19620);
nand UO_521 (O_521,N_19682,N_19614);
nor UO_522 (O_522,N_19736,N_19758);
or UO_523 (O_523,N_19941,N_19908);
nand UO_524 (O_524,N_19850,N_19661);
and UO_525 (O_525,N_19652,N_19873);
nor UO_526 (O_526,N_19908,N_19982);
nand UO_527 (O_527,N_19705,N_19771);
nor UO_528 (O_528,N_19881,N_19823);
xnor UO_529 (O_529,N_19744,N_19988);
nor UO_530 (O_530,N_19634,N_19637);
or UO_531 (O_531,N_19760,N_19990);
nand UO_532 (O_532,N_19871,N_19632);
nor UO_533 (O_533,N_19885,N_19821);
nor UO_534 (O_534,N_19718,N_19844);
nand UO_535 (O_535,N_19973,N_19862);
xnor UO_536 (O_536,N_19849,N_19998);
and UO_537 (O_537,N_19871,N_19729);
nor UO_538 (O_538,N_19731,N_19748);
xnor UO_539 (O_539,N_19937,N_19986);
nand UO_540 (O_540,N_19842,N_19963);
xnor UO_541 (O_541,N_19656,N_19688);
or UO_542 (O_542,N_19800,N_19882);
and UO_543 (O_543,N_19881,N_19736);
and UO_544 (O_544,N_19969,N_19747);
nor UO_545 (O_545,N_19832,N_19664);
xor UO_546 (O_546,N_19744,N_19751);
nor UO_547 (O_547,N_19610,N_19648);
and UO_548 (O_548,N_19881,N_19926);
nand UO_549 (O_549,N_19736,N_19903);
nand UO_550 (O_550,N_19629,N_19744);
and UO_551 (O_551,N_19758,N_19750);
nand UO_552 (O_552,N_19838,N_19950);
or UO_553 (O_553,N_19711,N_19661);
xor UO_554 (O_554,N_19615,N_19796);
xor UO_555 (O_555,N_19817,N_19706);
nor UO_556 (O_556,N_19769,N_19945);
xnor UO_557 (O_557,N_19721,N_19753);
and UO_558 (O_558,N_19968,N_19698);
nand UO_559 (O_559,N_19793,N_19766);
nor UO_560 (O_560,N_19904,N_19885);
and UO_561 (O_561,N_19607,N_19938);
or UO_562 (O_562,N_19628,N_19717);
xor UO_563 (O_563,N_19603,N_19820);
and UO_564 (O_564,N_19942,N_19925);
nor UO_565 (O_565,N_19717,N_19693);
nand UO_566 (O_566,N_19949,N_19776);
nand UO_567 (O_567,N_19763,N_19627);
and UO_568 (O_568,N_19868,N_19942);
nor UO_569 (O_569,N_19767,N_19736);
and UO_570 (O_570,N_19673,N_19923);
and UO_571 (O_571,N_19791,N_19892);
nor UO_572 (O_572,N_19795,N_19864);
or UO_573 (O_573,N_19854,N_19646);
or UO_574 (O_574,N_19946,N_19846);
nand UO_575 (O_575,N_19928,N_19865);
xor UO_576 (O_576,N_19866,N_19617);
xnor UO_577 (O_577,N_19889,N_19795);
xor UO_578 (O_578,N_19652,N_19947);
nand UO_579 (O_579,N_19983,N_19646);
and UO_580 (O_580,N_19730,N_19728);
nor UO_581 (O_581,N_19835,N_19777);
xor UO_582 (O_582,N_19970,N_19924);
nor UO_583 (O_583,N_19845,N_19888);
and UO_584 (O_584,N_19758,N_19610);
nor UO_585 (O_585,N_19984,N_19911);
or UO_586 (O_586,N_19671,N_19674);
nand UO_587 (O_587,N_19664,N_19776);
or UO_588 (O_588,N_19692,N_19936);
nand UO_589 (O_589,N_19638,N_19949);
and UO_590 (O_590,N_19797,N_19688);
and UO_591 (O_591,N_19693,N_19709);
and UO_592 (O_592,N_19808,N_19833);
or UO_593 (O_593,N_19849,N_19994);
xor UO_594 (O_594,N_19686,N_19684);
and UO_595 (O_595,N_19989,N_19791);
xnor UO_596 (O_596,N_19834,N_19662);
or UO_597 (O_597,N_19877,N_19621);
or UO_598 (O_598,N_19681,N_19671);
and UO_599 (O_599,N_19709,N_19859);
xor UO_600 (O_600,N_19677,N_19756);
nand UO_601 (O_601,N_19960,N_19633);
xnor UO_602 (O_602,N_19686,N_19636);
and UO_603 (O_603,N_19930,N_19640);
nor UO_604 (O_604,N_19602,N_19910);
nor UO_605 (O_605,N_19706,N_19718);
nor UO_606 (O_606,N_19619,N_19601);
or UO_607 (O_607,N_19691,N_19885);
nor UO_608 (O_608,N_19695,N_19772);
and UO_609 (O_609,N_19791,N_19816);
or UO_610 (O_610,N_19898,N_19919);
nor UO_611 (O_611,N_19930,N_19744);
nor UO_612 (O_612,N_19690,N_19820);
and UO_613 (O_613,N_19664,N_19938);
and UO_614 (O_614,N_19601,N_19658);
nor UO_615 (O_615,N_19897,N_19890);
xnor UO_616 (O_616,N_19724,N_19666);
xor UO_617 (O_617,N_19738,N_19846);
xor UO_618 (O_618,N_19796,N_19601);
or UO_619 (O_619,N_19633,N_19839);
and UO_620 (O_620,N_19899,N_19852);
nand UO_621 (O_621,N_19957,N_19788);
xor UO_622 (O_622,N_19807,N_19879);
or UO_623 (O_623,N_19948,N_19982);
xnor UO_624 (O_624,N_19846,N_19807);
nor UO_625 (O_625,N_19923,N_19674);
nor UO_626 (O_626,N_19727,N_19696);
and UO_627 (O_627,N_19926,N_19880);
or UO_628 (O_628,N_19905,N_19950);
nand UO_629 (O_629,N_19613,N_19909);
nand UO_630 (O_630,N_19972,N_19996);
and UO_631 (O_631,N_19680,N_19602);
nand UO_632 (O_632,N_19637,N_19758);
or UO_633 (O_633,N_19988,N_19611);
or UO_634 (O_634,N_19636,N_19941);
nor UO_635 (O_635,N_19635,N_19882);
and UO_636 (O_636,N_19942,N_19812);
xor UO_637 (O_637,N_19668,N_19669);
nor UO_638 (O_638,N_19832,N_19730);
or UO_639 (O_639,N_19921,N_19662);
and UO_640 (O_640,N_19693,N_19886);
and UO_641 (O_641,N_19801,N_19813);
and UO_642 (O_642,N_19738,N_19729);
or UO_643 (O_643,N_19658,N_19622);
xnor UO_644 (O_644,N_19676,N_19983);
and UO_645 (O_645,N_19901,N_19794);
nand UO_646 (O_646,N_19903,N_19621);
nor UO_647 (O_647,N_19771,N_19864);
nand UO_648 (O_648,N_19703,N_19749);
nor UO_649 (O_649,N_19957,N_19633);
or UO_650 (O_650,N_19797,N_19721);
and UO_651 (O_651,N_19902,N_19869);
xor UO_652 (O_652,N_19862,N_19971);
nor UO_653 (O_653,N_19825,N_19603);
or UO_654 (O_654,N_19615,N_19882);
or UO_655 (O_655,N_19608,N_19611);
and UO_656 (O_656,N_19944,N_19722);
or UO_657 (O_657,N_19999,N_19945);
nor UO_658 (O_658,N_19927,N_19824);
or UO_659 (O_659,N_19615,N_19789);
nand UO_660 (O_660,N_19981,N_19751);
nand UO_661 (O_661,N_19919,N_19794);
xor UO_662 (O_662,N_19857,N_19890);
nor UO_663 (O_663,N_19672,N_19794);
and UO_664 (O_664,N_19850,N_19705);
and UO_665 (O_665,N_19817,N_19886);
nor UO_666 (O_666,N_19714,N_19878);
nor UO_667 (O_667,N_19709,N_19606);
and UO_668 (O_668,N_19781,N_19620);
nor UO_669 (O_669,N_19781,N_19786);
nand UO_670 (O_670,N_19689,N_19640);
or UO_671 (O_671,N_19707,N_19778);
and UO_672 (O_672,N_19874,N_19854);
xor UO_673 (O_673,N_19693,N_19726);
and UO_674 (O_674,N_19676,N_19810);
xor UO_675 (O_675,N_19858,N_19978);
xnor UO_676 (O_676,N_19826,N_19764);
xor UO_677 (O_677,N_19720,N_19730);
nand UO_678 (O_678,N_19721,N_19670);
nand UO_679 (O_679,N_19639,N_19908);
xnor UO_680 (O_680,N_19823,N_19922);
nor UO_681 (O_681,N_19695,N_19981);
or UO_682 (O_682,N_19616,N_19626);
xor UO_683 (O_683,N_19727,N_19630);
nor UO_684 (O_684,N_19639,N_19628);
xor UO_685 (O_685,N_19631,N_19918);
nor UO_686 (O_686,N_19774,N_19684);
xnor UO_687 (O_687,N_19783,N_19714);
xor UO_688 (O_688,N_19639,N_19874);
xnor UO_689 (O_689,N_19904,N_19936);
nor UO_690 (O_690,N_19660,N_19778);
xnor UO_691 (O_691,N_19724,N_19670);
or UO_692 (O_692,N_19854,N_19612);
nor UO_693 (O_693,N_19988,N_19705);
nand UO_694 (O_694,N_19886,N_19779);
nor UO_695 (O_695,N_19714,N_19686);
nand UO_696 (O_696,N_19999,N_19754);
or UO_697 (O_697,N_19754,N_19873);
xnor UO_698 (O_698,N_19955,N_19848);
nor UO_699 (O_699,N_19659,N_19814);
xor UO_700 (O_700,N_19720,N_19983);
nand UO_701 (O_701,N_19623,N_19670);
xor UO_702 (O_702,N_19688,N_19849);
nor UO_703 (O_703,N_19693,N_19600);
and UO_704 (O_704,N_19704,N_19983);
or UO_705 (O_705,N_19983,N_19629);
nand UO_706 (O_706,N_19676,N_19817);
nand UO_707 (O_707,N_19677,N_19680);
or UO_708 (O_708,N_19999,N_19937);
nor UO_709 (O_709,N_19678,N_19994);
xor UO_710 (O_710,N_19721,N_19864);
nand UO_711 (O_711,N_19641,N_19608);
and UO_712 (O_712,N_19794,N_19671);
or UO_713 (O_713,N_19680,N_19919);
and UO_714 (O_714,N_19734,N_19906);
nor UO_715 (O_715,N_19642,N_19730);
nor UO_716 (O_716,N_19741,N_19671);
and UO_717 (O_717,N_19875,N_19822);
xor UO_718 (O_718,N_19840,N_19798);
nor UO_719 (O_719,N_19800,N_19801);
or UO_720 (O_720,N_19713,N_19791);
nand UO_721 (O_721,N_19795,N_19886);
nand UO_722 (O_722,N_19798,N_19977);
xnor UO_723 (O_723,N_19955,N_19699);
nand UO_724 (O_724,N_19855,N_19992);
nor UO_725 (O_725,N_19749,N_19636);
or UO_726 (O_726,N_19657,N_19624);
or UO_727 (O_727,N_19608,N_19673);
and UO_728 (O_728,N_19642,N_19904);
xnor UO_729 (O_729,N_19835,N_19749);
and UO_730 (O_730,N_19783,N_19631);
nand UO_731 (O_731,N_19986,N_19762);
nand UO_732 (O_732,N_19635,N_19861);
nand UO_733 (O_733,N_19646,N_19961);
xor UO_734 (O_734,N_19765,N_19992);
and UO_735 (O_735,N_19775,N_19757);
or UO_736 (O_736,N_19699,N_19841);
and UO_737 (O_737,N_19645,N_19641);
xnor UO_738 (O_738,N_19623,N_19651);
nor UO_739 (O_739,N_19924,N_19963);
xor UO_740 (O_740,N_19675,N_19699);
nand UO_741 (O_741,N_19778,N_19808);
and UO_742 (O_742,N_19762,N_19781);
xor UO_743 (O_743,N_19776,N_19976);
nand UO_744 (O_744,N_19680,N_19937);
nand UO_745 (O_745,N_19983,N_19829);
nand UO_746 (O_746,N_19810,N_19993);
nor UO_747 (O_747,N_19642,N_19923);
nand UO_748 (O_748,N_19916,N_19964);
or UO_749 (O_749,N_19650,N_19997);
nor UO_750 (O_750,N_19756,N_19874);
xnor UO_751 (O_751,N_19960,N_19733);
or UO_752 (O_752,N_19694,N_19642);
xnor UO_753 (O_753,N_19860,N_19606);
and UO_754 (O_754,N_19826,N_19607);
and UO_755 (O_755,N_19702,N_19784);
xor UO_756 (O_756,N_19694,N_19817);
xnor UO_757 (O_757,N_19658,N_19884);
nand UO_758 (O_758,N_19710,N_19877);
nor UO_759 (O_759,N_19784,N_19602);
xnor UO_760 (O_760,N_19863,N_19906);
and UO_761 (O_761,N_19989,N_19993);
nand UO_762 (O_762,N_19751,N_19722);
nor UO_763 (O_763,N_19750,N_19844);
nor UO_764 (O_764,N_19937,N_19936);
and UO_765 (O_765,N_19728,N_19792);
and UO_766 (O_766,N_19613,N_19713);
xnor UO_767 (O_767,N_19702,N_19805);
or UO_768 (O_768,N_19980,N_19746);
xnor UO_769 (O_769,N_19914,N_19779);
nand UO_770 (O_770,N_19726,N_19999);
or UO_771 (O_771,N_19671,N_19952);
or UO_772 (O_772,N_19870,N_19914);
xor UO_773 (O_773,N_19707,N_19982);
or UO_774 (O_774,N_19980,N_19749);
nand UO_775 (O_775,N_19902,N_19945);
xnor UO_776 (O_776,N_19962,N_19843);
and UO_777 (O_777,N_19602,N_19859);
nand UO_778 (O_778,N_19649,N_19765);
nor UO_779 (O_779,N_19657,N_19639);
or UO_780 (O_780,N_19908,N_19891);
or UO_781 (O_781,N_19664,N_19614);
and UO_782 (O_782,N_19695,N_19610);
or UO_783 (O_783,N_19622,N_19889);
nor UO_784 (O_784,N_19617,N_19791);
and UO_785 (O_785,N_19895,N_19890);
nand UO_786 (O_786,N_19664,N_19779);
nand UO_787 (O_787,N_19688,N_19816);
or UO_788 (O_788,N_19995,N_19949);
or UO_789 (O_789,N_19970,N_19936);
xnor UO_790 (O_790,N_19996,N_19700);
or UO_791 (O_791,N_19854,N_19729);
nor UO_792 (O_792,N_19986,N_19825);
or UO_793 (O_793,N_19784,N_19662);
or UO_794 (O_794,N_19892,N_19915);
or UO_795 (O_795,N_19782,N_19797);
or UO_796 (O_796,N_19618,N_19885);
and UO_797 (O_797,N_19993,N_19964);
xnor UO_798 (O_798,N_19938,N_19916);
or UO_799 (O_799,N_19873,N_19897);
and UO_800 (O_800,N_19987,N_19905);
or UO_801 (O_801,N_19931,N_19932);
or UO_802 (O_802,N_19827,N_19752);
xnor UO_803 (O_803,N_19643,N_19737);
nand UO_804 (O_804,N_19687,N_19815);
nor UO_805 (O_805,N_19734,N_19907);
or UO_806 (O_806,N_19906,N_19691);
nor UO_807 (O_807,N_19813,N_19803);
or UO_808 (O_808,N_19620,N_19619);
and UO_809 (O_809,N_19981,N_19881);
or UO_810 (O_810,N_19833,N_19741);
nor UO_811 (O_811,N_19933,N_19622);
nor UO_812 (O_812,N_19667,N_19754);
xor UO_813 (O_813,N_19992,N_19633);
nand UO_814 (O_814,N_19916,N_19666);
xor UO_815 (O_815,N_19858,N_19949);
or UO_816 (O_816,N_19871,N_19805);
or UO_817 (O_817,N_19701,N_19936);
xnor UO_818 (O_818,N_19700,N_19938);
nor UO_819 (O_819,N_19758,N_19993);
nor UO_820 (O_820,N_19761,N_19682);
or UO_821 (O_821,N_19694,N_19974);
nor UO_822 (O_822,N_19814,N_19783);
nand UO_823 (O_823,N_19975,N_19705);
nor UO_824 (O_824,N_19746,N_19705);
nor UO_825 (O_825,N_19848,N_19614);
and UO_826 (O_826,N_19898,N_19949);
nand UO_827 (O_827,N_19864,N_19692);
and UO_828 (O_828,N_19886,N_19618);
xor UO_829 (O_829,N_19962,N_19756);
xor UO_830 (O_830,N_19743,N_19738);
xnor UO_831 (O_831,N_19848,N_19824);
and UO_832 (O_832,N_19740,N_19765);
and UO_833 (O_833,N_19853,N_19993);
nand UO_834 (O_834,N_19991,N_19672);
nor UO_835 (O_835,N_19760,N_19660);
and UO_836 (O_836,N_19707,N_19716);
nand UO_837 (O_837,N_19856,N_19936);
nor UO_838 (O_838,N_19957,N_19742);
or UO_839 (O_839,N_19933,N_19949);
or UO_840 (O_840,N_19848,N_19985);
or UO_841 (O_841,N_19806,N_19605);
or UO_842 (O_842,N_19698,N_19753);
nand UO_843 (O_843,N_19630,N_19979);
or UO_844 (O_844,N_19628,N_19630);
and UO_845 (O_845,N_19737,N_19878);
nand UO_846 (O_846,N_19659,N_19923);
nor UO_847 (O_847,N_19672,N_19852);
or UO_848 (O_848,N_19824,N_19995);
xor UO_849 (O_849,N_19893,N_19616);
nor UO_850 (O_850,N_19776,N_19851);
nand UO_851 (O_851,N_19908,N_19707);
nand UO_852 (O_852,N_19904,N_19772);
nand UO_853 (O_853,N_19679,N_19684);
nor UO_854 (O_854,N_19839,N_19744);
nand UO_855 (O_855,N_19968,N_19879);
and UO_856 (O_856,N_19935,N_19842);
or UO_857 (O_857,N_19805,N_19984);
xnor UO_858 (O_858,N_19612,N_19924);
or UO_859 (O_859,N_19759,N_19710);
nor UO_860 (O_860,N_19951,N_19685);
nand UO_861 (O_861,N_19681,N_19757);
and UO_862 (O_862,N_19774,N_19931);
or UO_863 (O_863,N_19986,N_19746);
and UO_864 (O_864,N_19712,N_19998);
xnor UO_865 (O_865,N_19917,N_19766);
or UO_866 (O_866,N_19845,N_19711);
xnor UO_867 (O_867,N_19832,N_19928);
xor UO_868 (O_868,N_19820,N_19972);
nand UO_869 (O_869,N_19891,N_19662);
nand UO_870 (O_870,N_19901,N_19672);
and UO_871 (O_871,N_19841,N_19948);
xor UO_872 (O_872,N_19883,N_19841);
and UO_873 (O_873,N_19694,N_19708);
nor UO_874 (O_874,N_19809,N_19696);
xnor UO_875 (O_875,N_19862,N_19923);
nor UO_876 (O_876,N_19783,N_19823);
or UO_877 (O_877,N_19900,N_19808);
nor UO_878 (O_878,N_19642,N_19842);
nand UO_879 (O_879,N_19611,N_19890);
nor UO_880 (O_880,N_19763,N_19979);
and UO_881 (O_881,N_19720,N_19764);
xnor UO_882 (O_882,N_19938,N_19885);
xor UO_883 (O_883,N_19656,N_19635);
and UO_884 (O_884,N_19888,N_19914);
nand UO_885 (O_885,N_19921,N_19815);
nor UO_886 (O_886,N_19627,N_19749);
and UO_887 (O_887,N_19946,N_19632);
and UO_888 (O_888,N_19793,N_19808);
xnor UO_889 (O_889,N_19888,N_19784);
nor UO_890 (O_890,N_19707,N_19984);
or UO_891 (O_891,N_19833,N_19906);
nand UO_892 (O_892,N_19773,N_19689);
and UO_893 (O_893,N_19991,N_19890);
and UO_894 (O_894,N_19752,N_19873);
xnor UO_895 (O_895,N_19672,N_19953);
nand UO_896 (O_896,N_19973,N_19887);
and UO_897 (O_897,N_19681,N_19737);
and UO_898 (O_898,N_19949,N_19681);
nand UO_899 (O_899,N_19618,N_19904);
xnor UO_900 (O_900,N_19946,N_19612);
and UO_901 (O_901,N_19635,N_19740);
nor UO_902 (O_902,N_19912,N_19994);
or UO_903 (O_903,N_19628,N_19769);
nand UO_904 (O_904,N_19738,N_19640);
and UO_905 (O_905,N_19895,N_19659);
and UO_906 (O_906,N_19701,N_19707);
nand UO_907 (O_907,N_19829,N_19952);
xor UO_908 (O_908,N_19901,N_19991);
nor UO_909 (O_909,N_19771,N_19795);
and UO_910 (O_910,N_19651,N_19994);
and UO_911 (O_911,N_19700,N_19613);
nand UO_912 (O_912,N_19706,N_19962);
nand UO_913 (O_913,N_19931,N_19989);
or UO_914 (O_914,N_19996,N_19726);
xor UO_915 (O_915,N_19762,N_19675);
and UO_916 (O_916,N_19620,N_19726);
and UO_917 (O_917,N_19612,N_19801);
nor UO_918 (O_918,N_19789,N_19768);
nor UO_919 (O_919,N_19656,N_19720);
or UO_920 (O_920,N_19977,N_19776);
and UO_921 (O_921,N_19977,N_19657);
xnor UO_922 (O_922,N_19820,N_19852);
and UO_923 (O_923,N_19612,N_19619);
nand UO_924 (O_924,N_19825,N_19981);
nand UO_925 (O_925,N_19920,N_19824);
or UO_926 (O_926,N_19705,N_19699);
or UO_927 (O_927,N_19612,N_19935);
nor UO_928 (O_928,N_19633,N_19935);
nor UO_929 (O_929,N_19659,N_19906);
xnor UO_930 (O_930,N_19885,N_19873);
nand UO_931 (O_931,N_19831,N_19933);
or UO_932 (O_932,N_19814,N_19898);
nand UO_933 (O_933,N_19917,N_19931);
and UO_934 (O_934,N_19888,N_19819);
nand UO_935 (O_935,N_19761,N_19680);
xor UO_936 (O_936,N_19920,N_19626);
nand UO_937 (O_937,N_19929,N_19668);
xor UO_938 (O_938,N_19718,N_19662);
and UO_939 (O_939,N_19912,N_19976);
nor UO_940 (O_940,N_19844,N_19663);
and UO_941 (O_941,N_19791,N_19722);
xnor UO_942 (O_942,N_19855,N_19933);
or UO_943 (O_943,N_19934,N_19602);
or UO_944 (O_944,N_19781,N_19631);
nand UO_945 (O_945,N_19608,N_19619);
nand UO_946 (O_946,N_19695,N_19713);
and UO_947 (O_947,N_19748,N_19781);
xnor UO_948 (O_948,N_19950,N_19831);
and UO_949 (O_949,N_19677,N_19947);
nor UO_950 (O_950,N_19900,N_19758);
xnor UO_951 (O_951,N_19810,N_19756);
nor UO_952 (O_952,N_19918,N_19676);
nor UO_953 (O_953,N_19857,N_19620);
nor UO_954 (O_954,N_19917,N_19791);
or UO_955 (O_955,N_19681,N_19657);
and UO_956 (O_956,N_19752,N_19674);
xnor UO_957 (O_957,N_19700,N_19828);
nand UO_958 (O_958,N_19734,N_19744);
nor UO_959 (O_959,N_19872,N_19983);
xor UO_960 (O_960,N_19850,N_19840);
nand UO_961 (O_961,N_19700,N_19739);
and UO_962 (O_962,N_19874,N_19956);
nand UO_963 (O_963,N_19858,N_19930);
nand UO_964 (O_964,N_19837,N_19675);
or UO_965 (O_965,N_19810,N_19671);
or UO_966 (O_966,N_19710,N_19868);
nor UO_967 (O_967,N_19725,N_19811);
or UO_968 (O_968,N_19907,N_19934);
nor UO_969 (O_969,N_19861,N_19815);
nor UO_970 (O_970,N_19860,N_19805);
and UO_971 (O_971,N_19836,N_19884);
or UO_972 (O_972,N_19681,N_19936);
and UO_973 (O_973,N_19699,N_19603);
xor UO_974 (O_974,N_19675,N_19602);
nor UO_975 (O_975,N_19695,N_19653);
or UO_976 (O_976,N_19811,N_19796);
or UO_977 (O_977,N_19721,N_19724);
xor UO_978 (O_978,N_19621,N_19640);
and UO_979 (O_979,N_19800,N_19959);
nor UO_980 (O_980,N_19613,N_19778);
xnor UO_981 (O_981,N_19950,N_19674);
xor UO_982 (O_982,N_19621,N_19852);
nand UO_983 (O_983,N_19784,N_19940);
xor UO_984 (O_984,N_19850,N_19799);
or UO_985 (O_985,N_19830,N_19742);
and UO_986 (O_986,N_19809,N_19637);
and UO_987 (O_987,N_19936,N_19857);
or UO_988 (O_988,N_19934,N_19784);
and UO_989 (O_989,N_19865,N_19670);
nand UO_990 (O_990,N_19613,N_19628);
and UO_991 (O_991,N_19749,N_19718);
nor UO_992 (O_992,N_19938,N_19744);
or UO_993 (O_993,N_19809,N_19811);
or UO_994 (O_994,N_19849,N_19647);
xnor UO_995 (O_995,N_19733,N_19724);
or UO_996 (O_996,N_19689,N_19858);
nand UO_997 (O_997,N_19880,N_19654);
or UO_998 (O_998,N_19766,N_19843);
nor UO_999 (O_999,N_19671,N_19802);
nor UO_1000 (O_1000,N_19630,N_19710);
xnor UO_1001 (O_1001,N_19609,N_19741);
nor UO_1002 (O_1002,N_19903,N_19656);
nand UO_1003 (O_1003,N_19735,N_19925);
nand UO_1004 (O_1004,N_19630,N_19901);
xnor UO_1005 (O_1005,N_19674,N_19811);
nand UO_1006 (O_1006,N_19631,N_19954);
and UO_1007 (O_1007,N_19989,N_19788);
xor UO_1008 (O_1008,N_19939,N_19806);
nor UO_1009 (O_1009,N_19843,N_19907);
and UO_1010 (O_1010,N_19757,N_19759);
xor UO_1011 (O_1011,N_19660,N_19849);
and UO_1012 (O_1012,N_19923,N_19798);
and UO_1013 (O_1013,N_19863,N_19787);
nor UO_1014 (O_1014,N_19860,N_19653);
and UO_1015 (O_1015,N_19962,N_19758);
xnor UO_1016 (O_1016,N_19841,N_19806);
nor UO_1017 (O_1017,N_19834,N_19852);
or UO_1018 (O_1018,N_19637,N_19731);
nor UO_1019 (O_1019,N_19790,N_19745);
nand UO_1020 (O_1020,N_19732,N_19824);
and UO_1021 (O_1021,N_19918,N_19677);
nor UO_1022 (O_1022,N_19681,N_19877);
nand UO_1023 (O_1023,N_19681,N_19926);
and UO_1024 (O_1024,N_19650,N_19781);
and UO_1025 (O_1025,N_19845,N_19822);
xnor UO_1026 (O_1026,N_19847,N_19671);
and UO_1027 (O_1027,N_19879,N_19837);
or UO_1028 (O_1028,N_19748,N_19930);
nor UO_1029 (O_1029,N_19923,N_19729);
and UO_1030 (O_1030,N_19826,N_19970);
and UO_1031 (O_1031,N_19752,N_19879);
nand UO_1032 (O_1032,N_19700,N_19979);
xnor UO_1033 (O_1033,N_19696,N_19762);
or UO_1034 (O_1034,N_19990,N_19724);
or UO_1035 (O_1035,N_19784,N_19996);
or UO_1036 (O_1036,N_19602,N_19712);
xnor UO_1037 (O_1037,N_19677,N_19600);
and UO_1038 (O_1038,N_19869,N_19684);
nand UO_1039 (O_1039,N_19872,N_19839);
nor UO_1040 (O_1040,N_19672,N_19939);
and UO_1041 (O_1041,N_19977,N_19806);
and UO_1042 (O_1042,N_19842,N_19882);
nor UO_1043 (O_1043,N_19893,N_19921);
nand UO_1044 (O_1044,N_19921,N_19829);
and UO_1045 (O_1045,N_19955,N_19779);
or UO_1046 (O_1046,N_19866,N_19897);
and UO_1047 (O_1047,N_19855,N_19737);
xnor UO_1048 (O_1048,N_19819,N_19918);
nand UO_1049 (O_1049,N_19722,N_19941);
and UO_1050 (O_1050,N_19926,N_19904);
nand UO_1051 (O_1051,N_19971,N_19682);
nand UO_1052 (O_1052,N_19705,N_19831);
xnor UO_1053 (O_1053,N_19608,N_19746);
nor UO_1054 (O_1054,N_19747,N_19884);
and UO_1055 (O_1055,N_19650,N_19780);
xor UO_1056 (O_1056,N_19833,N_19609);
nand UO_1057 (O_1057,N_19715,N_19997);
and UO_1058 (O_1058,N_19959,N_19710);
xnor UO_1059 (O_1059,N_19660,N_19911);
or UO_1060 (O_1060,N_19920,N_19783);
nand UO_1061 (O_1061,N_19901,N_19629);
nor UO_1062 (O_1062,N_19735,N_19921);
and UO_1063 (O_1063,N_19728,N_19891);
or UO_1064 (O_1064,N_19866,N_19894);
or UO_1065 (O_1065,N_19648,N_19784);
xor UO_1066 (O_1066,N_19610,N_19959);
nand UO_1067 (O_1067,N_19958,N_19989);
or UO_1068 (O_1068,N_19821,N_19977);
nand UO_1069 (O_1069,N_19806,N_19922);
and UO_1070 (O_1070,N_19839,N_19791);
nor UO_1071 (O_1071,N_19970,N_19762);
nand UO_1072 (O_1072,N_19908,N_19638);
nand UO_1073 (O_1073,N_19836,N_19713);
or UO_1074 (O_1074,N_19704,N_19979);
or UO_1075 (O_1075,N_19695,N_19639);
xnor UO_1076 (O_1076,N_19697,N_19894);
nand UO_1077 (O_1077,N_19880,N_19922);
and UO_1078 (O_1078,N_19924,N_19642);
or UO_1079 (O_1079,N_19989,N_19794);
and UO_1080 (O_1080,N_19952,N_19981);
xor UO_1081 (O_1081,N_19640,N_19854);
xor UO_1082 (O_1082,N_19790,N_19997);
and UO_1083 (O_1083,N_19984,N_19627);
nand UO_1084 (O_1084,N_19763,N_19951);
xnor UO_1085 (O_1085,N_19761,N_19709);
and UO_1086 (O_1086,N_19730,N_19854);
nor UO_1087 (O_1087,N_19632,N_19852);
or UO_1088 (O_1088,N_19994,N_19711);
or UO_1089 (O_1089,N_19932,N_19638);
or UO_1090 (O_1090,N_19992,N_19872);
nor UO_1091 (O_1091,N_19871,N_19980);
nor UO_1092 (O_1092,N_19726,N_19841);
and UO_1093 (O_1093,N_19945,N_19762);
or UO_1094 (O_1094,N_19948,N_19666);
nand UO_1095 (O_1095,N_19804,N_19909);
or UO_1096 (O_1096,N_19910,N_19756);
or UO_1097 (O_1097,N_19714,N_19977);
xor UO_1098 (O_1098,N_19615,N_19949);
nor UO_1099 (O_1099,N_19654,N_19988);
nand UO_1100 (O_1100,N_19997,N_19857);
nand UO_1101 (O_1101,N_19706,N_19801);
and UO_1102 (O_1102,N_19829,N_19737);
and UO_1103 (O_1103,N_19672,N_19867);
and UO_1104 (O_1104,N_19667,N_19917);
xor UO_1105 (O_1105,N_19767,N_19635);
or UO_1106 (O_1106,N_19741,N_19801);
or UO_1107 (O_1107,N_19915,N_19661);
xnor UO_1108 (O_1108,N_19632,N_19851);
or UO_1109 (O_1109,N_19620,N_19814);
and UO_1110 (O_1110,N_19793,N_19607);
nand UO_1111 (O_1111,N_19685,N_19895);
and UO_1112 (O_1112,N_19873,N_19911);
xnor UO_1113 (O_1113,N_19689,N_19821);
nor UO_1114 (O_1114,N_19669,N_19634);
and UO_1115 (O_1115,N_19973,N_19765);
nand UO_1116 (O_1116,N_19915,N_19660);
nor UO_1117 (O_1117,N_19637,N_19721);
nand UO_1118 (O_1118,N_19727,N_19995);
nor UO_1119 (O_1119,N_19736,N_19783);
xnor UO_1120 (O_1120,N_19999,N_19963);
or UO_1121 (O_1121,N_19786,N_19958);
nand UO_1122 (O_1122,N_19775,N_19660);
nand UO_1123 (O_1123,N_19611,N_19910);
xnor UO_1124 (O_1124,N_19860,N_19762);
and UO_1125 (O_1125,N_19903,N_19677);
or UO_1126 (O_1126,N_19741,N_19798);
nand UO_1127 (O_1127,N_19836,N_19917);
or UO_1128 (O_1128,N_19618,N_19890);
nand UO_1129 (O_1129,N_19926,N_19968);
and UO_1130 (O_1130,N_19777,N_19762);
xor UO_1131 (O_1131,N_19702,N_19761);
xor UO_1132 (O_1132,N_19871,N_19944);
or UO_1133 (O_1133,N_19732,N_19612);
and UO_1134 (O_1134,N_19725,N_19637);
nand UO_1135 (O_1135,N_19938,N_19884);
xor UO_1136 (O_1136,N_19826,N_19799);
xnor UO_1137 (O_1137,N_19677,N_19861);
nor UO_1138 (O_1138,N_19786,N_19763);
and UO_1139 (O_1139,N_19673,N_19662);
nor UO_1140 (O_1140,N_19711,N_19998);
nor UO_1141 (O_1141,N_19669,N_19678);
or UO_1142 (O_1142,N_19697,N_19803);
xor UO_1143 (O_1143,N_19983,N_19685);
or UO_1144 (O_1144,N_19951,N_19741);
nand UO_1145 (O_1145,N_19847,N_19736);
nor UO_1146 (O_1146,N_19636,N_19831);
nand UO_1147 (O_1147,N_19682,N_19622);
nor UO_1148 (O_1148,N_19731,N_19843);
nor UO_1149 (O_1149,N_19658,N_19707);
xnor UO_1150 (O_1150,N_19919,N_19653);
nor UO_1151 (O_1151,N_19961,N_19962);
or UO_1152 (O_1152,N_19986,N_19946);
and UO_1153 (O_1153,N_19828,N_19752);
or UO_1154 (O_1154,N_19901,N_19839);
and UO_1155 (O_1155,N_19622,N_19939);
xnor UO_1156 (O_1156,N_19763,N_19838);
or UO_1157 (O_1157,N_19792,N_19928);
nand UO_1158 (O_1158,N_19628,N_19880);
or UO_1159 (O_1159,N_19750,N_19625);
xnor UO_1160 (O_1160,N_19937,N_19707);
nor UO_1161 (O_1161,N_19676,N_19963);
nand UO_1162 (O_1162,N_19638,N_19878);
xor UO_1163 (O_1163,N_19792,N_19626);
nand UO_1164 (O_1164,N_19680,N_19842);
or UO_1165 (O_1165,N_19891,N_19950);
xnor UO_1166 (O_1166,N_19610,N_19735);
nor UO_1167 (O_1167,N_19952,N_19618);
or UO_1168 (O_1168,N_19975,N_19912);
and UO_1169 (O_1169,N_19624,N_19725);
nand UO_1170 (O_1170,N_19982,N_19640);
xor UO_1171 (O_1171,N_19795,N_19725);
nor UO_1172 (O_1172,N_19700,N_19815);
nand UO_1173 (O_1173,N_19853,N_19630);
and UO_1174 (O_1174,N_19995,N_19925);
and UO_1175 (O_1175,N_19960,N_19729);
or UO_1176 (O_1176,N_19817,N_19922);
xor UO_1177 (O_1177,N_19603,N_19776);
and UO_1178 (O_1178,N_19629,N_19616);
xnor UO_1179 (O_1179,N_19608,N_19978);
nor UO_1180 (O_1180,N_19998,N_19991);
and UO_1181 (O_1181,N_19836,N_19645);
nand UO_1182 (O_1182,N_19860,N_19666);
and UO_1183 (O_1183,N_19816,N_19757);
nand UO_1184 (O_1184,N_19630,N_19739);
or UO_1185 (O_1185,N_19835,N_19633);
nor UO_1186 (O_1186,N_19917,N_19689);
nor UO_1187 (O_1187,N_19655,N_19712);
or UO_1188 (O_1188,N_19935,N_19798);
xor UO_1189 (O_1189,N_19607,N_19709);
nor UO_1190 (O_1190,N_19880,N_19886);
nor UO_1191 (O_1191,N_19998,N_19839);
or UO_1192 (O_1192,N_19748,N_19968);
and UO_1193 (O_1193,N_19810,N_19989);
nand UO_1194 (O_1194,N_19621,N_19792);
or UO_1195 (O_1195,N_19646,N_19616);
and UO_1196 (O_1196,N_19619,N_19690);
xor UO_1197 (O_1197,N_19698,N_19997);
nand UO_1198 (O_1198,N_19912,N_19817);
nand UO_1199 (O_1199,N_19824,N_19677);
nor UO_1200 (O_1200,N_19699,N_19956);
nor UO_1201 (O_1201,N_19753,N_19745);
nand UO_1202 (O_1202,N_19743,N_19873);
and UO_1203 (O_1203,N_19679,N_19754);
nor UO_1204 (O_1204,N_19986,N_19662);
nand UO_1205 (O_1205,N_19933,N_19993);
xor UO_1206 (O_1206,N_19762,N_19774);
xnor UO_1207 (O_1207,N_19664,N_19900);
nand UO_1208 (O_1208,N_19699,N_19846);
or UO_1209 (O_1209,N_19790,N_19750);
and UO_1210 (O_1210,N_19635,N_19713);
nand UO_1211 (O_1211,N_19736,N_19917);
xor UO_1212 (O_1212,N_19702,N_19856);
nor UO_1213 (O_1213,N_19619,N_19958);
nor UO_1214 (O_1214,N_19897,N_19734);
nand UO_1215 (O_1215,N_19743,N_19953);
xor UO_1216 (O_1216,N_19959,N_19755);
or UO_1217 (O_1217,N_19928,N_19902);
xnor UO_1218 (O_1218,N_19786,N_19911);
nor UO_1219 (O_1219,N_19608,N_19866);
xnor UO_1220 (O_1220,N_19916,N_19725);
nor UO_1221 (O_1221,N_19895,N_19699);
and UO_1222 (O_1222,N_19833,N_19715);
nor UO_1223 (O_1223,N_19711,N_19642);
or UO_1224 (O_1224,N_19976,N_19744);
nand UO_1225 (O_1225,N_19696,N_19918);
and UO_1226 (O_1226,N_19839,N_19799);
or UO_1227 (O_1227,N_19862,N_19670);
or UO_1228 (O_1228,N_19978,N_19719);
xor UO_1229 (O_1229,N_19822,N_19667);
and UO_1230 (O_1230,N_19863,N_19634);
nor UO_1231 (O_1231,N_19987,N_19862);
or UO_1232 (O_1232,N_19934,N_19740);
nand UO_1233 (O_1233,N_19835,N_19731);
or UO_1234 (O_1234,N_19750,N_19854);
xnor UO_1235 (O_1235,N_19641,N_19603);
and UO_1236 (O_1236,N_19648,N_19891);
and UO_1237 (O_1237,N_19828,N_19671);
nor UO_1238 (O_1238,N_19755,N_19832);
and UO_1239 (O_1239,N_19858,N_19822);
xnor UO_1240 (O_1240,N_19901,N_19960);
xor UO_1241 (O_1241,N_19823,N_19702);
or UO_1242 (O_1242,N_19771,N_19981);
nand UO_1243 (O_1243,N_19888,N_19758);
or UO_1244 (O_1244,N_19993,N_19934);
nand UO_1245 (O_1245,N_19701,N_19859);
or UO_1246 (O_1246,N_19888,N_19963);
nor UO_1247 (O_1247,N_19797,N_19600);
nor UO_1248 (O_1248,N_19814,N_19718);
nor UO_1249 (O_1249,N_19636,N_19710);
and UO_1250 (O_1250,N_19723,N_19692);
nor UO_1251 (O_1251,N_19933,N_19803);
or UO_1252 (O_1252,N_19897,N_19754);
and UO_1253 (O_1253,N_19776,N_19785);
and UO_1254 (O_1254,N_19763,N_19782);
nor UO_1255 (O_1255,N_19979,N_19613);
nand UO_1256 (O_1256,N_19689,N_19875);
or UO_1257 (O_1257,N_19911,N_19626);
or UO_1258 (O_1258,N_19823,N_19876);
xnor UO_1259 (O_1259,N_19988,N_19919);
xnor UO_1260 (O_1260,N_19632,N_19772);
or UO_1261 (O_1261,N_19829,N_19726);
or UO_1262 (O_1262,N_19744,N_19853);
and UO_1263 (O_1263,N_19678,N_19690);
nand UO_1264 (O_1264,N_19870,N_19806);
xnor UO_1265 (O_1265,N_19857,N_19882);
or UO_1266 (O_1266,N_19669,N_19835);
or UO_1267 (O_1267,N_19960,N_19879);
xnor UO_1268 (O_1268,N_19921,N_19729);
nor UO_1269 (O_1269,N_19655,N_19865);
xnor UO_1270 (O_1270,N_19862,N_19966);
and UO_1271 (O_1271,N_19781,N_19670);
and UO_1272 (O_1272,N_19964,N_19939);
nor UO_1273 (O_1273,N_19769,N_19756);
and UO_1274 (O_1274,N_19813,N_19610);
xnor UO_1275 (O_1275,N_19766,N_19607);
or UO_1276 (O_1276,N_19644,N_19901);
and UO_1277 (O_1277,N_19766,N_19618);
xor UO_1278 (O_1278,N_19795,N_19945);
nand UO_1279 (O_1279,N_19658,N_19963);
and UO_1280 (O_1280,N_19810,N_19875);
or UO_1281 (O_1281,N_19931,N_19699);
and UO_1282 (O_1282,N_19947,N_19811);
xnor UO_1283 (O_1283,N_19957,N_19738);
or UO_1284 (O_1284,N_19889,N_19737);
nand UO_1285 (O_1285,N_19958,N_19656);
xor UO_1286 (O_1286,N_19906,N_19649);
nand UO_1287 (O_1287,N_19987,N_19886);
and UO_1288 (O_1288,N_19920,N_19875);
and UO_1289 (O_1289,N_19928,N_19805);
nor UO_1290 (O_1290,N_19999,N_19711);
nor UO_1291 (O_1291,N_19659,N_19976);
xor UO_1292 (O_1292,N_19640,N_19762);
and UO_1293 (O_1293,N_19772,N_19849);
nor UO_1294 (O_1294,N_19647,N_19797);
nand UO_1295 (O_1295,N_19934,N_19902);
nor UO_1296 (O_1296,N_19987,N_19725);
or UO_1297 (O_1297,N_19941,N_19697);
xnor UO_1298 (O_1298,N_19817,N_19892);
and UO_1299 (O_1299,N_19653,N_19928);
nand UO_1300 (O_1300,N_19909,N_19775);
or UO_1301 (O_1301,N_19769,N_19624);
xnor UO_1302 (O_1302,N_19773,N_19618);
and UO_1303 (O_1303,N_19974,N_19942);
or UO_1304 (O_1304,N_19919,N_19888);
or UO_1305 (O_1305,N_19792,N_19945);
nand UO_1306 (O_1306,N_19951,N_19917);
nand UO_1307 (O_1307,N_19787,N_19980);
nor UO_1308 (O_1308,N_19854,N_19811);
and UO_1309 (O_1309,N_19850,N_19942);
nor UO_1310 (O_1310,N_19746,N_19855);
nor UO_1311 (O_1311,N_19687,N_19806);
and UO_1312 (O_1312,N_19642,N_19752);
nor UO_1313 (O_1313,N_19608,N_19679);
nor UO_1314 (O_1314,N_19970,N_19741);
and UO_1315 (O_1315,N_19659,N_19813);
nand UO_1316 (O_1316,N_19672,N_19835);
xor UO_1317 (O_1317,N_19618,N_19972);
nor UO_1318 (O_1318,N_19956,N_19670);
or UO_1319 (O_1319,N_19625,N_19890);
and UO_1320 (O_1320,N_19779,N_19830);
or UO_1321 (O_1321,N_19744,N_19659);
or UO_1322 (O_1322,N_19791,N_19633);
nand UO_1323 (O_1323,N_19634,N_19962);
or UO_1324 (O_1324,N_19835,N_19890);
xnor UO_1325 (O_1325,N_19672,N_19931);
nand UO_1326 (O_1326,N_19983,N_19758);
or UO_1327 (O_1327,N_19819,N_19897);
and UO_1328 (O_1328,N_19752,N_19976);
and UO_1329 (O_1329,N_19625,N_19925);
and UO_1330 (O_1330,N_19770,N_19623);
nor UO_1331 (O_1331,N_19632,N_19834);
or UO_1332 (O_1332,N_19635,N_19657);
xor UO_1333 (O_1333,N_19882,N_19606);
or UO_1334 (O_1334,N_19836,N_19861);
and UO_1335 (O_1335,N_19752,N_19952);
nor UO_1336 (O_1336,N_19707,N_19727);
and UO_1337 (O_1337,N_19653,N_19707);
or UO_1338 (O_1338,N_19663,N_19855);
or UO_1339 (O_1339,N_19623,N_19879);
nor UO_1340 (O_1340,N_19965,N_19732);
or UO_1341 (O_1341,N_19973,N_19992);
and UO_1342 (O_1342,N_19722,N_19776);
nor UO_1343 (O_1343,N_19966,N_19731);
or UO_1344 (O_1344,N_19644,N_19764);
nand UO_1345 (O_1345,N_19885,N_19829);
nor UO_1346 (O_1346,N_19662,N_19635);
or UO_1347 (O_1347,N_19683,N_19812);
or UO_1348 (O_1348,N_19648,N_19878);
or UO_1349 (O_1349,N_19613,N_19829);
nand UO_1350 (O_1350,N_19735,N_19764);
xnor UO_1351 (O_1351,N_19660,N_19736);
nor UO_1352 (O_1352,N_19709,N_19837);
or UO_1353 (O_1353,N_19888,N_19713);
or UO_1354 (O_1354,N_19648,N_19676);
nand UO_1355 (O_1355,N_19722,N_19748);
xnor UO_1356 (O_1356,N_19771,N_19868);
xnor UO_1357 (O_1357,N_19913,N_19991);
xnor UO_1358 (O_1358,N_19749,N_19960);
or UO_1359 (O_1359,N_19792,N_19757);
nor UO_1360 (O_1360,N_19839,N_19693);
nand UO_1361 (O_1361,N_19730,N_19776);
xor UO_1362 (O_1362,N_19649,N_19699);
and UO_1363 (O_1363,N_19971,N_19604);
and UO_1364 (O_1364,N_19838,N_19921);
or UO_1365 (O_1365,N_19979,N_19668);
nor UO_1366 (O_1366,N_19752,N_19665);
and UO_1367 (O_1367,N_19988,N_19675);
nand UO_1368 (O_1368,N_19938,N_19826);
nand UO_1369 (O_1369,N_19763,N_19669);
or UO_1370 (O_1370,N_19678,N_19624);
and UO_1371 (O_1371,N_19888,N_19773);
and UO_1372 (O_1372,N_19959,N_19668);
nor UO_1373 (O_1373,N_19936,N_19935);
nand UO_1374 (O_1374,N_19690,N_19709);
or UO_1375 (O_1375,N_19798,N_19903);
and UO_1376 (O_1376,N_19610,N_19933);
nor UO_1377 (O_1377,N_19794,N_19856);
and UO_1378 (O_1378,N_19986,N_19769);
nand UO_1379 (O_1379,N_19745,N_19760);
and UO_1380 (O_1380,N_19725,N_19727);
nor UO_1381 (O_1381,N_19943,N_19606);
nand UO_1382 (O_1382,N_19679,N_19717);
and UO_1383 (O_1383,N_19799,N_19881);
xor UO_1384 (O_1384,N_19833,N_19689);
or UO_1385 (O_1385,N_19992,N_19807);
and UO_1386 (O_1386,N_19875,N_19913);
nand UO_1387 (O_1387,N_19793,N_19886);
and UO_1388 (O_1388,N_19639,N_19608);
or UO_1389 (O_1389,N_19955,N_19786);
nand UO_1390 (O_1390,N_19827,N_19788);
and UO_1391 (O_1391,N_19616,N_19751);
xnor UO_1392 (O_1392,N_19633,N_19881);
nor UO_1393 (O_1393,N_19973,N_19695);
and UO_1394 (O_1394,N_19992,N_19757);
or UO_1395 (O_1395,N_19896,N_19605);
nor UO_1396 (O_1396,N_19751,N_19698);
xor UO_1397 (O_1397,N_19667,N_19676);
nor UO_1398 (O_1398,N_19604,N_19993);
xnor UO_1399 (O_1399,N_19744,N_19770);
or UO_1400 (O_1400,N_19749,N_19825);
nand UO_1401 (O_1401,N_19825,N_19873);
xor UO_1402 (O_1402,N_19919,N_19771);
xnor UO_1403 (O_1403,N_19716,N_19985);
nand UO_1404 (O_1404,N_19913,N_19960);
xor UO_1405 (O_1405,N_19994,N_19629);
nor UO_1406 (O_1406,N_19975,N_19788);
xnor UO_1407 (O_1407,N_19794,N_19660);
nand UO_1408 (O_1408,N_19971,N_19742);
xor UO_1409 (O_1409,N_19915,N_19905);
nor UO_1410 (O_1410,N_19706,N_19732);
xnor UO_1411 (O_1411,N_19679,N_19892);
nand UO_1412 (O_1412,N_19809,N_19872);
and UO_1413 (O_1413,N_19654,N_19755);
and UO_1414 (O_1414,N_19991,N_19772);
or UO_1415 (O_1415,N_19841,N_19712);
xnor UO_1416 (O_1416,N_19653,N_19621);
and UO_1417 (O_1417,N_19821,N_19790);
nor UO_1418 (O_1418,N_19886,N_19859);
xor UO_1419 (O_1419,N_19829,N_19787);
and UO_1420 (O_1420,N_19921,N_19917);
nand UO_1421 (O_1421,N_19807,N_19621);
and UO_1422 (O_1422,N_19628,N_19739);
or UO_1423 (O_1423,N_19607,N_19917);
nor UO_1424 (O_1424,N_19952,N_19738);
nor UO_1425 (O_1425,N_19705,N_19884);
and UO_1426 (O_1426,N_19909,N_19839);
nand UO_1427 (O_1427,N_19731,N_19633);
nand UO_1428 (O_1428,N_19906,N_19778);
or UO_1429 (O_1429,N_19762,N_19981);
nand UO_1430 (O_1430,N_19820,N_19966);
nand UO_1431 (O_1431,N_19903,N_19726);
nand UO_1432 (O_1432,N_19966,N_19828);
xnor UO_1433 (O_1433,N_19993,N_19926);
nor UO_1434 (O_1434,N_19652,N_19946);
or UO_1435 (O_1435,N_19645,N_19934);
or UO_1436 (O_1436,N_19661,N_19651);
xor UO_1437 (O_1437,N_19714,N_19838);
nand UO_1438 (O_1438,N_19954,N_19692);
xor UO_1439 (O_1439,N_19821,N_19887);
nor UO_1440 (O_1440,N_19638,N_19684);
xor UO_1441 (O_1441,N_19825,N_19784);
or UO_1442 (O_1442,N_19682,N_19749);
nor UO_1443 (O_1443,N_19868,N_19938);
or UO_1444 (O_1444,N_19801,N_19906);
or UO_1445 (O_1445,N_19797,N_19715);
and UO_1446 (O_1446,N_19621,N_19917);
nor UO_1447 (O_1447,N_19765,N_19776);
or UO_1448 (O_1448,N_19936,N_19913);
xnor UO_1449 (O_1449,N_19926,N_19818);
xnor UO_1450 (O_1450,N_19731,N_19825);
or UO_1451 (O_1451,N_19732,N_19772);
or UO_1452 (O_1452,N_19897,N_19635);
nor UO_1453 (O_1453,N_19693,N_19702);
xnor UO_1454 (O_1454,N_19614,N_19898);
or UO_1455 (O_1455,N_19655,N_19618);
or UO_1456 (O_1456,N_19798,N_19963);
nand UO_1457 (O_1457,N_19741,N_19768);
nor UO_1458 (O_1458,N_19967,N_19928);
nand UO_1459 (O_1459,N_19606,N_19602);
xnor UO_1460 (O_1460,N_19766,N_19966);
and UO_1461 (O_1461,N_19858,N_19824);
nand UO_1462 (O_1462,N_19605,N_19641);
nor UO_1463 (O_1463,N_19971,N_19957);
or UO_1464 (O_1464,N_19800,N_19692);
and UO_1465 (O_1465,N_19878,N_19852);
nor UO_1466 (O_1466,N_19801,N_19847);
or UO_1467 (O_1467,N_19792,N_19603);
xor UO_1468 (O_1468,N_19728,N_19890);
and UO_1469 (O_1469,N_19609,N_19843);
or UO_1470 (O_1470,N_19710,N_19771);
and UO_1471 (O_1471,N_19838,N_19664);
and UO_1472 (O_1472,N_19763,N_19881);
xnor UO_1473 (O_1473,N_19796,N_19910);
and UO_1474 (O_1474,N_19680,N_19974);
nand UO_1475 (O_1475,N_19883,N_19994);
xnor UO_1476 (O_1476,N_19759,N_19921);
nor UO_1477 (O_1477,N_19705,N_19665);
xor UO_1478 (O_1478,N_19701,N_19888);
or UO_1479 (O_1479,N_19749,N_19632);
and UO_1480 (O_1480,N_19656,N_19815);
nor UO_1481 (O_1481,N_19684,N_19752);
and UO_1482 (O_1482,N_19955,N_19921);
nor UO_1483 (O_1483,N_19983,N_19885);
nand UO_1484 (O_1484,N_19610,N_19608);
and UO_1485 (O_1485,N_19884,N_19706);
nor UO_1486 (O_1486,N_19786,N_19784);
and UO_1487 (O_1487,N_19635,N_19913);
nor UO_1488 (O_1488,N_19998,N_19655);
xor UO_1489 (O_1489,N_19675,N_19765);
nor UO_1490 (O_1490,N_19688,N_19696);
xor UO_1491 (O_1491,N_19959,N_19785);
nand UO_1492 (O_1492,N_19655,N_19980);
xnor UO_1493 (O_1493,N_19752,N_19850);
nor UO_1494 (O_1494,N_19618,N_19769);
and UO_1495 (O_1495,N_19687,N_19914);
and UO_1496 (O_1496,N_19606,N_19913);
and UO_1497 (O_1497,N_19799,N_19731);
nor UO_1498 (O_1498,N_19761,N_19940);
nor UO_1499 (O_1499,N_19708,N_19901);
or UO_1500 (O_1500,N_19749,N_19726);
nor UO_1501 (O_1501,N_19848,N_19749);
nor UO_1502 (O_1502,N_19696,N_19871);
nand UO_1503 (O_1503,N_19781,N_19789);
nor UO_1504 (O_1504,N_19730,N_19935);
or UO_1505 (O_1505,N_19698,N_19879);
nand UO_1506 (O_1506,N_19917,N_19772);
or UO_1507 (O_1507,N_19818,N_19955);
or UO_1508 (O_1508,N_19829,N_19786);
nand UO_1509 (O_1509,N_19977,N_19815);
nor UO_1510 (O_1510,N_19664,N_19805);
or UO_1511 (O_1511,N_19862,N_19619);
and UO_1512 (O_1512,N_19999,N_19639);
nor UO_1513 (O_1513,N_19809,N_19660);
and UO_1514 (O_1514,N_19926,N_19919);
or UO_1515 (O_1515,N_19617,N_19640);
or UO_1516 (O_1516,N_19774,N_19914);
xor UO_1517 (O_1517,N_19775,N_19788);
nand UO_1518 (O_1518,N_19655,N_19897);
nand UO_1519 (O_1519,N_19656,N_19602);
nand UO_1520 (O_1520,N_19778,N_19665);
nand UO_1521 (O_1521,N_19670,N_19634);
xor UO_1522 (O_1522,N_19937,N_19938);
xor UO_1523 (O_1523,N_19878,N_19970);
xor UO_1524 (O_1524,N_19615,N_19735);
and UO_1525 (O_1525,N_19734,N_19982);
nor UO_1526 (O_1526,N_19790,N_19694);
and UO_1527 (O_1527,N_19677,N_19768);
or UO_1528 (O_1528,N_19771,N_19791);
and UO_1529 (O_1529,N_19855,N_19715);
or UO_1530 (O_1530,N_19903,N_19869);
or UO_1531 (O_1531,N_19808,N_19926);
nand UO_1532 (O_1532,N_19783,N_19622);
or UO_1533 (O_1533,N_19792,N_19884);
or UO_1534 (O_1534,N_19917,N_19752);
and UO_1535 (O_1535,N_19685,N_19724);
xnor UO_1536 (O_1536,N_19774,N_19612);
nand UO_1537 (O_1537,N_19717,N_19946);
or UO_1538 (O_1538,N_19625,N_19955);
and UO_1539 (O_1539,N_19666,N_19703);
nor UO_1540 (O_1540,N_19864,N_19770);
nand UO_1541 (O_1541,N_19636,N_19808);
nand UO_1542 (O_1542,N_19946,N_19949);
nand UO_1543 (O_1543,N_19991,N_19883);
or UO_1544 (O_1544,N_19624,N_19910);
xnor UO_1545 (O_1545,N_19951,N_19768);
nand UO_1546 (O_1546,N_19817,N_19644);
nand UO_1547 (O_1547,N_19621,N_19772);
xnor UO_1548 (O_1548,N_19675,N_19766);
nand UO_1549 (O_1549,N_19885,N_19946);
or UO_1550 (O_1550,N_19753,N_19676);
or UO_1551 (O_1551,N_19834,N_19993);
and UO_1552 (O_1552,N_19820,N_19881);
and UO_1553 (O_1553,N_19634,N_19640);
and UO_1554 (O_1554,N_19988,N_19719);
nor UO_1555 (O_1555,N_19846,N_19653);
nor UO_1556 (O_1556,N_19873,N_19734);
nor UO_1557 (O_1557,N_19866,N_19712);
xor UO_1558 (O_1558,N_19748,N_19982);
xor UO_1559 (O_1559,N_19933,N_19924);
xor UO_1560 (O_1560,N_19863,N_19959);
and UO_1561 (O_1561,N_19647,N_19887);
and UO_1562 (O_1562,N_19730,N_19875);
xnor UO_1563 (O_1563,N_19849,N_19907);
xnor UO_1564 (O_1564,N_19600,N_19940);
nor UO_1565 (O_1565,N_19675,N_19617);
nand UO_1566 (O_1566,N_19787,N_19739);
and UO_1567 (O_1567,N_19995,N_19662);
and UO_1568 (O_1568,N_19835,N_19856);
or UO_1569 (O_1569,N_19639,N_19900);
xnor UO_1570 (O_1570,N_19818,N_19674);
nor UO_1571 (O_1571,N_19993,N_19764);
and UO_1572 (O_1572,N_19896,N_19935);
and UO_1573 (O_1573,N_19997,N_19663);
nand UO_1574 (O_1574,N_19843,N_19780);
nand UO_1575 (O_1575,N_19674,N_19698);
xor UO_1576 (O_1576,N_19860,N_19803);
or UO_1577 (O_1577,N_19885,N_19770);
nor UO_1578 (O_1578,N_19614,N_19973);
nor UO_1579 (O_1579,N_19914,N_19651);
or UO_1580 (O_1580,N_19684,N_19827);
nand UO_1581 (O_1581,N_19765,N_19825);
nor UO_1582 (O_1582,N_19965,N_19828);
or UO_1583 (O_1583,N_19994,N_19957);
nor UO_1584 (O_1584,N_19758,N_19895);
and UO_1585 (O_1585,N_19768,N_19777);
nand UO_1586 (O_1586,N_19951,N_19865);
nor UO_1587 (O_1587,N_19928,N_19837);
xor UO_1588 (O_1588,N_19864,N_19732);
or UO_1589 (O_1589,N_19671,N_19707);
or UO_1590 (O_1590,N_19976,N_19678);
or UO_1591 (O_1591,N_19978,N_19842);
xor UO_1592 (O_1592,N_19842,N_19916);
and UO_1593 (O_1593,N_19611,N_19786);
nand UO_1594 (O_1594,N_19840,N_19746);
or UO_1595 (O_1595,N_19810,N_19707);
nor UO_1596 (O_1596,N_19939,N_19738);
xor UO_1597 (O_1597,N_19678,N_19845);
or UO_1598 (O_1598,N_19808,N_19803);
and UO_1599 (O_1599,N_19960,N_19786);
nand UO_1600 (O_1600,N_19883,N_19727);
and UO_1601 (O_1601,N_19832,N_19798);
or UO_1602 (O_1602,N_19691,N_19967);
xnor UO_1603 (O_1603,N_19821,N_19949);
nand UO_1604 (O_1604,N_19643,N_19976);
xnor UO_1605 (O_1605,N_19878,N_19980);
or UO_1606 (O_1606,N_19964,N_19914);
xor UO_1607 (O_1607,N_19762,N_19991);
or UO_1608 (O_1608,N_19709,N_19885);
or UO_1609 (O_1609,N_19832,N_19670);
xnor UO_1610 (O_1610,N_19606,N_19807);
and UO_1611 (O_1611,N_19626,N_19657);
xnor UO_1612 (O_1612,N_19717,N_19859);
nand UO_1613 (O_1613,N_19678,N_19955);
or UO_1614 (O_1614,N_19800,N_19948);
xnor UO_1615 (O_1615,N_19668,N_19675);
nor UO_1616 (O_1616,N_19778,N_19711);
or UO_1617 (O_1617,N_19839,N_19919);
nor UO_1618 (O_1618,N_19945,N_19946);
xnor UO_1619 (O_1619,N_19694,N_19867);
nor UO_1620 (O_1620,N_19774,N_19663);
and UO_1621 (O_1621,N_19849,N_19675);
or UO_1622 (O_1622,N_19841,N_19904);
or UO_1623 (O_1623,N_19656,N_19997);
nand UO_1624 (O_1624,N_19824,N_19881);
and UO_1625 (O_1625,N_19918,N_19956);
or UO_1626 (O_1626,N_19924,N_19910);
nor UO_1627 (O_1627,N_19677,N_19899);
and UO_1628 (O_1628,N_19949,N_19678);
xnor UO_1629 (O_1629,N_19939,N_19951);
nand UO_1630 (O_1630,N_19992,N_19798);
and UO_1631 (O_1631,N_19693,N_19928);
nand UO_1632 (O_1632,N_19942,N_19921);
xnor UO_1633 (O_1633,N_19846,N_19691);
xnor UO_1634 (O_1634,N_19714,N_19966);
xor UO_1635 (O_1635,N_19851,N_19673);
and UO_1636 (O_1636,N_19814,N_19606);
xnor UO_1637 (O_1637,N_19609,N_19724);
xnor UO_1638 (O_1638,N_19977,N_19901);
xnor UO_1639 (O_1639,N_19858,N_19661);
or UO_1640 (O_1640,N_19727,N_19670);
or UO_1641 (O_1641,N_19625,N_19753);
nand UO_1642 (O_1642,N_19829,N_19773);
nor UO_1643 (O_1643,N_19846,N_19780);
or UO_1644 (O_1644,N_19980,N_19992);
and UO_1645 (O_1645,N_19921,N_19847);
nor UO_1646 (O_1646,N_19872,N_19634);
nand UO_1647 (O_1647,N_19670,N_19889);
or UO_1648 (O_1648,N_19747,N_19703);
or UO_1649 (O_1649,N_19696,N_19914);
nor UO_1650 (O_1650,N_19793,N_19985);
nor UO_1651 (O_1651,N_19991,N_19647);
nand UO_1652 (O_1652,N_19942,N_19859);
and UO_1653 (O_1653,N_19852,N_19780);
and UO_1654 (O_1654,N_19946,N_19719);
nor UO_1655 (O_1655,N_19731,N_19963);
nand UO_1656 (O_1656,N_19844,N_19876);
nand UO_1657 (O_1657,N_19677,N_19601);
and UO_1658 (O_1658,N_19915,N_19670);
xor UO_1659 (O_1659,N_19749,N_19763);
and UO_1660 (O_1660,N_19793,N_19935);
xor UO_1661 (O_1661,N_19719,N_19736);
nor UO_1662 (O_1662,N_19758,N_19978);
nand UO_1663 (O_1663,N_19781,N_19877);
and UO_1664 (O_1664,N_19747,N_19711);
nand UO_1665 (O_1665,N_19725,N_19814);
and UO_1666 (O_1666,N_19608,N_19825);
nor UO_1667 (O_1667,N_19895,N_19753);
xor UO_1668 (O_1668,N_19949,N_19967);
and UO_1669 (O_1669,N_19727,N_19969);
or UO_1670 (O_1670,N_19746,N_19803);
and UO_1671 (O_1671,N_19977,N_19953);
and UO_1672 (O_1672,N_19919,N_19729);
nand UO_1673 (O_1673,N_19750,N_19692);
nor UO_1674 (O_1674,N_19705,N_19743);
xor UO_1675 (O_1675,N_19795,N_19836);
nand UO_1676 (O_1676,N_19965,N_19604);
nand UO_1677 (O_1677,N_19624,N_19937);
nand UO_1678 (O_1678,N_19763,N_19761);
and UO_1679 (O_1679,N_19764,N_19750);
nor UO_1680 (O_1680,N_19950,N_19641);
xnor UO_1681 (O_1681,N_19878,N_19759);
xor UO_1682 (O_1682,N_19716,N_19761);
nand UO_1683 (O_1683,N_19825,N_19753);
nand UO_1684 (O_1684,N_19746,N_19946);
and UO_1685 (O_1685,N_19795,N_19838);
nor UO_1686 (O_1686,N_19944,N_19838);
nand UO_1687 (O_1687,N_19754,N_19856);
nor UO_1688 (O_1688,N_19745,N_19781);
nand UO_1689 (O_1689,N_19944,N_19880);
or UO_1690 (O_1690,N_19605,N_19733);
nor UO_1691 (O_1691,N_19796,N_19669);
nand UO_1692 (O_1692,N_19908,N_19725);
nand UO_1693 (O_1693,N_19731,N_19845);
xor UO_1694 (O_1694,N_19636,N_19751);
or UO_1695 (O_1695,N_19980,N_19911);
nand UO_1696 (O_1696,N_19962,N_19902);
xnor UO_1697 (O_1697,N_19606,N_19768);
and UO_1698 (O_1698,N_19725,N_19840);
xnor UO_1699 (O_1699,N_19714,N_19603);
nand UO_1700 (O_1700,N_19670,N_19660);
nor UO_1701 (O_1701,N_19718,N_19664);
nor UO_1702 (O_1702,N_19941,N_19721);
and UO_1703 (O_1703,N_19730,N_19840);
and UO_1704 (O_1704,N_19806,N_19738);
xor UO_1705 (O_1705,N_19760,N_19696);
and UO_1706 (O_1706,N_19916,N_19696);
or UO_1707 (O_1707,N_19973,N_19854);
and UO_1708 (O_1708,N_19748,N_19676);
and UO_1709 (O_1709,N_19792,N_19646);
xor UO_1710 (O_1710,N_19792,N_19687);
nand UO_1711 (O_1711,N_19755,N_19692);
or UO_1712 (O_1712,N_19830,N_19790);
nor UO_1713 (O_1713,N_19878,N_19789);
nor UO_1714 (O_1714,N_19606,N_19813);
and UO_1715 (O_1715,N_19910,N_19672);
and UO_1716 (O_1716,N_19982,N_19618);
nor UO_1717 (O_1717,N_19924,N_19601);
nand UO_1718 (O_1718,N_19856,N_19655);
nor UO_1719 (O_1719,N_19886,N_19750);
and UO_1720 (O_1720,N_19757,N_19963);
and UO_1721 (O_1721,N_19636,N_19884);
nor UO_1722 (O_1722,N_19808,N_19928);
xnor UO_1723 (O_1723,N_19858,N_19713);
nor UO_1724 (O_1724,N_19760,N_19927);
nor UO_1725 (O_1725,N_19976,N_19870);
and UO_1726 (O_1726,N_19843,N_19933);
or UO_1727 (O_1727,N_19915,N_19931);
nand UO_1728 (O_1728,N_19643,N_19857);
and UO_1729 (O_1729,N_19996,N_19770);
nand UO_1730 (O_1730,N_19793,N_19951);
nor UO_1731 (O_1731,N_19875,N_19975);
nand UO_1732 (O_1732,N_19778,N_19606);
nand UO_1733 (O_1733,N_19618,N_19880);
xnor UO_1734 (O_1734,N_19897,N_19924);
and UO_1735 (O_1735,N_19721,N_19892);
nand UO_1736 (O_1736,N_19607,N_19824);
xor UO_1737 (O_1737,N_19742,N_19686);
nand UO_1738 (O_1738,N_19837,N_19899);
nand UO_1739 (O_1739,N_19825,N_19865);
nor UO_1740 (O_1740,N_19681,N_19695);
xnor UO_1741 (O_1741,N_19724,N_19822);
nand UO_1742 (O_1742,N_19886,N_19986);
or UO_1743 (O_1743,N_19608,N_19788);
nor UO_1744 (O_1744,N_19886,N_19701);
nand UO_1745 (O_1745,N_19847,N_19692);
xor UO_1746 (O_1746,N_19979,N_19624);
or UO_1747 (O_1747,N_19706,N_19825);
xor UO_1748 (O_1748,N_19824,N_19853);
xnor UO_1749 (O_1749,N_19929,N_19945);
nand UO_1750 (O_1750,N_19922,N_19739);
or UO_1751 (O_1751,N_19633,N_19796);
nor UO_1752 (O_1752,N_19829,N_19895);
xor UO_1753 (O_1753,N_19975,N_19806);
and UO_1754 (O_1754,N_19737,N_19739);
nor UO_1755 (O_1755,N_19869,N_19967);
xor UO_1756 (O_1756,N_19835,N_19902);
and UO_1757 (O_1757,N_19863,N_19912);
nand UO_1758 (O_1758,N_19900,N_19909);
and UO_1759 (O_1759,N_19854,N_19883);
and UO_1760 (O_1760,N_19836,N_19823);
nor UO_1761 (O_1761,N_19794,N_19942);
and UO_1762 (O_1762,N_19991,N_19777);
nand UO_1763 (O_1763,N_19844,N_19809);
xnor UO_1764 (O_1764,N_19734,N_19659);
xnor UO_1765 (O_1765,N_19630,N_19629);
and UO_1766 (O_1766,N_19876,N_19635);
nor UO_1767 (O_1767,N_19782,N_19941);
nand UO_1768 (O_1768,N_19629,N_19618);
nand UO_1769 (O_1769,N_19684,N_19674);
and UO_1770 (O_1770,N_19668,N_19605);
or UO_1771 (O_1771,N_19805,N_19959);
and UO_1772 (O_1772,N_19834,N_19674);
nand UO_1773 (O_1773,N_19615,N_19944);
and UO_1774 (O_1774,N_19694,N_19794);
or UO_1775 (O_1775,N_19659,N_19995);
nand UO_1776 (O_1776,N_19794,N_19811);
or UO_1777 (O_1777,N_19965,N_19767);
nand UO_1778 (O_1778,N_19978,N_19658);
xnor UO_1779 (O_1779,N_19739,N_19909);
and UO_1780 (O_1780,N_19746,N_19958);
xor UO_1781 (O_1781,N_19749,N_19629);
nand UO_1782 (O_1782,N_19605,N_19945);
and UO_1783 (O_1783,N_19874,N_19633);
and UO_1784 (O_1784,N_19977,N_19894);
or UO_1785 (O_1785,N_19920,N_19740);
or UO_1786 (O_1786,N_19984,N_19889);
nor UO_1787 (O_1787,N_19613,N_19762);
nand UO_1788 (O_1788,N_19837,N_19947);
xnor UO_1789 (O_1789,N_19925,N_19845);
nand UO_1790 (O_1790,N_19697,N_19729);
nand UO_1791 (O_1791,N_19922,N_19665);
and UO_1792 (O_1792,N_19950,N_19966);
and UO_1793 (O_1793,N_19752,N_19657);
xor UO_1794 (O_1794,N_19652,N_19748);
and UO_1795 (O_1795,N_19890,N_19643);
nand UO_1796 (O_1796,N_19616,N_19847);
xnor UO_1797 (O_1797,N_19744,N_19719);
or UO_1798 (O_1798,N_19707,N_19907);
xor UO_1799 (O_1799,N_19793,N_19856);
xnor UO_1800 (O_1800,N_19835,N_19837);
or UO_1801 (O_1801,N_19680,N_19925);
or UO_1802 (O_1802,N_19723,N_19957);
xnor UO_1803 (O_1803,N_19692,N_19984);
xor UO_1804 (O_1804,N_19664,N_19642);
xor UO_1805 (O_1805,N_19821,N_19978);
nand UO_1806 (O_1806,N_19833,N_19937);
nor UO_1807 (O_1807,N_19819,N_19741);
nor UO_1808 (O_1808,N_19932,N_19993);
and UO_1809 (O_1809,N_19967,N_19953);
and UO_1810 (O_1810,N_19845,N_19729);
nor UO_1811 (O_1811,N_19840,N_19900);
nand UO_1812 (O_1812,N_19940,N_19914);
and UO_1813 (O_1813,N_19985,N_19892);
or UO_1814 (O_1814,N_19949,N_19754);
and UO_1815 (O_1815,N_19862,N_19621);
nand UO_1816 (O_1816,N_19763,N_19865);
nor UO_1817 (O_1817,N_19826,N_19683);
and UO_1818 (O_1818,N_19742,N_19897);
nand UO_1819 (O_1819,N_19981,N_19918);
and UO_1820 (O_1820,N_19709,N_19861);
xor UO_1821 (O_1821,N_19993,N_19880);
or UO_1822 (O_1822,N_19820,N_19744);
nand UO_1823 (O_1823,N_19863,N_19907);
and UO_1824 (O_1824,N_19838,N_19905);
xnor UO_1825 (O_1825,N_19987,N_19683);
nor UO_1826 (O_1826,N_19637,N_19675);
or UO_1827 (O_1827,N_19797,N_19633);
nand UO_1828 (O_1828,N_19829,N_19865);
nand UO_1829 (O_1829,N_19715,N_19969);
xnor UO_1830 (O_1830,N_19865,N_19827);
and UO_1831 (O_1831,N_19729,N_19818);
or UO_1832 (O_1832,N_19931,N_19765);
and UO_1833 (O_1833,N_19795,N_19785);
nand UO_1834 (O_1834,N_19643,N_19736);
nor UO_1835 (O_1835,N_19600,N_19729);
nor UO_1836 (O_1836,N_19831,N_19748);
and UO_1837 (O_1837,N_19993,N_19870);
nor UO_1838 (O_1838,N_19645,N_19992);
nor UO_1839 (O_1839,N_19655,N_19715);
or UO_1840 (O_1840,N_19936,N_19843);
or UO_1841 (O_1841,N_19775,N_19867);
nand UO_1842 (O_1842,N_19623,N_19760);
nand UO_1843 (O_1843,N_19954,N_19691);
xnor UO_1844 (O_1844,N_19667,N_19833);
xor UO_1845 (O_1845,N_19754,N_19862);
xor UO_1846 (O_1846,N_19966,N_19735);
or UO_1847 (O_1847,N_19986,N_19804);
or UO_1848 (O_1848,N_19706,N_19651);
nor UO_1849 (O_1849,N_19840,N_19886);
or UO_1850 (O_1850,N_19638,N_19618);
nor UO_1851 (O_1851,N_19782,N_19986);
xnor UO_1852 (O_1852,N_19701,N_19935);
nand UO_1853 (O_1853,N_19635,N_19972);
xnor UO_1854 (O_1854,N_19612,N_19910);
and UO_1855 (O_1855,N_19774,N_19824);
nand UO_1856 (O_1856,N_19718,N_19717);
nor UO_1857 (O_1857,N_19769,N_19891);
or UO_1858 (O_1858,N_19622,N_19665);
nand UO_1859 (O_1859,N_19892,N_19774);
xnor UO_1860 (O_1860,N_19898,N_19776);
nand UO_1861 (O_1861,N_19745,N_19772);
nand UO_1862 (O_1862,N_19984,N_19939);
or UO_1863 (O_1863,N_19669,N_19655);
xor UO_1864 (O_1864,N_19702,N_19642);
xor UO_1865 (O_1865,N_19724,N_19674);
nand UO_1866 (O_1866,N_19667,N_19885);
nand UO_1867 (O_1867,N_19934,N_19898);
or UO_1868 (O_1868,N_19639,N_19877);
nor UO_1869 (O_1869,N_19818,N_19716);
and UO_1870 (O_1870,N_19886,N_19946);
nor UO_1871 (O_1871,N_19695,N_19647);
xor UO_1872 (O_1872,N_19860,N_19875);
or UO_1873 (O_1873,N_19646,N_19706);
or UO_1874 (O_1874,N_19622,N_19612);
nand UO_1875 (O_1875,N_19726,N_19652);
nor UO_1876 (O_1876,N_19780,N_19979);
or UO_1877 (O_1877,N_19816,N_19655);
xor UO_1878 (O_1878,N_19758,N_19955);
or UO_1879 (O_1879,N_19805,N_19913);
or UO_1880 (O_1880,N_19602,N_19672);
xnor UO_1881 (O_1881,N_19682,N_19991);
xnor UO_1882 (O_1882,N_19938,N_19963);
nor UO_1883 (O_1883,N_19760,N_19732);
nand UO_1884 (O_1884,N_19925,N_19880);
nand UO_1885 (O_1885,N_19603,N_19818);
xnor UO_1886 (O_1886,N_19932,N_19721);
nor UO_1887 (O_1887,N_19933,N_19668);
nor UO_1888 (O_1888,N_19797,N_19790);
xnor UO_1889 (O_1889,N_19618,N_19786);
xnor UO_1890 (O_1890,N_19790,N_19722);
nor UO_1891 (O_1891,N_19604,N_19853);
nand UO_1892 (O_1892,N_19799,N_19941);
xnor UO_1893 (O_1893,N_19970,N_19679);
nand UO_1894 (O_1894,N_19675,N_19949);
nand UO_1895 (O_1895,N_19778,N_19672);
or UO_1896 (O_1896,N_19852,N_19760);
or UO_1897 (O_1897,N_19964,N_19834);
nand UO_1898 (O_1898,N_19651,N_19948);
or UO_1899 (O_1899,N_19972,N_19934);
xor UO_1900 (O_1900,N_19773,N_19831);
and UO_1901 (O_1901,N_19644,N_19981);
xnor UO_1902 (O_1902,N_19786,N_19624);
nand UO_1903 (O_1903,N_19806,N_19895);
xnor UO_1904 (O_1904,N_19654,N_19809);
xor UO_1905 (O_1905,N_19924,N_19956);
xnor UO_1906 (O_1906,N_19772,N_19636);
or UO_1907 (O_1907,N_19629,N_19854);
nand UO_1908 (O_1908,N_19776,N_19781);
xnor UO_1909 (O_1909,N_19863,N_19673);
or UO_1910 (O_1910,N_19884,N_19817);
nor UO_1911 (O_1911,N_19935,N_19808);
nand UO_1912 (O_1912,N_19902,N_19688);
xor UO_1913 (O_1913,N_19937,N_19988);
or UO_1914 (O_1914,N_19633,N_19806);
nand UO_1915 (O_1915,N_19913,N_19898);
nor UO_1916 (O_1916,N_19855,N_19980);
or UO_1917 (O_1917,N_19813,N_19832);
nand UO_1918 (O_1918,N_19939,N_19687);
xor UO_1919 (O_1919,N_19683,N_19982);
or UO_1920 (O_1920,N_19829,N_19924);
nor UO_1921 (O_1921,N_19739,N_19771);
nor UO_1922 (O_1922,N_19958,N_19733);
xor UO_1923 (O_1923,N_19823,N_19817);
nor UO_1924 (O_1924,N_19695,N_19924);
and UO_1925 (O_1925,N_19794,N_19970);
or UO_1926 (O_1926,N_19766,N_19604);
nand UO_1927 (O_1927,N_19635,N_19640);
or UO_1928 (O_1928,N_19716,N_19629);
or UO_1929 (O_1929,N_19778,N_19865);
nor UO_1930 (O_1930,N_19955,N_19672);
nand UO_1931 (O_1931,N_19877,N_19899);
and UO_1932 (O_1932,N_19860,N_19778);
nor UO_1933 (O_1933,N_19866,N_19630);
nand UO_1934 (O_1934,N_19820,N_19607);
nor UO_1935 (O_1935,N_19992,N_19744);
and UO_1936 (O_1936,N_19951,N_19808);
nand UO_1937 (O_1937,N_19795,N_19787);
or UO_1938 (O_1938,N_19752,N_19857);
nand UO_1939 (O_1939,N_19613,N_19704);
or UO_1940 (O_1940,N_19667,N_19812);
nor UO_1941 (O_1941,N_19910,N_19881);
nand UO_1942 (O_1942,N_19869,N_19839);
nand UO_1943 (O_1943,N_19986,N_19654);
nor UO_1944 (O_1944,N_19604,N_19906);
nor UO_1945 (O_1945,N_19785,N_19823);
nand UO_1946 (O_1946,N_19818,N_19725);
nand UO_1947 (O_1947,N_19970,N_19880);
xor UO_1948 (O_1948,N_19631,N_19628);
xnor UO_1949 (O_1949,N_19903,N_19949);
and UO_1950 (O_1950,N_19637,N_19975);
nor UO_1951 (O_1951,N_19781,N_19764);
nand UO_1952 (O_1952,N_19910,N_19610);
and UO_1953 (O_1953,N_19766,N_19864);
nand UO_1954 (O_1954,N_19712,N_19720);
and UO_1955 (O_1955,N_19875,N_19677);
xor UO_1956 (O_1956,N_19644,N_19815);
nand UO_1957 (O_1957,N_19688,N_19934);
xnor UO_1958 (O_1958,N_19969,N_19700);
and UO_1959 (O_1959,N_19972,N_19695);
nor UO_1960 (O_1960,N_19765,N_19955);
nor UO_1961 (O_1961,N_19636,N_19902);
nand UO_1962 (O_1962,N_19983,N_19849);
xnor UO_1963 (O_1963,N_19978,N_19656);
xnor UO_1964 (O_1964,N_19824,N_19930);
nor UO_1965 (O_1965,N_19937,N_19993);
or UO_1966 (O_1966,N_19629,N_19932);
or UO_1967 (O_1967,N_19704,N_19628);
or UO_1968 (O_1968,N_19937,N_19804);
and UO_1969 (O_1969,N_19876,N_19631);
xnor UO_1970 (O_1970,N_19853,N_19740);
or UO_1971 (O_1971,N_19605,N_19984);
and UO_1972 (O_1972,N_19606,N_19772);
nand UO_1973 (O_1973,N_19993,N_19802);
nand UO_1974 (O_1974,N_19927,N_19905);
nor UO_1975 (O_1975,N_19780,N_19753);
xnor UO_1976 (O_1976,N_19815,N_19978);
and UO_1977 (O_1977,N_19806,N_19691);
and UO_1978 (O_1978,N_19767,N_19843);
nand UO_1979 (O_1979,N_19866,N_19864);
xnor UO_1980 (O_1980,N_19747,N_19855);
xor UO_1981 (O_1981,N_19743,N_19848);
nand UO_1982 (O_1982,N_19692,N_19655);
and UO_1983 (O_1983,N_19765,N_19712);
or UO_1984 (O_1984,N_19979,N_19631);
nor UO_1985 (O_1985,N_19793,N_19637);
nor UO_1986 (O_1986,N_19791,N_19971);
and UO_1987 (O_1987,N_19780,N_19718);
nand UO_1988 (O_1988,N_19798,N_19901);
and UO_1989 (O_1989,N_19716,N_19791);
nor UO_1990 (O_1990,N_19872,N_19615);
xor UO_1991 (O_1991,N_19711,N_19627);
xnor UO_1992 (O_1992,N_19747,N_19775);
xnor UO_1993 (O_1993,N_19977,N_19681);
nor UO_1994 (O_1994,N_19712,N_19626);
nand UO_1995 (O_1995,N_19956,N_19999);
nor UO_1996 (O_1996,N_19885,N_19828);
nor UO_1997 (O_1997,N_19791,N_19891);
nand UO_1998 (O_1998,N_19951,N_19947);
and UO_1999 (O_1999,N_19862,N_19699);
or UO_2000 (O_2000,N_19830,N_19815);
nor UO_2001 (O_2001,N_19894,N_19743);
xnor UO_2002 (O_2002,N_19882,N_19861);
nor UO_2003 (O_2003,N_19934,N_19636);
or UO_2004 (O_2004,N_19701,N_19777);
xnor UO_2005 (O_2005,N_19853,N_19755);
and UO_2006 (O_2006,N_19671,N_19823);
and UO_2007 (O_2007,N_19732,N_19762);
xor UO_2008 (O_2008,N_19988,N_19995);
xnor UO_2009 (O_2009,N_19935,N_19729);
xor UO_2010 (O_2010,N_19838,N_19702);
xnor UO_2011 (O_2011,N_19959,N_19706);
nor UO_2012 (O_2012,N_19690,N_19911);
and UO_2013 (O_2013,N_19731,N_19647);
or UO_2014 (O_2014,N_19688,N_19978);
or UO_2015 (O_2015,N_19633,N_19663);
xor UO_2016 (O_2016,N_19666,N_19895);
nor UO_2017 (O_2017,N_19842,N_19879);
xor UO_2018 (O_2018,N_19959,N_19946);
or UO_2019 (O_2019,N_19788,N_19853);
nand UO_2020 (O_2020,N_19637,N_19991);
xnor UO_2021 (O_2021,N_19806,N_19668);
nand UO_2022 (O_2022,N_19656,N_19991);
xor UO_2023 (O_2023,N_19615,N_19957);
nor UO_2024 (O_2024,N_19615,N_19865);
or UO_2025 (O_2025,N_19809,N_19804);
xnor UO_2026 (O_2026,N_19810,N_19785);
nand UO_2027 (O_2027,N_19641,N_19635);
xor UO_2028 (O_2028,N_19666,N_19840);
nand UO_2029 (O_2029,N_19973,N_19627);
nand UO_2030 (O_2030,N_19780,N_19648);
or UO_2031 (O_2031,N_19972,N_19786);
xnor UO_2032 (O_2032,N_19713,N_19714);
xor UO_2033 (O_2033,N_19922,N_19992);
or UO_2034 (O_2034,N_19866,N_19707);
or UO_2035 (O_2035,N_19688,N_19643);
xnor UO_2036 (O_2036,N_19784,N_19862);
xor UO_2037 (O_2037,N_19976,N_19918);
and UO_2038 (O_2038,N_19867,N_19937);
or UO_2039 (O_2039,N_19825,N_19820);
nand UO_2040 (O_2040,N_19692,N_19794);
and UO_2041 (O_2041,N_19601,N_19976);
nor UO_2042 (O_2042,N_19865,N_19600);
xor UO_2043 (O_2043,N_19621,N_19754);
and UO_2044 (O_2044,N_19929,N_19604);
nor UO_2045 (O_2045,N_19712,N_19603);
nor UO_2046 (O_2046,N_19948,N_19976);
nor UO_2047 (O_2047,N_19815,N_19747);
or UO_2048 (O_2048,N_19658,N_19775);
nor UO_2049 (O_2049,N_19730,N_19805);
or UO_2050 (O_2050,N_19982,N_19774);
or UO_2051 (O_2051,N_19975,N_19921);
nor UO_2052 (O_2052,N_19975,N_19885);
nor UO_2053 (O_2053,N_19916,N_19744);
or UO_2054 (O_2054,N_19759,N_19857);
nor UO_2055 (O_2055,N_19657,N_19751);
or UO_2056 (O_2056,N_19999,N_19719);
nand UO_2057 (O_2057,N_19795,N_19932);
xor UO_2058 (O_2058,N_19837,N_19666);
nand UO_2059 (O_2059,N_19877,N_19912);
or UO_2060 (O_2060,N_19655,N_19757);
xor UO_2061 (O_2061,N_19728,N_19614);
or UO_2062 (O_2062,N_19615,N_19833);
nor UO_2063 (O_2063,N_19947,N_19862);
and UO_2064 (O_2064,N_19617,N_19945);
nand UO_2065 (O_2065,N_19649,N_19728);
nand UO_2066 (O_2066,N_19832,N_19630);
nor UO_2067 (O_2067,N_19843,N_19814);
and UO_2068 (O_2068,N_19942,N_19996);
xor UO_2069 (O_2069,N_19767,N_19682);
nand UO_2070 (O_2070,N_19875,N_19716);
or UO_2071 (O_2071,N_19771,N_19873);
or UO_2072 (O_2072,N_19970,N_19968);
or UO_2073 (O_2073,N_19882,N_19704);
and UO_2074 (O_2074,N_19713,N_19813);
nor UO_2075 (O_2075,N_19695,N_19974);
and UO_2076 (O_2076,N_19759,N_19808);
and UO_2077 (O_2077,N_19835,N_19639);
nand UO_2078 (O_2078,N_19650,N_19949);
nand UO_2079 (O_2079,N_19713,N_19784);
nand UO_2080 (O_2080,N_19856,N_19725);
nor UO_2081 (O_2081,N_19613,N_19969);
nor UO_2082 (O_2082,N_19912,N_19906);
nor UO_2083 (O_2083,N_19806,N_19971);
and UO_2084 (O_2084,N_19872,N_19662);
or UO_2085 (O_2085,N_19793,N_19903);
xor UO_2086 (O_2086,N_19979,N_19990);
nor UO_2087 (O_2087,N_19919,N_19660);
nand UO_2088 (O_2088,N_19608,N_19994);
nor UO_2089 (O_2089,N_19958,N_19611);
nand UO_2090 (O_2090,N_19767,N_19935);
and UO_2091 (O_2091,N_19860,N_19826);
and UO_2092 (O_2092,N_19751,N_19863);
nor UO_2093 (O_2093,N_19879,N_19806);
xnor UO_2094 (O_2094,N_19994,N_19894);
and UO_2095 (O_2095,N_19764,N_19886);
or UO_2096 (O_2096,N_19759,N_19797);
xnor UO_2097 (O_2097,N_19946,N_19769);
and UO_2098 (O_2098,N_19926,N_19638);
or UO_2099 (O_2099,N_19726,N_19792);
nand UO_2100 (O_2100,N_19645,N_19990);
or UO_2101 (O_2101,N_19943,N_19925);
or UO_2102 (O_2102,N_19975,N_19923);
nor UO_2103 (O_2103,N_19671,N_19963);
nand UO_2104 (O_2104,N_19843,N_19976);
nand UO_2105 (O_2105,N_19956,N_19798);
xnor UO_2106 (O_2106,N_19872,N_19898);
xnor UO_2107 (O_2107,N_19885,N_19962);
xnor UO_2108 (O_2108,N_19747,N_19780);
xnor UO_2109 (O_2109,N_19738,N_19768);
or UO_2110 (O_2110,N_19747,N_19853);
nor UO_2111 (O_2111,N_19753,N_19756);
nor UO_2112 (O_2112,N_19690,N_19794);
nand UO_2113 (O_2113,N_19966,N_19665);
or UO_2114 (O_2114,N_19836,N_19940);
and UO_2115 (O_2115,N_19627,N_19708);
or UO_2116 (O_2116,N_19964,N_19891);
xnor UO_2117 (O_2117,N_19952,N_19913);
xor UO_2118 (O_2118,N_19736,N_19838);
nand UO_2119 (O_2119,N_19943,N_19920);
xnor UO_2120 (O_2120,N_19746,N_19736);
or UO_2121 (O_2121,N_19981,N_19733);
and UO_2122 (O_2122,N_19665,N_19795);
and UO_2123 (O_2123,N_19945,N_19927);
nor UO_2124 (O_2124,N_19711,N_19825);
nand UO_2125 (O_2125,N_19990,N_19977);
nor UO_2126 (O_2126,N_19841,N_19817);
nor UO_2127 (O_2127,N_19913,N_19854);
nand UO_2128 (O_2128,N_19619,N_19740);
or UO_2129 (O_2129,N_19918,N_19768);
or UO_2130 (O_2130,N_19811,N_19828);
nor UO_2131 (O_2131,N_19836,N_19632);
xor UO_2132 (O_2132,N_19820,N_19750);
and UO_2133 (O_2133,N_19772,N_19699);
nand UO_2134 (O_2134,N_19640,N_19740);
and UO_2135 (O_2135,N_19887,N_19942);
xnor UO_2136 (O_2136,N_19677,N_19802);
or UO_2137 (O_2137,N_19658,N_19783);
nand UO_2138 (O_2138,N_19923,N_19733);
nand UO_2139 (O_2139,N_19708,N_19730);
or UO_2140 (O_2140,N_19897,N_19725);
xnor UO_2141 (O_2141,N_19999,N_19637);
xor UO_2142 (O_2142,N_19852,N_19966);
nor UO_2143 (O_2143,N_19915,N_19703);
nand UO_2144 (O_2144,N_19917,N_19738);
nor UO_2145 (O_2145,N_19746,N_19929);
xor UO_2146 (O_2146,N_19744,N_19794);
nand UO_2147 (O_2147,N_19731,N_19699);
nor UO_2148 (O_2148,N_19906,N_19758);
nand UO_2149 (O_2149,N_19723,N_19645);
and UO_2150 (O_2150,N_19621,N_19637);
nor UO_2151 (O_2151,N_19856,N_19666);
or UO_2152 (O_2152,N_19681,N_19617);
or UO_2153 (O_2153,N_19952,N_19868);
nor UO_2154 (O_2154,N_19823,N_19769);
or UO_2155 (O_2155,N_19908,N_19664);
or UO_2156 (O_2156,N_19836,N_19811);
or UO_2157 (O_2157,N_19945,N_19823);
nand UO_2158 (O_2158,N_19615,N_19783);
nor UO_2159 (O_2159,N_19870,N_19798);
or UO_2160 (O_2160,N_19866,N_19643);
xnor UO_2161 (O_2161,N_19977,N_19609);
nand UO_2162 (O_2162,N_19897,N_19620);
xnor UO_2163 (O_2163,N_19941,N_19730);
nor UO_2164 (O_2164,N_19878,N_19621);
or UO_2165 (O_2165,N_19637,N_19940);
or UO_2166 (O_2166,N_19701,N_19694);
xor UO_2167 (O_2167,N_19704,N_19743);
or UO_2168 (O_2168,N_19609,N_19974);
nand UO_2169 (O_2169,N_19789,N_19736);
nand UO_2170 (O_2170,N_19840,N_19949);
nor UO_2171 (O_2171,N_19759,N_19996);
xnor UO_2172 (O_2172,N_19801,N_19799);
and UO_2173 (O_2173,N_19746,N_19965);
or UO_2174 (O_2174,N_19991,N_19805);
xor UO_2175 (O_2175,N_19674,N_19989);
nor UO_2176 (O_2176,N_19788,N_19944);
and UO_2177 (O_2177,N_19601,N_19728);
nor UO_2178 (O_2178,N_19919,N_19800);
nor UO_2179 (O_2179,N_19947,N_19853);
nand UO_2180 (O_2180,N_19915,N_19643);
or UO_2181 (O_2181,N_19993,N_19762);
nand UO_2182 (O_2182,N_19726,N_19879);
and UO_2183 (O_2183,N_19664,N_19606);
nor UO_2184 (O_2184,N_19980,N_19982);
nand UO_2185 (O_2185,N_19692,N_19602);
nand UO_2186 (O_2186,N_19872,N_19818);
xnor UO_2187 (O_2187,N_19720,N_19913);
nand UO_2188 (O_2188,N_19942,N_19619);
nand UO_2189 (O_2189,N_19901,N_19738);
or UO_2190 (O_2190,N_19615,N_19617);
xor UO_2191 (O_2191,N_19992,N_19895);
nor UO_2192 (O_2192,N_19912,N_19812);
and UO_2193 (O_2193,N_19714,N_19852);
xnor UO_2194 (O_2194,N_19724,N_19766);
nand UO_2195 (O_2195,N_19850,N_19887);
xnor UO_2196 (O_2196,N_19710,N_19623);
nand UO_2197 (O_2197,N_19751,N_19607);
nor UO_2198 (O_2198,N_19933,N_19628);
or UO_2199 (O_2199,N_19938,N_19698);
nor UO_2200 (O_2200,N_19654,N_19942);
nand UO_2201 (O_2201,N_19725,N_19857);
or UO_2202 (O_2202,N_19627,N_19756);
and UO_2203 (O_2203,N_19931,N_19621);
or UO_2204 (O_2204,N_19727,N_19652);
nand UO_2205 (O_2205,N_19695,N_19910);
nor UO_2206 (O_2206,N_19809,N_19733);
nand UO_2207 (O_2207,N_19763,N_19876);
nor UO_2208 (O_2208,N_19940,N_19877);
nand UO_2209 (O_2209,N_19777,N_19891);
nor UO_2210 (O_2210,N_19658,N_19938);
or UO_2211 (O_2211,N_19724,N_19904);
nor UO_2212 (O_2212,N_19675,N_19660);
nor UO_2213 (O_2213,N_19725,N_19965);
or UO_2214 (O_2214,N_19602,N_19922);
xor UO_2215 (O_2215,N_19662,N_19655);
xor UO_2216 (O_2216,N_19670,N_19746);
nand UO_2217 (O_2217,N_19878,N_19879);
nand UO_2218 (O_2218,N_19608,N_19718);
and UO_2219 (O_2219,N_19605,N_19929);
and UO_2220 (O_2220,N_19722,N_19774);
or UO_2221 (O_2221,N_19956,N_19768);
nand UO_2222 (O_2222,N_19851,N_19828);
nor UO_2223 (O_2223,N_19682,N_19865);
or UO_2224 (O_2224,N_19730,N_19669);
xnor UO_2225 (O_2225,N_19665,N_19754);
and UO_2226 (O_2226,N_19814,N_19904);
or UO_2227 (O_2227,N_19802,N_19813);
or UO_2228 (O_2228,N_19907,N_19797);
nand UO_2229 (O_2229,N_19630,N_19730);
and UO_2230 (O_2230,N_19820,N_19697);
nand UO_2231 (O_2231,N_19679,N_19860);
nor UO_2232 (O_2232,N_19850,N_19933);
xnor UO_2233 (O_2233,N_19791,N_19724);
nand UO_2234 (O_2234,N_19702,N_19862);
or UO_2235 (O_2235,N_19809,N_19827);
nand UO_2236 (O_2236,N_19856,N_19737);
and UO_2237 (O_2237,N_19774,N_19771);
nand UO_2238 (O_2238,N_19619,N_19905);
or UO_2239 (O_2239,N_19676,N_19669);
or UO_2240 (O_2240,N_19845,N_19821);
or UO_2241 (O_2241,N_19789,N_19875);
or UO_2242 (O_2242,N_19985,N_19615);
nand UO_2243 (O_2243,N_19911,N_19957);
and UO_2244 (O_2244,N_19723,N_19715);
xnor UO_2245 (O_2245,N_19948,N_19647);
nor UO_2246 (O_2246,N_19971,N_19903);
or UO_2247 (O_2247,N_19715,N_19631);
xor UO_2248 (O_2248,N_19620,N_19818);
or UO_2249 (O_2249,N_19852,N_19904);
or UO_2250 (O_2250,N_19645,N_19999);
or UO_2251 (O_2251,N_19679,N_19784);
xor UO_2252 (O_2252,N_19835,N_19993);
xor UO_2253 (O_2253,N_19930,N_19648);
nor UO_2254 (O_2254,N_19943,N_19670);
and UO_2255 (O_2255,N_19794,N_19755);
and UO_2256 (O_2256,N_19951,N_19772);
or UO_2257 (O_2257,N_19777,N_19692);
nor UO_2258 (O_2258,N_19916,N_19873);
nand UO_2259 (O_2259,N_19969,N_19690);
xor UO_2260 (O_2260,N_19718,N_19760);
xor UO_2261 (O_2261,N_19603,N_19936);
nand UO_2262 (O_2262,N_19667,N_19774);
xor UO_2263 (O_2263,N_19985,N_19983);
nand UO_2264 (O_2264,N_19703,N_19988);
xor UO_2265 (O_2265,N_19832,N_19935);
and UO_2266 (O_2266,N_19925,N_19850);
and UO_2267 (O_2267,N_19730,N_19694);
nor UO_2268 (O_2268,N_19703,N_19686);
nor UO_2269 (O_2269,N_19646,N_19794);
and UO_2270 (O_2270,N_19745,N_19779);
xor UO_2271 (O_2271,N_19836,N_19942);
xor UO_2272 (O_2272,N_19747,N_19826);
nor UO_2273 (O_2273,N_19819,N_19697);
and UO_2274 (O_2274,N_19848,N_19722);
xnor UO_2275 (O_2275,N_19786,N_19620);
or UO_2276 (O_2276,N_19987,N_19626);
nand UO_2277 (O_2277,N_19934,N_19840);
or UO_2278 (O_2278,N_19828,N_19655);
or UO_2279 (O_2279,N_19961,N_19689);
nor UO_2280 (O_2280,N_19933,N_19627);
and UO_2281 (O_2281,N_19969,N_19664);
or UO_2282 (O_2282,N_19651,N_19749);
and UO_2283 (O_2283,N_19677,N_19905);
and UO_2284 (O_2284,N_19935,N_19723);
or UO_2285 (O_2285,N_19826,N_19784);
or UO_2286 (O_2286,N_19884,N_19863);
and UO_2287 (O_2287,N_19882,N_19693);
xor UO_2288 (O_2288,N_19956,N_19730);
nand UO_2289 (O_2289,N_19929,N_19775);
and UO_2290 (O_2290,N_19713,N_19921);
or UO_2291 (O_2291,N_19761,N_19861);
or UO_2292 (O_2292,N_19904,N_19889);
or UO_2293 (O_2293,N_19842,N_19934);
or UO_2294 (O_2294,N_19903,N_19912);
nor UO_2295 (O_2295,N_19872,N_19948);
or UO_2296 (O_2296,N_19635,N_19960);
or UO_2297 (O_2297,N_19672,N_19751);
and UO_2298 (O_2298,N_19602,N_19682);
nor UO_2299 (O_2299,N_19703,N_19850);
or UO_2300 (O_2300,N_19721,N_19608);
nor UO_2301 (O_2301,N_19860,N_19686);
or UO_2302 (O_2302,N_19671,N_19913);
or UO_2303 (O_2303,N_19813,N_19940);
or UO_2304 (O_2304,N_19837,N_19952);
nand UO_2305 (O_2305,N_19958,N_19783);
nand UO_2306 (O_2306,N_19961,N_19845);
xnor UO_2307 (O_2307,N_19622,N_19919);
or UO_2308 (O_2308,N_19762,N_19624);
xnor UO_2309 (O_2309,N_19602,N_19929);
nand UO_2310 (O_2310,N_19809,N_19927);
and UO_2311 (O_2311,N_19969,N_19814);
nor UO_2312 (O_2312,N_19813,N_19630);
and UO_2313 (O_2313,N_19966,N_19767);
or UO_2314 (O_2314,N_19835,N_19871);
nor UO_2315 (O_2315,N_19626,N_19990);
nor UO_2316 (O_2316,N_19775,N_19631);
nor UO_2317 (O_2317,N_19606,N_19827);
nor UO_2318 (O_2318,N_19986,N_19824);
nand UO_2319 (O_2319,N_19623,N_19672);
or UO_2320 (O_2320,N_19675,N_19891);
or UO_2321 (O_2321,N_19895,N_19879);
and UO_2322 (O_2322,N_19717,N_19855);
xnor UO_2323 (O_2323,N_19600,N_19922);
and UO_2324 (O_2324,N_19819,N_19879);
nand UO_2325 (O_2325,N_19625,N_19919);
nand UO_2326 (O_2326,N_19608,N_19733);
or UO_2327 (O_2327,N_19678,N_19975);
nor UO_2328 (O_2328,N_19925,N_19993);
xor UO_2329 (O_2329,N_19772,N_19804);
or UO_2330 (O_2330,N_19752,N_19958);
nand UO_2331 (O_2331,N_19640,N_19869);
nor UO_2332 (O_2332,N_19834,N_19730);
or UO_2333 (O_2333,N_19762,N_19888);
and UO_2334 (O_2334,N_19780,N_19635);
nor UO_2335 (O_2335,N_19986,N_19956);
and UO_2336 (O_2336,N_19982,N_19899);
nand UO_2337 (O_2337,N_19866,N_19801);
or UO_2338 (O_2338,N_19781,N_19686);
or UO_2339 (O_2339,N_19634,N_19988);
or UO_2340 (O_2340,N_19776,N_19852);
nand UO_2341 (O_2341,N_19637,N_19855);
nand UO_2342 (O_2342,N_19859,N_19652);
nand UO_2343 (O_2343,N_19831,N_19928);
or UO_2344 (O_2344,N_19777,N_19649);
xnor UO_2345 (O_2345,N_19814,N_19975);
nand UO_2346 (O_2346,N_19940,N_19676);
xnor UO_2347 (O_2347,N_19878,N_19689);
nand UO_2348 (O_2348,N_19846,N_19615);
or UO_2349 (O_2349,N_19880,N_19858);
and UO_2350 (O_2350,N_19910,N_19640);
and UO_2351 (O_2351,N_19727,N_19825);
nand UO_2352 (O_2352,N_19876,N_19807);
xor UO_2353 (O_2353,N_19733,N_19671);
and UO_2354 (O_2354,N_19927,N_19862);
xor UO_2355 (O_2355,N_19905,N_19824);
nor UO_2356 (O_2356,N_19696,N_19834);
and UO_2357 (O_2357,N_19607,N_19902);
and UO_2358 (O_2358,N_19898,N_19615);
xor UO_2359 (O_2359,N_19994,N_19773);
xnor UO_2360 (O_2360,N_19764,N_19976);
nand UO_2361 (O_2361,N_19854,N_19622);
or UO_2362 (O_2362,N_19722,N_19831);
nor UO_2363 (O_2363,N_19896,N_19794);
nor UO_2364 (O_2364,N_19672,N_19731);
nand UO_2365 (O_2365,N_19830,N_19618);
nor UO_2366 (O_2366,N_19956,N_19965);
xnor UO_2367 (O_2367,N_19693,N_19833);
or UO_2368 (O_2368,N_19728,N_19835);
xnor UO_2369 (O_2369,N_19671,N_19697);
and UO_2370 (O_2370,N_19846,N_19808);
or UO_2371 (O_2371,N_19743,N_19840);
xor UO_2372 (O_2372,N_19698,N_19903);
xor UO_2373 (O_2373,N_19852,N_19647);
nand UO_2374 (O_2374,N_19930,N_19776);
xor UO_2375 (O_2375,N_19712,N_19821);
and UO_2376 (O_2376,N_19731,N_19680);
or UO_2377 (O_2377,N_19967,N_19654);
nand UO_2378 (O_2378,N_19853,N_19790);
and UO_2379 (O_2379,N_19958,N_19638);
xnor UO_2380 (O_2380,N_19842,N_19703);
and UO_2381 (O_2381,N_19939,N_19860);
nand UO_2382 (O_2382,N_19727,N_19739);
nor UO_2383 (O_2383,N_19994,N_19975);
nor UO_2384 (O_2384,N_19744,N_19857);
nor UO_2385 (O_2385,N_19999,N_19955);
and UO_2386 (O_2386,N_19900,N_19825);
nor UO_2387 (O_2387,N_19893,N_19805);
or UO_2388 (O_2388,N_19851,N_19644);
and UO_2389 (O_2389,N_19806,N_19966);
xor UO_2390 (O_2390,N_19914,N_19978);
or UO_2391 (O_2391,N_19999,N_19784);
nand UO_2392 (O_2392,N_19683,N_19864);
nor UO_2393 (O_2393,N_19970,N_19803);
or UO_2394 (O_2394,N_19723,N_19919);
nor UO_2395 (O_2395,N_19639,N_19916);
and UO_2396 (O_2396,N_19873,N_19739);
nor UO_2397 (O_2397,N_19877,N_19760);
nand UO_2398 (O_2398,N_19712,N_19860);
or UO_2399 (O_2399,N_19885,N_19706);
and UO_2400 (O_2400,N_19705,N_19816);
nand UO_2401 (O_2401,N_19859,N_19713);
xor UO_2402 (O_2402,N_19700,N_19661);
nor UO_2403 (O_2403,N_19704,N_19605);
or UO_2404 (O_2404,N_19677,N_19714);
xor UO_2405 (O_2405,N_19757,N_19839);
or UO_2406 (O_2406,N_19654,N_19680);
xnor UO_2407 (O_2407,N_19850,N_19650);
nand UO_2408 (O_2408,N_19606,N_19930);
and UO_2409 (O_2409,N_19780,N_19892);
xnor UO_2410 (O_2410,N_19744,N_19803);
and UO_2411 (O_2411,N_19986,N_19919);
nand UO_2412 (O_2412,N_19769,N_19826);
nor UO_2413 (O_2413,N_19990,N_19615);
or UO_2414 (O_2414,N_19842,N_19956);
xnor UO_2415 (O_2415,N_19955,N_19771);
nand UO_2416 (O_2416,N_19918,N_19900);
or UO_2417 (O_2417,N_19838,N_19622);
xor UO_2418 (O_2418,N_19657,N_19677);
xnor UO_2419 (O_2419,N_19693,N_19655);
and UO_2420 (O_2420,N_19668,N_19882);
nand UO_2421 (O_2421,N_19934,N_19657);
nand UO_2422 (O_2422,N_19945,N_19998);
or UO_2423 (O_2423,N_19939,N_19805);
nor UO_2424 (O_2424,N_19623,N_19907);
nor UO_2425 (O_2425,N_19615,N_19657);
nand UO_2426 (O_2426,N_19832,N_19903);
or UO_2427 (O_2427,N_19837,N_19853);
nand UO_2428 (O_2428,N_19781,N_19760);
and UO_2429 (O_2429,N_19751,N_19649);
nor UO_2430 (O_2430,N_19767,N_19796);
and UO_2431 (O_2431,N_19874,N_19602);
nor UO_2432 (O_2432,N_19687,N_19644);
nor UO_2433 (O_2433,N_19733,N_19963);
nand UO_2434 (O_2434,N_19792,N_19660);
or UO_2435 (O_2435,N_19663,N_19809);
or UO_2436 (O_2436,N_19979,N_19638);
and UO_2437 (O_2437,N_19627,N_19946);
and UO_2438 (O_2438,N_19935,N_19665);
nand UO_2439 (O_2439,N_19604,N_19639);
nor UO_2440 (O_2440,N_19876,N_19885);
and UO_2441 (O_2441,N_19716,N_19692);
and UO_2442 (O_2442,N_19676,N_19937);
xnor UO_2443 (O_2443,N_19838,N_19776);
nand UO_2444 (O_2444,N_19728,N_19798);
nand UO_2445 (O_2445,N_19641,N_19971);
or UO_2446 (O_2446,N_19810,N_19754);
and UO_2447 (O_2447,N_19665,N_19693);
xor UO_2448 (O_2448,N_19773,N_19700);
nand UO_2449 (O_2449,N_19932,N_19684);
xor UO_2450 (O_2450,N_19865,N_19997);
xnor UO_2451 (O_2451,N_19673,N_19629);
nand UO_2452 (O_2452,N_19879,N_19692);
and UO_2453 (O_2453,N_19693,N_19754);
nor UO_2454 (O_2454,N_19797,N_19744);
and UO_2455 (O_2455,N_19733,N_19900);
nor UO_2456 (O_2456,N_19627,N_19819);
xnor UO_2457 (O_2457,N_19894,N_19972);
nor UO_2458 (O_2458,N_19967,N_19891);
and UO_2459 (O_2459,N_19972,N_19725);
nor UO_2460 (O_2460,N_19776,N_19710);
or UO_2461 (O_2461,N_19819,N_19639);
nor UO_2462 (O_2462,N_19704,N_19654);
xnor UO_2463 (O_2463,N_19698,N_19633);
xnor UO_2464 (O_2464,N_19605,N_19867);
and UO_2465 (O_2465,N_19767,N_19737);
and UO_2466 (O_2466,N_19613,N_19871);
nor UO_2467 (O_2467,N_19681,N_19786);
and UO_2468 (O_2468,N_19826,N_19653);
nor UO_2469 (O_2469,N_19730,N_19933);
and UO_2470 (O_2470,N_19895,N_19788);
nand UO_2471 (O_2471,N_19882,N_19907);
nor UO_2472 (O_2472,N_19855,N_19719);
nand UO_2473 (O_2473,N_19951,N_19946);
xor UO_2474 (O_2474,N_19679,N_19928);
nand UO_2475 (O_2475,N_19646,N_19906);
nand UO_2476 (O_2476,N_19816,N_19764);
nor UO_2477 (O_2477,N_19677,N_19748);
and UO_2478 (O_2478,N_19989,N_19909);
nor UO_2479 (O_2479,N_19992,N_19759);
nor UO_2480 (O_2480,N_19654,N_19726);
or UO_2481 (O_2481,N_19918,N_19711);
nor UO_2482 (O_2482,N_19652,N_19712);
nor UO_2483 (O_2483,N_19902,N_19892);
nand UO_2484 (O_2484,N_19628,N_19873);
and UO_2485 (O_2485,N_19988,N_19779);
xor UO_2486 (O_2486,N_19831,N_19887);
nand UO_2487 (O_2487,N_19809,N_19855);
nand UO_2488 (O_2488,N_19842,N_19810);
and UO_2489 (O_2489,N_19831,N_19629);
xnor UO_2490 (O_2490,N_19980,N_19860);
or UO_2491 (O_2491,N_19717,N_19961);
xnor UO_2492 (O_2492,N_19911,N_19860);
nand UO_2493 (O_2493,N_19865,N_19950);
xnor UO_2494 (O_2494,N_19688,N_19871);
xor UO_2495 (O_2495,N_19913,N_19790);
and UO_2496 (O_2496,N_19924,N_19670);
nand UO_2497 (O_2497,N_19613,N_19714);
or UO_2498 (O_2498,N_19745,N_19691);
xnor UO_2499 (O_2499,N_19627,N_19776);
endmodule