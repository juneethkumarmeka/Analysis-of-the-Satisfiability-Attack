module basic_2000_20000_2500_4_levels_5xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
or U0 (N_0,In_7,In_610);
nand U1 (N_1,In_1797,In_720);
nand U2 (N_2,In_103,In_135);
nand U3 (N_3,In_312,In_105);
nand U4 (N_4,In_1664,In_0);
and U5 (N_5,In_1551,In_1945);
nor U6 (N_6,In_1331,In_1299);
nor U7 (N_7,In_572,In_1944);
and U8 (N_8,In_1187,In_506);
and U9 (N_9,In_955,In_1203);
and U10 (N_10,In_447,In_1248);
nand U11 (N_11,In_782,In_1963);
and U12 (N_12,In_1296,In_232);
or U13 (N_13,In_1633,In_937);
and U14 (N_14,In_1029,In_939);
nor U15 (N_15,In_1795,In_405);
nand U16 (N_16,In_1863,In_695);
nor U17 (N_17,In_1267,In_79);
xnor U18 (N_18,In_1210,In_1337);
and U19 (N_19,In_1524,In_1098);
xnor U20 (N_20,In_1052,In_1993);
nor U21 (N_21,In_1458,In_846);
xor U22 (N_22,In_1449,In_1670);
and U23 (N_23,In_1720,In_806);
and U24 (N_24,In_1542,In_1058);
nor U25 (N_25,In_1149,In_1427);
nor U26 (N_26,In_755,In_1594);
and U27 (N_27,In_869,In_1107);
and U28 (N_28,In_1539,In_1439);
nor U29 (N_29,In_1703,In_1752);
or U30 (N_30,In_1915,In_345);
nand U31 (N_31,In_333,In_169);
nand U32 (N_32,In_314,In_228);
nand U33 (N_33,In_1657,In_1529);
xor U34 (N_34,In_1272,In_1475);
or U35 (N_35,In_663,In_1214);
or U36 (N_36,In_822,In_157);
or U37 (N_37,In_430,In_1634);
nand U38 (N_38,In_1489,In_1096);
nor U39 (N_39,In_868,In_863);
and U40 (N_40,In_1918,In_1216);
nand U41 (N_41,In_183,In_236);
xnor U42 (N_42,In_424,In_133);
nand U43 (N_43,In_366,In_1414);
and U44 (N_44,In_1951,In_1852);
nand U45 (N_45,In_1297,In_1485);
nor U46 (N_46,In_1603,In_1157);
nand U47 (N_47,In_1717,In_1048);
nand U48 (N_48,In_554,In_1082);
nor U49 (N_49,In_1511,In_1364);
or U50 (N_50,In_1249,In_1958);
nand U51 (N_51,In_1579,In_973);
nor U52 (N_52,In_828,In_1238);
nand U53 (N_53,In_1431,In_473);
nand U54 (N_54,In_947,In_684);
nand U55 (N_55,In_91,In_1229);
nand U56 (N_56,In_1146,In_248);
nor U57 (N_57,In_987,In_1114);
xor U58 (N_58,In_1936,In_1142);
or U59 (N_59,In_843,In_1365);
nand U60 (N_60,In_1665,In_1691);
nand U61 (N_61,In_485,In_1373);
or U62 (N_62,In_368,In_349);
nand U63 (N_63,In_1195,In_1921);
nand U64 (N_64,In_518,In_1970);
xnor U65 (N_65,In_53,In_390);
nand U66 (N_66,In_1332,In_998);
nor U67 (N_67,In_1042,In_1600);
nand U68 (N_68,In_34,In_626);
or U69 (N_69,In_989,In_700);
and U70 (N_70,In_871,In_662);
nand U71 (N_71,In_24,In_204);
nand U72 (N_72,In_1979,In_1748);
nand U73 (N_73,In_476,In_1252);
nand U74 (N_74,In_1695,In_1499);
nand U75 (N_75,In_1931,In_29);
nor U76 (N_76,In_218,In_1080);
and U77 (N_77,In_1192,In_1736);
and U78 (N_78,In_468,In_678);
and U79 (N_79,In_780,In_522);
nand U80 (N_80,In_654,In_1467);
nor U81 (N_81,In_928,In_694);
nor U82 (N_82,In_1160,In_605);
or U83 (N_83,In_840,In_798);
or U84 (N_84,In_205,In_1152);
or U85 (N_85,In_922,In_600);
nand U86 (N_86,In_643,In_1682);
or U87 (N_87,In_1770,In_1581);
nor U88 (N_88,In_294,In_1882);
or U89 (N_89,In_1158,In_951);
or U90 (N_90,In_211,In_1739);
nor U91 (N_91,In_1153,In_233);
and U92 (N_92,In_28,In_1487);
nor U93 (N_93,In_1630,In_1334);
xor U94 (N_94,In_593,In_1780);
and U95 (N_95,In_494,In_1803);
nand U96 (N_96,In_1286,In_1159);
nand U97 (N_97,In_882,In_83);
xor U98 (N_98,In_503,In_1909);
nand U99 (N_99,In_1023,In_725);
or U100 (N_100,In_817,In_1068);
nand U101 (N_101,In_172,In_875);
or U102 (N_102,In_1009,In_1729);
or U103 (N_103,In_1019,In_1517);
nor U104 (N_104,In_1340,In_724);
nand U105 (N_105,In_773,In_758);
nand U106 (N_106,In_265,In_216);
xor U107 (N_107,In_1399,In_243);
nor U108 (N_108,In_1593,In_1627);
or U109 (N_109,In_1441,In_1652);
or U110 (N_110,In_1523,In_1094);
nand U111 (N_111,In_877,In_693);
or U112 (N_112,In_1874,In_1805);
nor U113 (N_113,In_344,In_1710);
and U114 (N_114,In_1011,In_845);
nand U115 (N_115,In_1826,In_1434);
and U116 (N_116,In_1790,In_364);
and U117 (N_117,In_633,In_1424);
nand U118 (N_118,In_1911,In_1775);
and U119 (N_119,In_400,In_270);
nand U120 (N_120,In_1067,In_889);
nor U121 (N_121,In_1314,In_722);
nand U122 (N_122,In_1277,In_661);
nor U123 (N_123,In_1783,In_534);
nor U124 (N_124,In_909,In_866);
or U125 (N_125,In_1577,In_1135);
or U126 (N_126,In_1723,In_33);
nand U127 (N_127,In_844,In_331);
and U128 (N_128,In_713,In_1137);
or U129 (N_129,In_166,In_635);
nand U130 (N_130,In_730,In_335);
or U131 (N_131,In_792,In_523);
and U132 (N_132,In_1686,In_1347);
nand U133 (N_133,In_799,In_1794);
nor U134 (N_134,In_1541,In_1947);
and U135 (N_135,In_898,In_1389);
and U136 (N_136,In_379,In_1933);
nor U137 (N_137,In_1089,In_543);
nand U138 (N_138,In_1092,In_342);
nor U139 (N_139,In_1133,In_716);
or U140 (N_140,In_1645,In_1193);
nand U141 (N_141,In_824,In_289);
nor U142 (N_142,In_652,In_850);
nor U143 (N_143,In_1117,In_1779);
nor U144 (N_144,In_1932,In_1896);
nor U145 (N_145,In_36,In_1335);
or U146 (N_146,In_1853,In_326);
or U147 (N_147,In_224,In_1430);
and U148 (N_148,In_41,In_1900);
and U149 (N_149,In_329,In_252);
and U150 (N_150,In_639,In_1995);
nor U151 (N_151,In_1490,In_1377);
nand U152 (N_152,In_1698,In_1569);
nand U153 (N_153,In_1156,In_818);
nor U154 (N_154,In_1948,In_50);
nor U155 (N_155,In_1077,In_328);
and U156 (N_156,In_1255,In_659);
nor U157 (N_157,In_90,In_1385);
xnor U158 (N_158,In_1410,In_411);
and U159 (N_159,In_1671,In_549);
or U160 (N_160,In_321,In_147);
nand U161 (N_161,In_303,In_574);
or U162 (N_162,In_1582,In_1576);
and U163 (N_163,In_1323,In_1452);
and U164 (N_164,In_1525,In_3);
nand U165 (N_165,In_1804,In_247);
nand U166 (N_166,In_981,In_687);
nand U167 (N_167,In_1530,In_805);
xnor U168 (N_168,In_1837,In_1103);
nor U169 (N_169,In_1497,In_665);
nor U170 (N_170,In_201,In_681);
and U171 (N_171,In_1744,In_1250);
nand U172 (N_172,In_1880,In_1268);
and U173 (N_173,In_897,In_539);
nor U174 (N_174,In_222,In_508);
and U175 (N_175,In_1714,In_703);
nor U176 (N_176,In_1336,In_1139);
xor U177 (N_177,In_1599,In_1387);
nand U178 (N_178,In_1303,In_747);
nand U179 (N_179,In_1221,In_1181);
or U180 (N_180,In_640,In_1433);
nand U181 (N_181,In_346,In_1798);
and U182 (N_182,In_313,In_1);
nor U183 (N_183,In_207,In_848);
and U184 (N_184,In_491,In_182);
and U185 (N_185,In_1394,In_1680);
or U186 (N_186,In_590,In_1819);
nand U187 (N_187,In_766,In_258);
or U188 (N_188,In_1182,In_997);
nand U189 (N_189,In_786,In_1169);
or U190 (N_190,In_1086,In_778);
nor U191 (N_191,In_1763,In_1832);
or U192 (N_192,In_466,In_1376);
or U193 (N_193,In_448,In_790);
and U194 (N_194,In_477,In_1887);
nand U195 (N_195,In_203,In_884);
xor U196 (N_196,In_1526,In_1959);
nand U197 (N_197,In_1428,In_1064);
and U198 (N_198,In_402,In_414);
or U199 (N_199,In_569,In_791);
or U200 (N_200,In_1788,In_489);
or U201 (N_201,In_1285,In_1980);
xnor U202 (N_202,In_95,In_988);
nor U203 (N_203,In_919,In_407);
nor U204 (N_204,In_1417,In_1626);
and U205 (N_205,In_1493,In_337);
nor U206 (N_206,In_1534,In_1402);
nand U207 (N_207,In_1728,In_1586);
and U208 (N_208,In_16,In_1006);
nand U209 (N_209,In_647,In_1864);
or U210 (N_210,In_1623,In_691);
nand U211 (N_211,In_1491,In_679);
nor U212 (N_212,In_1359,In_999);
or U213 (N_213,In_154,In_1173);
or U214 (N_214,In_497,In_1590);
nand U215 (N_215,In_956,In_1785);
and U216 (N_216,In_308,In_1031);
nand U217 (N_217,In_1099,In_1999);
xnor U218 (N_218,In_271,In_1850);
nor U219 (N_219,In_1369,In_2);
or U220 (N_220,In_1507,In_556);
or U221 (N_221,In_890,In_580);
xor U222 (N_222,In_936,In_385);
nor U223 (N_223,In_195,In_958);
and U224 (N_224,In_1217,In_606);
nand U225 (N_225,In_1053,In_1243);
and U226 (N_226,In_474,In_212);
or U227 (N_227,In_1287,In_1609);
nor U228 (N_228,In_1848,In_1946);
nor U229 (N_229,In_1097,In_517);
and U230 (N_230,In_913,In_1190);
or U231 (N_231,In_860,In_1740);
or U232 (N_232,In_710,In_343);
or U233 (N_233,In_1806,In_607);
or U234 (N_234,In_904,In_1465);
or U235 (N_235,In_1624,In_980);
or U236 (N_236,In_878,In_1245);
or U237 (N_237,In_594,In_754);
and U238 (N_238,In_601,In_1119);
nand U239 (N_239,In_586,In_944);
and U240 (N_240,In_383,In_749);
nand U241 (N_241,In_1844,In_119);
nand U242 (N_242,In_1401,In_1547);
nor U243 (N_243,In_1591,In_1888);
nor U244 (N_244,In_370,In_1422);
or U245 (N_245,In_327,In_624);
and U246 (N_246,In_1201,In_759);
or U247 (N_247,In_1145,In_300);
nor U248 (N_248,In_393,In_1513);
and U249 (N_249,In_1165,In_736);
or U250 (N_250,In_1075,In_530);
and U251 (N_251,In_1321,In_969);
nor U252 (N_252,In_1765,In_961);
nor U253 (N_253,In_492,In_1261);
or U254 (N_254,In_571,In_301);
nand U255 (N_255,In_391,In_853);
nor U256 (N_256,In_1988,In_1189);
nand U257 (N_257,In_475,In_266);
nand U258 (N_258,In_1984,In_1057);
and U259 (N_259,In_1294,In_1715);
or U260 (N_260,In_1502,In_1903);
or U261 (N_261,In_283,In_1606);
xnor U262 (N_262,In_1416,In_916);
xor U263 (N_263,In_168,In_481);
or U264 (N_264,In_618,In_1725);
or U265 (N_265,In_42,In_1776);
nand U266 (N_266,In_1757,In_1202);
or U267 (N_267,In_309,In_398);
nor U268 (N_268,In_394,In_323);
and U269 (N_269,In_120,In_1104);
and U270 (N_270,In_583,In_1601);
nand U271 (N_271,In_1110,In_1350);
nand U272 (N_272,In_657,In_551);
nor U273 (N_273,In_765,In_1611);
nand U274 (N_274,In_102,In_597);
xnor U275 (N_275,In_1934,In_1998);
nor U276 (N_276,In_908,In_175);
and U277 (N_277,In_1025,In_1212);
nor U278 (N_278,In_1649,In_1178);
nand U279 (N_279,In_1544,In_471);
and U280 (N_280,In_748,In_1981);
nand U281 (N_281,In_1817,In_1102);
nor U282 (N_282,In_836,In_1111);
and U283 (N_283,In_1460,In_1127);
nand U284 (N_284,In_462,In_381);
or U285 (N_285,In_1629,In_1200);
nand U286 (N_286,In_1301,In_1300);
nand U287 (N_287,In_563,In_1307);
and U288 (N_288,In_267,In_535);
nand U289 (N_289,In_263,In_762);
and U290 (N_290,In_945,In_184);
or U291 (N_291,In_727,In_1901);
or U292 (N_292,In_1847,In_764);
and U293 (N_293,In_1587,In_1274);
nand U294 (N_294,In_1688,In_927);
and U295 (N_295,In_1237,In_1105);
xor U296 (N_296,In_311,In_953);
nor U297 (N_297,In_795,In_1760);
xor U298 (N_298,In_1907,In_1204);
nand U299 (N_299,In_753,In_1134);
or U300 (N_300,In_1069,In_1386);
nor U301 (N_301,In_99,In_905);
or U302 (N_302,In_1758,In_1010);
or U303 (N_303,In_1841,In_1043);
nand U304 (N_304,In_963,In_1235);
nor U305 (N_305,In_1503,In_1846);
nand U306 (N_306,In_1508,In_810);
or U307 (N_307,In_131,In_1681);
xnor U308 (N_308,In_1696,In_1141);
nand U309 (N_309,In_596,In_540);
and U310 (N_310,In_60,In_1793);
nor U311 (N_311,In_584,In_316);
and U312 (N_312,In_912,In_67);
nor U313 (N_313,In_1592,In_376);
or U314 (N_314,In_1028,In_153);
nor U315 (N_315,In_1398,In_1176);
nor U316 (N_316,In_1230,In_531);
or U317 (N_317,In_128,In_144);
and U318 (N_318,In_1573,In_1138);
and U319 (N_319,In_515,In_97);
nand U320 (N_320,In_996,In_670);
or U321 (N_321,In_63,In_340);
nand U322 (N_322,In_544,In_1749);
and U323 (N_323,In_1322,In_1381);
or U324 (N_324,In_92,In_1413);
nand U325 (N_325,In_1438,In_1085);
nor U326 (N_326,In_933,In_1676);
nor U327 (N_327,In_482,In_784);
nand U328 (N_328,In_1044,In_885);
or U329 (N_329,In_1355,In_1244);
or U330 (N_330,In_202,In_1213);
or U331 (N_331,In_1168,In_1483);
and U332 (N_332,In_1186,In_1435);
nor U333 (N_333,In_957,In_1083);
nand U334 (N_334,In_1128,In_75);
xnor U335 (N_335,In_76,In_432);
and U336 (N_336,In_1769,In_838);
and U337 (N_337,In_1310,In_760);
and U338 (N_338,In_1356,In_136);
nand U339 (N_339,In_851,In_1494);
or U340 (N_340,In_121,In_1822);
or U341 (N_341,In_1421,In_1861);
nand U342 (N_342,In_221,In_1997);
and U343 (N_343,In_1727,In_1589);
and U344 (N_344,In_1730,In_306);
and U345 (N_345,In_977,In_598);
and U346 (N_346,In_1650,In_1761);
or U347 (N_347,In_220,In_1578);
nor U348 (N_348,In_1488,In_1000);
xor U349 (N_349,In_739,In_1554);
and U350 (N_350,In_1563,In_1001);
and U351 (N_351,In_1407,In_1264);
and U352 (N_352,In_254,In_1408);
nor U353 (N_353,In_1718,In_752);
nor U354 (N_354,In_718,In_921);
nor U355 (N_355,In_1070,In_134);
nor U356 (N_356,In_1823,In_516);
nor U357 (N_357,In_1572,In_588);
xnor U358 (N_358,In_1943,In_815);
nor U359 (N_359,In_547,In_512);
nand U360 (N_360,In_1219,In_733);
nor U361 (N_361,In_1046,In_1692);
nor U362 (N_362,In_209,In_1093);
xnor U363 (N_363,In_113,In_71);
or U364 (N_364,In_353,In_1442);
and U365 (N_365,In_111,In_1669);
nor U366 (N_366,In_4,In_525);
nand U367 (N_367,In_809,In_1226);
xor U368 (N_368,In_1171,In_1802);
nand U369 (N_369,In_690,In_406);
nand U370 (N_370,In_613,In_743);
and U371 (N_371,In_1037,In_1050);
and U372 (N_372,In_188,In_1256);
and U373 (N_373,In_1234,In_219);
nand U374 (N_374,In_1942,In_100);
or U375 (N_375,In_826,In_533);
nand U376 (N_376,In_1353,In_416);
nand U377 (N_377,In_161,In_288);
nand U378 (N_378,In_979,In_49);
nor U379 (N_379,In_1527,In_861);
and U380 (N_380,In_1824,In_578);
or U381 (N_381,In_650,In_896);
and U382 (N_382,In_1866,In_1531);
nor U383 (N_383,In_1916,In_1521);
or U384 (N_384,In_284,In_1786);
and U385 (N_385,In_1782,In_1899);
and U386 (N_386,In_185,In_1668);
and U387 (N_387,In_1778,In_1810);
or U388 (N_388,In_1342,In_1625);
nand U389 (N_389,In_638,In_852);
nor U390 (N_390,In_318,In_1891);
or U391 (N_391,In_847,In_1196);
nor U392 (N_392,In_15,In_1233);
nor U393 (N_393,In_110,In_952);
nand U394 (N_394,In_1357,In_1172);
and U395 (N_395,In_305,In_1764);
nor U396 (N_396,In_1505,In_1170);
nor U397 (N_397,In_298,In_1358);
nor U398 (N_398,In_1370,In_341);
or U399 (N_399,In_373,In_438);
nand U400 (N_400,In_58,In_880);
and U401 (N_401,In_559,In_1716);
and U402 (N_402,In_472,In_1033);
or U403 (N_403,In_1838,In_245);
and U404 (N_404,In_622,In_627);
nand U405 (N_405,In_382,In_612);
or U406 (N_406,In_872,In_32);
nor U407 (N_407,In_445,In_903);
nor U408 (N_408,In_565,In_213);
or U409 (N_409,In_1878,In_1304);
or U410 (N_410,In_1712,In_23);
or U411 (N_411,In_357,In_292);
or U412 (N_412,In_1602,In_932);
nor U413 (N_413,In_257,In_1393);
and U414 (N_414,In_830,In_1054);
or U415 (N_415,In_8,In_277);
nand U416 (N_416,In_1528,In_275);
nand U417 (N_417,In_1024,In_1273);
or U418 (N_418,In_415,In_857);
nand U419 (N_419,In_116,In_1996);
or U420 (N_420,In_1078,In_1247);
nand U421 (N_421,In_708,In_967);
or U422 (N_422,In_1236,In_974);
xor U423 (N_423,In_47,In_486);
nand U424 (N_424,In_787,In_1124);
nor U425 (N_425,In_668,In_637);
and U426 (N_426,In_737,In_1132);
nor U427 (N_427,In_550,In_46);
nand U428 (N_428,In_1598,In_1150);
or U429 (N_429,In_1500,In_568);
and U430 (N_430,In_1095,In_673);
or U431 (N_431,In_1440,In_1191);
nand U432 (N_432,In_307,In_1584);
nand U433 (N_433,In_602,In_279);
nand U434 (N_434,In_1515,In_1477);
xor U435 (N_435,In_1608,In_719);
nand U436 (N_436,In_17,In_274);
or U437 (N_437,In_812,In_813);
nor U438 (N_438,In_1913,In_1320);
nand U439 (N_439,In_85,In_22);
xor U440 (N_440,In_196,In_163);
nor U441 (N_441,In_167,In_966);
nor U442 (N_442,In_575,In_591);
nand U443 (N_443,In_1045,In_1518);
nand U444 (N_444,In_1924,In_911);
or U445 (N_445,In_1374,In_801);
and U446 (N_446,In_867,In_802);
xor U447 (N_447,In_1890,In_841);
nor U448 (N_448,In_1978,In_104);
nand U449 (N_449,In_1557,In_1756);
and U450 (N_450,In_1546,In_285);
and U451 (N_451,In_500,In_1305);
nand U452 (N_452,In_976,In_545);
nor U453 (N_453,In_1858,In_165);
nor U454 (N_454,In_126,In_608);
nor U455 (N_455,In_1856,In_1767);
or U456 (N_456,In_1612,In_595);
and U457 (N_457,In_66,In_1506);
and U458 (N_458,In_803,In_1354);
or U459 (N_459,In_874,In_141);
nand U460 (N_460,In_237,In_1282);
nand U461 (N_461,In_1558,In_269);
xor U462 (N_462,In_155,In_653);
nand U463 (N_463,In_645,In_56);
xnor U464 (N_464,In_109,In_1595);
or U465 (N_465,In_660,In_1893);
and U466 (N_466,In_240,In_125);
xor U467 (N_467,In_1444,In_352);
xnor U468 (N_468,In_1813,In_1144);
or U469 (N_469,In_320,In_1112);
nand U470 (N_470,In_338,In_1708);
or U471 (N_471,In_1166,In_457);
nor U472 (N_472,In_1862,In_94);
xnor U473 (N_473,In_317,In_1621);
or U474 (N_474,In_62,In_621);
nand U475 (N_475,In_171,In_404);
nand U476 (N_476,In_210,In_907);
or U477 (N_477,In_672,In_498);
nor U478 (N_478,In_360,In_194);
nor U479 (N_479,In_1619,In_454);
nor U480 (N_480,In_1298,In_1352);
nor U481 (N_481,In_895,In_567);
and U482 (N_482,In_734,In_949);
xor U483 (N_483,In_774,In_355);
and U484 (N_484,In_1454,In_1063);
or U485 (N_485,In_1583,In_1648);
and U486 (N_486,In_1990,In_137);
nand U487 (N_487,In_1704,In_1091);
nand U488 (N_488,In_513,In_1205);
and U489 (N_489,In_1768,In_865);
nor U490 (N_490,In_671,In_1656);
and U491 (N_491,In_1291,In_985);
nor U492 (N_492,In_1361,In_483);
xnor U493 (N_493,In_1257,In_37);
or U494 (N_494,In_1071,In_127);
and U495 (N_495,In_1957,In_1251);
or U496 (N_496,In_656,In_881);
nor U497 (N_497,In_160,In_582);
or U498 (N_498,In_1923,In_1701);
and U499 (N_499,In_634,In_297);
or U500 (N_500,In_887,In_1533);
and U501 (N_501,In_655,In_1411);
or U502 (N_502,In_504,In_1362);
or U503 (N_503,In_408,In_763);
and U504 (N_504,In_1777,In_469);
xnor U505 (N_505,In_452,In_1163);
xor U506 (N_506,In_467,In_1318);
nand U507 (N_507,In_101,In_420);
nor U508 (N_508,In_1269,In_1655);
or U509 (N_509,In_145,In_1418);
xor U510 (N_510,In_1700,In_399);
nor U511 (N_511,In_1821,In_1426);
and U512 (N_512,In_499,In_625);
or U513 (N_513,In_244,In_1724);
nand U514 (N_514,In_1129,In_1892);
or U515 (N_515,In_1759,In_1496);
or U516 (N_516,In_1991,In_453);
and U517 (N_517,In_893,In_706);
and U518 (N_518,In_440,In_1906);
nor U519 (N_519,In_142,In_1384);
xor U520 (N_520,In_130,In_1131);
or U521 (N_521,In_1726,In_666);
nor U522 (N_522,In_64,In_1486);
nor U523 (N_523,In_1266,In_72);
or U524 (N_524,In_1719,In_1894);
nor U525 (N_525,In_883,In_1967);
nor U526 (N_526,In_1754,In_350);
nor U527 (N_527,In_45,In_732);
and U528 (N_528,In_1658,In_946);
nor U529 (N_529,In_1451,In_253);
xor U530 (N_530,In_528,In_675);
or U531 (N_531,In_555,In_1161);
nor U532 (N_532,In_422,In_1315);
and U533 (N_533,In_804,In_821);
nor U534 (N_534,In_686,In_359);
nand U535 (N_535,In_1631,In_837);
or U536 (N_536,In_367,In_1504);
and U537 (N_537,In_1855,In_975);
xor U538 (N_538,In_1185,In_570);
or U539 (N_539,In_831,In_39);
or U540 (N_540,In_234,In_1538);
xnor U541 (N_541,In_1140,In_771);
xnor U542 (N_542,In_1935,In_1868);
nor U543 (N_543,In_403,In_1781);
and U544 (N_544,In_1062,In_378);
nor U545 (N_545,In_1455,In_1972);
xnor U546 (N_546,In_480,In_1910);
nand U547 (N_547,In_1960,In_994);
nor U548 (N_548,In_524,In_1860);
nor U549 (N_549,In_1148,In_1406);
nand U550 (N_550,In_1620,In_1327);
and U551 (N_551,In_1641,In_938);
or U552 (N_552,In_1550,In_1755);
and U553 (N_553,In_1869,In_1747);
or U554 (N_554,In_1179,In_940);
nand U555 (N_555,In_1879,In_789);
or U556 (N_556,In_970,In_1812);
nor U557 (N_557,In_699,In_1450);
or U558 (N_558,In_375,In_395);
nor U559 (N_559,In_984,In_934);
nand U560 (N_560,In_456,In_1745);
and U561 (N_561,In_849,In_1733);
nand U562 (N_562,In_1690,In_461);
or U563 (N_563,In_579,In_1188);
nand U564 (N_564,In_636,In_1877);
nor U565 (N_565,In_332,In_823);
nor U566 (N_566,In_1125,In_410);
nor U567 (N_567,In_1930,In_1480);
nand U568 (N_568,In_1459,In_1328);
or U569 (N_569,In_351,In_1344);
nor U570 (N_570,In_1800,In_943);
nand U571 (N_571,In_1588,In_44);
nor U572 (N_572,In_705,In_1827);
and U573 (N_573,In_1929,In_1808);
nand U574 (N_574,In_238,In_1231);
xor U575 (N_575,In_761,In_1985);
nand U576 (N_576,In_1897,In_1343);
xor U577 (N_577,In_1270,In_1883);
and U578 (N_578,In_1457,In_619);
nand U579 (N_579,In_1616,In_777);
nand U580 (N_580,In_775,In_738);
or U581 (N_581,In_421,In_1478);
nor U582 (N_582,In_800,In_900);
nor U583 (N_583,In_1040,In_241);
and U584 (N_584,In_948,In_250);
or U585 (N_585,In_510,In_460);
or U586 (N_586,In_781,In_1618);
or U587 (N_587,In_746,In_1476);
nand U588 (N_588,In_1628,In_1865);
or U589 (N_589,In_698,In_1632);
or U590 (N_590,In_149,In_413);
and U591 (N_591,In_1743,In_1519);
nor U592 (N_592,In_1927,In_891);
or U593 (N_593,In_680,In_1642);
nand U594 (N_594,In_669,In_418);
nor U595 (N_595,In_1351,In_272);
nor U596 (N_596,In_1084,In_1319);
or U597 (N_597,In_918,In_1973);
nor U598 (N_598,In_971,In_1106);
nor U599 (N_599,In_1482,In_449);
nand U600 (N_600,In_978,In_1122);
xor U601 (N_601,In_1568,In_1481);
or U602 (N_602,In_519,In_129);
nand U603 (N_603,In_917,In_1312);
nand U604 (N_604,In_1076,In_1809);
and U605 (N_605,In_1843,In_1225);
nand U606 (N_606,In_1060,In_1675);
or U607 (N_607,In_1663,In_520);
nor U608 (N_608,In_59,In_862);
nand U609 (N_609,In_1820,In_757);
or U610 (N_610,In_688,In_490);
nor U611 (N_611,In_426,In_1056);
nand U612 (N_612,In_1938,In_1939);
xor U613 (N_613,In_1017,In_114);
nor U614 (N_614,In_702,In_365);
or U615 (N_615,In_1390,In_450);
nor U616 (N_616,In_158,In_162);
nor U617 (N_617,In_1789,In_1382);
xnor U618 (N_618,In_181,In_599);
nor U619 (N_619,In_721,In_1072);
nor U620 (N_620,In_1325,In_443);
nor U621 (N_621,In_1198,In_682);
or U622 (N_622,In_463,In_88);
nor U623 (N_623,In_57,In_1771);
nand U624 (N_624,In_538,In_926);
nor U625 (N_625,In_286,In_177);
or U626 (N_626,In_1516,In_742);
nor U627 (N_627,In_1952,In_1854);
xnor U628 (N_628,In_1693,In_1220);
nand U629 (N_629,In_152,In_729);
nand U630 (N_630,In_1065,In_1015);
nor U631 (N_631,In_1640,In_278);
or U632 (N_632,In_180,In_442);
or U633 (N_633,In_138,In_61);
xnor U634 (N_634,In_386,In_735);
nand U635 (N_635,In_514,In_18);
nor U636 (N_636,In_630,In_696);
and U637 (N_637,In_87,In_290);
nand U638 (N_638,In_1443,In_1654);
nor U639 (N_639,In_794,In_676);
nor U640 (N_640,In_914,In_683);
xor U641 (N_641,In_1562,In_1409);
nor U642 (N_642,In_797,In_1290);
or U643 (N_643,In_1684,In_1262);
nor U644 (N_644,In_139,In_74);
nand U645 (N_645,In_1047,In_1971);
or U646 (N_646,In_1143,In_1278);
and U647 (N_647,In_1734,In_1283);
or U648 (N_648,In_14,In_291);
and U649 (N_649,In_1961,In_935);
or U650 (N_650,In_1976,In_1073);
or U651 (N_651,In_1051,In_1026);
xnor U652 (N_652,In_1647,In_832);
nor U653 (N_653,In_1466,In_1575);
and U654 (N_654,In_964,In_1762);
and U655 (N_655,In_1925,In_479);
or U656 (N_656,In_1532,In_1520);
nand U657 (N_657,In_509,In_942);
and U658 (N_658,In_13,In_1711);
and U659 (N_659,In_1081,In_560);
and U660 (N_660,In_282,In_86);
or U661 (N_661,In_950,In_1501);
and U662 (N_662,In_929,In_151);
nor U663 (N_663,In_1677,In_1240);
or U664 (N_664,In_712,In_198);
nand U665 (N_665,In_1333,In_1271);
and U666 (N_666,In_615,In_577);
and U667 (N_667,In_779,In_427);
or U668 (N_668,In_1400,In_132);
or U669 (N_669,In_409,In_146);
nand U670 (N_670,In_431,In_1254);
and U671 (N_671,In_1032,In_363);
and U672 (N_672,In_1360,In_573);
or U673 (N_673,In_1136,In_496);
or U674 (N_674,In_1510,In_993);
and U675 (N_675,In_954,In_644);
and U676 (N_676,In_1842,In_40);
nor U677 (N_677,In_1992,In_664);
xnor U678 (N_678,In_1027,In_1989);
nor U679 (N_679,In_259,In_715);
and U680 (N_680,In_1836,In_1013);
or U681 (N_681,In_1367,In_1914);
or U682 (N_682,In_1155,In_159);
and U683 (N_683,In_1471,In_1937);
and U684 (N_684,In_1049,In_35);
nor U685 (N_685,In_1673,In_5);
nand U686 (N_686,In_347,In_959);
nor U687 (N_687,In_1694,In_192);
xor U688 (N_688,In_455,In_164);
nor U689 (N_689,In_894,In_505);
nand U690 (N_690,In_268,In_1741);
or U691 (N_691,In_1555,In_750);
or U692 (N_692,In_1831,In_1920);
nor U693 (N_693,In_1807,In_1473);
nand U694 (N_694,In_527,In_1895);
and U695 (N_695,In_704,In_1636);
nor U696 (N_696,In_542,In_1607);
nand U697 (N_697,In_150,In_667);
nor U698 (N_698,In_1545,In_261);
nand U699 (N_699,In_1121,In_384);
and U700 (N_700,In_1721,In_1873);
and U701 (N_701,In_299,In_1004);
xnor U702 (N_702,In_214,In_521);
and U703 (N_703,In_229,In_1801);
or U704 (N_704,In_1180,In_1368);
xor U705 (N_705,In_178,In_1919);
and U706 (N_706,In_1120,In_1570);
and U707 (N_707,In_273,In_436);
and U708 (N_708,In_769,In_112);
nand U709 (N_709,In_646,In_1666);
and U710 (N_710,In_1637,In_1002);
and U711 (N_711,In_1445,In_215);
nand U712 (N_712,In_1311,In_623);
xnor U713 (N_713,In_1295,In_281);
xor U714 (N_714,In_1977,In_6);
xor U715 (N_715,In_1383,In_1926);
or U716 (N_716,In_658,In_25);
nand U717 (N_717,In_1639,In_1549);
nor U718 (N_718,In_54,In_81);
and U719 (N_719,In_548,In_304);
or U720 (N_720,In_446,In_1683);
xor U721 (N_721,In_1662,In_731);
nand U722 (N_722,In_1397,In_1638);
or U723 (N_723,In_1548,In_614);
nor U724 (N_724,In_1116,In_9);
nor U725 (N_725,In_82,In_470);
xor U726 (N_726,In_1348,In_1420);
or U727 (N_727,In_1215,In_242);
or U728 (N_728,In_1151,In_217);
xnor U729 (N_729,In_552,In_558);
nor U730 (N_730,In_1090,In_1147);
nand U731 (N_731,In_689,In_84);
and U732 (N_732,In_310,In_931);
nor U733 (N_733,In_1751,In_1279);
or U734 (N_734,In_541,In_1326);
nor U735 (N_735,In_459,In_1206);
nand U736 (N_736,In_1284,In_879);
xnor U737 (N_737,In_1495,In_827);
nor U738 (N_738,In_628,In_1175);
or U739 (N_739,In_620,In_930);
nor U740 (N_740,In_235,In_1564);
nor U741 (N_741,In_435,In_1292);
and U742 (N_742,In_557,In_1905);
nand U743 (N_743,In_78,In_920);
xnor U744 (N_744,In_1209,In_537);
and U745 (N_745,In_1415,In_1969);
nand U746 (N_746,In_20,In_1419);
nand U747 (N_747,In_255,In_354);
or U748 (N_748,In_336,In_227);
nand U749 (N_749,In_876,In_1479);
xor U750 (N_750,In_429,In_697);
nand U751 (N_751,In_1674,In_1699);
nand U752 (N_752,In_186,In_19);
nor U753 (N_753,In_1613,In_1014);
or U754 (N_754,In_70,In_108);
or U755 (N_755,In_1543,In_315);
nand U756 (N_756,In_1660,In_1840);
xor U757 (N_757,In_1994,In_1537);
xor U758 (N_758,In_1020,In_1940);
nand U759 (N_759,In_1036,In_1941);
xor U760 (N_760,In_38,In_502);
nand U761 (N_761,In_68,In_1816);
and U762 (N_762,In_1258,In_1735);
xnor U763 (N_763,In_339,In_768);
nand U764 (N_764,In_1259,In_106);
or U765 (N_765,In_1388,In_651);
nor U766 (N_766,In_811,In_77);
nand U767 (N_767,In_1167,In_1512);
nor U768 (N_768,In_239,In_419);
or U769 (N_769,In_1742,In_1522);
and U770 (N_770,In_1514,In_589);
xnor U771 (N_771,In_1737,In_854);
or U772 (N_772,In_1366,In_808);
xor U773 (N_773,In_1329,In_27);
nand U774 (N_774,In_1912,In_21);
nor U775 (N_775,In_1707,In_1559);
nor U776 (N_776,In_199,In_770);
nand U777 (N_777,In_1346,In_200);
nand U778 (N_778,In_941,In_1184);
or U779 (N_779,In_51,In_293);
and U780 (N_780,In_208,In_1380);
and U781 (N_781,In_1713,In_1126);
or U782 (N_782,In_372,In_632);
or U783 (N_783,In_1197,In_858);
nor U784 (N_784,In_1339,In_1130);
xnor U785 (N_785,In_324,In_1222);
and U786 (N_786,In_296,In_325);
or U787 (N_787,In_1227,In_1306);
nand U788 (N_788,In_642,In_1034);
or U789 (N_789,In_711,In_807);
xnor U790 (N_790,In_98,In_191);
nand U791 (N_791,In_464,In_1302);
nor U792 (N_792,In_1242,In_1614);
nand U793 (N_793,In_536,In_43);
nand U794 (N_794,In_829,In_276);
xnor U795 (N_795,In_1571,In_728);
nand U796 (N_796,In_648,In_380);
and U797 (N_797,In_1833,In_870);
nand U798 (N_798,In_631,In_1975);
nor U799 (N_799,In_1317,In_1492);
xor U800 (N_800,In_65,In_1536);
xor U801 (N_801,In_1622,In_493);
nor U802 (N_802,In_1275,In_1635);
and U803 (N_803,In_89,In_1038);
nor U804 (N_804,In_1857,In_230);
and U805 (N_805,In_888,In_745);
nor U806 (N_806,In_1008,In_507);
or U807 (N_807,In_892,In_478);
nand U808 (N_808,In_1950,In_1766);
nor U809 (N_809,In_576,In_156);
and U810 (N_810,In_433,In_1851);
nand U811 (N_811,In_629,In_1395);
and U812 (N_812,In_709,In_225);
or U813 (N_813,In_1330,In_1118);
nor U814 (N_814,In_1705,In_990);
nand U815 (N_815,In_226,In_816);
or U816 (N_816,In_1061,In_69);
nand U817 (N_817,In_1574,In_1566);
nor U818 (N_818,In_187,In_1732);
nor U819 (N_819,In_1615,In_1829);
or U820 (N_820,In_1309,In_73);
and U821 (N_821,In_1041,In_1462);
or U822 (N_822,In_280,In_1239);
nand U823 (N_823,In_1100,In_744);
and U824 (N_824,In_319,In_1246);
xor U825 (N_825,In_179,In_1363);
and U826 (N_826,In_206,In_1610);
nand U827 (N_827,In_1974,In_1954);
xnor U828 (N_828,In_1289,In_295);
nand U829 (N_829,In_1241,In_1949);
nor U830 (N_830,In_417,In_1224);
nor U831 (N_831,In_856,In_611);
and U832 (N_832,In_115,In_1101);
and U833 (N_833,In_1689,In_1885);
and U834 (N_834,In_1432,In_1886);
or U835 (N_835,In_1345,In_55);
and U836 (N_836,In_425,In_1378);
and U837 (N_837,In_1814,In_1016);
or U838 (N_838,In_1651,In_1412);
nor U839 (N_839,In_1447,In_1884);
nand U840 (N_840,In_819,In_1953);
nor U841 (N_841,In_1055,In_434);
or U842 (N_842,In_1697,In_1162);
nor U843 (N_843,In_1774,In_260);
nand U844 (N_844,In_377,In_223);
and U845 (N_845,In_1109,In_995);
nand U846 (N_846,In_1253,In_529);
nor U847 (N_847,In_714,In_1474);
nor U848 (N_848,In_1667,In_1772);
or U849 (N_849,In_1498,In_302);
and U850 (N_850,In_173,In_1316);
nor U851 (N_851,In_1066,In_1556);
nor U852 (N_852,In_1661,In_617);
nor U853 (N_853,In_1375,In_1113);
and U854 (N_854,In_1372,In_1371);
xor U855 (N_855,In_1870,In_1709);
nor U856 (N_856,In_501,In_1313);
or U857 (N_857,In_902,In_1177);
and U858 (N_858,In_122,In_1552);
or U859 (N_859,In_1750,In_1643);
nor U860 (N_860,In_1685,In_1966);
and U861 (N_861,In_264,In_546);
and U862 (N_862,In_1902,In_1585);
or U863 (N_863,In_1379,In_11);
nor U864 (N_864,In_330,In_1818);
nor U865 (N_865,In_1722,In_1825);
nor U866 (N_866,In_1308,In_1871);
and U867 (N_867,In_170,In_1773);
nand U868 (N_868,In_561,In_776);
or U869 (N_869,In_726,In_1349);
or U870 (N_870,In_358,In_924);
nand U871 (N_871,In_140,In_923);
and U872 (N_872,In_1509,In_685);
nand U873 (N_873,In_717,In_1074);
nand U874 (N_874,In_1738,In_437);
nor U875 (N_875,In_616,In_1338);
nor U876 (N_876,In_1437,In_1199);
nor U877 (N_877,In_412,In_1799);
nand U878 (N_878,In_1260,In_1898);
nand U879 (N_879,In_1908,In_986);
nor U880 (N_880,In_1982,In_1208);
xor U881 (N_881,In_1962,In_1746);
nand U882 (N_882,In_1753,In_1604);
nor U883 (N_883,In_1553,In_251);
nor U884 (N_884,In_397,In_348);
or U885 (N_885,In_197,In_1881);
and U886 (N_886,In_873,In_1464);
nand U887 (N_887,In_374,In_532);
nor U888 (N_888,In_793,In_190);
and U889 (N_889,In_1845,In_52);
and U890 (N_890,In_701,In_1540);
or U891 (N_891,In_488,In_439);
or U892 (N_892,In_1453,In_1174);
or U893 (N_893,In_1469,In_1218);
or U894 (N_894,In_1280,In_1018);
xnor U895 (N_895,In_906,In_581);
nand U896 (N_896,In_1702,In_526);
or U897 (N_897,In_1672,In_834);
and U898 (N_898,In_756,In_1964);
nand U899 (N_899,In_1986,In_1859);
or U900 (N_900,In_1889,In_1108);
and U901 (N_901,In_1535,In_1456);
and U902 (N_902,In_820,In_859);
or U903 (N_903,In_1405,In_833);
and U904 (N_904,In_1706,In_965);
and U905 (N_905,In_1472,In_1470);
or U906 (N_906,In_1463,In_1875);
nor U907 (N_907,In_1423,In_707);
nor U908 (N_908,In_80,In_910);
xor U909 (N_909,In_1561,In_1079);
xnor U910 (N_910,In_1560,In_193);
or U911 (N_911,In_864,In_1228);
and U912 (N_912,In_1232,In_444);
nand U913 (N_913,In_723,In_1039);
nor U914 (N_914,In_1265,In_1030);
or U915 (N_915,In_972,In_1928);
and U916 (N_916,In_785,In_1436);
nand U917 (N_917,In_1183,In_562);
nor U918 (N_918,In_287,In_1983);
or U919 (N_919,In_991,In_1021);
xor U920 (N_920,In_1867,In_262);
or U921 (N_921,In_1956,In_189);
nor U922 (N_922,In_915,In_1815);
nor U923 (N_923,In_96,In_1687);
xnor U924 (N_924,In_839,In_1968);
nand U925 (N_925,In_1403,In_566);
nand U926 (N_926,In_587,In_458);
nor U927 (N_927,In_487,In_401);
or U928 (N_928,In_362,In_604);
nand U929 (N_929,In_641,In_1324);
and U930 (N_930,In_564,In_1792);
and U931 (N_931,In_925,In_246);
nand U932 (N_932,In_118,In_369);
nand U933 (N_933,In_962,In_796);
nand U934 (N_934,In_1839,In_176);
or U935 (N_935,In_1288,In_825);
nor U936 (N_936,In_674,In_1678);
nor U937 (N_937,In_1035,In_1404);
nor U938 (N_938,In_1164,In_767);
and U939 (N_939,In_1429,In_814);
or U940 (N_940,In_1849,In_1917);
and U941 (N_941,In_1605,In_361);
nand U942 (N_942,In_1644,In_1391);
nor U943 (N_943,In_1211,In_322);
or U944 (N_944,In_93,In_1276);
or U945 (N_945,In_1987,In_1835);
nor U946 (N_946,In_1617,In_1281);
nand U947 (N_947,In_1087,In_901);
or U948 (N_948,In_553,In_1461);
and U949 (N_949,In_465,In_1484);
nand U950 (N_950,In_148,In_107);
or U951 (N_951,In_1904,In_26);
nand U952 (N_952,In_1834,In_1811);
nand U953 (N_953,In_396,In_123);
nor U954 (N_954,In_249,In_1207);
and U955 (N_955,In_48,In_772);
nor U956 (N_956,In_842,In_1396);
nor U957 (N_957,In_788,In_983);
nor U958 (N_958,In_511,In_1872);
or U959 (N_959,In_12,In_1446);
nor U960 (N_960,In_388,In_1223);
xnor U961 (N_961,In_1007,In_751);
nor U962 (N_962,In_1005,In_1154);
and U963 (N_963,In_1876,In_1791);
nor U964 (N_964,In_1263,In_256);
nor U965 (N_965,In_124,In_484);
nand U966 (N_966,In_592,In_1830);
and U967 (N_967,In_1955,In_783);
nand U968 (N_968,In_1003,In_1731);
nor U969 (N_969,In_741,In_1653);
nor U970 (N_970,In_423,In_1341);
nor U971 (N_971,In_899,In_1784);
nand U972 (N_972,In_585,In_982);
or U973 (N_973,In_1293,In_1468);
nor U974 (N_974,In_231,In_356);
nor U975 (N_975,In_992,In_441);
and U976 (N_976,In_174,In_740);
nor U977 (N_977,In_428,In_603);
nor U978 (N_978,In_1059,In_1115);
or U979 (N_979,In_1787,In_495);
and U980 (N_980,In_1679,In_30);
or U981 (N_981,In_1965,In_677);
or U982 (N_982,In_387,In_143);
nand U983 (N_983,In_10,In_1828);
nor U984 (N_984,In_1596,In_371);
nor U985 (N_985,In_692,In_835);
nor U986 (N_986,In_334,In_389);
nor U987 (N_987,In_1796,In_1392);
or U988 (N_988,In_117,In_1646);
nand U989 (N_989,In_1448,In_609);
nand U990 (N_990,In_1922,In_1022);
or U991 (N_991,In_968,In_1012);
and U992 (N_992,In_1194,In_451);
nand U993 (N_993,In_1580,In_1425);
and U994 (N_994,In_960,In_392);
and U995 (N_995,In_855,In_1088);
or U996 (N_996,In_1123,In_31);
and U997 (N_997,In_1597,In_1565);
nand U998 (N_998,In_886,In_1567);
nor U999 (N_999,In_649,In_1659);
nor U1000 (N_1000,In_55,In_1714);
or U1001 (N_1001,In_1447,In_304);
nor U1002 (N_1002,In_626,In_533);
nand U1003 (N_1003,In_1747,In_1743);
or U1004 (N_1004,In_1921,In_1251);
and U1005 (N_1005,In_1685,In_27);
nand U1006 (N_1006,In_1869,In_1075);
and U1007 (N_1007,In_185,In_217);
nand U1008 (N_1008,In_402,In_74);
and U1009 (N_1009,In_1172,In_1929);
and U1010 (N_1010,In_1268,In_1892);
and U1011 (N_1011,In_1297,In_1216);
and U1012 (N_1012,In_1004,In_1861);
nand U1013 (N_1013,In_1174,In_1759);
nor U1014 (N_1014,In_1728,In_253);
and U1015 (N_1015,In_403,In_910);
nand U1016 (N_1016,In_821,In_1219);
or U1017 (N_1017,In_651,In_1400);
or U1018 (N_1018,In_415,In_1605);
xnor U1019 (N_1019,In_1185,In_1158);
nor U1020 (N_1020,In_101,In_1977);
and U1021 (N_1021,In_1145,In_1873);
xnor U1022 (N_1022,In_1956,In_463);
or U1023 (N_1023,In_991,In_594);
nor U1024 (N_1024,In_967,In_692);
xor U1025 (N_1025,In_772,In_938);
and U1026 (N_1026,In_307,In_541);
xor U1027 (N_1027,In_1560,In_1375);
or U1028 (N_1028,In_1685,In_1038);
nand U1029 (N_1029,In_1108,In_509);
and U1030 (N_1030,In_1149,In_1068);
or U1031 (N_1031,In_1000,In_1710);
and U1032 (N_1032,In_969,In_739);
xnor U1033 (N_1033,In_1424,In_871);
or U1034 (N_1034,In_1643,In_1892);
nand U1035 (N_1035,In_1775,In_376);
and U1036 (N_1036,In_221,In_96);
nor U1037 (N_1037,In_1085,In_198);
and U1038 (N_1038,In_1832,In_1333);
and U1039 (N_1039,In_138,In_1852);
and U1040 (N_1040,In_1098,In_1184);
or U1041 (N_1041,In_1254,In_739);
nor U1042 (N_1042,In_710,In_954);
nor U1043 (N_1043,In_946,In_892);
nand U1044 (N_1044,In_295,In_1507);
nor U1045 (N_1045,In_941,In_1512);
nand U1046 (N_1046,In_421,In_136);
nand U1047 (N_1047,In_620,In_1827);
or U1048 (N_1048,In_582,In_1185);
and U1049 (N_1049,In_300,In_896);
xor U1050 (N_1050,In_754,In_573);
and U1051 (N_1051,In_1953,In_689);
nor U1052 (N_1052,In_1831,In_1990);
nor U1053 (N_1053,In_318,In_1123);
and U1054 (N_1054,In_200,In_1308);
and U1055 (N_1055,In_291,In_1080);
nor U1056 (N_1056,In_1728,In_1681);
or U1057 (N_1057,In_1242,In_74);
nand U1058 (N_1058,In_593,In_991);
and U1059 (N_1059,In_1775,In_130);
and U1060 (N_1060,In_959,In_1247);
or U1061 (N_1061,In_1877,In_890);
nand U1062 (N_1062,In_829,In_1664);
and U1063 (N_1063,In_1904,In_649);
xor U1064 (N_1064,In_80,In_1824);
or U1065 (N_1065,In_1344,In_1778);
nand U1066 (N_1066,In_1510,In_1228);
and U1067 (N_1067,In_512,In_1519);
and U1068 (N_1068,In_552,In_392);
xor U1069 (N_1069,In_938,In_437);
nand U1070 (N_1070,In_89,In_69);
nor U1071 (N_1071,In_193,In_1696);
nor U1072 (N_1072,In_752,In_1078);
and U1073 (N_1073,In_1375,In_1499);
and U1074 (N_1074,In_1728,In_108);
nand U1075 (N_1075,In_961,In_1634);
or U1076 (N_1076,In_201,In_661);
xor U1077 (N_1077,In_1536,In_1502);
nand U1078 (N_1078,In_905,In_306);
and U1079 (N_1079,In_229,In_1750);
nor U1080 (N_1080,In_268,In_1841);
or U1081 (N_1081,In_1696,In_1346);
and U1082 (N_1082,In_1833,In_1318);
nand U1083 (N_1083,In_471,In_1568);
and U1084 (N_1084,In_114,In_417);
nor U1085 (N_1085,In_1869,In_792);
nor U1086 (N_1086,In_808,In_87);
xor U1087 (N_1087,In_457,In_667);
nor U1088 (N_1088,In_995,In_1759);
nor U1089 (N_1089,In_1496,In_83);
or U1090 (N_1090,In_1618,In_1009);
and U1091 (N_1091,In_1518,In_1795);
or U1092 (N_1092,In_1543,In_963);
or U1093 (N_1093,In_918,In_1709);
nand U1094 (N_1094,In_1006,In_457);
or U1095 (N_1095,In_1454,In_1368);
nor U1096 (N_1096,In_1042,In_1772);
nor U1097 (N_1097,In_769,In_614);
nor U1098 (N_1098,In_1599,In_1286);
or U1099 (N_1099,In_1793,In_181);
and U1100 (N_1100,In_548,In_1236);
nand U1101 (N_1101,In_1964,In_1873);
nand U1102 (N_1102,In_1421,In_986);
or U1103 (N_1103,In_269,In_258);
nand U1104 (N_1104,In_378,In_301);
nand U1105 (N_1105,In_315,In_1443);
nand U1106 (N_1106,In_1573,In_1845);
nor U1107 (N_1107,In_555,In_896);
and U1108 (N_1108,In_1539,In_838);
and U1109 (N_1109,In_1640,In_1159);
xor U1110 (N_1110,In_811,In_49);
nor U1111 (N_1111,In_546,In_1794);
nand U1112 (N_1112,In_860,In_942);
nand U1113 (N_1113,In_553,In_969);
xor U1114 (N_1114,In_159,In_854);
nor U1115 (N_1115,In_1372,In_289);
nor U1116 (N_1116,In_1464,In_1399);
nand U1117 (N_1117,In_1885,In_736);
or U1118 (N_1118,In_1192,In_1055);
and U1119 (N_1119,In_131,In_1939);
and U1120 (N_1120,In_1767,In_894);
nor U1121 (N_1121,In_1905,In_1766);
nand U1122 (N_1122,In_1784,In_1067);
nand U1123 (N_1123,In_1159,In_1726);
or U1124 (N_1124,In_295,In_820);
nand U1125 (N_1125,In_1968,In_1681);
nor U1126 (N_1126,In_710,In_1909);
nor U1127 (N_1127,In_1959,In_515);
nand U1128 (N_1128,In_530,In_1917);
and U1129 (N_1129,In_1877,In_997);
nand U1130 (N_1130,In_1559,In_1433);
nand U1131 (N_1131,In_654,In_339);
and U1132 (N_1132,In_643,In_1795);
or U1133 (N_1133,In_1223,In_1099);
nor U1134 (N_1134,In_207,In_279);
xor U1135 (N_1135,In_1697,In_1114);
or U1136 (N_1136,In_617,In_358);
and U1137 (N_1137,In_680,In_1937);
or U1138 (N_1138,In_779,In_526);
xnor U1139 (N_1139,In_345,In_1392);
and U1140 (N_1140,In_304,In_199);
nor U1141 (N_1141,In_1696,In_431);
nor U1142 (N_1142,In_1828,In_1100);
xor U1143 (N_1143,In_1446,In_1107);
nor U1144 (N_1144,In_1732,In_330);
nand U1145 (N_1145,In_428,In_1401);
or U1146 (N_1146,In_989,In_1913);
nor U1147 (N_1147,In_1481,In_689);
and U1148 (N_1148,In_306,In_1182);
or U1149 (N_1149,In_986,In_1108);
nor U1150 (N_1150,In_1938,In_283);
xor U1151 (N_1151,In_565,In_1963);
nor U1152 (N_1152,In_771,In_537);
and U1153 (N_1153,In_1193,In_166);
or U1154 (N_1154,In_247,In_430);
or U1155 (N_1155,In_342,In_110);
nand U1156 (N_1156,In_1905,In_355);
nor U1157 (N_1157,In_760,In_1994);
or U1158 (N_1158,In_378,In_658);
nand U1159 (N_1159,In_55,In_1335);
nand U1160 (N_1160,In_746,In_1713);
nor U1161 (N_1161,In_989,In_1288);
or U1162 (N_1162,In_855,In_1360);
or U1163 (N_1163,In_56,In_1870);
nor U1164 (N_1164,In_134,In_1453);
and U1165 (N_1165,In_38,In_1652);
and U1166 (N_1166,In_174,In_1400);
or U1167 (N_1167,In_1584,In_1829);
nor U1168 (N_1168,In_237,In_646);
and U1169 (N_1169,In_898,In_647);
or U1170 (N_1170,In_1562,In_1561);
nor U1171 (N_1171,In_549,In_1493);
xnor U1172 (N_1172,In_643,In_1425);
nand U1173 (N_1173,In_527,In_1899);
nand U1174 (N_1174,In_331,In_816);
nand U1175 (N_1175,In_304,In_217);
and U1176 (N_1176,In_1691,In_1696);
xnor U1177 (N_1177,In_714,In_1479);
nor U1178 (N_1178,In_738,In_547);
nor U1179 (N_1179,In_1395,In_737);
or U1180 (N_1180,In_1882,In_180);
xnor U1181 (N_1181,In_683,In_216);
nand U1182 (N_1182,In_992,In_1779);
or U1183 (N_1183,In_1030,In_1820);
or U1184 (N_1184,In_202,In_1303);
and U1185 (N_1185,In_1395,In_653);
or U1186 (N_1186,In_282,In_1493);
nand U1187 (N_1187,In_848,In_923);
xor U1188 (N_1188,In_472,In_922);
nor U1189 (N_1189,In_423,In_1113);
and U1190 (N_1190,In_177,In_1732);
and U1191 (N_1191,In_963,In_76);
xnor U1192 (N_1192,In_247,In_715);
xnor U1193 (N_1193,In_949,In_1601);
xnor U1194 (N_1194,In_1635,In_638);
or U1195 (N_1195,In_451,In_652);
nand U1196 (N_1196,In_1762,In_1295);
nor U1197 (N_1197,In_776,In_706);
or U1198 (N_1198,In_433,In_135);
nor U1199 (N_1199,In_1881,In_1107);
or U1200 (N_1200,In_491,In_351);
or U1201 (N_1201,In_317,In_270);
nand U1202 (N_1202,In_532,In_929);
or U1203 (N_1203,In_234,In_1898);
nor U1204 (N_1204,In_1020,In_802);
xnor U1205 (N_1205,In_1938,In_1447);
nor U1206 (N_1206,In_1189,In_194);
nor U1207 (N_1207,In_1870,In_808);
nand U1208 (N_1208,In_1698,In_620);
nand U1209 (N_1209,In_1139,In_118);
and U1210 (N_1210,In_1231,In_648);
nor U1211 (N_1211,In_1734,In_430);
nand U1212 (N_1212,In_46,In_1402);
nor U1213 (N_1213,In_1251,In_100);
nor U1214 (N_1214,In_685,In_2);
nand U1215 (N_1215,In_1818,In_362);
nor U1216 (N_1216,In_83,In_1174);
and U1217 (N_1217,In_444,In_478);
nor U1218 (N_1218,In_295,In_1912);
nor U1219 (N_1219,In_845,In_72);
or U1220 (N_1220,In_1759,In_316);
nand U1221 (N_1221,In_480,In_569);
nor U1222 (N_1222,In_1883,In_502);
or U1223 (N_1223,In_326,In_1140);
nor U1224 (N_1224,In_129,In_1460);
or U1225 (N_1225,In_1938,In_1083);
nor U1226 (N_1226,In_22,In_1233);
nor U1227 (N_1227,In_279,In_289);
or U1228 (N_1228,In_1129,In_1307);
or U1229 (N_1229,In_1379,In_586);
nand U1230 (N_1230,In_603,In_1506);
nand U1231 (N_1231,In_1140,In_206);
nand U1232 (N_1232,In_242,In_1227);
and U1233 (N_1233,In_431,In_945);
or U1234 (N_1234,In_183,In_710);
nor U1235 (N_1235,In_144,In_1348);
nor U1236 (N_1236,In_1477,In_368);
nand U1237 (N_1237,In_1581,In_79);
nand U1238 (N_1238,In_180,In_110);
nand U1239 (N_1239,In_74,In_894);
nor U1240 (N_1240,In_1447,In_384);
nand U1241 (N_1241,In_1413,In_1080);
and U1242 (N_1242,In_509,In_1727);
and U1243 (N_1243,In_737,In_1857);
nor U1244 (N_1244,In_458,In_1116);
and U1245 (N_1245,In_1838,In_1599);
and U1246 (N_1246,In_477,In_1366);
and U1247 (N_1247,In_1995,In_1166);
nor U1248 (N_1248,In_957,In_626);
or U1249 (N_1249,In_884,In_543);
and U1250 (N_1250,In_282,In_311);
and U1251 (N_1251,In_18,In_1965);
or U1252 (N_1252,In_722,In_1639);
and U1253 (N_1253,In_1841,In_754);
and U1254 (N_1254,In_1490,In_985);
nand U1255 (N_1255,In_1250,In_1806);
xor U1256 (N_1256,In_1874,In_1811);
nand U1257 (N_1257,In_593,In_6);
nand U1258 (N_1258,In_98,In_605);
nand U1259 (N_1259,In_1954,In_142);
or U1260 (N_1260,In_1672,In_748);
and U1261 (N_1261,In_495,In_1488);
or U1262 (N_1262,In_1014,In_123);
nand U1263 (N_1263,In_1060,In_1861);
nor U1264 (N_1264,In_1573,In_238);
nor U1265 (N_1265,In_592,In_1456);
nand U1266 (N_1266,In_1656,In_1648);
and U1267 (N_1267,In_255,In_1863);
or U1268 (N_1268,In_367,In_618);
or U1269 (N_1269,In_1816,In_1469);
nor U1270 (N_1270,In_1522,In_380);
nor U1271 (N_1271,In_562,In_144);
or U1272 (N_1272,In_401,In_1509);
nor U1273 (N_1273,In_546,In_395);
nor U1274 (N_1274,In_1420,In_559);
or U1275 (N_1275,In_228,In_1932);
or U1276 (N_1276,In_1632,In_435);
xor U1277 (N_1277,In_1206,In_721);
or U1278 (N_1278,In_1666,In_1112);
xor U1279 (N_1279,In_1477,In_1134);
nor U1280 (N_1280,In_602,In_223);
or U1281 (N_1281,In_1233,In_550);
or U1282 (N_1282,In_1656,In_912);
and U1283 (N_1283,In_1241,In_1523);
nor U1284 (N_1284,In_1554,In_1613);
and U1285 (N_1285,In_1922,In_1426);
nor U1286 (N_1286,In_883,In_1467);
and U1287 (N_1287,In_759,In_1896);
nand U1288 (N_1288,In_1409,In_1479);
xnor U1289 (N_1289,In_1905,In_1582);
and U1290 (N_1290,In_1035,In_792);
nor U1291 (N_1291,In_1913,In_1102);
nand U1292 (N_1292,In_75,In_131);
xnor U1293 (N_1293,In_412,In_1043);
nand U1294 (N_1294,In_434,In_1462);
and U1295 (N_1295,In_1458,In_1697);
or U1296 (N_1296,In_1286,In_1678);
or U1297 (N_1297,In_1260,In_585);
or U1298 (N_1298,In_406,In_1943);
nand U1299 (N_1299,In_1092,In_1239);
nor U1300 (N_1300,In_1190,In_1894);
or U1301 (N_1301,In_22,In_1128);
nand U1302 (N_1302,In_1929,In_1341);
or U1303 (N_1303,In_403,In_460);
or U1304 (N_1304,In_44,In_1459);
nor U1305 (N_1305,In_717,In_1459);
nand U1306 (N_1306,In_1859,In_1192);
and U1307 (N_1307,In_1391,In_1442);
or U1308 (N_1308,In_326,In_1392);
nor U1309 (N_1309,In_17,In_1705);
or U1310 (N_1310,In_975,In_1726);
nor U1311 (N_1311,In_1560,In_1195);
nor U1312 (N_1312,In_1523,In_659);
nand U1313 (N_1313,In_213,In_1036);
nand U1314 (N_1314,In_800,In_1051);
nand U1315 (N_1315,In_1659,In_827);
nor U1316 (N_1316,In_891,In_1200);
or U1317 (N_1317,In_1671,In_1575);
and U1318 (N_1318,In_920,In_1377);
and U1319 (N_1319,In_425,In_394);
nor U1320 (N_1320,In_1644,In_270);
and U1321 (N_1321,In_1326,In_442);
and U1322 (N_1322,In_1794,In_1275);
nand U1323 (N_1323,In_794,In_1574);
and U1324 (N_1324,In_996,In_736);
or U1325 (N_1325,In_1326,In_1684);
xor U1326 (N_1326,In_1963,In_221);
nand U1327 (N_1327,In_643,In_1803);
or U1328 (N_1328,In_1742,In_140);
nor U1329 (N_1329,In_1517,In_365);
or U1330 (N_1330,In_1357,In_691);
or U1331 (N_1331,In_5,In_1339);
or U1332 (N_1332,In_1460,In_1689);
xor U1333 (N_1333,In_1348,In_1845);
nand U1334 (N_1334,In_1226,In_745);
xor U1335 (N_1335,In_172,In_903);
and U1336 (N_1336,In_1283,In_1227);
and U1337 (N_1337,In_1214,In_185);
or U1338 (N_1338,In_940,In_973);
nand U1339 (N_1339,In_1005,In_281);
xor U1340 (N_1340,In_1730,In_951);
nand U1341 (N_1341,In_1943,In_1096);
nor U1342 (N_1342,In_1497,In_1170);
or U1343 (N_1343,In_249,In_356);
nor U1344 (N_1344,In_1279,In_73);
and U1345 (N_1345,In_1126,In_1969);
and U1346 (N_1346,In_1933,In_1128);
or U1347 (N_1347,In_372,In_976);
xor U1348 (N_1348,In_529,In_69);
nor U1349 (N_1349,In_355,In_821);
nor U1350 (N_1350,In_1203,In_1879);
or U1351 (N_1351,In_564,In_1676);
and U1352 (N_1352,In_873,In_520);
and U1353 (N_1353,In_713,In_1840);
xnor U1354 (N_1354,In_197,In_1085);
nor U1355 (N_1355,In_617,In_1925);
nor U1356 (N_1356,In_52,In_330);
xor U1357 (N_1357,In_1896,In_830);
or U1358 (N_1358,In_706,In_305);
and U1359 (N_1359,In_402,In_343);
nand U1360 (N_1360,In_644,In_33);
nor U1361 (N_1361,In_484,In_1527);
nor U1362 (N_1362,In_244,In_1196);
and U1363 (N_1363,In_1573,In_378);
or U1364 (N_1364,In_166,In_1346);
nand U1365 (N_1365,In_109,In_1248);
or U1366 (N_1366,In_1745,In_1292);
or U1367 (N_1367,In_108,In_472);
nor U1368 (N_1368,In_1675,In_132);
xor U1369 (N_1369,In_216,In_1227);
or U1370 (N_1370,In_1862,In_1011);
nand U1371 (N_1371,In_1399,In_1021);
nor U1372 (N_1372,In_316,In_1423);
nor U1373 (N_1373,In_982,In_1383);
nand U1374 (N_1374,In_1215,In_1733);
nor U1375 (N_1375,In_928,In_5);
or U1376 (N_1376,In_617,In_216);
nand U1377 (N_1377,In_1210,In_560);
and U1378 (N_1378,In_1789,In_1644);
nor U1379 (N_1379,In_804,In_1864);
or U1380 (N_1380,In_811,In_248);
and U1381 (N_1381,In_618,In_626);
nand U1382 (N_1382,In_318,In_867);
xnor U1383 (N_1383,In_975,In_84);
or U1384 (N_1384,In_1710,In_1391);
and U1385 (N_1385,In_1403,In_616);
nand U1386 (N_1386,In_148,In_1423);
nand U1387 (N_1387,In_599,In_676);
and U1388 (N_1388,In_528,In_452);
nor U1389 (N_1389,In_1849,In_1591);
nand U1390 (N_1390,In_376,In_708);
xor U1391 (N_1391,In_945,In_713);
and U1392 (N_1392,In_1717,In_157);
or U1393 (N_1393,In_239,In_426);
and U1394 (N_1394,In_1,In_449);
or U1395 (N_1395,In_591,In_499);
nor U1396 (N_1396,In_1526,In_103);
nand U1397 (N_1397,In_862,In_591);
nand U1398 (N_1398,In_1146,In_1754);
or U1399 (N_1399,In_1074,In_1899);
nand U1400 (N_1400,In_1412,In_1584);
xor U1401 (N_1401,In_1821,In_1977);
or U1402 (N_1402,In_1925,In_1966);
nor U1403 (N_1403,In_919,In_1824);
nand U1404 (N_1404,In_1916,In_371);
and U1405 (N_1405,In_235,In_1621);
or U1406 (N_1406,In_1674,In_810);
or U1407 (N_1407,In_347,In_1694);
or U1408 (N_1408,In_1458,In_829);
nor U1409 (N_1409,In_1177,In_802);
nand U1410 (N_1410,In_493,In_1534);
xor U1411 (N_1411,In_150,In_853);
nand U1412 (N_1412,In_1356,In_1303);
nor U1413 (N_1413,In_385,In_1974);
nand U1414 (N_1414,In_430,In_1222);
and U1415 (N_1415,In_1383,In_1646);
and U1416 (N_1416,In_1673,In_983);
xor U1417 (N_1417,In_1706,In_405);
xor U1418 (N_1418,In_404,In_1146);
and U1419 (N_1419,In_1463,In_720);
xnor U1420 (N_1420,In_1361,In_60);
nor U1421 (N_1421,In_885,In_738);
and U1422 (N_1422,In_475,In_980);
nor U1423 (N_1423,In_1163,In_773);
nand U1424 (N_1424,In_1077,In_488);
nor U1425 (N_1425,In_960,In_835);
or U1426 (N_1426,In_542,In_1422);
or U1427 (N_1427,In_793,In_857);
nor U1428 (N_1428,In_1381,In_1523);
and U1429 (N_1429,In_1100,In_453);
nand U1430 (N_1430,In_124,In_1749);
and U1431 (N_1431,In_18,In_715);
nor U1432 (N_1432,In_303,In_371);
nand U1433 (N_1433,In_814,In_1272);
nand U1434 (N_1434,In_758,In_1843);
and U1435 (N_1435,In_1141,In_336);
and U1436 (N_1436,In_176,In_850);
or U1437 (N_1437,In_1031,In_253);
nand U1438 (N_1438,In_1224,In_1617);
and U1439 (N_1439,In_339,In_926);
or U1440 (N_1440,In_1680,In_234);
nor U1441 (N_1441,In_746,In_1101);
nor U1442 (N_1442,In_641,In_1999);
and U1443 (N_1443,In_1752,In_727);
nor U1444 (N_1444,In_305,In_1151);
nor U1445 (N_1445,In_881,In_337);
or U1446 (N_1446,In_371,In_1827);
or U1447 (N_1447,In_312,In_316);
nand U1448 (N_1448,In_920,In_943);
nand U1449 (N_1449,In_1556,In_1759);
or U1450 (N_1450,In_1264,In_792);
nand U1451 (N_1451,In_1518,In_980);
or U1452 (N_1452,In_1642,In_482);
nand U1453 (N_1453,In_325,In_521);
nand U1454 (N_1454,In_1855,In_559);
nor U1455 (N_1455,In_506,In_530);
nand U1456 (N_1456,In_1051,In_1728);
xor U1457 (N_1457,In_1353,In_1752);
nor U1458 (N_1458,In_1094,In_868);
nor U1459 (N_1459,In_482,In_1387);
or U1460 (N_1460,In_1522,In_452);
nand U1461 (N_1461,In_179,In_1132);
or U1462 (N_1462,In_831,In_584);
nand U1463 (N_1463,In_1789,In_548);
nand U1464 (N_1464,In_1810,In_1683);
nor U1465 (N_1465,In_1444,In_1098);
nor U1466 (N_1466,In_1655,In_1732);
and U1467 (N_1467,In_409,In_989);
and U1468 (N_1468,In_118,In_1481);
or U1469 (N_1469,In_588,In_867);
nand U1470 (N_1470,In_646,In_1085);
nand U1471 (N_1471,In_593,In_1105);
and U1472 (N_1472,In_78,In_118);
nor U1473 (N_1473,In_793,In_424);
or U1474 (N_1474,In_964,In_13);
or U1475 (N_1475,In_1033,In_366);
and U1476 (N_1476,In_1758,In_1201);
nor U1477 (N_1477,In_135,In_229);
or U1478 (N_1478,In_1126,In_1859);
nor U1479 (N_1479,In_205,In_1231);
and U1480 (N_1480,In_22,In_1302);
nand U1481 (N_1481,In_799,In_1062);
or U1482 (N_1482,In_1528,In_134);
nor U1483 (N_1483,In_496,In_273);
or U1484 (N_1484,In_872,In_242);
and U1485 (N_1485,In_801,In_408);
and U1486 (N_1486,In_847,In_651);
nand U1487 (N_1487,In_702,In_179);
and U1488 (N_1488,In_1622,In_1991);
xnor U1489 (N_1489,In_741,In_937);
or U1490 (N_1490,In_512,In_764);
nand U1491 (N_1491,In_1723,In_1498);
xor U1492 (N_1492,In_1981,In_1224);
nand U1493 (N_1493,In_1318,In_1387);
and U1494 (N_1494,In_1165,In_855);
nand U1495 (N_1495,In_719,In_1044);
or U1496 (N_1496,In_672,In_651);
and U1497 (N_1497,In_1548,In_704);
or U1498 (N_1498,In_1424,In_953);
nor U1499 (N_1499,In_308,In_1664);
nand U1500 (N_1500,In_1640,In_1649);
nor U1501 (N_1501,In_1723,In_1883);
nand U1502 (N_1502,In_1564,In_300);
or U1503 (N_1503,In_1192,In_642);
or U1504 (N_1504,In_1739,In_1623);
nor U1505 (N_1505,In_1856,In_1285);
nand U1506 (N_1506,In_627,In_515);
nand U1507 (N_1507,In_653,In_1845);
nand U1508 (N_1508,In_1707,In_466);
or U1509 (N_1509,In_1031,In_669);
nor U1510 (N_1510,In_705,In_1433);
nor U1511 (N_1511,In_1554,In_273);
nand U1512 (N_1512,In_577,In_972);
xnor U1513 (N_1513,In_655,In_1045);
nand U1514 (N_1514,In_579,In_1086);
nor U1515 (N_1515,In_291,In_1288);
nor U1516 (N_1516,In_978,In_888);
or U1517 (N_1517,In_635,In_436);
xor U1518 (N_1518,In_560,In_286);
nand U1519 (N_1519,In_253,In_703);
nor U1520 (N_1520,In_1274,In_413);
or U1521 (N_1521,In_99,In_277);
nand U1522 (N_1522,In_1885,In_1592);
nor U1523 (N_1523,In_1036,In_7);
xnor U1524 (N_1524,In_638,In_307);
nand U1525 (N_1525,In_912,In_1369);
or U1526 (N_1526,In_829,In_1540);
or U1527 (N_1527,In_1157,In_1757);
and U1528 (N_1528,In_1032,In_1586);
nand U1529 (N_1529,In_1096,In_242);
and U1530 (N_1530,In_912,In_628);
nor U1531 (N_1531,In_1378,In_1337);
or U1532 (N_1532,In_1730,In_146);
xnor U1533 (N_1533,In_245,In_583);
nor U1534 (N_1534,In_689,In_876);
nand U1535 (N_1535,In_453,In_1446);
or U1536 (N_1536,In_412,In_1251);
xnor U1537 (N_1537,In_644,In_1749);
and U1538 (N_1538,In_180,In_735);
or U1539 (N_1539,In_1945,In_49);
and U1540 (N_1540,In_4,In_1527);
or U1541 (N_1541,In_653,In_555);
nand U1542 (N_1542,In_1885,In_333);
nor U1543 (N_1543,In_1204,In_1991);
or U1544 (N_1544,In_339,In_864);
nand U1545 (N_1545,In_1630,In_964);
or U1546 (N_1546,In_57,In_1777);
nand U1547 (N_1547,In_874,In_1342);
xor U1548 (N_1548,In_74,In_500);
xnor U1549 (N_1549,In_151,In_1592);
xnor U1550 (N_1550,In_107,In_464);
and U1551 (N_1551,In_1335,In_982);
nor U1552 (N_1552,In_1658,In_550);
nand U1553 (N_1553,In_1098,In_1134);
nor U1554 (N_1554,In_1360,In_973);
or U1555 (N_1555,In_729,In_1520);
nand U1556 (N_1556,In_261,In_1342);
nand U1557 (N_1557,In_1356,In_1714);
and U1558 (N_1558,In_103,In_1016);
and U1559 (N_1559,In_163,In_224);
nor U1560 (N_1560,In_1556,In_347);
or U1561 (N_1561,In_1276,In_1996);
or U1562 (N_1562,In_1819,In_1270);
and U1563 (N_1563,In_1956,In_426);
nand U1564 (N_1564,In_464,In_10);
or U1565 (N_1565,In_611,In_1533);
nor U1566 (N_1566,In_1833,In_33);
nand U1567 (N_1567,In_1667,In_1585);
or U1568 (N_1568,In_1424,In_1446);
nor U1569 (N_1569,In_300,In_1853);
and U1570 (N_1570,In_1663,In_817);
or U1571 (N_1571,In_1638,In_1869);
nand U1572 (N_1572,In_243,In_807);
xnor U1573 (N_1573,In_1433,In_507);
nor U1574 (N_1574,In_1300,In_1618);
or U1575 (N_1575,In_934,In_405);
or U1576 (N_1576,In_8,In_1021);
nor U1577 (N_1577,In_1208,In_683);
nand U1578 (N_1578,In_1126,In_1142);
nand U1579 (N_1579,In_381,In_733);
and U1580 (N_1580,In_1626,In_522);
nor U1581 (N_1581,In_61,In_1469);
or U1582 (N_1582,In_572,In_500);
or U1583 (N_1583,In_1532,In_1543);
or U1584 (N_1584,In_422,In_661);
nand U1585 (N_1585,In_1003,In_52);
xnor U1586 (N_1586,In_237,In_1176);
nor U1587 (N_1587,In_1113,In_27);
and U1588 (N_1588,In_1715,In_1182);
and U1589 (N_1589,In_1968,In_1778);
or U1590 (N_1590,In_381,In_378);
and U1591 (N_1591,In_482,In_1737);
and U1592 (N_1592,In_225,In_1896);
or U1593 (N_1593,In_1236,In_1326);
and U1594 (N_1594,In_1644,In_1003);
nand U1595 (N_1595,In_77,In_997);
xor U1596 (N_1596,In_1404,In_1456);
and U1597 (N_1597,In_1182,In_891);
and U1598 (N_1598,In_1996,In_625);
nand U1599 (N_1599,In_562,In_1663);
nor U1600 (N_1600,In_703,In_528);
nand U1601 (N_1601,In_136,In_1101);
nand U1602 (N_1602,In_1496,In_1701);
xor U1603 (N_1603,In_155,In_611);
nand U1604 (N_1604,In_1884,In_568);
xnor U1605 (N_1605,In_605,In_520);
or U1606 (N_1606,In_341,In_490);
nor U1607 (N_1607,In_553,In_463);
nor U1608 (N_1608,In_552,In_1983);
nor U1609 (N_1609,In_1099,In_273);
and U1610 (N_1610,In_1380,In_147);
nor U1611 (N_1611,In_1252,In_457);
and U1612 (N_1612,In_1819,In_1418);
or U1613 (N_1613,In_838,In_699);
nor U1614 (N_1614,In_919,In_1913);
or U1615 (N_1615,In_1439,In_985);
or U1616 (N_1616,In_355,In_229);
or U1617 (N_1617,In_505,In_75);
or U1618 (N_1618,In_266,In_325);
or U1619 (N_1619,In_1918,In_1177);
nor U1620 (N_1620,In_1444,In_1183);
and U1621 (N_1621,In_1058,In_747);
nor U1622 (N_1622,In_1297,In_349);
or U1623 (N_1623,In_1728,In_1147);
xnor U1624 (N_1624,In_1763,In_34);
nor U1625 (N_1625,In_48,In_1231);
xnor U1626 (N_1626,In_41,In_1743);
nor U1627 (N_1627,In_564,In_741);
or U1628 (N_1628,In_1578,In_1889);
nor U1629 (N_1629,In_890,In_880);
or U1630 (N_1630,In_1933,In_684);
nor U1631 (N_1631,In_42,In_1233);
xnor U1632 (N_1632,In_1566,In_417);
nand U1633 (N_1633,In_1414,In_1709);
or U1634 (N_1634,In_1665,In_866);
nor U1635 (N_1635,In_1189,In_585);
nand U1636 (N_1636,In_1276,In_1907);
nand U1637 (N_1637,In_980,In_1827);
and U1638 (N_1638,In_403,In_634);
or U1639 (N_1639,In_113,In_783);
xnor U1640 (N_1640,In_76,In_1548);
nor U1641 (N_1641,In_1918,In_1099);
and U1642 (N_1642,In_130,In_493);
and U1643 (N_1643,In_428,In_1544);
xnor U1644 (N_1644,In_546,In_430);
or U1645 (N_1645,In_342,In_1919);
xor U1646 (N_1646,In_691,In_860);
or U1647 (N_1647,In_1511,In_21);
or U1648 (N_1648,In_373,In_1572);
and U1649 (N_1649,In_435,In_1283);
and U1650 (N_1650,In_629,In_1334);
or U1651 (N_1651,In_986,In_532);
nand U1652 (N_1652,In_1042,In_583);
or U1653 (N_1653,In_1534,In_358);
nand U1654 (N_1654,In_1058,In_399);
nor U1655 (N_1655,In_1488,In_446);
nand U1656 (N_1656,In_248,In_66);
and U1657 (N_1657,In_451,In_1744);
or U1658 (N_1658,In_1586,In_1547);
xnor U1659 (N_1659,In_1435,In_594);
nor U1660 (N_1660,In_1097,In_1932);
nor U1661 (N_1661,In_549,In_1789);
nand U1662 (N_1662,In_1556,In_1768);
and U1663 (N_1663,In_505,In_1107);
and U1664 (N_1664,In_1643,In_1318);
and U1665 (N_1665,In_162,In_1431);
nand U1666 (N_1666,In_85,In_603);
nor U1667 (N_1667,In_274,In_1561);
and U1668 (N_1668,In_1074,In_1161);
or U1669 (N_1669,In_1171,In_122);
nand U1670 (N_1670,In_1177,In_1832);
nor U1671 (N_1671,In_5,In_1874);
and U1672 (N_1672,In_667,In_374);
nand U1673 (N_1673,In_1267,In_1889);
xor U1674 (N_1674,In_183,In_1461);
and U1675 (N_1675,In_206,In_385);
nor U1676 (N_1676,In_935,In_1776);
nor U1677 (N_1677,In_1217,In_1005);
nand U1678 (N_1678,In_510,In_107);
xor U1679 (N_1679,In_568,In_1201);
nand U1680 (N_1680,In_1199,In_873);
nor U1681 (N_1681,In_1260,In_228);
or U1682 (N_1682,In_1058,In_582);
nand U1683 (N_1683,In_1452,In_792);
xor U1684 (N_1684,In_171,In_480);
and U1685 (N_1685,In_695,In_1346);
xor U1686 (N_1686,In_685,In_1648);
nand U1687 (N_1687,In_609,In_1011);
or U1688 (N_1688,In_982,In_1366);
nor U1689 (N_1689,In_113,In_1700);
nor U1690 (N_1690,In_1094,In_1386);
nand U1691 (N_1691,In_827,In_871);
nand U1692 (N_1692,In_1083,In_232);
or U1693 (N_1693,In_574,In_595);
nor U1694 (N_1694,In_1150,In_405);
nor U1695 (N_1695,In_15,In_179);
nor U1696 (N_1696,In_1827,In_197);
or U1697 (N_1697,In_1443,In_1331);
or U1698 (N_1698,In_83,In_221);
and U1699 (N_1699,In_1233,In_215);
nor U1700 (N_1700,In_1554,In_1760);
and U1701 (N_1701,In_339,In_535);
and U1702 (N_1702,In_1279,In_1692);
nand U1703 (N_1703,In_723,In_1776);
nor U1704 (N_1704,In_414,In_966);
or U1705 (N_1705,In_1302,In_101);
nand U1706 (N_1706,In_1550,In_1240);
nor U1707 (N_1707,In_1537,In_1411);
and U1708 (N_1708,In_635,In_1751);
nand U1709 (N_1709,In_1372,In_341);
or U1710 (N_1710,In_101,In_1501);
or U1711 (N_1711,In_357,In_1);
nor U1712 (N_1712,In_790,In_1439);
and U1713 (N_1713,In_1128,In_1446);
xnor U1714 (N_1714,In_758,In_977);
or U1715 (N_1715,In_1633,In_1924);
nand U1716 (N_1716,In_136,In_1988);
and U1717 (N_1717,In_1867,In_1230);
nor U1718 (N_1718,In_76,In_166);
nand U1719 (N_1719,In_945,In_769);
and U1720 (N_1720,In_1344,In_1500);
and U1721 (N_1721,In_1408,In_1929);
nor U1722 (N_1722,In_177,In_456);
and U1723 (N_1723,In_213,In_287);
nor U1724 (N_1724,In_1145,In_232);
and U1725 (N_1725,In_467,In_44);
or U1726 (N_1726,In_514,In_1646);
and U1727 (N_1727,In_939,In_643);
nand U1728 (N_1728,In_353,In_604);
nand U1729 (N_1729,In_1717,In_439);
nor U1730 (N_1730,In_820,In_858);
nor U1731 (N_1731,In_1827,In_310);
or U1732 (N_1732,In_792,In_59);
nor U1733 (N_1733,In_1258,In_1531);
nor U1734 (N_1734,In_1733,In_160);
nor U1735 (N_1735,In_1071,In_449);
or U1736 (N_1736,In_1693,In_1418);
nor U1737 (N_1737,In_929,In_97);
nor U1738 (N_1738,In_637,In_1808);
and U1739 (N_1739,In_976,In_1551);
and U1740 (N_1740,In_504,In_15);
and U1741 (N_1741,In_1000,In_242);
or U1742 (N_1742,In_1211,In_1490);
or U1743 (N_1743,In_1656,In_1230);
or U1744 (N_1744,In_405,In_669);
xnor U1745 (N_1745,In_1457,In_1715);
xnor U1746 (N_1746,In_943,In_1878);
or U1747 (N_1747,In_1472,In_870);
or U1748 (N_1748,In_85,In_876);
and U1749 (N_1749,In_380,In_1768);
xnor U1750 (N_1750,In_493,In_638);
nand U1751 (N_1751,In_1498,In_42);
xnor U1752 (N_1752,In_1228,In_1989);
nor U1753 (N_1753,In_1617,In_877);
and U1754 (N_1754,In_1426,In_306);
and U1755 (N_1755,In_86,In_1146);
nor U1756 (N_1756,In_1761,In_1891);
nand U1757 (N_1757,In_73,In_607);
and U1758 (N_1758,In_1988,In_574);
and U1759 (N_1759,In_1648,In_1009);
nand U1760 (N_1760,In_444,In_183);
or U1761 (N_1761,In_335,In_448);
nand U1762 (N_1762,In_810,In_1953);
or U1763 (N_1763,In_844,In_1554);
and U1764 (N_1764,In_523,In_1236);
and U1765 (N_1765,In_840,In_977);
or U1766 (N_1766,In_1737,In_801);
and U1767 (N_1767,In_1777,In_644);
xor U1768 (N_1768,In_905,In_1841);
or U1769 (N_1769,In_162,In_609);
nand U1770 (N_1770,In_691,In_959);
or U1771 (N_1771,In_1818,In_1158);
nand U1772 (N_1772,In_607,In_718);
and U1773 (N_1773,In_132,In_413);
xor U1774 (N_1774,In_461,In_119);
nand U1775 (N_1775,In_1284,In_273);
and U1776 (N_1776,In_1225,In_381);
and U1777 (N_1777,In_475,In_1109);
nand U1778 (N_1778,In_689,In_367);
or U1779 (N_1779,In_1239,In_1219);
or U1780 (N_1780,In_1518,In_935);
and U1781 (N_1781,In_1273,In_1461);
xnor U1782 (N_1782,In_373,In_333);
nor U1783 (N_1783,In_76,In_266);
xnor U1784 (N_1784,In_655,In_659);
and U1785 (N_1785,In_1515,In_945);
nand U1786 (N_1786,In_1565,In_1260);
nand U1787 (N_1787,In_1207,In_132);
nand U1788 (N_1788,In_225,In_1405);
nor U1789 (N_1789,In_945,In_122);
nor U1790 (N_1790,In_1389,In_1960);
and U1791 (N_1791,In_150,In_1784);
nand U1792 (N_1792,In_1041,In_1610);
nand U1793 (N_1793,In_1285,In_96);
or U1794 (N_1794,In_1369,In_1379);
nand U1795 (N_1795,In_1141,In_1206);
xor U1796 (N_1796,In_502,In_614);
nor U1797 (N_1797,In_1376,In_514);
and U1798 (N_1798,In_246,In_634);
and U1799 (N_1799,In_784,In_586);
nand U1800 (N_1800,In_1046,In_1249);
xnor U1801 (N_1801,In_540,In_1749);
or U1802 (N_1802,In_681,In_1340);
nor U1803 (N_1803,In_992,In_1169);
and U1804 (N_1804,In_94,In_1032);
nand U1805 (N_1805,In_377,In_1804);
or U1806 (N_1806,In_1937,In_671);
nand U1807 (N_1807,In_1866,In_1182);
nor U1808 (N_1808,In_415,In_210);
or U1809 (N_1809,In_1062,In_783);
or U1810 (N_1810,In_1016,In_772);
nand U1811 (N_1811,In_1407,In_1855);
or U1812 (N_1812,In_102,In_1969);
or U1813 (N_1813,In_1224,In_1556);
nand U1814 (N_1814,In_896,In_1267);
nand U1815 (N_1815,In_657,In_780);
nor U1816 (N_1816,In_1935,In_1115);
and U1817 (N_1817,In_1540,In_1951);
or U1818 (N_1818,In_1310,In_846);
nor U1819 (N_1819,In_1583,In_1);
or U1820 (N_1820,In_319,In_1305);
nand U1821 (N_1821,In_385,In_16);
or U1822 (N_1822,In_401,In_1519);
nand U1823 (N_1823,In_1091,In_58);
nand U1824 (N_1824,In_1054,In_1367);
nor U1825 (N_1825,In_716,In_1136);
and U1826 (N_1826,In_1991,In_1207);
and U1827 (N_1827,In_1961,In_1084);
nand U1828 (N_1828,In_1221,In_170);
xor U1829 (N_1829,In_504,In_1049);
nand U1830 (N_1830,In_1589,In_1630);
nand U1831 (N_1831,In_1416,In_355);
xor U1832 (N_1832,In_1756,In_1056);
nand U1833 (N_1833,In_559,In_987);
nand U1834 (N_1834,In_927,In_1530);
or U1835 (N_1835,In_933,In_1070);
or U1836 (N_1836,In_1967,In_1341);
nor U1837 (N_1837,In_88,In_1400);
nor U1838 (N_1838,In_941,In_1332);
nor U1839 (N_1839,In_1027,In_1808);
nand U1840 (N_1840,In_939,In_1520);
nand U1841 (N_1841,In_1310,In_175);
nor U1842 (N_1842,In_785,In_1461);
or U1843 (N_1843,In_876,In_1538);
and U1844 (N_1844,In_1136,In_1055);
or U1845 (N_1845,In_255,In_66);
nor U1846 (N_1846,In_326,In_1033);
nand U1847 (N_1847,In_1674,In_1367);
or U1848 (N_1848,In_329,In_579);
and U1849 (N_1849,In_733,In_845);
xor U1850 (N_1850,In_94,In_1731);
or U1851 (N_1851,In_548,In_1317);
nor U1852 (N_1852,In_212,In_823);
nand U1853 (N_1853,In_1771,In_765);
and U1854 (N_1854,In_1286,In_1395);
xor U1855 (N_1855,In_1053,In_798);
nor U1856 (N_1856,In_654,In_1872);
nand U1857 (N_1857,In_1505,In_1973);
nand U1858 (N_1858,In_1144,In_1451);
or U1859 (N_1859,In_1022,In_1255);
and U1860 (N_1860,In_1886,In_815);
xor U1861 (N_1861,In_1175,In_1863);
nand U1862 (N_1862,In_1905,In_1642);
xor U1863 (N_1863,In_454,In_1364);
nand U1864 (N_1864,In_338,In_1446);
or U1865 (N_1865,In_1375,In_1369);
and U1866 (N_1866,In_1707,In_1362);
nor U1867 (N_1867,In_611,In_71);
nor U1868 (N_1868,In_535,In_602);
and U1869 (N_1869,In_1997,In_258);
or U1870 (N_1870,In_1480,In_131);
or U1871 (N_1871,In_50,In_901);
nand U1872 (N_1872,In_792,In_1507);
nor U1873 (N_1873,In_367,In_762);
and U1874 (N_1874,In_453,In_829);
or U1875 (N_1875,In_1558,In_749);
or U1876 (N_1876,In_847,In_376);
nand U1877 (N_1877,In_596,In_1523);
and U1878 (N_1878,In_1883,In_1431);
nand U1879 (N_1879,In_62,In_57);
xor U1880 (N_1880,In_1272,In_1442);
xnor U1881 (N_1881,In_1625,In_459);
nand U1882 (N_1882,In_1344,In_51);
and U1883 (N_1883,In_567,In_458);
nor U1884 (N_1884,In_1739,In_1415);
nand U1885 (N_1885,In_827,In_763);
or U1886 (N_1886,In_826,In_724);
or U1887 (N_1887,In_1925,In_223);
nor U1888 (N_1888,In_1394,In_1883);
xor U1889 (N_1889,In_1671,In_1130);
nand U1890 (N_1890,In_282,In_875);
nor U1891 (N_1891,In_471,In_1759);
xnor U1892 (N_1892,In_59,In_1011);
nand U1893 (N_1893,In_1516,In_116);
nor U1894 (N_1894,In_128,In_127);
or U1895 (N_1895,In_460,In_1884);
xnor U1896 (N_1896,In_1877,In_599);
and U1897 (N_1897,In_1198,In_1604);
nor U1898 (N_1898,In_1580,In_1807);
nor U1899 (N_1899,In_1251,In_663);
nand U1900 (N_1900,In_1877,In_656);
nor U1901 (N_1901,In_536,In_1419);
nor U1902 (N_1902,In_388,In_479);
or U1903 (N_1903,In_709,In_58);
nand U1904 (N_1904,In_1446,In_1837);
or U1905 (N_1905,In_1560,In_229);
nor U1906 (N_1906,In_1266,In_1599);
nor U1907 (N_1907,In_1342,In_1012);
or U1908 (N_1908,In_175,In_1995);
nand U1909 (N_1909,In_1471,In_1486);
nand U1910 (N_1910,In_1991,In_1289);
and U1911 (N_1911,In_936,In_394);
or U1912 (N_1912,In_1968,In_569);
xor U1913 (N_1913,In_285,In_1599);
or U1914 (N_1914,In_149,In_1981);
or U1915 (N_1915,In_835,In_1148);
xor U1916 (N_1916,In_1176,In_1309);
xnor U1917 (N_1917,In_833,In_1904);
nand U1918 (N_1918,In_1870,In_1727);
nor U1919 (N_1919,In_1343,In_191);
or U1920 (N_1920,In_1676,In_831);
nor U1921 (N_1921,In_713,In_1569);
xnor U1922 (N_1922,In_297,In_928);
nor U1923 (N_1923,In_1861,In_138);
and U1924 (N_1924,In_71,In_106);
nand U1925 (N_1925,In_1304,In_1314);
or U1926 (N_1926,In_364,In_374);
or U1927 (N_1927,In_935,In_1991);
or U1928 (N_1928,In_1365,In_140);
nand U1929 (N_1929,In_1749,In_1332);
nor U1930 (N_1930,In_170,In_1315);
nor U1931 (N_1931,In_1781,In_1668);
nor U1932 (N_1932,In_1669,In_1108);
or U1933 (N_1933,In_1769,In_1140);
xor U1934 (N_1934,In_723,In_794);
nand U1935 (N_1935,In_1701,In_1194);
or U1936 (N_1936,In_833,In_239);
or U1937 (N_1937,In_41,In_1776);
and U1938 (N_1938,In_1284,In_730);
and U1939 (N_1939,In_1823,In_1314);
or U1940 (N_1940,In_448,In_1291);
or U1941 (N_1941,In_1502,In_1704);
nand U1942 (N_1942,In_1153,In_101);
xnor U1943 (N_1943,In_1836,In_228);
and U1944 (N_1944,In_124,In_1895);
xnor U1945 (N_1945,In_1210,In_892);
nand U1946 (N_1946,In_200,In_1117);
nor U1947 (N_1947,In_1142,In_1966);
or U1948 (N_1948,In_1539,In_71);
or U1949 (N_1949,In_1382,In_1669);
and U1950 (N_1950,In_807,In_506);
and U1951 (N_1951,In_1586,In_291);
nand U1952 (N_1952,In_1290,In_478);
or U1953 (N_1953,In_646,In_451);
nand U1954 (N_1954,In_1923,In_751);
nor U1955 (N_1955,In_1358,In_919);
nand U1956 (N_1956,In_1065,In_272);
nand U1957 (N_1957,In_215,In_1226);
or U1958 (N_1958,In_1549,In_1881);
xnor U1959 (N_1959,In_809,In_1850);
nor U1960 (N_1960,In_641,In_604);
nor U1961 (N_1961,In_842,In_1988);
xnor U1962 (N_1962,In_1544,In_596);
nor U1963 (N_1963,In_115,In_709);
nand U1964 (N_1964,In_345,In_1502);
nor U1965 (N_1965,In_381,In_1851);
nand U1966 (N_1966,In_1109,In_494);
nand U1967 (N_1967,In_915,In_230);
nand U1968 (N_1968,In_1149,In_1835);
nand U1969 (N_1969,In_21,In_1697);
and U1970 (N_1970,In_903,In_897);
nand U1971 (N_1971,In_1603,In_1859);
nor U1972 (N_1972,In_1991,In_1217);
nor U1973 (N_1973,In_580,In_470);
and U1974 (N_1974,In_881,In_1369);
nor U1975 (N_1975,In_1882,In_328);
nand U1976 (N_1976,In_1014,In_1617);
nand U1977 (N_1977,In_1854,In_1409);
or U1978 (N_1978,In_1816,In_730);
or U1979 (N_1979,In_410,In_1918);
and U1980 (N_1980,In_1401,In_1367);
nand U1981 (N_1981,In_813,In_1888);
nor U1982 (N_1982,In_423,In_805);
and U1983 (N_1983,In_624,In_349);
nand U1984 (N_1984,In_1787,In_490);
nand U1985 (N_1985,In_1718,In_628);
and U1986 (N_1986,In_661,In_645);
nor U1987 (N_1987,In_52,In_190);
and U1988 (N_1988,In_1444,In_511);
nand U1989 (N_1989,In_561,In_974);
and U1990 (N_1990,In_640,In_1349);
nor U1991 (N_1991,In_563,In_1781);
nand U1992 (N_1992,In_756,In_293);
nand U1993 (N_1993,In_1943,In_680);
or U1994 (N_1994,In_313,In_1525);
nor U1995 (N_1995,In_368,In_1816);
nor U1996 (N_1996,In_1076,In_1781);
nor U1997 (N_1997,In_1098,In_1070);
nand U1998 (N_1998,In_1800,In_1269);
nand U1999 (N_1999,In_817,In_893);
nor U2000 (N_2000,In_1510,In_923);
and U2001 (N_2001,In_1594,In_1636);
nor U2002 (N_2002,In_974,In_1458);
and U2003 (N_2003,In_1128,In_1159);
and U2004 (N_2004,In_1324,In_510);
nand U2005 (N_2005,In_1397,In_1413);
or U2006 (N_2006,In_1641,In_874);
nand U2007 (N_2007,In_299,In_1664);
or U2008 (N_2008,In_47,In_1248);
nand U2009 (N_2009,In_582,In_1715);
or U2010 (N_2010,In_233,In_694);
or U2011 (N_2011,In_965,In_854);
or U2012 (N_2012,In_587,In_1750);
or U2013 (N_2013,In_1624,In_1671);
or U2014 (N_2014,In_1336,In_938);
nor U2015 (N_2015,In_252,In_1808);
nand U2016 (N_2016,In_914,In_203);
and U2017 (N_2017,In_22,In_1028);
or U2018 (N_2018,In_385,In_1496);
and U2019 (N_2019,In_551,In_624);
nor U2020 (N_2020,In_1041,In_980);
and U2021 (N_2021,In_237,In_140);
and U2022 (N_2022,In_1382,In_1068);
and U2023 (N_2023,In_801,In_29);
nand U2024 (N_2024,In_1275,In_1709);
nor U2025 (N_2025,In_801,In_1210);
nand U2026 (N_2026,In_951,In_1208);
or U2027 (N_2027,In_864,In_116);
and U2028 (N_2028,In_894,In_1799);
nor U2029 (N_2029,In_1477,In_1485);
or U2030 (N_2030,In_1813,In_1263);
nand U2031 (N_2031,In_1935,In_1545);
and U2032 (N_2032,In_148,In_1010);
xnor U2033 (N_2033,In_1834,In_1597);
nor U2034 (N_2034,In_1272,In_491);
or U2035 (N_2035,In_893,In_470);
or U2036 (N_2036,In_1281,In_1944);
nor U2037 (N_2037,In_1145,In_371);
or U2038 (N_2038,In_1996,In_1091);
nand U2039 (N_2039,In_133,In_78);
nand U2040 (N_2040,In_1915,In_621);
and U2041 (N_2041,In_1585,In_1316);
or U2042 (N_2042,In_1197,In_1724);
and U2043 (N_2043,In_882,In_1667);
xor U2044 (N_2044,In_195,In_1060);
nand U2045 (N_2045,In_217,In_935);
or U2046 (N_2046,In_908,In_1092);
and U2047 (N_2047,In_342,In_1482);
or U2048 (N_2048,In_1130,In_568);
or U2049 (N_2049,In_56,In_145);
nand U2050 (N_2050,In_1187,In_614);
xnor U2051 (N_2051,In_1321,In_1113);
and U2052 (N_2052,In_1452,In_1163);
or U2053 (N_2053,In_1197,In_9);
nor U2054 (N_2054,In_1369,In_1790);
and U2055 (N_2055,In_1779,In_248);
xor U2056 (N_2056,In_1710,In_1576);
or U2057 (N_2057,In_1075,In_168);
nand U2058 (N_2058,In_129,In_957);
xnor U2059 (N_2059,In_624,In_1288);
xor U2060 (N_2060,In_588,In_191);
or U2061 (N_2061,In_1007,In_1643);
and U2062 (N_2062,In_1910,In_1508);
nand U2063 (N_2063,In_1153,In_376);
and U2064 (N_2064,In_167,In_650);
nor U2065 (N_2065,In_1254,In_642);
nand U2066 (N_2066,In_1727,In_1043);
nand U2067 (N_2067,In_1833,In_1078);
nand U2068 (N_2068,In_1864,In_1042);
xor U2069 (N_2069,In_1063,In_1794);
or U2070 (N_2070,In_1729,In_936);
xor U2071 (N_2071,In_124,In_1183);
and U2072 (N_2072,In_1648,In_795);
nor U2073 (N_2073,In_1175,In_161);
nand U2074 (N_2074,In_1563,In_248);
xor U2075 (N_2075,In_130,In_342);
xnor U2076 (N_2076,In_773,In_1287);
or U2077 (N_2077,In_431,In_1647);
and U2078 (N_2078,In_539,In_1647);
and U2079 (N_2079,In_1442,In_1469);
xor U2080 (N_2080,In_1046,In_856);
and U2081 (N_2081,In_1189,In_1114);
nand U2082 (N_2082,In_1935,In_576);
nor U2083 (N_2083,In_311,In_1720);
and U2084 (N_2084,In_1833,In_1018);
or U2085 (N_2085,In_957,In_608);
nand U2086 (N_2086,In_1673,In_315);
nand U2087 (N_2087,In_1075,In_949);
nor U2088 (N_2088,In_1624,In_1272);
nand U2089 (N_2089,In_255,In_20);
nand U2090 (N_2090,In_1780,In_1385);
nand U2091 (N_2091,In_1832,In_11);
xor U2092 (N_2092,In_33,In_1144);
or U2093 (N_2093,In_1986,In_1740);
nor U2094 (N_2094,In_1702,In_884);
nor U2095 (N_2095,In_1637,In_1922);
nand U2096 (N_2096,In_15,In_100);
or U2097 (N_2097,In_819,In_137);
xnor U2098 (N_2098,In_322,In_1949);
or U2099 (N_2099,In_1641,In_1136);
and U2100 (N_2100,In_1294,In_1825);
nor U2101 (N_2101,In_1801,In_625);
and U2102 (N_2102,In_1435,In_666);
xnor U2103 (N_2103,In_106,In_536);
nand U2104 (N_2104,In_1809,In_1633);
nor U2105 (N_2105,In_324,In_483);
nand U2106 (N_2106,In_87,In_763);
or U2107 (N_2107,In_578,In_1121);
and U2108 (N_2108,In_735,In_536);
nand U2109 (N_2109,In_429,In_1271);
nor U2110 (N_2110,In_619,In_1594);
nand U2111 (N_2111,In_8,In_1550);
xor U2112 (N_2112,In_526,In_609);
nand U2113 (N_2113,In_1124,In_1567);
or U2114 (N_2114,In_1002,In_1716);
nor U2115 (N_2115,In_1458,In_1134);
or U2116 (N_2116,In_116,In_1352);
xnor U2117 (N_2117,In_1704,In_236);
nand U2118 (N_2118,In_1665,In_1934);
or U2119 (N_2119,In_1130,In_347);
or U2120 (N_2120,In_1163,In_1419);
and U2121 (N_2121,In_130,In_564);
nor U2122 (N_2122,In_206,In_623);
and U2123 (N_2123,In_687,In_1720);
nand U2124 (N_2124,In_293,In_968);
and U2125 (N_2125,In_1716,In_942);
nor U2126 (N_2126,In_1874,In_945);
xor U2127 (N_2127,In_246,In_244);
and U2128 (N_2128,In_374,In_1468);
nand U2129 (N_2129,In_61,In_399);
xor U2130 (N_2130,In_526,In_892);
xnor U2131 (N_2131,In_1545,In_1733);
nor U2132 (N_2132,In_1572,In_1186);
or U2133 (N_2133,In_242,In_1053);
or U2134 (N_2134,In_1195,In_366);
nand U2135 (N_2135,In_220,In_1477);
nand U2136 (N_2136,In_1509,In_1983);
or U2137 (N_2137,In_1264,In_1685);
or U2138 (N_2138,In_1271,In_1919);
and U2139 (N_2139,In_1408,In_1679);
nor U2140 (N_2140,In_1745,In_471);
nor U2141 (N_2141,In_454,In_13);
or U2142 (N_2142,In_1852,In_1943);
nor U2143 (N_2143,In_788,In_274);
nor U2144 (N_2144,In_984,In_804);
or U2145 (N_2145,In_1637,In_400);
nand U2146 (N_2146,In_1635,In_1317);
nor U2147 (N_2147,In_1300,In_561);
or U2148 (N_2148,In_1023,In_1478);
or U2149 (N_2149,In_1746,In_1425);
xor U2150 (N_2150,In_541,In_306);
or U2151 (N_2151,In_497,In_731);
nand U2152 (N_2152,In_219,In_1049);
nor U2153 (N_2153,In_994,In_1812);
xor U2154 (N_2154,In_915,In_1234);
xor U2155 (N_2155,In_1888,In_883);
nor U2156 (N_2156,In_1129,In_259);
nor U2157 (N_2157,In_519,In_1442);
nand U2158 (N_2158,In_1339,In_992);
or U2159 (N_2159,In_355,In_1183);
nor U2160 (N_2160,In_65,In_464);
nor U2161 (N_2161,In_70,In_447);
xnor U2162 (N_2162,In_1686,In_602);
or U2163 (N_2163,In_365,In_1493);
or U2164 (N_2164,In_834,In_646);
xnor U2165 (N_2165,In_710,In_1785);
and U2166 (N_2166,In_478,In_1236);
nor U2167 (N_2167,In_81,In_1631);
or U2168 (N_2168,In_1090,In_516);
and U2169 (N_2169,In_681,In_504);
and U2170 (N_2170,In_1641,In_1837);
nand U2171 (N_2171,In_769,In_937);
or U2172 (N_2172,In_1882,In_939);
nand U2173 (N_2173,In_820,In_992);
nor U2174 (N_2174,In_1145,In_22);
nor U2175 (N_2175,In_1740,In_450);
nand U2176 (N_2176,In_965,In_1078);
or U2177 (N_2177,In_509,In_1747);
or U2178 (N_2178,In_1483,In_1192);
nand U2179 (N_2179,In_51,In_1707);
nand U2180 (N_2180,In_1577,In_392);
and U2181 (N_2181,In_1593,In_1544);
nand U2182 (N_2182,In_912,In_1956);
nor U2183 (N_2183,In_1631,In_70);
xor U2184 (N_2184,In_426,In_89);
nand U2185 (N_2185,In_1171,In_1336);
nand U2186 (N_2186,In_1006,In_164);
nand U2187 (N_2187,In_1543,In_923);
and U2188 (N_2188,In_1745,In_495);
or U2189 (N_2189,In_98,In_910);
or U2190 (N_2190,In_1153,In_1678);
nand U2191 (N_2191,In_1860,In_583);
xnor U2192 (N_2192,In_66,In_131);
nand U2193 (N_2193,In_71,In_10);
nand U2194 (N_2194,In_1623,In_1122);
xnor U2195 (N_2195,In_707,In_325);
and U2196 (N_2196,In_1923,In_351);
nand U2197 (N_2197,In_1224,In_913);
nor U2198 (N_2198,In_588,In_1230);
and U2199 (N_2199,In_1998,In_1930);
nand U2200 (N_2200,In_1882,In_821);
or U2201 (N_2201,In_1799,In_889);
nor U2202 (N_2202,In_538,In_1702);
or U2203 (N_2203,In_627,In_1853);
nor U2204 (N_2204,In_1341,In_1185);
and U2205 (N_2205,In_156,In_918);
nor U2206 (N_2206,In_281,In_606);
nand U2207 (N_2207,In_334,In_370);
nand U2208 (N_2208,In_109,In_1367);
nor U2209 (N_2209,In_1339,In_1940);
nor U2210 (N_2210,In_49,In_1240);
and U2211 (N_2211,In_1648,In_1115);
xor U2212 (N_2212,In_559,In_1850);
and U2213 (N_2213,In_1698,In_608);
nand U2214 (N_2214,In_366,In_1513);
or U2215 (N_2215,In_1219,In_1736);
and U2216 (N_2216,In_541,In_169);
or U2217 (N_2217,In_942,In_1795);
xor U2218 (N_2218,In_820,In_318);
and U2219 (N_2219,In_370,In_199);
or U2220 (N_2220,In_986,In_1087);
or U2221 (N_2221,In_12,In_452);
and U2222 (N_2222,In_426,In_1077);
nand U2223 (N_2223,In_1649,In_1619);
nor U2224 (N_2224,In_601,In_481);
and U2225 (N_2225,In_771,In_855);
or U2226 (N_2226,In_302,In_234);
nand U2227 (N_2227,In_1663,In_1056);
nand U2228 (N_2228,In_176,In_1455);
nor U2229 (N_2229,In_1216,In_752);
xor U2230 (N_2230,In_1624,In_115);
xor U2231 (N_2231,In_947,In_1205);
nand U2232 (N_2232,In_1375,In_1889);
or U2233 (N_2233,In_1340,In_1519);
or U2234 (N_2234,In_1992,In_729);
or U2235 (N_2235,In_1162,In_757);
xor U2236 (N_2236,In_1894,In_1820);
nand U2237 (N_2237,In_569,In_623);
nand U2238 (N_2238,In_1129,In_1276);
nor U2239 (N_2239,In_797,In_1138);
nor U2240 (N_2240,In_4,In_414);
or U2241 (N_2241,In_1558,In_1402);
nor U2242 (N_2242,In_1328,In_616);
nor U2243 (N_2243,In_1488,In_1387);
nor U2244 (N_2244,In_1737,In_1719);
nand U2245 (N_2245,In_1077,In_1926);
nand U2246 (N_2246,In_1217,In_929);
nor U2247 (N_2247,In_707,In_332);
nor U2248 (N_2248,In_411,In_311);
and U2249 (N_2249,In_528,In_1782);
xor U2250 (N_2250,In_1843,In_1734);
or U2251 (N_2251,In_1972,In_1767);
and U2252 (N_2252,In_209,In_1490);
nor U2253 (N_2253,In_305,In_679);
nand U2254 (N_2254,In_1034,In_147);
and U2255 (N_2255,In_243,In_1610);
xor U2256 (N_2256,In_381,In_1179);
or U2257 (N_2257,In_1213,In_415);
and U2258 (N_2258,In_1254,In_842);
nor U2259 (N_2259,In_259,In_1445);
nor U2260 (N_2260,In_1019,In_797);
and U2261 (N_2261,In_196,In_1456);
xnor U2262 (N_2262,In_632,In_1507);
nor U2263 (N_2263,In_834,In_419);
xor U2264 (N_2264,In_1537,In_125);
nand U2265 (N_2265,In_1150,In_450);
xor U2266 (N_2266,In_267,In_171);
xnor U2267 (N_2267,In_1013,In_140);
and U2268 (N_2268,In_1812,In_235);
or U2269 (N_2269,In_1712,In_806);
or U2270 (N_2270,In_450,In_1623);
nand U2271 (N_2271,In_269,In_28);
or U2272 (N_2272,In_1278,In_1670);
and U2273 (N_2273,In_658,In_1315);
or U2274 (N_2274,In_263,In_1564);
and U2275 (N_2275,In_1779,In_1120);
nand U2276 (N_2276,In_1881,In_1087);
or U2277 (N_2277,In_682,In_422);
and U2278 (N_2278,In_943,In_1909);
nor U2279 (N_2279,In_964,In_1213);
xnor U2280 (N_2280,In_1271,In_1314);
nand U2281 (N_2281,In_940,In_325);
and U2282 (N_2282,In_157,In_1215);
and U2283 (N_2283,In_1928,In_1142);
nand U2284 (N_2284,In_132,In_1628);
or U2285 (N_2285,In_252,In_1221);
or U2286 (N_2286,In_1379,In_1629);
nand U2287 (N_2287,In_1148,In_522);
and U2288 (N_2288,In_780,In_639);
nand U2289 (N_2289,In_949,In_1016);
nor U2290 (N_2290,In_323,In_705);
nor U2291 (N_2291,In_634,In_513);
xnor U2292 (N_2292,In_252,In_1314);
nand U2293 (N_2293,In_1960,In_448);
and U2294 (N_2294,In_139,In_1992);
xnor U2295 (N_2295,In_1275,In_316);
or U2296 (N_2296,In_1509,In_26);
and U2297 (N_2297,In_681,In_1040);
nand U2298 (N_2298,In_814,In_870);
nor U2299 (N_2299,In_751,In_119);
nor U2300 (N_2300,In_215,In_920);
or U2301 (N_2301,In_891,In_1840);
and U2302 (N_2302,In_1447,In_1067);
and U2303 (N_2303,In_1357,In_639);
or U2304 (N_2304,In_1946,In_1591);
or U2305 (N_2305,In_845,In_1312);
nor U2306 (N_2306,In_1297,In_190);
and U2307 (N_2307,In_1283,In_315);
and U2308 (N_2308,In_1887,In_582);
nand U2309 (N_2309,In_478,In_273);
and U2310 (N_2310,In_1408,In_1853);
and U2311 (N_2311,In_652,In_153);
xor U2312 (N_2312,In_1422,In_782);
or U2313 (N_2313,In_1342,In_1974);
xnor U2314 (N_2314,In_548,In_1540);
or U2315 (N_2315,In_1777,In_1306);
and U2316 (N_2316,In_1435,In_1309);
nand U2317 (N_2317,In_440,In_205);
xor U2318 (N_2318,In_841,In_506);
or U2319 (N_2319,In_1988,In_1422);
xnor U2320 (N_2320,In_1738,In_880);
and U2321 (N_2321,In_1121,In_1142);
or U2322 (N_2322,In_516,In_165);
and U2323 (N_2323,In_884,In_822);
or U2324 (N_2324,In_255,In_368);
nand U2325 (N_2325,In_1342,In_1077);
or U2326 (N_2326,In_1629,In_356);
and U2327 (N_2327,In_1351,In_33);
and U2328 (N_2328,In_637,In_395);
nand U2329 (N_2329,In_1610,In_501);
and U2330 (N_2330,In_1811,In_1691);
nor U2331 (N_2331,In_1264,In_199);
nor U2332 (N_2332,In_133,In_1873);
and U2333 (N_2333,In_1281,In_1783);
nor U2334 (N_2334,In_593,In_1305);
nand U2335 (N_2335,In_1214,In_1773);
or U2336 (N_2336,In_708,In_1470);
and U2337 (N_2337,In_225,In_246);
nor U2338 (N_2338,In_674,In_708);
or U2339 (N_2339,In_1857,In_364);
nand U2340 (N_2340,In_1451,In_186);
nor U2341 (N_2341,In_1146,In_1114);
nor U2342 (N_2342,In_1368,In_1596);
or U2343 (N_2343,In_565,In_1898);
nor U2344 (N_2344,In_694,In_1712);
or U2345 (N_2345,In_1896,In_1229);
and U2346 (N_2346,In_954,In_825);
and U2347 (N_2347,In_1996,In_677);
nor U2348 (N_2348,In_969,In_1541);
nor U2349 (N_2349,In_1422,In_1258);
nor U2350 (N_2350,In_1392,In_163);
or U2351 (N_2351,In_66,In_497);
and U2352 (N_2352,In_251,In_1543);
and U2353 (N_2353,In_175,In_1317);
nor U2354 (N_2354,In_124,In_765);
nand U2355 (N_2355,In_83,In_1091);
nor U2356 (N_2356,In_1326,In_70);
and U2357 (N_2357,In_178,In_1337);
or U2358 (N_2358,In_33,In_874);
nor U2359 (N_2359,In_353,In_540);
and U2360 (N_2360,In_1141,In_716);
nor U2361 (N_2361,In_1170,In_36);
or U2362 (N_2362,In_820,In_640);
and U2363 (N_2363,In_973,In_1000);
nor U2364 (N_2364,In_1909,In_413);
nand U2365 (N_2365,In_551,In_423);
nand U2366 (N_2366,In_455,In_413);
nor U2367 (N_2367,In_1439,In_620);
nand U2368 (N_2368,In_869,In_1165);
and U2369 (N_2369,In_519,In_1971);
or U2370 (N_2370,In_145,In_344);
nand U2371 (N_2371,In_807,In_310);
or U2372 (N_2372,In_199,In_586);
xnor U2373 (N_2373,In_735,In_413);
and U2374 (N_2374,In_1230,In_1101);
nor U2375 (N_2375,In_1978,In_1727);
nor U2376 (N_2376,In_1896,In_1673);
and U2377 (N_2377,In_73,In_222);
or U2378 (N_2378,In_285,In_1973);
xor U2379 (N_2379,In_792,In_1810);
nor U2380 (N_2380,In_1240,In_113);
nor U2381 (N_2381,In_1272,In_261);
nor U2382 (N_2382,In_1884,In_571);
nand U2383 (N_2383,In_1194,In_797);
or U2384 (N_2384,In_429,In_146);
xor U2385 (N_2385,In_29,In_161);
and U2386 (N_2386,In_1655,In_526);
or U2387 (N_2387,In_1821,In_142);
nand U2388 (N_2388,In_822,In_1091);
nand U2389 (N_2389,In_1631,In_46);
or U2390 (N_2390,In_792,In_38);
nor U2391 (N_2391,In_457,In_1474);
nand U2392 (N_2392,In_800,In_1012);
or U2393 (N_2393,In_1934,In_899);
nand U2394 (N_2394,In_1966,In_543);
nor U2395 (N_2395,In_652,In_1115);
xnor U2396 (N_2396,In_816,In_1411);
nor U2397 (N_2397,In_1708,In_1458);
or U2398 (N_2398,In_1648,In_1546);
and U2399 (N_2399,In_1958,In_1949);
nor U2400 (N_2400,In_476,In_815);
and U2401 (N_2401,In_1896,In_1675);
and U2402 (N_2402,In_1074,In_1183);
nor U2403 (N_2403,In_595,In_947);
and U2404 (N_2404,In_1234,In_1799);
nor U2405 (N_2405,In_93,In_1952);
nor U2406 (N_2406,In_1999,In_1250);
nand U2407 (N_2407,In_1935,In_959);
and U2408 (N_2408,In_1027,In_1280);
nor U2409 (N_2409,In_1189,In_1178);
nor U2410 (N_2410,In_1712,In_1197);
and U2411 (N_2411,In_501,In_1364);
xor U2412 (N_2412,In_608,In_1623);
and U2413 (N_2413,In_294,In_550);
or U2414 (N_2414,In_62,In_1741);
or U2415 (N_2415,In_1445,In_1914);
or U2416 (N_2416,In_1723,In_334);
nand U2417 (N_2417,In_1047,In_1781);
or U2418 (N_2418,In_963,In_2);
or U2419 (N_2419,In_1386,In_1133);
and U2420 (N_2420,In_1676,In_1817);
or U2421 (N_2421,In_604,In_1095);
and U2422 (N_2422,In_596,In_1607);
nand U2423 (N_2423,In_1376,In_938);
nand U2424 (N_2424,In_1457,In_584);
and U2425 (N_2425,In_577,In_1733);
nand U2426 (N_2426,In_241,In_1883);
nand U2427 (N_2427,In_487,In_540);
and U2428 (N_2428,In_43,In_210);
or U2429 (N_2429,In_659,In_1996);
nor U2430 (N_2430,In_274,In_1283);
nor U2431 (N_2431,In_454,In_1380);
nor U2432 (N_2432,In_1141,In_1879);
nand U2433 (N_2433,In_1860,In_723);
nor U2434 (N_2434,In_1417,In_1067);
or U2435 (N_2435,In_1386,In_628);
xnor U2436 (N_2436,In_932,In_1773);
xor U2437 (N_2437,In_1358,In_935);
or U2438 (N_2438,In_1166,In_1410);
nor U2439 (N_2439,In_1149,In_885);
and U2440 (N_2440,In_333,In_1240);
or U2441 (N_2441,In_807,In_1415);
nand U2442 (N_2442,In_752,In_1978);
nand U2443 (N_2443,In_654,In_1260);
xor U2444 (N_2444,In_800,In_1627);
and U2445 (N_2445,In_247,In_235);
nor U2446 (N_2446,In_371,In_179);
nand U2447 (N_2447,In_548,In_240);
nor U2448 (N_2448,In_487,In_679);
or U2449 (N_2449,In_1566,In_1759);
nand U2450 (N_2450,In_77,In_156);
or U2451 (N_2451,In_661,In_1111);
and U2452 (N_2452,In_1297,In_1860);
nand U2453 (N_2453,In_104,In_920);
nand U2454 (N_2454,In_305,In_1968);
and U2455 (N_2455,In_1745,In_991);
and U2456 (N_2456,In_1452,In_1270);
and U2457 (N_2457,In_110,In_402);
nand U2458 (N_2458,In_326,In_549);
nand U2459 (N_2459,In_982,In_1346);
nand U2460 (N_2460,In_1871,In_501);
nor U2461 (N_2461,In_26,In_19);
or U2462 (N_2462,In_62,In_1551);
nand U2463 (N_2463,In_983,In_284);
or U2464 (N_2464,In_1066,In_1975);
nand U2465 (N_2465,In_1195,In_1833);
xor U2466 (N_2466,In_525,In_647);
or U2467 (N_2467,In_269,In_1423);
nand U2468 (N_2468,In_614,In_135);
or U2469 (N_2469,In_729,In_1241);
nor U2470 (N_2470,In_530,In_1935);
nor U2471 (N_2471,In_1747,In_640);
nor U2472 (N_2472,In_1479,In_261);
nor U2473 (N_2473,In_1858,In_359);
nand U2474 (N_2474,In_1579,In_561);
or U2475 (N_2475,In_984,In_1518);
or U2476 (N_2476,In_497,In_1249);
nor U2477 (N_2477,In_1,In_125);
nor U2478 (N_2478,In_675,In_1560);
nor U2479 (N_2479,In_896,In_485);
and U2480 (N_2480,In_699,In_249);
or U2481 (N_2481,In_780,In_191);
and U2482 (N_2482,In_1739,In_823);
nand U2483 (N_2483,In_1189,In_16);
nand U2484 (N_2484,In_1451,In_1367);
nand U2485 (N_2485,In_604,In_670);
or U2486 (N_2486,In_347,In_607);
or U2487 (N_2487,In_511,In_65);
nor U2488 (N_2488,In_581,In_1208);
nor U2489 (N_2489,In_51,In_1141);
nor U2490 (N_2490,In_548,In_1813);
nand U2491 (N_2491,In_993,In_864);
nand U2492 (N_2492,In_619,In_888);
or U2493 (N_2493,In_164,In_222);
and U2494 (N_2494,In_1299,In_1205);
nand U2495 (N_2495,In_624,In_1515);
xor U2496 (N_2496,In_364,In_1778);
nor U2497 (N_2497,In_906,In_1670);
nor U2498 (N_2498,In_1175,In_1454);
or U2499 (N_2499,In_349,In_10);
xnor U2500 (N_2500,In_1185,In_1099);
nor U2501 (N_2501,In_1447,In_901);
nand U2502 (N_2502,In_270,In_1825);
nand U2503 (N_2503,In_162,In_1605);
and U2504 (N_2504,In_1151,In_1816);
nor U2505 (N_2505,In_1025,In_1193);
or U2506 (N_2506,In_1030,In_693);
and U2507 (N_2507,In_1415,In_66);
nor U2508 (N_2508,In_250,In_347);
or U2509 (N_2509,In_1757,In_565);
nor U2510 (N_2510,In_35,In_564);
nand U2511 (N_2511,In_815,In_1354);
nand U2512 (N_2512,In_1137,In_1639);
nor U2513 (N_2513,In_938,In_230);
xor U2514 (N_2514,In_472,In_1145);
or U2515 (N_2515,In_485,In_12);
and U2516 (N_2516,In_1474,In_1102);
or U2517 (N_2517,In_1265,In_1648);
and U2518 (N_2518,In_1726,In_1569);
nor U2519 (N_2519,In_986,In_1682);
and U2520 (N_2520,In_384,In_407);
or U2521 (N_2521,In_1180,In_751);
nor U2522 (N_2522,In_1416,In_556);
or U2523 (N_2523,In_1852,In_1297);
and U2524 (N_2524,In_1776,In_1572);
or U2525 (N_2525,In_899,In_435);
nor U2526 (N_2526,In_1545,In_175);
and U2527 (N_2527,In_946,In_1908);
or U2528 (N_2528,In_308,In_729);
and U2529 (N_2529,In_1398,In_151);
and U2530 (N_2530,In_1719,In_1493);
or U2531 (N_2531,In_962,In_1205);
nor U2532 (N_2532,In_887,In_1429);
nor U2533 (N_2533,In_1290,In_1427);
or U2534 (N_2534,In_982,In_40);
or U2535 (N_2535,In_152,In_1307);
xnor U2536 (N_2536,In_1075,In_1252);
nor U2537 (N_2537,In_1048,In_163);
nand U2538 (N_2538,In_1146,In_1289);
nor U2539 (N_2539,In_110,In_1386);
or U2540 (N_2540,In_1341,In_674);
or U2541 (N_2541,In_289,In_322);
nor U2542 (N_2542,In_1829,In_1700);
and U2543 (N_2543,In_1768,In_668);
nor U2544 (N_2544,In_1317,In_1637);
xor U2545 (N_2545,In_1076,In_1197);
nor U2546 (N_2546,In_1310,In_1184);
or U2547 (N_2547,In_1401,In_193);
and U2548 (N_2548,In_1112,In_1684);
nor U2549 (N_2549,In_1335,In_1566);
nor U2550 (N_2550,In_854,In_1606);
and U2551 (N_2551,In_168,In_1891);
nand U2552 (N_2552,In_1874,In_1698);
nand U2553 (N_2553,In_1281,In_1250);
or U2554 (N_2554,In_365,In_784);
and U2555 (N_2555,In_1720,In_1959);
nor U2556 (N_2556,In_1303,In_1727);
or U2557 (N_2557,In_795,In_141);
nor U2558 (N_2558,In_262,In_1000);
and U2559 (N_2559,In_581,In_415);
nand U2560 (N_2560,In_238,In_737);
nand U2561 (N_2561,In_1765,In_716);
nor U2562 (N_2562,In_108,In_1893);
nand U2563 (N_2563,In_1603,In_164);
and U2564 (N_2564,In_1955,In_1483);
nor U2565 (N_2565,In_1394,In_976);
nand U2566 (N_2566,In_934,In_1775);
nand U2567 (N_2567,In_883,In_1040);
or U2568 (N_2568,In_394,In_812);
xnor U2569 (N_2569,In_1276,In_258);
nand U2570 (N_2570,In_179,In_24);
or U2571 (N_2571,In_800,In_40);
nand U2572 (N_2572,In_420,In_1410);
nand U2573 (N_2573,In_1244,In_1639);
or U2574 (N_2574,In_1652,In_895);
or U2575 (N_2575,In_1555,In_1260);
nand U2576 (N_2576,In_1792,In_1870);
nand U2577 (N_2577,In_1402,In_1435);
nor U2578 (N_2578,In_721,In_295);
or U2579 (N_2579,In_1452,In_468);
nand U2580 (N_2580,In_662,In_1094);
and U2581 (N_2581,In_1839,In_1763);
or U2582 (N_2582,In_1354,In_280);
or U2583 (N_2583,In_1749,In_1815);
or U2584 (N_2584,In_1796,In_1238);
nand U2585 (N_2585,In_564,In_1443);
nand U2586 (N_2586,In_1856,In_169);
and U2587 (N_2587,In_1505,In_1681);
nand U2588 (N_2588,In_1608,In_1556);
and U2589 (N_2589,In_1608,In_1244);
nand U2590 (N_2590,In_174,In_1279);
xor U2591 (N_2591,In_1027,In_635);
nand U2592 (N_2592,In_1868,In_720);
xor U2593 (N_2593,In_1586,In_80);
nor U2594 (N_2594,In_1639,In_1399);
or U2595 (N_2595,In_1111,In_1322);
nor U2596 (N_2596,In_1999,In_164);
and U2597 (N_2597,In_728,In_1489);
and U2598 (N_2598,In_1486,In_339);
nand U2599 (N_2599,In_172,In_1157);
nand U2600 (N_2600,In_1801,In_553);
nor U2601 (N_2601,In_1459,In_1444);
nor U2602 (N_2602,In_303,In_1767);
nand U2603 (N_2603,In_1947,In_130);
and U2604 (N_2604,In_182,In_1534);
nor U2605 (N_2605,In_86,In_316);
and U2606 (N_2606,In_283,In_1166);
nor U2607 (N_2607,In_1943,In_862);
nor U2608 (N_2608,In_1337,In_416);
and U2609 (N_2609,In_1370,In_1832);
or U2610 (N_2610,In_1153,In_1503);
or U2611 (N_2611,In_367,In_32);
or U2612 (N_2612,In_1567,In_275);
or U2613 (N_2613,In_1815,In_1089);
xor U2614 (N_2614,In_185,In_612);
and U2615 (N_2615,In_91,In_1743);
nor U2616 (N_2616,In_1704,In_1867);
xnor U2617 (N_2617,In_1609,In_1186);
and U2618 (N_2618,In_898,In_1822);
and U2619 (N_2619,In_1315,In_146);
or U2620 (N_2620,In_361,In_601);
nand U2621 (N_2621,In_91,In_663);
or U2622 (N_2622,In_710,In_1289);
or U2623 (N_2623,In_1827,In_1690);
nand U2624 (N_2624,In_1813,In_1049);
nor U2625 (N_2625,In_1487,In_1844);
nor U2626 (N_2626,In_843,In_1705);
or U2627 (N_2627,In_1675,In_1900);
or U2628 (N_2628,In_1262,In_700);
nor U2629 (N_2629,In_124,In_468);
xnor U2630 (N_2630,In_1988,In_514);
nor U2631 (N_2631,In_1715,In_1821);
or U2632 (N_2632,In_533,In_1109);
nor U2633 (N_2633,In_291,In_1857);
or U2634 (N_2634,In_1616,In_176);
and U2635 (N_2635,In_1294,In_979);
or U2636 (N_2636,In_344,In_1962);
nor U2637 (N_2637,In_609,In_600);
nand U2638 (N_2638,In_1593,In_1095);
and U2639 (N_2639,In_820,In_1121);
nor U2640 (N_2640,In_653,In_1252);
and U2641 (N_2641,In_787,In_937);
or U2642 (N_2642,In_1910,In_364);
or U2643 (N_2643,In_797,In_247);
or U2644 (N_2644,In_1853,In_1877);
nand U2645 (N_2645,In_1551,In_1673);
or U2646 (N_2646,In_112,In_1396);
nand U2647 (N_2647,In_478,In_1225);
nand U2648 (N_2648,In_1257,In_1563);
or U2649 (N_2649,In_792,In_1733);
nand U2650 (N_2650,In_30,In_759);
xnor U2651 (N_2651,In_1974,In_1688);
nand U2652 (N_2652,In_246,In_1872);
nor U2653 (N_2653,In_1956,In_1336);
nor U2654 (N_2654,In_1539,In_234);
xnor U2655 (N_2655,In_637,In_373);
nor U2656 (N_2656,In_963,In_1062);
and U2657 (N_2657,In_1617,In_1084);
and U2658 (N_2658,In_220,In_620);
nor U2659 (N_2659,In_1373,In_1569);
and U2660 (N_2660,In_623,In_700);
nand U2661 (N_2661,In_1795,In_1209);
or U2662 (N_2662,In_1271,In_1378);
nand U2663 (N_2663,In_1925,In_1933);
and U2664 (N_2664,In_296,In_1517);
and U2665 (N_2665,In_1555,In_455);
nor U2666 (N_2666,In_1055,In_526);
nor U2667 (N_2667,In_533,In_683);
and U2668 (N_2668,In_930,In_382);
and U2669 (N_2669,In_1649,In_1310);
or U2670 (N_2670,In_1649,In_1593);
nand U2671 (N_2671,In_738,In_1122);
nand U2672 (N_2672,In_1640,In_887);
nand U2673 (N_2673,In_1637,In_324);
xor U2674 (N_2674,In_1192,In_101);
or U2675 (N_2675,In_493,In_128);
nor U2676 (N_2676,In_1674,In_832);
and U2677 (N_2677,In_1542,In_1273);
xnor U2678 (N_2678,In_1917,In_1422);
and U2679 (N_2679,In_522,In_887);
nand U2680 (N_2680,In_199,In_866);
nor U2681 (N_2681,In_435,In_113);
nand U2682 (N_2682,In_492,In_944);
nor U2683 (N_2683,In_177,In_1910);
and U2684 (N_2684,In_1633,In_1979);
and U2685 (N_2685,In_1321,In_56);
nor U2686 (N_2686,In_1568,In_789);
nand U2687 (N_2687,In_1014,In_1427);
nand U2688 (N_2688,In_414,In_1261);
xnor U2689 (N_2689,In_365,In_475);
and U2690 (N_2690,In_478,In_707);
nor U2691 (N_2691,In_544,In_1498);
nand U2692 (N_2692,In_910,In_1251);
nand U2693 (N_2693,In_538,In_253);
nand U2694 (N_2694,In_1812,In_1660);
nor U2695 (N_2695,In_1879,In_516);
xor U2696 (N_2696,In_1752,In_1567);
nand U2697 (N_2697,In_1873,In_1784);
nand U2698 (N_2698,In_383,In_131);
xnor U2699 (N_2699,In_519,In_1047);
nand U2700 (N_2700,In_112,In_530);
nand U2701 (N_2701,In_1759,In_1400);
and U2702 (N_2702,In_1660,In_1056);
nor U2703 (N_2703,In_1909,In_1319);
and U2704 (N_2704,In_271,In_835);
nor U2705 (N_2705,In_1966,In_36);
and U2706 (N_2706,In_1757,In_1220);
nand U2707 (N_2707,In_860,In_1002);
and U2708 (N_2708,In_1750,In_787);
and U2709 (N_2709,In_1820,In_8);
nand U2710 (N_2710,In_630,In_1625);
and U2711 (N_2711,In_331,In_1872);
nor U2712 (N_2712,In_664,In_217);
and U2713 (N_2713,In_1392,In_1385);
nor U2714 (N_2714,In_814,In_1367);
xnor U2715 (N_2715,In_981,In_1584);
nand U2716 (N_2716,In_1502,In_0);
nand U2717 (N_2717,In_253,In_49);
and U2718 (N_2718,In_431,In_993);
nand U2719 (N_2719,In_1288,In_1410);
xor U2720 (N_2720,In_525,In_1663);
nand U2721 (N_2721,In_720,In_303);
or U2722 (N_2722,In_336,In_830);
nand U2723 (N_2723,In_1734,In_772);
nor U2724 (N_2724,In_1362,In_1930);
or U2725 (N_2725,In_146,In_385);
or U2726 (N_2726,In_1380,In_1395);
nand U2727 (N_2727,In_455,In_998);
nor U2728 (N_2728,In_1985,In_61);
and U2729 (N_2729,In_630,In_1448);
nand U2730 (N_2730,In_1091,In_1473);
or U2731 (N_2731,In_215,In_470);
and U2732 (N_2732,In_705,In_1704);
or U2733 (N_2733,In_216,In_670);
xor U2734 (N_2734,In_1213,In_1988);
nand U2735 (N_2735,In_543,In_944);
and U2736 (N_2736,In_26,In_1055);
and U2737 (N_2737,In_777,In_1574);
nor U2738 (N_2738,In_441,In_882);
nor U2739 (N_2739,In_1213,In_1944);
and U2740 (N_2740,In_273,In_1455);
or U2741 (N_2741,In_1507,In_1517);
and U2742 (N_2742,In_1203,In_1293);
nor U2743 (N_2743,In_1718,In_1372);
or U2744 (N_2744,In_1308,In_909);
nor U2745 (N_2745,In_38,In_1510);
and U2746 (N_2746,In_1556,In_177);
nand U2747 (N_2747,In_714,In_699);
nand U2748 (N_2748,In_1383,In_1956);
nand U2749 (N_2749,In_167,In_612);
nor U2750 (N_2750,In_1325,In_1487);
nor U2751 (N_2751,In_309,In_1634);
nor U2752 (N_2752,In_920,In_1301);
nor U2753 (N_2753,In_358,In_1249);
nand U2754 (N_2754,In_969,In_1151);
and U2755 (N_2755,In_1486,In_644);
nand U2756 (N_2756,In_1609,In_1997);
nor U2757 (N_2757,In_1917,In_1530);
and U2758 (N_2758,In_1849,In_1321);
and U2759 (N_2759,In_1763,In_1788);
or U2760 (N_2760,In_543,In_1241);
or U2761 (N_2761,In_437,In_1870);
or U2762 (N_2762,In_779,In_409);
nand U2763 (N_2763,In_978,In_1203);
and U2764 (N_2764,In_46,In_1456);
xnor U2765 (N_2765,In_760,In_1640);
nand U2766 (N_2766,In_1220,In_1674);
and U2767 (N_2767,In_472,In_1035);
nor U2768 (N_2768,In_444,In_1487);
and U2769 (N_2769,In_1621,In_1261);
or U2770 (N_2770,In_1542,In_285);
or U2771 (N_2771,In_102,In_311);
or U2772 (N_2772,In_1959,In_660);
or U2773 (N_2773,In_1374,In_1152);
nand U2774 (N_2774,In_252,In_1447);
nor U2775 (N_2775,In_928,In_181);
or U2776 (N_2776,In_1180,In_280);
or U2777 (N_2777,In_179,In_1582);
nand U2778 (N_2778,In_1039,In_500);
and U2779 (N_2779,In_380,In_590);
or U2780 (N_2780,In_432,In_271);
and U2781 (N_2781,In_311,In_1279);
or U2782 (N_2782,In_837,In_348);
nor U2783 (N_2783,In_1363,In_385);
or U2784 (N_2784,In_298,In_955);
or U2785 (N_2785,In_318,In_927);
nand U2786 (N_2786,In_923,In_1459);
nand U2787 (N_2787,In_1664,In_1636);
or U2788 (N_2788,In_237,In_1408);
and U2789 (N_2789,In_1204,In_360);
xnor U2790 (N_2790,In_590,In_749);
nor U2791 (N_2791,In_1391,In_1932);
nand U2792 (N_2792,In_1342,In_876);
or U2793 (N_2793,In_242,In_1482);
nor U2794 (N_2794,In_1914,In_986);
xnor U2795 (N_2795,In_922,In_527);
or U2796 (N_2796,In_1502,In_1984);
xnor U2797 (N_2797,In_324,In_1484);
or U2798 (N_2798,In_67,In_484);
nand U2799 (N_2799,In_123,In_256);
or U2800 (N_2800,In_16,In_1327);
or U2801 (N_2801,In_1950,In_1419);
xor U2802 (N_2802,In_1165,In_1698);
and U2803 (N_2803,In_775,In_1107);
nor U2804 (N_2804,In_1223,In_284);
or U2805 (N_2805,In_475,In_1460);
and U2806 (N_2806,In_883,In_529);
nor U2807 (N_2807,In_847,In_137);
nor U2808 (N_2808,In_1281,In_1071);
or U2809 (N_2809,In_1176,In_325);
and U2810 (N_2810,In_1990,In_1367);
and U2811 (N_2811,In_1192,In_27);
and U2812 (N_2812,In_881,In_1044);
or U2813 (N_2813,In_1615,In_1830);
and U2814 (N_2814,In_23,In_1319);
or U2815 (N_2815,In_489,In_1238);
nor U2816 (N_2816,In_603,In_1266);
nand U2817 (N_2817,In_1870,In_1600);
nand U2818 (N_2818,In_673,In_922);
or U2819 (N_2819,In_1830,In_1787);
or U2820 (N_2820,In_1144,In_79);
or U2821 (N_2821,In_1204,In_356);
and U2822 (N_2822,In_1729,In_701);
or U2823 (N_2823,In_1611,In_808);
and U2824 (N_2824,In_1308,In_393);
nor U2825 (N_2825,In_841,In_950);
or U2826 (N_2826,In_1022,In_708);
nand U2827 (N_2827,In_1364,In_855);
nand U2828 (N_2828,In_171,In_1743);
or U2829 (N_2829,In_1257,In_1009);
and U2830 (N_2830,In_1152,In_1590);
or U2831 (N_2831,In_1773,In_862);
or U2832 (N_2832,In_1761,In_416);
nand U2833 (N_2833,In_730,In_805);
nor U2834 (N_2834,In_1033,In_1540);
nor U2835 (N_2835,In_1920,In_647);
and U2836 (N_2836,In_13,In_473);
nand U2837 (N_2837,In_1700,In_1930);
or U2838 (N_2838,In_1355,In_549);
or U2839 (N_2839,In_605,In_892);
and U2840 (N_2840,In_1139,In_1599);
and U2841 (N_2841,In_1265,In_1107);
and U2842 (N_2842,In_1347,In_893);
and U2843 (N_2843,In_273,In_1638);
and U2844 (N_2844,In_1297,In_1160);
nand U2845 (N_2845,In_1725,In_1420);
nor U2846 (N_2846,In_1315,In_530);
nor U2847 (N_2847,In_358,In_953);
and U2848 (N_2848,In_165,In_1570);
nand U2849 (N_2849,In_1305,In_1987);
nor U2850 (N_2850,In_1518,In_169);
or U2851 (N_2851,In_1964,In_123);
and U2852 (N_2852,In_285,In_989);
or U2853 (N_2853,In_1237,In_559);
and U2854 (N_2854,In_1629,In_1224);
xnor U2855 (N_2855,In_323,In_280);
xor U2856 (N_2856,In_522,In_1271);
nand U2857 (N_2857,In_59,In_1990);
xor U2858 (N_2858,In_365,In_762);
nor U2859 (N_2859,In_577,In_1549);
nand U2860 (N_2860,In_1529,In_782);
nand U2861 (N_2861,In_497,In_1382);
and U2862 (N_2862,In_1608,In_1385);
or U2863 (N_2863,In_190,In_0);
nand U2864 (N_2864,In_986,In_633);
nand U2865 (N_2865,In_1790,In_771);
nor U2866 (N_2866,In_1929,In_1546);
nor U2867 (N_2867,In_999,In_361);
nand U2868 (N_2868,In_852,In_1644);
nor U2869 (N_2869,In_908,In_285);
and U2870 (N_2870,In_948,In_174);
nor U2871 (N_2871,In_1937,In_1829);
or U2872 (N_2872,In_160,In_1287);
or U2873 (N_2873,In_144,In_725);
and U2874 (N_2874,In_636,In_338);
nand U2875 (N_2875,In_1089,In_1153);
nor U2876 (N_2876,In_1681,In_363);
and U2877 (N_2877,In_841,In_471);
and U2878 (N_2878,In_1185,In_344);
nand U2879 (N_2879,In_374,In_83);
and U2880 (N_2880,In_1272,In_750);
nand U2881 (N_2881,In_96,In_296);
or U2882 (N_2882,In_957,In_1353);
xnor U2883 (N_2883,In_1602,In_1569);
nor U2884 (N_2884,In_1054,In_805);
or U2885 (N_2885,In_1467,In_1657);
and U2886 (N_2886,In_431,In_554);
and U2887 (N_2887,In_178,In_1776);
nor U2888 (N_2888,In_154,In_1740);
and U2889 (N_2889,In_1569,In_705);
nor U2890 (N_2890,In_906,In_283);
xnor U2891 (N_2891,In_1600,In_536);
or U2892 (N_2892,In_1504,In_604);
nor U2893 (N_2893,In_931,In_799);
or U2894 (N_2894,In_904,In_524);
nand U2895 (N_2895,In_1134,In_705);
or U2896 (N_2896,In_600,In_176);
and U2897 (N_2897,In_883,In_413);
xor U2898 (N_2898,In_422,In_1864);
nor U2899 (N_2899,In_364,In_486);
nor U2900 (N_2900,In_1749,In_1794);
nand U2901 (N_2901,In_1621,In_1191);
nand U2902 (N_2902,In_927,In_1745);
nor U2903 (N_2903,In_1722,In_1160);
nand U2904 (N_2904,In_1952,In_411);
xnor U2905 (N_2905,In_259,In_304);
nor U2906 (N_2906,In_496,In_1606);
nor U2907 (N_2907,In_1959,In_917);
and U2908 (N_2908,In_1313,In_293);
or U2909 (N_2909,In_415,In_963);
nand U2910 (N_2910,In_962,In_177);
nand U2911 (N_2911,In_1922,In_830);
or U2912 (N_2912,In_1914,In_28);
nor U2913 (N_2913,In_1705,In_840);
nor U2914 (N_2914,In_796,In_948);
nor U2915 (N_2915,In_1748,In_1003);
nor U2916 (N_2916,In_1145,In_670);
xor U2917 (N_2917,In_1582,In_1529);
nand U2918 (N_2918,In_465,In_1402);
nor U2919 (N_2919,In_847,In_1877);
and U2920 (N_2920,In_699,In_1363);
nor U2921 (N_2921,In_1154,In_86);
and U2922 (N_2922,In_39,In_1544);
nor U2923 (N_2923,In_486,In_9);
nand U2924 (N_2924,In_1254,In_1571);
nor U2925 (N_2925,In_965,In_796);
or U2926 (N_2926,In_39,In_1005);
nand U2927 (N_2927,In_1368,In_145);
nor U2928 (N_2928,In_573,In_1746);
nand U2929 (N_2929,In_1239,In_1601);
or U2930 (N_2930,In_257,In_1169);
nor U2931 (N_2931,In_898,In_669);
nand U2932 (N_2932,In_1057,In_419);
nand U2933 (N_2933,In_1679,In_981);
and U2934 (N_2934,In_67,In_179);
nor U2935 (N_2935,In_1696,In_1662);
or U2936 (N_2936,In_308,In_432);
or U2937 (N_2937,In_1439,In_1480);
or U2938 (N_2938,In_1930,In_1730);
nor U2939 (N_2939,In_901,In_1069);
nand U2940 (N_2940,In_658,In_954);
or U2941 (N_2941,In_1756,In_708);
or U2942 (N_2942,In_500,In_741);
or U2943 (N_2943,In_1429,In_1725);
and U2944 (N_2944,In_1739,In_1839);
nor U2945 (N_2945,In_1237,In_445);
or U2946 (N_2946,In_1745,In_526);
nor U2947 (N_2947,In_643,In_20);
and U2948 (N_2948,In_1341,In_1013);
nand U2949 (N_2949,In_1463,In_921);
nor U2950 (N_2950,In_144,In_245);
and U2951 (N_2951,In_391,In_263);
and U2952 (N_2952,In_1005,In_270);
nand U2953 (N_2953,In_1452,In_853);
and U2954 (N_2954,In_928,In_997);
or U2955 (N_2955,In_178,In_948);
nor U2956 (N_2956,In_1875,In_1784);
and U2957 (N_2957,In_250,In_1817);
or U2958 (N_2958,In_1639,In_1027);
and U2959 (N_2959,In_1007,In_1077);
and U2960 (N_2960,In_1339,In_1920);
and U2961 (N_2961,In_1701,In_361);
or U2962 (N_2962,In_1515,In_1955);
and U2963 (N_2963,In_451,In_279);
nor U2964 (N_2964,In_1691,In_1166);
nor U2965 (N_2965,In_747,In_733);
and U2966 (N_2966,In_1600,In_182);
nor U2967 (N_2967,In_635,In_119);
xor U2968 (N_2968,In_278,In_1560);
nor U2969 (N_2969,In_1325,In_1442);
nand U2970 (N_2970,In_1703,In_1198);
nand U2971 (N_2971,In_658,In_1176);
nand U2972 (N_2972,In_1674,In_217);
nand U2973 (N_2973,In_522,In_1554);
and U2974 (N_2974,In_1546,In_1772);
or U2975 (N_2975,In_1778,In_336);
or U2976 (N_2976,In_1459,In_1653);
nand U2977 (N_2977,In_1684,In_1536);
and U2978 (N_2978,In_1866,In_300);
and U2979 (N_2979,In_1367,In_788);
and U2980 (N_2980,In_7,In_1917);
nor U2981 (N_2981,In_459,In_238);
and U2982 (N_2982,In_775,In_1287);
xor U2983 (N_2983,In_892,In_1548);
or U2984 (N_2984,In_1752,In_1616);
and U2985 (N_2985,In_1943,In_1290);
and U2986 (N_2986,In_517,In_1291);
nand U2987 (N_2987,In_1972,In_1605);
nand U2988 (N_2988,In_1466,In_1385);
and U2989 (N_2989,In_843,In_382);
nor U2990 (N_2990,In_494,In_994);
and U2991 (N_2991,In_777,In_398);
and U2992 (N_2992,In_1374,In_382);
nor U2993 (N_2993,In_38,In_98);
nand U2994 (N_2994,In_942,In_1013);
or U2995 (N_2995,In_842,In_1175);
xnor U2996 (N_2996,In_111,In_943);
nand U2997 (N_2997,In_1293,In_986);
nand U2998 (N_2998,In_533,In_394);
or U2999 (N_2999,In_61,In_1768);
nor U3000 (N_3000,In_1278,In_685);
nor U3001 (N_3001,In_1395,In_1518);
and U3002 (N_3002,In_58,In_628);
nor U3003 (N_3003,In_1043,In_1115);
or U3004 (N_3004,In_271,In_1159);
or U3005 (N_3005,In_1350,In_1135);
and U3006 (N_3006,In_683,In_1152);
and U3007 (N_3007,In_1075,In_1424);
nor U3008 (N_3008,In_1047,In_881);
nor U3009 (N_3009,In_455,In_47);
xnor U3010 (N_3010,In_1168,In_1554);
nor U3011 (N_3011,In_605,In_1587);
nand U3012 (N_3012,In_1108,In_271);
nor U3013 (N_3013,In_1789,In_679);
and U3014 (N_3014,In_1526,In_920);
nand U3015 (N_3015,In_895,In_1358);
or U3016 (N_3016,In_125,In_528);
and U3017 (N_3017,In_637,In_784);
or U3018 (N_3018,In_1778,In_1017);
nand U3019 (N_3019,In_1556,In_401);
or U3020 (N_3020,In_1468,In_1407);
xnor U3021 (N_3021,In_1856,In_88);
and U3022 (N_3022,In_826,In_718);
and U3023 (N_3023,In_1545,In_1102);
nor U3024 (N_3024,In_808,In_352);
and U3025 (N_3025,In_1593,In_388);
or U3026 (N_3026,In_1693,In_276);
or U3027 (N_3027,In_1193,In_1109);
or U3028 (N_3028,In_131,In_303);
nor U3029 (N_3029,In_901,In_847);
nand U3030 (N_3030,In_1534,In_11);
and U3031 (N_3031,In_1664,In_958);
nor U3032 (N_3032,In_1440,In_1788);
nand U3033 (N_3033,In_5,In_1213);
and U3034 (N_3034,In_743,In_1035);
nor U3035 (N_3035,In_1602,In_1269);
and U3036 (N_3036,In_700,In_1103);
or U3037 (N_3037,In_562,In_1012);
xor U3038 (N_3038,In_198,In_173);
nor U3039 (N_3039,In_1975,In_248);
or U3040 (N_3040,In_153,In_746);
and U3041 (N_3041,In_758,In_1403);
xnor U3042 (N_3042,In_584,In_686);
and U3043 (N_3043,In_511,In_174);
nand U3044 (N_3044,In_350,In_1008);
nor U3045 (N_3045,In_682,In_180);
and U3046 (N_3046,In_480,In_1929);
or U3047 (N_3047,In_736,In_1870);
nor U3048 (N_3048,In_1657,In_953);
or U3049 (N_3049,In_1720,In_506);
nor U3050 (N_3050,In_1961,In_969);
and U3051 (N_3051,In_423,In_1540);
nor U3052 (N_3052,In_1403,In_577);
and U3053 (N_3053,In_739,In_1664);
and U3054 (N_3054,In_1308,In_374);
nor U3055 (N_3055,In_1183,In_1063);
and U3056 (N_3056,In_777,In_373);
nor U3057 (N_3057,In_264,In_689);
nand U3058 (N_3058,In_809,In_700);
nand U3059 (N_3059,In_1229,In_1478);
nand U3060 (N_3060,In_10,In_1342);
xnor U3061 (N_3061,In_159,In_642);
and U3062 (N_3062,In_1368,In_702);
or U3063 (N_3063,In_103,In_1844);
nand U3064 (N_3064,In_1672,In_418);
and U3065 (N_3065,In_620,In_1284);
nand U3066 (N_3066,In_729,In_1555);
and U3067 (N_3067,In_96,In_264);
xor U3068 (N_3068,In_1354,In_0);
nor U3069 (N_3069,In_884,In_388);
or U3070 (N_3070,In_50,In_1628);
and U3071 (N_3071,In_846,In_1469);
nor U3072 (N_3072,In_326,In_1648);
nor U3073 (N_3073,In_1419,In_1082);
or U3074 (N_3074,In_904,In_1099);
nor U3075 (N_3075,In_926,In_963);
nand U3076 (N_3076,In_1658,In_1962);
or U3077 (N_3077,In_1149,In_693);
and U3078 (N_3078,In_1589,In_759);
or U3079 (N_3079,In_1939,In_1158);
xnor U3080 (N_3080,In_857,In_475);
and U3081 (N_3081,In_1923,In_1008);
or U3082 (N_3082,In_1847,In_630);
nor U3083 (N_3083,In_922,In_1795);
nand U3084 (N_3084,In_1426,In_1674);
or U3085 (N_3085,In_1762,In_1516);
nand U3086 (N_3086,In_1222,In_1409);
or U3087 (N_3087,In_99,In_703);
nand U3088 (N_3088,In_213,In_762);
and U3089 (N_3089,In_1735,In_778);
nand U3090 (N_3090,In_662,In_384);
nor U3091 (N_3091,In_139,In_1779);
nand U3092 (N_3092,In_1430,In_719);
nand U3093 (N_3093,In_662,In_371);
or U3094 (N_3094,In_437,In_102);
and U3095 (N_3095,In_698,In_26);
nor U3096 (N_3096,In_1054,In_518);
nor U3097 (N_3097,In_1163,In_1316);
nand U3098 (N_3098,In_860,In_1071);
nor U3099 (N_3099,In_1662,In_1994);
and U3100 (N_3100,In_1061,In_1649);
and U3101 (N_3101,In_1107,In_1220);
or U3102 (N_3102,In_1425,In_1314);
and U3103 (N_3103,In_659,In_1135);
xnor U3104 (N_3104,In_1538,In_531);
and U3105 (N_3105,In_682,In_197);
or U3106 (N_3106,In_986,In_1735);
nor U3107 (N_3107,In_304,In_1661);
nand U3108 (N_3108,In_1961,In_1150);
nand U3109 (N_3109,In_1787,In_363);
and U3110 (N_3110,In_428,In_1609);
and U3111 (N_3111,In_460,In_628);
or U3112 (N_3112,In_570,In_282);
nor U3113 (N_3113,In_1770,In_1750);
nor U3114 (N_3114,In_854,In_1468);
nor U3115 (N_3115,In_1877,In_800);
nor U3116 (N_3116,In_1692,In_112);
or U3117 (N_3117,In_500,In_118);
nand U3118 (N_3118,In_976,In_1925);
or U3119 (N_3119,In_1088,In_1245);
and U3120 (N_3120,In_1726,In_994);
or U3121 (N_3121,In_1779,In_1250);
nand U3122 (N_3122,In_1278,In_1726);
nand U3123 (N_3123,In_857,In_77);
and U3124 (N_3124,In_286,In_1078);
nand U3125 (N_3125,In_1750,In_342);
or U3126 (N_3126,In_756,In_445);
and U3127 (N_3127,In_226,In_814);
nand U3128 (N_3128,In_1480,In_557);
nor U3129 (N_3129,In_825,In_1731);
or U3130 (N_3130,In_1080,In_1264);
nand U3131 (N_3131,In_1350,In_1938);
and U3132 (N_3132,In_1250,In_902);
nor U3133 (N_3133,In_490,In_1034);
or U3134 (N_3134,In_181,In_367);
nor U3135 (N_3135,In_127,In_858);
or U3136 (N_3136,In_1426,In_1562);
and U3137 (N_3137,In_1772,In_1666);
or U3138 (N_3138,In_58,In_556);
and U3139 (N_3139,In_1898,In_1946);
nor U3140 (N_3140,In_519,In_1158);
and U3141 (N_3141,In_174,In_1108);
or U3142 (N_3142,In_1975,In_1233);
nand U3143 (N_3143,In_1554,In_1968);
xor U3144 (N_3144,In_1891,In_803);
xor U3145 (N_3145,In_216,In_1307);
nand U3146 (N_3146,In_1009,In_1098);
or U3147 (N_3147,In_958,In_121);
nor U3148 (N_3148,In_1395,In_979);
or U3149 (N_3149,In_1810,In_866);
nand U3150 (N_3150,In_428,In_1439);
xor U3151 (N_3151,In_504,In_207);
and U3152 (N_3152,In_1683,In_34);
nor U3153 (N_3153,In_585,In_1033);
or U3154 (N_3154,In_1144,In_1876);
nor U3155 (N_3155,In_239,In_446);
or U3156 (N_3156,In_1076,In_865);
nand U3157 (N_3157,In_1460,In_528);
nand U3158 (N_3158,In_895,In_46);
nand U3159 (N_3159,In_747,In_403);
nor U3160 (N_3160,In_1100,In_647);
and U3161 (N_3161,In_1518,In_1534);
nor U3162 (N_3162,In_1654,In_843);
nand U3163 (N_3163,In_1230,In_1675);
xnor U3164 (N_3164,In_602,In_1942);
nand U3165 (N_3165,In_630,In_30);
nand U3166 (N_3166,In_1603,In_1172);
xor U3167 (N_3167,In_995,In_1447);
nand U3168 (N_3168,In_413,In_822);
and U3169 (N_3169,In_1024,In_1496);
nand U3170 (N_3170,In_1347,In_1658);
or U3171 (N_3171,In_727,In_975);
xor U3172 (N_3172,In_408,In_1964);
xor U3173 (N_3173,In_483,In_545);
nor U3174 (N_3174,In_593,In_616);
or U3175 (N_3175,In_1751,In_605);
or U3176 (N_3176,In_1263,In_1050);
or U3177 (N_3177,In_605,In_1979);
xor U3178 (N_3178,In_1929,In_505);
xnor U3179 (N_3179,In_140,In_1505);
xnor U3180 (N_3180,In_381,In_1233);
or U3181 (N_3181,In_1487,In_770);
or U3182 (N_3182,In_1938,In_1517);
nor U3183 (N_3183,In_1270,In_683);
or U3184 (N_3184,In_886,In_357);
nor U3185 (N_3185,In_660,In_1689);
nor U3186 (N_3186,In_1770,In_79);
and U3187 (N_3187,In_130,In_492);
xnor U3188 (N_3188,In_1956,In_1648);
and U3189 (N_3189,In_1842,In_1257);
and U3190 (N_3190,In_1210,In_1606);
nand U3191 (N_3191,In_686,In_1969);
and U3192 (N_3192,In_796,In_903);
and U3193 (N_3193,In_150,In_103);
nand U3194 (N_3194,In_157,In_388);
and U3195 (N_3195,In_174,In_576);
nor U3196 (N_3196,In_1276,In_741);
and U3197 (N_3197,In_78,In_480);
xnor U3198 (N_3198,In_493,In_464);
nor U3199 (N_3199,In_526,In_137);
nand U3200 (N_3200,In_391,In_1230);
nand U3201 (N_3201,In_65,In_838);
nor U3202 (N_3202,In_1988,In_1425);
and U3203 (N_3203,In_1221,In_580);
or U3204 (N_3204,In_835,In_134);
nand U3205 (N_3205,In_877,In_298);
nor U3206 (N_3206,In_1527,In_737);
xor U3207 (N_3207,In_1857,In_1708);
and U3208 (N_3208,In_920,In_784);
nand U3209 (N_3209,In_193,In_916);
nor U3210 (N_3210,In_1377,In_1594);
nor U3211 (N_3211,In_177,In_203);
and U3212 (N_3212,In_352,In_387);
and U3213 (N_3213,In_521,In_1190);
nand U3214 (N_3214,In_1128,In_1297);
nor U3215 (N_3215,In_633,In_1725);
and U3216 (N_3216,In_982,In_402);
nand U3217 (N_3217,In_157,In_1458);
and U3218 (N_3218,In_1640,In_34);
nand U3219 (N_3219,In_941,In_833);
and U3220 (N_3220,In_1021,In_543);
nor U3221 (N_3221,In_1027,In_525);
and U3222 (N_3222,In_1713,In_101);
nor U3223 (N_3223,In_1503,In_1877);
or U3224 (N_3224,In_1232,In_773);
xor U3225 (N_3225,In_1848,In_376);
and U3226 (N_3226,In_1007,In_951);
or U3227 (N_3227,In_942,In_1020);
nand U3228 (N_3228,In_711,In_793);
nand U3229 (N_3229,In_1321,In_1855);
and U3230 (N_3230,In_1926,In_915);
nand U3231 (N_3231,In_1761,In_1350);
and U3232 (N_3232,In_1711,In_1643);
or U3233 (N_3233,In_397,In_1779);
or U3234 (N_3234,In_1919,In_1532);
nand U3235 (N_3235,In_1215,In_63);
and U3236 (N_3236,In_477,In_620);
and U3237 (N_3237,In_621,In_480);
and U3238 (N_3238,In_895,In_413);
or U3239 (N_3239,In_1792,In_998);
nor U3240 (N_3240,In_1894,In_744);
nor U3241 (N_3241,In_577,In_24);
and U3242 (N_3242,In_1617,In_540);
nand U3243 (N_3243,In_1426,In_456);
and U3244 (N_3244,In_327,In_31);
or U3245 (N_3245,In_1668,In_1592);
or U3246 (N_3246,In_20,In_834);
and U3247 (N_3247,In_1291,In_828);
nor U3248 (N_3248,In_1596,In_880);
or U3249 (N_3249,In_343,In_297);
and U3250 (N_3250,In_1914,In_1836);
nand U3251 (N_3251,In_26,In_1141);
and U3252 (N_3252,In_1239,In_727);
nor U3253 (N_3253,In_735,In_811);
xnor U3254 (N_3254,In_1084,In_1339);
and U3255 (N_3255,In_121,In_1950);
nand U3256 (N_3256,In_500,In_710);
and U3257 (N_3257,In_1665,In_676);
and U3258 (N_3258,In_1773,In_1089);
and U3259 (N_3259,In_1925,In_1969);
nor U3260 (N_3260,In_936,In_1486);
xor U3261 (N_3261,In_322,In_1492);
and U3262 (N_3262,In_1827,In_326);
and U3263 (N_3263,In_1774,In_726);
nand U3264 (N_3264,In_1966,In_197);
or U3265 (N_3265,In_793,In_944);
nand U3266 (N_3266,In_1639,In_321);
and U3267 (N_3267,In_1678,In_56);
nor U3268 (N_3268,In_1493,In_1765);
nand U3269 (N_3269,In_1319,In_1220);
nand U3270 (N_3270,In_575,In_628);
and U3271 (N_3271,In_912,In_1999);
or U3272 (N_3272,In_422,In_1271);
and U3273 (N_3273,In_104,In_158);
or U3274 (N_3274,In_1875,In_319);
nand U3275 (N_3275,In_812,In_207);
nand U3276 (N_3276,In_1842,In_470);
and U3277 (N_3277,In_1988,In_989);
and U3278 (N_3278,In_1973,In_59);
xor U3279 (N_3279,In_119,In_1460);
and U3280 (N_3280,In_1830,In_1806);
nand U3281 (N_3281,In_388,In_1860);
nand U3282 (N_3282,In_244,In_433);
and U3283 (N_3283,In_354,In_506);
nor U3284 (N_3284,In_709,In_1180);
nand U3285 (N_3285,In_603,In_1593);
xor U3286 (N_3286,In_1425,In_1309);
nor U3287 (N_3287,In_520,In_247);
and U3288 (N_3288,In_1914,In_177);
or U3289 (N_3289,In_555,In_734);
nor U3290 (N_3290,In_541,In_1716);
and U3291 (N_3291,In_801,In_1289);
nand U3292 (N_3292,In_584,In_780);
nor U3293 (N_3293,In_1598,In_1567);
xnor U3294 (N_3294,In_1153,In_414);
nor U3295 (N_3295,In_1307,In_1050);
nor U3296 (N_3296,In_1798,In_1737);
and U3297 (N_3297,In_110,In_1322);
nor U3298 (N_3298,In_916,In_1213);
or U3299 (N_3299,In_1961,In_910);
and U3300 (N_3300,In_948,In_1449);
and U3301 (N_3301,In_1354,In_291);
xnor U3302 (N_3302,In_521,In_58);
nand U3303 (N_3303,In_1853,In_1677);
and U3304 (N_3304,In_996,In_133);
xnor U3305 (N_3305,In_734,In_525);
or U3306 (N_3306,In_418,In_1925);
nor U3307 (N_3307,In_211,In_971);
nand U3308 (N_3308,In_749,In_1774);
nor U3309 (N_3309,In_1321,In_1319);
or U3310 (N_3310,In_1500,In_854);
and U3311 (N_3311,In_340,In_452);
nand U3312 (N_3312,In_1439,In_488);
and U3313 (N_3313,In_21,In_690);
or U3314 (N_3314,In_1185,In_1312);
and U3315 (N_3315,In_1217,In_53);
or U3316 (N_3316,In_1684,In_1758);
nor U3317 (N_3317,In_888,In_786);
or U3318 (N_3318,In_1363,In_588);
nor U3319 (N_3319,In_482,In_564);
and U3320 (N_3320,In_1637,In_503);
or U3321 (N_3321,In_1063,In_334);
and U3322 (N_3322,In_924,In_1896);
and U3323 (N_3323,In_1336,In_1036);
and U3324 (N_3324,In_1454,In_383);
and U3325 (N_3325,In_1164,In_36);
xor U3326 (N_3326,In_1640,In_830);
and U3327 (N_3327,In_579,In_210);
or U3328 (N_3328,In_489,In_173);
and U3329 (N_3329,In_1202,In_1190);
nor U3330 (N_3330,In_1872,In_1991);
or U3331 (N_3331,In_562,In_230);
and U3332 (N_3332,In_1877,In_1691);
or U3333 (N_3333,In_785,In_15);
or U3334 (N_3334,In_1945,In_1769);
nor U3335 (N_3335,In_398,In_56);
and U3336 (N_3336,In_183,In_766);
and U3337 (N_3337,In_1512,In_382);
nand U3338 (N_3338,In_1796,In_563);
nor U3339 (N_3339,In_909,In_728);
nand U3340 (N_3340,In_1264,In_1190);
nand U3341 (N_3341,In_1811,In_859);
and U3342 (N_3342,In_1335,In_656);
xnor U3343 (N_3343,In_1056,In_1571);
nand U3344 (N_3344,In_114,In_1236);
and U3345 (N_3345,In_1367,In_393);
and U3346 (N_3346,In_1597,In_482);
or U3347 (N_3347,In_976,In_1126);
or U3348 (N_3348,In_919,In_1725);
or U3349 (N_3349,In_889,In_1362);
and U3350 (N_3350,In_654,In_1989);
nand U3351 (N_3351,In_867,In_549);
or U3352 (N_3352,In_1901,In_1637);
nand U3353 (N_3353,In_816,In_1275);
nand U3354 (N_3354,In_1028,In_459);
or U3355 (N_3355,In_750,In_1060);
nand U3356 (N_3356,In_856,In_1743);
and U3357 (N_3357,In_1255,In_599);
nor U3358 (N_3358,In_332,In_271);
and U3359 (N_3359,In_205,In_1387);
and U3360 (N_3360,In_275,In_1583);
nor U3361 (N_3361,In_86,In_928);
nand U3362 (N_3362,In_1827,In_1895);
nor U3363 (N_3363,In_176,In_1040);
or U3364 (N_3364,In_1120,In_956);
and U3365 (N_3365,In_445,In_114);
nor U3366 (N_3366,In_139,In_778);
nor U3367 (N_3367,In_1519,In_1898);
nand U3368 (N_3368,In_1207,In_762);
or U3369 (N_3369,In_440,In_1989);
or U3370 (N_3370,In_15,In_1682);
nand U3371 (N_3371,In_1606,In_337);
nor U3372 (N_3372,In_1870,In_691);
nor U3373 (N_3373,In_1307,In_1996);
and U3374 (N_3374,In_1638,In_873);
or U3375 (N_3375,In_1058,In_1913);
nand U3376 (N_3376,In_1133,In_1253);
and U3377 (N_3377,In_1542,In_651);
nor U3378 (N_3378,In_818,In_1487);
or U3379 (N_3379,In_1017,In_1838);
nand U3380 (N_3380,In_561,In_25);
nor U3381 (N_3381,In_1277,In_535);
nand U3382 (N_3382,In_447,In_1255);
or U3383 (N_3383,In_184,In_1853);
or U3384 (N_3384,In_1903,In_1689);
nor U3385 (N_3385,In_416,In_1440);
nor U3386 (N_3386,In_104,In_1695);
and U3387 (N_3387,In_725,In_560);
nor U3388 (N_3388,In_1535,In_1299);
nor U3389 (N_3389,In_1498,In_1900);
or U3390 (N_3390,In_1370,In_1092);
or U3391 (N_3391,In_295,In_301);
nor U3392 (N_3392,In_505,In_1208);
or U3393 (N_3393,In_853,In_51);
nor U3394 (N_3394,In_1280,In_1998);
or U3395 (N_3395,In_1218,In_1697);
and U3396 (N_3396,In_1566,In_572);
or U3397 (N_3397,In_1251,In_961);
and U3398 (N_3398,In_478,In_914);
and U3399 (N_3399,In_1894,In_700);
and U3400 (N_3400,In_1844,In_1623);
or U3401 (N_3401,In_928,In_1830);
xnor U3402 (N_3402,In_1623,In_1288);
or U3403 (N_3403,In_1187,In_1933);
nor U3404 (N_3404,In_521,In_1383);
and U3405 (N_3405,In_1312,In_398);
or U3406 (N_3406,In_1859,In_263);
or U3407 (N_3407,In_413,In_810);
or U3408 (N_3408,In_389,In_1173);
nor U3409 (N_3409,In_1724,In_1699);
nor U3410 (N_3410,In_125,In_1261);
or U3411 (N_3411,In_334,In_613);
nor U3412 (N_3412,In_1731,In_1213);
or U3413 (N_3413,In_617,In_227);
xor U3414 (N_3414,In_1053,In_84);
nand U3415 (N_3415,In_1537,In_1769);
nor U3416 (N_3416,In_136,In_1607);
nor U3417 (N_3417,In_41,In_22);
nor U3418 (N_3418,In_675,In_1654);
nor U3419 (N_3419,In_1714,In_1073);
and U3420 (N_3420,In_157,In_1520);
nor U3421 (N_3421,In_1154,In_1698);
or U3422 (N_3422,In_1757,In_1271);
xor U3423 (N_3423,In_972,In_1831);
and U3424 (N_3424,In_602,In_1735);
or U3425 (N_3425,In_760,In_327);
nor U3426 (N_3426,In_845,In_350);
nand U3427 (N_3427,In_365,In_1237);
and U3428 (N_3428,In_1879,In_313);
and U3429 (N_3429,In_458,In_1055);
nand U3430 (N_3430,In_1646,In_1156);
nand U3431 (N_3431,In_569,In_971);
nor U3432 (N_3432,In_1757,In_1149);
or U3433 (N_3433,In_149,In_264);
nand U3434 (N_3434,In_1830,In_1734);
or U3435 (N_3435,In_797,In_1769);
xor U3436 (N_3436,In_279,In_1134);
and U3437 (N_3437,In_365,In_1863);
nand U3438 (N_3438,In_752,In_372);
nor U3439 (N_3439,In_1868,In_947);
nand U3440 (N_3440,In_374,In_1703);
and U3441 (N_3441,In_52,In_1699);
nand U3442 (N_3442,In_1978,In_218);
xor U3443 (N_3443,In_1800,In_1572);
and U3444 (N_3444,In_884,In_537);
or U3445 (N_3445,In_962,In_579);
and U3446 (N_3446,In_1483,In_1637);
xnor U3447 (N_3447,In_1581,In_688);
and U3448 (N_3448,In_196,In_443);
nand U3449 (N_3449,In_386,In_78);
or U3450 (N_3450,In_397,In_351);
and U3451 (N_3451,In_1197,In_1722);
or U3452 (N_3452,In_1120,In_808);
nor U3453 (N_3453,In_979,In_730);
and U3454 (N_3454,In_185,In_68);
nor U3455 (N_3455,In_497,In_286);
and U3456 (N_3456,In_1816,In_969);
nor U3457 (N_3457,In_555,In_518);
and U3458 (N_3458,In_724,In_1531);
xor U3459 (N_3459,In_631,In_164);
nand U3460 (N_3460,In_528,In_983);
and U3461 (N_3461,In_1386,In_132);
nor U3462 (N_3462,In_1978,In_833);
and U3463 (N_3463,In_1929,In_6);
nand U3464 (N_3464,In_807,In_1063);
xor U3465 (N_3465,In_1195,In_679);
and U3466 (N_3466,In_990,In_370);
nor U3467 (N_3467,In_796,In_165);
nand U3468 (N_3468,In_1224,In_289);
and U3469 (N_3469,In_1976,In_1601);
and U3470 (N_3470,In_1020,In_949);
or U3471 (N_3471,In_38,In_851);
nor U3472 (N_3472,In_1052,In_1733);
nand U3473 (N_3473,In_1520,In_522);
or U3474 (N_3474,In_1529,In_1867);
and U3475 (N_3475,In_864,In_1577);
nor U3476 (N_3476,In_294,In_1762);
nor U3477 (N_3477,In_576,In_458);
nand U3478 (N_3478,In_1642,In_648);
or U3479 (N_3479,In_1194,In_1151);
nor U3480 (N_3480,In_822,In_1665);
nor U3481 (N_3481,In_228,In_657);
or U3482 (N_3482,In_481,In_387);
nor U3483 (N_3483,In_1005,In_794);
nor U3484 (N_3484,In_728,In_969);
nor U3485 (N_3485,In_1969,In_800);
nand U3486 (N_3486,In_439,In_1732);
nor U3487 (N_3487,In_276,In_283);
nand U3488 (N_3488,In_275,In_1503);
nand U3489 (N_3489,In_1805,In_513);
and U3490 (N_3490,In_1484,In_69);
nor U3491 (N_3491,In_1117,In_1755);
and U3492 (N_3492,In_1528,In_1544);
or U3493 (N_3493,In_1065,In_1865);
nand U3494 (N_3494,In_1685,In_657);
xor U3495 (N_3495,In_1269,In_1110);
and U3496 (N_3496,In_937,In_141);
and U3497 (N_3497,In_644,In_145);
nand U3498 (N_3498,In_1793,In_1104);
or U3499 (N_3499,In_33,In_777);
and U3500 (N_3500,In_987,In_1734);
xor U3501 (N_3501,In_1369,In_1144);
nor U3502 (N_3502,In_286,In_707);
or U3503 (N_3503,In_1520,In_974);
nand U3504 (N_3504,In_1606,In_1461);
or U3505 (N_3505,In_136,In_1860);
nand U3506 (N_3506,In_1756,In_1497);
and U3507 (N_3507,In_1016,In_1758);
or U3508 (N_3508,In_1321,In_1284);
xor U3509 (N_3509,In_6,In_880);
nor U3510 (N_3510,In_129,In_1588);
xnor U3511 (N_3511,In_1222,In_1660);
or U3512 (N_3512,In_893,In_461);
or U3513 (N_3513,In_1384,In_439);
or U3514 (N_3514,In_873,In_846);
or U3515 (N_3515,In_102,In_852);
and U3516 (N_3516,In_1754,In_1741);
or U3517 (N_3517,In_12,In_48);
or U3518 (N_3518,In_481,In_1189);
and U3519 (N_3519,In_1418,In_549);
or U3520 (N_3520,In_1623,In_1360);
and U3521 (N_3521,In_1072,In_872);
and U3522 (N_3522,In_1240,In_1136);
nor U3523 (N_3523,In_1667,In_283);
and U3524 (N_3524,In_1071,In_702);
and U3525 (N_3525,In_627,In_1003);
or U3526 (N_3526,In_451,In_1658);
or U3527 (N_3527,In_1845,In_1875);
nand U3528 (N_3528,In_400,In_411);
or U3529 (N_3529,In_1403,In_201);
or U3530 (N_3530,In_1855,In_1797);
nand U3531 (N_3531,In_818,In_693);
and U3532 (N_3532,In_338,In_1705);
or U3533 (N_3533,In_99,In_468);
and U3534 (N_3534,In_1392,In_498);
or U3535 (N_3535,In_748,In_1394);
nand U3536 (N_3536,In_330,In_629);
and U3537 (N_3537,In_1363,In_305);
nor U3538 (N_3538,In_71,In_1953);
and U3539 (N_3539,In_1815,In_1742);
and U3540 (N_3540,In_1646,In_1954);
xor U3541 (N_3541,In_1400,In_547);
nor U3542 (N_3542,In_947,In_1340);
nor U3543 (N_3543,In_1851,In_1861);
nor U3544 (N_3544,In_1645,In_1135);
and U3545 (N_3545,In_421,In_286);
nor U3546 (N_3546,In_633,In_136);
or U3547 (N_3547,In_78,In_467);
and U3548 (N_3548,In_867,In_394);
nand U3549 (N_3549,In_118,In_722);
nand U3550 (N_3550,In_1332,In_1929);
or U3551 (N_3551,In_1990,In_370);
xnor U3552 (N_3552,In_1797,In_1762);
and U3553 (N_3553,In_1965,In_1028);
nand U3554 (N_3554,In_967,In_518);
and U3555 (N_3555,In_974,In_807);
nor U3556 (N_3556,In_1576,In_1026);
nand U3557 (N_3557,In_336,In_862);
and U3558 (N_3558,In_1186,In_239);
xnor U3559 (N_3559,In_1484,In_1420);
or U3560 (N_3560,In_1082,In_1738);
nand U3561 (N_3561,In_1615,In_23);
or U3562 (N_3562,In_439,In_594);
nor U3563 (N_3563,In_615,In_1935);
and U3564 (N_3564,In_1768,In_60);
nand U3565 (N_3565,In_1799,In_983);
nand U3566 (N_3566,In_681,In_526);
nor U3567 (N_3567,In_1691,In_272);
nor U3568 (N_3568,In_632,In_428);
nor U3569 (N_3569,In_1477,In_624);
or U3570 (N_3570,In_358,In_1050);
or U3571 (N_3571,In_1201,In_882);
xor U3572 (N_3572,In_1313,In_1861);
and U3573 (N_3573,In_1854,In_1676);
or U3574 (N_3574,In_374,In_1439);
nor U3575 (N_3575,In_421,In_461);
or U3576 (N_3576,In_1804,In_1227);
and U3577 (N_3577,In_1383,In_1291);
or U3578 (N_3578,In_181,In_175);
nand U3579 (N_3579,In_1129,In_1342);
or U3580 (N_3580,In_1442,In_1863);
nor U3581 (N_3581,In_1498,In_999);
or U3582 (N_3582,In_493,In_544);
xnor U3583 (N_3583,In_1076,In_96);
nand U3584 (N_3584,In_782,In_1783);
or U3585 (N_3585,In_769,In_705);
and U3586 (N_3586,In_872,In_1830);
and U3587 (N_3587,In_1730,In_446);
nand U3588 (N_3588,In_964,In_360);
or U3589 (N_3589,In_41,In_1670);
nor U3590 (N_3590,In_970,In_307);
nand U3591 (N_3591,In_1453,In_734);
nor U3592 (N_3592,In_1769,In_1323);
and U3593 (N_3593,In_223,In_1874);
nor U3594 (N_3594,In_1774,In_507);
and U3595 (N_3595,In_248,In_1596);
nor U3596 (N_3596,In_1520,In_320);
or U3597 (N_3597,In_718,In_1033);
or U3598 (N_3598,In_1822,In_1364);
and U3599 (N_3599,In_482,In_1604);
nor U3600 (N_3600,In_1270,In_449);
and U3601 (N_3601,In_1210,In_306);
nand U3602 (N_3602,In_555,In_1670);
or U3603 (N_3603,In_828,In_1297);
nand U3604 (N_3604,In_951,In_609);
nor U3605 (N_3605,In_1806,In_868);
nand U3606 (N_3606,In_935,In_826);
nand U3607 (N_3607,In_813,In_816);
or U3608 (N_3608,In_1289,In_398);
nand U3609 (N_3609,In_1213,In_279);
and U3610 (N_3610,In_1225,In_966);
and U3611 (N_3611,In_654,In_653);
nand U3612 (N_3612,In_243,In_1505);
nor U3613 (N_3613,In_517,In_1904);
nand U3614 (N_3614,In_813,In_461);
nand U3615 (N_3615,In_1416,In_251);
nand U3616 (N_3616,In_1064,In_1078);
and U3617 (N_3617,In_1454,In_1363);
or U3618 (N_3618,In_823,In_992);
xnor U3619 (N_3619,In_244,In_41);
and U3620 (N_3620,In_244,In_657);
nand U3621 (N_3621,In_1809,In_169);
nand U3622 (N_3622,In_1137,In_1584);
xnor U3623 (N_3623,In_1814,In_1975);
nand U3624 (N_3624,In_407,In_1145);
or U3625 (N_3625,In_336,In_1293);
and U3626 (N_3626,In_258,In_636);
nor U3627 (N_3627,In_1893,In_981);
nor U3628 (N_3628,In_48,In_1130);
nor U3629 (N_3629,In_1125,In_79);
nor U3630 (N_3630,In_120,In_988);
and U3631 (N_3631,In_1409,In_1303);
and U3632 (N_3632,In_1120,In_71);
nand U3633 (N_3633,In_908,In_229);
or U3634 (N_3634,In_425,In_297);
nor U3635 (N_3635,In_1711,In_711);
nor U3636 (N_3636,In_102,In_1540);
or U3637 (N_3637,In_1206,In_1838);
and U3638 (N_3638,In_1050,In_674);
nor U3639 (N_3639,In_1924,In_1272);
and U3640 (N_3640,In_1762,In_936);
and U3641 (N_3641,In_1248,In_1202);
xor U3642 (N_3642,In_1913,In_913);
and U3643 (N_3643,In_1591,In_1261);
nor U3644 (N_3644,In_746,In_548);
and U3645 (N_3645,In_675,In_1645);
or U3646 (N_3646,In_386,In_1993);
and U3647 (N_3647,In_1663,In_1475);
or U3648 (N_3648,In_1766,In_1669);
and U3649 (N_3649,In_1844,In_178);
xor U3650 (N_3650,In_1835,In_1953);
nor U3651 (N_3651,In_1472,In_1343);
or U3652 (N_3652,In_1775,In_30);
or U3653 (N_3653,In_5,In_1251);
nor U3654 (N_3654,In_1942,In_1357);
nand U3655 (N_3655,In_1651,In_50);
nand U3656 (N_3656,In_1825,In_1318);
or U3657 (N_3657,In_1447,In_1426);
and U3658 (N_3658,In_1555,In_512);
nand U3659 (N_3659,In_1133,In_1245);
or U3660 (N_3660,In_1465,In_113);
or U3661 (N_3661,In_1380,In_1583);
and U3662 (N_3662,In_322,In_1265);
or U3663 (N_3663,In_91,In_472);
nor U3664 (N_3664,In_462,In_1365);
nand U3665 (N_3665,In_456,In_1781);
nor U3666 (N_3666,In_93,In_1644);
and U3667 (N_3667,In_1614,In_1552);
xor U3668 (N_3668,In_1926,In_1534);
and U3669 (N_3669,In_58,In_923);
or U3670 (N_3670,In_589,In_1307);
or U3671 (N_3671,In_1589,In_43);
nand U3672 (N_3672,In_19,In_1959);
nand U3673 (N_3673,In_1342,In_298);
xor U3674 (N_3674,In_70,In_1315);
and U3675 (N_3675,In_835,In_1370);
nor U3676 (N_3676,In_283,In_125);
or U3677 (N_3677,In_303,In_795);
xor U3678 (N_3678,In_1805,In_1880);
and U3679 (N_3679,In_380,In_441);
and U3680 (N_3680,In_1740,In_481);
or U3681 (N_3681,In_448,In_4);
and U3682 (N_3682,In_774,In_1952);
or U3683 (N_3683,In_439,In_978);
or U3684 (N_3684,In_128,In_1936);
and U3685 (N_3685,In_680,In_548);
or U3686 (N_3686,In_1515,In_1582);
or U3687 (N_3687,In_1013,In_567);
nand U3688 (N_3688,In_1988,In_1321);
xor U3689 (N_3689,In_1400,In_82);
and U3690 (N_3690,In_342,In_195);
nor U3691 (N_3691,In_1082,In_1255);
and U3692 (N_3692,In_1855,In_979);
and U3693 (N_3693,In_498,In_1569);
nand U3694 (N_3694,In_1608,In_1135);
or U3695 (N_3695,In_752,In_1113);
or U3696 (N_3696,In_815,In_250);
xor U3697 (N_3697,In_46,In_81);
or U3698 (N_3698,In_1757,In_1921);
or U3699 (N_3699,In_253,In_167);
nand U3700 (N_3700,In_739,In_669);
or U3701 (N_3701,In_355,In_1438);
nand U3702 (N_3702,In_1057,In_1161);
nand U3703 (N_3703,In_1961,In_953);
nor U3704 (N_3704,In_1758,In_1024);
nor U3705 (N_3705,In_586,In_79);
and U3706 (N_3706,In_219,In_1875);
nor U3707 (N_3707,In_1344,In_668);
and U3708 (N_3708,In_331,In_1223);
and U3709 (N_3709,In_1713,In_751);
nand U3710 (N_3710,In_339,In_1988);
or U3711 (N_3711,In_1026,In_807);
or U3712 (N_3712,In_1952,In_181);
nor U3713 (N_3713,In_646,In_496);
xor U3714 (N_3714,In_945,In_77);
and U3715 (N_3715,In_936,In_633);
nor U3716 (N_3716,In_1668,In_754);
nor U3717 (N_3717,In_310,In_239);
nor U3718 (N_3718,In_1844,In_848);
xnor U3719 (N_3719,In_471,In_1872);
or U3720 (N_3720,In_24,In_1091);
and U3721 (N_3721,In_1708,In_1775);
and U3722 (N_3722,In_1499,In_455);
nand U3723 (N_3723,In_251,In_1773);
or U3724 (N_3724,In_1169,In_946);
xor U3725 (N_3725,In_816,In_444);
and U3726 (N_3726,In_1672,In_375);
or U3727 (N_3727,In_1654,In_1838);
and U3728 (N_3728,In_872,In_779);
and U3729 (N_3729,In_1705,In_380);
or U3730 (N_3730,In_972,In_1031);
nor U3731 (N_3731,In_108,In_1911);
or U3732 (N_3732,In_868,In_1902);
or U3733 (N_3733,In_241,In_347);
nand U3734 (N_3734,In_1560,In_1543);
nand U3735 (N_3735,In_533,In_1112);
and U3736 (N_3736,In_186,In_1965);
and U3737 (N_3737,In_682,In_400);
nand U3738 (N_3738,In_399,In_1115);
and U3739 (N_3739,In_595,In_635);
nand U3740 (N_3740,In_1572,In_16);
or U3741 (N_3741,In_678,In_312);
or U3742 (N_3742,In_580,In_1281);
or U3743 (N_3743,In_183,In_1450);
nand U3744 (N_3744,In_1320,In_1337);
nor U3745 (N_3745,In_908,In_758);
and U3746 (N_3746,In_317,In_732);
and U3747 (N_3747,In_1370,In_76);
nor U3748 (N_3748,In_651,In_723);
nand U3749 (N_3749,In_1643,In_1002);
nand U3750 (N_3750,In_1267,In_72);
and U3751 (N_3751,In_1865,In_1235);
or U3752 (N_3752,In_1507,In_54);
and U3753 (N_3753,In_1179,In_1694);
and U3754 (N_3754,In_1772,In_569);
nand U3755 (N_3755,In_1671,In_1386);
or U3756 (N_3756,In_406,In_869);
or U3757 (N_3757,In_1829,In_1245);
or U3758 (N_3758,In_448,In_229);
nand U3759 (N_3759,In_588,In_632);
nand U3760 (N_3760,In_1572,In_1384);
or U3761 (N_3761,In_1919,In_1646);
nor U3762 (N_3762,In_242,In_1429);
and U3763 (N_3763,In_417,In_1493);
xor U3764 (N_3764,In_728,In_1573);
and U3765 (N_3765,In_1172,In_1860);
nor U3766 (N_3766,In_796,In_516);
nor U3767 (N_3767,In_999,In_1325);
and U3768 (N_3768,In_557,In_870);
nand U3769 (N_3769,In_1480,In_1314);
and U3770 (N_3770,In_329,In_1670);
and U3771 (N_3771,In_832,In_1262);
nor U3772 (N_3772,In_569,In_1479);
or U3773 (N_3773,In_334,In_278);
or U3774 (N_3774,In_129,In_165);
nor U3775 (N_3775,In_650,In_867);
nand U3776 (N_3776,In_1773,In_200);
xnor U3777 (N_3777,In_689,In_375);
nand U3778 (N_3778,In_1676,In_295);
and U3779 (N_3779,In_216,In_1285);
nor U3780 (N_3780,In_415,In_1862);
nand U3781 (N_3781,In_1397,In_1254);
nand U3782 (N_3782,In_94,In_1401);
or U3783 (N_3783,In_1778,In_1669);
or U3784 (N_3784,In_1959,In_1387);
and U3785 (N_3785,In_342,In_1357);
nor U3786 (N_3786,In_860,In_1301);
nor U3787 (N_3787,In_794,In_1662);
and U3788 (N_3788,In_301,In_852);
nor U3789 (N_3789,In_805,In_1223);
nor U3790 (N_3790,In_1357,In_1811);
and U3791 (N_3791,In_424,In_273);
nand U3792 (N_3792,In_1956,In_1729);
nand U3793 (N_3793,In_724,In_1559);
nor U3794 (N_3794,In_1445,In_1389);
or U3795 (N_3795,In_354,In_998);
xor U3796 (N_3796,In_1015,In_1878);
nand U3797 (N_3797,In_139,In_1308);
nor U3798 (N_3798,In_161,In_1959);
nand U3799 (N_3799,In_1119,In_944);
nor U3800 (N_3800,In_128,In_669);
or U3801 (N_3801,In_981,In_1422);
nand U3802 (N_3802,In_634,In_1372);
nor U3803 (N_3803,In_1695,In_1035);
nand U3804 (N_3804,In_1967,In_678);
nand U3805 (N_3805,In_1829,In_1751);
or U3806 (N_3806,In_825,In_510);
nor U3807 (N_3807,In_828,In_122);
xor U3808 (N_3808,In_1862,In_657);
and U3809 (N_3809,In_1221,In_1002);
or U3810 (N_3810,In_318,In_492);
xnor U3811 (N_3811,In_1991,In_825);
nand U3812 (N_3812,In_1189,In_1837);
and U3813 (N_3813,In_1700,In_1973);
or U3814 (N_3814,In_1131,In_1682);
and U3815 (N_3815,In_1932,In_1933);
nand U3816 (N_3816,In_1054,In_1418);
nand U3817 (N_3817,In_1953,In_242);
nand U3818 (N_3818,In_1309,In_773);
nand U3819 (N_3819,In_1087,In_369);
or U3820 (N_3820,In_1684,In_1491);
or U3821 (N_3821,In_17,In_1262);
or U3822 (N_3822,In_1459,In_489);
nand U3823 (N_3823,In_1312,In_1926);
and U3824 (N_3824,In_516,In_1906);
nand U3825 (N_3825,In_1510,In_1936);
xor U3826 (N_3826,In_776,In_558);
or U3827 (N_3827,In_1980,In_1913);
or U3828 (N_3828,In_1897,In_480);
nor U3829 (N_3829,In_1749,In_817);
or U3830 (N_3830,In_1055,In_1878);
nor U3831 (N_3831,In_1768,In_946);
xnor U3832 (N_3832,In_1724,In_1352);
and U3833 (N_3833,In_389,In_1776);
or U3834 (N_3834,In_785,In_86);
and U3835 (N_3835,In_753,In_1877);
and U3836 (N_3836,In_103,In_439);
or U3837 (N_3837,In_1558,In_58);
xor U3838 (N_3838,In_1047,In_754);
nor U3839 (N_3839,In_1631,In_1800);
and U3840 (N_3840,In_262,In_472);
and U3841 (N_3841,In_873,In_1253);
and U3842 (N_3842,In_1984,In_1309);
nand U3843 (N_3843,In_551,In_410);
or U3844 (N_3844,In_1475,In_601);
and U3845 (N_3845,In_609,In_925);
and U3846 (N_3846,In_747,In_1023);
or U3847 (N_3847,In_1260,In_1655);
or U3848 (N_3848,In_348,In_1043);
nor U3849 (N_3849,In_925,In_859);
or U3850 (N_3850,In_1504,In_1932);
nor U3851 (N_3851,In_516,In_1564);
nor U3852 (N_3852,In_1337,In_299);
nand U3853 (N_3853,In_1369,In_1290);
and U3854 (N_3854,In_1255,In_193);
nor U3855 (N_3855,In_112,In_1034);
xor U3856 (N_3856,In_1818,In_178);
or U3857 (N_3857,In_811,In_891);
or U3858 (N_3858,In_1201,In_981);
nand U3859 (N_3859,In_1648,In_1375);
nand U3860 (N_3860,In_1988,In_1271);
and U3861 (N_3861,In_372,In_1);
and U3862 (N_3862,In_1819,In_628);
or U3863 (N_3863,In_666,In_294);
nor U3864 (N_3864,In_1861,In_645);
nand U3865 (N_3865,In_1641,In_989);
and U3866 (N_3866,In_222,In_344);
and U3867 (N_3867,In_46,In_1118);
xor U3868 (N_3868,In_259,In_431);
or U3869 (N_3869,In_1256,In_413);
nor U3870 (N_3870,In_1879,In_961);
and U3871 (N_3871,In_1088,In_1743);
nor U3872 (N_3872,In_979,In_1524);
xnor U3873 (N_3873,In_1661,In_1780);
or U3874 (N_3874,In_128,In_957);
nor U3875 (N_3875,In_1242,In_108);
xnor U3876 (N_3876,In_1674,In_1102);
nand U3877 (N_3877,In_506,In_727);
or U3878 (N_3878,In_866,In_1585);
nor U3879 (N_3879,In_1645,In_1182);
nor U3880 (N_3880,In_131,In_1332);
nor U3881 (N_3881,In_292,In_1068);
nand U3882 (N_3882,In_768,In_342);
or U3883 (N_3883,In_889,In_122);
and U3884 (N_3884,In_1421,In_1679);
nor U3885 (N_3885,In_181,In_198);
xnor U3886 (N_3886,In_1820,In_1761);
and U3887 (N_3887,In_184,In_193);
or U3888 (N_3888,In_29,In_1668);
nand U3889 (N_3889,In_1447,In_470);
xnor U3890 (N_3890,In_881,In_1111);
nand U3891 (N_3891,In_1819,In_777);
xnor U3892 (N_3892,In_1564,In_870);
nor U3893 (N_3893,In_516,In_1773);
and U3894 (N_3894,In_1555,In_1471);
or U3895 (N_3895,In_696,In_1590);
nor U3896 (N_3896,In_1980,In_250);
xnor U3897 (N_3897,In_1440,In_1225);
or U3898 (N_3898,In_645,In_1834);
xnor U3899 (N_3899,In_1578,In_1408);
and U3900 (N_3900,In_1093,In_139);
nor U3901 (N_3901,In_1812,In_1083);
nand U3902 (N_3902,In_106,In_654);
and U3903 (N_3903,In_574,In_1086);
nand U3904 (N_3904,In_1908,In_53);
or U3905 (N_3905,In_1988,In_690);
and U3906 (N_3906,In_148,In_754);
and U3907 (N_3907,In_669,In_1908);
or U3908 (N_3908,In_17,In_512);
nand U3909 (N_3909,In_1659,In_1238);
and U3910 (N_3910,In_1542,In_1934);
nand U3911 (N_3911,In_105,In_1175);
nor U3912 (N_3912,In_282,In_133);
nand U3913 (N_3913,In_533,In_629);
nor U3914 (N_3914,In_1300,In_493);
and U3915 (N_3915,In_646,In_272);
and U3916 (N_3916,In_1962,In_1476);
nor U3917 (N_3917,In_1889,In_1979);
nor U3918 (N_3918,In_740,In_1628);
xnor U3919 (N_3919,In_779,In_566);
or U3920 (N_3920,In_1168,In_5);
and U3921 (N_3921,In_1895,In_697);
and U3922 (N_3922,In_1504,In_1374);
nor U3923 (N_3923,In_1345,In_1408);
nor U3924 (N_3924,In_1701,In_681);
nor U3925 (N_3925,In_1893,In_1668);
and U3926 (N_3926,In_460,In_1646);
nand U3927 (N_3927,In_13,In_1912);
or U3928 (N_3928,In_363,In_1439);
or U3929 (N_3929,In_1032,In_869);
nor U3930 (N_3930,In_678,In_764);
nor U3931 (N_3931,In_617,In_1645);
nor U3932 (N_3932,In_1821,In_1894);
nand U3933 (N_3933,In_558,In_1747);
nor U3934 (N_3934,In_954,In_1683);
or U3935 (N_3935,In_1563,In_328);
and U3936 (N_3936,In_1971,In_1175);
or U3937 (N_3937,In_235,In_1210);
or U3938 (N_3938,In_289,In_31);
nor U3939 (N_3939,In_90,In_764);
nor U3940 (N_3940,In_47,In_1563);
and U3941 (N_3941,In_392,In_132);
nor U3942 (N_3942,In_66,In_1077);
nand U3943 (N_3943,In_1189,In_7);
nand U3944 (N_3944,In_768,In_561);
nand U3945 (N_3945,In_1184,In_1568);
or U3946 (N_3946,In_1687,In_1156);
nand U3947 (N_3947,In_1374,In_1386);
nor U3948 (N_3948,In_325,In_1971);
nor U3949 (N_3949,In_170,In_627);
nand U3950 (N_3950,In_560,In_13);
nand U3951 (N_3951,In_166,In_1908);
or U3952 (N_3952,In_1357,In_73);
nand U3953 (N_3953,In_1191,In_266);
and U3954 (N_3954,In_448,In_1961);
xor U3955 (N_3955,In_1301,In_49);
nand U3956 (N_3956,In_879,In_231);
or U3957 (N_3957,In_915,In_1421);
and U3958 (N_3958,In_235,In_49);
or U3959 (N_3959,In_1514,In_855);
and U3960 (N_3960,In_1259,In_392);
and U3961 (N_3961,In_617,In_1570);
nand U3962 (N_3962,In_1748,In_1133);
or U3963 (N_3963,In_654,In_206);
nor U3964 (N_3964,In_948,In_6);
xor U3965 (N_3965,In_1563,In_738);
and U3966 (N_3966,In_262,In_1536);
nand U3967 (N_3967,In_741,In_1583);
nor U3968 (N_3968,In_1683,In_1020);
and U3969 (N_3969,In_523,In_1009);
and U3970 (N_3970,In_1693,In_196);
or U3971 (N_3971,In_224,In_876);
nor U3972 (N_3972,In_150,In_1726);
xor U3973 (N_3973,In_1922,In_1793);
nand U3974 (N_3974,In_1222,In_100);
or U3975 (N_3975,In_1474,In_357);
xor U3976 (N_3976,In_219,In_1254);
nand U3977 (N_3977,In_1339,In_834);
nor U3978 (N_3978,In_1478,In_81);
and U3979 (N_3979,In_1087,In_455);
nand U3980 (N_3980,In_11,In_546);
nand U3981 (N_3981,In_20,In_1225);
nor U3982 (N_3982,In_1599,In_93);
and U3983 (N_3983,In_801,In_1490);
nand U3984 (N_3984,In_850,In_871);
xnor U3985 (N_3985,In_1791,In_1742);
or U3986 (N_3986,In_1262,In_1916);
nor U3987 (N_3987,In_1538,In_1787);
or U3988 (N_3988,In_262,In_1240);
and U3989 (N_3989,In_1421,In_1987);
nor U3990 (N_3990,In_272,In_31);
nand U3991 (N_3991,In_214,In_346);
xor U3992 (N_3992,In_1476,In_1924);
nor U3993 (N_3993,In_241,In_73);
or U3994 (N_3994,In_666,In_180);
and U3995 (N_3995,In_835,In_893);
nor U3996 (N_3996,In_1261,In_1575);
and U3997 (N_3997,In_430,In_972);
nor U3998 (N_3998,In_1835,In_429);
or U3999 (N_3999,In_358,In_285);
nor U4000 (N_4000,In_161,In_693);
nand U4001 (N_4001,In_1822,In_1994);
or U4002 (N_4002,In_1125,In_533);
and U4003 (N_4003,In_907,In_494);
and U4004 (N_4004,In_1317,In_64);
xor U4005 (N_4005,In_1706,In_452);
nand U4006 (N_4006,In_1360,In_1203);
nand U4007 (N_4007,In_248,In_1430);
or U4008 (N_4008,In_878,In_1008);
nand U4009 (N_4009,In_898,In_1815);
nand U4010 (N_4010,In_1886,In_607);
nand U4011 (N_4011,In_973,In_432);
and U4012 (N_4012,In_286,In_1940);
nor U4013 (N_4013,In_334,In_1431);
and U4014 (N_4014,In_1727,In_1954);
or U4015 (N_4015,In_218,In_353);
or U4016 (N_4016,In_684,In_1816);
and U4017 (N_4017,In_1281,In_1369);
or U4018 (N_4018,In_63,In_1281);
xor U4019 (N_4019,In_449,In_1082);
nand U4020 (N_4020,In_1567,In_483);
nor U4021 (N_4021,In_279,In_469);
and U4022 (N_4022,In_330,In_60);
nor U4023 (N_4023,In_372,In_1617);
nand U4024 (N_4024,In_281,In_1569);
xnor U4025 (N_4025,In_1513,In_1232);
and U4026 (N_4026,In_799,In_1733);
or U4027 (N_4027,In_1767,In_180);
or U4028 (N_4028,In_526,In_29);
or U4029 (N_4029,In_1365,In_353);
or U4030 (N_4030,In_1500,In_34);
nor U4031 (N_4031,In_319,In_821);
nor U4032 (N_4032,In_594,In_1502);
nand U4033 (N_4033,In_973,In_47);
nor U4034 (N_4034,In_638,In_590);
xor U4035 (N_4035,In_442,In_611);
nand U4036 (N_4036,In_1223,In_230);
or U4037 (N_4037,In_1082,In_844);
nand U4038 (N_4038,In_675,In_451);
xor U4039 (N_4039,In_1843,In_98);
nand U4040 (N_4040,In_559,In_704);
and U4041 (N_4041,In_927,In_1964);
nand U4042 (N_4042,In_865,In_711);
and U4043 (N_4043,In_1914,In_82);
nand U4044 (N_4044,In_1809,In_1705);
and U4045 (N_4045,In_240,In_1989);
nand U4046 (N_4046,In_255,In_1238);
nor U4047 (N_4047,In_251,In_484);
nand U4048 (N_4048,In_1225,In_407);
nand U4049 (N_4049,In_169,In_1271);
nor U4050 (N_4050,In_1863,In_765);
nor U4051 (N_4051,In_139,In_1324);
and U4052 (N_4052,In_1995,In_890);
or U4053 (N_4053,In_1918,In_892);
nor U4054 (N_4054,In_886,In_1229);
nor U4055 (N_4055,In_1700,In_1221);
or U4056 (N_4056,In_1881,In_853);
or U4057 (N_4057,In_689,In_111);
nor U4058 (N_4058,In_299,In_62);
nor U4059 (N_4059,In_246,In_1671);
or U4060 (N_4060,In_1890,In_149);
nor U4061 (N_4061,In_93,In_686);
nor U4062 (N_4062,In_390,In_359);
and U4063 (N_4063,In_1317,In_1544);
or U4064 (N_4064,In_1852,In_386);
nor U4065 (N_4065,In_1176,In_970);
nand U4066 (N_4066,In_770,In_1760);
or U4067 (N_4067,In_276,In_1092);
nor U4068 (N_4068,In_565,In_275);
and U4069 (N_4069,In_1160,In_1284);
or U4070 (N_4070,In_959,In_299);
nor U4071 (N_4071,In_891,In_1857);
nand U4072 (N_4072,In_284,In_340);
nand U4073 (N_4073,In_893,In_349);
nor U4074 (N_4074,In_284,In_1474);
or U4075 (N_4075,In_794,In_796);
nand U4076 (N_4076,In_212,In_126);
or U4077 (N_4077,In_325,In_254);
nor U4078 (N_4078,In_1245,In_1218);
and U4079 (N_4079,In_784,In_398);
and U4080 (N_4080,In_454,In_1154);
nor U4081 (N_4081,In_1630,In_85);
or U4082 (N_4082,In_112,In_728);
nand U4083 (N_4083,In_178,In_954);
nor U4084 (N_4084,In_1093,In_321);
nor U4085 (N_4085,In_1052,In_98);
nand U4086 (N_4086,In_1460,In_1148);
and U4087 (N_4087,In_1170,In_1023);
nor U4088 (N_4088,In_896,In_578);
nor U4089 (N_4089,In_18,In_434);
or U4090 (N_4090,In_508,In_1726);
or U4091 (N_4091,In_1537,In_1293);
xnor U4092 (N_4092,In_470,In_1222);
and U4093 (N_4093,In_1862,In_843);
nand U4094 (N_4094,In_788,In_320);
or U4095 (N_4095,In_350,In_1553);
xor U4096 (N_4096,In_1501,In_152);
and U4097 (N_4097,In_1735,In_1955);
nand U4098 (N_4098,In_704,In_1918);
nor U4099 (N_4099,In_196,In_1222);
nand U4100 (N_4100,In_1008,In_587);
or U4101 (N_4101,In_1142,In_374);
and U4102 (N_4102,In_879,In_645);
nor U4103 (N_4103,In_1101,In_1297);
or U4104 (N_4104,In_139,In_1792);
nor U4105 (N_4105,In_1249,In_1306);
or U4106 (N_4106,In_1227,In_609);
and U4107 (N_4107,In_1164,In_1516);
and U4108 (N_4108,In_150,In_1354);
xor U4109 (N_4109,In_1793,In_1907);
nand U4110 (N_4110,In_1096,In_1860);
nand U4111 (N_4111,In_984,In_1670);
and U4112 (N_4112,In_7,In_1001);
or U4113 (N_4113,In_369,In_850);
or U4114 (N_4114,In_1048,In_734);
or U4115 (N_4115,In_222,In_1779);
nor U4116 (N_4116,In_605,In_1606);
nand U4117 (N_4117,In_991,In_1153);
nand U4118 (N_4118,In_174,In_1790);
nor U4119 (N_4119,In_1041,In_1667);
and U4120 (N_4120,In_1281,In_824);
and U4121 (N_4121,In_41,In_1946);
or U4122 (N_4122,In_483,In_1969);
nor U4123 (N_4123,In_876,In_890);
nand U4124 (N_4124,In_1043,In_1815);
and U4125 (N_4125,In_840,In_707);
and U4126 (N_4126,In_636,In_1099);
nand U4127 (N_4127,In_784,In_1855);
and U4128 (N_4128,In_1532,In_951);
nor U4129 (N_4129,In_1161,In_605);
and U4130 (N_4130,In_1084,In_1934);
or U4131 (N_4131,In_225,In_936);
nor U4132 (N_4132,In_739,In_1182);
or U4133 (N_4133,In_1826,In_368);
and U4134 (N_4134,In_1315,In_1337);
nor U4135 (N_4135,In_1616,In_1028);
xnor U4136 (N_4136,In_680,In_988);
or U4137 (N_4137,In_1388,In_1426);
or U4138 (N_4138,In_757,In_64);
nor U4139 (N_4139,In_1734,In_1426);
and U4140 (N_4140,In_1235,In_1234);
nor U4141 (N_4141,In_441,In_75);
nand U4142 (N_4142,In_293,In_1732);
xor U4143 (N_4143,In_1734,In_1454);
nor U4144 (N_4144,In_655,In_1935);
nand U4145 (N_4145,In_181,In_312);
or U4146 (N_4146,In_925,In_712);
or U4147 (N_4147,In_819,In_1079);
nand U4148 (N_4148,In_1277,In_350);
nor U4149 (N_4149,In_1413,In_1089);
and U4150 (N_4150,In_1096,In_326);
nand U4151 (N_4151,In_360,In_460);
and U4152 (N_4152,In_1939,In_49);
and U4153 (N_4153,In_182,In_1389);
and U4154 (N_4154,In_1645,In_1786);
nor U4155 (N_4155,In_483,In_1634);
and U4156 (N_4156,In_573,In_1376);
nand U4157 (N_4157,In_350,In_741);
and U4158 (N_4158,In_54,In_1653);
and U4159 (N_4159,In_1838,In_635);
or U4160 (N_4160,In_1274,In_1571);
and U4161 (N_4161,In_1062,In_1326);
nor U4162 (N_4162,In_1547,In_991);
nor U4163 (N_4163,In_1469,In_490);
or U4164 (N_4164,In_554,In_584);
or U4165 (N_4165,In_1908,In_685);
and U4166 (N_4166,In_855,In_910);
nor U4167 (N_4167,In_1787,In_695);
nand U4168 (N_4168,In_870,In_1369);
xnor U4169 (N_4169,In_63,In_4);
nand U4170 (N_4170,In_1881,In_1469);
or U4171 (N_4171,In_504,In_1565);
nor U4172 (N_4172,In_546,In_1418);
or U4173 (N_4173,In_67,In_1657);
or U4174 (N_4174,In_1981,In_1833);
nand U4175 (N_4175,In_1137,In_1875);
xor U4176 (N_4176,In_1184,In_803);
nand U4177 (N_4177,In_1303,In_1666);
and U4178 (N_4178,In_1855,In_230);
nor U4179 (N_4179,In_1976,In_988);
nand U4180 (N_4180,In_70,In_1048);
nor U4181 (N_4181,In_590,In_1112);
xor U4182 (N_4182,In_1235,In_181);
and U4183 (N_4183,In_1590,In_1523);
nand U4184 (N_4184,In_794,In_567);
and U4185 (N_4185,In_1959,In_812);
or U4186 (N_4186,In_623,In_1101);
nor U4187 (N_4187,In_1698,In_423);
and U4188 (N_4188,In_998,In_1652);
and U4189 (N_4189,In_1020,In_252);
nor U4190 (N_4190,In_1016,In_967);
or U4191 (N_4191,In_1633,In_1240);
nand U4192 (N_4192,In_1679,In_274);
and U4193 (N_4193,In_505,In_785);
nor U4194 (N_4194,In_463,In_957);
and U4195 (N_4195,In_507,In_1832);
nand U4196 (N_4196,In_1427,In_1725);
and U4197 (N_4197,In_534,In_1532);
nand U4198 (N_4198,In_1304,In_740);
and U4199 (N_4199,In_486,In_22);
or U4200 (N_4200,In_1897,In_1139);
nor U4201 (N_4201,In_1999,In_1048);
and U4202 (N_4202,In_832,In_1452);
and U4203 (N_4203,In_423,In_631);
and U4204 (N_4204,In_1464,In_1109);
nand U4205 (N_4205,In_525,In_999);
or U4206 (N_4206,In_608,In_463);
nor U4207 (N_4207,In_1878,In_1110);
nand U4208 (N_4208,In_960,In_881);
nor U4209 (N_4209,In_1958,In_919);
xnor U4210 (N_4210,In_1909,In_978);
or U4211 (N_4211,In_827,In_1645);
and U4212 (N_4212,In_1071,In_1003);
nand U4213 (N_4213,In_1145,In_334);
nor U4214 (N_4214,In_892,In_1599);
nand U4215 (N_4215,In_747,In_1212);
or U4216 (N_4216,In_79,In_73);
or U4217 (N_4217,In_44,In_1125);
nor U4218 (N_4218,In_779,In_556);
nor U4219 (N_4219,In_443,In_1982);
nor U4220 (N_4220,In_1014,In_1401);
nor U4221 (N_4221,In_1627,In_1257);
nor U4222 (N_4222,In_851,In_1879);
and U4223 (N_4223,In_1447,In_1012);
nand U4224 (N_4224,In_704,In_110);
and U4225 (N_4225,In_1402,In_1796);
nand U4226 (N_4226,In_842,In_880);
and U4227 (N_4227,In_1967,In_1196);
nand U4228 (N_4228,In_1193,In_600);
nor U4229 (N_4229,In_882,In_1940);
nand U4230 (N_4230,In_1294,In_1933);
or U4231 (N_4231,In_306,In_866);
and U4232 (N_4232,In_528,In_1661);
and U4233 (N_4233,In_176,In_1126);
and U4234 (N_4234,In_1778,In_1722);
nor U4235 (N_4235,In_1641,In_1836);
and U4236 (N_4236,In_1208,In_754);
nor U4237 (N_4237,In_533,In_1261);
or U4238 (N_4238,In_1074,In_822);
or U4239 (N_4239,In_340,In_1361);
and U4240 (N_4240,In_1920,In_934);
nand U4241 (N_4241,In_190,In_1892);
nor U4242 (N_4242,In_1229,In_318);
or U4243 (N_4243,In_102,In_720);
or U4244 (N_4244,In_12,In_39);
and U4245 (N_4245,In_240,In_947);
or U4246 (N_4246,In_672,In_1929);
and U4247 (N_4247,In_1945,In_393);
nand U4248 (N_4248,In_301,In_1252);
and U4249 (N_4249,In_1803,In_244);
nand U4250 (N_4250,In_765,In_716);
or U4251 (N_4251,In_427,In_991);
or U4252 (N_4252,In_511,In_496);
xor U4253 (N_4253,In_1466,In_107);
or U4254 (N_4254,In_1731,In_1649);
nor U4255 (N_4255,In_170,In_1055);
or U4256 (N_4256,In_726,In_1604);
or U4257 (N_4257,In_1604,In_1263);
xnor U4258 (N_4258,In_412,In_764);
or U4259 (N_4259,In_1985,In_316);
nand U4260 (N_4260,In_180,In_527);
nand U4261 (N_4261,In_815,In_1466);
nor U4262 (N_4262,In_512,In_849);
nand U4263 (N_4263,In_1218,In_332);
nor U4264 (N_4264,In_1072,In_148);
and U4265 (N_4265,In_1126,In_1316);
and U4266 (N_4266,In_1027,In_1062);
nor U4267 (N_4267,In_500,In_471);
or U4268 (N_4268,In_1607,In_1547);
nor U4269 (N_4269,In_437,In_745);
and U4270 (N_4270,In_544,In_600);
and U4271 (N_4271,In_1761,In_1567);
or U4272 (N_4272,In_582,In_1341);
and U4273 (N_4273,In_1332,In_1943);
nand U4274 (N_4274,In_937,In_1851);
nand U4275 (N_4275,In_862,In_1472);
nand U4276 (N_4276,In_190,In_549);
or U4277 (N_4277,In_1428,In_720);
and U4278 (N_4278,In_772,In_338);
and U4279 (N_4279,In_1232,In_388);
nand U4280 (N_4280,In_1735,In_1288);
nor U4281 (N_4281,In_942,In_1448);
and U4282 (N_4282,In_1793,In_1521);
and U4283 (N_4283,In_514,In_1151);
nor U4284 (N_4284,In_1333,In_742);
xor U4285 (N_4285,In_1796,In_397);
and U4286 (N_4286,In_1019,In_1726);
or U4287 (N_4287,In_36,In_243);
nand U4288 (N_4288,In_266,In_526);
nor U4289 (N_4289,In_1425,In_1748);
nand U4290 (N_4290,In_146,In_252);
xor U4291 (N_4291,In_1146,In_802);
and U4292 (N_4292,In_1935,In_860);
or U4293 (N_4293,In_285,In_818);
nand U4294 (N_4294,In_718,In_1148);
nand U4295 (N_4295,In_1988,In_1436);
nor U4296 (N_4296,In_1255,In_819);
nand U4297 (N_4297,In_1483,In_1525);
xor U4298 (N_4298,In_524,In_748);
nand U4299 (N_4299,In_554,In_895);
or U4300 (N_4300,In_234,In_1873);
xor U4301 (N_4301,In_1165,In_420);
or U4302 (N_4302,In_7,In_965);
or U4303 (N_4303,In_1168,In_1505);
or U4304 (N_4304,In_917,In_1941);
xnor U4305 (N_4305,In_202,In_907);
and U4306 (N_4306,In_1729,In_1531);
or U4307 (N_4307,In_1618,In_541);
nor U4308 (N_4308,In_1585,In_284);
nand U4309 (N_4309,In_1492,In_681);
xnor U4310 (N_4310,In_216,In_645);
nand U4311 (N_4311,In_1954,In_1892);
and U4312 (N_4312,In_924,In_945);
or U4313 (N_4313,In_243,In_50);
nor U4314 (N_4314,In_1725,In_676);
nor U4315 (N_4315,In_1557,In_647);
or U4316 (N_4316,In_1644,In_1226);
nor U4317 (N_4317,In_487,In_936);
nor U4318 (N_4318,In_599,In_70);
and U4319 (N_4319,In_1537,In_952);
and U4320 (N_4320,In_96,In_976);
nand U4321 (N_4321,In_1988,In_51);
xnor U4322 (N_4322,In_171,In_328);
nor U4323 (N_4323,In_1699,In_1650);
nand U4324 (N_4324,In_936,In_338);
xor U4325 (N_4325,In_710,In_1739);
nand U4326 (N_4326,In_1905,In_1071);
and U4327 (N_4327,In_1605,In_1876);
nand U4328 (N_4328,In_1339,In_410);
or U4329 (N_4329,In_785,In_1384);
and U4330 (N_4330,In_505,In_1900);
nand U4331 (N_4331,In_594,In_367);
or U4332 (N_4332,In_99,In_1587);
or U4333 (N_4333,In_893,In_1103);
nor U4334 (N_4334,In_965,In_131);
nor U4335 (N_4335,In_1865,In_612);
xor U4336 (N_4336,In_597,In_1102);
and U4337 (N_4337,In_255,In_377);
nor U4338 (N_4338,In_472,In_1131);
and U4339 (N_4339,In_1808,In_404);
and U4340 (N_4340,In_1061,In_1692);
or U4341 (N_4341,In_1840,In_121);
nor U4342 (N_4342,In_789,In_86);
nand U4343 (N_4343,In_1283,In_759);
nand U4344 (N_4344,In_1218,In_235);
nand U4345 (N_4345,In_417,In_1868);
nor U4346 (N_4346,In_1883,In_1352);
nor U4347 (N_4347,In_562,In_1995);
or U4348 (N_4348,In_1261,In_370);
or U4349 (N_4349,In_1729,In_1804);
or U4350 (N_4350,In_714,In_1064);
xnor U4351 (N_4351,In_756,In_559);
and U4352 (N_4352,In_1247,In_1305);
nor U4353 (N_4353,In_1573,In_650);
nor U4354 (N_4354,In_295,In_1423);
nand U4355 (N_4355,In_848,In_416);
or U4356 (N_4356,In_925,In_8);
or U4357 (N_4357,In_310,In_740);
and U4358 (N_4358,In_1472,In_285);
or U4359 (N_4359,In_171,In_604);
and U4360 (N_4360,In_1412,In_776);
nor U4361 (N_4361,In_1739,In_24);
nor U4362 (N_4362,In_518,In_1555);
or U4363 (N_4363,In_1983,In_443);
nand U4364 (N_4364,In_661,In_1313);
or U4365 (N_4365,In_1777,In_984);
and U4366 (N_4366,In_323,In_1319);
xor U4367 (N_4367,In_1926,In_518);
and U4368 (N_4368,In_509,In_1066);
and U4369 (N_4369,In_944,In_184);
or U4370 (N_4370,In_356,In_1300);
nand U4371 (N_4371,In_407,In_227);
nor U4372 (N_4372,In_1914,In_1677);
nand U4373 (N_4373,In_682,In_1852);
nor U4374 (N_4374,In_541,In_867);
and U4375 (N_4375,In_1790,In_1206);
nand U4376 (N_4376,In_577,In_1129);
and U4377 (N_4377,In_1692,In_1651);
xnor U4378 (N_4378,In_685,In_535);
and U4379 (N_4379,In_1546,In_1836);
and U4380 (N_4380,In_1020,In_1564);
nor U4381 (N_4381,In_277,In_1933);
and U4382 (N_4382,In_1386,In_1044);
nor U4383 (N_4383,In_1557,In_1268);
nor U4384 (N_4384,In_1297,In_1087);
nor U4385 (N_4385,In_1189,In_385);
and U4386 (N_4386,In_1262,In_1260);
nor U4387 (N_4387,In_1191,In_1897);
nor U4388 (N_4388,In_874,In_1490);
xor U4389 (N_4389,In_861,In_1734);
and U4390 (N_4390,In_973,In_1490);
nor U4391 (N_4391,In_1015,In_1217);
or U4392 (N_4392,In_360,In_513);
nor U4393 (N_4393,In_344,In_1765);
nand U4394 (N_4394,In_119,In_770);
nand U4395 (N_4395,In_538,In_733);
xor U4396 (N_4396,In_1927,In_1477);
or U4397 (N_4397,In_1041,In_1219);
or U4398 (N_4398,In_154,In_1192);
and U4399 (N_4399,In_1686,In_1238);
and U4400 (N_4400,In_488,In_344);
xnor U4401 (N_4401,In_806,In_1379);
xnor U4402 (N_4402,In_518,In_282);
and U4403 (N_4403,In_928,In_1227);
and U4404 (N_4404,In_999,In_1213);
xnor U4405 (N_4405,In_1675,In_1955);
nor U4406 (N_4406,In_800,In_1496);
or U4407 (N_4407,In_1660,In_640);
nand U4408 (N_4408,In_1195,In_293);
nor U4409 (N_4409,In_672,In_832);
nor U4410 (N_4410,In_1342,In_578);
or U4411 (N_4411,In_479,In_1481);
and U4412 (N_4412,In_1035,In_137);
nand U4413 (N_4413,In_1129,In_866);
xnor U4414 (N_4414,In_692,In_1949);
or U4415 (N_4415,In_1849,In_1082);
nor U4416 (N_4416,In_617,In_1506);
nor U4417 (N_4417,In_632,In_1553);
or U4418 (N_4418,In_947,In_65);
nand U4419 (N_4419,In_1654,In_1494);
nand U4420 (N_4420,In_956,In_1223);
and U4421 (N_4421,In_1465,In_777);
nor U4422 (N_4422,In_1381,In_425);
or U4423 (N_4423,In_298,In_1936);
nand U4424 (N_4424,In_1345,In_1935);
and U4425 (N_4425,In_649,In_148);
nand U4426 (N_4426,In_792,In_745);
or U4427 (N_4427,In_815,In_1871);
nor U4428 (N_4428,In_1110,In_860);
xor U4429 (N_4429,In_518,In_1771);
and U4430 (N_4430,In_1526,In_797);
nand U4431 (N_4431,In_368,In_535);
nand U4432 (N_4432,In_229,In_991);
and U4433 (N_4433,In_1662,In_869);
xor U4434 (N_4434,In_177,In_1365);
or U4435 (N_4435,In_173,In_931);
nand U4436 (N_4436,In_23,In_114);
and U4437 (N_4437,In_1908,In_1823);
or U4438 (N_4438,In_1658,In_978);
nand U4439 (N_4439,In_1097,In_1095);
nand U4440 (N_4440,In_481,In_644);
or U4441 (N_4441,In_1451,In_868);
and U4442 (N_4442,In_615,In_58);
or U4443 (N_4443,In_1974,In_155);
and U4444 (N_4444,In_59,In_784);
and U4445 (N_4445,In_1997,In_484);
nand U4446 (N_4446,In_1613,In_1005);
nand U4447 (N_4447,In_1811,In_1442);
xor U4448 (N_4448,In_57,In_264);
nor U4449 (N_4449,In_1566,In_1237);
xor U4450 (N_4450,In_383,In_1988);
nand U4451 (N_4451,In_1552,In_960);
and U4452 (N_4452,In_699,In_1328);
and U4453 (N_4453,In_1968,In_288);
or U4454 (N_4454,In_966,In_1192);
nand U4455 (N_4455,In_1230,In_1219);
nand U4456 (N_4456,In_61,In_541);
nor U4457 (N_4457,In_1610,In_898);
or U4458 (N_4458,In_454,In_1153);
nor U4459 (N_4459,In_302,In_1217);
and U4460 (N_4460,In_1568,In_450);
and U4461 (N_4461,In_1134,In_679);
nor U4462 (N_4462,In_1853,In_1940);
or U4463 (N_4463,In_591,In_306);
nor U4464 (N_4464,In_964,In_1821);
and U4465 (N_4465,In_1362,In_1646);
nand U4466 (N_4466,In_1052,In_1932);
nand U4467 (N_4467,In_1202,In_1236);
or U4468 (N_4468,In_458,In_76);
xnor U4469 (N_4469,In_12,In_976);
or U4470 (N_4470,In_676,In_870);
nor U4471 (N_4471,In_778,In_17);
nor U4472 (N_4472,In_1429,In_736);
and U4473 (N_4473,In_54,In_594);
or U4474 (N_4474,In_1912,In_996);
nand U4475 (N_4475,In_104,In_1677);
and U4476 (N_4476,In_583,In_1646);
nor U4477 (N_4477,In_631,In_1276);
nand U4478 (N_4478,In_1239,In_1505);
nor U4479 (N_4479,In_1314,In_56);
or U4480 (N_4480,In_1218,In_920);
nor U4481 (N_4481,In_1054,In_1218);
nor U4482 (N_4482,In_1187,In_1540);
and U4483 (N_4483,In_773,In_564);
or U4484 (N_4484,In_679,In_1855);
or U4485 (N_4485,In_1225,In_789);
nor U4486 (N_4486,In_1592,In_682);
or U4487 (N_4487,In_1204,In_842);
and U4488 (N_4488,In_374,In_92);
nor U4489 (N_4489,In_1454,In_418);
xnor U4490 (N_4490,In_334,In_307);
and U4491 (N_4491,In_1709,In_303);
nand U4492 (N_4492,In_1900,In_646);
or U4493 (N_4493,In_1588,In_235);
or U4494 (N_4494,In_368,In_137);
or U4495 (N_4495,In_455,In_931);
nand U4496 (N_4496,In_707,In_1472);
nand U4497 (N_4497,In_891,In_1714);
nand U4498 (N_4498,In_1051,In_1202);
and U4499 (N_4499,In_1067,In_744);
nand U4500 (N_4500,In_984,In_1895);
and U4501 (N_4501,In_1014,In_1632);
or U4502 (N_4502,In_1382,In_559);
nor U4503 (N_4503,In_1662,In_1897);
or U4504 (N_4504,In_326,In_126);
xor U4505 (N_4505,In_1239,In_1116);
nand U4506 (N_4506,In_1700,In_1342);
nor U4507 (N_4507,In_1867,In_1155);
or U4508 (N_4508,In_1694,In_1176);
or U4509 (N_4509,In_689,In_1818);
and U4510 (N_4510,In_964,In_224);
nand U4511 (N_4511,In_1468,In_1190);
nand U4512 (N_4512,In_20,In_69);
nor U4513 (N_4513,In_87,In_835);
and U4514 (N_4514,In_1820,In_1619);
and U4515 (N_4515,In_45,In_1521);
and U4516 (N_4516,In_1599,In_1729);
and U4517 (N_4517,In_1628,In_746);
or U4518 (N_4518,In_1163,In_1272);
or U4519 (N_4519,In_945,In_1171);
xor U4520 (N_4520,In_599,In_817);
and U4521 (N_4521,In_530,In_476);
nor U4522 (N_4522,In_653,In_648);
nor U4523 (N_4523,In_1473,In_1667);
nand U4524 (N_4524,In_741,In_1411);
or U4525 (N_4525,In_687,In_1757);
xnor U4526 (N_4526,In_1158,In_701);
xor U4527 (N_4527,In_396,In_89);
or U4528 (N_4528,In_839,In_106);
nand U4529 (N_4529,In_1017,In_1253);
nor U4530 (N_4530,In_1938,In_1933);
and U4531 (N_4531,In_1739,In_1524);
or U4532 (N_4532,In_1563,In_1086);
or U4533 (N_4533,In_1767,In_1194);
and U4534 (N_4534,In_1502,In_1118);
or U4535 (N_4535,In_1341,In_957);
nor U4536 (N_4536,In_271,In_640);
nand U4537 (N_4537,In_236,In_1806);
or U4538 (N_4538,In_187,In_1797);
and U4539 (N_4539,In_944,In_192);
and U4540 (N_4540,In_1532,In_177);
nor U4541 (N_4541,In_912,In_160);
nor U4542 (N_4542,In_1137,In_620);
or U4543 (N_4543,In_719,In_441);
nor U4544 (N_4544,In_450,In_26);
nand U4545 (N_4545,In_38,In_99);
nor U4546 (N_4546,In_1020,In_1211);
or U4547 (N_4547,In_1356,In_1828);
or U4548 (N_4548,In_1267,In_1516);
or U4549 (N_4549,In_1141,In_403);
and U4550 (N_4550,In_694,In_1408);
and U4551 (N_4551,In_306,In_934);
and U4552 (N_4552,In_313,In_131);
xnor U4553 (N_4553,In_1425,In_1684);
nor U4554 (N_4554,In_1722,In_1216);
or U4555 (N_4555,In_182,In_1856);
and U4556 (N_4556,In_1548,In_590);
nor U4557 (N_4557,In_935,In_1993);
or U4558 (N_4558,In_555,In_60);
or U4559 (N_4559,In_295,In_1298);
and U4560 (N_4560,In_141,In_1239);
nor U4561 (N_4561,In_490,In_1106);
nand U4562 (N_4562,In_118,In_298);
nor U4563 (N_4563,In_1008,In_400);
nor U4564 (N_4564,In_838,In_599);
nand U4565 (N_4565,In_1440,In_1277);
nor U4566 (N_4566,In_165,In_1768);
nand U4567 (N_4567,In_1779,In_1639);
nor U4568 (N_4568,In_1665,In_386);
xnor U4569 (N_4569,In_347,In_1723);
or U4570 (N_4570,In_1602,In_575);
and U4571 (N_4571,In_1384,In_1714);
and U4572 (N_4572,In_46,In_1341);
or U4573 (N_4573,In_561,In_607);
or U4574 (N_4574,In_916,In_1055);
and U4575 (N_4575,In_545,In_343);
nor U4576 (N_4576,In_641,In_1983);
or U4577 (N_4577,In_1858,In_1115);
and U4578 (N_4578,In_322,In_572);
nand U4579 (N_4579,In_1890,In_1113);
and U4580 (N_4580,In_1198,In_1160);
nor U4581 (N_4581,In_167,In_111);
nor U4582 (N_4582,In_1553,In_12);
nand U4583 (N_4583,In_57,In_708);
or U4584 (N_4584,In_339,In_97);
and U4585 (N_4585,In_766,In_901);
or U4586 (N_4586,In_1353,In_1930);
nor U4587 (N_4587,In_1216,In_1050);
nand U4588 (N_4588,In_1213,In_1992);
nor U4589 (N_4589,In_1518,In_52);
and U4590 (N_4590,In_592,In_1322);
nand U4591 (N_4591,In_1517,In_1546);
nand U4592 (N_4592,In_1561,In_227);
and U4593 (N_4593,In_1945,In_335);
or U4594 (N_4594,In_786,In_1705);
and U4595 (N_4595,In_298,In_1270);
xor U4596 (N_4596,In_1722,In_652);
nand U4597 (N_4597,In_1990,In_1163);
and U4598 (N_4598,In_518,In_1329);
and U4599 (N_4599,In_223,In_1693);
or U4600 (N_4600,In_1127,In_956);
nand U4601 (N_4601,In_1119,In_1069);
nand U4602 (N_4602,In_639,In_1394);
nor U4603 (N_4603,In_1770,In_375);
or U4604 (N_4604,In_1770,In_815);
or U4605 (N_4605,In_1404,In_585);
nor U4606 (N_4606,In_1765,In_1250);
or U4607 (N_4607,In_63,In_419);
nor U4608 (N_4608,In_270,In_1646);
xor U4609 (N_4609,In_229,In_1636);
xor U4610 (N_4610,In_1198,In_321);
nand U4611 (N_4611,In_785,In_1500);
nor U4612 (N_4612,In_741,In_1708);
nor U4613 (N_4613,In_268,In_862);
and U4614 (N_4614,In_1890,In_1891);
nor U4615 (N_4615,In_1169,In_1477);
and U4616 (N_4616,In_674,In_121);
or U4617 (N_4617,In_618,In_1726);
nor U4618 (N_4618,In_1309,In_991);
xor U4619 (N_4619,In_1019,In_1294);
nor U4620 (N_4620,In_545,In_1507);
or U4621 (N_4621,In_912,In_811);
nor U4622 (N_4622,In_1625,In_380);
xnor U4623 (N_4623,In_1580,In_1928);
nor U4624 (N_4624,In_1102,In_726);
and U4625 (N_4625,In_887,In_483);
xnor U4626 (N_4626,In_715,In_33);
nand U4627 (N_4627,In_217,In_1416);
and U4628 (N_4628,In_807,In_677);
nand U4629 (N_4629,In_283,In_374);
nand U4630 (N_4630,In_1816,In_382);
xnor U4631 (N_4631,In_1823,In_223);
and U4632 (N_4632,In_677,In_1877);
nor U4633 (N_4633,In_1701,In_942);
and U4634 (N_4634,In_378,In_1106);
or U4635 (N_4635,In_634,In_1599);
nor U4636 (N_4636,In_676,In_1401);
nor U4637 (N_4637,In_58,In_793);
or U4638 (N_4638,In_704,In_1437);
or U4639 (N_4639,In_640,In_217);
or U4640 (N_4640,In_896,In_148);
nor U4641 (N_4641,In_618,In_100);
and U4642 (N_4642,In_516,In_1743);
and U4643 (N_4643,In_414,In_1251);
and U4644 (N_4644,In_651,In_265);
and U4645 (N_4645,In_762,In_1250);
and U4646 (N_4646,In_372,In_1200);
or U4647 (N_4647,In_934,In_484);
or U4648 (N_4648,In_489,In_1478);
and U4649 (N_4649,In_326,In_724);
nand U4650 (N_4650,In_1042,In_1790);
nand U4651 (N_4651,In_115,In_567);
and U4652 (N_4652,In_1523,In_461);
and U4653 (N_4653,In_308,In_1080);
or U4654 (N_4654,In_1766,In_179);
or U4655 (N_4655,In_563,In_186);
nor U4656 (N_4656,In_1141,In_1812);
nand U4657 (N_4657,In_365,In_1474);
or U4658 (N_4658,In_676,In_529);
and U4659 (N_4659,In_516,In_897);
and U4660 (N_4660,In_1233,In_801);
nor U4661 (N_4661,In_1578,In_637);
or U4662 (N_4662,In_224,In_218);
xor U4663 (N_4663,In_785,In_720);
or U4664 (N_4664,In_860,In_1488);
and U4665 (N_4665,In_1313,In_1730);
and U4666 (N_4666,In_335,In_1017);
or U4667 (N_4667,In_728,In_1507);
nor U4668 (N_4668,In_1050,In_1092);
nor U4669 (N_4669,In_1381,In_420);
or U4670 (N_4670,In_1972,In_1616);
or U4671 (N_4671,In_1891,In_88);
nor U4672 (N_4672,In_576,In_1306);
nand U4673 (N_4673,In_1376,In_1011);
and U4674 (N_4674,In_1421,In_1580);
nand U4675 (N_4675,In_779,In_229);
nand U4676 (N_4676,In_564,In_1572);
or U4677 (N_4677,In_1302,In_1818);
or U4678 (N_4678,In_574,In_182);
or U4679 (N_4679,In_1840,In_1070);
and U4680 (N_4680,In_113,In_345);
or U4681 (N_4681,In_1803,In_1983);
nand U4682 (N_4682,In_683,In_813);
nor U4683 (N_4683,In_577,In_759);
and U4684 (N_4684,In_69,In_1412);
nor U4685 (N_4685,In_166,In_358);
nor U4686 (N_4686,In_734,In_1972);
and U4687 (N_4687,In_247,In_1758);
nor U4688 (N_4688,In_1936,In_304);
xnor U4689 (N_4689,In_893,In_1637);
or U4690 (N_4690,In_877,In_20);
nor U4691 (N_4691,In_373,In_1830);
nor U4692 (N_4692,In_1899,In_802);
nand U4693 (N_4693,In_1604,In_1503);
or U4694 (N_4694,In_984,In_174);
nor U4695 (N_4695,In_662,In_957);
and U4696 (N_4696,In_22,In_869);
nor U4697 (N_4697,In_518,In_719);
xnor U4698 (N_4698,In_871,In_501);
nand U4699 (N_4699,In_653,In_1569);
nor U4700 (N_4700,In_684,In_1412);
nor U4701 (N_4701,In_1668,In_1689);
or U4702 (N_4702,In_610,In_848);
nand U4703 (N_4703,In_940,In_1160);
or U4704 (N_4704,In_954,In_460);
or U4705 (N_4705,In_847,In_152);
xnor U4706 (N_4706,In_1783,In_1265);
or U4707 (N_4707,In_901,In_306);
and U4708 (N_4708,In_265,In_1261);
nand U4709 (N_4709,In_1434,In_663);
nand U4710 (N_4710,In_1631,In_21);
nor U4711 (N_4711,In_1590,In_1369);
or U4712 (N_4712,In_1923,In_779);
nor U4713 (N_4713,In_43,In_1299);
nand U4714 (N_4714,In_851,In_618);
or U4715 (N_4715,In_840,In_182);
and U4716 (N_4716,In_1072,In_1181);
nand U4717 (N_4717,In_590,In_1370);
nand U4718 (N_4718,In_1574,In_1239);
or U4719 (N_4719,In_947,In_438);
nor U4720 (N_4720,In_1177,In_860);
or U4721 (N_4721,In_1464,In_431);
and U4722 (N_4722,In_1930,In_356);
nand U4723 (N_4723,In_662,In_150);
nor U4724 (N_4724,In_629,In_1988);
nor U4725 (N_4725,In_580,In_1597);
and U4726 (N_4726,In_604,In_842);
xnor U4727 (N_4727,In_1987,In_1316);
or U4728 (N_4728,In_398,In_1833);
nor U4729 (N_4729,In_449,In_1134);
nor U4730 (N_4730,In_534,In_76);
nor U4731 (N_4731,In_347,In_1687);
nor U4732 (N_4732,In_801,In_752);
or U4733 (N_4733,In_600,In_1712);
nor U4734 (N_4734,In_162,In_462);
xor U4735 (N_4735,In_282,In_1938);
and U4736 (N_4736,In_277,In_763);
and U4737 (N_4737,In_1685,In_1070);
nor U4738 (N_4738,In_1934,In_1482);
xnor U4739 (N_4739,In_1436,In_288);
nor U4740 (N_4740,In_1126,In_325);
xor U4741 (N_4741,In_1306,In_145);
or U4742 (N_4742,In_1087,In_1874);
nor U4743 (N_4743,In_7,In_1371);
nand U4744 (N_4744,In_1210,In_1520);
nand U4745 (N_4745,In_1865,In_733);
nor U4746 (N_4746,In_1006,In_1998);
or U4747 (N_4747,In_780,In_1422);
nor U4748 (N_4748,In_1676,In_1905);
nor U4749 (N_4749,In_982,In_50);
or U4750 (N_4750,In_461,In_1832);
or U4751 (N_4751,In_864,In_1954);
or U4752 (N_4752,In_1954,In_302);
or U4753 (N_4753,In_725,In_688);
nand U4754 (N_4754,In_1126,In_172);
xnor U4755 (N_4755,In_458,In_1844);
or U4756 (N_4756,In_1115,In_1818);
nand U4757 (N_4757,In_394,In_933);
nand U4758 (N_4758,In_1230,In_1985);
or U4759 (N_4759,In_181,In_908);
and U4760 (N_4760,In_373,In_585);
nor U4761 (N_4761,In_961,In_1303);
and U4762 (N_4762,In_48,In_1433);
and U4763 (N_4763,In_1210,In_434);
nand U4764 (N_4764,In_1481,In_1756);
or U4765 (N_4765,In_1350,In_1762);
nand U4766 (N_4766,In_1830,In_1536);
and U4767 (N_4767,In_1179,In_710);
and U4768 (N_4768,In_221,In_516);
nand U4769 (N_4769,In_721,In_1631);
and U4770 (N_4770,In_521,In_1047);
nand U4771 (N_4771,In_214,In_1616);
nand U4772 (N_4772,In_1842,In_1198);
or U4773 (N_4773,In_1728,In_42);
and U4774 (N_4774,In_1763,In_1261);
or U4775 (N_4775,In_1374,In_1046);
nor U4776 (N_4776,In_509,In_931);
or U4777 (N_4777,In_23,In_1346);
or U4778 (N_4778,In_1238,In_206);
and U4779 (N_4779,In_706,In_951);
and U4780 (N_4780,In_1257,In_450);
and U4781 (N_4781,In_931,In_1275);
xor U4782 (N_4782,In_681,In_378);
and U4783 (N_4783,In_360,In_228);
and U4784 (N_4784,In_1767,In_217);
and U4785 (N_4785,In_1807,In_126);
nor U4786 (N_4786,In_1158,In_1521);
nand U4787 (N_4787,In_873,In_1548);
nand U4788 (N_4788,In_668,In_993);
xor U4789 (N_4789,In_1311,In_366);
and U4790 (N_4790,In_950,In_1368);
and U4791 (N_4791,In_1568,In_1762);
nor U4792 (N_4792,In_1230,In_1009);
nand U4793 (N_4793,In_223,In_1813);
or U4794 (N_4794,In_1305,In_1335);
xor U4795 (N_4795,In_1252,In_614);
or U4796 (N_4796,In_1125,In_623);
nand U4797 (N_4797,In_598,In_1314);
or U4798 (N_4798,In_212,In_840);
xor U4799 (N_4799,In_31,In_90);
or U4800 (N_4800,In_1682,In_1880);
xnor U4801 (N_4801,In_770,In_729);
or U4802 (N_4802,In_864,In_727);
xor U4803 (N_4803,In_1687,In_1501);
and U4804 (N_4804,In_1685,In_81);
and U4805 (N_4805,In_820,In_305);
nand U4806 (N_4806,In_1135,In_81);
and U4807 (N_4807,In_747,In_1034);
nand U4808 (N_4808,In_1269,In_1413);
xnor U4809 (N_4809,In_411,In_1486);
nor U4810 (N_4810,In_1877,In_260);
nor U4811 (N_4811,In_1342,In_943);
and U4812 (N_4812,In_281,In_1022);
and U4813 (N_4813,In_1819,In_1587);
nor U4814 (N_4814,In_1870,In_370);
and U4815 (N_4815,In_1774,In_1561);
nand U4816 (N_4816,In_943,In_429);
nand U4817 (N_4817,In_902,In_435);
nor U4818 (N_4818,In_1845,In_1761);
xnor U4819 (N_4819,In_1950,In_822);
nand U4820 (N_4820,In_979,In_1387);
and U4821 (N_4821,In_1797,In_1692);
or U4822 (N_4822,In_1616,In_1824);
nor U4823 (N_4823,In_845,In_26);
xor U4824 (N_4824,In_1715,In_562);
and U4825 (N_4825,In_810,In_386);
nand U4826 (N_4826,In_902,In_1151);
or U4827 (N_4827,In_258,In_1254);
nand U4828 (N_4828,In_1861,In_982);
nor U4829 (N_4829,In_709,In_391);
xor U4830 (N_4830,In_522,In_1877);
xnor U4831 (N_4831,In_1622,In_918);
nand U4832 (N_4832,In_268,In_1608);
and U4833 (N_4833,In_1192,In_240);
or U4834 (N_4834,In_632,In_845);
nand U4835 (N_4835,In_1708,In_464);
nand U4836 (N_4836,In_1881,In_1861);
and U4837 (N_4837,In_1516,In_1140);
nand U4838 (N_4838,In_1228,In_1779);
nand U4839 (N_4839,In_797,In_1910);
nand U4840 (N_4840,In_511,In_859);
nor U4841 (N_4841,In_1018,In_1053);
or U4842 (N_4842,In_1731,In_959);
or U4843 (N_4843,In_1292,In_273);
and U4844 (N_4844,In_1631,In_1213);
nor U4845 (N_4845,In_349,In_278);
and U4846 (N_4846,In_1571,In_448);
nand U4847 (N_4847,In_932,In_232);
or U4848 (N_4848,In_746,In_1218);
nand U4849 (N_4849,In_123,In_1502);
or U4850 (N_4850,In_1998,In_1396);
xnor U4851 (N_4851,In_1231,In_930);
or U4852 (N_4852,In_604,In_2);
xnor U4853 (N_4853,In_679,In_762);
or U4854 (N_4854,In_1783,In_766);
or U4855 (N_4855,In_85,In_23);
nor U4856 (N_4856,In_386,In_1753);
xnor U4857 (N_4857,In_1647,In_1633);
or U4858 (N_4858,In_263,In_1493);
or U4859 (N_4859,In_248,In_1279);
nor U4860 (N_4860,In_1042,In_1734);
xor U4861 (N_4861,In_1000,In_1239);
and U4862 (N_4862,In_13,In_1204);
nor U4863 (N_4863,In_651,In_904);
nor U4864 (N_4864,In_1570,In_1469);
or U4865 (N_4865,In_267,In_840);
and U4866 (N_4866,In_1444,In_1920);
and U4867 (N_4867,In_1349,In_1924);
nand U4868 (N_4868,In_1755,In_762);
or U4869 (N_4869,In_1555,In_33);
nor U4870 (N_4870,In_1205,In_623);
or U4871 (N_4871,In_1358,In_699);
or U4872 (N_4872,In_448,In_130);
and U4873 (N_4873,In_738,In_787);
or U4874 (N_4874,In_60,In_781);
nor U4875 (N_4875,In_79,In_1530);
or U4876 (N_4876,In_57,In_352);
and U4877 (N_4877,In_1076,In_1399);
nand U4878 (N_4878,In_452,In_930);
and U4879 (N_4879,In_1686,In_703);
or U4880 (N_4880,In_647,In_633);
or U4881 (N_4881,In_270,In_825);
and U4882 (N_4882,In_754,In_944);
xor U4883 (N_4883,In_1331,In_983);
nand U4884 (N_4884,In_1327,In_1424);
nand U4885 (N_4885,In_648,In_237);
xor U4886 (N_4886,In_470,In_148);
and U4887 (N_4887,In_264,In_1907);
and U4888 (N_4888,In_399,In_819);
nand U4889 (N_4889,In_1083,In_1142);
nor U4890 (N_4890,In_1078,In_1782);
nand U4891 (N_4891,In_1911,In_1437);
and U4892 (N_4892,In_1452,In_1427);
nor U4893 (N_4893,In_209,In_627);
and U4894 (N_4894,In_696,In_716);
nor U4895 (N_4895,In_1739,In_1084);
or U4896 (N_4896,In_886,In_138);
nor U4897 (N_4897,In_1296,In_1519);
nor U4898 (N_4898,In_366,In_152);
nand U4899 (N_4899,In_941,In_614);
or U4900 (N_4900,In_1198,In_1576);
nor U4901 (N_4901,In_720,In_46);
nor U4902 (N_4902,In_272,In_205);
and U4903 (N_4903,In_531,In_1385);
and U4904 (N_4904,In_4,In_1808);
or U4905 (N_4905,In_1798,In_1495);
nand U4906 (N_4906,In_51,In_1383);
nor U4907 (N_4907,In_534,In_1182);
or U4908 (N_4908,In_52,In_1145);
or U4909 (N_4909,In_1651,In_840);
and U4910 (N_4910,In_1347,In_764);
nor U4911 (N_4911,In_964,In_522);
nor U4912 (N_4912,In_1113,In_778);
or U4913 (N_4913,In_1392,In_456);
or U4914 (N_4914,In_1475,In_1906);
or U4915 (N_4915,In_916,In_1134);
nand U4916 (N_4916,In_691,In_448);
and U4917 (N_4917,In_751,In_692);
xor U4918 (N_4918,In_587,In_249);
xnor U4919 (N_4919,In_908,In_643);
and U4920 (N_4920,In_1678,In_1493);
xnor U4921 (N_4921,In_1684,In_176);
and U4922 (N_4922,In_1222,In_122);
nor U4923 (N_4923,In_139,In_1591);
and U4924 (N_4924,In_1805,In_26);
xor U4925 (N_4925,In_1186,In_546);
nor U4926 (N_4926,In_998,In_334);
or U4927 (N_4927,In_897,In_52);
or U4928 (N_4928,In_640,In_1765);
nor U4929 (N_4929,In_1973,In_1349);
nand U4930 (N_4930,In_1945,In_342);
nand U4931 (N_4931,In_52,In_1707);
xor U4932 (N_4932,In_219,In_857);
nor U4933 (N_4933,In_1939,In_1454);
xor U4934 (N_4934,In_1092,In_1765);
nor U4935 (N_4935,In_384,In_1474);
or U4936 (N_4936,In_917,In_1982);
nand U4937 (N_4937,In_377,In_1473);
xnor U4938 (N_4938,In_1944,In_1641);
nor U4939 (N_4939,In_453,In_212);
or U4940 (N_4940,In_1079,In_873);
xor U4941 (N_4941,In_1446,In_918);
nand U4942 (N_4942,In_1892,In_556);
and U4943 (N_4943,In_164,In_1049);
nand U4944 (N_4944,In_641,In_35);
nor U4945 (N_4945,In_7,In_1472);
or U4946 (N_4946,In_1982,In_1267);
nand U4947 (N_4947,In_151,In_613);
nand U4948 (N_4948,In_1696,In_1083);
nor U4949 (N_4949,In_943,In_588);
nor U4950 (N_4950,In_712,In_1972);
nand U4951 (N_4951,In_176,In_611);
nand U4952 (N_4952,In_252,In_354);
nor U4953 (N_4953,In_491,In_287);
nand U4954 (N_4954,In_207,In_957);
nand U4955 (N_4955,In_1822,In_399);
nor U4956 (N_4956,In_1681,In_443);
xor U4957 (N_4957,In_1964,In_251);
nand U4958 (N_4958,In_1898,In_1661);
nor U4959 (N_4959,In_773,In_124);
and U4960 (N_4960,In_1807,In_444);
or U4961 (N_4961,In_244,In_383);
and U4962 (N_4962,In_1143,In_1490);
nor U4963 (N_4963,In_755,In_1202);
nand U4964 (N_4964,In_810,In_1724);
or U4965 (N_4965,In_455,In_1995);
nand U4966 (N_4966,In_1768,In_1713);
nand U4967 (N_4967,In_1380,In_233);
xnor U4968 (N_4968,In_1326,In_1271);
nor U4969 (N_4969,In_133,In_259);
nor U4970 (N_4970,In_1156,In_343);
or U4971 (N_4971,In_1639,In_1695);
nand U4972 (N_4972,In_1216,In_1147);
xor U4973 (N_4973,In_251,In_1982);
nor U4974 (N_4974,In_480,In_641);
xnor U4975 (N_4975,In_1261,In_348);
nand U4976 (N_4976,In_410,In_1459);
nor U4977 (N_4977,In_1230,In_1641);
nand U4978 (N_4978,In_1213,In_661);
nor U4979 (N_4979,In_920,In_1467);
xnor U4980 (N_4980,In_1769,In_152);
nand U4981 (N_4981,In_1259,In_1543);
or U4982 (N_4982,In_133,In_1812);
and U4983 (N_4983,In_1037,In_254);
and U4984 (N_4984,In_1375,In_805);
and U4985 (N_4985,In_1279,In_1237);
and U4986 (N_4986,In_1470,In_1336);
and U4987 (N_4987,In_499,In_55);
nor U4988 (N_4988,In_1073,In_619);
nand U4989 (N_4989,In_670,In_1336);
nand U4990 (N_4990,In_1500,In_197);
and U4991 (N_4991,In_2,In_1468);
and U4992 (N_4992,In_83,In_672);
or U4993 (N_4993,In_1322,In_0);
nand U4994 (N_4994,In_1008,In_1530);
nor U4995 (N_4995,In_339,In_896);
and U4996 (N_4996,In_596,In_1326);
nand U4997 (N_4997,In_481,In_1115);
and U4998 (N_4998,In_472,In_1103);
or U4999 (N_4999,In_1139,In_749);
and U5000 (N_5000,N_2071,N_4397);
or U5001 (N_5001,N_1846,N_1580);
and U5002 (N_5002,N_4848,N_481);
or U5003 (N_5003,N_342,N_4745);
nand U5004 (N_5004,N_1543,N_2966);
nor U5005 (N_5005,N_1293,N_1077);
nor U5006 (N_5006,N_492,N_4838);
nor U5007 (N_5007,N_2494,N_1786);
or U5008 (N_5008,N_2160,N_2302);
xnor U5009 (N_5009,N_2876,N_2839);
nor U5010 (N_5010,N_4663,N_1715);
nor U5011 (N_5011,N_530,N_3318);
nand U5012 (N_5012,N_3244,N_4067);
and U5013 (N_5013,N_2848,N_4279);
xor U5014 (N_5014,N_3414,N_3493);
or U5015 (N_5015,N_21,N_732);
or U5016 (N_5016,N_887,N_3246);
or U5017 (N_5017,N_4594,N_979);
and U5018 (N_5018,N_4018,N_1894);
nand U5019 (N_5019,N_1214,N_2522);
and U5020 (N_5020,N_852,N_1874);
or U5021 (N_5021,N_484,N_678);
nand U5022 (N_5022,N_895,N_738);
xor U5023 (N_5023,N_1609,N_3187);
or U5024 (N_5024,N_265,N_646);
or U5025 (N_5025,N_2884,N_4189);
xor U5026 (N_5026,N_3810,N_1112);
and U5027 (N_5027,N_1722,N_2279);
nor U5028 (N_5028,N_64,N_4247);
nor U5029 (N_5029,N_2491,N_1171);
or U5030 (N_5030,N_1016,N_4572);
xnor U5031 (N_5031,N_1213,N_3739);
and U5032 (N_5032,N_3823,N_3879);
nor U5033 (N_5033,N_1931,N_4181);
and U5034 (N_5034,N_2691,N_3293);
or U5035 (N_5035,N_2252,N_1091);
xor U5036 (N_5036,N_313,N_296);
and U5037 (N_5037,N_3849,N_805);
nor U5038 (N_5038,N_1225,N_894);
and U5039 (N_5039,N_3807,N_92);
nor U5040 (N_5040,N_904,N_4358);
or U5041 (N_5041,N_4539,N_4041);
nand U5042 (N_5042,N_1517,N_723);
nand U5043 (N_5043,N_3356,N_2157);
and U5044 (N_5044,N_1992,N_1051);
nand U5045 (N_5045,N_713,N_4007);
and U5046 (N_5046,N_1397,N_1706);
or U5047 (N_5047,N_4778,N_3088);
nand U5048 (N_5048,N_1649,N_3133);
nor U5049 (N_5049,N_4868,N_387);
nor U5050 (N_5050,N_3222,N_185);
nor U5051 (N_5051,N_1446,N_4609);
or U5052 (N_5052,N_4537,N_3421);
nor U5053 (N_5053,N_639,N_90);
nand U5054 (N_5054,N_4031,N_3047);
nor U5055 (N_5055,N_4385,N_3330);
and U5056 (N_5056,N_3142,N_4055);
nor U5057 (N_5057,N_4000,N_2283);
or U5058 (N_5058,N_2878,N_599);
or U5059 (N_5059,N_4200,N_2274);
and U5060 (N_5060,N_2891,N_178);
and U5061 (N_5061,N_2076,N_1210);
and U5062 (N_5062,N_4507,N_2762);
nand U5063 (N_5063,N_4448,N_2168);
nand U5064 (N_5064,N_3043,N_3007);
and U5065 (N_5065,N_2391,N_1761);
nor U5066 (N_5066,N_3144,N_4175);
nor U5067 (N_5067,N_238,N_16);
nor U5068 (N_5068,N_793,N_877);
nand U5069 (N_5069,N_2176,N_3382);
or U5070 (N_5070,N_1119,N_951);
and U5071 (N_5071,N_1848,N_4850);
nor U5072 (N_5072,N_1364,N_3727);
and U5073 (N_5073,N_2204,N_3484);
and U5074 (N_5074,N_4938,N_2575);
xnor U5075 (N_5075,N_1508,N_1297);
or U5076 (N_5076,N_2577,N_4694);
xnor U5077 (N_5077,N_690,N_1177);
nor U5078 (N_5078,N_2368,N_2965);
nor U5079 (N_5079,N_794,N_1962);
and U5080 (N_5080,N_4268,N_2447);
or U5081 (N_5081,N_4015,N_2505);
xnor U5082 (N_5082,N_2899,N_3358);
or U5083 (N_5083,N_3510,N_982);
and U5084 (N_5084,N_2284,N_33);
or U5085 (N_5085,N_2944,N_4080);
nand U5086 (N_5086,N_2515,N_4599);
nor U5087 (N_5087,N_3982,N_1548);
nand U5088 (N_5088,N_1778,N_1680);
nand U5089 (N_5089,N_1861,N_2041);
nor U5090 (N_5090,N_1797,N_1132);
or U5091 (N_5091,N_493,N_916);
and U5092 (N_5092,N_3756,N_883);
nor U5093 (N_5093,N_4008,N_2692);
or U5094 (N_5094,N_4482,N_2195);
and U5095 (N_5095,N_485,N_1940);
nor U5096 (N_5096,N_3277,N_2758);
and U5097 (N_5097,N_548,N_4280);
nand U5098 (N_5098,N_4973,N_2625);
nand U5099 (N_5099,N_4731,N_4050);
nand U5100 (N_5100,N_3126,N_4149);
and U5101 (N_5101,N_661,N_2266);
or U5102 (N_5102,N_176,N_2665);
and U5103 (N_5103,N_4430,N_2904);
nor U5104 (N_5104,N_753,N_366);
or U5105 (N_5105,N_4330,N_1551);
nand U5106 (N_5106,N_1138,N_557);
nor U5107 (N_5107,N_4378,N_4263);
nor U5108 (N_5108,N_1737,N_2148);
or U5109 (N_5109,N_491,N_496);
or U5110 (N_5110,N_174,N_2272);
and U5111 (N_5111,N_3605,N_1445);
nor U5112 (N_5112,N_514,N_1866);
or U5113 (N_5113,N_1929,N_3056);
nand U5114 (N_5114,N_3262,N_2054);
nor U5115 (N_5115,N_2753,N_330);
nor U5116 (N_5116,N_2267,N_98);
nor U5117 (N_5117,N_2450,N_669);
and U5118 (N_5118,N_2591,N_1053);
nand U5119 (N_5119,N_2930,N_3919);
nor U5120 (N_5120,N_349,N_2630);
or U5121 (N_5121,N_2210,N_3641);
or U5122 (N_5122,N_4056,N_2622);
nor U5123 (N_5123,N_4986,N_2580);
nand U5124 (N_5124,N_2261,N_3113);
nor U5125 (N_5125,N_1862,N_1350);
nor U5126 (N_5126,N_4390,N_4554);
and U5127 (N_5127,N_4216,N_329);
and U5128 (N_5128,N_3508,N_4472);
or U5129 (N_5129,N_3909,N_453);
xor U5130 (N_5130,N_4042,N_2962);
nand U5131 (N_5131,N_2896,N_3184);
or U5132 (N_5132,N_1566,N_2241);
or U5133 (N_5133,N_4628,N_3370);
or U5134 (N_5134,N_1329,N_2156);
nor U5135 (N_5135,N_72,N_61);
or U5136 (N_5136,N_889,N_93);
or U5137 (N_5137,N_4260,N_134);
nand U5138 (N_5138,N_4952,N_1174);
and U5139 (N_5139,N_2929,N_4089);
nand U5140 (N_5140,N_2439,N_4436);
or U5141 (N_5141,N_702,N_2420);
nor U5142 (N_5142,N_2513,N_3538);
or U5143 (N_5143,N_4338,N_3865);
xnor U5144 (N_5144,N_928,N_3032);
xor U5145 (N_5145,N_4084,N_766);
or U5146 (N_5146,N_3264,N_3512);
nand U5147 (N_5147,N_4556,N_4934);
xor U5148 (N_5148,N_222,N_2048);
nor U5149 (N_5149,N_3681,N_2928);
or U5150 (N_5150,N_440,N_3939);
and U5151 (N_5151,N_1443,N_912);
nor U5152 (N_5152,N_3403,N_3758);
nor U5153 (N_5153,N_2932,N_3532);
xor U5154 (N_5154,N_107,N_1011);
or U5155 (N_5155,N_328,N_1315);
and U5156 (N_5156,N_223,N_1842);
and U5157 (N_5157,N_4913,N_1414);
and U5158 (N_5158,N_2704,N_3904);
and U5159 (N_5159,N_3416,N_1105);
or U5160 (N_5160,N_3906,N_2178);
and U5161 (N_5161,N_1759,N_1195);
nand U5162 (N_5162,N_716,N_4682);
and U5163 (N_5163,N_1673,N_4037);
xor U5164 (N_5164,N_2804,N_778);
and U5165 (N_5165,N_4760,N_1153);
nand U5166 (N_5166,N_1700,N_2998);
or U5167 (N_5167,N_3520,N_1663);
xnor U5168 (N_5168,N_3721,N_688);
or U5169 (N_5169,N_763,N_685);
nor U5170 (N_5170,N_1512,N_4907);
or U5171 (N_5171,N_2767,N_255);
nor U5172 (N_5172,N_4292,N_1253);
nor U5173 (N_5173,N_1304,N_252);
or U5174 (N_5174,N_3082,N_2280);
and U5175 (N_5175,N_1176,N_1659);
nand U5176 (N_5176,N_124,N_4684);
and U5177 (N_5177,N_3579,N_106);
and U5178 (N_5178,N_1328,N_2258);
nand U5179 (N_5179,N_3519,N_3123);
nor U5180 (N_5180,N_866,N_3655);
and U5181 (N_5181,N_2708,N_4874);
xor U5182 (N_5182,N_1560,N_3443);
nand U5183 (N_5183,N_2816,N_3846);
nor U5184 (N_5184,N_3021,N_551);
nand U5185 (N_5185,N_603,N_1028);
and U5186 (N_5186,N_4066,N_360);
or U5187 (N_5187,N_3434,N_1758);
nand U5188 (N_5188,N_4719,N_1671);
xnor U5189 (N_5189,N_4862,N_2886);
or U5190 (N_5190,N_3192,N_2189);
or U5191 (N_5191,N_2674,N_52);
and U5192 (N_5192,N_869,N_3339);
nand U5193 (N_5193,N_4163,N_2065);
and U5194 (N_5194,N_17,N_3291);
or U5195 (N_5195,N_3881,N_1198);
and U5196 (N_5196,N_377,N_3299);
nor U5197 (N_5197,N_2444,N_500);
or U5198 (N_5198,N_1475,N_1170);
nor U5199 (N_5199,N_4075,N_2217);
nor U5200 (N_5200,N_3576,N_2590);
nand U5201 (N_5201,N_3866,N_1974);
nor U5202 (N_5202,N_3535,N_47);
nand U5203 (N_5203,N_959,N_2012);
and U5204 (N_5204,N_1411,N_3516);
and U5205 (N_5205,N_1074,N_3542);
and U5206 (N_5206,N_2776,N_428);
and U5207 (N_5207,N_526,N_4304);
nor U5208 (N_5208,N_3357,N_1937);
or U5209 (N_5209,N_3303,N_4111);
nand U5210 (N_5210,N_4869,N_987);
or U5211 (N_5211,N_3011,N_2943);
xnor U5212 (N_5212,N_4409,N_1242);
or U5213 (N_5213,N_1157,N_1608);
and U5214 (N_5214,N_1025,N_2564);
nor U5215 (N_5215,N_2750,N_2378);
or U5216 (N_5216,N_239,N_2737);
and U5217 (N_5217,N_1020,N_4708);
or U5218 (N_5218,N_4735,N_1882);
or U5219 (N_5219,N_4846,N_573);
nor U5220 (N_5220,N_1977,N_3102);
and U5221 (N_5221,N_962,N_2990);
nand U5222 (N_5222,N_821,N_282);
and U5223 (N_5223,N_721,N_1597);
or U5224 (N_5224,N_36,N_1793);
nand U5225 (N_5225,N_1779,N_2166);
nand U5226 (N_5226,N_1914,N_3664);
and U5227 (N_5227,N_2655,N_991);
nor U5228 (N_5228,N_1628,N_679);
and U5229 (N_5229,N_3517,N_520);
xnor U5230 (N_5230,N_4927,N_774);
nor U5231 (N_5231,N_2764,N_1622);
nor U5232 (N_5232,N_3350,N_592);
or U5233 (N_5233,N_3136,N_2291);
or U5234 (N_5234,N_3433,N_318);
nand U5235 (N_5235,N_1979,N_4212);
or U5236 (N_5236,N_3861,N_4267);
nand U5237 (N_5237,N_2561,N_2756);
or U5238 (N_5238,N_272,N_4027);
and U5239 (N_5239,N_3966,N_2861);
and U5240 (N_5240,N_1325,N_2187);
nand U5241 (N_5241,N_3341,N_658);
and U5242 (N_5242,N_1924,N_2730);
nor U5243 (N_5243,N_1764,N_849);
nor U5244 (N_5244,N_2104,N_1172);
nor U5245 (N_5245,N_466,N_3023);
and U5246 (N_5246,N_3957,N_1235);
or U5247 (N_5247,N_1535,N_2752);
or U5248 (N_5248,N_3199,N_3111);
xnor U5249 (N_5249,N_3951,N_260);
nor U5250 (N_5250,N_4843,N_1504);
and U5251 (N_5251,N_4053,N_3623);
nor U5252 (N_5252,N_1086,N_1031);
nand U5253 (N_5253,N_2047,N_2094);
xnor U5254 (N_5254,N_1377,N_3014);
and U5255 (N_5255,N_1623,N_1239);
nor U5256 (N_5256,N_3980,N_2654);
and U5257 (N_5257,N_1807,N_3301);
nor U5258 (N_5258,N_4833,N_1431);
nand U5259 (N_5259,N_159,N_4106);
nor U5260 (N_5260,N_1209,N_4389);
nand U5261 (N_5261,N_3566,N_3220);
nand U5262 (N_5262,N_1744,N_192);
or U5263 (N_5263,N_2853,N_4286);
nor U5264 (N_5264,N_4820,N_970);
and U5265 (N_5265,N_1143,N_2480);
and U5266 (N_5266,N_1194,N_950);
or U5267 (N_5267,N_668,N_3630);
and U5268 (N_5268,N_4231,N_1173);
nor U5269 (N_5269,N_2374,N_2710);
nor U5270 (N_5270,N_4091,N_352);
nand U5271 (N_5271,N_3560,N_795);
nor U5272 (N_5272,N_459,N_86);
and U5273 (N_5273,N_4418,N_2285);
nand U5274 (N_5274,N_4151,N_4196);
nand U5275 (N_5275,N_335,N_2954);
or U5276 (N_5276,N_1524,N_2511);
nand U5277 (N_5277,N_4650,N_2842);
nor U5278 (N_5278,N_3698,N_2413);
xor U5279 (N_5279,N_762,N_3811);
and U5280 (N_5280,N_2847,N_3009);
nand U5281 (N_5281,N_473,N_2989);
nand U5282 (N_5282,N_1252,N_1741);
nand U5283 (N_5283,N_4514,N_1952);
and U5284 (N_5284,N_3680,N_1332);
and U5285 (N_5285,N_2091,N_2733);
and U5286 (N_5286,N_2735,N_3965);
nand U5287 (N_5287,N_2819,N_1349);
and U5288 (N_5288,N_3294,N_1326);
nand U5289 (N_5289,N_4328,N_1234);
nor U5290 (N_5290,N_1573,N_1709);
or U5291 (N_5291,N_3628,N_399);
and U5292 (N_5292,N_1955,N_2489);
xor U5293 (N_5293,N_60,N_731);
nand U5294 (N_5294,N_4690,N_2530);
and U5295 (N_5295,N_3608,N_1830);
or U5296 (N_5296,N_4699,N_3798);
nand U5297 (N_5297,N_1643,N_3132);
or U5298 (N_5298,N_4274,N_3027);
nor U5299 (N_5299,N_2974,N_3254);
or U5300 (N_5300,N_553,N_1228);
xor U5301 (N_5301,N_4816,N_4798);
nor U5302 (N_5302,N_524,N_2873);
or U5303 (N_5303,N_1685,N_2020);
or U5304 (N_5304,N_1481,N_433);
or U5305 (N_5305,N_1531,N_4542);
xnor U5306 (N_5306,N_376,N_1688);
and U5307 (N_5307,N_4481,N_4256);
xor U5308 (N_5308,N_2823,N_1059);
nor U5309 (N_5309,N_4275,N_3033);
and U5310 (N_5310,N_3208,N_882);
or U5311 (N_5311,N_1571,N_2508);
xor U5312 (N_5312,N_1405,N_784);
xor U5313 (N_5313,N_2996,N_4533);
and U5314 (N_5314,N_944,N_1787);
or U5315 (N_5315,N_3168,N_4179);
nand U5316 (N_5316,N_3494,N_4425);
nor U5317 (N_5317,N_2199,N_4380);
or U5318 (N_5318,N_2152,N_1676);
nand U5319 (N_5319,N_1,N_1092);
xnor U5320 (N_5320,N_2414,N_2438);
nor U5321 (N_5321,N_1220,N_2820);
xor U5322 (N_5322,N_2544,N_3381);
nand U5323 (N_5323,N_3828,N_2009);
nor U5324 (N_5324,N_3467,N_3896);
nand U5325 (N_5325,N_3961,N_1054);
and U5326 (N_5326,N_2402,N_123);
or U5327 (N_5327,N_1868,N_2607);
and U5328 (N_5328,N_2711,N_1378);
and U5329 (N_5329,N_1283,N_943);
nand U5330 (N_5330,N_1646,N_4184);
xor U5331 (N_5331,N_2549,N_1627);
nor U5332 (N_5332,N_604,N_4616);
xnor U5333 (N_5333,N_3352,N_2229);
nor U5334 (N_5334,N_2163,N_1229);
and U5335 (N_5335,N_990,N_1544);
nand U5336 (N_5336,N_3448,N_3633);
and U5337 (N_5337,N_2906,N_4800);
nor U5338 (N_5338,N_546,N_2595);
or U5339 (N_5339,N_129,N_2358);
and U5340 (N_5340,N_2640,N_1746);
or U5341 (N_5341,N_43,N_3120);
or U5342 (N_5342,N_3504,N_2782);
or U5343 (N_5343,N_4023,N_615);
nand U5344 (N_5344,N_2066,N_735);
nand U5345 (N_5345,N_2526,N_1907);
nand U5346 (N_5346,N_2507,N_2850);
nand U5347 (N_5347,N_475,N_4432);
or U5348 (N_5348,N_3789,N_2614);
nand U5349 (N_5349,N_809,N_4736);
or U5350 (N_5350,N_3592,N_1030);
or U5351 (N_5351,N_4815,N_4420);
or U5352 (N_5352,N_3976,N_51);
and U5353 (N_5353,N_4667,N_1191);
nor U5354 (N_5354,N_4717,N_644);
or U5355 (N_5355,N_300,N_2723);
nor U5356 (N_5356,N_1811,N_2393);
nor U5357 (N_5357,N_4543,N_3039);
or U5358 (N_5358,N_4152,N_4924);
and U5359 (N_5359,N_1975,N_280);
nor U5360 (N_5360,N_4364,N_1612);
nand U5361 (N_5361,N_1376,N_2275);
and U5362 (N_5362,N_1389,N_4227);
and U5363 (N_5363,N_3938,N_2572);
nand U5364 (N_5364,N_4474,N_3999);
nand U5365 (N_5365,N_2372,N_4326);
and U5366 (N_5366,N_4726,N_933);
and U5367 (N_5367,N_1547,N_2308);
and U5368 (N_5368,N_2798,N_3327);
or U5369 (N_5369,N_528,N_100);
nand U5370 (N_5370,N_1967,N_1873);
or U5371 (N_5371,N_3872,N_243);
nor U5372 (N_5372,N_2881,N_2057);
nor U5373 (N_5373,N_2390,N_1179);
nand U5374 (N_5374,N_257,N_2821);
nor U5375 (N_5375,N_1614,N_631);
and U5376 (N_5376,N_4153,N_4547);
nand U5377 (N_5377,N_1262,N_1367);
nand U5378 (N_5378,N_3243,N_4693);
or U5379 (N_5379,N_2942,N_2858);
nor U5380 (N_5380,N_1447,N_2073);
nand U5381 (N_5381,N_3239,N_3114);
and U5382 (N_5382,N_3620,N_606);
or U5383 (N_5383,N_2589,N_1841);
nand U5384 (N_5384,N_836,N_523);
and U5385 (N_5385,N_39,N_2827);
nor U5386 (N_5386,N_3321,N_2060);
and U5387 (N_5387,N_4947,N_3399);
xor U5388 (N_5388,N_323,N_4320);
or U5389 (N_5389,N_594,N_2791);
nand U5390 (N_5390,N_2338,N_4264);
nor U5391 (N_5391,N_4306,N_297);
nor U5392 (N_5392,N_2901,N_4112);
and U5393 (N_5393,N_146,N_4413);
or U5394 (N_5394,N_3745,N_4892);
or U5395 (N_5395,N_2290,N_1847);
xor U5396 (N_5396,N_2602,N_911);
or U5397 (N_5397,N_4787,N_2112);
and U5398 (N_5398,N_2613,N_2101);
or U5399 (N_5399,N_3559,N_4128);
or U5400 (N_5400,N_2606,N_4764);
or U5401 (N_5401,N_2574,N_2181);
xor U5402 (N_5402,N_2637,N_256);
nand U5403 (N_5403,N_3224,N_2880);
or U5404 (N_5404,N_755,N_2223);
xnor U5405 (N_5405,N_182,N_3479);
nand U5406 (N_5406,N_1027,N_346);
nor U5407 (N_5407,N_1392,N_4329);
or U5408 (N_5408,N_4435,N_4520);
nor U5409 (N_5409,N_609,N_3128);
nand U5410 (N_5410,N_2656,N_1887);
nand U5411 (N_5411,N_4315,N_4896);
nand U5412 (N_5412,N_204,N_1363);
and U5413 (N_5413,N_3840,N_789);
nor U5414 (N_5414,N_2330,N_1561);
nand U5415 (N_5415,N_1660,N_4174);
and U5416 (N_5416,N_1985,N_544);
or U5417 (N_5417,N_3549,N_1775);
nor U5418 (N_5418,N_3127,N_3492);
nor U5419 (N_5419,N_874,N_3932);
nor U5420 (N_5420,N_3635,N_1564);
nand U5421 (N_5421,N_810,N_2231);
nor U5422 (N_5422,N_2714,N_2153);
xnor U5423 (N_5423,N_3986,N_4394);
nor U5424 (N_5424,N_2927,N_1558);
nand U5425 (N_5425,N_2300,N_3686);
nand U5426 (N_5426,N_2415,N_1581);
nor U5427 (N_5427,N_435,N_2978);
nand U5428 (N_5428,N_4297,N_1464);
nor U5429 (N_5429,N_3835,N_4826);
or U5430 (N_5430,N_3310,N_3086);
or U5431 (N_5431,N_4071,N_455);
xnor U5432 (N_5432,N_2785,N_1279);
nand U5433 (N_5433,N_2545,N_3972);
and U5434 (N_5434,N_4573,N_101);
nand U5435 (N_5435,N_4352,N_1870);
or U5436 (N_5436,N_3445,N_1617);
or U5437 (N_5437,N_456,N_4747);
and U5438 (N_5438,N_1588,N_2844);
or U5439 (N_5439,N_3060,N_2409);
or U5440 (N_5440,N_3665,N_2841);
or U5441 (N_5441,N_817,N_3687);
xnor U5442 (N_5442,N_3984,N_4950);
nor U5443 (N_5443,N_4853,N_1653);
nand U5444 (N_5444,N_1259,N_4489);
nor U5445 (N_5445,N_4376,N_3129);
xor U5446 (N_5446,N_4491,N_4598);
nand U5447 (N_5447,N_4773,N_2395);
or U5448 (N_5448,N_2198,N_1875);
nand U5449 (N_5449,N_152,N_4351);
nand U5450 (N_5450,N_541,N_3697);
nor U5451 (N_5451,N_2225,N_1600);
or U5452 (N_5452,N_2509,N_474);
or U5453 (N_5453,N_35,N_3019);
nor U5454 (N_5454,N_1904,N_1347);
nor U5455 (N_5455,N_4444,N_1060);
or U5456 (N_5456,N_4642,N_2812);
and U5457 (N_5457,N_1274,N_2038);
and U5458 (N_5458,N_2578,N_1125);
or U5459 (N_5459,N_1458,N_1452);
or U5460 (N_5460,N_992,N_4508);
and U5461 (N_5461,N_2611,N_1750);
nor U5462 (N_5462,N_4725,N_3631);
nor U5463 (N_5463,N_3273,N_830);
and U5464 (N_5464,N_3931,N_162);
and U5465 (N_5465,N_4878,N_550);
and U5466 (N_5466,N_1169,N_3545);
and U5467 (N_5467,N_2011,N_1034);
xor U5468 (N_5468,N_4946,N_3831);
nand U5469 (N_5469,N_1287,N_3118);
and U5470 (N_5470,N_2389,N_3981);
and U5471 (N_5471,N_2803,N_1751);
and U5472 (N_5472,N_3695,N_3228);
or U5473 (N_5473,N_4812,N_2641);
xnor U5474 (N_5474,N_655,N_2158);
and U5475 (N_5475,N_785,N_4570);
nor U5476 (N_5476,N_2353,N_4225);
and U5477 (N_5477,N_4829,N_1017);
or U5478 (N_5478,N_2422,N_1386);
and U5479 (N_5479,N_4568,N_3042);
nand U5480 (N_5480,N_4632,N_3511);
nor U5481 (N_5481,N_863,N_156);
nor U5482 (N_5482,N_4377,N_4847);
nand U5483 (N_5483,N_3718,N_1845);
xnor U5484 (N_5484,N_3107,N_23);
nand U5485 (N_5485,N_3567,N_3477);
or U5486 (N_5486,N_2986,N_2893);
and U5487 (N_5487,N_3200,N_3441);
and U5488 (N_5488,N_2396,N_3967);
nor U5489 (N_5489,N_2793,N_940);
nor U5490 (N_5490,N_46,N_4269);
nor U5491 (N_5491,N_2155,N_2994);
nand U5492 (N_5492,N_1007,N_2727);
nand U5493 (N_5493,N_2428,N_4375);
nor U5494 (N_5494,N_3376,N_2565);
nor U5495 (N_5495,N_1886,N_1471);
nor U5496 (N_5496,N_2007,N_2492);
xnor U5497 (N_5497,N_1880,N_2242);
nor U5498 (N_5498,N_1231,N_2837);
and U5499 (N_5499,N_4503,N_2889);
nor U5500 (N_5500,N_4550,N_1040);
nand U5501 (N_5501,N_2119,N_4318);
nand U5502 (N_5502,N_3,N_3805);
or U5503 (N_5503,N_315,N_1161);
or U5504 (N_5504,N_4365,N_2695);
nand U5505 (N_5505,N_2616,N_4388);
nor U5506 (N_5506,N_1439,N_3730);
and U5507 (N_5507,N_891,N_3689);
and U5508 (N_5508,N_258,N_1805);
nor U5509 (N_5509,N_2669,N_783);
nand U5510 (N_5510,N_2035,N_3780);
nand U5511 (N_5511,N_2352,N_1047);
nor U5512 (N_5512,N_4257,N_4794);
or U5513 (N_5513,N_127,N_4500);
nor U5514 (N_5514,N_2021,N_571);
or U5515 (N_5515,N_2581,N_3112);
or U5516 (N_5516,N_749,N_1144);
or U5517 (N_5517,N_4767,N_1549);
xor U5518 (N_5518,N_3912,N_2317);
or U5519 (N_5519,N_2096,N_4064);
xor U5520 (N_5520,N_3505,N_1897);
nor U5521 (N_5521,N_3052,N_3736);
nand U5522 (N_5522,N_4334,N_2310);
xnor U5523 (N_5523,N_2594,N_1237);
nand U5524 (N_5524,N_838,N_4368);
nor U5525 (N_5525,N_408,N_1180);
nand U5526 (N_5526,N_1240,N_611);
nor U5527 (N_5527,N_1920,N_1592);
nand U5528 (N_5528,N_4655,N_4856);
or U5529 (N_5529,N_2760,N_2008);
and U5530 (N_5530,N_2462,N_137);
and U5531 (N_5531,N_2754,N_3279);
nand U5532 (N_5532,N_3252,N_1067);
xnor U5533 (N_5533,N_325,N_42);
and U5534 (N_5534,N_1356,N_2835);
or U5535 (N_5535,N_3958,N_872);
nand U5536 (N_5536,N_4929,N_4631);
or U5537 (N_5537,N_4587,N_2945);
or U5538 (N_5538,N_3474,N_1533);
or U5539 (N_5539,N_4811,N_2672);
nand U5540 (N_5540,N_3284,N_216);
nor U5541 (N_5541,N_4047,N_627);
xor U5542 (N_5542,N_3365,N_2551);
and U5543 (N_5543,N_2934,N_291);
xor U5544 (N_5544,N_1440,N_170);
and U5545 (N_5545,N_4545,N_4440);
nor U5546 (N_5546,N_3160,N_490);
nand U5547 (N_5547,N_4635,N_3234);
nor U5548 (N_5548,N_4958,N_1619);
nor U5549 (N_5549,N_4657,N_126);
nor U5550 (N_5550,N_4917,N_4975);
xor U5551 (N_5551,N_3034,N_831);
nand U5552 (N_5552,N_3833,N_4859);
or U5553 (N_5553,N_4697,N_498);
or U5554 (N_5554,N_2221,N_2787);
and U5555 (N_5555,N_3459,N_0);
or U5556 (N_5556,N_230,N_3922);
nand U5557 (N_5557,N_3719,N_2133);
or U5558 (N_5558,N_4093,N_2766);
and U5559 (N_5559,N_3953,N_3994);
nor U5560 (N_5560,N_3629,N_3764);
or U5561 (N_5561,N_1090,N_1233);
nor U5562 (N_5562,N_4741,N_1681);
or U5563 (N_5563,N_1745,N_1365);
and U5564 (N_5564,N_2180,N_3159);
nand U5565 (N_5565,N_4224,N_3067);
nand U5566 (N_5566,N_741,N_2362);
nand U5567 (N_5567,N_1410,N_2397);
and U5568 (N_5568,N_4516,N_3152);
nor U5569 (N_5569,N_3073,N_30);
or U5570 (N_5570,N_2755,N_1522);
or U5571 (N_5571,N_3379,N_3525);
nand U5572 (N_5572,N_2288,N_2465);
nor U5573 (N_5573,N_2829,N_4442);
nand U5574 (N_5574,N_2859,N_4701);
nor U5575 (N_5575,N_476,N_1124);
nand U5576 (N_5576,N_2681,N_1687);
and U5577 (N_5577,N_2446,N_2087);
or U5578 (N_5578,N_2468,N_2140);
or U5579 (N_5579,N_3170,N_4678);
and U5580 (N_5580,N_1012,N_4981);
nor U5581 (N_5581,N_483,N_4670);
and U5582 (N_5582,N_3457,N_3647);
nand U5583 (N_5583,N_2024,N_233);
or U5584 (N_5584,N_3900,N_2874);
or U5585 (N_5585,N_3729,N_719);
nand U5586 (N_5586,N_2722,N_1110);
xnor U5587 (N_5587,N_3225,N_1383);
nor U5588 (N_5588,N_4781,N_988);
nor U5589 (N_5589,N_1678,N_922);
and U5590 (N_5590,N_1918,N_3640);
or U5591 (N_5591,N_286,N_3563);
or U5592 (N_5592,N_2110,N_2851);
nor U5593 (N_5593,N_3916,N_2629);
nand U5594 (N_5594,N_4190,N_1528);
and U5595 (N_5595,N_4202,N_4531);
and U5596 (N_5596,N_429,N_121);
nand U5597 (N_5597,N_736,N_3911);
nor U5598 (N_5598,N_3028,N_2271);
nor U5599 (N_5599,N_3097,N_3400);
nor U5600 (N_5600,N_4087,N_1721);
and U5601 (N_5601,N_2502,N_1344);
nand U5602 (N_5602,N_2603,N_2650);
and U5603 (N_5603,N_3612,N_1461);
and U5604 (N_5604,N_1728,N_1545);
and U5605 (N_5605,N_84,N_1441);
and U5606 (N_5606,N_1435,N_1714);
nand U5607 (N_5607,N_4817,N_2124);
and U5608 (N_5608,N_4369,N_4169);
nand U5609 (N_5609,N_3308,N_777);
nor U5610 (N_5610,N_2437,N_4459);
nor U5611 (N_5611,N_4965,N_3547);
and U5612 (N_5612,N_3012,N_4894);
nand U5613 (N_5613,N_4423,N_3808);
nor U5614 (N_5614,N_2014,N_4831);
or U5615 (N_5615,N_1296,N_3838);
and U5616 (N_5616,N_2405,N_3733);
nor U5617 (N_5617,N_4998,N_3240);
nand U5618 (N_5618,N_919,N_513);
nor U5619 (N_5619,N_3925,N_1419);
nand U5620 (N_5620,N_4845,N_4569);
and U5621 (N_5621,N_3848,N_1944);
or U5622 (N_5622,N_4808,N_600);
nor U5623 (N_5623,N_3354,N_197);
or U5624 (N_5624,N_3929,N_3531);
nor U5625 (N_5625,N_1205,N_1416);
nor U5626 (N_5626,N_3749,N_326);
nand U5627 (N_5627,N_2908,N_2618);
and U5628 (N_5628,N_1695,N_24);
or U5629 (N_5629,N_2486,N_800);
nor U5630 (N_5630,N_1217,N_3177);
and U5631 (N_5631,N_4393,N_2418);
or U5632 (N_5632,N_3219,N_4766);
and U5633 (N_5633,N_1388,N_2089);
nor U5634 (N_5634,N_1485,N_1345);
nor U5635 (N_5635,N_3461,N_3431);
nand U5636 (N_5636,N_198,N_1661);
nor U5637 (N_5637,N_19,N_2277);
nand U5638 (N_5638,N_3117,N_744);
and U5639 (N_5639,N_1605,N_210);
nor U5640 (N_5640,N_1518,N_1361);
nand U5641 (N_5641,N_4779,N_3776);
nor U5642 (N_5642,N_4830,N_3820);
xor U5643 (N_5643,N_4367,N_1506);
nor U5644 (N_5644,N_2537,N_4526);
and U5645 (N_5645,N_3338,N_1334);
xor U5646 (N_5646,N_3794,N_3533);
or U5647 (N_5647,N_472,N_1683);
or U5648 (N_5648,N_2001,N_4252);
and U5649 (N_5649,N_386,N_3229);
nand U5650 (N_5650,N_2512,N_3008);
or U5651 (N_5651,N_1703,N_2293);
nor U5652 (N_5652,N_3070,N_3393);
nand U5653 (N_5653,N_4502,N_2686);
and U5654 (N_5654,N_4399,N_3218);
nand U5655 (N_5655,N_930,N_1822);
nor U5656 (N_5656,N_4198,N_2729);
and U5657 (N_5657,N_2678,N_4422);
nand U5658 (N_5658,N_2987,N_3543);
nor U5659 (N_5659,N_4470,N_692);
or U5660 (N_5660,N_3439,N_4158);
or U5661 (N_5661,N_3137,N_2458);
or U5662 (N_5662,N_2624,N_3332);
nor U5663 (N_5663,N_3387,N_3134);
nor U5664 (N_5664,N_317,N_4221);
or U5665 (N_5665,N_3935,N_1099);
or U5666 (N_5666,N_2188,N_4032);
xnor U5667 (N_5667,N_2740,N_1407);
xnor U5668 (N_5668,N_1883,N_4914);
or U5669 (N_5669,N_3369,N_4461);
or U5670 (N_5670,N_1465,N_4928);
nor U5671 (N_5671,N_1483,N_2312);
xnor U5672 (N_5672,N_1765,N_4123);
or U5673 (N_5673,N_1820,N_2619);
nor U5674 (N_5674,N_3139,N_4649);
nand U5675 (N_5675,N_2456,N_4121);
nor U5676 (N_5676,N_1829,N_1819);
or U5677 (N_5677,N_2097,N_4108);
nor U5678 (N_5678,N_3713,N_166);
or U5679 (N_5679,N_740,N_3478);
nor U5680 (N_5680,N_3205,N_1359);
nor U5681 (N_5681,N_95,N_2126);
and U5682 (N_5682,N_799,N_4879);
or U5683 (N_5683,N_1973,N_1519);
xnor U5684 (N_5684,N_4824,N_2318);
and U5685 (N_5685,N_507,N_2424);
or U5686 (N_5686,N_4925,N_3526);
and U5687 (N_5687,N_724,N_3195);
and U5688 (N_5688,N_1831,N_1082);
xor U5689 (N_5689,N_3905,N_4722);
nand U5690 (N_5690,N_2497,N_3682);
xnor U5691 (N_5691,N_649,N_3515);
xnor U5692 (N_5692,N_2554,N_215);
and U5693 (N_5693,N_353,N_1833);
and U5694 (N_5694,N_3684,N_2751);
xnor U5695 (N_5695,N_4206,N_1712);
xor U5696 (N_5696,N_3973,N_1199);
nor U5697 (N_5697,N_4792,N_2324);
and U5698 (N_5698,N_3410,N_518);
nand U5699 (N_5699,N_3261,N_955);
nand U5700 (N_5700,N_2197,N_920);
nor U5701 (N_5701,N_4211,N_4881);
and U5702 (N_5702,N_4076,N_1792);
or U5703 (N_5703,N_3882,N_1804);
nor U5704 (N_5704,N_923,N_1263);
xor U5705 (N_5705,N_1008,N_752);
or U5706 (N_5706,N_1454,N_3748);
and U5707 (N_5707,N_4937,N_4737);
nand U5708 (N_5708,N_4234,N_4723);
nor U5709 (N_5709,N_2963,N_2863);
nand U5710 (N_5710,N_1154,N_589);
and U5711 (N_5711,N_2958,N_947);
or U5712 (N_5712,N_3162,N_3452);
and U5713 (N_5713,N_2540,N_1720);
or U5714 (N_5714,N_4501,N_1269);
xnor U5715 (N_5715,N_2442,N_4178);
nor U5716 (N_5716,N_539,N_1885);
or U5717 (N_5717,N_2067,N_1651);
or U5718 (N_5718,N_67,N_967);
or U5719 (N_5719,N_3180,N_3489);
or U5720 (N_5720,N_2170,N_2081);
nand U5721 (N_5721,N_1893,N_70);
and U5722 (N_5722,N_2196,N_2682);
xnor U5723 (N_5723,N_4104,N_1254);
xor U5724 (N_5724,N_3844,N_4733);
nand U5725 (N_5725,N_3143,N_3245);
and U5726 (N_5726,N_2202,N_841);
and U5727 (N_5727,N_899,N_4113);
and U5728 (N_5728,N_1800,N_2778);
and U5729 (N_5729,N_4691,N_1479);
or U5730 (N_5730,N_105,N_2765);
nor U5731 (N_5731,N_4715,N_660);
nor U5732 (N_5732,N_4475,N_1286);
nand U5733 (N_5733,N_4494,N_4827);
or U5734 (N_5734,N_2918,N_3890);
xnor U5735 (N_5735,N_4777,N_1003);
nand U5736 (N_5736,N_4517,N_537);
nand U5737 (N_5737,N_1756,N_707);
or U5738 (N_5738,N_4659,N_827);
nor U5739 (N_5739,N_3423,N_4322);
nand U5740 (N_5740,N_357,N_2404);
and U5741 (N_5741,N_2287,N_1064);
and U5742 (N_5742,N_3606,N_3472);
nand U5743 (N_5743,N_4916,N_4966);
nor U5744 (N_5744,N_3071,N_402);
or U5745 (N_5745,N_2980,N_1667);
nor U5746 (N_5746,N_141,N_2072);
nand U5747 (N_5747,N_1537,N_4382);
nor U5748 (N_5748,N_2015,N_2969);
or U5749 (N_5749,N_4317,N_2685);
nand U5750 (N_5750,N_1631,N_3743);
and U5751 (N_5751,N_4450,N_4945);
or U5752 (N_5752,N_4012,N_1311);
and U5753 (N_5753,N_4528,N_3425);
and U5754 (N_5754,N_142,N_3903);
or U5755 (N_5755,N_2772,N_2728);
and U5756 (N_5756,N_253,N_1836);
and U5757 (N_5757,N_1682,N_4386);
nor U5758 (N_5758,N_250,N_1050);
xnor U5759 (N_5759,N_3928,N_2323);
or U5760 (N_5760,N_3232,N_3600);
xor U5761 (N_5761,N_2913,N_2843);
and U5762 (N_5762,N_818,N_2218);
and U5763 (N_5763,N_3038,N_2488);
nor U5764 (N_5764,N_1585,N_2316);
and U5765 (N_5765,N_547,N_512);
nand U5766 (N_5766,N_4643,N_1930);
or U5767 (N_5767,N_2547,N_212);
and U5768 (N_5768,N_4170,N_1488);
or U5769 (N_5769,N_254,N_4751);
nor U5770 (N_5770,N_1859,N_213);
nor U5771 (N_5771,N_2870,N_562);
xnor U5772 (N_5772,N_1236,N_245);
nand U5773 (N_5773,N_2626,N_1035);
xnor U5774 (N_5774,N_148,N_4464);
nor U5775 (N_5775,N_4930,N_4654);
and U5776 (N_5776,N_3814,N_2260);
or U5777 (N_5777,N_4828,N_3757);
and U5778 (N_5778,N_1360,N_902);
nor U5779 (N_5779,N_698,N_1593);
or U5780 (N_5780,N_284,N_2933);
and U5781 (N_5781,N_4939,N_316);
nand U5782 (N_5782,N_2448,N_2115);
nor U5783 (N_5783,N_438,N_4707);
or U5784 (N_5784,N_4797,N_4834);
xnor U5785 (N_5785,N_1155,N_773);
nor U5786 (N_5786,N_2805,N_1318);
and U5787 (N_5787,N_2387,N_2777);
nand U5788 (N_5788,N_1969,N_1532);
or U5789 (N_5789,N_1539,N_3089);
nand U5790 (N_5790,N_2745,N_3394);
or U5791 (N_5791,N_1965,N_4744);
nand U5792 (N_5792,N_359,N_791);
nand U5793 (N_5793,N_4126,N_69);
and U5794 (N_5794,N_3658,N_1999);
and U5795 (N_5795,N_351,N_4085);
and U5796 (N_5796,N_2371,N_1498);
and U5797 (N_5797,N_3728,N_1601);
and U5798 (N_5798,N_931,N_140);
nand U5799 (N_5799,N_343,N_1557);
or U5800 (N_5800,N_2142,N_2278);
nand U5801 (N_5801,N_1158,N_914);
xor U5802 (N_5802,N_3621,N_1579);
nand U5803 (N_5803,N_3875,N_2083);
nand U5804 (N_5804,N_4255,N_1939);
xnor U5805 (N_5805,N_823,N_3215);
nor U5806 (N_5806,N_3969,N_2172);
or U5807 (N_5807,N_764,N_4361);
nor U5808 (N_5808,N_3233,N_1832);
nand U5809 (N_5809,N_1226,N_3979);
or U5810 (N_5810,N_120,N_4384);
or U5811 (N_5811,N_1768,N_2106);
and U5812 (N_5812,N_704,N_2715);
and U5813 (N_5813,N_391,N_3722);
and U5814 (N_5814,N_1338,N_1986);
or U5815 (N_5815,N_3213,N_4486);
or U5816 (N_5816,N_3589,N_2905);
nand U5817 (N_5817,N_2524,N_3701);
nor U5818 (N_5818,N_1207,N_3417);
xnor U5819 (N_5819,N_3570,N_1806);
or U5820 (N_5820,N_3275,N_4220);
and U5821 (N_5821,N_1062,N_3197);
nand U5822 (N_5822,N_502,N_2634);
xor U5823 (N_5823,N_2085,N_2599);
nor U5824 (N_5824,N_1818,N_2451);
nand U5825 (N_5825,N_3300,N_154);
or U5826 (N_5826,N_1844,N_2852);
nor U5827 (N_5827,N_648,N_2705);
xor U5828 (N_5828,N_613,N_18);
nor U5829 (N_5829,N_4045,N_770);
or U5830 (N_5830,N_4003,N_4611);
nor U5831 (N_5831,N_78,N_853);
or U5832 (N_5832,N_3242,N_2212);
or U5833 (N_5833,N_4086,N_269);
nand U5834 (N_5834,N_3314,N_1096);
nor U5835 (N_5835,N_3305,N_4465);
nor U5836 (N_5836,N_2800,N_2113);
or U5837 (N_5837,N_80,N_3770);
or U5838 (N_5838,N_1903,N_1669);
nor U5839 (N_5839,N_1625,N_281);
nand U5840 (N_5840,N_4120,N_3346);
or U5841 (N_5841,N_2457,N_4312);
and U5842 (N_5842,N_2294,N_3059);
or U5843 (N_5843,N_3853,N_828);
and U5844 (N_5844,N_1038,N_3573);
nand U5845 (N_5845,N_385,N_1654);
nand U5846 (N_5846,N_3288,N_4905);
or U5847 (N_5847,N_1372,N_2584);
and U5848 (N_5848,N_671,N_3720);
nand U5849 (N_5849,N_3883,N_4316);
nand U5850 (N_5850,N_403,N_1708);
nor U5851 (N_5851,N_2167,N_2721);
and U5852 (N_5852,N_3652,N_1736);
nand U5853 (N_5853,N_595,N_4872);
nor U5854 (N_5854,N_382,N_2660);
and U5855 (N_5855,N_4984,N_1648);
nor U5856 (N_5856,N_2566,N_1291);
and U5857 (N_5857,N_1570,N_1988);
or U5858 (N_5858,N_2445,N_2327);
or U5859 (N_5859,N_714,N_1621);
nand U5860 (N_5860,N_2548,N_1686);
or U5861 (N_5861,N_4983,N_2898);
nor U5862 (N_5862,N_1295,N_839);
and U5863 (N_5863,N_4201,N_3380);
nor U5864 (N_5864,N_2909,N_4176);
nand U5865 (N_5865,N_2757,N_4566);
nor U5866 (N_5866,N_3788,N_4530);
or U5867 (N_5867,N_4861,N_4783);
or U5868 (N_5868,N_2449,N_1029);
xor U5869 (N_5869,N_581,N_4070);
nand U5870 (N_5870,N_426,N_276);
and U5871 (N_5871,N_3773,N_2175);
nand U5872 (N_5872,N_1004,N_591);
nor U5873 (N_5873,N_3391,N_3201);
nand U5874 (N_5874,N_1121,N_4496);
and U5875 (N_5875,N_1324,N_3292);
or U5876 (N_5876,N_3761,N_3590);
nand U5877 (N_5877,N_4029,N_290);
and U5878 (N_5878,N_3654,N_1642);
or U5879 (N_5879,N_2407,N_1635);
xnor U5880 (N_5880,N_1436,N_3022);
and U5881 (N_5881,N_708,N_1908);
and U5882 (N_5882,N_4685,N_516);
or U5883 (N_5883,N_2895,N_4090);
or U5884 (N_5884,N_4497,N_3594);
or U5885 (N_5885,N_3179,N_1456);
and U5886 (N_5886,N_125,N_619);
and U5887 (N_5887,N_1701,N_1509);
nor U5888 (N_5888,N_4044,N_4974);
nor U5889 (N_5889,N_4051,N_1423);
nor U5890 (N_5890,N_4311,N_4493);
xor U5891 (N_5891,N_1511,N_932);
xor U5892 (N_5892,N_4634,N_293);
nor U5893 (N_5893,N_3259,N_626);
nand U5894 (N_5894,N_775,N_4613);
nand U5895 (N_5895,N_986,N_2773);
xnor U5896 (N_5896,N_865,N_1470);
nand U5897 (N_5897,N_3029,N_4416);
nand U5898 (N_5898,N_3285,N_642);
nor U5899 (N_5899,N_2997,N_4063);
or U5900 (N_5900,N_1319,N_368);
nor U5901 (N_5901,N_697,N_4802);
or U5902 (N_5902,N_2459,N_4327);
or U5903 (N_5903,N_3353,N_758);
and U5904 (N_5904,N_479,N_4452);
and U5905 (N_5905,N_394,N_1662);
nor U5906 (N_5906,N_1618,N_3747);
nor U5907 (N_5907,N_2683,N_4046);
nand U5908 (N_5908,N_2807,N_3298);
and U5909 (N_5909,N_3782,N_1632);
nand U5910 (N_5910,N_4898,N_3161);
or U5911 (N_5911,N_322,N_3265);
xor U5912 (N_5912,N_4471,N_3396);
nand U5913 (N_5913,N_2171,N_4696);
and U5914 (N_5914,N_1838,N_3790);
nor U5915 (N_5915,N_1493,N_2309);
xnor U5916 (N_5916,N_4990,N_2779);
nor U5917 (N_5917,N_2058,N_434);
and U5918 (N_5918,N_540,N_2479);
and U5919 (N_5919,N_371,N_722);
and U5920 (N_5920,N_4592,N_1895);
nand U5921 (N_5921,N_3985,N_3307);
nand U5922 (N_5922,N_577,N_3328);
nor U5923 (N_5923,N_26,N_2460);
and U5924 (N_5924,N_3878,N_3666);
or U5925 (N_5925,N_2725,N_2952);
xnor U5926 (N_5926,N_321,N_6);
and U5927 (N_5927,N_1773,N_119);
or U5928 (N_5928,N_871,N_4727);
nor U5929 (N_5929,N_4025,N_2443);
or U5930 (N_5930,N_1644,N_2538);
or U5931 (N_5931,N_20,N_437);
and U5932 (N_5932,N_3037,N_2004);
or U5933 (N_5933,N_4236,N_634);
and U5934 (N_5934,N_3447,N_2657);
or U5935 (N_5935,N_2833,N_1717);
and U5936 (N_5936,N_1769,N_2410);
or U5937 (N_5937,N_494,N_4836);
and U5938 (N_5938,N_2078,N_856);
nand U5939 (N_5939,N_1401,N_407);
or U5940 (N_5940,N_2576,N_925);
nor U5941 (N_5941,N_1834,N_3250);
and U5942 (N_5942,N_1943,N_1529);
xnor U5943 (N_5943,N_2516,N_3995);
nand U5944 (N_5944,N_3717,N_3669);
nor U5945 (N_5945,N_545,N_2775);
xor U5946 (N_5946,N_2063,N_3852);
and U5947 (N_5947,N_3436,N_4265);
nand U5948 (N_5948,N_1398,N_651);
nor U5949 (N_5949,N_833,N_3119);
nor U5950 (N_5950,N_4724,N_2230);
and U5951 (N_5951,N_3068,N_983);
or U5952 (N_5952,N_3315,N_957);
or U5953 (N_5953,N_1433,N_1193);
and U5954 (N_5954,N_686,N_2875);
or U5955 (N_5955,N_361,N_2441);
nor U5956 (N_5956,N_3926,N_1947);
and U5957 (N_5957,N_27,N_3411);
nand U5958 (N_5958,N_3509,N_1553);
xor U5959 (N_5959,N_4796,N_4062);
and U5960 (N_5960,N_3642,N_1474);
or U5961 (N_5961,N_3868,N_1089);
nor U5962 (N_5962,N_4193,N_3430);
nor U5963 (N_5963,N_946,N_3101);
nor U5964 (N_5964,N_2070,N_672);
nor U5965 (N_5965,N_1577,N_3738);
xnor U5966 (N_5966,N_1990,N_1080);
and U5967 (N_5967,N_139,N_2888);
nor U5968 (N_5968,N_2671,N_1527);
or U5969 (N_5969,N_908,N_4374);
or U5970 (N_5970,N_623,N_4487);
nand U5971 (N_5971,N_2154,N_3017);
or U5972 (N_5972,N_2939,N_4017);
and U5973 (N_5973,N_3797,N_2882);
xor U5974 (N_5974,N_1337,N_653);
nor U5975 (N_5975,N_1057,N_971);
and U5976 (N_5976,N_3700,N_3286);
and U5977 (N_5977,N_2164,N_4441);
xor U5978 (N_5978,N_767,N_4729);
xor U5979 (N_5979,N_2469,N_2523);
nor U5980 (N_5980,N_2357,N_1113);
nand U5981 (N_5981,N_1373,N_4887);
and U5982 (N_5982,N_4458,N_980);
xnor U5983 (N_5983,N_71,N_981);
and U5984 (N_5984,N_3138,N_3786);
nor U5985 (N_5985,N_1586,N_2961);
nor U5986 (N_5986,N_3320,N_1182);
nand U5987 (N_5987,N_109,N_601);
and U5988 (N_5988,N_3049,N_2086);
or U5989 (N_5989,N_765,N_3856);
nor U5990 (N_5990,N_4291,N_4014);
and U5991 (N_5991,N_2601,N_2670);
and U5992 (N_5992,N_907,N_3675);
nand U5993 (N_5993,N_3740,N_179);
xor U5994 (N_5994,N_4963,N_4583);
nand U5995 (N_5995,N_274,N_993);
nor U5996 (N_5996,N_131,N_4333);
and U5997 (N_5997,N_1938,N_1183);
nand U5998 (N_5998,N_470,N_3793);
or U5999 (N_5999,N_1052,N_1200);
xnor U6000 (N_6000,N_2,N_2638);
nor U6001 (N_6001,N_2247,N_2315);
nor U6002 (N_6002,N_206,N_2319);
xnor U6003 (N_6003,N_1739,N_1948);
and U6004 (N_6004,N_381,N_4426);
or U6005 (N_6005,N_195,N_2579);
or U6006 (N_6006,N_832,N_242);
xnor U6007 (N_6007,N_4692,N_4932);
or U6008 (N_6008,N_3446,N_4743);
or U6009 (N_6009,N_4102,N_3760);
or U6010 (N_6010,N_1534,N_1087);
xor U6011 (N_6011,N_4347,N_2049);
nor U6012 (N_6012,N_2628,N_4506);
nand U6013 (N_6013,N_2652,N_956);
and U6014 (N_6014,N_2748,N_2481);
and U6015 (N_6015,N_2377,N_4864);
and U6016 (N_6016,N_4532,N_1102);
xor U6017 (N_6017,N_3954,N_4770);
and U6018 (N_6018,N_2587,N_4370);
and U6019 (N_6019,N_3778,N_2718);
nor U6020 (N_6020,N_94,N_128);
or U6021 (N_6021,N_1698,N_1260);
or U6022 (N_6022,N_961,N_4107);
or U6023 (N_6023,N_2364,N_4354);
and U6024 (N_6024,N_2194,N_3540);
nand U6025 (N_6025,N_3432,N_3869);
nand U6026 (N_6026,N_4412,N_3813);
or U6027 (N_6027,N_4340,N_2401);
nand U6028 (N_6028,N_3876,N_1302);
or U6029 (N_6029,N_4301,N_383);
or U6030 (N_6030,N_2824,N_2228);
or U6031 (N_6031,N_921,N_3312);
nor U6032 (N_6032,N_3998,N_3349);
nand U6033 (N_6033,N_1569,N_4119);
or U6034 (N_6034,N_375,N_674);
and U6035 (N_6035,N_1404,N_843);
or U6036 (N_6036,N_211,N_2550);
or U6037 (N_6037,N_782,N_2542);
nand U6038 (N_6038,N_2417,N_542);
nor U6039 (N_6039,N_4979,N_3977);
and U6040 (N_6040,N_2129,N_4580);
xor U6041 (N_6041,N_1864,N_3768);
or U6042 (N_6042,N_1181,N_1665);
nor U6043 (N_6043,N_3148,N_3836);
and U6044 (N_6044,N_3806,N_3165);
xnor U6045 (N_6045,N_3582,N_1380);
nand U6046 (N_6046,N_2030,N_4058);
or U6047 (N_6047,N_1951,N_2568);
or U6048 (N_6048,N_4283,N_2703);
nand U6049 (N_6049,N_3947,N_4092);
nand U6050 (N_6050,N_1387,N_3822);
nand U6051 (N_6051,N_3774,N_3829);
nor U6052 (N_6052,N_4681,N_1307);
nand U6053 (N_6053,N_3024,N_4703);
nand U6054 (N_6054,N_2661,N_905);
nor U6055 (N_6055,N_1689,N_1196);
and U6056 (N_6056,N_2268,N_3480);
and U6057 (N_6057,N_4060,N_4626);
nor U6058 (N_6058,N_4171,N_3407);
and U6059 (N_6059,N_2956,N_2034);
nand U6060 (N_6060,N_701,N_2046);
nor U6061 (N_6061,N_1696,N_3690);
nand U6062 (N_6062,N_4579,N_1972);
nand U6063 (N_6063,N_3950,N_41);
nand U6064 (N_6064,N_331,N_4081);
nor U6065 (N_6065,N_2506,N_3611);
nor U6066 (N_6066,N_2474,N_2658);
nand U6067 (N_6067,N_1591,N_3742);
and U6068 (N_6068,N_637,N_130);
nand U6069 (N_6069,N_2620,N_4309);
nor U6070 (N_6070,N_25,N_4117);
or U6071 (N_6071,N_4355,N_4602);
and U6072 (N_6072,N_449,N_4607);
nand U6073 (N_6073,N_718,N_3667);
nor U6074 (N_6074,N_57,N_1159);
nand U6075 (N_6075,N_1523,N_1257);
nand U6076 (N_6076,N_1899,N_3050);
nor U6077 (N_6077,N_3424,N_4504);
or U6078 (N_6078,N_3440,N_3915);
nor U6079 (N_6079,N_3040,N_4339);
nor U6080 (N_6080,N_4035,N_3676);
or U6081 (N_6081,N_3386,N_172);
nand U6082 (N_6082,N_2388,N_2709);
or U6083 (N_6083,N_4167,N_3862);
nand U6084 (N_6084,N_1850,N_2141);
xor U6085 (N_6085,N_703,N_1891);
nor U6086 (N_6086,N_304,N_448);
nand U6087 (N_6087,N_2563,N_4282);
nand U6088 (N_6088,N_2286,N_2662);
xnor U6089 (N_6089,N_4155,N_3688);
nand U6090 (N_6090,N_4209,N_1438);
nor U6091 (N_6091,N_3753,N_3231);
and U6092 (N_6092,N_3108,N_3946);
and U6093 (N_6093,N_83,N_4734);
nand U6094 (N_6094,N_9,N_63);
or U6095 (N_6095,N_3116,N_1137);
nand U6096 (N_6096,N_2864,N_4555);
and U6097 (N_6097,N_1629,N_3671);
or U6098 (N_6098,N_3373,N_3371);
nor U6099 (N_6099,N_3834,N_1005);
nand U6100 (N_6100,N_4590,N_3752);
xnor U6101 (N_6101,N_231,N_3886);
or U6102 (N_6102,N_2647,N_2701);
nand U6103 (N_6103,N_1449,N_745);
and U6104 (N_6104,N_416,N_3920);
and U6105 (N_6105,N_3734,N_2645);
nand U6106 (N_6106,N_1780,N_824);
xnor U6107 (N_6107,N_2653,N_854);
nor U6108 (N_6108,N_2857,N_3645);
xor U6109 (N_6109,N_4230,N_617);
nand U6110 (N_6110,N_3895,N_2050);
nand U6111 (N_6111,N_1166,N_3098);
and U6112 (N_6112,N_1078,N_405);
and U6113 (N_6113,N_3156,N_341);
nor U6114 (N_6114,N_3412,N_96);
xor U6115 (N_6115,N_3413,N_3258);
xnor U6116 (N_6116,N_2817,N_859);
or U6117 (N_6117,N_4314,N_976);
and U6118 (N_6118,N_3817,N_425);
nor U6119 (N_6119,N_689,N_2539);
nor U6120 (N_6120,N_2051,N_802);
nand U6121 (N_6121,N_3051,N_1303);
nand U6122 (N_6122,N_4782,N_3157);
and U6123 (N_6123,N_696,N_699);
nand U6124 (N_6124,N_4656,N_2573);
and U6125 (N_6125,N_2558,N_4324);
nor U6126 (N_6126,N_4296,N_3610);
and U6127 (N_6127,N_3247,N_1285);
or U6128 (N_6128,N_1996,N_3194);
and U6129 (N_6129,N_1515,N_1852);
or U6130 (N_6130,N_1926,N_3544);
or U6131 (N_6131,N_1261,N_4138);
and U6132 (N_6132,N_3109,N_2075);
nor U6133 (N_6133,N_2731,N_389);
nor U6134 (N_6134,N_1503,N_2135);
nor U6135 (N_6135,N_373,N_4589);
xnor U6136 (N_6136,N_4646,N_2712);
xnor U6137 (N_6137,N_886,N_2381);
nor U6138 (N_6138,N_4381,N_910);
xor U6139 (N_6139,N_715,N_3171);
xnor U6140 (N_6140,N_183,N_1860);
nor U6141 (N_6141,N_467,N_15);
nor U6142 (N_6142,N_1984,N_4166);
nand U6143 (N_6143,N_4529,N_4730);
or U6144 (N_6144,N_4299,N_4350);
or U6145 (N_6145,N_4162,N_2560);
xnor U6146 (N_6146,N_3048,N_4116);
or U6147 (N_6147,N_117,N_3072);
and U6148 (N_6148,N_1716,N_1742);
xnor U6149 (N_6149,N_3135,N_1163);
nand U6150 (N_6150,N_2425,N_554);
or U6151 (N_6151,N_3940,N_457);
nand U6152 (N_6152,N_1674,N_1115);
or U6153 (N_6153,N_3945,N_4515);
nand U6154 (N_6154,N_1590,N_1536);
nor U6155 (N_6155,N_1322,N_2333);
and U6156 (N_6156,N_2983,N_2609);
and U6157 (N_6157,N_1754,N_2761);
and U6158 (N_6158,N_1032,N_4644);
and U6159 (N_6159,N_3418,N_3841);
or U6160 (N_6160,N_743,N_1753);
xnor U6161 (N_6161,N_2107,N_2789);
nor U6162 (N_6162,N_519,N_2894);
and U6163 (N_6163,N_395,N_927);
and U6164 (N_6164,N_73,N_2343);
or U6165 (N_6165,N_596,N_4600);
nand U6166 (N_6166,N_4906,N_1968);
and U6167 (N_6167,N_12,N_1116);
or U6168 (N_6168,N_1010,N_3054);
or U6169 (N_6169,N_1374,N_3921);
and U6170 (N_6170,N_3937,N_1111);
and U6171 (N_6171,N_3574,N_2336);
nor U6172 (N_6172,N_3267,N_4793);
and U6173 (N_6173,N_3673,N_188);
or U6174 (N_6174,N_2354,N_3483);
or U6175 (N_6175,N_4742,N_2868);
xor U6176 (N_6176,N_4137,N_3296);
xor U6177 (N_6177,N_4522,N_1900);
or U6178 (N_6178,N_3366,N_3005);
or U6179 (N_6179,N_4187,N_1425);
nand U6180 (N_6180,N_2784,N_3280);
nor U6181 (N_6181,N_3271,N_4857);
nand U6182 (N_6182,N_3473,N_2025);
nor U6183 (N_6183,N_848,N_163);
nor U6184 (N_6184,N_3031,N_4313);
nor U6185 (N_6185,N_1784,N_3843);
xnor U6186 (N_6186,N_2519,N_1140);
nor U6187 (N_6187,N_4443,N_4028);
or U6188 (N_6188,N_3221,N_2535);
xnor U6189 (N_6189,N_989,N_4970);
and U6190 (N_6190,N_1413,N_4784);
nor U6191 (N_6191,N_3615,N_2747);
xnor U6192 (N_6192,N_4790,N_1355);
and U6193 (N_6193,N_4218,N_4954);
and U6194 (N_6194,N_4010,N_2454);
or U6195 (N_6195,N_1933,N_4910);
nand U6196 (N_6196,N_1266,N_4341);
and U6197 (N_6197,N_355,N_1141);
nor U6198 (N_6198,N_3364,N_3754);
xor U6199 (N_6199,N_2355,N_1542);
nor U6200 (N_6200,N_1915,N_2136);
and U6201 (N_6201,N_319,N_1370);
nor U6202 (N_6202,N_4637,N_574);
nor U6203 (N_6203,N_534,N_964);
or U6204 (N_6204,N_3503,N_289);
nand U6205 (N_6205,N_460,N_798);
xnor U6206 (N_6206,N_2306,N_4210);
or U6207 (N_6207,N_3827,N_2281);
nand U6208 (N_6208,N_3859,N_2043);
nand U6209 (N_6209,N_1782,N_4277);
xor U6210 (N_6210,N_203,N_4889);
or U6211 (N_6211,N_1655,N_2010);
nand U6212 (N_6212,N_3978,N_362);
or U6213 (N_6213,N_996,N_1095);
nand U6214 (N_6214,N_2452,N_3763);
nor U6215 (N_6215,N_4513,N_1484);
nor U6216 (N_6216,N_2940,N_2912);
nand U6217 (N_6217,N_1272,N_1574);
nand U6218 (N_6218,N_4904,N_787);
and U6219 (N_6219,N_3619,N_1727);
or U6220 (N_6220,N_3313,N_3518);
nor U6221 (N_6221,N_3030,N_2525);
or U6222 (N_6222,N_1783,N_3779);
and U6223 (N_6223,N_1009,N_3577);
nor U6224 (N_6224,N_2255,N_711);
nor U6225 (N_6225,N_662,N_1290);
and U6226 (N_6226,N_1424,N_65);
nand U6227 (N_6227,N_4552,N_973);
and U6228 (N_6228,N_3317,N_169);
or U6229 (N_6229,N_2596,N_477);
and U6230 (N_6230,N_694,N_4140);
and U6231 (N_6231,N_4803,N_2123);
xnor U6232 (N_6232,N_2659,N_4099);
or U6233 (N_6233,N_4584,N_4485);
nor U6234 (N_6234,N_4837,N_3962);
nand U6235 (N_6235,N_4971,N_411);
nand U6236 (N_6236,N_4940,N_1353);
and U6237 (N_6237,N_1473,N_1343);
xor U6238 (N_6238,N_1227,N_2375);
or U6239 (N_6239,N_2321,N_4059);
nor U6240 (N_6240,N_1409,N_3839);
nand U6241 (N_6241,N_4804,N_4332);
and U6242 (N_6242,N_4462,N_4305);
nand U6243 (N_6243,N_3304,N_173);
and U6244 (N_6244,N_4004,N_384);
nand U6245 (N_6245,N_3603,N_1384);
xor U6246 (N_6246,N_4226,N_3429);
nor U6247 (N_6247,N_1489,N_397);
or U6248 (N_6248,N_207,N_4706);
or U6249 (N_6249,N_3491,N_334);
and U6250 (N_6250,N_4668,N_4246);
and U6251 (N_6251,N_3818,N_2887);
or U6252 (N_6252,N_1385,N_4295);
xor U6253 (N_6253,N_3173,N_1559);
and U6254 (N_6254,N_1964,N_2103);
and U6255 (N_6255,N_1072,N_1877);
xor U6256 (N_6256,N_1645,N_3586);
or U6257 (N_6257,N_4969,N_3644);
nor U6258 (N_6258,N_3226,N_3125);
xor U6259 (N_6259,N_4446,N_3901);
and U6260 (N_6260,N_737,N_3898);
and U6261 (N_6261,N_1911,N_1763);
nand U6262 (N_6262,N_2593,N_2746);
nor U6263 (N_6263,N_3458,N_934);
xnor U6264 (N_6264,N_1247,N_710);
nor U6265 (N_6265,N_3064,N_4245);
xor U6266 (N_6266,N_3337,N_454);
xor U6267 (N_6267,N_3485,N_3236);
xnor U6268 (N_6268,N_4801,N_2334);
nand U6269 (N_6269,N_196,N_2056);
and U6270 (N_6270,N_4173,N_913);
or U6271 (N_6271,N_997,N_2623);
nor U6272 (N_6272,N_2477,N_728);
xnor U6273 (N_6273,N_3670,N_1691);
nand U6274 (N_6274,N_3435,N_2282);
nor U6275 (N_6275,N_1555,N_3158);
nor U6276 (N_6276,N_675,N_3389);
or U6277 (N_6277,N_4371,N_677);
nand U6278 (N_6278,N_873,N_3427);
or U6279 (N_6279,N_1037,N_307);
and U6280 (N_6280,N_4410,N_2475);
nand U6281 (N_6281,N_3426,N_4789);
nand U6282 (N_6282,N_62,N_880);
and U6283 (N_6283,N_972,N_4908);
nor U6284 (N_6284,N_1268,N_22);
or U6285 (N_6285,N_3548,N_1960);
nand U6286 (N_6286,N_3186,N_2687);
or U6287 (N_6287,N_4078,N_4242);
nor U6288 (N_6288,N_3847,N_3913);
xnor U6289 (N_6289,N_10,N_1184);
or U6290 (N_6290,N_3333,N_91);
nor U6291 (N_6291,N_4160,N_2822);
nand U6292 (N_6292,N_1925,N_761);
nor U6293 (N_6293,N_4098,N_2209);
nand U6294 (N_6294,N_4867,N_3845);
nand U6295 (N_6295,N_423,N_3877);
nand U6296 (N_6296,N_2053,N_2831);
nor U6297 (N_6297,N_3653,N_2879);
nand U6298 (N_6298,N_1913,N_3335);
nor U6299 (N_6299,N_2297,N_3065);
or U6300 (N_6300,N_4150,N_469);
and U6301 (N_6301,N_251,N_4996);
and U6302 (N_6302,N_2005,N_143);
or U6303 (N_6303,N_165,N_2222);
nor U6304 (N_6304,N_3731,N_85);
nor U6305 (N_6305,N_2184,N_1437);
and U6306 (N_6306,N_4748,N_4956);
nor U6307 (N_6307,N_111,N_2503);
nor U6308 (N_6308,N_3181,N_691);
and U6309 (N_6309,N_618,N_2632);
or U6310 (N_6310,N_3715,N_4118);
and U6311 (N_6311,N_2914,N_40);
nor U6312 (N_6312,N_1693,N_1065);
nor U6313 (N_6313,N_4849,N_3130);
nor U6314 (N_6314,N_4704,N_3062);
nand U6315 (N_6315,N_4941,N_2790);
or U6316 (N_6316,N_1957,N_1075);
xor U6317 (N_6317,N_4030,N_1827);
or U6318 (N_6318,N_1061,N_917);
nand U6319 (N_6319,N_1133,N_2936);
nand U6320 (N_6320,N_2398,N_1469);
or U6321 (N_6321,N_1497,N_2931);
xnor U6322 (N_6322,N_4213,N_4563);
nor U6323 (N_6323,N_3196,N_2322);
nor U6324 (N_6324,N_4172,N_244);
nand U6325 (N_6325,N_3626,N_4043);
xnor U6326 (N_6326,N_1390,N_1241);
nor U6327 (N_6327,N_1238,N_1084);
or U6328 (N_6328,N_4780,N_3475);
or U6329 (N_6329,N_3914,N_2337);
nand U6330 (N_6330,N_4079,N_3002);
nand U6331 (N_6331,N_115,N_1912);
or U6332 (N_6332,N_388,N_4854);
nand U6333 (N_6333,N_1666,N_3522);
nor U6334 (N_6334,N_4835,N_404);
nor U6335 (N_6335,N_1106,N_1906);
and U6336 (N_6336,N_580,N_1070);
and U6337 (N_6337,N_1048,N_3963);
or U6338 (N_6338,N_3781,N_486);
and U6339 (N_6339,N_575,N_2646);
or U6340 (N_6340,N_3351,N_3555);
nand U6341 (N_6341,N_1898,N_1277);
nand U6342 (N_6342,N_228,N_4944);
and U6343 (N_6343,N_4294,N_4125);
nor U6344 (N_6344,N_1690,N_4310);
or U6345 (N_6345,N_1776,N_4484);
nor U6346 (N_6346,N_3372,N_193);
and U6347 (N_6347,N_3602,N_2984);
nor U6348 (N_6348,N_116,N_2869);
or U6349 (N_6349,N_2111,N_1013);
or U6350 (N_6350,N_2694,N_3557);
and U6351 (N_6351,N_2464,N_2003);
or U6352 (N_6352,N_607,N_2667);
and U6353 (N_6353,N_3571,N_3057);
and U6354 (N_6354,N_4759,N_1610);
nor U6355 (N_6355,N_2421,N_3151);
and U6356 (N_6356,N_2501,N_2455);
nand U6357 (N_6357,N_2504,N_3857);
nor U6358 (N_6358,N_1791,N_4321);
nor U6359 (N_6359,N_2159,N_1118);
and U6360 (N_6360,N_4387,N_3887);
nand U6361 (N_6361,N_1139,N_4624);
nor U6362 (N_6362,N_4135,N_768);
or U6363 (N_6363,N_3249,N_746);
nand U6364 (N_6364,N_4968,N_1998);
xor U6365 (N_6365,N_332,N_308);
nor U6366 (N_6366,N_2960,N_4480);
and U6367 (N_6367,N_2531,N_2483);
nand U6368 (N_6368,N_3336,N_2871);
xor U6369 (N_6369,N_3705,N_4325);
nand U6370 (N_6370,N_2232,N_509);
nand U6371 (N_6371,N_4686,N_2394);
nand U6372 (N_6372,N_2068,N_4403);
or U6373 (N_6373,N_4972,N_270);
or U6374 (N_6374,N_161,N_2555);
nor U6375 (N_6375,N_3302,N_2092);
or U6376 (N_6376,N_4307,N_1434);
nor U6377 (N_6377,N_3257,N_4009);
and U6378 (N_6378,N_968,N_3075);
and U6379 (N_6379,N_2059,N_3263);
nand U6380 (N_6380,N_4926,N_2840);
or U6381 (N_6381,N_2431,N_3355);
or U6382 (N_6382,N_1393,N_1499);
nor U6383 (N_6383,N_3453,N_2518);
nor U6384 (N_6384,N_4366,N_1056);
and U6385 (N_6385,N_3238,N_4405);
and U6386 (N_6386,N_3342,N_556);
or U6387 (N_6387,N_1412,N_4618);
nand U6388 (N_6388,N_1781,N_2400);
nor U6389 (N_6389,N_936,N_1232);
and U6390 (N_6390,N_4541,N_1366);
nand U6391 (N_6391,N_3837,N_3534);
nor U6392 (N_6392,N_3596,N_1215);
and U6393 (N_6393,N_593,N_1909);
and U6394 (N_6394,N_1164,N_2631);
and U6395 (N_6395,N_2808,N_4344);
nor U6396 (N_6396,N_2892,N_527);
or U6397 (N_6397,N_4271,N_4884);
or U6398 (N_6398,N_224,N_419);
nand U6399 (N_6399,N_1713,N_4571);
and U6400 (N_6400,N_2289,N_2995);
and U6401 (N_6401,N_4454,N_3319);
nor U6402 (N_6402,N_2689,N_1477);
nor U6403 (N_6403,N_1556,N_3367);
nor U6404 (N_6404,N_2055,N_421);
and U6405 (N_6405,N_4746,N_488);
and U6406 (N_6406,N_3383,N_1097);
and U6407 (N_6407,N_2018,N_4142);
nor U6408 (N_6408,N_2299,N_3270);
nand U6409 (N_6409,N_1857,N_4931);
or U6410 (N_6410,N_2675,N_3578);
nand U6411 (N_6411,N_4034,N_1265);
nand U6412 (N_6412,N_2426,N_3785);
or U6413 (N_6413,N_1076,N_4400);
nor U6414 (N_6414,N_2150,N_4342);
nand U6415 (N_6415,N_4712,N_2074);
nand U6416 (N_6416,N_2597,N_2244);
or U6417 (N_6417,N_1826,N_44);
or U6418 (N_6418,N_2250,N_4876);
and U6419 (N_6419,N_4148,N_3036);
and U6420 (N_6420,N_3639,N_2985);
nor U6421 (N_6421,N_81,N_4840);
xnor U6422 (N_6422,N_3732,N_312);
or U6423 (N_6423,N_522,N_1288);
or U6424 (N_6424,N_3777,N_2935);
and U6425 (N_6425,N_2553,N_2621);
and U6426 (N_6426,N_941,N_2205);
nand U6427 (N_6427,N_3894,N_635);
nand U6428 (N_6428,N_4617,N_4919);
nor U6429 (N_6429,N_2828,N_3943);
or U6430 (N_6430,N_2254,N_3712);
xnor U6431 (N_6431,N_4885,N_1162);
nor U6432 (N_6432,N_3405,N_3607);
or U6433 (N_6433,N_3860,N_3000);
nand U6434 (N_6434,N_2970,N_1755);
nor U6435 (N_6435,N_4622,N_1280);
xor U6436 (N_6436,N_4038,N_4024);
or U6437 (N_6437,N_3490,N_3960);
nor U6438 (N_6438,N_3944,N_2095);
and U6439 (N_6439,N_235,N_347);
or U6440 (N_6440,N_3408,N_3622);
nor U6441 (N_6441,N_4546,N_3150);
nand U6442 (N_6442,N_2214,N_2433);
or U6443 (N_6443,N_1526,N_103);
nor U6444 (N_6444,N_4629,N_112);
and U6445 (N_6445,N_445,N_82);
nand U6446 (N_6446,N_885,N_1104);
nor U6447 (N_6447,N_1825,N_4832);
nand U6448 (N_6448,N_2249,N_1516);
and U6449 (N_6449,N_2534,N_1408);
or U6450 (N_6450,N_4040,N_1884);
xor U6451 (N_6451,N_4992,N_3826);
or U6452 (N_6452,N_2045,N_3281);
and U6453 (N_6453,N_378,N_264);
and U6454 (N_6454,N_2017,N_1371);
nor U6455 (N_6455,N_4769,N_431);
nand U6456 (N_6456,N_3704,N_2919);
nand U6457 (N_6457,N_4964,N_924);
or U6458 (N_6458,N_2818,N_667);
nand U6459 (N_6459,N_2907,N_3637);
xnor U6460 (N_6460,N_536,N_1221);
nand U6461 (N_6461,N_4630,N_867);
nor U6462 (N_6462,N_444,N_2644);
nor U6463 (N_6463,N_555,N_4445);
nor U6464 (N_6464,N_2016,N_1731);
nand U6465 (N_6465,N_1934,N_3971);
nand U6466 (N_6466,N_4586,N_2937);
and U6467 (N_6467,N_1151,N_4995);
nor U6468 (N_6468,N_2769,N_4511);
or U6469 (N_6469,N_673,N_1300);
or U6470 (N_6470,N_462,N_1735);
nor U6471 (N_6471,N_4855,N_4077);
and U6472 (N_6472,N_3864,N_2781);
and U6473 (N_6473,N_337,N_3663);
nor U6474 (N_6474,N_4414,N_4191);
or U6475 (N_6475,N_3398,N_4161);
nand U6476 (N_6476,N_1492,N_4337);
and U6477 (N_6477,N_4133,N_4105);
xor U6478 (N_6478,N_2917,N_901);
and U6479 (N_6479,N_3385,N_1896);
or U6480 (N_6480,N_3085,N_2890);
nand U6481 (N_6481,N_1809,N_3211);
and U6482 (N_6482,N_2484,N_3295);
nor U6483 (N_6483,N_1046,N_3802);
and U6484 (N_6484,N_974,N_4761);
nand U6485 (N_6485,N_4451,N_1336);
or U6486 (N_6486,N_1582,N_2201);
or U6487 (N_6487,N_1770,N_436);
and U6488 (N_6488,N_2052,N_666);
and U6489 (N_6489,N_2872,N_3146);
nand U6490 (N_6490,N_2226,N_3495);
or U6491 (N_6491,N_2386,N_3941);
xor U6492 (N_6492,N_3451,N_846);
nor U6493 (N_6493,N_3235,N_345);
or U6494 (N_6494,N_1243,N_249);
or U6495 (N_6495,N_1186,N_2741);
nand U6496 (N_6496,N_4254,N_3636);
xor U6497 (N_6497,N_189,N_2528);
nor U6498 (N_6498,N_4527,N_2453);
nor U6499 (N_6499,N_4521,N_4641);
and U6500 (N_6500,N_995,N_2440);
nor U6501 (N_6501,N_797,N_965);
nand U6502 (N_6502,N_1916,N_167);
nor U6503 (N_6503,N_3880,N_720);
nor U6504 (N_6504,N_1738,N_2248);
and U6505 (N_6505,N_221,N_3858);
nor U6506 (N_6506,N_2759,N_4476);
and U6507 (N_6507,N_311,N_2186);
nand U6508 (N_6508,N_4392,N_1362);
or U6509 (N_6509,N_780,N_2716);
xor U6510 (N_6510,N_4900,N_2403);
and U6511 (N_6511,N_978,N_582);
or U6512 (N_6512,N_614,N_1855);
nand U6513 (N_6513,N_1928,N_2643);
or U6514 (N_6514,N_2236,N_1604);
nor U6515 (N_6515,N_949,N_14);
nand U6516 (N_6516,N_464,N_1093);
nor U6517 (N_6517,N_278,N_398);
xnor U6518 (N_6518,N_511,N_3514);
or U6519 (N_6519,N_3572,N_2471);
nor U6520 (N_6520,N_2102,N_180);
and U6521 (N_6521,N_1292,N_77);
or U6522 (N_6522,N_3083,N_4429);
nor U6523 (N_6523,N_2174,N_1734);
xor U6524 (N_6524,N_2946,N_2239);
nand U6525 (N_6525,N_4921,N_1697);
nor U6526 (N_6526,N_2077,N_2520);
and U6527 (N_6527,N_647,N_1346);
nor U6528 (N_6528,N_4710,N_463);
or U6529 (N_6529,N_1808,N_4728);
or U6530 (N_6530,N_4591,N_3006);
xor U6531 (N_6531,N_4866,N_4953);
nand U6532 (N_6532,N_2546,N_3182);
and U6533 (N_6533,N_499,N_2588);
nor U6534 (N_6534,N_3464,N_1740);
and U6535 (N_6535,N_1224,N_3923);
and U6536 (N_6536,N_4258,N_1538);
and U6537 (N_6537,N_2788,N_525);
and U6538 (N_6538,N_2029,N_4883);
or U6539 (N_6539,N_636,N_2478);
nor U6540 (N_6540,N_181,N_1249);
nand U6541 (N_6541,N_3884,N_1167);
and U6542 (N_6542,N_441,N_4072);
or U6543 (N_6543,N_1853,N_2836);
nand U6544 (N_6544,N_4463,N_4762);
xnor U6545 (N_6545,N_4978,N_2825);
nor U6546 (N_6546,N_4195,N_1490);
nor U6547 (N_6547,N_2276,N_3867);
or U6548 (N_6548,N_1599,N_3583);
nor U6549 (N_6549,N_3710,N_4049);
nor U6550 (N_6550,N_1954,N_3668);
nor U6551 (N_6551,N_4466,N_4262);
nand U6552 (N_6552,N_50,N_88);
or U6553 (N_6553,N_2356,N_305);
and U6554 (N_6554,N_2237,N_3955);
nand U6555 (N_6555,N_505,N_3104);
nor U6556 (N_6556,N_3632,N_2739);
nand U6557 (N_6557,N_3750,N_2615);
nor U6558 (N_6558,N_4349,N_858);
and U6559 (N_6559,N_1801,N_969);
nor U6560 (N_6560,N_3918,N_3362);
or U6561 (N_6561,N_3588,N_1725);
nor U6562 (N_6562,N_2090,N_1073);
nand U6563 (N_6563,N_1487,N_3456);
nor U6564 (N_6564,N_3502,N_1014);
or U6565 (N_6565,N_2392,N_1230);
or U6566 (N_6566,N_3466,N_1602);
xnor U6567 (N_6567,N_4159,N_4615);
nand U6568 (N_6568,N_3217,N_890);
xnor U6569 (N_6569,N_2774,N_1472);
or U6570 (N_6570,N_1418,N_1218);
nor U6571 (N_6571,N_579,N_835);
nand U6572 (N_6572,N_4240,N_1950);
and U6573 (N_6573,N_3166,N_4750);
or U6574 (N_6574,N_4013,N_3149);
nor U6575 (N_6575,N_4825,N_3707);
nand U6576 (N_6576,N_4509,N_4920);
nor U6577 (N_6577,N_3716,N_3618);
nor U6578 (N_6578,N_54,N_2796);
xnor U6579 (N_6579,N_2259,N_4490);
and U6580 (N_6580,N_310,N_1813);
and U6581 (N_6581,N_327,N_4205);
nor U6582 (N_6582,N_2957,N_3016);
and U6583 (N_6583,N_3552,N_266);
nor U6584 (N_6584,N_1510,N_4994);
or U6585 (N_6585,N_1854,N_1354);
and U6586 (N_6586,N_549,N_4290);
nand U6587 (N_6587,N_471,N_4512);
and U6588 (N_6588,N_3528,N_3322);
nor U6589 (N_6589,N_1902,N_837);
xnor U6590 (N_6590,N_4839,N_4238);
and U6591 (N_6591,N_538,N_2795);
and U6592 (N_6592,N_3169,N_4967);
nand U6593 (N_6593,N_2541,N_1575);
nand U6594 (N_6594,N_2006,N_237);
and U6595 (N_6595,N_2860,N_147);
and U6596 (N_6596,N_4564,N_1391);
nand U6597 (N_6597,N_1101,N_4136);
or U6598 (N_6598,N_2369,N_135);
xor U6599 (N_6599,N_1088,N_939);
nor U6600 (N_6600,N_3174,N_1006);
nand U6601 (N_6601,N_640,N_1306);
or U6602 (N_6602,N_3787,N_4942);
xnor U6603 (N_6603,N_1201,N_1150);
nand U6604 (N_6604,N_4518,N_1584);
or U6605 (N_6605,N_2977,N_4415);
nand U6606 (N_6606,N_2000,N_417);
or U6607 (N_6607,N_2120,N_875);
nor U6608 (N_6608,N_2742,N_1507);
xnor U6609 (N_6609,N_2367,N_3609);
xnor U6610 (N_6610,N_2380,N_3140);
or U6611 (N_6611,N_3212,N_4877);
nor U6612 (N_6612,N_4597,N_3227);
nand U6613 (N_6613,N_1921,N_2273);
nand U6614 (N_6614,N_1640,N_4065);
nand U6615 (N_6615,N_153,N_3077);
and U6616 (N_6616,N_4757,N_3741);
nand U6617 (N_6617,N_808,N_2552);
or U6618 (N_6618,N_563,N_1839);
xnor U6619 (N_6619,N_984,N_3465);
xnor U6620 (N_6620,N_2724,N_3706);
nor U6621 (N_6621,N_1772,N_1015);
nand U6622 (N_6622,N_3564,N_2023);
or U6623 (N_6623,N_4373,N_531);
nor U6624 (N_6624,N_1956,N_3801);
nor U6625 (N_6625,N_1023,N_3470);
nor U6626 (N_6626,N_1340,N_2185);
nor U6627 (N_6627,N_2036,N_3223);
and U6628 (N_6628,N_268,N_2224);
and U6629 (N_6629,N_3988,N_2938);
or U6630 (N_6630,N_4022,N_4402);
or U6631 (N_6631,N_4899,N_2794);
nor U6632 (N_6632,N_3568,N_2265);
or U6633 (N_6633,N_3378,N_1244);
nand U6634 (N_6634,N_4980,N_739);
and U6635 (N_6635,N_857,N_1637);
or U6636 (N_6636,N_4288,N_2706);
or U6637 (N_6637,N_4871,N_2569);
or U6638 (N_6638,N_2411,N_3530);
or U6639 (N_6639,N_1321,N_220);
nor U6640 (N_6640,N_4233,N_1606);
nor U6641 (N_6641,N_3251,N_4614);
xor U6642 (N_6642,N_2211,N_2768);
nand U6643 (N_6643,N_4721,N_1810);
nor U6644 (N_6644,N_4575,N_4431);
and U6645 (N_6645,N_1108,N_4909);
and U6646 (N_6646,N_4353,N_3507);
nor U6647 (N_6647,N_363,N_4988);
nor U6648 (N_6648,N_4648,N_3679);
and U6649 (N_6649,N_3084,N_2536);
nor U6650 (N_6650,N_687,N_4822);
or U6651 (N_6651,N_1041,N_4888);
nor U6652 (N_6652,N_3792,N_610);
nor U6653 (N_6653,N_2430,N_1466);
nand U6654 (N_6654,N_4933,N_4469);
and U6655 (N_6655,N_4114,N_4131);
and U6656 (N_6656,N_2206,N_4139);
nor U6657 (N_6657,N_1394,N_1981);
nand U6658 (N_6658,N_3141,N_3762);
nor U6659 (N_6659,N_4923,N_3997);
nand U6660 (N_6660,N_1684,N_900);
nand U6661 (N_6661,N_1872,N_3870);
or U6662 (N_6662,N_4902,N_2127);
xnor U6663 (N_6663,N_811,N_2264);
xnor U6664 (N_6664,N_2304,N_2233);
nor U6665 (N_6665,N_3460,N_2673);
nand U6666 (N_6666,N_3816,N_1357);
nor U6667 (N_6667,N_2780,N_788);
nor U6668 (N_6668,N_4052,N_2191);
nor U6669 (N_6669,N_1317,N_1941);
nand U6670 (N_6670,N_4188,N_3575);
nand U6671 (N_6671,N_3948,N_4239);
nor U6672 (N_6672,N_79,N_4841);
nand U6673 (N_6673,N_3500,N_177);
and U6674 (N_6674,N_747,N_4999);
and U6675 (N_6675,N_4951,N_356);
or U6676 (N_6676,N_1094,N_4585);
and U6677 (N_6677,N_1442,N_354);
xor U6678 (N_6678,N_1871,N_1185);
nand U6679 (N_6679,N_1927,N_3323);
xor U6680 (N_6680,N_3309,N_4623);
nor U6681 (N_6681,N_3496,N_2707);
nand U6682 (N_6682,N_4165,N_751);
or U6683 (N_6683,N_34,N_2192);
nand U6684 (N_6684,N_218,N_3771);
or U6685 (N_6685,N_633,N_4229);
nand U6686 (N_6686,N_878,N_3442);
nand U6687 (N_6687,N_4753,N_2373);
and U6688 (N_6688,N_1876,N_2130);
nor U6689 (N_6689,N_3402,N_3080);
nor U6690 (N_6690,N_199,N_1245);
nor U6691 (N_6691,N_1795,N_2436);
nand U6692 (N_6692,N_3604,N_1460);
or U6693 (N_6693,N_4360,N_1837);
or U6694 (N_6694,N_3651,N_4019);
xnor U6695 (N_6695,N_643,N_1369);
nor U6696 (N_6696,N_3949,N_2026);
and U6697 (N_6697,N_1358,N_4664);
nand U6698 (N_6698,N_295,N_2147);
nor U6699 (N_6699,N_1211,N_1289);
nor U6700 (N_6700,N_1021,N_4540);
nor U6701 (N_6701,N_2517,N_2376);
nor U6702 (N_6702,N_4976,N_3842);
or U6703 (N_6703,N_2726,N_1616);
nor U6704 (N_6704,N_3045,N_533);
and U6705 (N_6705,N_4763,N_2350);
or U6706 (N_6706,N_3420,N_2256);
nor U6707 (N_6707,N_2529,N_4219);
or U6708 (N_6708,N_1403,N_4164);
and U6709 (N_6709,N_3287,N_4775);
or U6710 (N_6710,N_826,N_1160);
or U6711 (N_6711,N_2925,N_3751);
nand U6712 (N_6712,N_4127,N_1429);
and U6713 (N_6713,N_132,N_2903);
or U6714 (N_6714,N_4498,N_3885);
xor U6715 (N_6715,N_840,N_3983);
nor U6716 (N_6716,N_3593,N_2346);
or U6717 (N_6717,N_1595,N_338);
nand U6718 (N_6718,N_4372,N_1212);
or U6719 (N_6719,N_1044,N_4259);
and U6720 (N_6720,N_1995,N_4989);
nor U6721 (N_6721,N_2301,N_2329);
nand U6722 (N_6722,N_1888,N_4303);
or U6723 (N_6723,N_1480,N_3529);
and U6724 (N_6724,N_175,N_4651);
and U6725 (N_6725,N_1476,N_1821);
xor U6726 (N_6726,N_2207,N_3415);
and U6727 (N_6727,N_149,N_3274);
and U6728 (N_6728,N_4680,N_3537);
and U6729 (N_6729,N_2799,N_4638);
nand U6730 (N_6730,N_1723,N_4447);
nor U6731 (N_6731,N_219,N_3026);
nor U6732 (N_6732,N_4244,N_4285);
and U6733 (N_6733,N_4039,N_365);
xnor U6734 (N_6734,N_4809,N_4658);
nand U6735 (N_6735,N_2108,N_4718);
xnor U6736 (N_6736,N_439,N_144);
nor U6737 (N_6737,N_2556,N_2326);
or U6738 (N_6738,N_3899,N_4194);
xor U6739 (N_6739,N_888,N_4675);
nor U6740 (N_6740,N_2080,N_4666);
and U6741 (N_6741,N_1554,N_442);
nand U6742 (N_6742,N_4943,N_2763);
xnor U6743 (N_6743,N_3419,N_1175);
nand U6744 (N_6744,N_267,N_3053);
nor U6745 (N_6745,N_4891,N_684);
and U6746 (N_6746,N_3488,N_4987);
or U6747 (N_6747,N_2360,N_3703);
xnor U6748 (N_6748,N_3952,N_2105);
or U6749 (N_6749,N_1520,N_4335);
nor U6750 (N_6750,N_515,N_1766);
nand U6751 (N_6751,N_4756,N_2349);
and U6752 (N_6752,N_2636,N_4204);
nor U6753 (N_6753,N_1284,N_4396);
or U6754 (N_6754,N_1382,N_3775);
nand U6755 (N_6755,N_320,N_3696);
xor U6756 (N_6756,N_2543,N_938);
and U6757 (N_6757,N_3598,N_3746);
and U6758 (N_6758,N_1970,N_2098);
nor U6759 (N_6759,N_2227,N_1747);
and U6760 (N_6760,N_4677,N_145);
and U6761 (N_6761,N_4581,N_717);
xnor U6762 (N_6762,N_918,N_2022);
nand U6763 (N_6763,N_28,N_2792);
and U6764 (N_6764,N_234,N_3660);
nor U6765 (N_6765,N_3202,N_2967);
xor U6766 (N_6766,N_501,N_2608);
and U6767 (N_6767,N_1152,N_3290);
nand U6768 (N_6768,N_3803,N_1462);
nand U6769 (N_6769,N_4438,N_2383);
nor U6770 (N_6770,N_2385,N_4021);
or U6771 (N_6771,N_292,N_1130);
xnor U6772 (N_6772,N_4911,N_157);
and U6773 (N_6773,N_3970,N_590);
or U6774 (N_6774,N_3001,N_4401);
nor U6775 (N_6775,N_3087,N_3659);
xor U6776 (N_6776,N_1858,N_1039);
nor U6777 (N_6777,N_3917,N_560);
nand U6778 (N_6778,N_564,N_616);
and U6779 (N_6779,N_430,N_4499);
or U6780 (N_6780,N_4610,N_1583);
and U6781 (N_6781,N_4094,N_168);
nor U6782 (N_6782,N_1692,N_4061);
nor U6783 (N_6783,N_3601,N_3167);
nand U6784 (N_6784,N_3942,N_482);
nor U6785 (N_6785,N_4115,N_4709);
or U6786 (N_6786,N_2351,N_2013);
nand U6787 (N_6787,N_1565,N_4026);
and U6788 (N_6788,N_3340,N_3968);
xor U6789 (N_6789,N_2811,N_1993);
xor U6790 (N_6790,N_4562,N_1282);
or U6791 (N_6791,N_1333,N_288);
nor U6792 (N_6792,N_4362,N_3854);
or U6793 (N_6793,N_1652,N_3809);
nand U6794 (N_6794,N_3283,N_2600);
nor U6795 (N_6795,N_1567,N_2680);
and U6796 (N_6796,N_654,N_247);
or U6797 (N_6797,N_4596,N_4177);
and U6798 (N_6798,N_1961,N_4557);
nor U6799 (N_6799,N_1932,N_583);
nand U6800 (N_6800,N_1278,N_3737);
nor U6801 (N_6801,N_3648,N_2348);
nand U6802 (N_6802,N_2482,N_1971);
or U6803 (N_6803,N_1426,N_1341);
and U6804 (N_6804,N_4606,N_620);
nor U6805 (N_6805,N_3061,N_1203);
nor U6806 (N_6806,N_3013,N_2379);
and U6807 (N_6807,N_4525,N_942);
nand U6808 (N_6808,N_2213,N_3650);
and U6809 (N_6809,N_4348,N_4739);
and U6810 (N_6810,N_3581,N_2697);
nand U6811 (N_6811,N_1491,N_2679);
and U6812 (N_6812,N_3551,N_3975);
and U6813 (N_6813,N_4560,N_4129);
or U6814 (N_6814,N_4215,N_3377);
or U6815 (N_6815,N_712,N_2487);
and U6816 (N_6816,N_4669,N_1788);
nand U6817 (N_6817,N_104,N_409);
nand U6818 (N_6818,N_2340,N_4453);
xnor U6819 (N_6819,N_3799,N_4222);
xor U6820 (N_6820,N_1978,N_4434);
nand U6821 (N_6821,N_2215,N_227);
xnor U6822 (N_6822,N_1729,N_3209);
and U6823 (N_6823,N_4467,N_2586);
nor U6824 (N_6824,N_2432,N_4576);
or U6825 (N_6825,N_822,N_1835);
nor U6826 (N_6826,N_4154,N_1724);
and U6827 (N_6827,N_3334,N_1719);
and U6828 (N_6828,N_1330,N_3934);
xnor U6829 (N_6829,N_3154,N_3614);
or U6830 (N_6830,N_3649,N_578);
nor U6831 (N_6831,N_4143,N_4289);
nand U6832 (N_6832,N_2585,N_2240);
xor U6833 (N_6833,N_3830,N_1146);
nor U6834 (N_6834,N_2412,N_4713);
and U6835 (N_6835,N_3892,N_1641);
or U6836 (N_6836,N_3345,N_2993);
nor U6837 (N_6837,N_1482,N_4652);
nor U6838 (N_6838,N_4821,N_2311);
xnor U6839 (N_6839,N_4752,N_2061);
or U6840 (N_6840,N_4662,N_3539);
or U6841 (N_6841,N_1267,N_4732);
xor U6842 (N_6842,N_3454,N_3278);
xnor U6843 (N_6843,N_110,N_2037);
or U6844 (N_6844,N_1135,N_1276);
nand U6845 (N_6845,N_1281,N_2959);
nor U6846 (N_6846,N_3105,N_2183);
nand U6847 (N_6847,N_779,N_4424);
xor U6848 (N_6848,N_3627,N_3597);
or U6849 (N_6849,N_285,N_2182);
and U6850 (N_6850,N_645,N_4538);
and U6851 (N_6851,N_3025,N_4740);
or U6852 (N_6852,N_75,N_4006);
nand U6853 (N_6853,N_186,N_2219);
nand U6854 (N_6854,N_2144,N_3889);
xnor U6855 (N_6855,N_4595,N_4398);
nor U6856 (N_6856,N_2981,N_3176);
nor U6857 (N_6857,N_443,N_2809);
nand U6858 (N_6858,N_4814,N_150);
nand U6859 (N_6859,N_2910,N_3580);
or U6860 (N_6860,N_4961,N_3343);
and U6861 (N_6861,N_74,N_465);
and U6862 (N_6862,N_535,N_3657);
nor U6863 (N_6863,N_3873,N_2193);
or U6864 (N_6864,N_4186,N_2328);
nand U6865 (N_6865,N_3772,N_2797);
and U6866 (N_6866,N_1248,N_3375);
or U6867 (N_6867,N_102,N_3175);
xnor U6868 (N_6868,N_3824,N_138);
nand U6869 (N_6869,N_1707,N_2617);
nor U6870 (N_6870,N_1148,N_4346);
and U6871 (N_6871,N_769,N_3851);
and U6872 (N_6872,N_2648,N_3316);
nand U6873 (N_6873,N_909,N_2320);
and U6874 (N_6874,N_3595,N_4182);
or U6875 (N_6875,N_1704,N_4805);
nand U6876 (N_6876,N_2082,N_1415);
nand U6877 (N_6877,N_4567,N_8);
nand U6878 (N_6878,N_3624,N_1994);
or U6879 (N_6879,N_1563,N_1752);
or U6880 (N_6880,N_3546,N_1022);
nand U6881 (N_6881,N_4036,N_2736);
nand U6882 (N_6882,N_3924,N_2738);
nor U6883 (N_6883,N_4122,N_2921);
xor U6884 (N_6884,N_1541,N_622);
nand U6885 (N_6885,N_3153,N_680);
or U6886 (N_6886,N_3638,N_11);
nand U6887 (N_6887,N_3360,N_4772);
or U6888 (N_6888,N_4578,N_898);
and U6889 (N_6889,N_2856,N_915);
and U6890 (N_6890,N_510,N_2570);
nor U6891 (N_6891,N_960,N_194);
nand U6892 (N_6892,N_4057,N_3188);
or U6893 (N_6893,N_3634,N_4873);
and U6894 (N_6894,N_1762,N_568);
or U6895 (N_6895,N_1122,N_570);
nor U6896 (N_6896,N_3726,N_4918);
or U6897 (N_6897,N_480,N_1256);
and U6898 (N_6898,N_2363,N_2500);
and U6899 (N_6899,N_3815,N_3183);
and U6900 (N_6900,N_1045,N_3428);
nand U6901 (N_6901,N_4185,N_414);
nor U6902 (N_6902,N_4818,N_2332);
nand U6903 (N_6903,N_1100,N_1310);
nor U6904 (N_6904,N_1521,N_2382);
or U6905 (N_6905,N_58,N_781);
or U6906 (N_6906,N_1540,N_3463);
nor U6907 (N_6907,N_1049,N_2866);
nand U6908 (N_6908,N_4,N_1314);
xnor U6909 (N_6909,N_372,N_3348);
nand U6910 (N_6910,N_4860,N_56);
and U6911 (N_6911,N_4810,N_1760);
nor U6912 (N_6912,N_3910,N_1402);
nand U6913 (N_6913,N_133,N_3871);
nand U6914 (N_6914,N_3795,N_792);
nor U6915 (N_6915,N_2490,N_1656);
nand U6916 (N_6916,N_2902,N_1204);
nor U6917 (N_6917,N_4561,N_730);
and U6918 (N_6918,N_3297,N_2832);
or U6919 (N_6919,N_1018,N_3812);
nand U6920 (N_6920,N_1613,N_97);
nor U6921 (N_6921,N_4661,N_4633);
nor U6922 (N_6922,N_2975,N_1705);
or U6923 (N_6923,N_1863,N_3020);
nand U6924 (N_6924,N_4535,N_2370);
nand U6925 (N_6925,N_569,N_4519);
nor U6926 (N_6926,N_1208,N_1342);
nor U6927 (N_6927,N_1422,N_2345);
nor U6928 (N_6928,N_3164,N_4433);
or U6929 (N_6929,N_4676,N_529);
and U6930 (N_6930,N_2702,N_2801);
nand U6931 (N_6931,N_424,N_2143);
or U6932 (N_6932,N_4993,N_2717);
nand U6933 (N_6933,N_4156,N_2885);
xnor U6934 (N_6934,N_4421,N_184);
and U6935 (N_6935,N_4395,N_4627);
and U6936 (N_6936,N_1615,N_3409);
nor U6937 (N_6937,N_2649,N_4020);
and U6938 (N_6938,N_4510,N_3513);
or U6939 (N_6939,N_1748,N_1299);
xor U6940 (N_6940,N_1922,N_3693);
nand U6941 (N_6941,N_1823,N_2033);
nand U6942 (N_6942,N_632,N_1919);
or U6943 (N_6943,N_4199,N_2948);
or U6944 (N_6944,N_2109,N_1079);
and U6945 (N_6945,N_3121,N_2361);
or U6946 (N_6946,N_1258,N_1136);
nor U6947 (N_6947,N_350,N_4168);
nor U6948 (N_6948,N_2610,N_3210);
nor U6949 (N_6949,N_1494,N_1149);
nand U6950 (N_6950,N_2521,N_3800);
or U6951 (N_6951,N_1320,N_420);
nand U6952 (N_6952,N_998,N_1348);
xor U6953 (N_6953,N_1935,N_2941);
nor U6954 (N_6954,N_3744,N_271);
or U6955 (N_6955,N_815,N_1270);
or U6956 (N_6956,N_864,N_29);
or U6957 (N_6957,N_2419,N_374);
nor U6958 (N_6958,N_3163,N_1298);
or U6959 (N_6959,N_225,N_727);
nand U6960 (N_6960,N_2028,N_2734);
and U6961 (N_6961,N_3959,N_3237);
and U6962 (N_6962,N_4363,N_1178);
nor U6963 (N_6963,N_4647,N_4096);
or U6964 (N_6964,N_695,N_2125);
nand U6965 (N_6965,N_202,N_4407);
nor U6966 (N_6966,N_803,N_2423);
or U6967 (N_6967,N_1840,N_4665);
and U6968 (N_6968,N_390,N_3524);
and U6969 (N_6969,N_2838,N_2635);
nor U6970 (N_6970,N_4146,N_1936);
xor U6971 (N_6971,N_367,N_1789);
or U6972 (N_6972,N_3095,N_3455);
nor U6973 (N_6973,N_4997,N_750);
or U6974 (N_6974,N_1222,N_4893);
and U6975 (N_6975,N_559,N_1966);
or U6976 (N_6976,N_4620,N_4134);
and U6977 (N_6977,N_3992,N_3003);
nor U6978 (N_6978,N_4791,N_820);
nand U6979 (N_6979,N_4890,N_1814);
nand U6980 (N_6980,N_4786,N_2427);
or U6981 (N_6981,N_1421,N_2032);
nor U6982 (N_6982,N_3585,N_59);
or U6983 (N_6983,N_3076,N_452);
and U6984 (N_6984,N_1495,N_2684);
nor U6985 (N_6985,N_2700,N_3974);
nor U6986 (N_6986,N_3255,N_4865);
nand U6987 (N_6987,N_1905,N_1190);
nor U6988 (N_6988,N_340,N_1500);
xor U6989 (N_6989,N_1576,N_4711);
xnor U6990 (N_6990,N_786,N_3662);
nand U6991 (N_6991,N_4192,N_3587);
nand U6992 (N_6992,N_3241,N_813);
and U6993 (N_6993,N_3691,N_1849);
nand U6994 (N_6994,N_994,N_324);
nand U6995 (N_6995,N_3406,N_4130);
or U6996 (N_6996,N_3269,N_2991);
and U6997 (N_6997,N_608,N_948);
and U6998 (N_6998,N_756,N_657);
nand U6999 (N_6999,N_3521,N_4144);
xor U7000 (N_7000,N_369,N_468);
or U7001 (N_7001,N_1867,N_2627);
xor U7002 (N_7002,N_1120,N_2473);
and U7003 (N_7003,N_884,N_1815);
or U7004 (N_7004,N_2973,N_3565);
nor U7005 (N_7005,N_4608,N_588);
xnor U7006 (N_7006,N_4852,N_171);
nand U7007 (N_7007,N_4915,N_68);
or U7008 (N_7008,N_3131,N_3206);
nand U7009 (N_7009,N_954,N_1068);
or U7010 (N_7010,N_1187,N_4214);
and U7011 (N_7011,N_3311,N_410);
or U7012 (N_7012,N_2245,N_4101);
nor U7013 (N_7013,N_1275,N_1305);
and U7014 (N_7014,N_298,N_621);
or U7015 (N_7015,N_1633,N_1702);
nand U7016 (N_7016,N_1312,N_344);
and U7017 (N_7017,N_38,N_2583);
and U7018 (N_7018,N_1019,N_4203);
nand U7019 (N_7019,N_2002,N_1624);
nand U7020 (N_7020,N_3482,N_1114);
and U7021 (N_7021,N_3497,N_2246);
nand U7022 (N_7022,N_2532,N_844);
nand U7023 (N_7023,N_1657,N_935);
nand U7024 (N_7024,N_3907,N_2732);
or U7025 (N_7025,N_4559,N_776);
or U7026 (N_7026,N_4875,N_850);
xnor U7027 (N_7027,N_2633,N_1000);
or U7028 (N_7028,N_558,N_1976);
and U7029 (N_7029,N_506,N_3189);
nand U7030 (N_7030,N_1546,N_2605);
nand U7031 (N_7031,N_2039,N_2498);
nand U7032 (N_7032,N_2331,N_1798);
and U7033 (N_7033,N_4700,N_816);
and U7034 (N_7034,N_2131,N_4823);
and U7035 (N_7035,N_1192,N_1987);
and U7036 (N_7036,N_725,N_89);
xor U7037 (N_7037,N_1026,N_2463);
nand U7038 (N_7038,N_248,N_4524);
or U7039 (N_7039,N_1399,N_4293);
nor U7040 (N_7040,N_487,N_3993);
nor U7041 (N_7041,N_1450,N_4674);
or U7042 (N_7042,N_4005,N_1828);
nor U7043 (N_7043,N_2666,N_2408);
nand U7044 (N_7044,N_2971,N_348);
nor U7045 (N_7045,N_1375,N_1055);
nor U7046 (N_7046,N_2169,N_299);
or U7047 (N_7047,N_4982,N_567);
or U7048 (N_7048,N_3708,N_587);
and U7049 (N_7049,N_273,N_2826);
or U7050 (N_7050,N_2384,N_860);
and U7051 (N_7051,N_3759,N_1878);
nor U7052 (N_7052,N_1083,N_277);
or U7053 (N_7053,N_3902,N_4639);
xor U7054 (N_7054,N_2950,N_2664);
nand U7055 (N_7055,N_4068,N_4488);
and U7056 (N_7056,N_1147,N_2220);
nand U7057 (N_7057,N_847,N_4492);
xor U7058 (N_7058,N_2598,N_4357);
nor U7059 (N_7059,N_1997,N_122);
and U7060 (N_7060,N_4755,N_3891);
nand U7061 (N_7061,N_214,N_99);
and U7062 (N_7062,N_4478,N_4197);
nand U7063 (N_7063,N_4319,N_1552);
and U7064 (N_7064,N_2845,N_2093);
and U7065 (N_7065,N_259,N_3058);
nand U7066 (N_7066,N_3527,N_1206);
and U7067 (N_7067,N_3041,N_3099);
or U7068 (N_7068,N_1406,N_2813);
or U7069 (N_7069,N_4281,N_3092);
or U7070 (N_7070,N_3625,N_999);
nor U7071 (N_7071,N_3015,N_4477);
and U7072 (N_7072,N_2696,N_4795);
and U7073 (N_7073,N_3392,N_855);
nand U7074 (N_7074,N_1309,N_3081);
nand U7075 (N_7075,N_2313,N_3004);
and U7076 (N_7076,N_1339,N_3172);
nor U7077 (N_7077,N_4549,N_1530);
and U7078 (N_7078,N_1794,N_597);
nor U7079 (N_7079,N_3989,N_2642);
nor U7080 (N_7080,N_4886,N_517);
nor U7081 (N_7081,N_4495,N_3927);
or U7082 (N_7082,N_1718,N_31);
nor U7083 (N_7083,N_3203,N_985);
or U7084 (N_7084,N_552,N_2562);
or U7085 (N_7085,N_4565,N_693);
or U7086 (N_7086,N_2132,N_1796);
or U7087 (N_7087,N_2719,N_4391);
nand U7088 (N_7088,N_977,N_158);
nand U7089 (N_7089,N_2416,N_4863);
nand U7090 (N_7090,N_2926,N_2145);
or U7091 (N_7091,N_400,N_406);
nor U7092 (N_7092,N_2253,N_3266);
xnor U7093 (N_7093,N_3765,N_2342);
nor U7094 (N_7094,N_2916,N_2117);
and U7095 (N_7095,N_2122,N_3683);
nand U7096 (N_7096,N_4679,N_2923);
or U7097 (N_7097,N_4807,N_2138);
nand U7098 (N_7098,N_1945,N_4544);
xnor U7099 (N_7099,N_3216,N_1879);
or U7100 (N_7100,N_3145,N_1308);
or U7101 (N_7101,N_4858,N_897);
nand U7102 (N_7102,N_209,N_2877);
nor U7103 (N_7103,N_4439,N_503);
xnor U7104 (N_7104,N_1478,N_1033);
or U7105 (N_7105,N_4082,N_3711);
and U7106 (N_7106,N_4897,N_427);
nor U7107 (N_7107,N_576,N_2920);
or U7108 (N_7108,N_733,N_2128);
and U7109 (N_7109,N_1881,N_1757);
and U7110 (N_7110,N_401,N_1743);
xnor U7111 (N_7111,N_4455,N_4673);
or U7112 (N_7112,N_1942,N_396);
or U7113 (N_7113,N_3930,N_3506);
nand U7114 (N_7114,N_1670,N_2951);
xor U7115 (N_7115,N_4132,N_3044);
nor U7116 (N_7116,N_3735,N_461);
and U7117 (N_7117,N_4880,N_2949);
nor U7118 (N_7118,N_4577,N_3103);
xor U7119 (N_7119,N_2651,N_3272);
nor U7120 (N_7120,N_2151,N_2234);
and U7121 (N_7121,N_393,N_663);
and U7122 (N_7122,N_3326,N_4457);
nand U7123 (N_7123,N_4870,N_3646);
nor U7124 (N_7124,N_2435,N_4331);
nand U7125 (N_7125,N_4278,N_241);
or U7126 (N_7126,N_4208,N_1331);
or U7127 (N_7127,N_2314,N_1107);
nor U7128 (N_7128,N_586,N_4774);
and U7129 (N_7129,N_861,N_4147);
nor U7130 (N_7130,N_1129,N_1496);
nand U7131 (N_7131,N_3122,N_333);
and U7132 (N_7132,N_1165,N_652);
or U7133 (N_7133,N_602,N_1699);
nor U7134 (N_7134,N_2510,N_2307);
nand U7135 (N_7135,N_1594,N_1771);
or U7136 (N_7136,N_4534,N_2208);
nand U7137 (N_7137,N_3469,N_4553);
and U7138 (N_7138,N_3874,N_1568);
nor U7139 (N_7139,N_1946,N_4359);
or U7140 (N_7140,N_3462,N_2924);
and U7141 (N_7141,N_2406,N_3010);
and U7142 (N_7142,N_2676,N_926);
xor U7143 (N_7143,N_681,N_2347);
nand U7144 (N_7144,N_1058,N_7);
or U7145 (N_7145,N_4985,N_757);
and U7146 (N_7146,N_1335,N_3363);
or U7147 (N_7147,N_4785,N_963);
nand U7148 (N_7148,N_2027,N_2429);
nor U7149 (N_7149,N_1216,N_3268);
or U7150 (N_7150,N_2571,N_532);
xnor U7151 (N_7151,N_4253,N_2814);
xnor U7152 (N_7152,N_709,N_4936);
nor U7153 (N_7153,N_4110,N_659);
nor U7154 (N_7154,N_303,N_3438);
and U7155 (N_7155,N_3437,N_1134);
nand U7156 (N_7156,N_1505,N_676);
and U7157 (N_7157,N_1066,N_2514);
or U7158 (N_7158,N_53,N_4217);
or U7159 (N_7159,N_4428,N_4411);
nor U7160 (N_7160,N_450,N_2114);
nand U7161 (N_7161,N_2146,N_1327);
nor U7162 (N_7162,N_3093,N_1127);
nand U7163 (N_7163,N_4383,N_585);
xor U7164 (N_7164,N_3692,N_1639);
and U7165 (N_7165,N_3796,N_246);
and U7166 (N_7166,N_1313,N_4851);
nor U7167 (N_7167,N_814,N_670);
and U7168 (N_7168,N_641,N_1255);
nor U7169 (N_7169,N_3990,N_1156);
or U7170 (N_7170,N_2771,N_2263);
and U7171 (N_7171,N_2900,N_4959);
or U7172 (N_7172,N_4223,N_656);
or U7173 (N_7173,N_806,N_3276);
or U7174 (N_7174,N_3444,N_4601);
and U7175 (N_7175,N_1963,N_4145);
nand U7176 (N_7176,N_1002,N_2802);
nor U7177 (N_7177,N_2854,N_1455);
nor U7178 (N_7178,N_1790,N_2262);
nor U7179 (N_7179,N_3449,N_1430);
nand U7180 (N_7180,N_2592,N_1749);
nor U7181 (N_7181,N_4604,N_1448);
nor U7182 (N_7182,N_862,N_5);
or U7183 (N_7183,N_3936,N_3155);
xnor U7184 (N_7184,N_1572,N_2849);
and U7185 (N_7185,N_2269,N_3191);
nor U7186 (N_7186,N_4248,N_2499);
xor U7187 (N_7187,N_1246,N_1063);
nand U7188 (N_7188,N_3554,N_1145);
or U7189 (N_7189,N_2972,N_4776);
and U7190 (N_7190,N_240,N_4948);
nor U7191 (N_7191,N_45,N_392);
nand U7192 (N_7192,N_742,N_4912);
xnor U7193 (N_7193,N_4636,N_1467);
and U7194 (N_7194,N_2806,N_263);
and U7195 (N_7195,N_4100,N_3562);
and U7196 (N_7196,N_2235,N_1587);
and U7197 (N_7197,N_628,N_2134);
nand U7198 (N_7198,N_790,N_1459);
and U7199 (N_7199,N_561,N_3256);
nand U7200 (N_7200,N_2883,N_2815);
or U7201 (N_7201,N_1069,N_2911);
nand U7202 (N_7202,N_2834,N_1677);
nand U7203 (N_7203,N_336,N_4266);
and U7204 (N_7204,N_892,N_3282);
nand U7205 (N_7205,N_1889,N_3499);
or U7206 (N_7206,N_1774,N_262);
and U7207 (N_7207,N_3672,N_572);
nor U7208 (N_7208,N_4460,N_4261);
and U7209 (N_7209,N_1042,N_4001);
and U7210 (N_7210,N_2292,N_379);
nor U7211 (N_7211,N_952,N_3018);
nand U7212 (N_7212,N_801,N_605);
or U7213 (N_7213,N_4437,N_2559);
nor U7214 (N_7214,N_3850,N_4765);
or U7215 (N_7215,N_226,N_1126);
and U7216 (N_7216,N_2084,N_3784);
nor U7217 (N_7217,N_1024,N_754);
xor U7218 (N_7218,N_2688,N_1223);
or U7219 (N_7219,N_3248,N_3486);
and U7220 (N_7220,N_339,N_2964);
nor U7221 (N_7221,N_3855,N_3100);
or U7222 (N_7222,N_4523,N_1869);
xnor U7223 (N_7223,N_3783,N_4241);
nand U7224 (N_7224,N_3553,N_1607);
or U7225 (N_7225,N_4083,N_4345);
and U7226 (N_7226,N_164,N_3616);
xnor U7227 (N_7227,N_3678,N_2042);
and U7228 (N_7228,N_190,N_1949);
nand U7229 (N_7229,N_2663,N_665);
or U7230 (N_7230,N_37,N_108);
nand U7231 (N_7231,N_4323,N_3723);
nand U7232 (N_7232,N_4069,N_3096);
and U7233 (N_7233,N_2693,N_287);
and U7234 (N_7234,N_3359,N_294);
or U7235 (N_7235,N_261,N_929);
or U7236 (N_7236,N_301,N_4882);
xnor U7237 (N_7237,N_3991,N_1128);
nor U7238 (N_7238,N_302,N_380);
or U7239 (N_7239,N_2238,N_1598);
nor U7240 (N_7240,N_2915,N_819);
nor U7241 (N_7241,N_4625,N_2069);
and U7242 (N_7242,N_4250,N_3550);
xor U7243 (N_7243,N_4483,N_4033);
nor U7244 (N_7244,N_4640,N_1658);
nand U7245 (N_7245,N_2846,N_2955);
nand U7246 (N_7246,N_1991,N_2897);
nor U7247 (N_7247,N_236,N_495);
nand U7248 (N_7248,N_4671,N_3091);
or U7249 (N_7249,N_1197,N_1983);
nand U7250 (N_7250,N_3501,N_845);
xor U7251 (N_7251,N_1982,N_893);
or U7252 (N_7252,N_3361,N_879);
or U7253 (N_7253,N_4551,N_4955);
nand U7254 (N_7254,N_4473,N_2862);
or U7255 (N_7255,N_1036,N_3198);
nor U7256 (N_7256,N_2713,N_4683);
nand U7257 (N_7257,N_4695,N_1668);
nor U7258 (N_7258,N_2470,N_1273);
or U7259 (N_7259,N_759,N_726);
and U7260 (N_7260,N_2557,N_4588);
nand U7261 (N_7261,N_3344,N_208);
nor U7262 (N_7262,N_1578,N_2339);
or U7263 (N_7263,N_1417,N_497);
and U7264 (N_7264,N_1395,N_3106);
or U7265 (N_7265,N_76,N_1611);
xor U7266 (N_7266,N_1679,N_364);
nor U7267 (N_7267,N_4302,N_3422);
or U7268 (N_7268,N_4237,N_4619);
and U7269 (N_7269,N_683,N_2668);
or U7270 (N_7270,N_4276,N_1323);
and U7271 (N_7271,N_4449,N_3724);
nand U7272 (N_7272,N_1865,N_4901);
nand U7273 (N_7273,N_2359,N_3656);
nor U7274 (N_7274,N_2325,N_201);
nor U7275 (N_7275,N_2298,N_1043);
nand U7276 (N_7276,N_3599,N_868);
nor U7277 (N_7277,N_1168,N_4270);
xnor U7278 (N_7278,N_1634,N_3541);
nand U7279 (N_7279,N_4228,N_3079);
nand U7280 (N_7280,N_3124,N_2335);
and U7281 (N_7281,N_504,N_113);
or U7282 (N_7282,N_4356,N_2485);
and U7283 (N_7283,N_3066,N_451);
or U7284 (N_7284,N_3214,N_1219);
and U7285 (N_7285,N_4960,N_4180);
nand U7286 (N_7286,N_3617,N_3397);
or U7287 (N_7287,N_804,N_2079);
nand U7288 (N_7288,N_160,N_958);
nand U7289 (N_7289,N_2830,N_705);
or U7290 (N_7290,N_2495,N_2720);
and U7291 (N_7291,N_4300,N_4672);
or U7292 (N_7292,N_2743,N_4308);
and U7293 (N_7293,N_3591,N_3325);
nor U7294 (N_7294,N_2461,N_279);
nor U7295 (N_7295,N_4813,N_4768);
and U7296 (N_7296,N_2744,N_4406);
or U7297 (N_7297,N_4991,N_3404);
nand U7298 (N_7298,N_1189,N_1432);
or U7299 (N_7299,N_3090,N_1251);
or U7300 (N_7300,N_136,N_447);
or U7301 (N_7301,N_3996,N_1264);
and U7302 (N_7302,N_2062,N_4207);
xor U7303 (N_7303,N_422,N_1589);
nand U7304 (N_7304,N_3401,N_2203);
and U7305 (N_7305,N_3523,N_4788);
or U7306 (N_7306,N_4048,N_1843);
nand U7307 (N_7307,N_1301,N_4819);
or U7308 (N_7308,N_1444,N_4799);
nor U7309 (N_7309,N_1638,N_478);
nor U7310 (N_7310,N_2149,N_1620);
and U7311 (N_7311,N_4095,N_2434);
nand U7312 (N_7312,N_3347,N_2612);
or U7313 (N_7313,N_1368,N_1799);
and U7314 (N_7314,N_1502,N_3324);
nor U7315 (N_7315,N_1109,N_584);
nand U7316 (N_7316,N_66,N_3702);
nor U7317 (N_7317,N_229,N_1923);
and U7318 (N_7318,N_275,N_4124);
and U7319 (N_7319,N_2922,N_4771);
nand U7320 (N_7320,N_3253,N_4417);
xor U7321 (N_7321,N_771,N_3699);
nand U7322 (N_7322,N_2251,N_2677);
or U7323 (N_7323,N_3933,N_4603);
and U7324 (N_7324,N_4002,N_4621);
xor U7325 (N_7325,N_1694,N_4272);
and U7326 (N_7326,N_4088,N_896);
xor U7327 (N_7327,N_4935,N_1630);
nor U7328 (N_7328,N_1098,N_2366);
nor U7329 (N_7329,N_734,N_2476);
nand U7330 (N_7330,N_638,N_1428);
and U7331 (N_7331,N_834,N_3069);
nor U7332 (N_7332,N_3115,N_3714);
and U7333 (N_7333,N_1396,N_2690);
nor U7334 (N_7334,N_3987,N_4404);
nor U7335 (N_7335,N_2466,N_4427);
xor U7336 (N_7336,N_2999,N_3190);
nand U7337 (N_7337,N_4536,N_3306);
nand U7338 (N_7338,N_3832,N_937);
nand U7339 (N_7339,N_1117,N_1486);
or U7340 (N_7340,N_2582,N_1785);
nor U7341 (N_7341,N_4612,N_4141);
nand U7342 (N_7342,N_664,N_4689);
and U7343 (N_7343,N_1626,N_4593);
nor U7344 (N_7344,N_3055,N_4016);
or U7345 (N_7345,N_1562,N_49);
or U7346 (N_7346,N_650,N_700);
nand U7347 (N_7347,N_2161,N_1453);
nor U7348 (N_7348,N_4754,N_1103);
nand U7349 (N_7349,N_1802,N_13);
or U7350 (N_7350,N_1732,N_3558);
nand U7351 (N_7351,N_2031,N_1513);
or U7352 (N_7352,N_682,N_2982);
or U7353 (N_7353,N_1352,N_3569);
nor U7354 (N_7354,N_2947,N_796);
nor U7355 (N_7355,N_3178,N_4957);
nand U7356 (N_7356,N_2749,N_3661);
and U7357 (N_7357,N_1726,N_2064);
nor U7358 (N_7358,N_1733,N_1892);
nand U7359 (N_7359,N_3825,N_1316);
or U7360 (N_7360,N_4653,N_4251);
or U7361 (N_7361,N_1550,N_4408);
xor U7362 (N_7362,N_3388,N_1890);
xnor U7363 (N_7363,N_3767,N_32);
nand U7364 (N_7364,N_1131,N_1959);
and U7365 (N_7365,N_1294,N_2044);
and U7366 (N_7366,N_2303,N_4157);
nor U7367 (N_7367,N_4705,N_3498);
and U7368 (N_7368,N_309,N_812);
nand U7369 (N_7369,N_508,N_4702);
or U7370 (N_7370,N_3897,N_3094);
nor U7371 (N_7371,N_975,N_3046);
nand U7372 (N_7372,N_4419,N_4687);
nand U7373 (N_7373,N_953,N_1451);
xnor U7374 (N_7374,N_3613,N_2988);
and U7375 (N_7375,N_4558,N_118);
nand U7376 (N_7376,N_2976,N_966);
nor U7377 (N_7377,N_870,N_2979);
nor U7378 (N_7378,N_4379,N_232);
or U7379 (N_7379,N_2200,N_4698);
nand U7380 (N_7380,N_3074,N_3374);
nand U7381 (N_7381,N_598,N_1085);
and U7382 (N_7382,N_2992,N_3450);
and U7383 (N_7383,N_1142,N_2019);
nor U7384 (N_7384,N_625,N_2699);
or U7385 (N_7385,N_4903,N_3471);
and U7386 (N_7386,N_3110,N_3384);
or U7387 (N_7387,N_1910,N_4806);
nor U7388 (N_7388,N_3766,N_1650);
or U7389 (N_7389,N_1647,N_1468);
or U7390 (N_7390,N_155,N_1711);
and U7391 (N_7391,N_3468,N_2165);
or U7392 (N_7392,N_114,N_1856);
or U7393 (N_7393,N_2243,N_1901);
nor U7394 (N_7394,N_4716,N_200);
nor U7395 (N_7395,N_4183,N_630);
nand U7396 (N_7396,N_3395,N_1989);
nand U7397 (N_7397,N_2867,N_3476);
and U7398 (N_7398,N_4011,N_772);
or U7399 (N_7399,N_3230,N_2472);
or U7400 (N_7400,N_1188,N_2783);
and U7401 (N_7401,N_4738,N_3821);
or U7402 (N_7402,N_370,N_4103);
or U7403 (N_7403,N_446,N_2100);
nand U7404 (N_7404,N_3893,N_1420);
and U7405 (N_7405,N_2493,N_3193);
nand U7406 (N_7406,N_881,N_748);
nor U7407 (N_7407,N_4054,N_3769);
nor U7408 (N_7408,N_1514,N_2496);
xnor U7409 (N_7409,N_760,N_1250);
and U7410 (N_7410,N_3755,N_1675);
xnor U7411 (N_7411,N_2190,N_2344);
xor U7412 (N_7412,N_2855,N_4109);
and U7413 (N_7413,N_4842,N_3643);
and U7414 (N_7414,N_4468,N_829);
nor U7415 (N_7415,N_3888,N_1672);
or U7416 (N_7416,N_3331,N_2257);
nor U7417 (N_7417,N_1071,N_2173);
or U7418 (N_7418,N_1917,N_3536);
and U7419 (N_7419,N_3390,N_4962);
nand U7420 (N_7420,N_191,N_706);
xnor U7421 (N_7421,N_4582,N_2116);
and U7422 (N_7422,N_1817,N_2295);
or U7423 (N_7423,N_1271,N_2040);
or U7424 (N_7424,N_4758,N_521);
or U7425 (N_7425,N_2770,N_4749);
nor U7426 (N_7426,N_729,N_314);
or U7427 (N_7427,N_2162,N_2365);
nand U7428 (N_7428,N_2953,N_4273);
or U7429 (N_7429,N_1730,N_3908);
and U7430 (N_7430,N_807,N_2810);
xnor U7431 (N_7431,N_432,N_412);
and U7432 (N_7432,N_3584,N_358);
or U7433 (N_7433,N_3260,N_2139);
or U7434 (N_7434,N_1202,N_1123);
nand U7435 (N_7435,N_3694,N_4284);
or U7436 (N_7436,N_4895,N_3063);
and U7437 (N_7437,N_3677,N_1664);
nand U7438 (N_7438,N_3207,N_3481);
xor U7439 (N_7439,N_825,N_876);
and U7440 (N_7440,N_2968,N_1777);
or U7441 (N_7441,N_1001,N_1351);
nor U7442 (N_7442,N_1816,N_4287);
or U7443 (N_7443,N_48,N_4456);
and U7444 (N_7444,N_2179,N_1953);
nor U7445 (N_7445,N_3204,N_2216);
nor U7446 (N_7446,N_2088,N_1636);
nand U7447 (N_7447,N_2467,N_283);
xnor U7448 (N_7448,N_3804,N_3863);
and U7449 (N_7449,N_3709,N_3289);
nor U7450 (N_7450,N_624,N_306);
xnor U7451 (N_7451,N_1980,N_2341);
or U7452 (N_7452,N_3035,N_1958);
nand U7453 (N_7453,N_187,N_3561);
and U7454 (N_7454,N_151,N_3147);
and U7455 (N_7455,N_489,N_1457);
or U7456 (N_7456,N_1803,N_1824);
nor U7457 (N_7457,N_4505,N_2296);
nand U7458 (N_7458,N_2121,N_565);
nor U7459 (N_7459,N_2118,N_1525);
or U7460 (N_7460,N_4844,N_4249);
nand U7461 (N_7461,N_629,N_4574);
nor U7462 (N_7462,N_3685,N_4922);
or U7463 (N_7463,N_1381,N_4605);
nor U7464 (N_7464,N_1427,N_4660);
and U7465 (N_7465,N_2270,N_413);
and U7466 (N_7466,N_566,N_3185);
nand U7467 (N_7467,N_945,N_205);
nand U7468 (N_7468,N_1379,N_2137);
nand U7469 (N_7469,N_4479,N_2865);
and U7470 (N_7470,N_3956,N_458);
and U7471 (N_7471,N_4073,N_2639);
nor U7472 (N_7472,N_4645,N_1812);
nand U7473 (N_7473,N_906,N_1596);
nand U7474 (N_7474,N_4343,N_3964);
nand U7475 (N_7475,N_3078,N_1463);
nor U7476 (N_7476,N_4243,N_4235);
nand U7477 (N_7477,N_415,N_2099);
nand U7478 (N_7478,N_1081,N_1603);
xnor U7479 (N_7479,N_87,N_612);
xor U7480 (N_7480,N_3368,N_3791);
nor U7481 (N_7481,N_4548,N_903);
nor U7482 (N_7482,N_543,N_4949);
nand U7483 (N_7483,N_1400,N_1501);
xor U7484 (N_7484,N_2567,N_2399);
or U7485 (N_7485,N_4232,N_4720);
or U7486 (N_7486,N_3556,N_4977);
or U7487 (N_7487,N_1767,N_418);
or U7488 (N_7488,N_4688,N_3725);
or U7489 (N_7489,N_2533,N_3329);
nand U7490 (N_7490,N_4074,N_2527);
or U7491 (N_7491,N_1851,N_851);
nor U7492 (N_7492,N_4097,N_2305);
and U7493 (N_7493,N_4298,N_4714);
or U7494 (N_7494,N_2604,N_2698);
and U7495 (N_7495,N_1710,N_2177);
nor U7496 (N_7496,N_55,N_2786);
or U7497 (N_7497,N_217,N_4336);
or U7498 (N_7498,N_842,N_3674);
nor U7499 (N_7499,N_3487,N_3819);
and U7500 (N_7500,N_1322,N_202);
and U7501 (N_7501,N_3830,N_4680);
and U7502 (N_7502,N_4892,N_3359);
nor U7503 (N_7503,N_25,N_2382);
or U7504 (N_7504,N_1815,N_158);
xor U7505 (N_7505,N_4319,N_4322);
nor U7506 (N_7506,N_4304,N_3364);
nor U7507 (N_7507,N_2199,N_4909);
nand U7508 (N_7508,N_151,N_2678);
xor U7509 (N_7509,N_318,N_237);
nor U7510 (N_7510,N_2740,N_3698);
and U7511 (N_7511,N_2703,N_2740);
and U7512 (N_7512,N_378,N_3997);
and U7513 (N_7513,N_2669,N_797);
or U7514 (N_7514,N_2808,N_3629);
nand U7515 (N_7515,N_1942,N_402);
nand U7516 (N_7516,N_2111,N_3088);
or U7517 (N_7517,N_4376,N_4107);
nand U7518 (N_7518,N_1790,N_1794);
nand U7519 (N_7519,N_4584,N_2117);
or U7520 (N_7520,N_3042,N_4842);
and U7521 (N_7521,N_4824,N_385);
xor U7522 (N_7522,N_557,N_2398);
nand U7523 (N_7523,N_4035,N_3607);
nand U7524 (N_7524,N_2891,N_3647);
or U7525 (N_7525,N_218,N_4211);
nand U7526 (N_7526,N_1306,N_3990);
nand U7527 (N_7527,N_1695,N_178);
or U7528 (N_7528,N_1940,N_3260);
and U7529 (N_7529,N_1881,N_4085);
and U7530 (N_7530,N_3886,N_3913);
or U7531 (N_7531,N_239,N_356);
nand U7532 (N_7532,N_276,N_4549);
and U7533 (N_7533,N_3844,N_1829);
and U7534 (N_7534,N_1756,N_1157);
and U7535 (N_7535,N_3208,N_4753);
nand U7536 (N_7536,N_2463,N_1154);
nand U7537 (N_7537,N_1887,N_638);
nand U7538 (N_7538,N_1872,N_4109);
nor U7539 (N_7539,N_965,N_2764);
nor U7540 (N_7540,N_1952,N_2048);
and U7541 (N_7541,N_3753,N_1198);
nor U7542 (N_7542,N_680,N_302);
nand U7543 (N_7543,N_4074,N_1985);
nor U7544 (N_7544,N_245,N_4784);
xnor U7545 (N_7545,N_1253,N_2240);
or U7546 (N_7546,N_4202,N_627);
nor U7547 (N_7547,N_471,N_3274);
or U7548 (N_7548,N_1630,N_4200);
or U7549 (N_7549,N_2439,N_2353);
nand U7550 (N_7550,N_2885,N_617);
and U7551 (N_7551,N_1481,N_4922);
nor U7552 (N_7552,N_4542,N_533);
nor U7553 (N_7553,N_2178,N_2571);
nor U7554 (N_7554,N_3467,N_3394);
nand U7555 (N_7555,N_4820,N_1363);
xor U7556 (N_7556,N_4867,N_3741);
nor U7557 (N_7557,N_871,N_2134);
nand U7558 (N_7558,N_372,N_2995);
or U7559 (N_7559,N_4815,N_3015);
nor U7560 (N_7560,N_1512,N_3892);
nor U7561 (N_7561,N_4192,N_1571);
nor U7562 (N_7562,N_4664,N_2855);
nand U7563 (N_7563,N_499,N_3945);
nand U7564 (N_7564,N_4393,N_1114);
nand U7565 (N_7565,N_3731,N_2084);
nand U7566 (N_7566,N_1383,N_2511);
or U7567 (N_7567,N_1028,N_1159);
nor U7568 (N_7568,N_67,N_4388);
nand U7569 (N_7569,N_4409,N_3010);
and U7570 (N_7570,N_2310,N_2794);
xnor U7571 (N_7571,N_3295,N_3890);
or U7572 (N_7572,N_3893,N_3214);
nand U7573 (N_7573,N_4373,N_1588);
nor U7574 (N_7574,N_2470,N_1183);
and U7575 (N_7575,N_1398,N_4015);
or U7576 (N_7576,N_4852,N_3346);
xor U7577 (N_7577,N_4275,N_499);
nand U7578 (N_7578,N_507,N_923);
nand U7579 (N_7579,N_299,N_4002);
nand U7580 (N_7580,N_3462,N_2050);
or U7581 (N_7581,N_3993,N_2472);
nor U7582 (N_7582,N_2915,N_1928);
xnor U7583 (N_7583,N_850,N_2809);
xnor U7584 (N_7584,N_1767,N_4963);
nand U7585 (N_7585,N_4023,N_1930);
or U7586 (N_7586,N_4368,N_1431);
nand U7587 (N_7587,N_4936,N_1385);
or U7588 (N_7588,N_531,N_47);
nor U7589 (N_7589,N_2388,N_2219);
nand U7590 (N_7590,N_2984,N_4367);
nand U7591 (N_7591,N_124,N_2494);
nor U7592 (N_7592,N_1384,N_2174);
and U7593 (N_7593,N_2909,N_3866);
nor U7594 (N_7594,N_1149,N_1477);
and U7595 (N_7595,N_137,N_2864);
or U7596 (N_7596,N_4538,N_3083);
xor U7597 (N_7597,N_2259,N_1790);
xor U7598 (N_7598,N_4072,N_4821);
or U7599 (N_7599,N_2078,N_3688);
nand U7600 (N_7600,N_4995,N_3317);
or U7601 (N_7601,N_2098,N_918);
and U7602 (N_7602,N_245,N_3541);
or U7603 (N_7603,N_980,N_2071);
and U7604 (N_7604,N_986,N_4282);
nor U7605 (N_7605,N_1684,N_2429);
nand U7606 (N_7606,N_1727,N_4746);
xnor U7607 (N_7607,N_2379,N_4282);
xor U7608 (N_7608,N_3264,N_2453);
or U7609 (N_7609,N_4733,N_3957);
xnor U7610 (N_7610,N_4030,N_1790);
or U7611 (N_7611,N_1817,N_4175);
and U7612 (N_7612,N_4529,N_4057);
and U7613 (N_7613,N_973,N_1827);
nor U7614 (N_7614,N_4368,N_1737);
or U7615 (N_7615,N_2595,N_2997);
nor U7616 (N_7616,N_2206,N_1210);
nand U7617 (N_7617,N_1412,N_1180);
or U7618 (N_7618,N_1243,N_1416);
nand U7619 (N_7619,N_3289,N_2770);
or U7620 (N_7620,N_623,N_480);
xor U7621 (N_7621,N_4156,N_2199);
nor U7622 (N_7622,N_1218,N_1713);
xnor U7623 (N_7623,N_2487,N_4345);
and U7624 (N_7624,N_3396,N_3673);
or U7625 (N_7625,N_2954,N_1475);
xnor U7626 (N_7626,N_1070,N_74);
and U7627 (N_7627,N_4204,N_123);
nand U7628 (N_7628,N_3978,N_2851);
nand U7629 (N_7629,N_3866,N_112);
and U7630 (N_7630,N_2855,N_2352);
nor U7631 (N_7631,N_4038,N_4640);
and U7632 (N_7632,N_4474,N_3026);
and U7633 (N_7633,N_4291,N_2376);
nand U7634 (N_7634,N_1011,N_3721);
and U7635 (N_7635,N_900,N_1845);
xor U7636 (N_7636,N_3103,N_3742);
nor U7637 (N_7637,N_3414,N_4538);
or U7638 (N_7638,N_1206,N_2440);
nor U7639 (N_7639,N_3369,N_1448);
nor U7640 (N_7640,N_2920,N_1433);
and U7641 (N_7641,N_3865,N_2205);
nor U7642 (N_7642,N_1194,N_2030);
or U7643 (N_7643,N_1183,N_571);
nor U7644 (N_7644,N_4533,N_522);
or U7645 (N_7645,N_4511,N_4590);
nor U7646 (N_7646,N_3895,N_1607);
and U7647 (N_7647,N_176,N_1746);
or U7648 (N_7648,N_4638,N_2521);
nand U7649 (N_7649,N_311,N_3885);
xnor U7650 (N_7650,N_1499,N_41);
nand U7651 (N_7651,N_3050,N_4119);
and U7652 (N_7652,N_3849,N_2522);
and U7653 (N_7653,N_2455,N_4487);
or U7654 (N_7654,N_1761,N_2825);
or U7655 (N_7655,N_3135,N_3335);
or U7656 (N_7656,N_1597,N_2376);
and U7657 (N_7657,N_319,N_218);
nand U7658 (N_7658,N_1351,N_2785);
nor U7659 (N_7659,N_436,N_4913);
nor U7660 (N_7660,N_859,N_1413);
or U7661 (N_7661,N_4142,N_4355);
and U7662 (N_7662,N_4915,N_3297);
or U7663 (N_7663,N_407,N_3189);
nand U7664 (N_7664,N_3152,N_4634);
or U7665 (N_7665,N_649,N_125);
and U7666 (N_7666,N_2733,N_2554);
nor U7667 (N_7667,N_1862,N_1879);
nor U7668 (N_7668,N_1164,N_2461);
and U7669 (N_7669,N_734,N_533);
nor U7670 (N_7670,N_2996,N_4324);
or U7671 (N_7671,N_4279,N_4266);
xnor U7672 (N_7672,N_4038,N_2106);
or U7673 (N_7673,N_458,N_2741);
nor U7674 (N_7674,N_3262,N_2341);
nand U7675 (N_7675,N_1954,N_3771);
or U7676 (N_7676,N_3526,N_3010);
nand U7677 (N_7677,N_1774,N_1591);
and U7678 (N_7678,N_3298,N_3750);
xnor U7679 (N_7679,N_3167,N_3098);
xnor U7680 (N_7680,N_3176,N_63);
nand U7681 (N_7681,N_1952,N_4370);
or U7682 (N_7682,N_630,N_347);
nor U7683 (N_7683,N_2013,N_4926);
and U7684 (N_7684,N_28,N_3836);
and U7685 (N_7685,N_3596,N_2587);
nand U7686 (N_7686,N_3298,N_1929);
nand U7687 (N_7687,N_3646,N_3513);
xor U7688 (N_7688,N_1203,N_564);
and U7689 (N_7689,N_4700,N_1382);
nor U7690 (N_7690,N_2077,N_12);
xnor U7691 (N_7691,N_499,N_567);
or U7692 (N_7692,N_2228,N_4763);
or U7693 (N_7693,N_3940,N_3589);
nor U7694 (N_7694,N_379,N_3081);
nor U7695 (N_7695,N_4442,N_983);
xor U7696 (N_7696,N_2673,N_545);
nor U7697 (N_7697,N_4351,N_2946);
or U7698 (N_7698,N_4371,N_3233);
or U7699 (N_7699,N_2838,N_2305);
and U7700 (N_7700,N_4707,N_2291);
nor U7701 (N_7701,N_4590,N_1690);
and U7702 (N_7702,N_4855,N_4299);
nor U7703 (N_7703,N_365,N_4779);
and U7704 (N_7704,N_2766,N_2318);
nor U7705 (N_7705,N_3507,N_3924);
nor U7706 (N_7706,N_4992,N_210);
nand U7707 (N_7707,N_4112,N_2572);
nor U7708 (N_7708,N_496,N_1404);
and U7709 (N_7709,N_3712,N_444);
nor U7710 (N_7710,N_3437,N_4297);
and U7711 (N_7711,N_2403,N_723);
xor U7712 (N_7712,N_1769,N_4412);
or U7713 (N_7713,N_2244,N_2053);
or U7714 (N_7714,N_3551,N_1103);
nor U7715 (N_7715,N_4811,N_3693);
and U7716 (N_7716,N_42,N_3138);
or U7717 (N_7717,N_2975,N_4134);
nor U7718 (N_7718,N_2884,N_4676);
and U7719 (N_7719,N_1102,N_4844);
nor U7720 (N_7720,N_3285,N_3905);
nor U7721 (N_7721,N_197,N_1254);
or U7722 (N_7722,N_4663,N_690);
or U7723 (N_7723,N_4063,N_4332);
and U7724 (N_7724,N_446,N_750);
nand U7725 (N_7725,N_519,N_3588);
and U7726 (N_7726,N_4510,N_243);
nand U7727 (N_7727,N_1480,N_4025);
nor U7728 (N_7728,N_3710,N_1708);
nand U7729 (N_7729,N_4547,N_4274);
and U7730 (N_7730,N_2259,N_4058);
or U7731 (N_7731,N_1518,N_2656);
xor U7732 (N_7732,N_989,N_21);
xor U7733 (N_7733,N_2762,N_635);
xor U7734 (N_7734,N_3293,N_223);
nand U7735 (N_7735,N_2255,N_1059);
nand U7736 (N_7736,N_4367,N_3086);
or U7737 (N_7737,N_894,N_3393);
xnor U7738 (N_7738,N_3681,N_3989);
or U7739 (N_7739,N_1574,N_2288);
and U7740 (N_7740,N_3867,N_4601);
and U7741 (N_7741,N_3334,N_1372);
and U7742 (N_7742,N_1791,N_4600);
and U7743 (N_7743,N_3129,N_1372);
or U7744 (N_7744,N_264,N_4249);
and U7745 (N_7745,N_3077,N_3184);
or U7746 (N_7746,N_4993,N_1266);
and U7747 (N_7747,N_4683,N_3399);
nor U7748 (N_7748,N_2107,N_2660);
nor U7749 (N_7749,N_3223,N_1083);
nand U7750 (N_7750,N_3503,N_766);
xnor U7751 (N_7751,N_4815,N_2723);
and U7752 (N_7752,N_3750,N_2359);
nor U7753 (N_7753,N_3119,N_184);
nor U7754 (N_7754,N_3485,N_2529);
or U7755 (N_7755,N_1888,N_1349);
xnor U7756 (N_7756,N_263,N_25);
and U7757 (N_7757,N_1329,N_343);
or U7758 (N_7758,N_722,N_469);
nor U7759 (N_7759,N_380,N_4066);
or U7760 (N_7760,N_1580,N_1694);
nand U7761 (N_7761,N_4015,N_732);
or U7762 (N_7762,N_81,N_50);
nor U7763 (N_7763,N_4954,N_2479);
and U7764 (N_7764,N_200,N_1195);
or U7765 (N_7765,N_4719,N_1198);
xor U7766 (N_7766,N_310,N_4090);
and U7767 (N_7767,N_2676,N_2132);
nand U7768 (N_7768,N_2440,N_451);
or U7769 (N_7769,N_4317,N_3870);
nor U7770 (N_7770,N_4474,N_1093);
nor U7771 (N_7771,N_3789,N_1867);
nor U7772 (N_7772,N_842,N_3927);
nand U7773 (N_7773,N_4405,N_1518);
nand U7774 (N_7774,N_410,N_1355);
nor U7775 (N_7775,N_291,N_3026);
and U7776 (N_7776,N_4447,N_1232);
nor U7777 (N_7777,N_4898,N_2698);
or U7778 (N_7778,N_2764,N_885);
or U7779 (N_7779,N_51,N_2647);
nand U7780 (N_7780,N_1529,N_2683);
and U7781 (N_7781,N_4636,N_2451);
and U7782 (N_7782,N_3404,N_1153);
nand U7783 (N_7783,N_1624,N_4869);
nand U7784 (N_7784,N_562,N_2792);
and U7785 (N_7785,N_495,N_2355);
or U7786 (N_7786,N_4536,N_3606);
nor U7787 (N_7787,N_565,N_2733);
nor U7788 (N_7788,N_4644,N_2700);
xnor U7789 (N_7789,N_783,N_2751);
or U7790 (N_7790,N_4877,N_2148);
nor U7791 (N_7791,N_1406,N_1694);
xor U7792 (N_7792,N_2599,N_3480);
nand U7793 (N_7793,N_1868,N_4067);
nand U7794 (N_7794,N_4572,N_388);
and U7795 (N_7795,N_2573,N_2301);
xor U7796 (N_7796,N_2705,N_479);
or U7797 (N_7797,N_301,N_1427);
and U7798 (N_7798,N_1124,N_3012);
nor U7799 (N_7799,N_3625,N_2653);
nand U7800 (N_7800,N_866,N_3794);
or U7801 (N_7801,N_4665,N_3218);
and U7802 (N_7802,N_4357,N_28);
and U7803 (N_7803,N_4130,N_331);
or U7804 (N_7804,N_3322,N_2588);
and U7805 (N_7805,N_4050,N_2787);
and U7806 (N_7806,N_57,N_116);
nor U7807 (N_7807,N_3766,N_3160);
nand U7808 (N_7808,N_4262,N_4208);
nand U7809 (N_7809,N_2391,N_2164);
nand U7810 (N_7810,N_4799,N_1761);
nand U7811 (N_7811,N_3609,N_965);
nand U7812 (N_7812,N_2284,N_3280);
or U7813 (N_7813,N_2621,N_777);
nand U7814 (N_7814,N_4955,N_1207);
nor U7815 (N_7815,N_4396,N_2421);
and U7816 (N_7816,N_788,N_463);
nor U7817 (N_7817,N_2463,N_658);
nor U7818 (N_7818,N_374,N_1476);
or U7819 (N_7819,N_211,N_1311);
nor U7820 (N_7820,N_378,N_494);
or U7821 (N_7821,N_2441,N_4086);
or U7822 (N_7822,N_2095,N_3093);
or U7823 (N_7823,N_1911,N_4359);
and U7824 (N_7824,N_3485,N_3949);
nor U7825 (N_7825,N_1591,N_4645);
or U7826 (N_7826,N_815,N_4539);
nand U7827 (N_7827,N_2086,N_2452);
and U7828 (N_7828,N_4108,N_2263);
or U7829 (N_7829,N_3201,N_1660);
nor U7830 (N_7830,N_4420,N_1186);
xnor U7831 (N_7831,N_4907,N_2411);
or U7832 (N_7832,N_2718,N_709);
xor U7833 (N_7833,N_2807,N_710);
or U7834 (N_7834,N_1626,N_1785);
xor U7835 (N_7835,N_1150,N_804);
nand U7836 (N_7836,N_1474,N_1166);
nor U7837 (N_7837,N_4027,N_4172);
nor U7838 (N_7838,N_4033,N_3521);
or U7839 (N_7839,N_3461,N_942);
nor U7840 (N_7840,N_4040,N_1531);
and U7841 (N_7841,N_4484,N_2551);
or U7842 (N_7842,N_998,N_1728);
or U7843 (N_7843,N_3845,N_574);
nand U7844 (N_7844,N_811,N_4322);
and U7845 (N_7845,N_3352,N_248);
nor U7846 (N_7846,N_3724,N_4240);
and U7847 (N_7847,N_2750,N_1673);
and U7848 (N_7848,N_4405,N_3855);
nand U7849 (N_7849,N_2533,N_2660);
nor U7850 (N_7850,N_1187,N_1956);
or U7851 (N_7851,N_4184,N_1668);
or U7852 (N_7852,N_979,N_1041);
or U7853 (N_7853,N_4852,N_417);
and U7854 (N_7854,N_4876,N_1663);
and U7855 (N_7855,N_3182,N_1009);
nand U7856 (N_7856,N_3365,N_1851);
and U7857 (N_7857,N_2124,N_1266);
xnor U7858 (N_7858,N_1283,N_207);
and U7859 (N_7859,N_1344,N_3200);
and U7860 (N_7860,N_4578,N_839);
xnor U7861 (N_7861,N_1045,N_1629);
or U7862 (N_7862,N_3477,N_3601);
or U7863 (N_7863,N_2639,N_1800);
nand U7864 (N_7864,N_3859,N_2761);
nor U7865 (N_7865,N_3179,N_409);
xor U7866 (N_7866,N_1380,N_1903);
and U7867 (N_7867,N_4322,N_1130);
nand U7868 (N_7868,N_2936,N_1089);
or U7869 (N_7869,N_3528,N_539);
nor U7870 (N_7870,N_231,N_485);
nand U7871 (N_7871,N_884,N_2475);
or U7872 (N_7872,N_2892,N_4123);
or U7873 (N_7873,N_3350,N_2383);
or U7874 (N_7874,N_2402,N_4536);
nand U7875 (N_7875,N_3633,N_3079);
or U7876 (N_7876,N_3661,N_1808);
nand U7877 (N_7877,N_36,N_2518);
nor U7878 (N_7878,N_2234,N_948);
and U7879 (N_7879,N_2904,N_1465);
nand U7880 (N_7880,N_1754,N_3613);
nor U7881 (N_7881,N_4680,N_3938);
or U7882 (N_7882,N_1037,N_2505);
or U7883 (N_7883,N_4567,N_4718);
and U7884 (N_7884,N_4369,N_4298);
nor U7885 (N_7885,N_4660,N_3491);
and U7886 (N_7886,N_2424,N_2481);
nor U7887 (N_7887,N_3712,N_3309);
and U7888 (N_7888,N_479,N_1802);
nand U7889 (N_7889,N_4197,N_4243);
xnor U7890 (N_7890,N_2840,N_845);
and U7891 (N_7891,N_2611,N_1220);
or U7892 (N_7892,N_3743,N_806);
and U7893 (N_7893,N_3935,N_3539);
nor U7894 (N_7894,N_42,N_2143);
and U7895 (N_7895,N_4354,N_2251);
and U7896 (N_7896,N_858,N_912);
nand U7897 (N_7897,N_924,N_4258);
or U7898 (N_7898,N_2837,N_1736);
and U7899 (N_7899,N_4,N_4730);
nand U7900 (N_7900,N_4885,N_1797);
nor U7901 (N_7901,N_4556,N_4920);
nand U7902 (N_7902,N_3585,N_1215);
nor U7903 (N_7903,N_3886,N_4488);
or U7904 (N_7904,N_2959,N_2524);
and U7905 (N_7905,N_1027,N_3567);
or U7906 (N_7906,N_1346,N_3633);
nor U7907 (N_7907,N_4634,N_456);
nand U7908 (N_7908,N_3650,N_2030);
or U7909 (N_7909,N_2793,N_3426);
nor U7910 (N_7910,N_2820,N_3382);
and U7911 (N_7911,N_3382,N_3529);
or U7912 (N_7912,N_2286,N_4018);
xnor U7913 (N_7913,N_1763,N_4769);
or U7914 (N_7914,N_1381,N_2052);
nand U7915 (N_7915,N_3764,N_2388);
and U7916 (N_7916,N_1673,N_3263);
and U7917 (N_7917,N_4207,N_77);
and U7918 (N_7918,N_2788,N_2108);
nor U7919 (N_7919,N_4692,N_3900);
and U7920 (N_7920,N_1374,N_4635);
and U7921 (N_7921,N_1172,N_3697);
nor U7922 (N_7922,N_2235,N_2137);
or U7923 (N_7923,N_3523,N_3366);
and U7924 (N_7924,N_4573,N_3522);
and U7925 (N_7925,N_158,N_4366);
and U7926 (N_7926,N_4403,N_2631);
nor U7927 (N_7927,N_2990,N_1470);
or U7928 (N_7928,N_452,N_987);
nor U7929 (N_7929,N_4564,N_4021);
nand U7930 (N_7930,N_2599,N_1307);
nand U7931 (N_7931,N_1150,N_2283);
nor U7932 (N_7932,N_1014,N_605);
nor U7933 (N_7933,N_3133,N_3007);
nand U7934 (N_7934,N_3249,N_2844);
xnor U7935 (N_7935,N_2926,N_1197);
nand U7936 (N_7936,N_179,N_3730);
or U7937 (N_7937,N_662,N_3028);
and U7938 (N_7938,N_3299,N_2638);
nor U7939 (N_7939,N_4352,N_788);
nor U7940 (N_7940,N_3234,N_3556);
or U7941 (N_7941,N_1707,N_4680);
xor U7942 (N_7942,N_2130,N_1699);
and U7943 (N_7943,N_3372,N_4281);
nor U7944 (N_7944,N_218,N_1322);
and U7945 (N_7945,N_3209,N_1183);
nor U7946 (N_7946,N_1735,N_2632);
nor U7947 (N_7947,N_3242,N_3440);
and U7948 (N_7948,N_226,N_2111);
and U7949 (N_7949,N_2512,N_2688);
nand U7950 (N_7950,N_899,N_1991);
nor U7951 (N_7951,N_2122,N_3962);
and U7952 (N_7952,N_4357,N_267);
nand U7953 (N_7953,N_3886,N_4066);
and U7954 (N_7954,N_736,N_4385);
and U7955 (N_7955,N_2290,N_4458);
nand U7956 (N_7956,N_3885,N_1123);
nor U7957 (N_7957,N_3978,N_4296);
or U7958 (N_7958,N_872,N_3854);
xor U7959 (N_7959,N_1258,N_4244);
nor U7960 (N_7960,N_1223,N_1088);
nand U7961 (N_7961,N_4259,N_4612);
or U7962 (N_7962,N_4751,N_2868);
and U7963 (N_7963,N_4734,N_3544);
and U7964 (N_7964,N_4304,N_1993);
nor U7965 (N_7965,N_3229,N_4672);
or U7966 (N_7966,N_4560,N_4014);
or U7967 (N_7967,N_4610,N_2885);
xor U7968 (N_7968,N_731,N_1209);
and U7969 (N_7969,N_3174,N_1412);
nand U7970 (N_7970,N_2684,N_3643);
or U7971 (N_7971,N_523,N_2957);
and U7972 (N_7972,N_1031,N_749);
or U7973 (N_7973,N_4267,N_1437);
nor U7974 (N_7974,N_3025,N_2264);
or U7975 (N_7975,N_3194,N_1190);
xor U7976 (N_7976,N_3988,N_4113);
and U7977 (N_7977,N_296,N_2870);
nor U7978 (N_7978,N_2690,N_2166);
or U7979 (N_7979,N_3065,N_580);
nor U7980 (N_7980,N_2188,N_2398);
or U7981 (N_7981,N_1343,N_2788);
and U7982 (N_7982,N_1425,N_4272);
or U7983 (N_7983,N_726,N_2047);
or U7984 (N_7984,N_2656,N_4541);
xnor U7985 (N_7985,N_3176,N_1500);
or U7986 (N_7986,N_3303,N_2118);
and U7987 (N_7987,N_1151,N_3894);
and U7988 (N_7988,N_243,N_1485);
nand U7989 (N_7989,N_1838,N_4646);
or U7990 (N_7990,N_1476,N_1100);
nor U7991 (N_7991,N_1298,N_3098);
nor U7992 (N_7992,N_366,N_1387);
nor U7993 (N_7993,N_3214,N_4108);
and U7994 (N_7994,N_4328,N_4704);
nor U7995 (N_7995,N_4722,N_941);
nand U7996 (N_7996,N_1956,N_523);
and U7997 (N_7997,N_4554,N_1778);
nor U7998 (N_7998,N_2581,N_2070);
and U7999 (N_7999,N_3768,N_1446);
nand U8000 (N_8000,N_173,N_2841);
and U8001 (N_8001,N_1671,N_2891);
nor U8002 (N_8002,N_793,N_3545);
nand U8003 (N_8003,N_4639,N_790);
and U8004 (N_8004,N_1252,N_3088);
nor U8005 (N_8005,N_296,N_1337);
or U8006 (N_8006,N_3509,N_2258);
nor U8007 (N_8007,N_984,N_2019);
or U8008 (N_8008,N_3526,N_1273);
nor U8009 (N_8009,N_3649,N_2423);
nand U8010 (N_8010,N_4093,N_187);
nor U8011 (N_8011,N_2774,N_2010);
xor U8012 (N_8012,N_4045,N_4816);
and U8013 (N_8013,N_1767,N_4313);
or U8014 (N_8014,N_4499,N_961);
nor U8015 (N_8015,N_1778,N_2853);
or U8016 (N_8016,N_655,N_932);
nor U8017 (N_8017,N_3950,N_4927);
xnor U8018 (N_8018,N_2555,N_3867);
and U8019 (N_8019,N_4261,N_3513);
nand U8020 (N_8020,N_1656,N_2401);
nor U8021 (N_8021,N_1805,N_1459);
and U8022 (N_8022,N_341,N_1582);
and U8023 (N_8023,N_46,N_2103);
and U8024 (N_8024,N_1319,N_1188);
or U8025 (N_8025,N_4509,N_3075);
nand U8026 (N_8026,N_4651,N_3096);
or U8027 (N_8027,N_3999,N_3362);
nor U8028 (N_8028,N_685,N_998);
or U8029 (N_8029,N_2240,N_4116);
nor U8030 (N_8030,N_1117,N_557);
or U8031 (N_8031,N_4652,N_623);
or U8032 (N_8032,N_1871,N_3739);
nand U8033 (N_8033,N_1589,N_770);
and U8034 (N_8034,N_2363,N_3740);
nand U8035 (N_8035,N_4884,N_3580);
or U8036 (N_8036,N_2431,N_3467);
and U8037 (N_8037,N_3839,N_4808);
nand U8038 (N_8038,N_2442,N_4765);
or U8039 (N_8039,N_4348,N_337);
nand U8040 (N_8040,N_837,N_2426);
nand U8041 (N_8041,N_3726,N_458);
or U8042 (N_8042,N_1922,N_2839);
nand U8043 (N_8043,N_308,N_2711);
and U8044 (N_8044,N_890,N_2692);
xnor U8045 (N_8045,N_1920,N_1381);
or U8046 (N_8046,N_4091,N_2191);
and U8047 (N_8047,N_3662,N_2482);
nor U8048 (N_8048,N_1121,N_3575);
and U8049 (N_8049,N_4959,N_4845);
and U8050 (N_8050,N_868,N_2913);
and U8051 (N_8051,N_451,N_3570);
xor U8052 (N_8052,N_4217,N_933);
and U8053 (N_8053,N_862,N_4929);
nand U8054 (N_8054,N_216,N_3403);
nor U8055 (N_8055,N_3367,N_4113);
or U8056 (N_8056,N_4882,N_3581);
nor U8057 (N_8057,N_2196,N_4148);
nand U8058 (N_8058,N_164,N_447);
xnor U8059 (N_8059,N_3415,N_3318);
and U8060 (N_8060,N_105,N_4934);
or U8061 (N_8061,N_3999,N_521);
and U8062 (N_8062,N_1546,N_2178);
or U8063 (N_8063,N_4777,N_2107);
nor U8064 (N_8064,N_802,N_3796);
nor U8065 (N_8065,N_3386,N_4910);
nand U8066 (N_8066,N_4031,N_4987);
nand U8067 (N_8067,N_1001,N_1891);
or U8068 (N_8068,N_4126,N_2401);
nor U8069 (N_8069,N_3838,N_2669);
nand U8070 (N_8070,N_763,N_283);
or U8071 (N_8071,N_2813,N_3788);
and U8072 (N_8072,N_2690,N_936);
xnor U8073 (N_8073,N_1079,N_3434);
nor U8074 (N_8074,N_629,N_3335);
nor U8075 (N_8075,N_2583,N_396);
nor U8076 (N_8076,N_4731,N_2504);
or U8077 (N_8077,N_64,N_3648);
and U8078 (N_8078,N_1253,N_4050);
nor U8079 (N_8079,N_4098,N_4988);
or U8080 (N_8080,N_682,N_816);
or U8081 (N_8081,N_4209,N_4279);
nand U8082 (N_8082,N_83,N_1306);
xor U8083 (N_8083,N_1129,N_1279);
nor U8084 (N_8084,N_3040,N_4838);
nor U8085 (N_8085,N_3915,N_4281);
nand U8086 (N_8086,N_4171,N_3206);
xor U8087 (N_8087,N_3210,N_3213);
nor U8088 (N_8088,N_3503,N_2456);
and U8089 (N_8089,N_4954,N_2522);
nand U8090 (N_8090,N_4473,N_3045);
or U8091 (N_8091,N_4576,N_4769);
and U8092 (N_8092,N_510,N_2294);
or U8093 (N_8093,N_239,N_89);
nand U8094 (N_8094,N_2017,N_1084);
or U8095 (N_8095,N_3209,N_2281);
or U8096 (N_8096,N_1821,N_3593);
or U8097 (N_8097,N_331,N_3208);
nor U8098 (N_8098,N_1557,N_1586);
nor U8099 (N_8099,N_1195,N_262);
nor U8100 (N_8100,N_623,N_737);
or U8101 (N_8101,N_3356,N_2813);
xor U8102 (N_8102,N_3545,N_3544);
nand U8103 (N_8103,N_3183,N_1964);
nor U8104 (N_8104,N_4290,N_532);
or U8105 (N_8105,N_2490,N_4011);
xnor U8106 (N_8106,N_2760,N_1768);
or U8107 (N_8107,N_1422,N_783);
or U8108 (N_8108,N_1156,N_4138);
nand U8109 (N_8109,N_1069,N_1402);
nor U8110 (N_8110,N_1827,N_686);
or U8111 (N_8111,N_721,N_105);
nor U8112 (N_8112,N_756,N_1550);
and U8113 (N_8113,N_2490,N_1197);
nor U8114 (N_8114,N_2087,N_4256);
xnor U8115 (N_8115,N_2016,N_4524);
nand U8116 (N_8116,N_3833,N_1236);
or U8117 (N_8117,N_764,N_2114);
nor U8118 (N_8118,N_2099,N_80);
nor U8119 (N_8119,N_4737,N_1019);
or U8120 (N_8120,N_2113,N_4341);
or U8121 (N_8121,N_3113,N_263);
nand U8122 (N_8122,N_2609,N_136);
nor U8123 (N_8123,N_471,N_4815);
nand U8124 (N_8124,N_1882,N_1707);
and U8125 (N_8125,N_2809,N_3281);
nor U8126 (N_8126,N_1420,N_2200);
nand U8127 (N_8127,N_1356,N_1550);
xnor U8128 (N_8128,N_4443,N_1355);
xor U8129 (N_8129,N_267,N_1753);
or U8130 (N_8130,N_3378,N_3830);
nand U8131 (N_8131,N_4971,N_1543);
and U8132 (N_8132,N_4465,N_193);
and U8133 (N_8133,N_4771,N_3995);
nand U8134 (N_8134,N_4916,N_3943);
or U8135 (N_8135,N_1253,N_4837);
nand U8136 (N_8136,N_824,N_3826);
nor U8137 (N_8137,N_4422,N_569);
and U8138 (N_8138,N_1482,N_4978);
nand U8139 (N_8139,N_1121,N_4484);
nand U8140 (N_8140,N_2747,N_3765);
or U8141 (N_8141,N_1246,N_567);
nand U8142 (N_8142,N_1810,N_802);
and U8143 (N_8143,N_558,N_1649);
nand U8144 (N_8144,N_3487,N_3889);
nand U8145 (N_8145,N_1130,N_2010);
or U8146 (N_8146,N_91,N_875);
or U8147 (N_8147,N_1260,N_1625);
nand U8148 (N_8148,N_4429,N_424);
or U8149 (N_8149,N_4253,N_2428);
or U8150 (N_8150,N_976,N_3437);
and U8151 (N_8151,N_1288,N_4752);
nand U8152 (N_8152,N_4652,N_4273);
nand U8153 (N_8153,N_2899,N_1006);
nor U8154 (N_8154,N_1060,N_131);
and U8155 (N_8155,N_2439,N_3269);
and U8156 (N_8156,N_1838,N_4778);
nand U8157 (N_8157,N_3186,N_207);
or U8158 (N_8158,N_2458,N_2385);
nand U8159 (N_8159,N_1572,N_1588);
xnor U8160 (N_8160,N_1041,N_3798);
xnor U8161 (N_8161,N_3459,N_4901);
and U8162 (N_8162,N_741,N_2451);
nor U8163 (N_8163,N_2288,N_2262);
xnor U8164 (N_8164,N_269,N_2118);
nand U8165 (N_8165,N_1262,N_928);
and U8166 (N_8166,N_3426,N_4333);
xnor U8167 (N_8167,N_4919,N_90);
and U8168 (N_8168,N_3314,N_2697);
nor U8169 (N_8169,N_1756,N_1069);
or U8170 (N_8170,N_4840,N_3180);
or U8171 (N_8171,N_249,N_4244);
nand U8172 (N_8172,N_852,N_1250);
or U8173 (N_8173,N_2528,N_2275);
nor U8174 (N_8174,N_3022,N_4937);
and U8175 (N_8175,N_3384,N_2252);
nor U8176 (N_8176,N_1066,N_1355);
nor U8177 (N_8177,N_596,N_1417);
and U8178 (N_8178,N_3828,N_2030);
and U8179 (N_8179,N_2052,N_1834);
nand U8180 (N_8180,N_1142,N_3866);
xnor U8181 (N_8181,N_893,N_3079);
nor U8182 (N_8182,N_713,N_1167);
xor U8183 (N_8183,N_3167,N_48);
nand U8184 (N_8184,N_2322,N_4821);
and U8185 (N_8185,N_4792,N_364);
or U8186 (N_8186,N_4031,N_3444);
and U8187 (N_8187,N_1522,N_2883);
or U8188 (N_8188,N_2136,N_4645);
and U8189 (N_8189,N_162,N_4532);
or U8190 (N_8190,N_4273,N_3068);
or U8191 (N_8191,N_4315,N_3870);
or U8192 (N_8192,N_2746,N_3201);
or U8193 (N_8193,N_2221,N_1699);
xor U8194 (N_8194,N_4815,N_1121);
or U8195 (N_8195,N_3234,N_3630);
and U8196 (N_8196,N_4795,N_640);
nand U8197 (N_8197,N_1836,N_3248);
xnor U8198 (N_8198,N_4776,N_1853);
or U8199 (N_8199,N_13,N_2668);
nor U8200 (N_8200,N_2026,N_4950);
nor U8201 (N_8201,N_2845,N_1396);
nand U8202 (N_8202,N_4682,N_311);
or U8203 (N_8203,N_4501,N_2226);
and U8204 (N_8204,N_57,N_321);
xor U8205 (N_8205,N_807,N_3749);
or U8206 (N_8206,N_1951,N_4583);
nand U8207 (N_8207,N_834,N_3619);
nor U8208 (N_8208,N_4118,N_4830);
nor U8209 (N_8209,N_3005,N_1781);
nor U8210 (N_8210,N_4697,N_457);
xor U8211 (N_8211,N_303,N_4411);
or U8212 (N_8212,N_2052,N_1748);
and U8213 (N_8213,N_4026,N_2176);
or U8214 (N_8214,N_2821,N_3117);
or U8215 (N_8215,N_3586,N_2687);
nand U8216 (N_8216,N_1865,N_2885);
nor U8217 (N_8217,N_1300,N_4098);
nor U8218 (N_8218,N_2094,N_1665);
nor U8219 (N_8219,N_1436,N_2092);
nand U8220 (N_8220,N_2011,N_3934);
nand U8221 (N_8221,N_4444,N_2317);
and U8222 (N_8222,N_4515,N_927);
or U8223 (N_8223,N_843,N_3218);
and U8224 (N_8224,N_967,N_2870);
nand U8225 (N_8225,N_683,N_1736);
and U8226 (N_8226,N_2560,N_4835);
and U8227 (N_8227,N_198,N_4988);
nor U8228 (N_8228,N_4712,N_3609);
or U8229 (N_8229,N_4707,N_3145);
or U8230 (N_8230,N_1011,N_995);
and U8231 (N_8231,N_4923,N_1966);
or U8232 (N_8232,N_1587,N_699);
or U8233 (N_8233,N_595,N_3487);
nor U8234 (N_8234,N_1867,N_1866);
and U8235 (N_8235,N_1198,N_1451);
nor U8236 (N_8236,N_2394,N_3972);
nor U8237 (N_8237,N_506,N_1756);
nand U8238 (N_8238,N_1535,N_4216);
nor U8239 (N_8239,N_3165,N_1374);
and U8240 (N_8240,N_4449,N_473);
nor U8241 (N_8241,N_936,N_4309);
nand U8242 (N_8242,N_1280,N_770);
xnor U8243 (N_8243,N_767,N_4388);
nand U8244 (N_8244,N_1583,N_3901);
nor U8245 (N_8245,N_3871,N_471);
nor U8246 (N_8246,N_4803,N_3640);
nor U8247 (N_8247,N_4779,N_2115);
nand U8248 (N_8248,N_2578,N_1121);
xor U8249 (N_8249,N_1839,N_2284);
nor U8250 (N_8250,N_895,N_1960);
nand U8251 (N_8251,N_1205,N_130);
or U8252 (N_8252,N_1463,N_3281);
and U8253 (N_8253,N_979,N_725);
xor U8254 (N_8254,N_4804,N_4507);
or U8255 (N_8255,N_3777,N_2620);
or U8256 (N_8256,N_1168,N_2160);
nor U8257 (N_8257,N_4541,N_1018);
nor U8258 (N_8258,N_4560,N_606);
nor U8259 (N_8259,N_245,N_4470);
nand U8260 (N_8260,N_4448,N_334);
nand U8261 (N_8261,N_3909,N_1917);
nand U8262 (N_8262,N_568,N_3941);
xnor U8263 (N_8263,N_4839,N_3153);
nand U8264 (N_8264,N_2771,N_969);
nor U8265 (N_8265,N_2768,N_2993);
or U8266 (N_8266,N_4433,N_766);
nor U8267 (N_8267,N_427,N_3628);
nor U8268 (N_8268,N_4151,N_2067);
and U8269 (N_8269,N_403,N_192);
nand U8270 (N_8270,N_2412,N_1599);
nor U8271 (N_8271,N_821,N_4066);
xor U8272 (N_8272,N_1963,N_3046);
nor U8273 (N_8273,N_2136,N_8);
nor U8274 (N_8274,N_4249,N_4520);
nand U8275 (N_8275,N_57,N_474);
and U8276 (N_8276,N_1547,N_165);
nor U8277 (N_8277,N_4928,N_2703);
nand U8278 (N_8278,N_784,N_1013);
nand U8279 (N_8279,N_1342,N_4949);
nor U8280 (N_8280,N_505,N_2356);
xnor U8281 (N_8281,N_435,N_4184);
xnor U8282 (N_8282,N_1223,N_1413);
and U8283 (N_8283,N_4700,N_3327);
and U8284 (N_8284,N_4350,N_1900);
nand U8285 (N_8285,N_2584,N_1186);
nand U8286 (N_8286,N_2743,N_3337);
nand U8287 (N_8287,N_3126,N_55);
xnor U8288 (N_8288,N_876,N_1943);
and U8289 (N_8289,N_1093,N_109);
xor U8290 (N_8290,N_3961,N_1019);
and U8291 (N_8291,N_425,N_132);
or U8292 (N_8292,N_3808,N_20);
nand U8293 (N_8293,N_1767,N_2226);
or U8294 (N_8294,N_3900,N_2050);
and U8295 (N_8295,N_4140,N_3163);
nand U8296 (N_8296,N_3900,N_566);
or U8297 (N_8297,N_1655,N_1523);
and U8298 (N_8298,N_3193,N_13);
nor U8299 (N_8299,N_60,N_151);
nor U8300 (N_8300,N_3198,N_4541);
or U8301 (N_8301,N_883,N_4126);
nor U8302 (N_8302,N_3516,N_2741);
nand U8303 (N_8303,N_3585,N_2301);
and U8304 (N_8304,N_824,N_4144);
and U8305 (N_8305,N_2543,N_3910);
xnor U8306 (N_8306,N_4476,N_1261);
nand U8307 (N_8307,N_3115,N_1331);
xnor U8308 (N_8308,N_2593,N_4538);
nand U8309 (N_8309,N_4439,N_3069);
nand U8310 (N_8310,N_1678,N_2081);
nor U8311 (N_8311,N_4711,N_1492);
or U8312 (N_8312,N_1012,N_716);
nor U8313 (N_8313,N_259,N_1557);
nand U8314 (N_8314,N_3629,N_1614);
nand U8315 (N_8315,N_2413,N_3256);
or U8316 (N_8316,N_3281,N_4963);
nand U8317 (N_8317,N_209,N_385);
or U8318 (N_8318,N_513,N_198);
nand U8319 (N_8319,N_1115,N_4394);
and U8320 (N_8320,N_807,N_2321);
nand U8321 (N_8321,N_3247,N_2411);
nor U8322 (N_8322,N_1834,N_1574);
nand U8323 (N_8323,N_3566,N_874);
xnor U8324 (N_8324,N_1765,N_1514);
xnor U8325 (N_8325,N_929,N_2548);
or U8326 (N_8326,N_1162,N_1134);
and U8327 (N_8327,N_2693,N_1655);
or U8328 (N_8328,N_176,N_1199);
or U8329 (N_8329,N_3632,N_1800);
xnor U8330 (N_8330,N_2583,N_4294);
nor U8331 (N_8331,N_845,N_2929);
nor U8332 (N_8332,N_2513,N_3305);
nor U8333 (N_8333,N_3538,N_3742);
nor U8334 (N_8334,N_4505,N_3497);
and U8335 (N_8335,N_704,N_4200);
and U8336 (N_8336,N_1892,N_3280);
and U8337 (N_8337,N_4293,N_2095);
or U8338 (N_8338,N_1459,N_3627);
nor U8339 (N_8339,N_2035,N_4308);
nor U8340 (N_8340,N_3451,N_4991);
nand U8341 (N_8341,N_3915,N_1763);
and U8342 (N_8342,N_2380,N_489);
xor U8343 (N_8343,N_4852,N_2414);
nand U8344 (N_8344,N_2232,N_4892);
nand U8345 (N_8345,N_312,N_1967);
xor U8346 (N_8346,N_737,N_781);
nand U8347 (N_8347,N_3023,N_856);
nor U8348 (N_8348,N_2422,N_4767);
or U8349 (N_8349,N_2652,N_2634);
and U8350 (N_8350,N_2982,N_2008);
nor U8351 (N_8351,N_1932,N_4817);
nor U8352 (N_8352,N_4846,N_940);
and U8353 (N_8353,N_4313,N_352);
or U8354 (N_8354,N_162,N_476);
or U8355 (N_8355,N_1917,N_1807);
nand U8356 (N_8356,N_3443,N_351);
nand U8357 (N_8357,N_169,N_3341);
or U8358 (N_8358,N_3957,N_4621);
nor U8359 (N_8359,N_1584,N_4330);
or U8360 (N_8360,N_4534,N_4266);
or U8361 (N_8361,N_1649,N_1595);
or U8362 (N_8362,N_2874,N_3496);
nor U8363 (N_8363,N_1958,N_588);
and U8364 (N_8364,N_1150,N_4698);
or U8365 (N_8365,N_2307,N_2853);
xnor U8366 (N_8366,N_134,N_1615);
and U8367 (N_8367,N_1188,N_1770);
or U8368 (N_8368,N_4289,N_302);
and U8369 (N_8369,N_3984,N_1154);
nand U8370 (N_8370,N_951,N_3910);
or U8371 (N_8371,N_4405,N_3771);
nor U8372 (N_8372,N_3525,N_2841);
nand U8373 (N_8373,N_2296,N_3540);
nor U8374 (N_8374,N_2184,N_2005);
and U8375 (N_8375,N_799,N_4036);
xnor U8376 (N_8376,N_207,N_3828);
and U8377 (N_8377,N_4547,N_2842);
or U8378 (N_8378,N_4117,N_4979);
nand U8379 (N_8379,N_1075,N_3166);
nand U8380 (N_8380,N_3764,N_4465);
nor U8381 (N_8381,N_731,N_1023);
and U8382 (N_8382,N_4749,N_2166);
or U8383 (N_8383,N_1974,N_543);
or U8384 (N_8384,N_1460,N_3980);
or U8385 (N_8385,N_2322,N_3041);
or U8386 (N_8386,N_3624,N_3705);
nor U8387 (N_8387,N_4401,N_396);
nand U8388 (N_8388,N_679,N_2738);
nor U8389 (N_8389,N_1110,N_4271);
nand U8390 (N_8390,N_2751,N_124);
xnor U8391 (N_8391,N_4618,N_3287);
or U8392 (N_8392,N_661,N_4803);
nor U8393 (N_8393,N_1405,N_1734);
nor U8394 (N_8394,N_4927,N_1534);
nor U8395 (N_8395,N_2787,N_4075);
nor U8396 (N_8396,N_1020,N_3100);
or U8397 (N_8397,N_2099,N_1201);
nor U8398 (N_8398,N_3222,N_2526);
and U8399 (N_8399,N_4615,N_4511);
or U8400 (N_8400,N_1500,N_2179);
xor U8401 (N_8401,N_263,N_2355);
and U8402 (N_8402,N_4392,N_3105);
or U8403 (N_8403,N_1709,N_3443);
nor U8404 (N_8404,N_3364,N_622);
or U8405 (N_8405,N_3133,N_4123);
or U8406 (N_8406,N_1887,N_4455);
nor U8407 (N_8407,N_4943,N_589);
nor U8408 (N_8408,N_4617,N_1030);
or U8409 (N_8409,N_4680,N_1055);
or U8410 (N_8410,N_4901,N_630);
nand U8411 (N_8411,N_3028,N_4670);
nand U8412 (N_8412,N_1187,N_4682);
or U8413 (N_8413,N_3194,N_3920);
nor U8414 (N_8414,N_2464,N_4137);
nand U8415 (N_8415,N_4450,N_1570);
nand U8416 (N_8416,N_3932,N_2271);
nand U8417 (N_8417,N_4333,N_3814);
nor U8418 (N_8418,N_2769,N_1658);
xor U8419 (N_8419,N_311,N_2016);
xor U8420 (N_8420,N_3065,N_2269);
and U8421 (N_8421,N_2199,N_4379);
nor U8422 (N_8422,N_290,N_2281);
and U8423 (N_8423,N_4893,N_3990);
nor U8424 (N_8424,N_1566,N_1552);
xnor U8425 (N_8425,N_3943,N_4434);
and U8426 (N_8426,N_946,N_4075);
nor U8427 (N_8427,N_1779,N_1775);
xnor U8428 (N_8428,N_3551,N_2142);
or U8429 (N_8429,N_4430,N_1350);
nand U8430 (N_8430,N_3046,N_3374);
nor U8431 (N_8431,N_4852,N_2348);
or U8432 (N_8432,N_4971,N_1207);
or U8433 (N_8433,N_2182,N_529);
nor U8434 (N_8434,N_1323,N_1259);
nor U8435 (N_8435,N_4271,N_3394);
and U8436 (N_8436,N_4010,N_3860);
nand U8437 (N_8437,N_2035,N_2503);
and U8438 (N_8438,N_161,N_2146);
and U8439 (N_8439,N_980,N_3465);
and U8440 (N_8440,N_1510,N_2453);
nor U8441 (N_8441,N_616,N_3927);
or U8442 (N_8442,N_3684,N_4476);
or U8443 (N_8443,N_1261,N_1727);
nand U8444 (N_8444,N_2324,N_3403);
nand U8445 (N_8445,N_4777,N_508);
and U8446 (N_8446,N_4012,N_2463);
nand U8447 (N_8447,N_2902,N_4187);
or U8448 (N_8448,N_4409,N_842);
xor U8449 (N_8449,N_3562,N_4103);
and U8450 (N_8450,N_3894,N_2691);
nor U8451 (N_8451,N_518,N_9);
nand U8452 (N_8452,N_3290,N_3075);
xor U8453 (N_8453,N_4164,N_2044);
nand U8454 (N_8454,N_2901,N_4503);
or U8455 (N_8455,N_3906,N_2673);
nand U8456 (N_8456,N_963,N_892);
nand U8457 (N_8457,N_4452,N_1055);
nand U8458 (N_8458,N_136,N_741);
xor U8459 (N_8459,N_3756,N_284);
and U8460 (N_8460,N_1765,N_3358);
nor U8461 (N_8461,N_3664,N_2485);
nand U8462 (N_8462,N_3254,N_549);
xnor U8463 (N_8463,N_3277,N_4332);
and U8464 (N_8464,N_1385,N_3327);
nor U8465 (N_8465,N_1579,N_799);
or U8466 (N_8466,N_1797,N_1259);
or U8467 (N_8467,N_2289,N_485);
xnor U8468 (N_8468,N_227,N_415);
nor U8469 (N_8469,N_1764,N_3241);
and U8470 (N_8470,N_3452,N_1328);
nand U8471 (N_8471,N_390,N_4150);
or U8472 (N_8472,N_1364,N_1990);
nand U8473 (N_8473,N_3560,N_3937);
or U8474 (N_8474,N_947,N_1996);
or U8475 (N_8475,N_3701,N_1525);
xnor U8476 (N_8476,N_4186,N_4253);
and U8477 (N_8477,N_3323,N_4041);
or U8478 (N_8478,N_1589,N_70);
or U8479 (N_8479,N_3227,N_2062);
or U8480 (N_8480,N_4085,N_1532);
or U8481 (N_8481,N_3264,N_3171);
or U8482 (N_8482,N_657,N_4073);
nor U8483 (N_8483,N_2394,N_2412);
nor U8484 (N_8484,N_3500,N_3580);
nor U8485 (N_8485,N_3484,N_1005);
nor U8486 (N_8486,N_29,N_1495);
or U8487 (N_8487,N_2903,N_4584);
nor U8488 (N_8488,N_1370,N_1713);
xnor U8489 (N_8489,N_4018,N_3854);
nor U8490 (N_8490,N_470,N_4486);
nor U8491 (N_8491,N_3486,N_2936);
or U8492 (N_8492,N_2607,N_869);
nor U8493 (N_8493,N_1579,N_1068);
or U8494 (N_8494,N_1487,N_4889);
or U8495 (N_8495,N_690,N_2030);
nand U8496 (N_8496,N_2753,N_4680);
xnor U8497 (N_8497,N_1145,N_62);
xnor U8498 (N_8498,N_1071,N_3146);
nand U8499 (N_8499,N_4120,N_2525);
nor U8500 (N_8500,N_1923,N_2793);
nor U8501 (N_8501,N_27,N_3110);
nand U8502 (N_8502,N_639,N_4368);
and U8503 (N_8503,N_1160,N_1563);
and U8504 (N_8504,N_3032,N_3660);
or U8505 (N_8505,N_1532,N_1816);
nor U8506 (N_8506,N_1505,N_3320);
and U8507 (N_8507,N_4506,N_2192);
or U8508 (N_8508,N_1011,N_3728);
nand U8509 (N_8509,N_3245,N_475);
nand U8510 (N_8510,N_4398,N_2365);
nand U8511 (N_8511,N_2346,N_304);
and U8512 (N_8512,N_4207,N_2426);
and U8513 (N_8513,N_3251,N_4063);
nand U8514 (N_8514,N_3441,N_220);
nand U8515 (N_8515,N_2261,N_3728);
nand U8516 (N_8516,N_4335,N_2806);
or U8517 (N_8517,N_3660,N_1789);
or U8518 (N_8518,N_1639,N_1256);
nor U8519 (N_8519,N_4983,N_1152);
and U8520 (N_8520,N_4193,N_2229);
nand U8521 (N_8521,N_1017,N_956);
and U8522 (N_8522,N_1085,N_280);
nor U8523 (N_8523,N_3850,N_2877);
or U8524 (N_8524,N_3268,N_3683);
and U8525 (N_8525,N_773,N_3105);
nand U8526 (N_8526,N_4123,N_1502);
and U8527 (N_8527,N_2654,N_989);
or U8528 (N_8528,N_4345,N_173);
nand U8529 (N_8529,N_4722,N_3772);
or U8530 (N_8530,N_2259,N_929);
nand U8531 (N_8531,N_1711,N_3308);
xor U8532 (N_8532,N_872,N_4656);
nor U8533 (N_8533,N_598,N_4640);
xor U8534 (N_8534,N_3874,N_3210);
or U8535 (N_8535,N_2466,N_2870);
nor U8536 (N_8536,N_1678,N_3911);
nor U8537 (N_8537,N_760,N_3952);
or U8538 (N_8538,N_1431,N_4884);
xor U8539 (N_8539,N_923,N_1835);
xor U8540 (N_8540,N_4871,N_1189);
xnor U8541 (N_8541,N_475,N_897);
xnor U8542 (N_8542,N_3746,N_2902);
or U8543 (N_8543,N_3675,N_747);
nor U8544 (N_8544,N_3515,N_104);
nand U8545 (N_8545,N_4706,N_477);
or U8546 (N_8546,N_1266,N_817);
nor U8547 (N_8547,N_3520,N_297);
or U8548 (N_8548,N_1469,N_539);
xor U8549 (N_8549,N_2429,N_2243);
nor U8550 (N_8550,N_2711,N_2599);
nand U8551 (N_8551,N_4838,N_411);
and U8552 (N_8552,N_4484,N_1652);
or U8553 (N_8553,N_2313,N_4604);
nor U8554 (N_8554,N_2327,N_676);
and U8555 (N_8555,N_4461,N_3382);
and U8556 (N_8556,N_1219,N_1341);
nand U8557 (N_8557,N_1325,N_2604);
and U8558 (N_8558,N_3387,N_2541);
or U8559 (N_8559,N_890,N_1652);
nor U8560 (N_8560,N_3848,N_3547);
nand U8561 (N_8561,N_2826,N_2280);
nor U8562 (N_8562,N_1557,N_2913);
and U8563 (N_8563,N_1057,N_4878);
nand U8564 (N_8564,N_4695,N_2667);
or U8565 (N_8565,N_858,N_3012);
and U8566 (N_8566,N_4720,N_2745);
and U8567 (N_8567,N_2789,N_4819);
nor U8568 (N_8568,N_354,N_2791);
xor U8569 (N_8569,N_986,N_1501);
xor U8570 (N_8570,N_3332,N_3787);
and U8571 (N_8571,N_553,N_1705);
or U8572 (N_8572,N_100,N_2149);
xnor U8573 (N_8573,N_452,N_3587);
nand U8574 (N_8574,N_2693,N_1450);
nand U8575 (N_8575,N_763,N_4220);
and U8576 (N_8576,N_4087,N_165);
or U8577 (N_8577,N_140,N_16);
or U8578 (N_8578,N_3374,N_3695);
or U8579 (N_8579,N_137,N_2621);
and U8580 (N_8580,N_2984,N_4514);
nand U8581 (N_8581,N_4162,N_3186);
nor U8582 (N_8582,N_1732,N_4582);
and U8583 (N_8583,N_368,N_3035);
nand U8584 (N_8584,N_3838,N_2956);
nor U8585 (N_8585,N_336,N_2254);
or U8586 (N_8586,N_1136,N_2100);
nor U8587 (N_8587,N_2927,N_1868);
or U8588 (N_8588,N_1032,N_4456);
nand U8589 (N_8589,N_3595,N_490);
and U8590 (N_8590,N_556,N_2998);
xnor U8591 (N_8591,N_4144,N_1699);
nor U8592 (N_8592,N_1665,N_2519);
nor U8593 (N_8593,N_1425,N_2595);
nand U8594 (N_8594,N_4444,N_1463);
and U8595 (N_8595,N_474,N_4935);
or U8596 (N_8596,N_2674,N_1867);
or U8597 (N_8597,N_2222,N_2574);
nand U8598 (N_8598,N_2455,N_6);
nor U8599 (N_8599,N_4766,N_1881);
and U8600 (N_8600,N_4944,N_4851);
xnor U8601 (N_8601,N_2181,N_4778);
or U8602 (N_8602,N_2518,N_1532);
xnor U8603 (N_8603,N_554,N_2791);
and U8604 (N_8604,N_3043,N_3048);
or U8605 (N_8605,N_4609,N_3497);
and U8606 (N_8606,N_3697,N_3964);
nand U8607 (N_8607,N_4008,N_3672);
and U8608 (N_8608,N_2167,N_198);
and U8609 (N_8609,N_4068,N_2279);
and U8610 (N_8610,N_1380,N_3779);
xnor U8611 (N_8611,N_438,N_4536);
nor U8612 (N_8612,N_2115,N_2186);
nor U8613 (N_8613,N_651,N_364);
nor U8614 (N_8614,N_3291,N_4024);
nor U8615 (N_8615,N_2237,N_436);
nor U8616 (N_8616,N_47,N_1932);
nor U8617 (N_8617,N_1732,N_3421);
or U8618 (N_8618,N_2403,N_3427);
nor U8619 (N_8619,N_4811,N_3867);
nor U8620 (N_8620,N_3536,N_4768);
xnor U8621 (N_8621,N_1667,N_4070);
xnor U8622 (N_8622,N_4448,N_2712);
and U8623 (N_8623,N_2716,N_3311);
and U8624 (N_8624,N_4848,N_3088);
xor U8625 (N_8625,N_3727,N_3033);
nor U8626 (N_8626,N_3569,N_3615);
and U8627 (N_8627,N_4493,N_2116);
and U8628 (N_8628,N_1745,N_3128);
nand U8629 (N_8629,N_1526,N_1138);
nor U8630 (N_8630,N_1611,N_1131);
and U8631 (N_8631,N_4820,N_4418);
or U8632 (N_8632,N_1542,N_872);
nand U8633 (N_8633,N_3902,N_1027);
nand U8634 (N_8634,N_3673,N_122);
xnor U8635 (N_8635,N_720,N_815);
or U8636 (N_8636,N_1190,N_250);
and U8637 (N_8637,N_724,N_531);
or U8638 (N_8638,N_1812,N_1507);
xor U8639 (N_8639,N_1260,N_4547);
nand U8640 (N_8640,N_2014,N_259);
or U8641 (N_8641,N_824,N_2722);
or U8642 (N_8642,N_2823,N_347);
xnor U8643 (N_8643,N_2128,N_2301);
or U8644 (N_8644,N_1385,N_1388);
and U8645 (N_8645,N_3062,N_1255);
or U8646 (N_8646,N_2967,N_4264);
or U8647 (N_8647,N_2881,N_3721);
nor U8648 (N_8648,N_164,N_290);
or U8649 (N_8649,N_404,N_724);
and U8650 (N_8650,N_873,N_3032);
nor U8651 (N_8651,N_2661,N_4847);
nor U8652 (N_8652,N_178,N_3116);
and U8653 (N_8653,N_2636,N_440);
nand U8654 (N_8654,N_3923,N_4263);
and U8655 (N_8655,N_2601,N_3122);
nand U8656 (N_8656,N_4227,N_1238);
nand U8657 (N_8657,N_2201,N_474);
and U8658 (N_8658,N_4190,N_3224);
xor U8659 (N_8659,N_366,N_672);
or U8660 (N_8660,N_1883,N_4618);
nand U8661 (N_8661,N_4672,N_3262);
or U8662 (N_8662,N_4546,N_175);
nor U8663 (N_8663,N_3897,N_3788);
or U8664 (N_8664,N_1511,N_102);
and U8665 (N_8665,N_325,N_670);
nand U8666 (N_8666,N_3701,N_3458);
xor U8667 (N_8667,N_586,N_795);
nor U8668 (N_8668,N_49,N_1296);
nand U8669 (N_8669,N_3838,N_1824);
nand U8670 (N_8670,N_3241,N_449);
xor U8671 (N_8671,N_1278,N_2007);
nor U8672 (N_8672,N_471,N_1253);
and U8673 (N_8673,N_4094,N_4613);
nand U8674 (N_8674,N_469,N_204);
nand U8675 (N_8675,N_1424,N_55);
and U8676 (N_8676,N_1185,N_439);
nand U8677 (N_8677,N_4278,N_3607);
nand U8678 (N_8678,N_914,N_1594);
or U8679 (N_8679,N_2200,N_88);
nand U8680 (N_8680,N_381,N_1193);
nor U8681 (N_8681,N_4440,N_601);
or U8682 (N_8682,N_3901,N_666);
or U8683 (N_8683,N_3052,N_1634);
nor U8684 (N_8684,N_2706,N_1032);
or U8685 (N_8685,N_1065,N_2405);
or U8686 (N_8686,N_2694,N_4288);
nand U8687 (N_8687,N_2512,N_2134);
and U8688 (N_8688,N_4994,N_4935);
or U8689 (N_8689,N_519,N_1540);
and U8690 (N_8690,N_1081,N_516);
nor U8691 (N_8691,N_1507,N_1128);
or U8692 (N_8692,N_340,N_1959);
nor U8693 (N_8693,N_4267,N_175);
and U8694 (N_8694,N_926,N_712);
nand U8695 (N_8695,N_1157,N_701);
or U8696 (N_8696,N_2183,N_204);
or U8697 (N_8697,N_4076,N_4275);
or U8698 (N_8698,N_2652,N_377);
and U8699 (N_8699,N_4830,N_1246);
nand U8700 (N_8700,N_530,N_2387);
or U8701 (N_8701,N_787,N_4115);
or U8702 (N_8702,N_633,N_3671);
nor U8703 (N_8703,N_3566,N_3809);
or U8704 (N_8704,N_4035,N_1010);
xor U8705 (N_8705,N_2438,N_2643);
nor U8706 (N_8706,N_58,N_3500);
nor U8707 (N_8707,N_758,N_3696);
nor U8708 (N_8708,N_2948,N_904);
nand U8709 (N_8709,N_3691,N_3283);
nor U8710 (N_8710,N_700,N_2598);
nand U8711 (N_8711,N_3329,N_1284);
or U8712 (N_8712,N_1119,N_3531);
nor U8713 (N_8713,N_165,N_3139);
nand U8714 (N_8714,N_3693,N_2893);
nand U8715 (N_8715,N_3561,N_1402);
and U8716 (N_8716,N_1389,N_3024);
nor U8717 (N_8717,N_3651,N_1447);
nor U8718 (N_8718,N_264,N_489);
or U8719 (N_8719,N_4403,N_4924);
or U8720 (N_8720,N_4425,N_2481);
nor U8721 (N_8721,N_1728,N_370);
nor U8722 (N_8722,N_2142,N_1017);
or U8723 (N_8723,N_4059,N_4887);
nor U8724 (N_8724,N_2106,N_2830);
xor U8725 (N_8725,N_3147,N_3660);
nand U8726 (N_8726,N_4817,N_2776);
and U8727 (N_8727,N_3742,N_2591);
nor U8728 (N_8728,N_2069,N_205);
or U8729 (N_8729,N_1126,N_455);
nand U8730 (N_8730,N_557,N_1730);
or U8731 (N_8731,N_2614,N_4036);
nor U8732 (N_8732,N_3813,N_4111);
or U8733 (N_8733,N_94,N_3110);
nor U8734 (N_8734,N_4794,N_3612);
and U8735 (N_8735,N_3585,N_3681);
or U8736 (N_8736,N_2708,N_90);
and U8737 (N_8737,N_3687,N_4932);
and U8738 (N_8738,N_1222,N_335);
nor U8739 (N_8739,N_58,N_3435);
nand U8740 (N_8740,N_2592,N_591);
nor U8741 (N_8741,N_3105,N_1904);
nand U8742 (N_8742,N_3076,N_846);
or U8743 (N_8743,N_2149,N_2987);
nand U8744 (N_8744,N_2299,N_3036);
and U8745 (N_8745,N_1073,N_3341);
and U8746 (N_8746,N_4603,N_3082);
and U8747 (N_8747,N_4077,N_1766);
or U8748 (N_8748,N_2143,N_4789);
nor U8749 (N_8749,N_155,N_2807);
xor U8750 (N_8750,N_4225,N_3698);
nand U8751 (N_8751,N_4122,N_458);
nand U8752 (N_8752,N_51,N_2934);
nor U8753 (N_8753,N_1917,N_229);
nor U8754 (N_8754,N_1379,N_1787);
and U8755 (N_8755,N_699,N_4877);
nor U8756 (N_8756,N_2918,N_4093);
or U8757 (N_8757,N_302,N_135);
and U8758 (N_8758,N_204,N_3781);
and U8759 (N_8759,N_1641,N_1967);
or U8760 (N_8760,N_1855,N_1376);
or U8761 (N_8761,N_2149,N_1511);
nor U8762 (N_8762,N_1712,N_804);
nand U8763 (N_8763,N_1550,N_533);
or U8764 (N_8764,N_3878,N_869);
nor U8765 (N_8765,N_2286,N_3025);
and U8766 (N_8766,N_117,N_452);
nand U8767 (N_8767,N_2309,N_1590);
nor U8768 (N_8768,N_3370,N_1434);
and U8769 (N_8769,N_1603,N_2913);
and U8770 (N_8770,N_1202,N_4627);
nor U8771 (N_8771,N_968,N_2253);
nand U8772 (N_8772,N_3956,N_389);
nand U8773 (N_8773,N_3067,N_4715);
xnor U8774 (N_8774,N_2004,N_2732);
and U8775 (N_8775,N_3235,N_3448);
nand U8776 (N_8776,N_4100,N_2406);
and U8777 (N_8777,N_553,N_3029);
or U8778 (N_8778,N_1809,N_3752);
and U8779 (N_8779,N_4968,N_3393);
and U8780 (N_8780,N_1007,N_4310);
and U8781 (N_8781,N_1552,N_672);
or U8782 (N_8782,N_809,N_4199);
nand U8783 (N_8783,N_2431,N_4799);
nor U8784 (N_8784,N_2383,N_2122);
nor U8785 (N_8785,N_2728,N_1889);
or U8786 (N_8786,N_2299,N_3835);
and U8787 (N_8787,N_450,N_4450);
and U8788 (N_8788,N_3584,N_1218);
nor U8789 (N_8789,N_4728,N_404);
xor U8790 (N_8790,N_731,N_4075);
nand U8791 (N_8791,N_1400,N_2883);
and U8792 (N_8792,N_2125,N_185);
nor U8793 (N_8793,N_4042,N_4904);
nor U8794 (N_8794,N_1909,N_886);
and U8795 (N_8795,N_806,N_506);
xor U8796 (N_8796,N_3425,N_1683);
or U8797 (N_8797,N_1777,N_1212);
nand U8798 (N_8798,N_3483,N_4952);
or U8799 (N_8799,N_1377,N_2726);
or U8800 (N_8800,N_1228,N_2679);
xor U8801 (N_8801,N_3061,N_4239);
or U8802 (N_8802,N_2321,N_3050);
nor U8803 (N_8803,N_1312,N_1618);
or U8804 (N_8804,N_4010,N_772);
nand U8805 (N_8805,N_3695,N_2739);
or U8806 (N_8806,N_2499,N_28);
or U8807 (N_8807,N_749,N_4793);
and U8808 (N_8808,N_1717,N_4481);
or U8809 (N_8809,N_240,N_2187);
nand U8810 (N_8810,N_3819,N_2400);
nor U8811 (N_8811,N_2966,N_997);
and U8812 (N_8812,N_2416,N_4878);
xnor U8813 (N_8813,N_1665,N_1404);
and U8814 (N_8814,N_867,N_3844);
or U8815 (N_8815,N_4806,N_4655);
and U8816 (N_8816,N_2341,N_4398);
or U8817 (N_8817,N_3397,N_2121);
nand U8818 (N_8818,N_4952,N_1863);
nand U8819 (N_8819,N_3749,N_4621);
nand U8820 (N_8820,N_2065,N_4148);
xnor U8821 (N_8821,N_2434,N_875);
nand U8822 (N_8822,N_3350,N_1933);
or U8823 (N_8823,N_1679,N_93);
xor U8824 (N_8824,N_4369,N_4733);
xor U8825 (N_8825,N_4739,N_305);
or U8826 (N_8826,N_4981,N_677);
or U8827 (N_8827,N_336,N_4344);
and U8828 (N_8828,N_4834,N_3956);
and U8829 (N_8829,N_2132,N_3750);
nor U8830 (N_8830,N_3392,N_1337);
and U8831 (N_8831,N_535,N_3270);
xnor U8832 (N_8832,N_1454,N_3641);
nor U8833 (N_8833,N_2397,N_1430);
nor U8834 (N_8834,N_3996,N_1816);
and U8835 (N_8835,N_1048,N_4644);
xnor U8836 (N_8836,N_1752,N_2030);
nor U8837 (N_8837,N_2214,N_1052);
nor U8838 (N_8838,N_3144,N_1224);
or U8839 (N_8839,N_4005,N_4800);
nor U8840 (N_8840,N_220,N_428);
nor U8841 (N_8841,N_4689,N_1794);
nand U8842 (N_8842,N_4032,N_4482);
nand U8843 (N_8843,N_4920,N_2108);
nor U8844 (N_8844,N_1794,N_2693);
and U8845 (N_8845,N_3046,N_4966);
or U8846 (N_8846,N_3377,N_2000);
and U8847 (N_8847,N_397,N_1804);
nor U8848 (N_8848,N_609,N_3042);
or U8849 (N_8849,N_2320,N_1777);
and U8850 (N_8850,N_1464,N_1792);
or U8851 (N_8851,N_2996,N_3277);
or U8852 (N_8852,N_3030,N_203);
and U8853 (N_8853,N_730,N_85);
or U8854 (N_8854,N_4506,N_2434);
nand U8855 (N_8855,N_94,N_282);
and U8856 (N_8856,N_3835,N_1634);
nor U8857 (N_8857,N_3354,N_2703);
nor U8858 (N_8858,N_2873,N_3152);
xnor U8859 (N_8859,N_1242,N_2413);
and U8860 (N_8860,N_3127,N_62);
and U8861 (N_8861,N_661,N_2332);
or U8862 (N_8862,N_3431,N_711);
nand U8863 (N_8863,N_1030,N_4476);
or U8864 (N_8864,N_3183,N_761);
and U8865 (N_8865,N_4261,N_3365);
nand U8866 (N_8866,N_623,N_1923);
nor U8867 (N_8867,N_4118,N_534);
or U8868 (N_8868,N_2260,N_3859);
nand U8869 (N_8869,N_1890,N_1540);
or U8870 (N_8870,N_3052,N_1097);
nand U8871 (N_8871,N_3131,N_1337);
and U8872 (N_8872,N_4770,N_1594);
nand U8873 (N_8873,N_1657,N_484);
or U8874 (N_8874,N_759,N_238);
xnor U8875 (N_8875,N_1892,N_4768);
or U8876 (N_8876,N_2433,N_4345);
or U8877 (N_8877,N_3856,N_3127);
or U8878 (N_8878,N_2977,N_2626);
or U8879 (N_8879,N_199,N_479);
or U8880 (N_8880,N_4550,N_4994);
nor U8881 (N_8881,N_1857,N_2609);
and U8882 (N_8882,N_3889,N_1979);
nand U8883 (N_8883,N_2494,N_4824);
and U8884 (N_8884,N_34,N_3008);
nand U8885 (N_8885,N_3942,N_1968);
nor U8886 (N_8886,N_3348,N_1776);
nand U8887 (N_8887,N_4448,N_4262);
nand U8888 (N_8888,N_1586,N_3009);
nor U8889 (N_8889,N_1426,N_20);
nand U8890 (N_8890,N_1809,N_1965);
nor U8891 (N_8891,N_42,N_1096);
nor U8892 (N_8892,N_3066,N_1034);
nand U8893 (N_8893,N_3462,N_2843);
xor U8894 (N_8894,N_3858,N_4956);
xnor U8895 (N_8895,N_419,N_2382);
or U8896 (N_8896,N_541,N_4243);
or U8897 (N_8897,N_2658,N_3427);
xnor U8898 (N_8898,N_4268,N_3690);
and U8899 (N_8899,N_452,N_4156);
or U8900 (N_8900,N_4786,N_3596);
xor U8901 (N_8901,N_995,N_1466);
nand U8902 (N_8902,N_7,N_3226);
and U8903 (N_8903,N_3640,N_2368);
and U8904 (N_8904,N_3683,N_4348);
nor U8905 (N_8905,N_1346,N_3467);
and U8906 (N_8906,N_1551,N_3050);
nor U8907 (N_8907,N_1530,N_3897);
nor U8908 (N_8908,N_3411,N_353);
xnor U8909 (N_8909,N_2425,N_4821);
or U8910 (N_8910,N_1464,N_2889);
and U8911 (N_8911,N_3495,N_2389);
nand U8912 (N_8912,N_2068,N_1925);
and U8913 (N_8913,N_2589,N_3091);
and U8914 (N_8914,N_1804,N_1499);
nor U8915 (N_8915,N_3022,N_2448);
and U8916 (N_8916,N_1416,N_1061);
or U8917 (N_8917,N_4658,N_3301);
nor U8918 (N_8918,N_3361,N_3651);
xor U8919 (N_8919,N_4328,N_4152);
nor U8920 (N_8920,N_397,N_1096);
nand U8921 (N_8921,N_4940,N_1711);
or U8922 (N_8922,N_3813,N_1363);
or U8923 (N_8923,N_2132,N_4025);
nand U8924 (N_8924,N_4204,N_1356);
or U8925 (N_8925,N_3653,N_1798);
or U8926 (N_8926,N_2653,N_3253);
and U8927 (N_8927,N_4475,N_4164);
or U8928 (N_8928,N_989,N_2870);
xnor U8929 (N_8929,N_1514,N_3905);
nand U8930 (N_8930,N_3021,N_3058);
nand U8931 (N_8931,N_470,N_1345);
or U8932 (N_8932,N_4669,N_1156);
or U8933 (N_8933,N_3237,N_849);
nand U8934 (N_8934,N_1747,N_3687);
and U8935 (N_8935,N_4680,N_1990);
and U8936 (N_8936,N_4642,N_4444);
or U8937 (N_8937,N_1761,N_3017);
nor U8938 (N_8938,N_3012,N_949);
xnor U8939 (N_8939,N_1867,N_240);
and U8940 (N_8940,N_1456,N_2892);
and U8941 (N_8941,N_122,N_3392);
nor U8942 (N_8942,N_3743,N_1337);
or U8943 (N_8943,N_3953,N_1360);
xor U8944 (N_8944,N_2717,N_4179);
and U8945 (N_8945,N_51,N_121);
nor U8946 (N_8946,N_1727,N_3340);
nor U8947 (N_8947,N_3938,N_3882);
xor U8948 (N_8948,N_3597,N_2159);
and U8949 (N_8949,N_4563,N_3327);
nand U8950 (N_8950,N_2248,N_3292);
nor U8951 (N_8951,N_2834,N_2245);
nor U8952 (N_8952,N_2275,N_2213);
and U8953 (N_8953,N_4328,N_2382);
and U8954 (N_8954,N_3033,N_2433);
or U8955 (N_8955,N_3019,N_4468);
or U8956 (N_8956,N_4813,N_3567);
nor U8957 (N_8957,N_3575,N_4932);
and U8958 (N_8958,N_1016,N_3051);
nor U8959 (N_8959,N_101,N_4851);
nor U8960 (N_8960,N_2930,N_2580);
nand U8961 (N_8961,N_4738,N_247);
nor U8962 (N_8962,N_1548,N_1227);
or U8963 (N_8963,N_3652,N_523);
nand U8964 (N_8964,N_4244,N_4568);
nor U8965 (N_8965,N_1691,N_3692);
or U8966 (N_8966,N_3233,N_2680);
or U8967 (N_8967,N_1236,N_1447);
nand U8968 (N_8968,N_71,N_4606);
nor U8969 (N_8969,N_3038,N_3902);
xnor U8970 (N_8970,N_2138,N_4101);
xor U8971 (N_8971,N_4879,N_940);
nor U8972 (N_8972,N_778,N_3982);
and U8973 (N_8973,N_2550,N_398);
or U8974 (N_8974,N_3403,N_4985);
xnor U8975 (N_8975,N_3703,N_1778);
or U8976 (N_8976,N_4746,N_4867);
or U8977 (N_8977,N_1847,N_249);
and U8978 (N_8978,N_4873,N_4783);
and U8979 (N_8979,N_4153,N_2711);
and U8980 (N_8980,N_796,N_1725);
or U8981 (N_8981,N_4696,N_2591);
and U8982 (N_8982,N_3374,N_2657);
and U8983 (N_8983,N_3024,N_4745);
and U8984 (N_8984,N_282,N_2865);
or U8985 (N_8985,N_2688,N_2694);
and U8986 (N_8986,N_777,N_1554);
or U8987 (N_8987,N_4836,N_786);
and U8988 (N_8988,N_3342,N_3644);
nor U8989 (N_8989,N_992,N_4988);
nand U8990 (N_8990,N_1188,N_1713);
or U8991 (N_8991,N_2103,N_3708);
nor U8992 (N_8992,N_1137,N_535);
nand U8993 (N_8993,N_632,N_4220);
nand U8994 (N_8994,N_4169,N_4099);
nor U8995 (N_8995,N_3369,N_2522);
nor U8996 (N_8996,N_4862,N_2936);
and U8997 (N_8997,N_3743,N_1207);
xnor U8998 (N_8998,N_327,N_261);
nor U8999 (N_8999,N_1468,N_4757);
and U9000 (N_9000,N_3226,N_4545);
nand U9001 (N_9001,N_3663,N_18);
and U9002 (N_9002,N_1193,N_1908);
and U9003 (N_9003,N_2618,N_965);
xnor U9004 (N_9004,N_1591,N_927);
nand U9005 (N_9005,N_1960,N_843);
and U9006 (N_9006,N_3991,N_3338);
nand U9007 (N_9007,N_3253,N_4794);
and U9008 (N_9008,N_3359,N_2808);
and U9009 (N_9009,N_1568,N_2404);
nor U9010 (N_9010,N_4580,N_1076);
nand U9011 (N_9011,N_1436,N_400);
nand U9012 (N_9012,N_2412,N_2461);
nor U9013 (N_9013,N_3821,N_3794);
nor U9014 (N_9014,N_4255,N_2607);
and U9015 (N_9015,N_2792,N_574);
and U9016 (N_9016,N_3900,N_945);
xor U9017 (N_9017,N_1073,N_2027);
nand U9018 (N_9018,N_3446,N_4452);
and U9019 (N_9019,N_985,N_3822);
nor U9020 (N_9020,N_2366,N_2194);
nor U9021 (N_9021,N_1563,N_1557);
and U9022 (N_9022,N_99,N_4819);
and U9023 (N_9023,N_541,N_736);
or U9024 (N_9024,N_3248,N_3938);
or U9025 (N_9025,N_995,N_1522);
xnor U9026 (N_9026,N_3209,N_3513);
nor U9027 (N_9027,N_3101,N_4627);
xnor U9028 (N_9028,N_3442,N_3984);
or U9029 (N_9029,N_4461,N_667);
or U9030 (N_9030,N_2056,N_4127);
and U9031 (N_9031,N_1549,N_3409);
and U9032 (N_9032,N_2311,N_2061);
nor U9033 (N_9033,N_4229,N_2937);
nand U9034 (N_9034,N_614,N_2223);
and U9035 (N_9035,N_4987,N_3201);
nor U9036 (N_9036,N_4148,N_4485);
or U9037 (N_9037,N_1482,N_2356);
nand U9038 (N_9038,N_2098,N_4960);
nor U9039 (N_9039,N_2736,N_425);
or U9040 (N_9040,N_3428,N_1637);
and U9041 (N_9041,N_1718,N_1397);
and U9042 (N_9042,N_1004,N_4656);
and U9043 (N_9043,N_24,N_3376);
nor U9044 (N_9044,N_2325,N_3149);
and U9045 (N_9045,N_2336,N_1553);
xor U9046 (N_9046,N_552,N_2073);
and U9047 (N_9047,N_3062,N_731);
nand U9048 (N_9048,N_845,N_4908);
or U9049 (N_9049,N_3490,N_835);
xor U9050 (N_9050,N_2072,N_1396);
nor U9051 (N_9051,N_1926,N_4672);
xnor U9052 (N_9052,N_1112,N_694);
nand U9053 (N_9053,N_1728,N_802);
or U9054 (N_9054,N_2062,N_3763);
or U9055 (N_9055,N_3580,N_2893);
or U9056 (N_9056,N_4026,N_211);
and U9057 (N_9057,N_2402,N_1558);
or U9058 (N_9058,N_1116,N_372);
nor U9059 (N_9059,N_2381,N_1893);
nand U9060 (N_9060,N_2796,N_1053);
or U9061 (N_9061,N_2268,N_2177);
or U9062 (N_9062,N_1536,N_4130);
nor U9063 (N_9063,N_4731,N_36);
nand U9064 (N_9064,N_2952,N_4594);
nor U9065 (N_9065,N_4721,N_1575);
or U9066 (N_9066,N_3759,N_4196);
xnor U9067 (N_9067,N_1922,N_2614);
nand U9068 (N_9068,N_1210,N_1256);
and U9069 (N_9069,N_3525,N_4279);
nand U9070 (N_9070,N_829,N_1404);
nand U9071 (N_9071,N_2057,N_923);
and U9072 (N_9072,N_1382,N_380);
or U9073 (N_9073,N_3292,N_1302);
nor U9074 (N_9074,N_4383,N_2585);
xor U9075 (N_9075,N_1937,N_3842);
and U9076 (N_9076,N_1010,N_3682);
nor U9077 (N_9077,N_4319,N_1492);
nand U9078 (N_9078,N_2226,N_4007);
and U9079 (N_9079,N_918,N_3005);
or U9080 (N_9080,N_1149,N_1064);
nand U9081 (N_9081,N_3512,N_530);
or U9082 (N_9082,N_4511,N_1162);
xor U9083 (N_9083,N_1298,N_1443);
and U9084 (N_9084,N_2111,N_4941);
and U9085 (N_9085,N_3781,N_1181);
and U9086 (N_9086,N_900,N_4970);
xor U9087 (N_9087,N_1341,N_3704);
and U9088 (N_9088,N_2915,N_1234);
or U9089 (N_9089,N_324,N_1125);
nand U9090 (N_9090,N_202,N_2976);
nand U9091 (N_9091,N_2829,N_1909);
xnor U9092 (N_9092,N_4857,N_3804);
nor U9093 (N_9093,N_1549,N_1404);
nor U9094 (N_9094,N_1636,N_2242);
nor U9095 (N_9095,N_587,N_456);
nand U9096 (N_9096,N_4575,N_543);
nor U9097 (N_9097,N_2827,N_1155);
xor U9098 (N_9098,N_3878,N_3924);
nand U9099 (N_9099,N_3171,N_4309);
nor U9100 (N_9100,N_2121,N_3698);
nor U9101 (N_9101,N_2382,N_3205);
and U9102 (N_9102,N_3271,N_1056);
xnor U9103 (N_9103,N_2909,N_2203);
xnor U9104 (N_9104,N_1948,N_2179);
and U9105 (N_9105,N_4252,N_1167);
nor U9106 (N_9106,N_1767,N_3454);
and U9107 (N_9107,N_2964,N_349);
nand U9108 (N_9108,N_1423,N_474);
nor U9109 (N_9109,N_653,N_3246);
xnor U9110 (N_9110,N_1522,N_361);
nand U9111 (N_9111,N_4240,N_4994);
nand U9112 (N_9112,N_3805,N_3365);
nand U9113 (N_9113,N_1560,N_727);
and U9114 (N_9114,N_1728,N_2851);
or U9115 (N_9115,N_1277,N_4374);
nor U9116 (N_9116,N_4812,N_1384);
or U9117 (N_9117,N_3991,N_2411);
nand U9118 (N_9118,N_4584,N_1786);
or U9119 (N_9119,N_231,N_2741);
or U9120 (N_9120,N_61,N_904);
and U9121 (N_9121,N_1895,N_2358);
nand U9122 (N_9122,N_4505,N_4923);
and U9123 (N_9123,N_1601,N_744);
nand U9124 (N_9124,N_4482,N_1974);
nor U9125 (N_9125,N_4723,N_4780);
nor U9126 (N_9126,N_48,N_4590);
nand U9127 (N_9127,N_4140,N_983);
xnor U9128 (N_9128,N_4,N_4416);
nor U9129 (N_9129,N_2580,N_2257);
nor U9130 (N_9130,N_4955,N_1226);
nor U9131 (N_9131,N_4922,N_2429);
nand U9132 (N_9132,N_2593,N_1010);
and U9133 (N_9133,N_4557,N_971);
nor U9134 (N_9134,N_2910,N_3841);
and U9135 (N_9135,N_1037,N_1165);
and U9136 (N_9136,N_951,N_1152);
nand U9137 (N_9137,N_716,N_2804);
and U9138 (N_9138,N_4943,N_3229);
nor U9139 (N_9139,N_3041,N_4082);
or U9140 (N_9140,N_3226,N_3199);
nor U9141 (N_9141,N_3590,N_3644);
nor U9142 (N_9142,N_2805,N_627);
or U9143 (N_9143,N_4859,N_3593);
nor U9144 (N_9144,N_4708,N_2436);
nor U9145 (N_9145,N_498,N_3451);
nand U9146 (N_9146,N_4277,N_3929);
nor U9147 (N_9147,N_4823,N_4746);
nor U9148 (N_9148,N_972,N_1377);
and U9149 (N_9149,N_4646,N_1295);
or U9150 (N_9150,N_2993,N_67);
and U9151 (N_9151,N_1294,N_4165);
nor U9152 (N_9152,N_4133,N_1156);
or U9153 (N_9153,N_2022,N_4334);
and U9154 (N_9154,N_4112,N_4378);
or U9155 (N_9155,N_48,N_264);
nand U9156 (N_9156,N_3537,N_933);
nor U9157 (N_9157,N_1058,N_1644);
nor U9158 (N_9158,N_3425,N_2479);
xor U9159 (N_9159,N_510,N_4703);
nor U9160 (N_9160,N_1356,N_4909);
xor U9161 (N_9161,N_2445,N_784);
xor U9162 (N_9162,N_2411,N_4169);
and U9163 (N_9163,N_4679,N_205);
xor U9164 (N_9164,N_1077,N_653);
or U9165 (N_9165,N_3555,N_1309);
nor U9166 (N_9166,N_4713,N_1360);
and U9167 (N_9167,N_984,N_670);
xor U9168 (N_9168,N_2417,N_2999);
nor U9169 (N_9169,N_2901,N_1548);
nand U9170 (N_9170,N_3909,N_1757);
or U9171 (N_9171,N_1399,N_2007);
nand U9172 (N_9172,N_580,N_1622);
nor U9173 (N_9173,N_3968,N_3771);
and U9174 (N_9174,N_3678,N_786);
or U9175 (N_9175,N_845,N_4242);
nand U9176 (N_9176,N_4714,N_2979);
or U9177 (N_9177,N_2690,N_3351);
nand U9178 (N_9178,N_544,N_1799);
nor U9179 (N_9179,N_1793,N_1506);
or U9180 (N_9180,N_2734,N_1903);
xor U9181 (N_9181,N_700,N_422);
nand U9182 (N_9182,N_2442,N_2106);
nor U9183 (N_9183,N_436,N_3526);
and U9184 (N_9184,N_4820,N_1362);
xnor U9185 (N_9185,N_3889,N_2582);
or U9186 (N_9186,N_2447,N_1549);
and U9187 (N_9187,N_111,N_3352);
or U9188 (N_9188,N_660,N_2071);
or U9189 (N_9189,N_1319,N_4176);
and U9190 (N_9190,N_1194,N_4026);
nor U9191 (N_9191,N_4587,N_2785);
nor U9192 (N_9192,N_45,N_1346);
or U9193 (N_9193,N_3194,N_500);
xnor U9194 (N_9194,N_237,N_1892);
nor U9195 (N_9195,N_1587,N_1293);
or U9196 (N_9196,N_3556,N_2058);
nand U9197 (N_9197,N_2283,N_2803);
nand U9198 (N_9198,N_1223,N_864);
and U9199 (N_9199,N_4499,N_3435);
and U9200 (N_9200,N_3643,N_3023);
or U9201 (N_9201,N_2604,N_851);
nor U9202 (N_9202,N_722,N_4678);
nor U9203 (N_9203,N_693,N_945);
or U9204 (N_9204,N_332,N_2376);
and U9205 (N_9205,N_3998,N_2389);
nand U9206 (N_9206,N_3849,N_3171);
and U9207 (N_9207,N_2275,N_4107);
or U9208 (N_9208,N_1015,N_2460);
xnor U9209 (N_9209,N_2819,N_1102);
and U9210 (N_9210,N_4053,N_2823);
nand U9211 (N_9211,N_1863,N_4894);
nor U9212 (N_9212,N_3494,N_2215);
nor U9213 (N_9213,N_1418,N_2166);
xor U9214 (N_9214,N_1923,N_1553);
nand U9215 (N_9215,N_1965,N_1339);
and U9216 (N_9216,N_2104,N_2846);
nand U9217 (N_9217,N_3636,N_3070);
xor U9218 (N_9218,N_2296,N_708);
and U9219 (N_9219,N_546,N_4135);
or U9220 (N_9220,N_12,N_3064);
and U9221 (N_9221,N_4551,N_182);
nand U9222 (N_9222,N_685,N_2883);
and U9223 (N_9223,N_1754,N_3871);
or U9224 (N_9224,N_3496,N_4761);
nand U9225 (N_9225,N_4822,N_1235);
nor U9226 (N_9226,N_2459,N_89);
or U9227 (N_9227,N_2025,N_1956);
or U9228 (N_9228,N_3913,N_488);
or U9229 (N_9229,N_4831,N_995);
nand U9230 (N_9230,N_4970,N_1216);
nor U9231 (N_9231,N_3390,N_2445);
nand U9232 (N_9232,N_2445,N_854);
nor U9233 (N_9233,N_4360,N_4517);
nand U9234 (N_9234,N_2448,N_1341);
nand U9235 (N_9235,N_4152,N_3338);
and U9236 (N_9236,N_1140,N_3767);
or U9237 (N_9237,N_4892,N_2869);
nand U9238 (N_9238,N_175,N_2893);
nor U9239 (N_9239,N_779,N_1956);
nor U9240 (N_9240,N_506,N_3222);
and U9241 (N_9241,N_131,N_4140);
nor U9242 (N_9242,N_1286,N_170);
nor U9243 (N_9243,N_2745,N_97);
and U9244 (N_9244,N_1943,N_4377);
and U9245 (N_9245,N_2820,N_3364);
or U9246 (N_9246,N_2514,N_2206);
or U9247 (N_9247,N_1722,N_3178);
nor U9248 (N_9248,N_2619,N_2991);
xor U9249 (N_9249,N_2459,N_143);
nand U9250 (N_9250,N_788,N_4559);
and U9251 (N_9251,N_3910,N_3974);
and U9252 (N_9252,N_2476,N_1065);
and U9253 (N_9253,N_2178,N_4279);
nand U9254 (N_9254,N_1314,N_1539);
nand U9255 (N_9255,N_403,N_3153);
nand U9256 (N_9256,N_4843,N_873);
nor U9257 (N_9257,N_4736,N_2002);
nor U9258 (N_9258,N_3110,N_1143);
nand U9259 (N_9259,N_234,N_2396);
nand U9260 (N_9260,N_1472,N_2024);
and U9261 (N_9261,N_4341,N_3979);
nor U9262 (N_9262,N_2979,N_4016);
or U9263 (N_9263,N_1442,N_4847);
and U9264 (N_9264,N_454,N_3094);
or U9265 (N_9265,N_506,N_1737);
and U9266 (N_9266,N_1521,N_2229);
or U9267 (N_9267,N_4584,N_4324);
nand U9268 (N_9268,N_3864,N_4284);
and U9269 (N_9269,N_617,N_4083);
nor U9270 (N_9270,N_4582,N_157);
and U9271 (N_9271,N_3452,N_3890);
nand U9272 (N_9272,N_2378,N_3122);
nand U9273 (N_9273,N_2323,N_1719);
and U9274 (N_9274,N_4162,N_4939);
nand U9275 (N_9275,N_3628,N_3239);
nand U9276 (N_9276,N_4242,N_4235);
and U9277 (N_9277,N_2786,N_2772);
nand U9278 (N_9278,N_2543,N_3427);
nand U9279 (N_9279,N_3088,N_3490);
and U9280 (N_9280,N_3530,N_1154);
or U9281 (N_9281,N_2791,N_1820);
nand U9282 (N_9282,N_4745,N_2619);
nor U9283 (N_9283,N_1692,N_110);
or U9284 (N_9284,N_410,N_3186);
xor U9285 (N_9285,N_199,N_2240);
nand U9286 (N_9286,N_721,N_596);
or U9287 (N_9287,N_4287,N_1606);
or U9288 (N_9288,N_4637,N_4975);
or U9289 (N_9289,N_3237,N_3277);
xnor U9290 (N_9290,N_1620,N_3946);
nand U9291 (N_9291,N_3572,N_4370);
nor U9292 (N_9292,N_687,N_4663);
nand U9293 (N_9293,N_1058,N_1249);
or U9294 (N_9294,N_3561,N_4103);
or U9295 (N_9295,N_4365,N_482);
nand U9296 (N_9296,N_4917,N_1142);
or U9297 (N_9297,N_2541,N_1989);
xor U9298 (N_9298,N_194,N_4377);
nor U9299 (N_9299,N_1365,N_4758);
or U9300 (N_9300,N_938,N_2489);
or U9301 (N_9301,N_617,N_9);
nand U9302 (N_9302,N_4508,N_465);
nor U9303 (N_9303,N_1668,N_820);
or U9304 (N_9304,N_1310,N_4063);
nor U9305 (N_9305,N_1643,N_3108);
nor U9306 (N_9306,N_404,N_904);
nand U9307 (N_9307,N_3027,N_2068);
or U9308 (N_9308,N_3880,N_4383);
xor U9309 (N_9309,N_510,N_2605);
xnor U9310 (N_9310,N_2934,N_3376);
nand U9311 (N_9311,N_4465,N_4367);
nand U9312 (N_9312,N_3698,N_2170);
nand U9313 (N_9313,N_4092,N_4011);
nor U9314 (N_9314,N_3428,N_3025);
nand U9315 (N_9315,N_3402,N_2285);
and U9316 (N_9316,N_495,N_3133);
nand U9317 (N_9317,N_1157,N_778);
or U9318 (N_9318,N_2232,N_3920);
nand U9319 (N_9319,N_4533,N_4339);
xnor U9320 (N_9320,N_3813,N_4776);
xnor U9321 (N_9321,N_150,N_1993);
nand U9322 (N_9322,N_3387,N_4271);
nor U9323 (N_9323,N_3625,N_4646);
nand U9324 (N_9324,N_4250,N_965);
nand U9325 (N_9325,N_3228,N_2978);
nor U9326 (N_9326,N_3847,N_586);
xnor U9327 (N_9327,N_1830,N_67);
and U9328 (N_9328,N_1998,N_488);
nor U9329 (N_9329,N_4033,N_1337);
xnor U9330 (N_9330,N_351,N_781);
or U9331 (N_9331,N_469,N_4457);
nand U9332 (N_9332,N_4859,N_1349);
nor U9333 (N_9333,N_3875,N_139);
or U9334 (N_9334,N_1701,N_527);
and U9335 (N_9335,N_3833,N_4713);
or U9336 (N_9336,N_2163,N_3635);
and U9337 (N_9337,N_4696,N_2438);
nor U9338 (N_9338,N_4550,N_3572);
and U9339 (N_9339,N_3898,N_359);
xor U9340 (N_9340,N_1732,N_1095);
and U9341 (N_9341,N_2495,N_1242);
xnor U9342 (N_9342,N_3201,N_511);
or U9343 (N_9343,N_3436,N_4020);
or U9344 (N_9344,N_3121,N_2892);
nand U9345 (N_9345,N_1422,N_3386);
or U9346 (N_9346,N_3435,N_3543);
nor U9347 (N_9347,N_4421,N_2814);
nor U9348 (N_9348,N_3728,N_3990);
and U9349 (N_9349,N_1364,N_3348);
or U9350 (N_9350,N_1609,N_4905);
and U9351 (N_9351,N_2071,N_4834);
nor U9352 (N_9352,N_2370,N_1762);
or U9353 (N_9353,N_2499,N_3500);
nor U9354 (N_9354,N_1847,N_1856);
nor U9355 (N_9355,N_3234,N_3775);
or U9356 (N_9356,N_366,N_382);
or U9357 (N_9357,N_2018,N_4377);
nor U9358 (N_9358,N_2153,N_1813);
and U9359 (N_9359,N_4527,N_2272);
xor U9360 (N_9360,N_1302,N_3320);
or U9361 (N_9361,N_3736,N_2854);
or U9362 (N_9362,N_3850,N_1428);
xnor U9363 (N_9363,N_4096,N_2165);
nand U9364 (N_9364,N_3546,N_4842);
and U9365 (N_9365,N_1437,N_4542);
nand U9366 (N_9366,N_4435,N_3796);
and U9367 (N_9367,N_4632,N_4201);
xor U9368 (N_9368,N_4348,N_4584);
xor U9369 (N_9369,N_4167,N_319);
nand U9370 (N_9370,N_276,N_3858);
or U9371 (N_9371,N_2314,N_3897);
nand U9372 (N_9372,N_776,N_527);
xor U9373 (N_9373,N_778,N_3049);
and U9374 (N_9374,N_4927,N_4452);
and U9375 (N_9375,N_3974,N_259);
or U9376 (N_9376,N_3971,N_103);
nor U9377 (N_9377,N_2837,N_4891);
xnor U9378 (N_9378,N_1352,N_36);
or U9379 (N_9379,N_3860,N_1228);
or U9380 (N_9380,N_985,N_147);
nor U9381 (N_9381,N_3466,N_4762);
xor U9382 (N_9382,N_4241,N_4755);
and U9383 (N_9383,N_766,N_2645);
and U9384 (N_9384,N_1819,N_1716);
xor U9385 (N_9385,N_2352,N_979);
nor U9386 (N_9386,N_4229,N_4126);
nand U9387 (N_9387,N_1907,N_4838);
or U9388 (N_9388,N_2045,N_2529);
nor U9389 (N_9389,N_2625,N_1395);
xor U9390 (N_9390,N_2781,N_130);
nand U9391 (N_9391,N_4116,N_1004);
and U9392 (N_9392,N_2447,N_1252);
nand U9393 (N_9393,N_343,N_3262);
or U9394 (N_9394,N_3794,N_4899);
or U9395 (N_9395,N_1525,N_290);
or U9396 (N_9396,N_179,N_4767);
nor U9397 (N_9397,N_2826,N_1992);
and U9398 (N_9398,N_1372,N_4668);
and U9399 (N_9399,N_2339,N_491);
or U9400 (N_9400,N_607,N_1532);
and U9401 (N_9401,N_2582,N_1651);
or U9402 (N_9402,N_3625,N_2256);
nand U9403 (N_9403,N_1449,N_2101);
and U9404 (N_9404,N_1570,N_2887);
or U9405 (N_9405,N_3482,N_3475);
or U9406 (N_9406,N_457,N_760);
nand U9407 (N_9407,N_4068,N_4200);
or U9408 (N_9408,N_189,N_850);
nand U9409 (N_9409,N_4849,N_3074);
xnor U9410 (N_9410,N_2941,N_321);
or U9411 (N_9411,N_1787,N_3148);
or U9412 (N_9412,N_646,N_1648);
nand U9413 (N_9413,N_1264,N_4930);
nor U9414 (N_9414,N_4122,N_737);
nand U9415 (N_9415,N_4085,N_2625);
or U9416 (N_9416,N_3745,N_4873);
nor U9417 (N_9417,N_486,N_3868);
and U9418 (N_9418,N_4122,N_2786);
or U9419 (N_9419,N_3022,N_2710);
nand U9420 (N_9420,N_4649,N_4485);
and U9421 (N_9421,N_1364,N_4527);
or U9422 (N_9422,N_1534,N_4053);
nor U9423 (N_9423,N_4157,N_851);
nor U9424 (N_9424,N_2050,N_1623);
nand U9425 (N_9425,N_651,N_850);
xor U9426 (N_9426,N_2678,N_4708);
nand U9427 (N_9427,N_4791,N_1739);
and U9428 (N_9428,N_4887,N_4118);
and U9429 (N_9429,N_2346,N_3554);
or U9430 (N_9430,N_4483,N_3579);
or U9431 (N_9431,N_3051,N_1188);
or U9432 (N_9432,N_3701,N_4917);
xnor U9433 (N_9433,N_4853,N_1519);
or U9434 (N_9434,N_3635,N_2753);
nand U9435 (N_9435,N_378,N_3336);
and U9436 (N_9436,N_4222,N_237);
xnor U9437 (N_9437,N_3124,N_2293);
and U9438 (N_9438,N_2636,N_4783);
or U9439 (N_9439,N_3520,N_1143);
and U9440 (N_9440,N_4070,N_1264);
and U9441 (N_9441,N_1125,N_4832);
or U9442 (N_9442,N_1265,N_2040);
xnor U9443 (N_9443,N_4025,N_4747);
and U9444 (N_9444,N_657,N_1096);
and U9445 (N_9445,N_1686,N_703);
and U9446 (N_9446,N_2847,N_178);
nand U9447 (N_9447,N_2042,N_4963);
or U9448 (N_9448,N_633,N_3268);
or U9449 (N_9449,N_3422,N_2306);
nor U9450 (N_9450,N_3544,N_2357);
nor U9451 (N_9451,N_1729,N_3204);
or U9452 (N_9452,N_2754,N_4844);
or U9453 (N_9453,N_758,N_3742);
and U9454 (N_9454,N_3455,N_4424);
and U9455 (N_9455,N_3565,N_1850);
nor U9456 (N_9456,N_1348,N_4697);
or U9457 (N_9457,N_2098,N_123);
xor U9458 (N_9458,N_4106,N_4738);
nor U9459 (N_9459,N_1753,N_2157);
nor U9460 (N_9460,N_841,N_4390);
or U9461 (N_9461,N_3743,N_3352);
nor U9462 (N_9462,N_4471,N_1664);
and U9463 (N_9463,N_1819,N_1238);
xor U9464 (N_9464,N_2214,N_4962);
nand U9465 (N_9465,N_3459,N_4148);
xnor U9466 (N_9466,N_1830,N_2555);
and U9467 (N_9467,N_563,N_4874);
xnor U9468 (N_9468,N_4205,N_4923);
and U9469 (N_9469,N_2393,N_4858);
or U9470 (N_9470,N_2336,N_2867);
or U9471 (N_9471,N_3725,N_1400);
nor U9472 (N_9472,N_2178,N_4673);
xnor U9473 (N_9473,N_1274,N_314);
and U9474 (N_9474,N_1763,N_2182);
nand U9475 (N_9475,N_4350,N_3308);
xor U9476 (N_9476,N_3716,N_636);
or U9477 (N_9477,N_3205,N_4109);
or U9478 (N_9478,N_665,N_901);
and U9479 (N_9479,N_2496,N_1841);
or U9480 (N_9480,N_1690,N_2728);
or U9481 (N_9481,N_4689,N_4124);
and U9482 (N_9482,N_1664,N_1778);
xor U9483 (N_9483,N_267,N_1555);
nand U9484 (N_9484,N_1476,N_2124);
nand U9485 (N_9485,N_455,N_3052);
and U9486 (N_9486,N_2255,N_3561);
or U9487 (N_9487,N_2929,N_4975);
or U9488 (N_9488,N_3036,N_199);
nor U9489 (N_9489,N_4835,N_3097);
or U9490 (N_9490,N_2548,N_1671);
xor U9491 (N_9491,N_1668,N_781);
nand U9492 (N_9492,N_4887,N_2368);
xnor U9493 (N_9493,N_3565,N_2004);
and U9494 (N_9494,N_3483,N_4727);
xnor U9495 (N_9495,N_1337,N_4668);
and U9496 (N_9496,N_394,N_2970);
and U9497 (N_9497,N_2764,N_4324);
or U9498 (N_9498,N_3035,N_254);
or U9499 (N_9499,N_3,N_1841);
xor U9500 (N_9500,N_2108,N_4844);
nor U9501 (N_9501,N_1593,N_3451);
nand U9502 (N_9502,N_2769,N_3726);
or U9503 (N_9503,N_763,N_2464);
and U9504 (N_9504,N_2160,N_4350);
nand U9505 (N_9505,N_2740,N_4071);
xnor U9506 (N_9506,N_4140,N_4228);
or U9507 (N_9507,N_3692,N_3393);
nor U9508 (N_9508,N_4308,N_953);
nand U9509 (N_9509,N_3106,N_1599);
nor U9510 (N_9510,N_536,N_4249);
and U9511 (N_9511,N_1976,N_2308);
xnor U9512 (N_9512,N_1840,N_2456);
or U9513 (N_9513,N_3448,N_4725);
nand U9514 (N_9514,N_2383,N_1398);
nor U9515 (N_9515,N_2669,N_1759);
nand U9516 (N_9516,N_2752,N_412);
and U9517 (N_9517,N_780,N_3686);
or U9518 (N_9518,N_3482,N_2902);
nor U9519 (N_9519,N_2360,N_1641);
nor U9520 (N_9520,N_1809,N_2746);
and U9521 (N_9521,N_658,N_2260);
nand U9522 (N_9522,N_2711,N_4913);
nand U9523 (N_9523,N_3529,N_2958);
nand U9524 (N_9524,N_931,N_179);
or U9525 (N_9525,N_1684,N_434);
nand U9526 (N_9526,N_521,N_715);
nand U9527 (N_9527,N_4196,N_4844);
xor U9528 (N_9528,N_4262,N_1416);
and U9529 (N_9529,N_3455,N_3527);
and U9530 (N_9530,N_3916,N_2567);
nor U9531 (N_9531,N_1432,N_619);
xnor U9532 (N_9532,N_3921,N_1220);
xnor U9533 (N_9533,N_89,N_2371);
and U9534 (N_9534,N_1577,N_1178);
nor U9535 (N_9535,N_1283,N_3960);
nand U9536 (N_9536,N_2716,N_934);
nor U9537 (N_9537,N_2108,N_4091);
and U9538 (N_9538,N_4768,N_3951);
and U9539 (N_9539,N_987,N_4483);
nor U9540 (N_9540,N_3237,N_1303);
and U9541 (N_9541,N_1582,N_1346);
nand U9542 (N_9542,N_4158,N_3711);
nand U9543 (N_9543,N_600,N_1223);
nand U9544 (N_9544,N_2326,N_2046);
nand U9545 (N_9545,N_3031,N_1971);
or U9546 (N_9546,N_4754,N_293);
or U9547 (N_9547,N_4993,N_4835);
and U9548 (N_9548,N_2227,N_2602);
nand U9549 (N_9549,N_1769,N_4846);
nand U9550 (N_9550,N_258,N_1830);
nand U9551 (N_9551,N_2039,N_195);
and U9552 (N_9552,N_313,N_2050);
or U9553 (N_9553,N_886,N_3403);
nand U9554 (N_9554,N_515,N_646);
nor U9555 (N_9555,N_977,N_3456);
nand U9556 (N_9556,N_4782,N_2689);
nand U9557 (N_9557,N_3614,N_2270);
or U9558 (N_9558,N_1396,N_3428);
and U9559 (N_9559,N_4477,N_591);
and U9560 (N_9560,N_702,N_3008);
and U9561 (N_9561,N_4634,N_4480);
nand U9562 (N_9562,N_1373,N_1190);
and U9563 (N_9563,N_1335,N_4710);
nand U9564 (N_9564,N_2352,N_273);
or U9565 (N_9565,N_3497,N_3148);
nor U9566 (N_9566,N_4219,N_197);
nor U9567 (N_9567,N_3291,N_4347);
or U9568 (N_9568,N_4341,N_115);
or U9569 (N_9569,N_1221,N_4692);
nor U9570 (N_9570,N_4886,N_4223);
nand U9571 (N_9571,N_3021,N_2508);
nor U9572 (N_9572,N_3891,N_1443);
xor U9573 (N_9573,N_689,N_2162);
nor U9574 (N_9574,N_1863,N_2902);
and U9575 (N_9575,N_249,N_2875);
nor U9576 (N_9576,N_1102,N_709);
or U9577 (N_9577,N_1522,N_3274);
and U9578 (N_9578,N_2574,N_4939);
nor U9579 (N_9579,N_4052,N_1291);
nor U9580 (N_9580,N_3163,N_4832);
and U9581 (N_9581,N_3633,N_1718);
nor U9582 (N_9582,N_2135,N_1562);
nand U9583 (N_9583,N_3117,N_3325);
or U9584 (N_9584,N_4585,N_4816);
and U9585 (N_9585,N_3993,N_44);
nor U9586 (N_9586,N_3083,N_236);
nand U9587 (N_9587,N_4100,N_2063);
nand U9588 (N_9588,N_2033,N_2628);
xor U9589 (N_9589,N_839,N_456);
nand U9590 (N_9590,N_2600,N_1804);
nand U9591 (N_9591,N_738,N_923);
or U9592 (N_9592,N_4017,N_4299);
nand U9593 (N_9593,N_4058,N_3372);
nor U9594 (N_9594,N_4361,N_874);
nand U9595 (N_9595,N_80,N_3542);
nor U9596 (N_9596,N_2870,N_1361);
nand U9597 (N_9597,N_685,N_2780);
and U9598 (N_9598,N_3413,N_4139);
nand U9599 (N_9599,N_149,N_44);
and U9600 (N_9600,N_4349,N_4879);
nor U9601 (N_9601,N_3261,N_1226);
nor U9602 (N_9602,N_4357,N_612);
nor U9603 (N_9603,N_2289,N_3309);
nor U9604 (N_9604,N_4961,N_851);
nor U9605 (N_9605,N_4602,N_1119);
nor U9606 (N_9606,N_2531,N_3327);
nand U9607 (N_9607,N_4020,N_4423);
or U9608 (N_9608,N_1549,N_4144);
or U9609 (N_9609,N_342,N_3758);
nor U9610 (N_9610,N_2538,N_2081);
xor U9611 (N_9611,N_3363,N_810);
or U9612 (N_9612,N_1693,N_2486);
and U9613 (N_9613,N_3708,N_2804);
xnor U9614 (N_9614,N_3422,N_1359);
or U9615 (N_9615,N_3404,N_1519);
nor U9616 (N_9616,N_37,N_2286);
or U9617 (N_9617,N_557,N_3573);
nor U9618 (N_9618,N_1478,N_934);
or U9619 (N_9619,N_3699,N_4583);
nor U9620 (N_9620,N_4135,N_2707);
nand U9621 (N_9621,N_811,N_2448);
nor U9622 (N_9622,N_819,N_4153);
nor U9623 (N_9623,N_563,N_3812);
nor U9624 (N_9624,N_4289,N_4424);
or U9625 (N_9625,N_1811,N_1061);
and U9626 (N_9626,N_3386,N_3621);
and U9627 (N_9627,N_4727,N_2642);
or U9628 (N_9628,N_3240,N_1427);
and U9629 (N_9629,N_2218,N_425);
nand U9630 (N_9630,N_3935,N_2221);
xnor U9631 (N_9631,N_460,N_2521);
xnor U9632 (N_9632,N_2972,N_1291);
or U9633 (N_9633,N_3771,N_1001);
nand U9634 (N_9634,N_3294,N_1656);
and U9635 (N_9635,N_3689,N_1224);
and U9636 (N_9636,N_4435,N_3639);
and U9637 (N_9637,N_825,N_3557);
xor U9638 (N_9638,N_1800,N_2946);
nor U9639 (N_9639,N_3872,N_634);
and U9640 (N_9640,N_4725,N_1892);
and U9641 (N_9641,N_2897,N_3755);
nor U9642 (N_9642,N_981,N_3377);
or U9643 (N_9643,N_4023,N_2988);
and U9644 (N_9644,N_3040,N_1267);
nor U9645 (N_9645,N_434,N_3389);
nor U9646 (N_9646,N_1265,N_1361);
nor U9647 (N_9647,N_917,N_205);
or U9648 (N_9648,N_4841,N_3942);
nor U9649 (N_9649,N_4918,N_1531);
and U9650 (N_9650,N_2465,N_4545);
and U9651 (N_9651,N_1743,N_2014);
and U9652 (N_9652,N_3231,N_2032);
or U9653 (N_9653,N_4324,N_2441);
nor U9654 (N_9654,N_912,N_591);
nand U9655 (N_9655,N_4363,N_1415);
and U9656 (N_9656,N_1485,N_1889);
xor U9657 (N_9657,N_1726,N_4402);
or U9658 (N_9658,N_3007,N_936);
nand U9659 (N_9659,N_4368,N_2348);
nor U9660 (N_9660,N_198,N_2749);
nor U9661 (N_9661,N_3520,N_1434);
nor U9662 (N_9662,N_1467,N_1269);
or U9663 (N_9663,N_3071,N_1426);
or U9664 (N_9664,N_4065,N_3315);
or U9665 (N_9665,N_4205,N_2398);
and U9666 (N_9666,N_3734,N_4670);
nand U9667 (N_9667,N_1862,N_2028);
or U9668 (N_9668,N_4558,N_2702);
nor U9669 (N_9669,N_4247,N_1494);
nand U9670 (N_9670,N_2767,N_1901);
and U9671 (N_9671,N_513,N_4087);
or U9672 (N_9672,N_2608,N_4654);
nor U9673 (N_9673,N_4336,N_1802);
xor U9674 (N_9674,N_1118,N_3682);
and U9675 (N_9675,N_257,N_1392);
xor U9676 (N_9676,N_2837,N_4623);
or U9677 (N_9677,N_3296,N_4300);
nand U9678 (N_9678,N_119,N_2198);
and U9679 (N_9679,N_1430,N_4620);
or U9680 (N_9680,N_1904,N_395);
or U9681 (N_9681,N_4705,N_3807);
nand U9682 (N_9682,N_2706,N_398);
nor U9683 (N_9683,N_384,N_999);
or U9684 (N_9684,N_1641,N_2991);
nand U9685 (N_9685,N_551,N_3354);
and U9686 (N_9686,N_200,N_1408);
and U9687 (N_9687,N_3117,N_1663);
nor U9688 (N_9688,N_3319,N_2432);
nor U9689 (N_9689,N_4416,N_692);
and U9690 (N_9690,N_717,N_1687);
or U9691 (N_9691,N_4051,N_58);
and U9692 (N_9692,N_3035,N_4792);
nand U9693 (N_9693,N_4794,N_2070);
and U9694 (N_9694,N_2675,N_3137);
xor U9695 (N_9695,N_4738,N_2270);
nor U9696 (N_9696,N_3790,N_1648);
or U9697 (N_9697,N_760,N_891);
nand U9698 (N_9698,N_2828,N_4694);
or U9699 (N_9699,N_816,N_906);
nor U9700 (N_9700,N_2905,N_4607);
nand U9701 (N_9701,N_323,N_2464);
and U9702 (N_9702,N_2769,N_2015);
nand U9703 (N_9703,N_4972,N_416);
or U9704 (N_9704,N_1230,N_2326);
nor U9705 (N_9705,N_1055,N_809);
xnor U9706 (N_9706,N_2576,N_3268);
nand U9707 (N_9707,N_1685,N_1669);
or U9708 (N_9708,N_1299,N_4139);
and U9709 (N_9709,N_1970,N_4793);
or U9710 (N_9710,N_3181,N_3833);
nor U9711 (N_9711,N_958,N_2087);
nand U9712 (N_9712,N_4335,N_1685);
nand U9713 (N_9713,N_4144,N_4000);
nor U9714 (N_9714,N_4011,N_3999);
and U9715 (N_9715,N_2812,N_1582);
and U9716 (N_9716,N_517,N_3440);
or U9717 (N_9717,N_4259,N_682);
or U9718 (N_9718,N_3293,N_1059);
nand U9719 (N_9719,N_1006,N_1286);
xnor U9720 (N_9720,N_3284,N_1661);
xor U9721 (N_9721,N_4620,N_2775);
nor U9722 (N_9722,N_816,N_2091);
or U9723 (N_9723,N_2835,N_3121);
nor U9724 (N_9724,N_92,N_804);
nand U9725 (N_9725,N_1265,N_276);
nand U9726 (N_9726,N_3890,N_2366);
or U9727 (N_9727,N_2113,N_1728);
and U9728 (N_9728,N_383,N_3684);
nor U9729 (N_9729,N_2462,N_3836);
and U9730 (N_9730,N_2194,N_2205);
nor U9731 (N_9731,N_2521,N_2216);
nor U9732 (N_9732,N_2585,N_2923);
or U9733 (N_9733,N_2117,N_4639);
or U9734 (N_9734,N_4603,N_2887);
nor U9735 (N_9735,N_4222,N_559);
nor U9736 (N_9736,N_1074,N_2224);
or U9737 (N_9737,N_1001,N_1075);
nand U9738 (N_9738,N_1128,N_2816);
or U9739 (N_9739,N_636,N_3930);
nand U9740 (N_9740,N_3571,N_4888);
nand U9741 (N_9741,N_2476,N_1458);
nor U9742 (N_9742,N_3212,N_2390);
and U9743 (N_9743,N_1414,N_3708);
nand U9744 (N_9744,N_1814,N_2944);
and U9745 (N_9745,N_2349,N_4978);
nor U9746 (N_9746,N_2892,N_3588);
nand U9747 (N_9747,N_2166,N_4678);
xor U9748 (N_9748,N_1985,N_4115);
nor U9749 (N_9749,N_3455,N_434);
xnor U9750 (N_9750,N_2525,N_576);
xnor U9751 (N_9751,N_1129,N_4052);
nor U9752 (N_9752,N_751,N_4111);
and U9753 (N_9753,N_4180,N_3610);
nor U9754 (N_9754,N_2330,N_2655);
and U9755 (N_9755,N_3965,N_2351);
or U9756 (N_9756,N_3964,N_344);
or U9757 (N_9757,N_4021,N_1956);
nand U9758 (N_9758,N_1384,N_4001);
or U9759 (N_9759,N_2268,N_2672);
nor U9760 (N_9760,N_897,N_2289);
and U9761 (N_9761,N_380,N_4162);
or U9762 (N_9762,N_2191,N_873);
nand U9763 (N_9763,N_1105,N_3141);
nand U9764 (N_9764,N_906,N_4862);
nor U9765 (N_9765,N_4060,N_2185);
nor U9766 (N_9766,N_3306,N_3189);
and U9767 (N_9767,N_2034,N_2795);
xor U9768 (N_9768,N_3678,N_1491);
nand U9769 (N_9769,N_2830,N_1322);
and U9770 (N_9770,N_4353,N_1595);
xor U9771 (N_9771,N_1502,N_1850);
or U9772 (N_9772,N_2617,N_1040);
xor U9773 (N_9773,N_1146,N_3048);
nor U9774 (N_9774,N_3846,N_462);
xnor U9775 (N_9775,N_3054,N_362);
and U9776 (N_9776,N_274,N_2130);
or U9777 (N_9777,N_72,N_4507);
nor U9778 (N_9778,N_54,N_4960);
or U9779 (N_9779,N_1481,N_2098);
or U9780 (N_9780,N_4246,N_4624);
and U9781 (N_9781,N_2404,N_2014);
nand U9782 (N_9782,N_547,N_3952);
nand U9783 (N_9783,N_554,N_2122);
and U9784 (N_9784,N_79,N_3766);
xor U9785 (N_9785,N_3218,N_4419);
nor U9786 (N_9786,N_4020,N_1928);
and U9787 (N_9787,N_4824,N_2956);
or U9788 (N_9788,N_52,N_4052);
or U9789 (N_9789,N_4119,N_1878);
xor U9790 (N_9790,N_4314,N_4540);
or U9791 (N_9791,N_693,N_3890);
or U9792 (N_9792,N_457,N_2799);
xnor U9793 (N_9793,N_4335,N_4373);
or U9794 (N_9794,N_2870,N_3501);
or U9795 (N_9795,N_603,N_2640);
nor U9796 (N_9796,N_3941,N_1654);
or U9797 (N_9797,N_3592,N_4907);
nand U9798 (N_9798,N_815,N_2874);
xnor U9799 (N_9799,N_331,N_3702);
nand U9800 (N_9800,N_1009,N_4292);
and U9801 (N_9801,N_3173,N_4902);
or U9802 (N_9802,N_2589,N_642);
or U9803 (N_9803,N_366,N_4957);
nor U9804 (N_9804,N_1836,N_2709);
nor U9805 (N_9805,N_4517,N_3092);
or U9806 (N_9806,N_4839,N_1116);
nand U9807 (N_9807,N_362,N_667);
xor U9808 (N_9808,N_2081,N_3866);
or U9809 (N_9809,N_1432,N_2807);
xnor U9810 (N_9810,N_1550,N_2195);
xor U9811 (N_9811,N_340,N_4032);
and U9812 (N_9812,N_2251,N_3965);
and U9813 (N_9813,N_4672,N_687);
and U9814 (N_9814,N_4003,N_3188);
xnor U9815 (N_9815,N_220,N_2062);
nand U9816 (N_9816,N_4049,N_590);
nor U9817 (N_9817,N_1285,N_1020);
nor U9818 (N_9818,N_552,N_3636);
nor U9819 (N_9819,N_1280,N_125);
nand U9820 (N_9820,N_1675,N_2989);
or U9821 (N_9821,N_3757,N_1716);
and U9822 (N_9822,N_2999,N_2698);
and U9823 (N_9823,N_4950,N_960);
nand U9824 (N_9824,N_1856,N_4351);
nor U9825 (N_9825,N_536,N_2688);
nor U9826 (N_9826,N_3579,N_1486);
nand U9827 (N_9827,N_1162,N_3030);
or U9828 (N_9828,N_801,N_525);
or U9829 (N_9829,N_3759,N_1153);
or U9830 (N_9830,N_2076,N_3229);
and U9831 (N_9831,N_1642,N_4038);
nand U9832 (N_9832,N_2473,N_3588);
and U9833 (N_9833,N_3332,N_311);
nand U9834 (N_9834,N_313,N_3388);
or U9835 (N_9835,N_3990,N_2416);
and U9836 (N_9836,N_2681,N_3435);
nand U9837 (N_9837,N_1006,N_1914);
and U9838 (N_9838,N_3898,N_2081);
or U9839 (N_9839,N_4715,N_4004);
and U9840 (N_9840,N_1954,N_4771);
nand U9841 (N_9841,N_4579,N_4167);
or U9842 (N_9842,N_1281,N_4249);
or U9843 (N_9843,N_861,N_1703);
and U9844 (N_9844,N_4594,N_4631);
xnor U9845 (N_9845,N_2508,N_1881);
or U9846 (N_9846,N_3704,N_1497);
xnor U9847 (N_9847,N_2395,N_4011);
nand U9848 (N_9848,N_783,N_4119);
and U9849 (N_9849,N_4370,N_2218);
nand U9850 (N_9850,N_4683,N_3005);
nor U9851 (N_9851,N_543,N_2920);
and U9852 (N_9852,N_3796,N_3909);
nand U9853 (N_9853,N_4127,N_1693);
nand U9854 (N_9854,N_1151,N_3521);
nor U9855 (N_9855,N_1420,N_604);
nand U9856 (N_9856,N_1025,N_3875);
or U9857 (N_9857,N_4547,N_3910);
nor U9858 (N_9858,N_3314,N_4681);
and U9859 (N_9859,N_4746,N_447);
nor U9860 (N_9860,N_4666,N_500);
nand U9861 (N_9861,N_4567,N_2780);
and U9862 (N_9862,N_911,N_2709);
nor U9863 (N_9863,N_4922,N_4093);
or U9864 (N_9864,N_1391,N_2559);
xnor U9865 (N_9865,N_527,N_995);
xnor U9866 (N_9866,N_4502,N_3486);
or U9867 (N_9867,N_421,N_1754);
nor U9868 (N_9868,N_4215,N_2017);
or U9869 (N_9869,N_454,N_1562);
and U9870 (N_9870,N_593,N_1549);
nor U9871 (N_9871,N_2299,N_1275);
and U9872 (N_9872,N_112,N_3984);
nor U9873 (N_9873,N_2428,N_597);
and U9874 (N_9874,N_1252,N_3767);
nor U9875 (N_9875,N_1868,N_3693);
or U9876 (N_9876,N_1203,N_169);
or U9877 (N_9877,N_342,N_4265);
and U9878 (N_9878,N_4509,N_4335);
nor U9879 (N_9879,N_3534,N_4576);
and U9880 (N_9880,N_827,N_2815);
or U9881 (N_9881,N_1690,N_3416);
nor U9882 (N_9882,N_1263,N_4620);
and U9883 (N_9883,N_2666,N_1893);
nor U9884 (N_9884,N_2996,N_2584);
and U9885 (N_9885,N_1661,N_4909);
nor U9886 (N_9886,N_3799,N_4025);
nand U9887 (N_9887,N_3087,N_4460);
and U9888 (N_9888,N_2037,N_4205);
nand U9889 (N_9889,N_1104,N_1941);
nor U9890 (N_9890,N_3810,N_2834);
and U9891 (N_9891,N_856,N_1160);
nand U9892 (N_9892,N_390,N_4277);
nand U9893 (N_9893,N_4727,N_2157);
nand U9894 (N_9894,N_3049,N_3515);
nor U9895 (N_9895,N_1063,N_728);
nor U9896 (N_9896,N_4869,N_4242);
or U9897 (N_9897,N_903,N_4529);
nand U9898 (N_9898,N_1868,N_1001);
or U9899 (N_9899,N_2363,N_818);
nor U9900 (N_9900,N_1211,N_3471);
or U9901 (N_9901,N_3862,N_645);
or U9902 (N_9902,N_1458,N_3144);
nor U9903 (N_9903,N_4505,N_1092);
and U9904 (N_9904,N_1353,N_547);
nand U9905 (N_9905,N_2869,N_3302);
nand U9906 (N_9906,N_3621,N_1938);
nor U9907 (N_9907,N_4067,N_3790);
nand U9908 (N_9908,N_1410,N_4533);
nor U9909 (N_9909,N_743,N_2175);
and U9910 (N_9910,N_1160,N_632);
nand U9911 (N_9911,N_836,N_2748);
nand U9912 (N_9912,N_1240,N_1520);
nor U9913 (N_9913,N_2027,N_2879);
nor U9914 (N_9914,N_671,N_4087);
nor U9915 (N_9915,N_4542,N_3363);
nor U9916 (N_9916,N_1801,N_195);
nand U9917 (N_9917,N_1027,N_87);
nor U9918 (N_9918,N_1858,N_354);
and U9919 (N_9919,N_1251,N_1052);
nand U9920 (N_9920,N_2614,N_66);
nor U9921 (N_9921,N_533,N_519);
and U9922 (N_9922,N_2812,N_2323);
nand U9923 (N_9923,N_3030,N_1100);
nand U9924 (N_9924,N_2788,N_76);
and U9925 (N_9925,N_3107,N_3293);
nand U9926 (N_9926,N_760,N_4181);
nand U9927 (N_9927,N_2775,N_2075);
nor U9928 (N_9928,N_2291,N_4946);
nor U9929 (N_9929,N_2291,N_1503);
or U9930 (N_9930,N_1794,N_1320);
nand U9931 (N_9931,N_322,N_2950);
or U9932 (N_9932,N_620,N_847);
or U9933 (N_9933,N_3144,N_3955);
or U9934 (N_9934,N_1494,N_1627);
nor U9935 (N_9935,N_732,N_1813);
and U9936 (N_9936,N_1631,N_3213);
xnor U9937 (N_9937,N_4096,N_2355);
nor U9938 (N_9938,N_1627,N_716);
and U9939 (N_9939,N_1893,N_3933);
and U9940 (N_9940,N_2042,N_1874);
nand U9941 (N_9941,N_2185,N_4544);
nand U9942 (N_9942,N_4769,N_4631);
or U9943 (N_9943,N_3435,N_2868);
and U9944 (N_9944,N_4577,N_2635);
and U9945 (N_9945,N_2123,N_3885);
nor U9946 (N_9946,N_1785,N_3468);
nor U9947 (N_9947,N_894,N_4532);
xor U9948 (N_9948,N_1940,N_1762);
or U9949 (N_9949,N_1623,N_3133);
and U9950 (N_9950,N_2580,N_1500);
nor U9951 (N_9951,N_2810,N_3148);
nor U9952 (N_9952,N_801,N_3400);
nand U9953 (N_9953,N_3265,N_172);
and U9954 (N_9954,N_4227,N_1764);
and U9955 (N_9955,N_1032,N_1574);
nand U9956 (N_9956,N_2146,N_361);
or U9957 (N_9957,N_981,N_1999);
and U9958 (N_9958,N_2218,N_845);
nand U9959 (N_9959,N_1204,N_1368);
or U9960 (N_9960,N_3950,N_2465);
nand U9961 (N_9961,N_4876,N_692);
or U9962 (N_9962,N_643,N_4708);
nor U9963 (N_9963,N_4849,N_1181);
or U9964 (N_9964,N_1680,N_1508);
nand U9965 (N_9965,N_1600,N_3356);
nor U9966 (N_9966,N_4050,N_1941);
nor U9967 (N_9967,N_581,N_2792);
or U9968 (N_9968,N_2039,N_3647);
nand U9969 (N_9969,N_2526,N_4123);
and U9970 (N_9970,N_3962,N_4577);
and U9971 (N_9971,N_382,N_4277);
nor U9972 (N_9972,N_4410,N_512);
or U9973 (N_9973,N_3746,N_3851);
nor U9974 (N_9974,N_3173,N_4007);
nand U9975 (N_9975,N_1702,N_2343);
or U9976 (N_9976,N_1511,N_1480);
nor U9977 (N_9977,N_3592,N_2416);
nor U9978 (N_9978,N_964,N_1005);
or U9979 (N_9979,N_4785,N_4816);
nor U9980 (N_9980,N_3793,N_3911);
or U9981 (N_9981,N_2225,N_1489);
or U9982 (N_9982,N_964,N_2505);
nand U9983 (N_9983,N_2007,N_646);
and U9984 (N_9984,N_1044,N_1566);
nand U9985 (N_9985,N_482,N_4495);
nand U9986 (N_9986,N_3954,N_2355);
nand U9987 (N_9987,N_3797,N_4987);
or U9988 (N_9988,N_3296,N_1885);
xor U9989 (N_9989,N_3508,N_2106);
nor U9990 (N_9990,N_3257,N_150);
nor U9991 (N_9991,N_3777,N_2914);
and U9992 (N_9992,N_1382,N_4369);
or U9993 (N_9993,N_4331,N_2024);
nor U9994 (N_9994,N_2903,N_3404);
nand U9995 (N_9995,N_56,N_419);
xor U9996 (N_9996,N_3840,N_276);
or U9997 (N_9997,N_1670,N_2730);
or U9998 (N_9998,N_3157,N_3339);
and U9999 (N_9999,N_544,N_3175);
nor U10000 (N_10000,N_9727,N_9456);
xnor U10001 (N_10001,N_6856,N_5720);
nor U10002 (N_10002,N_6353,N_9846);
nor U10003 (N_10003,N_8151,N_8605);
nor U10004 (N_10004,N_8708,N_9520);
or U10005 (N_10005,N_8138,N_8173);
and U10006 (N_10006,N_7726,N_6022);
nor U10007 (N_10007,N_5005,N_6386);
or U10008 (N_10008,N_5625,N_7647);
nand U10009 (N_10009,N_6109,N_5498);
and U10010 (N_10010,N_6595,N_9207);
and U10011 (N_10011,N_5163,N_8130);
xnor U10012 (N_10012,N_7294,N_9004);
and U10013 (N_10013,N_8457,N_8816);
xor U10014 (N_10014,N_6147,N_9031);
nor U10015 (N_10015,N_5143,N_7886);
and U10016 (N_10016,N_7917,N_9042);
and U10017 (N_10017,N_9548,N_8882);
nand U10018 (N_10018,N_5310,N_8110);
nor U10019 (N_10019,N_8132,N_7575);
and U10020 (N_10020,N_6451,N_5859);
or U10021 (N_10021,N_6062,N_6668);
nor U10022 (N_10022,N_6910,N_7202);
nor U10023 (N_10023,N_5097,N_8383);
nand U10024 (N_10024,N_6343,N_8848);
nor U10025 (N_10025,N_8154,N_9326);
xnor U10026 (N_10026,N_5892,N_9802);
nor U10027 (N_10027,N_6435,N_7203);
nand U10028 (N_10028,N_7687,N_7504);
and U10029 (N_10029,N_7474,N_6963);
or U10030 (N_10030,N_7734,N_8849);
or U10031 (N_10031,N_6696,N_7162);
or U10032 (N_10032,N_8956,N_8612);
nor U10033 (N_10033,N_6646,N_5004);
and U10034 (N_10034,N_6321,N_6145);
nor U10035 (N_10035,N_9881,N_9787);
and U10036 (N_10036,N_5386,N_6490);
nor U10037 (N_10037,N_6962,N_7441);
nor U10038 (N_10038,N_5381,N_5201);
or U10039 (N_10039,N_6123,N_7234);
or U10040 (N_10040,N_5624,N_7088);
nor U10041 (N_10041,N_9280,N_5900);
nand U10042 (N_10042,N_9109,N_9128);
nor U10043 (N_10043,N_5454,N_6291);
nand U10044 (N_10044,N_5278,N_7761);
nor U10045 (N_10045,N_7823,N_9510);
nand U10046 (N_10046,N_7115,N_8021);
and U10047 (N_10047,N_6748,N_6342);
xor U10048 (N_10048,N_5594,N_8720);
nor U10049 (N_10049,N_8675,N_8996);
and U10050 (N_10050,N_9062,N_6400);
nand U10051 (N_10051,N_8325,N_7850);
xor U10052 (N_10052,N_8009,N_7952);
nor U10053 (N_10053,N_5123,N_8390);
xor U10054 (N_10054,N_8868,N_9779);
nand U10055 (N_10055,N_5877,N_7336);
and U10056 (N_10056,N_7978,N_8976);
or U10057 (N_10057,N_7292,N_9001);
nand U10058 (N_10058,N_8087,N_9960);
nand U10059 (N_10059,N_8806,N_7262);
nor U10060 (N_10060,N_7833,N_6607);
or U10061 (N_10061,N_8229,N_8749);
or U10062 (N_10062,N_6102,N_5939);
xnor U10063 (N_10063,N_9474,N_9139);
and U10064 (N_10064,N_7308,N_6887);
and U10065 (N_10065,N_6609,N_8224);
nor U10066 (N_10066,N_5506,N_5880);
or U10067 (N_10067,N_6279,N_9038);
nand U10068 (N_10068,N_5951,N_5073);
xor U10069 (N_10069,N_8760,N_5826);
and U10070 (N_10070,N_6011,N_8198);
nor U10071 (N_10071,N_8845,N_8312);
and U10072 (N_10072,N_8447,N_7724);
xnor U10073 (N_10073,N_6903,N_6048);
nor U10074 (N_10074,N_5179,N_9496);
xor U10075 (N_10075,N_9978,N_5623);
nor U10076 (N_10076,N_5745,N_9718);
nand U10077 (N_10077,N_7072,N_5103);
xor U10078 (N_10078,N_6169,N_9417);
nand U10079 (N_10079,N_7044,N_9805);
or U10080 (N_10080,N_9200,N_5340);
nor U10081 (N_10081,N_9276,N_6705);
xor U10082 (N_10082,N_9756,N_8250);
nand U10083 (N_10083,N_8997,N_8425);
nand U10084 (N_10084,N_5161,N_5964);
nor U10085 (N_10085,N_6805,N_8354);
or U10086 (N_10086,N_9052,N_7869);
and U10087 (N_10087,N_6710,N_5799);
and U10088 (N_10088,N_8435,N_8501);
or U10089 (N_10089,N_5582,N_8431);
or U10090 (N_10090,N_7852,N_6923);
nor U10091 (N_10091,N_5070,N_8945);
or U10092 (N_10092,N_8367,N_9007);
nand U10093 (N_10093,N_7080,N_9986);
and U10094 (N_10094,N_8498,N_5936);
nor U10095 (N_10095,N_5490,N_5879);
nand U10096 (N_10096,N_6175,N_7641);
nand U10097 (N_10097,N_9219,N_7851);
nand U10098 (N_10098,N_7009,N_7168);
or U10099 (N_10099,N_9041,N_8243);
nand U10100 (N_10100,N_6704,N_6822);
or U10101 (N_10101,N_7540,N_9317);
xnor U10102 (N_10102,N_6706,N_9675);
nor U10103 (N_10103,N_5062,N_9695);
or U10104 (N_10104,N_8264,N_8799);
nor U10105 (N_10105,N_9201,N_7493);
nand U10106 (N_10106,N_6876,N_6749);
and U10107 (N_10107,N_7967,N_5831);
nor U10108 (N_10108,N_6171,N_5300);
or U10109 (N_10109,N_5586,N_5916);
and U10110 (N_10110,N_6128,N_5301);
nor U10111 (N_10111,N_9858,N_5296);
or U10112 (N_10112,N_9735,N_5861);
nand U10113 (N_10113,N_8938,N_9610);
nand U10114 (N_10114,N_7274,N_8871);
or U10115 (N_10115,N_5651,N_5178);
and U10116 (N_10116,N_7882,N_7587);
nor U10117 (N_10117,N_6211,N_9240);
xnor U10118 (N_10118,N_9059,N_6701);
and U10119 (N_10119,N_6674,N_8893);
nand U10120 (N_10120,N_9151,N_8558);
nor U10121 (N_10121,N_5711,N_7569);
nor U10122 (N_10122,N_9889,N_8271);
or U10123 (N_10123,N_7145,N_7943);
or U10124 (N_10124,N_6335,N_6208);
nand U10125 (N_10125,N_8106,N_6070);
nor U10126 (N_10126,N_9975,N_8049);
nand U10127 (N_10127,N_9566,N_8208);
and U10128 (N_10128,N_6469,N_7327);
or U10129 (N_10129,N_5653,N_6257);
nand U10130 (N_10130,N_8793,N_6232);
and U10131 (N_10131,N_7206,N_9601);
nor U10132 (N_10132,N_8278,N_5121);
or U10133 (N_10133,N_9776,N_5126);
nand U10134 (N_10134,N_6076,N_9751);
or U10135 (N_10135,N_9167,N_9183);
nand U10136 (N_10136,N_6454,N_8571);
or U10137 (N_10137,N_8112,N_6734);
and U10138 (N_10138,N_9034,N_9998);
nand U10139 (N_10139,N_9150,N_7856);
or U10140 (N_10140,N_5215,N_8769);
nand U10141 (N_10141,N_9341,N_6301);
and U10142 (N_10142,N_6154,N_9110);
and U10143 (N_10143,N_7273,N_9574);
or U10144 (N_10144,N_6543,N_6085);
nand U10145 (N_10145,N_7400,N_6954);
and U10146 (N_10146,N_5714,N_5687);
nor U10147 (N_10147,N_7176,N_7134);
nand U10148 (N_10148,N_9364,N_8966);
nor U10149 (N_10149,N_6014,N_5489);
or U10150 (N_10150,N_6453,N_7981);
and U10151 (N_10151,N_6026,N_6883);
or U10152 (N_10152,N_6336,N_6006);
nor U10153 (N_10153,N_8975,N_5503);
and U10154 (N_10154,N_6639,N_6266);
nand U10155 (N_10155,N_7874,N_9943);
and U10156 (N_10156,N_9852,N_6645);
nand U10157 (N_10157,N_5098,N_8531);
and U10158 (N_10158,N_6666,N_9782);
or U10159 (N_10159,N_9262,N_9270);
nor U10160 (N_10160,N_6605,N_5652);
and U10161 (N_10161,N_5117,N_5459);
nand U10162 (N_10162,N_8702,N_7713);
nor U10163 (N_10163,N_8485,N_8314);
xor U10164 (N_10164,N_7759,N_8929);
and U10165 (N_10165,N_6261,N_6957);
xnor U10166 (N_10166,N_7419,N_8281);
nand U10167 (N_10167,N_9656,N_9467);
xor U10168 (N_10168,N_5311,N_6806);
and U10169 (N_10169,N_6796,N_7577);
nand U10170 (N_10170,N_5365,N_7029);
nor U10171 (N_10171,N_8574,N_6235);
and U10172 (N_10172,N_7602,N_5344);
nor U10173 (N_10173,N_8023,N_8445);
and U10174 (N_10174,N_9106,N_9265);
nand U10175 (N_10175,N_8292,N_5703);
nand U10176 (N_10176,N_5313,N_9550);
nand U10177 (N_10177,N_8918,N_5085);
nor U10178 (N_10178,N_8458,N_6206);
or U10179 (N_10179,N_8861,N_8565);
or U10180 (N_10180,N_9230,N_9893);
nand U10181 (N_10181,N_5578,N_5061);
and U10182 (N_10182,N_6551,N_6745);
and U10183 (N_10183,N_6428,N_6873);
nor U10184 (N_10184,N_7220,N_5698);
and U10185 (N_10185,N_6452,N_6479);
and U10186 (N_10186,N_9382,N_7824);
or U10187 (N_10187,N_6729,N_6383);
nor U10188 (N_10188,N_5959,N_8274);
or U10189 (N_10189,N_7762,N_5554);
and U10190 (N_10190,N_8785,N_8873);
nor U10191 (N_10191,N_8895,N_7857);
nand U10192 (N_10192,N_7418,N_5522);
nor U10193 (N_10193,N_9728,N_8905);
nand U10194 (N_10194,N_5003,N_6731);
nor U10195 (N_10195,N_5999,N_7460);
nand U10196 (N_10196,N_8294,N_5963);
or U10197 (N_10197,N_8883,N_7486);
xor U10198 (N_10198,N_9285,N_6000);
nand U10199 (N_10199,N_8872,N_8640);
nand U10200 (N_10200,N_7076,N_6976);
or U10201 (N_10201,N_9238,N_8419);
or U10202 (N_10202,N_7579,N_8520);
and U10203 (N_10203,N_8546,N_9775);
xnor U10204 (N_10204,N_7456,N_5280);
nand U10205 (N_10205,N_8624,N_7298);
xor U10206 (N_10206,N_5952,N_6449);
nor U10207 (N_10207,N_7254,N_5142);
and U10208 (N_10208,N_7370,N_6567);
or U10209 (N_10209,N_9416,N_5518);
xor U10210 (N_10210,N_5596,N_5798);
or U10211 (N_10211,N_8363,N_6462);
nand U10212 (N_10212,N_7074,N_6699);
and U10213 (N_10213,N_6135,N_7470);
nor U10214 (N_10214,N_5835,N_7958);
or U10215 (N_10215,N_6267,N_9414);
xnor U10216 (N_10216,N_7702,N_9153);
nor U10217 (N_10217,N_7535,N_8006);
xor U10218 (N_10218,N_5746,N_9103);
and U10219 (N_10219,N_5707,N_8045);
or U10220 (N_10220,N_8638,N_5661);
xnor U10221 (N_10221,N_7838,N_7281);
and U10222 (N_10222,N_9259,N_7064);
nor U10223 (N_10223,N_6970,N_7496);
nor U10224 (N_10224,N_6925,N_8223);
nand U10225 (N_10225,N_9247,N_7223);
and U10226 (N_10226,N_5740,N_8747);
or U10227 (N_10227,N_7306,N_7123);
and U10228 (N_10228,N_9147,N_9901);
and U10229 (N_10229,N_9622,N_7586);
or U10230 (N_10230,N_9730,N_7159);
or U10231 (N_10231,N_5497,N_8575);
nor U10232 (N_10232,N_6759,N_7037);
or U10233 (N_10233,N_8300,N_8542);
nor U10234 (N_10234,N_5620,N_8832);
nand U10235 (N_10235,N_9292,N_7240);
or U10236 (N_10236,N_7478,N_8601);
and U10237 (N_10237,N_8668,N_9168);
and U10238 (N_10238,N_8682,N_7337);
or U10239 (N_10239,N_7790,N_8762);
nand U10240 (N_10240,N_8074,N_7097);
nor U10241 (N_10241,N_5317,N_5241);
nand U10242 (N_10242,N_5760,N_6634);
and U10243 (N_10243,N_8742,N_6861);
nor U10244 (N_10244,N_6496,N_7127);
and U10245 (N_10245,N_8954,N_6224);
xor U10246 (N_10246,N_5332,N_9919);
and U10247 (N_10247,N_9921,N_6590);
or U10248 (N_10248,N_9323,N_7816);
nor U10249 (N_10249,N_7841,N_6942);
xnor U10250 (N_10250,N_9941,N_7356);
and U10251 (N_10251,N_6139,N_6108);
nand U10252 (N_10252,N_9969,N_9729);
and U10253 (N_10253,N_7495,N_8101);
nand U10254 (N_10254,N_6849,N_7099);
and U10255 (N_10255,N_8355,N_6306);
xor U10256 (N_10256,N_7484,N_7126);
nor U10257 (N_10257,N_9376,N_7949);
nor U10258 (N_10258,N_6867,N_7572);
and U10259 (N_10259,N_8568,N_6010);
or U10260 (N_10260,N_7578,N_9555);
nand U10261 (N_10261,N_7238,N_6637);
or U10262 (N_10262,N_9545,N_8672);
nand U10263 (N_10263,N_8261,N_8228);
or U10264 (N_10264,N_9268,N_5791);
nor U10265 (N_10265,N_9928,N_7321);
or U10266 (N_10266,N_5523,N_5309);
and U10267 (N_10267,N_6176,N_7897);
and U10268 (N_10268,N_5286,N_5854);
nand U10269 (N_10269,N_9359,N_6052);
and U10270 (N_10270,N_8662,N_6756);
nor U10271 (N_10271,N_9436,N_9434);
and U10272 (N_10272,N_9489,N_5391);
or U10273 (N_10273,N_6036,N_6236);
or U10274 (N_10274,N_7196,N_7753);
xnor U10275 (N_10275,N_7883,N_6552);
nor U10276 (N_10276,N_7564,N_9632);
and U10277 (N_10277,N_7335,N_6544);
and U10278 (N_10278,N_6524,N_9018);
nor U10279 (N_10279,N_8296,N_9012);
or U10280 (N_10280,N_5750,N_6845);
nor U10281 (N_10281,N_7342,N_7073);
nor U10282 (N_10282,N_9029,N_5823);
xnor U10283 (N_10283,N_7230,N_5992);
nor U10284 (N_10284,N_9408,N_8540);
nand U10285 (N_10285,N_5853,N_5084);
xor U10286 (N_10286,N_6960,N_8851);
nor U10287 (N_10287,N_8986,N_6564);
and U10288 (N_10288,N_7678,N_9182);
or U10289 (N_10289,N_9249,N_7039);
nor U10290 (N_10290,N_5099,N_5864);
xnor U10291 (N_10291,N_8761,N_6278);
or U10292 (N_10292,N_9892,N_6127);
xor U10293 (N_10293,N_9469,N_9596);
nor U10294 (N_10294,N_9391,N_9942);
nor U10295 (N_10295,N_9372,N_9816);
or U10296 (N_10296,N_6142,N_6602);
nand U10297 (N_10297,N_7027,N_9711);
nand U10298 (N_10298,N_7170,N_9304);
or U10299 (N_10299,N_6791,N_8239);
and U10300 (N_10300,N_9066,N_7235);
nand U10301 (N_10301,N_5599,N_9368);
and U10302 (N_10302,N_8071,N_8468);
and U10303 (N_10303,N_7032,N_6376);
and U10304 (N_10304,N_5326,N_8187);
or U10305 (N_10305,N_6906,N_9768);
or U10306 (N_10306,N_8920,N_7588);
nand U10307 (N_10307,N_5800,N_7275);
and U10308 (N_10308,N_5060,N_8414);
and U10309 (N_10309,N_7511,N_8024);
nor U10310 (N_10310,N_8470,N_9169);
nor U10311 (N_10311,N_9360,N_8897);
nand U10312 (N_10312,N_7889,N_9646);
nor U10313 (N_10313,N_6156,N_7807);
nand U10314 (N_10314,N_7314,N_8989);
and U10315 (N_10315,N_5270,N_7006);
or U10316 (N_10316,N_7545,N_5415);
nand U10317 (N_10317,N_5355,N_7430);
and U10318 (N_10318,N_6684,N_5263);
nor U10319 (N_10319,N_9196,N_9314);
nand U10320 (N_10320,N_6021,N_5485);
xor U10321 (N_10321,N_6083,N_7218);
or U10322 (N_10322,N_8040,N_9203);
nand U10323 (N_10323,N_8356,N_7876);
xor U10324 (N_10324,N_6017,N_8763);
nand U10325 (N_10325,N_8788,N_6272);
nand U10326 (N_10326,N_8674,N_8155);
or U10327 (N_10327,N_8225,N_5588);
or U10328 (N_10328,N_6019,N_6095);
nor U10329 (N_10329,N_7835,N_7596);
and U10330 (N_10330,N_6725,N_5010);
nand U10331 (N_10331,N_8273,N_6831);
xnor U10332 (N_10332,N_8634,N_8691);
nor U10333 (N_10333,N_6928,N_6106);
and U10334 (N_10334,N_6559,N_6242);
or U10335 (N_10335,N_7182,N_6364);
nor U10336 (N_10336,N_8705,N_6506);
nor U10337 (N_10337,N_7503,N_9322);
nor U10338 (N_10338,N_9965,N_7185);
nor U10339 (N_10339,N_8766,N_9275);
nand U10340 (N_10340,N_9309,N_5185);
or U10341 (N_10341,N_6565,N_8734);
and U10342 (N_10342,N_9984,N_8815);
or U10343 (N_10343,N_6866,N_7506);
and U10344 (N_10344,N_6483,N_5150);
nor U10345 (N_10345,N_6892,N_5530);
nand U10346 (N_10346,N_6037,N_8140);
nor U10347 (N_10347,N_5100,N_9896);
nor U10348 (N_10348,N_5922,N_7873);
nor U10349 (N_10349,N_6061,N_7911);
or U10350 (N_10350,N_7737,N_8898);
nor U10351 (N_10351,N_6986,N_7174);
and U10352 (N_10352,N_5763,N_7605);
and U10353 (N_10353,N_8245,N_8283);
xor U10354 (N_10354,N_5133,N_7390);
nand U10355 (N_10355,N_5040,N_8860);
nor U10356 (N_10356,N_8592,N_7243);
or U10357 (N_10357,N_6297,N_6445);
nand U10358 (N_10358,N_8216,N_6541);
nor U10359 (N_10359,N_9696,N_5574);
and U10360 (N_10360,N_8259,N_7249);
and U10361 (N_10361,N_9698,N_8660);
and U10362 (N_10362,N_5896,N_7936);
and U10363 (N_10363,N_7854,N_6038);
and U10364 (N_10364,N_9152,N_8538);
nand U10365 (N_10365,N_6440,N_5167);
and U10366 (N_10366,N_5205,N_7119);
nand U10367 (N_10367,N_6471,N_7760);
and U10368 (N_10368,N_9124,N_7973);
and U10369 (N_10369,N_7861,N_6687);
nor U10370 (N_10370,N_6511,N_9022);
and U10371 (N_10371,N_9594,N_7532);
or U10372 (N_10372,N_5820,N_8203);
nand U10373 (N_10373,N_8964,N_9184);
and U10374 (N_10374,N_6498,N_5604);
nor U10375 (N_10375,N_7423,N_9180);
nand U10376 (N_10376,N_8331,N_6217);
and U10377 (N_10377,N_8569,N_8548);
nand U10378 (N_10378,N_5954,N_7698);
nor U10379 (N_10379,N_7515,N_7160);
or U10380 (N_10380,N_9880,N_9754);
and U10381 (N_10381,N_8948,N_7498);
or U10382 (N_10382,N_9466,N_7646);
or U10383 (N_10383,N_6254,N_5284);
nor U10384 (N_10384,N_9424,N_5375);
nand U10385 (N_10385,N_8089,N_7584);
nor U10386 (N_10386,N_6537,N_8376);
nor U10387 (N_10387,N_7132,N_6884);
nor U10388 (N_10388,N_6346,N_5684);
nand U10389 (N_10389,N_7693,N_6165);
and U10390 (N_10390,N_7431,N_8516);
nand U10391 (N_10391,N_9983,N_9624);
and U10392 (N_10392,N_5742,N_6041);
nand U10393 (N_10393,N_8344,N_9949);
or U10394 (N_10394,N_6717,N_6079);
and U10395 (N_10395,N_5568,N_9017);
and U10396 (N_10396,N_9433,N_9840);
nand U10397 (N_10397,N_5719,N_7694);
and U10398 (N_10398,N_6895,N_5514);
nor U10399 (N_10399,N_8545,N_9597);
and U10400 (N_10400,N_5507,N_7962);
nand U10401 (N_10401,N_9287,N_5079);
nor U10402 (N_10402,N_9166,N_6881);
and U10403 (N_10403,N_8577,N_5076);
and U10404 (N_10404,N_7058,N_6111);
nor U10405 (N_10405,N_8163,N_9327);
xnor U10406 (N_10406,N_8267,N_5676);
and U10407 (N_10407,N_6130,N_5700);
xor U10408 (N_10408,N_6509,N_5156);
and U10409 (N_10409,N_9218,N_8126);
xnor U10410 (N_10410,N_8553,N_9536);
nand U10411 (N_10411,N_8329,N_7165);
or U10412 (N_10412,N_5119,N_6081);
or U10413 (N_10413,N_7556,N_5109);
or U10414 (N_10414,N_9916,N_9120);
nor U10415 (N_10415,N_5524,N_7499);
or U10416 (N_10416,N_6458,N_6007);
nand U10417 (N_10417,N_7214,N_9388);
nand U10418 (N_10418,N_9811,N_8217);
and U10419 (N_10419,N_6003,N_6890);
nand U10420 (N_10420,N_7517,N_9927);
and U10421 (N_10421,N_7628,N_7591);
xor U10422 (N_10422,N_9819,N_6616);
xor U10423 (N_10423,N_9633,N_9158);
nor U10424 (N_10424,N_6988,N_7666);
xor U10425 (N_10425,N_9641,N_9366);
or U10426 (N_10426,N_9873,N_9838);
or U10427 (N_10427,N_8035,N_5790);
nor U10428 (N_10428,N_5370,N_9707);
nand U10429 (N_10429,N_9132,N_9692);
or U10430 (N_10430,N_5267,N_6276);
xnor U10431 (N_10431,N_7339,N_7771);
or U10432 (N_10432,N_6885,N_5087);
nand U10433 (N_10433,N_7297,N_8387);
nor U10434 (N_10434,N_8215,N_5536);
or U10435 (N_10435,N_7283,N_6456);
xor U10436 (N_10436,N_6525,N_6514);
or U10437 (N_10437,N_9407,N_6655);
or U10438 (N_10438,N_6055,N_9485);
or U10439 (N_10439,N_6878,N_8384);
nor U10440 (N_10440,N_5632,N_7410);
or U10441 (N_10441,N_6025,N_5670);
nor U10442 (N_10442,N_9334,N_5449);
nor U10443 (N_10443,N_5838,N_8725);
and U10444 (N_10444,N_5047,N_5140);
nor U10445 (N_10445,N_7960,N_7963);
nand U10446 (N_10446,N_7216,N_5909);
nor U10447 (N_10447,N_8263,N_6863);
nand U10448 (N_10448,N_7386,N_7346);
nand U10449 (N_10449,N_6797,N_8654);
or U10450 (N_10450,N_8805,N_7795);
and U10451 (N_10451,N_6122,N_8214);
nor U10452 (N_10452,N_6329,N_5890);
nand U10453 (N_10453,N_8098,N_5442);
xor U10454 (N_10454,N_7828,N_8491);
and U10455 (N_10455,N_9300,N_9278);
or U10456 (N_10456,N_6377,N_7246);
and U10457 (N_10457,N_9325,N_6819);
nand U10458 (N_10458,N_8235,N_8181);
nand U10459 (N_10459,N_9712,N_9387);
xnor U10460 (N_10460,N_5072,N_7043);
and U10461 (N_10461,N_5945,N_9908);
nor U10462 (N_10462,N_9529,N_6094);
xnor U10463 (N_10463,N_9856,N_5077);
nand U10464 (N_10464,N_6961,N_8679);
and U10465 (N_10465,N_7451,N_8656);
or U10466 (N_10466,N_9934,N_6898);
nand U10467 (N_10467,N_7231,N_9912);
nor U10468 (N_10468,N_9784,N_7950);
nor U10469 (N_10469,N_5553,N_9229);
xnor U10470 (N_10470,N_9206,N_9330);
nand U10471 (N_10471,N_5755,N_7580);
nor U10472 (N_10472,N_6653,N_8099);
nand U10473 (N_10473,N_8527,N_5775);
xnor U10474 (N_10474,N_5701,N_9263);
nor U10475 (N_10475,N_5222,N_6947);
nand U10476 (N_10476,N_5146,N_7658);
xor U10477 (N_10477,N_7065,N_5028);
nand U10478 (N_10478,N_6741,N_9758);
nor U10479 (N_10479,N_6966,N_9140);
nand U10480 (N_10480,N_7796,N_9410);
or U10481 (N_10481,N_5034,N_5783);
or U10482 (N_10482,N_7059,N_5247);
and U10483 (N_10483,N_7625,N_9046);
or U10484 (N_10484,N_6042,N_9740);
nor U10485 (N_10485,N_9484,N_5086);
or U10486 (N_10486,N_6173,N_9188);
nor U10487 (N_10487,N_9832,N_7681);
and U10488 (N_10488,N_8960,N_9839);
nor U10489 (N_10489,N_6218,N_8765);
nor U10490 (N_10490,N_6584,N_8276);
xnor U10491 (N_10491,N_7383,N_6628);
nand U10492 (N_10492,N_9264,N_9156);
nand U10493 (N_10493,N_8870,N_7002);
or U10494 (N_10494,N_7905,N_9697);
nand U10495 (N_10495,N_7371,N_5390);
or U10496 (N_10496,N_8505,N_7539);
and U10497 (N_10497,N_6210,N_6691);
and U10498 (N_10498,N_7514,N_7933);
nor U10499 (N_10499,N_6040,N_8051);
nand U10500 (N_10500,N_5232,N_8330);
and U10501 (N_10501,N_5525,N_9352);
nor U10502 (N_10502,N_8703,N_6913);
and U10503 (N_10503,N_5682,N_9035);
nand U10504 (N_10504,N_7751,N_6916);
and U10505 (N_10505,N_9405,N_6434);
nor U10506 (N_10506,N_8484,N_9232);
and U10507 (N_10507,N_7806,N_7426);
nand U10508 (N_10508,N_6592,N_5323);
or U10509 (N_10509,N_7643,N_5373);
xnor U10510 (N_10510,N_5056,N_6613);
nor U10511 (N_10511,N_7750,N_5812);
nor U10512 (N_10512,N_5333,N_7974);
or U10513 (N_10513,N_6922,N_5195);
or U10514 (N_10514,N_9195,N_5515);
or U10515 (N_10515,N_5316,N_7060);
and U10516 (N_10516,N_8737,N_7604);
nor U10517 (N_10517,N_9621,N_9260);
and U10518 (N_10518,N_8333,N_7593);
and U10519 (N_10519,N_5276,N_5006);
nand U10520 (N_10520,N_7502,N_6547);
nor U10521 (N_10521,N_8533,N_9592);
nand U10522 (N_10522,N_5942,N_8518);
nor U10523 (N_10523,N_5226,N_5902);
nand U10524 (N_10524,N_6415,N_6110);
nand U10525 (N_10525,N_5932,N_7045);
or U10526 (N_10526,N_6358,N_8910);
nand U10527 (N_10527,N_7033,N_6854);
nand U10528 (N_10528,N_8752,N_7287);
or U10529 (N_10529,N_5279,N_8979);
and U10530 (N_10530,N_9884,N_8562);
xor U10531 (N_10531,N_5731,N_7420);
xnor U10532 (N_10532,N_9910,N_6665);
and U10533 (N_10533,N_5000,N_8921);
and U10534 (N_10534,N_6308,N_9674);
xor U10535 (N_10535,N_5581,N_6880);
nor U10536 (N_10536,N_8730,N_5184);
nor U10537 (N_10537,N_6669,N_9453);
xnor U10538 (N_10538,N_8395,N_8196);
nor U10539 (N_10539,N_6065,N_9149);
xor U10540 (N_10540,N_7524,N_9159);
nor U10541 (N_10541,N_6812,N_7928);
and U10542 (N_10542,N_8421,N_5631);
xor U10543 (N_10543,N_5403,N_7815);
and U10544 (N_10544,N_6814,N_5855);
nor U10545 (N_10545,N_6656,N_8459);
or U10546 (N_10546,N_8886,N_5659);
and U10547 (N_10547,N_6050,N_5752);
xnor U10548 (N_10548,N_9048,N_8370);
nor U10549 (N_10549,N_5175,N_9138);
nor U10550 (N_10550,N_8687,N_9464);
and U10551 (N_10551,N_9398,N_7573);
nor U10552 (N_10552,N_6658,N_5532);
nand U10553 (N_10553,N_9186,N_5400);
and U10554 (N_10554,N_5242,N_6535);
and U10555 (N_10555,N_5621,N_5245);
or U10556 (N_10556,N_8404,N_8326);
and U10557 (N_10557,N_9720,N_7599);
nand U10558 (N_10558,N_8050,N_7408);
nor U10559 (N_10559,N_5235,N_9631);
and U10560 (N_10560,N_7369,N_8590);
nand U10561 (N_10561,N_7541,N_7161);
and U10562 (N_10562,N_9807,N_5686);
and U10563 (N_10563,N_5937,N_7725);
nor U10564 (N_10564,N_8256,N_7712);
nand U10565 (N_10565,N_9305,N_9693);
or U10566 (N_10566,N_6993,N_5776);
and U10567 (N_10567,N_7270,N_8022);
nand U10568 (N_10568,N_6493,N_5974);
nand U10569 (N_10569,N_6926,N_5730);
or U10570 (N_10570,N_7895,N_5152);
xor U10571 (N_10571,N_6968,N_8809);
nand U10572 (N_10572,N_8136,N_8949);
nor U10573 (N_10573,N_5063,N_6736);
or U10574 (N_10574,N_5642,N_9385);
and U10575 (N_10575,N_7697,N_6792);
xor U10576 (N_10576,N_9972,N_8563);
or U10577 (N_10577,N_9743,N_6461);
nand U10578 (N_10578,N_8014,N_8507);
or U10579 (N_10579,N_9664,N_8567);
nor U10580 (N_10580,N_5948,N_8836);
nand U10581 (N_10581,N_7862,N_6443);
nor U10582 (N_10582,N_8128,N_7067);
nand U10583 (N_10583,N_7334,N_6004);
xnor U10584 (N_10584,N_8664,N_9241);
nand U10585 (N_10585,N_8364,N_9449);
nand U10586 (N_10586,N_9461,N_9008);
or U10587 (N_10587,N_8255,N_7312);
nor U10588 (N_10588,N_6549,N_9216);
nand U10589 (N_10589,N_5264,N_8145);
and U10590 (N_10590,N_7610,N_5451);
and U10591 (N_10591,N_8443,N_7379);
or U10592 (N_10592,N_6783,N_5327);
xnor U10593 (N_10593,N_7849,N_6527);
nor U10594 (N_10594,N_6804,N_9377);
or U10595 (N_10595,N_7241,N_6894);
nand U10596 (N_10596,N_5261,N_7972);
nand U10597 (N_10597,N_7295,N_8653);
nand U10598 (N_10598,N_6188,N_7380);
nand U10599 (N_10599,N_7347,N_8880);
or U10600 (N_10600,N_8811,N_6871);
nor U10601 (N_10601,N_8651,N_6522);
nand U10602 (N_10602,N_5105,N_5848);
xnor U10603 (N_10603,N_9797,N_9825);
or U10604 (N_10604,N_6994,N_6582);
or U10605 (N_10605,N_7146,N_9459);
and U10606 (N_10606,N_8598,N_5425);
or U10607 (N_10607,N_6585,N_5811);
nor U10608 (N_10608,N_5706,N_6432);
xor U10609 (N_10609,N_6572,N_7859);
xnor U10610 (N_10610,N_9131,N_6816);
nor U10611 (N_10611,N_7887,N_5899);
or U10612 (N_10612,N_9723,N_8896);
or U10613 (N_10613,N_9888,N_8671);
and U10614 (N_10614,N_6712,N_9676);
nand U10615 (N_10615,N_5124,N_6889);
nand U10616 (N_10616,N_6781,N_7105);
and U10617 (N_10617,N_9468,N_7909);
nand U10618 (N_10618,N_6588,N_9311);
and U10619 (N_10619,N_7880,N_7330);
nor U10620 (N_10620,N_8814,N_6626);
or U10621 (N_10621,N_9477,N_6760);
nand U10622 (N_10622,N_6893,N_6072);
nand U10623 (N_10623,N_7867,N_6991);
xor U10624 (N_10624,N_6395,N_6793);
or U10625 (N_10625,N_8504,N_5411);
nand U10626 (N_10626,N_8923,N_9506);
nand U10627 (N_10627,N_9640,N_7497);
nor U10628 (N_10628,N_8299,N_7332);
and U10629 (N_10629,N_8125,N_9629);
and U10630 (N_10630,N_7147,N_7232);
nor U10631 (N_10631,N_7018,N_7233);
nand U10632 (N_10632,N_9878,N_9465);
or U10633 (N_10633,N_5627,N_8655);
or U10634 (N_10634,N_6396,N_6480);
and U10635 (N_10635,N_8750,N_6846);
nand U10636 (N_10636,N_7141,N_8095);
nand U10637 (N_10637,N_8134,N_7583);
or U10638 (N_10638,N_7530,N_8974);
xnor U10639 (N_10639,N_9613,N_7565);
xnor U10640 (N_10640,N_7138,N_5101);
xnor U10641 (N_10641,N_6502,N_9088);
and U10642 (N_10642,N_7075,N_5444);
nand U10643 (N_10643,N_8442,N_8047);
nor U10644 (N_10644,N_7742,N_9423);
or U10645 (N_10645,N_6251,N_5722);
nor U10646 (N_10646,N_7208,N_5850);
nand U10647 (N_10647,N_7717,N_5697);
nor U10648 (N_10648,N_7582,N_6350);
and U10649 (N_10649,N_6505,N_9689);
nand U10650 (N_10650,N_8988,N_9899);
nand U10651 (N_10651,N_6788,N_7839);
nand U10652 (N_10652,N_5944,N_7597);
nand U10653 (N_10653,N_5510,N_9905);
or U10654 (N_10654,N_6911,N_8609);
or U10655 (N_10655,N_5325,N_5176);
and U10656 (N_10656,N_5765,N_7526);
or U10657 (N_10657,N_8578,N_7549);
nand U10658 (N_10658,N_6870,N_5867);
nand U10659 (N_10659,N_5387,N_5299);
nor U10660 (N_10660,N_6651,N_5735);
nand U10661 (N_10661,N_6627,N_6990);
nor U10662 (N_10662,N_9144,N_7527);
or U10663 (N_10663,N_7038,N_6391);
nand U10664 (N_10664,N_6345,N_5772);
and U10665 (N_10665,N_8347,N_9722);
nand U10666 (N_10666,N_7285,N_6977);
nand U10667 (N_10667,N_6753,N_7925);
or U10668 (N_10668,N_9853,N_7756);
xor U10669 (N_10669,N_7617,N_6492);
and U10670 (N_10670,N_6408,N_9071);
xnor U10671 (N_10671,N_8557,N_8581);
nand U10672 (N_10672,N_5273,N_9806);
or U10673 (N_10673,N_8328,N_6802);
and U10674 (N_10674,N_8402,N_7931);
nand U10675 (N_10675,N_5757,N_7155);
or U10676 (N_10676,N_8764,N_9988);
and U10677 (N_10677,N_6374,N_5359);
or U10678 (N_10678,N_7663,N_6548);
or U10679 (N_10679,N_9721,N_5508);
and U10680 (N_10680,N_9021,N_9137);
nand U10681 (N_10681,N_8361,N_7427);
and U10682 (N_10682,N_8603,N_6028);
nor U10683 (N_10683,N_9061,N_6937);
and U10684 (N_10684,N_7103,N_7810);
or U10685 (N_10685,N_5956,N_6930);
xor U10686 (N_10686,N_9361,N_8617);
and U10687 (N_10687,N_7091,N_7505);
nand U10688 (N_10688,N_9991,N_5913);
and U10689 (N_10689,N_9836,N_7660);
nand U10690 (N_10690,N_5452,N_7153);
nor U10691 (N_10691,N_6093,N_5605);
nor U10692 (N_10692,N_8589,N_7843);
and U10693 (N_10693,N_6641,N_7108);
or U10694 (N_10694,N_9024,N_5845);
nor U10695 (N_10695,N_7429,N_8768);
nand U10696 (N_10696,N_7868,N_8962);
nand U10697 (N_10697,N_7461,N_7634);
nor U10698 (N_10698,N_7636,N_8607);
nor U10699 (N_10699,N_7537,N_9190);
xnor U10700 (N_10700,N_8279,N_6409);
or U10701 (N_10701,N_9231,N_8194);
nor U10702 (N_10702,N_5792,N_8062);
and U10703 (N_10703,N_9279,N_7227);
and U10704 (N_10704,N_9351,N_9559);
nor U10705 (N_10705,N_6596,N_5940);
or U10706 (N_10706,N_8282,N_5438);
or U10707 (N_10707,N_5493,N_5288);
and U10708 (N_10708,N_9296,N_9576);
nand U10709 (N_10709,N_6611,N_7344);
and U10710 (N_10710,N_6694,N_8791);
or U10711 (N_10711,N_5015,N_7436);
nand U10712 (N_10712,N_8091,N_7078);
or U10713 (N_10713,N_8184,N_7585);
xor U10714 (N_10714,N_9123,N_6231);
nand U10715 (N_10715,N_6836,N_6832);
xor U10716 (N_10716,N_9673,N_7326);
or U10717 (N_10717,N_9223,N_7831);
or U10718 (N_10718,N_6470,N_9302);
and U10719 (N_10719,N_8179,N_7005);
xor U10720 (N_10720,N_8736,N_7749);
nand U10721 (N_10721,N_5960,N_5613);
or U10722 (N_10722,N_6478,N_7789);
nor U10723 (N_10723,N_6546,N_9487);
nand U10724 (N_10724,N_8758,N_6398);
nor U10725 (N_10725,N_6735,N_6333);
nor U10726 (N_10726,N_8461,N_8639);
nand U10727 (N_10727,N_9141,N_5437);
nor U10728 (N_10728,N_5095,N_5663);
or U10729 (N_10729,N_9809,N_9513);
or U10730 (N_10730,N_8175,N_8351);
nand U10731 (N_10731,N_5748,N_6045);
and U10732 (N_10732,N_5862,N_7809);
or U10733 (N_10733,N_9245,N_7507);
nor U10734 (N_10734,N_6047,N_6270);
nand U10735 (N_10735,N_5782,N_5614);
and U10736 (N_10736,N_9073,N_8432);
and U10737 (N_10737,N_8258,N_7411);
or U10738 (N_10738,N_7477,N_6303);
or U10739 (N_10739,N_6539,N_7299);
or U10740 (N_10740,N_9737,N_6837);
xnor U10741 (N_10741,N_7779,N_6245);
nor U10742 (N_10742,N_8585,N_7083);
nor U10743 (N_10743,N_7070,N_6233);
nand U10744 (N_10744,N_6624,N_5088);
nand U10745 (N_10745,N_6344,N_7425);
nand U10746 (N_10746,N_7276,N_9375);
nand U10747 (N_10747,N_7964,N_5996);
nand U10748 (N_10748,N_5918,N_6681);
nand U10749 (N_10749,N_5115,N_5406);
nor U10750 (N_10750,N_9766,N_9750);
and U10751 (N_10751,N_6284,N_6891);
or U10752 (N_10752,N_5329,N_6517);
nor U10753 (N_10753,N_7997,N_8602);
or U10754 (N_10754,N_9482,N_9346);
nor U10755 (N_10755,N_7047,N_6808);
nand U10756 (N_10756,N_5367,N_7102);
or U10757 (N_10757,N_5131,N_5306);
nand U10758 (N_10758,N_5339,N_8316);
and U10759 (N_10759,N_9982,N_7094);
nand U10760 (N_10760,N_9774,N_6629);
or U10761 (N_10761,N_7359,N_8348);
and U10762 (N_10762,N_8774,N_6859);
or U10763 (N_10763,N_8260,N_8928);
and U10764 (N_10764,N_8365,N_9006);
or U10765 (N_10765,N_8127,N_8797);
and U10766 (N_10766,N_6101,N_9651);
or U10767 (N_10767,N_5542,N_6520);
or U10768 (N_10768,N_8751,N_5412);
nand U10769 (N_10769,N_9614,N_5383);
or U10770 (N_10770,N_7908,N_5841);
or U10771 (N_10771,N_7457,N_7152);
nor U10772 (N_10772,N_7898,N_7137);
or U10773 (N_10773,N_6203,N_6155);
nand U10774 (N_10774,N_6779,N_6179);
nand U10775 (N_10775,N_8232,N_7228);
nor U10776 (N_10776,N_8452,N_5566);
or U10777 (N_10777,N_7848,N_8972);
nand U10778 (N_10778,N_5303,N_9504);
xor U10779 (N_10779,N_5059,N_7388);
nor U10780 (N_10780,N_7343,N_9913);
or U10781 (N_10781,N_6795,N_5870);
nand U10782 (N_10782,N_7212,N_9220);
nand U10783 (N_10783,N_5818,N_7066);
nor U10784 (N_10784,N_9662,N_5693);
nand U10785 (N_10785,N_7020,N_6113);
xor U10786 (N_10786,N_5419,N_6464);
nand U10787 (N_10787,N_6689,N_5749);
nor U10788 (N_10788,N_8036,N_6838);
nand U10789 (N_10789,N_7403,N_5194);
or U10790 (N_10790,N_7554,N_6675);
nor U10791 (N_10791,N_8532,N_5116);
nand U10792 (N_10792,N_9929,N_8642);
and U10793 (N_10793,N_5860,N_5607);
nor U10794 (N_10794,N_6230,N_5418);
and U10795 (N_10795,N_5708,N_8500);
and U10796 (N_10796,N_6356,N_8366);
and U10797 (N_10797,N_5979,N_8393);
or U10798 (N_10798,N_5849,N_6186);
or U10799 (N_10799,N_7305,N_6737);
and U10800 (N_10800,N_8479,N_9212);
or U10801 (N_10801,N_9870,N_5935);
nand U10802 (N_10802,N_9002,N_7547);
nor U10803 (N_10803,N_7594,N_8016);
nor U10804 (N_10804,N_8427,N_8667);
and U10805 (N_10805,N_8637,N_6719);
and U10806 (N_10806,N_7310,N_6888);
nor U10807 (N_10807,N_5218,N_8927);
nand U10808 (N_10808,N_7668,N_5696);
nand U10809 (N_10809,N_7864,N_6600);
and U10810 (N_10810,N_8242,N_7015);
nand U10811 (N_10811,N_8453,N_7387);
and U10812 (N_10812,N_8171,N_6148);
nand U10813 (N_10813,N_5120,N_7258);
and U10814 (N_10814,N_5612,N_7819);
and U10815 (N_10815,N_6643,N_6697);
and U10816 (N_10816,N_5162,N_5985);
nand U10817 (N_10817,N_5029,N_8576);
and U10818 (N_10818,N_5576,N_6786);
nor U10819 (N_10819,N_5038,N_9626);
xnor U10820 (N_10820,N_7559,N_9842);
or U10821 (N_10821,N_9412,N_6950);
nand U10822 (N_10822,N_6780,N_6900);
nand U10823 (N_10823,N_6310,N_8345);
or U10824 (N_10824,N_9028,N_8462);
nand U10825 (N_10825,N_5914,N_9914);
nand U10826 (N_10826,N_5832,N_8152);
nor U10827 (N_10827,N_8646,N_9185);
nor U10828 (N_10828,N_5713,N_7368);
or U10829 (N_10829,N_6657,N_9741);
or U10830 (N_10830,N_7180,N_6562);
and U10831 (N_10831,N_5281,N_8000);
or U10832 (N_10832,N_5254,N_7466);
xor U10833 (N_10833,N_5587,N_9625);
nor U10834 (N_10834,N_9682,N_5947);
or U10835 (N_10835,N_6800,N_9618);
or U10836 (N_10836,N_9527,N_7878);
and U10837 (N_10837,N_8221,N_6422);
xnor U10838 (N_10838,N_6388,N_5894);
xnor U10839 (N_10839,N_9554,N_9511);
and U10840 (N_10840,N_8288,N_5461);
and U10841 (N_10841,N_9850,N_7444);
and U10842 (N_10842,N_6240,N_5857);
nand U10843 (N_10843,N_6035,N_9938);
or U10844 (N_10844,N_8075,N_7399);
and U10845 (N_10845,N_5609,N_5216);
or U10846 (N_10846,N_6436,N_6180);
nand U10847 (N_10847,N_9688,N_9657);
or U10848 (N_10848,N_7193,N_8359);
nand U10849 (N_10849,N_5884,N_7440);
nand U10850 (N_10850,N_6143,N_9976);
nor U10851 (N_10851,N_8801,N_7494);
nor U10852 (N_10852,N_5957,N_6421);
nand U10853 (N_10853,N_7221,N_8027);
nand U10854 (N_10854,N_6181,N_8002);
nor U10855 (N_10855,N_5468,N_5074);
nor U10856 (N_10856,N_7699,N_5243);
and U10857 (N_10857,N_5973,N_7261);
nor U10858 (N_10858,N_9274,N_5738);
and U10859 (N_10859,N_5924,N_6381);
xor U10860 (N_10860,N_9963,N_8854);
xor U10861 (N_10861,N_8549,N_7521);
xor U10862 (N_10862,N_7272,N_5083);
and U10863 (N_10863,N_8696,N_5595);
nand U10864 (N_10864,N_9442,N_7309);
nor U10865 (N_10865,N_5118,N_8564);
nor U10866 (N_10866,N_5572,N_5920);
nor U10867 (N_10867,N_8775,N_9032);
or U10868 (N_10868,N_7454,N_5626);
and U10869 (N_10869,N_6201,N_9493);
nand U10870 (N_10870,N_5842,N_8841);
and U10871 (N_10871,N_8440,N_9810);
nor U10872 (N_10872,N_7183,N_7035);
or U10873 (N_10873,N_8249,N_9861);
nor U10874 (N_10874,N_6757,N_8965);
nor U10875 (N_10875,N_5177,N_6099);
nor U10876 (N_10876,N_7455,N_9102);
xnor U10877 (N_10877,N_7803,N_6935);
nand U10878 (N_10878,N_5337,N_5808);
nand U10879 (N_10879,N_9125,N_7836);
and U10880 (N_10880,N_9374,N_8912);
or U10881 (N_10881,N_9956,N_9063);
nand U10882 (N_10882,N_9997,N_6747);
and U10883 (N_10883,N_6197,N_7490);
nor U10884 (N_10884,N_7934,N_8285);
xor U10885 (N_10885,N_8608,N_6465);
nor U10886 (N_10886,N_5780,N_5463);
or U10887 (N_10887,N_9402,N_8064);
and U10888 (N_10888,N_6292,N_7114);
and U10889 (N_10889,N_7210,N_7595);
nand U10890 (N_10890,N_6733,N_5492);
nor U10891 (N_10891,N_6882,N_6738);
and U10892 (N_10892,N_5560,N_5851);
nor U10893 (N_10893,N_8894,N_6053);
and U10894 (N_10894,N_7129,N_5134);
nor U10895 (N_10895,N_8186,N_5837);
and U10896 (N_10896,N_6425,N_5809);
nor U10897 (N_10897,N_7784,N_7680);
and U10898 (N_10898,N_5484,N_5840);
nor U10899 (N_10899,N_7645,N_7229);
or U10900 (N_10900,N_6104,N_9009);
and U10901 (N_10901,N_5282,N_6571);
and U10902 (N_10902,N_5549,N_6196);
or U10903 (N_10903,N_7858,N_8983);
or U10904 (N_10904,N_8754,N_9898);
or U10905 (N_10905,N_5336,N_6074);
nor U10906 (N_10906,N_7792,N_7516);
nor U10907 (N_10907,N_9454,N_8206);
and U10908 (N_10908,N_5796,N_5371);
nand U10909 (N_10909,N_9427,N_5725);
nor U10910 (N_10910,N_8185,N_9748);
or U10911 (N_10911,N_9087,N_5151);
and U10912 (N_10912,N_5377,N_9649);
or U10913 (N_10913,N_6401,N_9968);
nor U10914 (N_10914,N_8746,N_8838);
nor U10915 (N_10915,N_6341,N_6262);
and U10916 (N_10916,N_7893,N_6207);
nor U10917 (N_10917,N_8195,N_7955);
and U10918 (N_10918,N_5949,N_9331);
or U10919 (N_10919,N_8908,N_6494);
nand U10920 (N_10920,N_5350,N_5829);
nand U10921 (N_10921,N_6785,N_9660);
and U10922 (N_10922,N_6667,N_7277);
nand U10923 (N_10923,N_7919,N_5223);
nor U10924 (N_10924,N_8233,N_7609);
and U10925 (N_10925,N_9401,N_5874);
or U10926 (N_10926,N_7286,N_6472);
nor U10927 (N_10927,N_8034,N_9866);
or U10928 (N_10928,N_6518,N_8102);
and U10929 (N_10929,N_6351,N_9495);
nor U10930 (N_10930,N_9733,N_5557);
xnor U10931 (N_10931,N_9332,N_5758);
and U10932 (N_10932,N_5033,N_5091);
nand U10933 (N_10933,N_5885,N_6482);
nand U10934 (N_10934,N_5923,N_8931);
xnor U10935 (N_10935,N_9419,N_8265);
or U10936 (N_10936,N_6216,N_9985);
nand U10937 (N_10937,N_7290,N_8149);
xor U10938 (N_10938,N_7443,N_8744);
nor U10939 (N_10939,N_8628,N_8313);
nor U10940 (N_10940,N_6214,N_8197);
and U10941 (N_10941,N_5168,N_6380);
xor U10942 (N_10942,N_9053,N_7891);
or U10943 (N_10943,N_9239,N_9516);
xor U10944 (N_10944,N_7378,N_6711);
nor U10945 (N_10945,N_7288,N_9307);
nor U10946 (N_10946,N_6286,N_6817);
and U10947 (N_10947,N_6153,N_5656);
nor U10948 (N_10948,N_6252,N_5778);
nor U10949 (N_10949,N_8808,N_7500);
and U10950 (N_10950,N_6362,N_7965);
xor U10951 (N_10951,N_9977,N_6931);
xor U10952 (N_10952,N_8287,N_6919);
or U10953 (N_10953,N_6116,N_9406);
nor U10954 (N_10954,N_5392,N_7951);
or U10955 (N_10955,N_7488,N_7659);
and U10956 (N_10956,N_7637,N_6933);
nor U10957 (N_10957,N_5617,N_9479);
or U10958 (N_10958,N_5396,N_9762);
nand U10959 (N_10959,N_8985,N_8951);
or U10960 (N_10960,N_5655,N_7686);
nand U10961 (N_10961,N_5283,N_5253);
nand U10962 (N_10962,N_6855,N_9512);
or U10963 (N_10963,N_8066,N_7608);
xor U10964 (N_10964,N_8403,N_8297);
and U10965 (N_10965,N_7729,N_7612);
nand U10966 (N_10966,N_8482,N_7772);
xnor U10967 (N_10967,N_8757,N_8042);
xor U10968 (N_10968,N_8738,N_8020);
and U10969 (N_10969,N_5446,N_7944);
nor U10970 (N_10970,N_6826,N_5224);
nor U10971 (N_10971,N_8901,N_6683);
nor U10972 (N_10972,N_7082,N_9273);
nor U10973 (N_10973,N_6289,N_6501);
xor U10974 (N_10974,N_5440,N_8026);
and U10975 (N_10975,N_6912,N_9650);
or U10976 (N_10976,N_6500,N_9100);
nand U10977 (N_10977,N_5203,N_5618);
nor U10978 (N_10978,N_6803,N_5876);
and U10979 (N_10979,N_7096,N_6790);
nand U10980 (N_10980,N_6959,N_6059);
xor U10981 (N_10981,N_9069,N_6172);
nand U10982 (N_10982,N_5597,N_7708);
and U10983 (N_10983,N_5335,N_5266);
and U10984 (N_10984,N_8980,N_8977);
or U10985 (N_10985,N_8476,N_6625);
or U10986 (N_10986,N_9386,N_5058);
or U10987 (N_10987,N_9478,N_5093);
and U10988 (N_10988,N_9498,N_6523);
nand U10989 (N_10989,N_8327,N_9324);
or U10990 (N_10990,N_8322,N_9255);
xor U10991 (N_10991,N_5071,N_5673);
or U10992 (N_10992,N_8107,N_6566);
nor U10993 (N_10993,N_7613,N_5519);
nand U10994 (N_10994,N_7323,N_7969);
and U10995 (N_10995,N_9452,N_8823);
or U10996 (N_10996,N_8222,N_9936);
nand U10997 (N_10997,N_8967,N_6743);
nand U10998 (N_10998,N_9146,N_8209);
nor U10999 (N_10999,N_9155,N_5183);
and U11000 (N_11000,N_7520,N_7329);
nand U11001 (N_11001,N_5807,N_5402);
nor U11002 (N_11002,N_7189,N_8692);
nor U11003 (N_11003,N_5925,N_9663);
and U11004 (N_11004,N_8852,N_9283);
nor U11005 (N_11005,N_9854,N_8506);
or U11006 (N_11006,N_5368,N_6063);
or U11007 (N_11007,N_5559,N_8591);
and U11008 (N_11008,N_8884,N_6051);
and U11009 (N_11009,N_8380,N_5533);
and U11010 (N_11010,N_9290,N_9600);
or U11011 (N_11011,N_5212,N_7236);
or U11012 (N_11012,N_9282,N_5643);
or U11013 (N_11013,N_8004,N_8611);
or U11014 (N_11014,N_6295,N_8694);
and U11015 (N_11015,N_9871,N_7322);
nand U11016 (N_11016,N_5526,N_9894);
or U11017 (N_11017,N_9242,N_7394);
and U11018 (N_11018,N_5565,N_9857);
nor U11019 (N_11019,N_5501,N_9710);
or U11020 (N_11020,N_8745,N_8689);
nor U11021 (N_11021,N_6827,N_9044);
nand U11022 (N_11022,N_9561,N_5575);
nand U11023 (N_11023,N_6739,N_6751);
xor U11024 (N_11024,N_8067,N_9057);
and U11025 (N_11025,N_9148,N_7769);
and U11026 (N_11026,N_6222,N_8587);
and U11027 (N_11027,N_6608,N_6538);
and U11028 (N_11028,N_7382,N_7333);
nor U11029 (N_11029,N_9683,N_6583);
nand U11030 (N_11030,N_8663,N_5672);
or U11031 (N_11031,N_8771,N_6877);
xnor U11032 (N_11032,N_6124,N_7665);
or U11033 (N_11033,N_9546,N_7316);
or U11034 (N_11034,N_7226,N_8550);
or U11035 (N_11035,N_5255,N_9476);
xor U11036 (N_11036,N_6504,N_5990);
nor U11037 (N_11037,N_6247,N_8029);
and U11038 (N_11038,N_5970,N_6120);
xor U11039 (N_11039,N_7331,N_9107);
or U11040 (N_11040,N_5883,N_5647);
or U11041 (N_11041,N_8247,N_7820);
and U11042 (N_11042,N_8610,N_8105);
nor U11043 (N_11043,N_5080,N_9752);
or U11044 (N_11044,N_9016,N_5664);
xnor U11045 (N_11045,N_5089,N_6529);
and U11046 (N_11046,N_7987,N_9420);
and U11047 (N_11047,N_6369,N_8397);
or U11048 (N_11048,N_6427,N_5137);
and U11049 (N_11049,N_5991,N_9686);
xnor U11050 (N_11050,N_7130,N_8295);
and U11051 (N_11051,N_5675,N_5122);
nor U11052 (N_11052,N_9687,N_9885);
and U11053 (N_11053,N_9931,N_7902);
xor U11054 (N_11054,N_9534,N_5721);
nand U11055 (N_11055,N_5768,N_8596);
nor U11056 (N_11056,N_9347,N_7448);
nand U11057 (N_11057,N_7553,N_6690);
nand U11058 (N_11058,N_8773,N_9443);
nor U11059 (N_11059,N_5051,N_8786);
or U11060 (N_11060,N_9950,N_9724);
nor U11061 (N_11061,N_7463,N_8341);
nor U11062 (N_11062,N_7389,N_8973);
xor U11063 (N_11063,N_8513,N_7811);
and U11064 (N_11064,N_9800,N_6507);
and U11065 (N_11065,N_9562,N_7519);
xnor U11066 (N_11066,N_8969,N_7946);
and U11067 (N_11067,N_7904,N_7437);
and U11068 (N_11068,N_8812,N_9639);
nor U11069 (N_11069,N_7068,N_9702);
nand U11070 (N_11070,N_6973,N_7611);
nand U11071 (N_11071,N_9425,N_8415);
nand U11072 (N_11072,N_5677,N_6630);
nor U11073 (N_11073,N_6185,N_7763);
nand U11074 (N_11074,N_5531,N_5981);
and U11075 (N_11075,N_8298,N_8780);
nand U11076 (N_11076,N_7093,N_9267);
or U11077 (N_11077,N_5234,N_8670);
or U11078 (N_11078,N_8936,N_8275);
or U11079 (N_11079,N_5138,N_8556);
or U11080 (N_11080,N_8840,N_9635);
nand U11081 (N_11081,N_6489,N_5821);
and U11082 (N_11082,N_8119,N_8497);
nor U11083 (N_11083,N_6399,N_8600);
and U11084 (N_11084,N_8859,N_7621);
nand U11085 (N_11085,N_5219,N_8420);
xor U11086 (N_11086,N_5983,N_8514);
and U11087 (N_11087,N_7022,N_6754);
or U11088 (N_11088,N_9491,N_9494);
or U11089 (N_11089,N_7657,N_6354);
and U11090 (N_11090,N_6902,N_8623);
xor U11091 (N_11091,N_6940,N_8053);
xnor U11092 (N_11092,N_5727,N_5157);
and U11093 (N_11093,N_9170,N_7271);
xnor U11094 (N_11094,N_8284,N_8544);
nand U11095 (N_11095,N_9583,N_8741);
nor U11096 (N_11096,N_8017,N_8189);
nand U11097 (N_11097,N_5736,N_8621);
nor U11098 (N_11098,N_6987,N_7117);
or U11099 (N_11099,N_5154,N_8647);
or U11100 (N_11100,N_9603,N_7568);
nand U11101 (N_11101,N_8211,N_7730);
nor U11102 (N_11102,N_7534,N_5346);
xor U11103 (N_11103,N_7748,N_8635);
nor U11104 (N_11104,N_6032,N_5431);
nand U11105 (N_11105,N_7722,N_9636);
or U11106 (N_11106,N_9903,N_9213);
and U11107 (N_11107,N_6521,N_9333);
nand U11108 (N_11108,N_7642,N_6801);
or U11109 (N_11109,N_8137,N_7352);
nand U11110 (N_11110,N_5702,N_5308);
nor U11111 (N_11111,N_8992,N_6168);
nor U11112 (N_11112,N_8269,N_9093);
nor U11113 (N_11113,N_5362,N_6137);
nor U11114 (N_11114,N_8733,N_7198);
nor U11115 (N_11115,N_7458,N_8141);
and U11116 (N_11116,N_5836,N_8236);
or U11117 (N_11117,N_7452,N_7268);
xor U11118 (N_11118,N_9515,N_7671);
nor U11119 (N_11119,N_5478,N_9257);
nand U11120 (N_11120,N_9411,N_5094);
or U11121 (N_11121,N_6721,N_6975);
nand U11122 (N_11122,N_7614,N_9235);
or U11123 (N_11123,N_5766,N_9773);
nand U11124 (N_11124,N_5511,N_8994);
nor U11125 (N_11125,N_6361,N_6141);
and U11126 (N_11126,N_8698,N_5527);
nand U11127 (N_11127,N_5354,N_5236);
or U11128 (N_11128,N_8438,N_8248);
nor U11129 (N_11129,N_8077,N_7409);
or U11130 (N_11130,N_7652,N_6126);
or U11131 (N_11131,N_8391,N_7866);
and U11132 (N_11132,N_9318,N_5654);
xnor U11133 (N_11133,N_6927,N_8320);
nand U11134 (N_11134,N_7319,N_6899);
nand U11135 (N_11135,N_5287,N_6244);
nor U11136 (N_11136,N_8728,N_5641);
nand U11137 (N_11137,N_8906,N_7435);
nor U11138 (N_11138,N_6515,N_9795);
and U11139 (N_11139,N_8874,N_7247);
nor U11140 (N_11140,N_7338,N_5921);
nand U11141 (N_11141,N_7416,N_5516);
and U11142 (N_11142,N_7745,N_9604);
or U11143 (N_11143,N_9343,N_5787);
nand U11144 (N_11144,N_6088,N_9404);
nor U11145 (N_11145,N_9767,N_7529);
nand U11146 (N_11146,N_9497,N_5035);
or U11147 (N_11147,N_9701,N_9547);
nor U11148 (N_11148,N_9072,N_8290);
xor U11149 (N_11149,N_8052,N_7245);
nor U11150 (N_11150,N_7669,N_7827);
and U11151 (N_11151,N_6073,N_5496);
nand U11152 (N_11152,N_9005,N_9295);
or U11153 (N_11153,N_7282,N_9178);
nor U11154 (N_11154,N_8399,N_7267);
xor U11155 (N_11155,N_8038,N_5520);
xor U11156 (N_11156,N_9358,N_5905);
and U11157 (N_11157,N_5897,N_5509);
xnor U11158 (N_11158,N_5513,N_9579);
xor U11159 (N_11159,N_7877,N_8582);
xnor U11160 (N_11160,N_9996,N_6835);
nor U11161 (N_11161,N_8846,N_8083);
and U11162 (N_11162,N_9438,N_7101);
nor U11163 (N_11163,N_6402,N_6766);
or U11164 (N_11164,N_9926,N_7966);
or U11165 (N_11165,N_9197,N_5054);
xnor U11166 (N_11166,N_5052,N_7690);
nand U11167 (N_11167,N_5025,N_9179);
nand U11168 (N_11168,N_5471,N_8865);
or U11169 (N_11169,N_5754,N_6614);
nor U11170 (N_11170,N_5965,N_7293);
or U11171 (N_11171,N_6580,N_5473);
or U11172 (N_11172,N_5781,N_5462);
nor U11173 (N_11173,N_5580,N_9075);
xor U11174 (N_11174,N_5602,N_9771);
nand U11175 (N_11175,N_9142,N_6886);
xnor U11176 (N_11176,N_9585,N_9261);
or U11177 (N_11177,N_8396,N_7194);
nor U11178 (N_11178,N_8560,N_8123);
nor U11179 (N_11179,N_9500,N_8524);
xor U11180 (N_11180,N_6375,N_9726);
and U11181 (N_11181,N_8121,N_8844);
nor U11182 (N_11182,N_9715,N_7453);
and U11183 (N_11183,N_7778,N_9429);
and U11184 (N_11184,N_9435,N_8237);
nand U11185 (N_11185,N_7473,N_8676);
or U11186 (N_11186,N_9580,N_7892);
or U11187 (N_11187,N_9911,N_5669);
and U11188 (N_11188,N_5966,N_7561);
xor U11189 (N_11189,N_8781,N_7079);
nand U11190 (N_11190,N_9951,N_7421);
nor U11191 (N_11191,N_5795,N_9523);
nand U11192 (N_11192,N_8477,N_7300);
or U11193 (N_11193,N_5055,N_8350);
and U11194 (N_11194,N_8573,N_5220);
or U11195 (N_11195,N_5667,N_7927);
and U11196 (N_11196,N_9770,N_5843);
and U11197 (N_11197,N_9749,N_8059);
nand U11198 (N_11198,N_5376,N_8999);
or U11199 (N_11199,N_6293,N_9671);
or U11200 (N_11200,N_6030,N_6182);
or U11201 (N_11201,N_5315,N_5814);
nor U11202 (N_11202,N_9014,N_8541);
and U11203 (N_11203,N_8244,N_9094);
or U11204 (N_11204,N_9637,N_9369);
and U11205 (N_11205,N_8707,N_9582);
and U11206 (N_11206,N_7910,N_9457);
or U11207 (N_11207,N_6417,N_6446);
nor U11208 (N_11208,N_8666,N_8338);
or U11209 (N_11209,N_9400,N_9521);
and U11210 (N_11210,N_9678,N_9081);
nor U11211 (N_11211,N_6663,N_5764);
nand U11212 (N_11212,N_7567,N_7173);
or U11213 (N_11213,N_9879,N_7222);
nand U11214 (N_11214,N_9441,N_6221);
nand U11215 (N_11215,N_8729,N_7624);
xnor U11216 (N_11216,N_8804,N_7324);
nor U11217 (N_11217,N_5272,N_6390);
or U11218 (N_11218,N_7397,N_5388);
and U11219 (N_11219,N_8650,N_6946);
and U11220 (N_11220,N_6140,N_7640);
and U11221 (N_11221,N_9915,N_7191);
xor U11222 (N_11222,N_8659,N_7802);
and U11223 (N_11223,N_9224,N_5321);
and U11224 (N_11224,N_5543,N_7050);
nand U11225 (N_11225,N_9532,N_8270);
nor U11226 (N_11226,N_6281,N_5428);
nand U11227 (N_11227,N_9834,N_8360);
xor U11228 (N_11228,N_6932,N_8770);
or U11229 (N_11229,N_7865,N_5548);
nand U11230 (N_11230,N_6774,N_7590);
nor U11231 (N_11231,N_9253,N_8060);
nor U11232 (N_11232,N_8614,N_7538);
or U11233 (N_11233,N_9753,N_5410);
nor U11234 (N_11234,N_9658,N_7683);
and U11235 (N_11235,N_9043,N_6269);
or U11236 (N_11236,N_7142,N_9946);
xnor U11237 (N_11237,N_8148,N_9812);
xnor U11238 (N_11238,N_7178,N_9460);
or U11239 (N_11239,N_8495,N_6330);
nor U11240 (N_11240,N_8496,N_8821);
and U11241 (N_11241,N_7829,N_7471);
and U11242 (N_11242,N_5066,N_6776);
nor U11243 (N_11243,N_5634,N_5881);
and U11244 (N_11244,N_6952,N_5978);
nand U11245 (N_11245,N_6166,N_9394);
nor U11246 (N_11246,N_5166,N_5064);
xnor U11247 (N_11247,N_9680,N_5969);
nand U11248 (N_11248,N_6707,N_9979);
nand U11249 (N_11249,N_6300,N_7464);
nand U11250 (N_11250,N_5044,N_9133);
and U11251 (N_11251,N_8740,N_6320);
and U11252 (N_11252,N_8318,N_7720);
nand U11253 (N_11253,N_5558,N_8412);
nor U11254 (N_11254,N_9611,N_9373);
nor U11255 (N_11255,N_9462,N_9299);
or U11256 (N_11256,N_6146,N_7476);
or U11257 (N_11257,N_8334,N_8124);
xnor U11258 (N_11258,N_9575,N_6129);
or U11259 (N_11259,N_9392,N_7840);
or U11260 (N_11260,N_5529,N_5801);
nand U11261 (N_11261,N_6312,N_6441);
nand U11262 (N_11262,N_7122,N_5380);
or U11263 (N_11263,N_7401,N_5244);
or U11264 (N_11264,N_7777,N_6799);
xnor U11265 (N_11265,N_6259,N_7406);
and U11266 (N_11266,N_5414,N_8686);
nor U11267 (N_11267,N_8028,N_6953);
and U11268 (N_11268,N_9193,N_9353);
or U11269 (N_11269,N_8789,N_6620);
nor U11270 (N_11270,N_9355,N_5225);
nor U11271 (N_11271,N_6397,N_7469);
and U11272 (N_11272,N_7989,N_7655);
or U11273 (N_11273,N_8078,N_5169);
or U11274 (N_11274,N_6075,N_5259);
or U11275 (N_11275,N_8858,N_6348);
nand U11276 (N_11276,N_7351,N_5962);
nor U11277 (N_11277,N_5709,N_7396);
nand U11278 (N_11278,N_8069,N_8210);
and U11279 (N_11279,N_6152,N_8842);
and U11280 (N_11280,N_7465,N_8379);
nor U11281 (N_11281,N_6193,N_8685);
nor U11282 (N_11282,N_9115,N_8118);
nor U11283 (N_11283,N_6512,N_9818);
nand U11284 (N_11284,N_6327,N_7607);
or U11285 (N_11285,N_7169,N_7325);
or U11286 (N_11286,N_9599,N_5668);
nand U11287 (N_11287,N_6670,N_6828);
and U11288 (N_11288,N_7144,N_8830);
or U11289 (N_11289,N_5239,N_8411);
and U11290 (N_11290,N_5571,N_7845);
nand U11291 (N_11291,N_7328,N_5824);
xnor U11292 (N_11292,N_6298,N_7797);
nor U11293 (N_11293,N_5540,N_7903);
nor U11294 (N_11294,N_7242,N_8887);
nand U11295 (N_11295,N_6787,N_8726);
and U11296 (N_11296,N_7480,N_6964);
and U11297 (N_11297,N_6442,N_9101);
and U11298 (N_11298,N_8559,N_7280);
and U11299 (N_11299,N_8863,N_7721);
nor U11300 (N_11300,N_9233,N_7000);
or U11301 (N_11301,N_6239,N_8940);
or U11302 (N_11302,N_8711,N_7714);
and U11303 (N_11303,N_7248,N_9403);
or U11304 (N_11304,N_7361,N_7536);
and U11305 (N_11305,N_8515,N_6324);
nor U11306 (N_11306,N_9541,N_8831);
or U11307 (N_11307,N_8177,N_8834);
and U11308 (N_11308,N_6770,N_7957);
and U11309 (N_11309,N_5153,N_9011);
nor U11310 (N_11310,N_9505,N_7061);
xnor U11311 (N_11311,N_7785,N_5774);
xor U11312 (N_11312,N_7225,N_6640);
and U11313 (N_11313,N_7650,N_5173);
nand U11314 (N_11314,N_5155,N_7727);
nor U11315 (N_11315,N_5430,N_7770);
nor U11316 (N_11316,N_6578,N_5535);
nor U11317 (N_11317,N_9821,N_7735);
xnor U11318 (N_11318,N_5456,N_8018);
or U11319 (N_11319,N_8782,N_5399);
nand U11320 (N_11320,N_7164,N_6260);
or U11321 (N_11321,N_6307,N_6532);
or U11322 (N_11322,N_8855,N_9828);
and U11323 (N_11323,N_5149,N_5603);
nor U11324 (N_11324,N_6237,N_9822);
nor U11325 (N_11325,N_5082,N_8088);
nor U11326 (N_11326,N_5638,N_9294);
or U11327 (N_11327,N_5221,N_6938);
nand U11328 (N_11328,N_9890,N_8826);
or U11329 (N_11329,N_7626,N_7550);
or U11330 (N_11330,N_6429,N_6905);
nor U11331 (N_11331,N_7181,N_8454);
and U11332 (N_11332,N_9508,N_5980);
nand U11333 (N_11333,N_6495,N_7414);
nor U11334 (N_11334,N_5078,N_5277);
nand U11335 (N_11335,N_9897,N_6762);
nor U11336 (N_11336,N_9379,N_7528);
and U11337 (N_11337,N_8862,N_8183);
nand U11338 (N_11338,N_7821,N_9390);
and U11339 (N_11339,N_9342,N_9483);
or U11340 (N_11340,N_6029,N_9272);
and U11341 (N_11341,N_8529,N_9868);
or U11342 (N_11342,N_6243,N_9990);
nor U11343 (N_11343,N_7695,N_8090);
nand U11344 (N_11344,N_7148,N_5771);
nand U11345 (N_11345,N_6773,N_7817);
nand U11346 (N_11346,N_8530,N_6579);
or U11347 (N_11347,N_6724,N_9623);
or U11348 (N_11348,N_8041,N_7462);
nor U11349 (N_11349,N_8202,N_6992);
nand U11350 (N_11350,N_9086,N_9440);
and U11351 (N_11351,N_9947,N_8517);
and U11352 (N_11352,N_5032,N_9553);
and U11353 (N_11353,N_7920,N_8594);
and U11354 (N_11354,N_9370,N_8352);
nand U11355 (N_11355,N_8170,N_7377);
or U11356 (N_11356,N_5743,N_8463);
nor U11357 (N_11357,N_8904,N_7566);
nor U11358 (N_11358,N_5958,N_5679);
nand U11359 (N_11359,N_6969,N_7926);
and U11360 (N_11360,N_8241,N_6662);
and U11361 (N_11361,N_6839,N_7837);
and U11362 (N_11362,N_9833,N_6740);
nor U11363 (N_11363,N_9992,N_7832);
or U11364 (N_11364,N_5683,N_7049);
nand U11365 (N_11365,N_5360,N_9310);
nor U11366 (N_11366,N_9475,N_5457);
nand U11367 (N_11367,N_6419,N_6167);
or U11368 (N_11368,N_9619,N_6929);
and U11369 (N_11369,N_7209,N_7940);
or U11370 (N_11370,N_8622,N_5546);
nor U11371 (N_11371,N_6187,N_7016);
or U11372 (N_11372,N_6558,N_6475);
and U11373 (N_11373,N_5021,N_9872);
nand U11374 (N_11374,N_6680,N_7253);
or U11375 (N_11375,N_6248,N_6405);
and U11376 (N_11376,N_8226,N_9616);
or U11377 (N_11377,N_9573,N_6778);
or U11378 (N_11378,N_6848,N_8649);
nor U11379 (N_11379,N_9251,N_6437);
and U11380 (N_11380,N_7034,N_8133);
or U11381 (N_11381,N_9126,N_7140);
or U11382 (N_11382,N_5767,N_9067);
or U11383 (N_11383,N_7139,N_5013);
nand U11384 (N_11384,N_5319,N_6982);
and U11385 (N_11385,N_6777,N_5172);
or U11386 (N_11386,N_6768,N_9567);
and U11387 (N_11387,N_8684,N_8321);
and U11388 (N_11388,N_8336,N_9967);
and U11389 (N_11389,N_6138,N_7707);
and U11390 (N_11390,N_5988,N_8251);
nor U11391 (N_11391,N_7348,N_7244);
and U11392 (N_11392,N_6516,N_6177);
and U11393 (N_11393,N_9617,N_5031);
or U11394 (N_11394,N_5026,N_9544);
and U11395 (N_11395,N_5307,N_9902);
nor U11396 (N_11396,N_5724,N_8423);
nand U11397 (N_11397,N_9518,N_7667);
or U11398 (N_11398,N_9841,N_5314);
nand U11399 (N_11399,N_7250,N_8739);
nand U11400 (N_11400,N_9444,N_8706);
and U11401 (N_11401,N_8456,N_5813);
nor U11402 (N_11402,N_5256,N_9845);
or U11403 (N_11403,N_5128,N_7733);
nand U11404 (N_11404,N_5828,N_9027);
and U11405 (N_11405,N_9531,N_5141);
nor U11406 (N_11406,N_6678,N_9076);
nand U11407 (N_11407,N_5692,N_9634);
nand U11408 (N_11408,N_6018,N_5260);
nand U11409 (N_11409,N_7679,N_9129);
and U11410 (N_11410,N_9492,N_8033);
xor U11411 (N_11411,N_6533,N_8864);
nor U11412 (N_11412,N_5784,N_8963);
nor U11413 (N_11413,N_8339,N_6576);
xor U11414 (N_11414,N_7158,N_8238);
nor U11415 (N_11415,N_5467,N_9136);
or U11416 (N_11416,N_6318,N_8410);
nand U11417 (N_11417,N_8372,N_6151);
or U11418 (N_11418,N_9209,N_8480);
nand U11419 (N_11419,N_8579,N_7373);
or U11420 (N_11420,N_8131,N_7357);
and U11421 (N_11421,N_6647,N_8464);
or U11422 (N_11422,N_9157,N_8998);
and U11423 (N_11423,N_7648,N_6746);
or U11424 (N_11424,N_6708,N_6955);
nand U11425 (N_11425,N_6423,N_8850);
nor U11426 (N_11426,N_8103,N_9638);
xor U11427 (N_11427,N_9792,N_9019);
nor U11428 (N_11428,N_8227,N_9590);
nor U11429 (N_11429,N_5521,N_7630);
or U11430 (N_11430,N_8481,N_5041);
or U11431 (N_11431,N_7315,N_6170);
or U11432 (N_11432,N_5777,N_9591);
nand U11433 (N_11433,N_5426,N_6924);
and U11434 (N_11434,N_8147,N_5971);
nand U11435 (N_11435,N_7042,N_7340);
nor U11436 (N_11436,N_6033,N_5424);
nand U11437 (N_11437,N_5872,N_9962);
or U11438 (N_11438,N_7870,N_9348);
nor U11439 (N_11439,N_7111,N_5364);
nor U11440 (N_11440,N_9615,N_7995);
nor U11441 (N_11441,N_9328,N_5213);
nand U11442 (N_11442,N_9801,N_8857);
nand U11443 (N_11443,N_8353,N_8627);
xor U11444 (N_11444,N_6430,N_6715);
nor U11445 (N_11445,N_5420,N_8618);
nand U11446 (N_11446,N_7576,N_6241);
nor U11447 (N_11447,N_7808,N_7054);
nor U11448 (N_11448,N_6046,N_8357);
nand U11449 (N_11449,N_8502,N_8819);
and U11450 (N_11450,N_8909,N_5458);
and U11451 (N_11451,N_6750,N_5585);
and U11452 (N_11452,N_8434,N_7914);
nand U11453 (N_11453,N_9108,N_8025);
nand U11454 (N_11454,N_5237,N_8159);
or U11455 (N_11455,N_8957,N_5658);
nand U11456 (N_11456,N_5579,N_6450);
nand U11457 (N_11457,N_9344,N_9691);
and U11458 (N_11458,N_5470,N_9096);
or U11459 (N_11459,N_7544,N_6149);
nor U11460 (N_11460,N_7776,N_8407);
xnor U11461 (N_11461,N_8613,N_7740);
nand U11462 (N_11462,N_8597,N_9705);
nand U11463 (N_11463,N_8375,N_9648);
xor U11464 (N_11464,N_7187,N_6107);
nor U11465 (N_11465,N_8394,N_7184);
or U11466 (N_11466,N_8593,N_9337);
nor U11467 (N_11467,N_6132,N_8246);
or U11468 (N_11468,N_9160,N_6542);
nand U11469 (N_11469,N_9308,N_5528);
nor U11470 (N_11470,N_9747,N_9539);
and U11471 (N_11471,N_7948,N_9882);
and U11472 (N_11472,N_8681,N_8837);
and U11473 (N_11473,N_7135,N_8081);
or U11474 (N_11474,N_8418,N_9448);
nand U11475 (N_11475,N_5102,N_8450);
or U11476 (N_11476,N_9731,N_5502);
nor U11477 (N_11477,N_5290,N_9876);
nor U11478 (N_11478,N_8068,N_7491);
or U11479 (N_11479,N_6202,N_7252);
nor U11480 (N_11480,N_9451,N_9003);
nor U11481 (N_11481,N_5067,N_6204);
or U11482 (N_11482,N_6574,N_8732);
or U11483 (N_11483,N_5500,N_5665);
nand U11484 (N_11484,N_8301,N_5762);
xor U11485 (N_11485,N_6843,N_6587);
and U11486 (N_11486,N_8643,N_6865);
nand U11487 (N_11487,N_6989,N_9189);
and U11488 (N_11488,N_7685,N_6264);
nand U11489 (N_11489,N_5285,N_7706);
nor U11490 (N_11490,N_6090,N_8389);
and U11491 (N_11491,N_5561,N_6594);
or U11492 (N_11492,N_6874,N_6338);
or U11493 (N_11493,N_5009,N_9225);
and U11494 (N_11494,N_5997,N_7163);
and U11495 (N_11495,N_6720,N_8483);
xnor U11496 (N_11496,N_5053,N_5995);
or U11497 (N_11497,N_6997,N_5384);
nor U11498 (N_11498,N_6486,N_6534);
nand U11499 (N_11499,N_8636,N_8406);
nor U11500 (N_11500,N_6672,N_7558);
nor U11501 (N_11501,N_5113,N_6908);
nor U11502 (N_11502,N_7563,N_8104);
and U11503 (N_11503,N_5610,N_9316);
or U11504 (N_11504,N_8426,N_9940);
or U11505 (N_11505,N_6897,N_7204);
nand U11506 (N_11506,N_8451,N_7087);
and U11507 (N_11507,N_5262,N_5289);
nand U11508 (N_11508,N_9907,N_7048);
and U11509 (N_11509,N_6606,N_7291);
nor U11510 (N_11510,N_6125,N_6632);
or U11511 (N_11511,N_6958,N_6956);
xor U11512 (N_11512,N_6761,N_7259);
or U11513 (N_11513,N_9329,N_8065);
or U11514 (N_11514,N_9084,N_8084);
and U11515 (N_11515,N_5159,N_9605);
nor U11516 (N_11516,N_8460,N_6322);
nor U11517 (N_11517,N_8212,N_6439);
and U11518 (N_11518,N_5737,N_8695);
nand U11519 (N_11519,N_8306,N_9860);
nor U11520 (N_11520,N_7885,N_6412);
or U11521 (N_11521,N_7812,N_8950);
and U11522 (N_11522,N_9769,N_5356);
nand U11523 (N_11523,N_8824,N_5907);
nand U11524 (N_11524,N_8315,N_6917);
xor U11525 (N_11525,N_6540,N_9421);
nand U11526 (N_11526,N_6136,N_8755);
nand U11527 (N_11527,N_8280,N_8080);
xor U11528 (N_11528,N_7318,N_6555);
xor U11529 (N_11529,N_7649,N_9862);
nand U11530 (N_11530,N_7251,N_9306);
nor U11531 (N_11531,N_7071,N_6057);
xor U11532 (N_11532,N_5482,N_6904);
nand U11533 (N_11533,N_9932,N_6044);
or U11534 (N_11534,N_7143,N_5443);
and U11535 (N_11535,N_8157,N_6619);
nand U11536 (N_11536,N_7428,N_7475);
and U11537 (N_11537,N_9557,N_9437);
nor U11538 (N_11538,N_5695,N_5422);
nand U11539 (N_11539,N_8800,N_6459);
or U11540 (N_11540,N_8311,N_8595);
nand U11541 (N_11541,N_7195,N_5908);
nor U11542 (N_11542,N_8727,N_6998);
and U11543 (N_11543,N_6782,N_7548);
nand U11544 (N_11544,N_8143,N_7023);
or U11545 (N_11545,N_9430,N_9739);
and U11546 (N_11546,N_7842,N_5938);
nand U11547 (N_11547,N_9097,N_8478);
nor U11548 (N_11548,N_7766,N_8492);
or U11549 (N_11549,N_6769,N_9030);
and U11550 (N_11550,N_6406,N_6728);
or U11551 (N_11551,N_5570,N_9569);
nand U11552 (N_11552,N_8934,N_6393);
nor U11553 (N_11553,N_8192,N_5494);
nand U11554 (N_11554,N_8958,N_5104);
and U11555 (N_11555,N_5534,N_7149);
or U11556 (N_11556,N_9791,N_7483);
nand U11557 (N_11557,N_5715,N_9552);
nor U11558 (N_11558,N_6271,N_7615);
nand U11559 (N_11559,N_7716,N_5545);
nor U11560 (N_11560,N_9025,N_5739);
or U11561 (N_11561,N_6965,N_9796);
nor U11562 (N_11562,N_7533,N_8677);
nor U11563 (N_11563,N_9577,N_6114);
and U11564 (N_11564,N_7977,N_9490);
nand U11565 (N_11565,N_7627,N_5688);
or U11566 (N_11566,N_7172,N_8683);
nor U11567 (N_11567,N_6526,N_7302);
nor U11568 (N_11568,N_6413,N_6403);
nand U11569 (N_11569,N_6424,N_5681);
nand U11570 (N_11570,N_8817,N_5312);
or U11571 (N_11571,N_9793,N_8993);
nand U11572 (N_11572,N_6225,N_6316);
or U11573 (N_11573,N_5075,N_7937);
nand U11574 (N_11574,N_7744,N_9595);
nand U11575 (N_11575,N_7363,N_9670);
nor U11576 (N_11576,N_5830,N_8743);
and U11577 (N_11577,N_7805,N_8795);
or U11578 (N_11578,N_9154,N_8048);
and U11579 (N_11579,N_5378,N_7063);
nand U11580 (N_11580,N_5888,N_8570);
xor U11581 (N_11581,N_6918,N_9426);
or U11582 (N_11582,N_5629,N_6742);
nand U11583 (N_11583,N_9654,N_7644);
or U11584 (N_11584,N_6868,N_7439);
nor U11585 (N_11585,N_7133,N_7916);
or U11586 (N_11586,N_9064,N_7482);
nor U11587 (N_11587,N_9652,N_9507);
or U11588 (N_11588,N_9023,N_7980);
or U11589 (N_11589,N_5024,N_9204);
or U11590 (N_11590,N_7215,N_9874);
nor U11591 (N_11591,N_7109,N_5551);
nand U11592 (N_11592,N_9653,N_9681);
and U11593 (N_11593,N_9945,N_8509);
xnor U11594 (N_11594,N_9761,N_5046);
nor U11595 (N_11595,N_9070,N_7367);
xnor U11596 (N_11596,N_7896,N_7890);
and U11597 (N_11597,N_6767,N_9221);
xor U11598 (N_11598,N_6016,N_9530);
xor U11599 (N_11599,N_6557,N_9198);
and U11600 (N_11600,N_6385,N_9798);
or U11601 (N_11601,N_9886,N_8620);
xor U11602 (N_11602,N_7166,N_5106);
nor U11603 (N_11603,N_9644,N_9909);
and U11604 (N_11604,N_9065,N_7131);
and U11605 (N_11605,N_9399,N_8240);
nand U11606 (N_11606,N_7092,N_7998);
nor U11607 (N_11607,N_9524,N_6581);
or U11608 (N_11608,N_5435,N_7684);
and U11609 (N_11609,N_5432,N_8709);
nor U11610 (N_11610,N_9381,N_9987);
or U11611 (N_11611,N_6349,N_6209);
or U11612 (N_11612,N_9286,N_7814);
nor U11613 (N_11613,N_7601,N_7345);
nor U11614 (N_11614,N_8405,N_5723);
and U11615 (N_11615,N_6191,N_7935);
xor U11616 (N_11616,N_7106,N_6513);
or U11617 (N_11617,N_7764,N_5487);
xor U11618 (N_11618,N_9105,N_7542);
nor U11619 (N_11619,N_9237,N_5455);
or U11620 (N_11620,N_6631,N_8699);
nand U11621 (N_11621,N_6133,N_8822);
nor U11622 (N_11622,N_7688,N_5345);
and U11623 (N_11623,N_6194,N_9666);
or U11624 (N_11624,N_9522,N_6068);
nor U11625 (N_11625,N_7008,N_6481);
or U11626 (N_11626,N_8332,N_6378);
xnor U11627 (N_11627,N_6192,N_5291);
nand U11628 (N_11628,N_8001,N_7818);
nor U11629 (N_11629,N_8109,N_7543);
nor U11630 (N_11630,N_9271,N_7923);
and U11631 (N_11631,N_8783,N_7355);
and U11632 (N_11632,N_7012,N_7899);
nor U11633 (N_11633,N_5382,N_7510);
nor U11634 (N_11634,N_8193,N_7661);
nand U11635 (N_11635,N_5512,N_8310);
nor U11636 (N_11636,N_5476,N_7052);
and U11637 (N_11637,N_6112,N_8400);
xnor U11638 (N_11638,N_8955,N_8408);
nand U11639 (N_11639,N_8935,N_8335);
or U11640 (N_11640,N_5699,N_9121);
nor U11641 (N_11641,N_7289,N_7459);
or U11642 (N_11642,N_5967,N_7053);
nand U11643 (N_11643,N_9713,N_8055);
nor U11644 (N_11644,N_5228,N_9565);
or U11645 (N_11645,N_7913,N_8475);
nand U11646 (N_11646,N_6660,N_9744);
or U11647 (N_11647,N_9384,N_6323);
nand U11648 (N_11648,N_5238,N_8680);
xnor U11649 (N_11649,N_6686,N_5998);
xnor U11650 (N_11650,N_5619,N_9356);
and U11651 (N_11651,N_6648,N_6091);
nor U11652 (N_11652,N_9020,N_8721);
nand U11653 (N_11653,N_6360,N_5869);
xor U11654 (N_11654,N_9288,N_9995);
xnor U11655 (N_11655,N_7993,N_9312);
and U11656 (N_11656,N_7056,N_5915);
nor U11657 (N_11657,N_5366,N_9803);
or U11658 (N_11658,N_7113,N_9904);
nand U11659 (N_11659,N_6654,N_7395);
nand U11660 (N_11660,N_8907,N_9642);
xor U11661 (N_11661,N_6860,N_9760);
nand U11662 (N_11662,N_8723,N_9714);
nand U11663 (N_11663,N_7924,N_6326);
nor U11664 (N_11664,N_8665,N_7279);
xor U11665 (N_11665,N_9503,N_6077);
nor U11666 (N_11666,N_8599,N_9742);
nor U11667 (N_11667,N_7124,N_9869);
and U11668 (N_11668,N_7040,N_7481);
and U11669 (N_11669,N_6159,N_5747);
or U11670 (N_11670,N_8941,N_6943);
nand U11671 (N_11671,N_8658,N_7674);
and U11672 (N_11672,N_7598,N_7907);
nand U11673 (N_11673,N_7472,N_9672);
or U11674 (N_11674,N_9321,N_8586);
or U11675 (N_11675,N_9700,N_5401);
xor U11676 (N_11676,N_5555,N_7509);
nand U11677 (N_11677,N_7307,N_9078);
nand U11678 (N_11678,N_6200,N_5646);
nand U11679 (N_11679,N_5662,N_6317);
and U11680 (N_11680,N_8735,N_9297);
nor U11681 (N_11681,N_6695,N_9933);
or U11682 (N_11682,N_8984,N_7014);
nor U11683 (N_11683,N_6598,N_8111);
nor U11684 (N_11684,N_9572,N_7107);
or U11685 (N_11685,N_6996,N_5148);
or U11686 (N_11686,N_8466,N_6253);
and U11687 (N_11687,N_7982,N_9040);
or U11688 (N_11688,N_7875,N_6205);
and U11689 (N_11689,N_9944,N_8523);
and U11690 (N_11690,N_6285,N_6830);
nand U11691 (N_11691,N_7562,N_8489);
or U11692 (N_11692,N_8293,N_7046);
and U11693 (N_11693,N_9192,N_5248);
nand U11694 (N_11694,N_5756,N_6457);
or U11695 (N_11695,N_8304,N_8378);
nand U11696 (N_11696,N_9113,N_8669);
nor U11697 (N_11697,N_9214,N_5227);
nor U11698 (N_11698,N_7446,N_9099);
nand U11699 (N_11699,N_7424,N_6995);
and U11700 (N_11700,N_9266,N_8008);
and U11701 (N_11701,N_9254,N_5834);
and U11702 (N_11702,N_7774,N_6305);
nand U11703 (N_11703,N_7036,N_7311);
and U11704 (N_11704,N_7084,N_9339);
or U11705 (N_11705,N_8716,N_7057);
nand U11706 (N_11706,N_5592,N_7151);
and U11707 (N_11707,N_7715,N_8917);
or U11708 (N_11708,N_9409,N_5147);
nor U11709 (N_11709,N_6433,N_8031);
nand U11710 (N_11710,N_8947,N_9824);
nor U11711 (N_11711,N_7570,N_5929);
or U11712 (N_11712,N_5846,N_9277);
nand U11713 (N_11713,N_6967,N_9111);
and U11714 (N_11714,N_9127,N_8875);
and U11715 (N_11715,N_8058,N_5357);
nand U11716 (N_11716,N_5977,N_6612);
nand U11717 (N_11717,N_7010,N_7392);
or U11718 (N_11718,N_6024,N_9957);
and U11719 (N_11719,N_6809,N_6852);
nor U11720 (N_11720,N_5436,N_7237);
nand U11721 (N_11721,N_5637,N_9165);
nor U11722 (N_11722,N_6610,N_5298);
nand U11723 (N_11723,N_6096,N_5505);
or U11724 (N_11724,N_9095,N_5372);
nand U11725 (N_11725,N_7932,N_5833);
nand U11726 (N_11726,N_7128,N_7959);
or U11727 (N_11727,N_5342,N_5027);
nand U11728 (N_11728,N_9813,N_9935);
nor U11729 (N_11729,N_9528,N_7434);
nand U11730 (N_11730,N_7629,N_7557);
or U11731 (N_11731,N_9859,N_6067);
and U11732 (N_11732,N_5292,N_9176);
nor U11733 (N_11733,N_6703,N_9830);
and U11734 (N_11734,N_7939,N_6726);
and U11735 (N_11735,N_5483,N_7104);
and U11736 (N_11736,N_9395,N_7783);
and U11737 (N_11737,N_8753,N_8180);
xor U11738 (N_11738,N_8204,N_9303);
and U11739 (N_11739,N_7719,N_8718);
and U11740 (N_11740,N_8876,N_5447);
xnor U11741 (N_11741,N_5186,N_7017);
xnor U11742 (N_11742,N_6331,N_6586);
or U11743 (N_11743,N_8792,N_8902);
xor U11744 (N_11744,N_5611,N_9284);
and U11745 (N_11745,N_5404,N_6008);
or U11746 (N_11746,N_7692,N_5803);
or U11747 (N_11747,N_7985,N_5322);
nor U11748 (N_11748,N_9817,N_7632);
or U11749 (N_11749,N_6228,N_8120);
nand U11750 (N_11750,N_5852,N_8892);
or U11751 (N_11751,N_5541,N_5019);
or U11752 (N_11752,N_7768,N_8168);
nor U11753 (N_11753,N_6664,N_8937);
xor U11754 (N_11754,N_8572,N_9269);
and U11755 (N_11755,N_9191,N_7979);
nor U11756 (N_11756,N_5734,N_6823);
nand U11757 (N_11757,N_6642,N_5567);
nor U11758 (N_11758,N_6163,N_9080);
and U11759 (N_11759,N_6039,N_5972);
nor U11760 (N_11760,N_9849,N_6071);
nor U11761 (N_11761,N_8866,N_8511);
and U11762 (N_11762,N_8430,N_6314);
and U11763 (N_11763,N_8307,N_7970);
or U11764 (N_11764,N_7013,N_9716);
and U11765 (N_11765,N_5408,N_5394);
and U11766 (N_11766,N_5304,N_7900);
nor U11767 (N_11767,N_8583,N_9345);
nor U11768 (N_11768,N_8448,N_7638);
nand U11769 (N_11769,N_6387,N_7205);
nand U11770 (N_11770,N_6589,N_9161);
nor U11771 (N_11771,N_9447,N_9013);
xor U11772 (N_11772,N_5397,N_7154);
or U11773 (N_11773,N_5600,N_8818);
nand U11774 (N_11774,N_6484,N_5901);
and U11775 (N_11775,N_6426,N_9745);
and U11776 (N_11776,N_9844,N_6879);
nor U11777 (N_11777,N_9335,N_7747);
and U11778 (N_11778,N_5445,N_7929);
or U11779 (N_11779,N_7358,N_8767);
nor U11780 (N_11780,N_8190,N_8135);
or U11781 (N_11781,N_8798,N_9098);
xor U11782 (N_11782,N_5180,N_9540);
or U11783 (N_11783,N_9679,N_5591);
and U11784 (N_11784,N_5293,N_9827);
nand U11785 (N_11785,N_9887,N_6355);
nor U11786 (N_11786,N_8490,N_7915);
and U11787 (N_11787,N_7412,N_7736);
and U11788 (N_11788,N_7853,N_6685);
nor U11789 (N_11789,N_6089,N_9952);
nor U11790 (N_11790,N_9732,N_5358);
and U11791 (N_11791,N_8554,N_6005);
and U11792 (N_11792,N_9719,N_7757);
xor U11793 (N_11793,N_6215,N_5453);
and U11794 (N_11794,N_5671,N_9058);
nor U11795 (N_11795,N_5644,N_9367);
or U11796 (N_11796,N_7826,N_5297);
and U11797 (N_11797,N_5016,N_7384);
nor U11798 (N_11798,N_5773,N_5210);
xnor U11799 (N_11799,N_8657,N_6692);
nand U11800 (N_11800,N_8835,N_9588);
or U11801 (N_11801,N_5895,N_7350);
and U11802 (N_11802,N_7788,N_7320);
nor U11803 (N_11803,N_8899,N_9630);
and U11804 (N_11804,N_6842,N_5374);
and U11805 (N_11805,N_7175,N_7953);
and U11806 (N_11806,N_7635,N_5552);
nor U11807 (N_11807,N_6315,N_7364);
and U11808 (N_11808,N_9939,N_8911);
or U11809 (N_11809,N_7999,N_8919);
nor U11810 (N_11810,N_6060,N_5130);
nand U11811 (N_11811,N_9891,N_5726);
xor U11812 (N_11812,N_5968,N_6296);
nor U11813 (N_11813,N_6755,N_8439);
and U11814 (N_11814,N_8369,N_5268);
or U11815 (N_11815,N_5132,N_5416);
or U11816 (N_11816,N_5926,N_9814);
or U11817 (N_11817,N_8719,N_8982);
or U11818 (N_11818,N_7672,N_9999);
or U11819 (N_11819,N_9340,N_7754);
nor U11820 (N_11820,N_9717,N_5049);
and U11821 (N_11821,N_5819,N_8534);
nor U11822 (N_11822,N_8156,N_5230);
nor U11823 (N_11823,N_5252,N_9226);
and U11824 (N_11824,N_5385,N_8522);
nand U11825 (N_11825,N_9517,N_8833);
or U11826 (N_11826,N_9799,N_6474);
nand U11827 (N_11827,N_8167,N_8924);
nand U11828 (N_11828,N_8254,N_9250);
nand U11829 (N_11829,N_9365,N_7531);
nand U11830 (N_11830,N_9514,N_9116);
or U11831 (N_11831,N_8444,N_8843);
xnor U11832 (N_11832,N_8323,N_9130);
and U11833 (N_11833,N_5645,N_5111);
nand U11834 (N_11834,N_9584,N_5839);
nor U11835 (N_11835,N_9199,N_9293);
nor U11836 (N_11836,N_6255,N_6275);
and U11837 (N_11837,N_8604,N_9612);
nor U11838 (N_11838,N_5328,N_9234);
xor U11839 (N_11839,N_6622,N_6468);
xnor U11840 (N_11840,N_7110,N_7025);
and U11841 (N_11841,N_6431,N_7417);
and U11842 (N_11842,N_6370,N_8704);
xnor U11843 (N_11843,N_9481,N_8888);
or U11844 (N_11844,N_9349,N_5274);
and U11845 (N_11845,N_8172,N_8813);
nand U11846 (N_11846,N_6288,N_9397);
xnor U11847 (N_11847,N_5170,N_6034);
nor U11848 (N_11848,N_6416,N_6162);
nor U11849 (N_11849,N_7765,N_8253);
or U11850 (N_11850,N_8381,N_6730);
nor U11851 (N_11851,N_9669,N_8205);
and U11852 (N_11852,N_6199,N_7731);
nor U11853 (N_11853,N_7200,N_6789);
nand U11854 (N_11854,N_9047,N_6227);
nand U11855 (N_11855,N_6049,N_6635);
and U11856 (N_11856,N_6054,N_8257);
or U11857 (N_11857,N_6487,N_8925);
nand U11858 (N_11858,N_8115,N_7571);
xor U11859 (N_11859,N_9458,N_5158);
nor U11860 (N_11860,N_8385,N_8082);
or U11861 (N_11861,N_7362,N_5989);
nor U11862 (N_11862,N_9525,N_9092);
or U11863 (N_11863,N_8037,N_6829);
nor U11864 (N_11864,N_7100,N_6078);
and U11865 (N_11865,N_7284,N_9205);
and U11866 (N_11866,N_5547,N_6304);
or U11867 (N_11867,N_7689,N_9542);
and U11868 (N_11868,N_7217,N_5448);
or U11869 (N_11869,N_7620,N_5204);
xnor U11870 (N_11870,N_5434,N_7024);
xor U11871 (N_11871,N_5295,N_6934);
or U11872 (N_11872,N_6418,N_6164);
nor U11873 (N_11873,N_5318,N_5919);
xnor U11874 (N_11874,N_6392,N_9177);
and U11875 (N_11875,N_6723,N_8308);
or U11876 (N_11876,N_5348,N_5712);
or U11877 (N_11877,N_9163,N_8437);
nor U11878 (N_11878,N_8388,N_9777);
nand U11879 (N_11879,N_9289,N_9074);
and U11880 (N_11880,N_8493,N_7525);
nor U11881 (N_11881,N_7442,N_5802);
xnor U11882 (N_11882,N_5349,N_5491);
nand U11883 (N_11883,N_7167,N_6659);
nand U11884 (N_11884,N_5817,N_7968);
nand U11885 (N_11885,N_9627,N_5933);
nor U11886 (N_11886,N_6294,N_6531);
nor U11887 (N_11887,N_8630,N_6319);
nor U11888 (N_11888,N_6189,N_5615);
and U11889 (N_11889,N_6914,N_8343);
xor U11890 (N_11890,N_7353,N_9804);
and U11891 (N_11891,N_9677,N_8829);
or U11892 (N_11892,N_9175,N_7739);
or U11893 (N_11893,N_5887,N_9432);
nand U11894 (N_11894,N_9655,N_9971);
and U11895 (N_11895,N_9380,N_8900);
nor U11896 (N_11896,N_7654,N_6716);
nand U11897 (N_11897,N_7001,N_6274);
nand U11898 (N_11898,N_7479,N_6563);
nor U11899 (N_11899,N_7019,N_6763);
nor U11900 (N_11900,N_8968,N_7574);
nor U11901 (N_11901,N_6491,N_6983);
nand U11902 (N_11902,N_7278,N_5904);
nor U11903 (N_11903,N_7432,N_5107);
nor U11904 (N_11904,N_7077,N_9301);
and U11905 (N_11905,N_7879,N_7523);
and U11906 (N_11906,N_8230,N_9563);
or U11907 (N_11907,N_6644,N_7081);
nand U11908 (N_11908,N_5649,N_6009);
xnor U11909 (N_11909,N_7822,N_9706);
nor U11910 (N_11910,N_5334,N_6352);
xor U11911 (N_11911,N_6528,N_9236);
nand U11912 (N_11912,N_5794,N_5577);
nor U11913 (N_11913,N_8778,N_9393);
and U11914 (N_11914,N_8096,N_8362);
nand U11915 (N_11915,N_9396,N_7415);
or U11916 (N_11916,N_6688,N_8790);
and U11917 (N_11917,N_6258,N_6623);
nand U11918 (N_11918,N_5733,N_5361);
and U11919 (N_11919,N_6105,N_9918);
or U11920 (N_11920,N_5573,N_7239);
or U11921 (N_11921,N_8978,N_9535);
and U11922 (N_11922,N_8013,N_5630);
or U11923 (N_11923,N_6948,N_9068);
and U11924 (N_11924,N_6984,N_5666);
and U11925 (N_11925,N_8644,N_9725);
nor U11926 (N_11926,N_9470,N_6223);
xnor U11927 (N_11927,N_7954,N_9598);
or U11928 (N_11928,N_7365,N_8915);
nand U11929 (N_11929,N_6031,N_8286);
and U11930 (N_11930,N_7263,N_7213);
xnor U11931 (N_11931,N_5550,N_7555);
nor U11932 (N_11932,N_8392,N_7786);
or U11933 (N_11933,N_8820,N_8398);
and U11934 (N_11934,N_8952,N_6460);
and U11935 (N_11935,N_7653,N_5927);
nand U11936 (N_11936,N_5398,N_9608);
nand U11937 (N_11937,N_8057,N_8701);
or U11938 (N_11938,N_8494,N_9602);
nand U11939 (N_11939,N_9704,N_8158);
and U11940 (N_11940,N_6411,N_7011);
or U11941 (N_11941,N_6603,N_5197);
nand U11942 (N_11942,N_6650,N_7860);
nand U11943 (N_11943,N_5036,N_7405);
or U11944 (N_11944,N_5810,N_9228);
nand U11945 (N_11945,N_5030,N_5022);
and U11946 (N_11946,N_6575,N_9509);
xor U11947 (N_11947,N_6012,N_8584);
nand U11948 (N_11948,N_6290,N_7560);
and U11949 (N_11949,N_5008,N_8526);
nor U11950 (N_11950,N_9661,N_6545);
nand U11951 (N_11951,N_8039,N_8827);
and U11952 (N_11952,N_9455,N_6862);
nand U11953 (N_11953,N_5718,N_8200);
or U11954 (N_11954,N_8207,N_8946);
nand U11955 (N_11955,N_9970,N_5950);
nor U11956 (N_11956,N_8712,N_6043);
and U11957 (N_11957,N_5007,N_7941);
nor U11958 (N_11958,N_8566,N_5982);
xor U11959 (N_11959,N_9568,N_8847);
nand U11960 (N_11960,N_6220,N_8867);
xor U11961 (N_11961,N_5873,N_8061);
or U11962 (N_11962,N_5955,N_6853);
and U11963 (N_11963,N_6325,N_7945);
nor U11964 (N_11964,N_8776,N_5209);
and U11965 (N_11965,N_8015,N_7971);
and U11966 (N_11966,N_9848,N_5789);
xnor U11967 (N_11967,N_8916,N_7691);
nand U11968 (N_11968,N_5331,N_6372);
nor U11969 (N_11969,N_5622,N_9413);
and U11970 (N_11970,N_5407,N_6713);
nand U11971 (N_11971,N_5231,N_6679);
nand U11972 (N_11972,N_6944,N_8891);
nand U11973 (N_11973,N_5198,N_7402);
nand U11974 (N_11974,N_9319,N_7793);
or U11975 (N_11975,N_8488,N_7179);
and U11976 (N_11976,N_6150,N_5108);
nor U11977 (N_11977,N_6553,N_5797);
nand U11978 (N_11978,N_7703,N_9256);
or U11979 (N_11979,N_5504,N_6499);
and U11980 (N_11980,N_8961,N_7799);
or U11981 (N_11981,N_5943,N_7303);
and U11982 (N_11982,N_7413,N_9778);
nand U11983 (N_11983,N_6178,N_8092);
nand U11984 (N_11984,N_7051,N_5657);
nand U11985 (N_11985,N_8182,N_5804);
and U11986 (N_11986,N_7467,N_8878);
or U11987 (N_11987,N_7447,N_6340);
nor U11988 (N_11988,N_5751,N_6569);
nor U11989 (N_11989,N_8645,N_7732);
and U11990 (N_11990,N_7090,N_8441);
nor U11991 (N_11991,N_9808,N_9865);
and U11992 (N_11992,N_9958,N_5488);
or U11993 (N_11993,N_5911,N_6337);
or U11994 (N_11994,N_6311,N_8536);
nor U11995 (N_11995,N_5793,N_8201);
or U11996 (N_11996,N_9000,N_9222);
nor U11997 (N_11997,N_5761,N_9684);
and U11998 (N_11998,N_6250,N_6485);
nor U11999 (N_11999,N_6082,N_8349);
nand U12000 (N_12000,N_7639,N_5208);
nand U12001 (N_12001,N_9472,N_8346);
nor U12002 (N_12002,N_8913,N_7211);
nor U12003 (N_12003,N_5856,N_7372);
nand U12004 (N_12004,N_8011,N_5906);
and U12005 (N_12005,N_5685,N_5868);
and U12006 (N_12006,N_9010,N_5816);
xor U12007 (N_12007,N_5257,N_7701);
or U12008 (N_12008,N_8922,N_8164);
or U12009 (N_12009,N_6593,N_6638);
nand U12010 (N_12010,N_8519,N_8825);
or U12011 (N_12011,N_7710,N_5538);
and U12012 (N_12012,N_5636,N_9851);
nand U12013 (N_12013,N_6368,N_5744);
nand U12014 (N_12014,N_9558,N_9694);
or U12015 (N_12015,N_8555,N_7069);
nand U12016 (N_12016,N_5903,N_7055);
nor U12017 (N_12017,N_9593,N_7186);
or U12018 (N_12018,N_5057,N_6064);
nand U12019 (N_12019,N_5182,N_8012);
nor U12020 (N_12020,N_6536,N_7947);
nand U12021 (N_12021,N_6949,N_8176);
nand U12022 (N_12022,N_7704,N_6821);
nor U12023 (N_12023,N_9082,N_8386);
nor U12024 (N_12024,N_9054,N_8503);
or U12025 (N_12025,N_9033,N_7618);
nor U12026 (N_12026,N_5441,N_7758);
and U12027 (N_12027,N_6134,N_8471);
nor U12028 (N_12028,N_7622,N_6373);
and U12029 (N_12029,N_9162,N_9118);
or U12030 (N_12030,N_8108,N_5135);
and U12031 (N_12031,N_6119,N_9578);
nand U12032 (N_12032,N_7489,N_5092);
nand U12033 (N_12033,N_8358,N_8885);
and U12034 (N_12034,N_6302,N_8616);
and U12035 (N_12035,N_7983,N_6213);
nor U12036 (N_12036,N_7633,N_6972);
and U12037 (N_12037,N_6869,N_7007);
and U12038 (N_12038,N_8673,N_9089);
nand U12039 (N_12039,N_6732,N_6661);
nor U12040 (N_12040,N_5674,N_9993);
nor U12041 (N_12041,N_9606,N_8508);
or U12042 (N_12042,N_9667,N_7188);
and U12043 (N_12043,N_9863,N_5495);
nor U12044 (N_12044,N_9039,N_9734);
xor U12045 (N_12045,N_7675,N_7830);
or U12046 (N_12046,N_9783,N_9488);
and U12047 (N_12047,N_9037,N_7317);
or U12048 (N_12048,N_6510,N_5691);
nor U12049 (N_12049,N_9533,N_6945);
and U12050 (N_12050,N_8146,N_8305);
or U12051 (N_12051,N_7984,N_7975);
nand U12052 (N_12052,N_8113,N_8641);
or U12053 (N_12053,N_7711,N_5389);
nor U12054 (N_12054,N_7825,N_6844);
nor U12055 (N_12055,N_8213,N_7741);
or U12056 (N_12056,N_9815,N_6601);
and U12057 (N_12057,N_9135,N_6020);
nor U12058 (N_12058,N_5164,N_7487);
nand U12059 (N_12059,N_9117,N_9194);
and U12060 (N_12060,N_5275,N_9173);
nand U12061 (N_12061,N_5608,N_5421);
nor U12062 (N_12062,N_9248,N_6463);
nand U12063 (N_12063,N_8003,N_5606);
nand U12064 (N_12064,N_7095,N_9422);
or U12065 (N_12065,N_5351,N_5562);
nand U12066 (N_12066,N_8191,N_8417);
xnor U12067 (N_12067,N_5427,N_7619);
and U12068 (N_12068,N_6698,N_6229);
xor U12069 (N_12069,N_9056,N_7894);
and U12070 (N_12070,N_7581,N_8632);
xnor U12071 (N_12071,N_7794,N_8890);
or U12072 (N_12072,N_8856,N_6971);
or U12073 (N_12073,N_9114,N_7775);
and U12074 (N_12074,N_6618,N_8094);
or U12075 (N_12075,N_5779,N_6824);
and U12076 (N_12076,N_9083,N_8521);
and U12077 (N_12077,N_6473,N_8166);
xnor U12078 (N_12078,N_6939,N_6407);
nand U12079 (N_12079,N_5569,N_8731);
and U12080 (N_12080,N_5886,N_7026);
nand U12081 (N_12081,N_6673,N_8810);
or U12082 (N_12082,N_6158,N_8150);
or U12083 (N_12083,N_8070,N_6084);
and U12084 (N_12084,N_8631,N_6621);
xnor U12085 (N_12085,N_7888,N_5759);
nor U12086 (N_12086,N_6332,N_8063);
and U12087 (N_12087,N_9973,N_6901);
and U12088 (N_12088,N_6100,N_8588);
and U12089 (N_12089,N_9357,N_6023);
and U12090 (N_12090,N_7804,N_9336);
nor U12091 (N_12091,N_5353,N_7682);
xnor U12092 (N_12092,N_5341,N_6056);
xor U12093 (N_12093,N_9499,N_6604);
nand U12094 (N_12094,N_9502,N_6087);
xor U12095 (N_12095,N_5882,N_5889);
and U12096 (N_12096,N_5324,N_8971);
nand U12097 (N_12097,N_8072,N_6722);
or U12098 (N_12098,N_9036,N_8317);
or U12099 (N_12099,N_9446,N_9112);
and U12100 (N_12100,N_8528,N_8552);
and U12101 (N_12101,N_9486,N_8449);
nor U12102 (N_12102,N_8465,N_8787);
or U12103 (N_12103,N_9026,N_9826);
or U12104 (N_12104,N_6410,N_5680);
or U12105 (N_12105,N_6263,N_5753);
xnor U12106 (N_12106,N_5065,N_6058);
or U12107 (N_12107,N_5480,N_5639);
nand U12108 (N_12108,N_7433,N_6212);
nor U12109 (N_12109,N_5481,N_9350);
xnor U12110 (N_12110,N_8093,N_8252);
nor U12111 (N_12111,N_8839,N_8097);
nand U12112 (N_12112,N_9647,N_9556);
and U12113 (N_12113,N_8076,N_8474);
nor U12114 (N_12114,N_8139,N_5584);
xor U12115 (N_12115,N_7728,N_8926);
xnor U12116 (N_12116,N_9837,N_9085);
or U12117 (N_12117,N_9780,N_8903);
nand U12118 (N_12118,N_7606,N_9291);
and U12119 (N_12119,N_9415,N_6951);
and U12120 (N_12120,N_8342,N_5628);
or U12121 (N_12121,N_5741,N_5258);
or U12122 (N_12122,N_5069,N_6794);
and U12123 (N_12123,N_5020,N_6560);
or U12124 (N_12124,N_7150,N_6313);
or U12125 (N_12125,N_8291,N_8995);
or U12126 (N_12126,N_8056,N_7813);
nand U12127 (N_12127,N_5934,N_9389);
or U12128 (N_12128,N_5946,N_6920);
nand U12129 (N_12129,N_6367,N_5993);
xor U12130 (N_12130,N_5770,N_7700);
or U12131 (N_12131,N_7918,N_6700);
nor U12132 (N_12132,N_5878,N_9077);
or U12133 (N_12133,N_7374,N_5590);
or U12134 (N_12134,N_6280,N_6702);
nand U12135 (N_12135,N_6833,N_5465);
or U12136 (N_12136,N_8377,N_6909);
nand U12137 (N_12137,N_6477,N_7912);
nand U12138 (N_12138,N_5171,N_5785);
or U12139 (N_12139,N_9786,N_5660);
nand U12140 (N_12140,N_6282,N_6771);
or U12141 (N_12141,N_5192,N_8268);
nor U12142 (N_12142,N_6981,N_5200);
and U12143 (N_12143,N_9708,N_8981);
or U12144 (N_12144,N_6497,N_6256);
nor U12145 (N_12145,N_7304,N_6384);
nor U12146 (N_12146,N_8543,N_7834);
and U12147 (N_12147,N_9790,N_7120);
and U12148 (N_12148,N_9855,N_7266);
xor U12149 (N_12149,N_9586,N_9690);
or U12150 (N_12150,N_6765,N_7341);
nand U12151 (N_12151,N_9246,N_9549);
nand U12152 (N_12152,N_9974,N_6834);
or U12153 (N_12153,N_9354,N_7922);
or U12154 (N_12154,N_9645,N_7256);
or U12155 (N_12155,N_5710,N_8939);
nand U12156 (N_12156,N_7930,N_7881);
nor U12157 (N_12157,N_8697,N_9378);
nor U12158 (N_12158,N_8144,N_9210);
xor U12159 (N_12159,N_7207,N_9668);
xor U12160 (N_12160,N_8551,N_6599);
xnor U12161 (N_12161,N_7485,N_9736);
and U12162 (N_12162,N_8759,N_7450);
nand U12163 (N_12163,N_5405,N_9091);
nand U12164 (N_12164,N_8371,N_5716);
and U12165 (N_12165,N_9875,N_8877);
and U12166 (N_12166,N_5395,N_9843);
nand U12167 (N_12167,N_6015,N_5144);
nand U12168 (N_12168,N_7118,N_5953);
nor U12169 (N_12169,N_9980,N_9788);
nand U12170 (N_12170,N_5589,N_7906);
and U12171 (N_12171,N_6287,N_7156);
and U12172 (N_12172,N_8779,N_8722);
or U12173 (N_12173,N_6872,N_9428);
nor U12174 (N_12174,N_5844,N_9122);
or U12175 (N_12175,N_6714,N_6226);
or U12176 (N_12176,N_8930,N_9738);
xor U12177 (N_12177,N_6561,N_8382);
nor U12178 (N_12178,N_5039,N_9362);
nand U12179 (N_12179,N_5206,N_6455);
or U12180 (N_12180,N_5202,N_5822);
and U12181 (N_12181,N_6508,N_7219);
nand U12182 (N_12182,N_6556,N_5863);
nand U12183 (N_12183,N_8879,N_5635);
nand U12184 (N_12184,N_9174,N_7662);
xor U12185 (N_12185,N_5466,N_9609);
or U12186 (N_12186,N_5474,N_5788);
and U12187 (N_12187,N_7884,N_8881);
nand U12188 (N_12188,N_8777,N_8473);
or U12189 (N_12189,N_6161,N_5891);
nand U12190 (N_12190,N_7996,N_9338);
nand U12191 (N_12191,N_9501,N_5250);
or U12192 (N_12192,N_8889,N_7518);
xnor U12193 (N_12193,N_5544,N_6633);
xnor U12194 (N_12194,N_7313,N_5786);
xor U12195 (N_12195,N_7422,N_8991);
nor U12196 (N_12196,N_9134,N_5460);
nand U12197 (N_12197,N_6519,N_7449);
xnor U12198 (N_12198,N_8633,N_6978);
or U12199 (N_12199,N_8005,N_6097);
or U12200 (N_12200,N_6941,N_5081);
or U12201 (N_12201,N_6238,N_9954);
and U12202 (N_12202,N_6709,N_6144);
xnor U12203 (N_12203,N_6117,N_6764);
or U12204 (N_12204,N_6121,N_6815);
or U12205 (N_12205,N_6915,N_9055);
or U12206 (N_12206,N_8807,N_8007);
or U12207 (N_12207,N_7354,N_7767);
nor U12208 (N_12208,N_9243,N_7381);
or U12209 (N_12209,N_8032,N_9785);
nand U12210 (N_12210,N_5110,N_8724);
and U12211 (N_12211,N_6727,N_7600);
nand U12212 (N_12212,N_7552,N_9383);
and U12213 (N_12213,N_7551,N_7522);
and U12214 (N_12214,N_8030,N_6999);
nand U12215 (N_12215,N_6249,N_5827);
nand U12216 (N_12216,N_8629,N_9439);
or U12217 (N_12217,N_5433,N_9480);
nor U12218 (N_12218,N_6718,N_5193);
and U12219 (N_12219,N_8303,N_6371);
xnor U12220 (N_12220,N_6334,N_8142);
nand U12221 (N_12221,N_5689,N_7021);
nand U12222 (N_12222,N_9090,N_6896);
or U12223 (N_12223,N_5450,N_5190);
or U12224 (N_12224,N_5705,N_6002);
or U12225 (N_12225,N_9104,N_7986);
nand U12226 (N_12226,N_7171,N_9659);
or U12227 (N_12227,N_9551,N_6069);
nor U12228 (N_12228,N_6772,N_9964);
or U12229 (N_12229,N_9820,N_7746);
nor U12230 (N_12230,N_6807,N_9202);
or U12231 (N_12231,N_9450,N_8262);
nor U12232 (N_12232,N_6979,N_6466);
xor U12233 (N_12233,N_5472,N_7677);
nor U12234 (N_12234,N_8853,N_9746);
or U12235 (N_12235,N_5910,N_6591);
and U12236 (N_12236,N_5096,N_7031);
nand U12237 (N_12237,N_7738,N_8043);
xnor U12238 (N_12238,N_7988,N_9571);
or U12239 (N_12239,N_6810,N_9570);
nor U12240 (N_12240,N_9538,N_6420);
nand U12241 (N_12241,N_9628,N_7801);
nand U12242 (N_12242,N_5048,N_6752);
or U12243 (N_12243,N_7098,N_6875);
nor U12244 (N_12244,N_5125,N_8990);
and U12245 (N_12245,N_6265,N_7991);
xnor U12246 (N_12246,N_7990,N_7616);
and U12247 (N_12247,N_7260,N_5732);
or U12248 (N_12248,N_9315,N_7512);
and U12249 (N_12249,N_8796,N_5050);
nor U12250 (N_12250,N_9925,N_5265);
nand U12251 (N_12251,N_9917,N_7723);
and U12252 (N_12252,N_9519,N_5014);
or U12253 (N_12253,N_6174,N_6404);
nor U12254 (N_12254,N_6299,N_6677);
nor U12255 (N_12255,N_5188,N_9959);
or U12256 (N_12256,N_5517,N_7438);
and U12257 (N_12257,N_9864,N_5001);
xnor U12258 (N_12258,N_9587,N_7781);
xnor U12259 (N_12259,N_9463,N_5825);
and U12260 (N_12260,N_8472,N_6488);
and U12261 (N_12261,N_9526,N_7855);
or U12262 (N_12262,N_5012,N_5479);
and U12263 (N_12263,N_5439,N_9924);
nand U12264 (N_12264,N_7086,N_9298);
nand U12265 (N_12265,N_9564,N_7199);
nor U12266 (N_12266,N_5912,N_5616);
and U12267 (N_12267,N_5343,N_5068);
nand U12268 (N_12268,N_6001,N_9045);
nor U12269 (N_12269,N_6615,N_9835);
nor U12270 (N_12270,N_5018,N_7136);
and U12271 (N_12271,N_8319,N_7116);
nand U12272 (N_12272,N_6573,N_8160);
nor U12273 (N_12273,N_5305,N_5160);
and U12274 (N_12274,N_9703,N_9473);
or U12275 (N_12275,N_8054,N_7743);
nor U12276 (N_12276,N_8525,N_5211);
xnor U12277 (N_12277,N_8455,N_8079);
nor U12278 (N_12278,N_5187,N_6246);
nand U12279 (N_12279,N_8772,N_8374);
nand U12280 (N_12280,N_6086,N_5564);
or U12281 (N_12281,N_9643,N_5633);
nor U12282 (N_12282,N_5320,N_5563);
and U12283 (N_12283,N_8539,N_9049);
and U12284 (N_12284,N_9847,N_5986);
and U12285 (N_12285,N_6784,N_8510);
nor U12286 (N_12286,N_7938,N_7112);
nor U12287 (N_12287,N_8987,N_8652);
nor U12288 (N_12288,N_6530,N_6847);
and U12289 (N_12289,N_7994,N_8046);
or U12290 (N_12290,N_6366,N_5486);
and U12291 (N_12291,N_7992,N_5136);
or U12292 (N_12292,N_5363,N_8436);
and U12293 (N_12293,N_8953,N_8625);
and U12294 (N_12294,N_5648,N_6985);
nand U12295 (N_12295,N_5815,N_8122);
nand U12296 (N_12296,N_9537,N_8277);
and U12297 (N_12297,N_9948,N_8413);
or U12298 (N_12298,N_6080,N_5961);
and U12299 (N_12299,N_7041,N_6131);
nor U12300 (N_12300,N_8199,N_9831);
nand U12301 (N_12301,N_9543,N_6283);
nor U12302 (N_12302,N_7787,N_6758);
and U12303 (N_12303,N_5593,N_8688);
nand U12304 (N_12304,N_9015,N_8784);
and U12305 (N_12305,N_6098,N_5975);
nand U12306 (N_12306,N_6339,N_5042);
nor U12307 (N_12307,N_9211,N_8433);
or U12308 (N_12308,N_7780,N_7872);
and U12309 (N_12309,N_9922,N_7847);
and U12310 (N_12310,N_6347,N_8234);
nor U12311 (N_12311,N_9050,N_9895);
and U12312 (N_12312,N_8169,N_6857);
nor U12313 (N_12313,N_5246,N_8678);
nor U12314 (N_12314,N_8869,N_7265);
xnor U12315 (N_12315,N_7656,N_7501);
nand U12316 (N_12316,N_5893,N_6974);
nand U12317 (N_12317,N_5847,N_5464);
nor U12318 (N_12318,N_8114,N_7651);
and U12319 (N_12319,N_5347,N_6577);
nand U12320 (N_12320,N_6118,N_6448);
or U12321 (N_12321,N_7508,N_5043);
nand U12322 (N_12322,N_5806,N_9281);
or U12323 (N_12323,N_5045,N_7407);
nand U12324 (N_12324,N_7264,N_8943);
or U12325 (N_12325,N_9320,N_9581);
nand U12326 (N_12326,N_5866,N_5987);
nor U12327 (N_12327,N_6027,N_7445);
and U12328 (N_12328,N_6858,N_6554);
and U12329 (N_12329,N_6309,N_6394);
nor U12330 (N_12330,N_8373,N_8487);
xnor U12331 (N_12331,N_5002,N_5249);
or U12332 (N_12332,N_6066,N_8429);
nand U12333 (N_12333,N_8340,N_6447);
nand U12334 (N_12334,N_8606,N_5139);
and U12335 (N_12335,N_5583,N_6273);
or U12336 (N_12336,N_9794,N_5976);
nand U12337 (N_12337,N_9906,N_5417);
and U12338 (N_12338,N_9981,N_6503);
nand U12339 (N_12339,N_5294,N_5475);
and U12340 (N_12340,N_5037,N_5338);
xnor U12341 (N_12341,N_8914,N_9823);
nor U12342 (N_12342,N_8690,N_5174);
nand U12343 (N_12343,N_8165,N_8580);
nand U12344 (N_12344,N_5728,N_5931);
nor U12345 (N_12345,N_6382,N_5023);
or U12346 (N_12346,N_9227,N_8942);
or U12347 (N_12347,N_6921,N_6476);
nor U12348 (N_12348,N_7391,N_8409);
nor U12349 (N_12349,N_6103,N_8794);
and U12350 (N_12350,N_9709,N_7085);
or U12351 (N_12351,N_8302,N_8178);
nand U12352 (N_12352,N_7376,N_7631);
nand U12353 (N_12353,N_5196,N_9759);
xor U12354 (N_12354,N_8401,N_6850);
or U12355 (N_12355,N_5694,N_8100);
xor U12356 (N_12356,N_8932,N_7664);
nor U12357 (N_12357,N_9953,N_7375);
or U12358 (N_12358,N_7798,N_5199);
or U12359 (N_12359,N_9172,N_8368);
or U12360 (N_12360,N_7942,N_6570);
nor U12361 (N_12361,N_5704,N_5127);
and U12362 (N_12362,N_6568,N_8073);
nand U12363 (N_12363,N_5017,N_6359);
nor U12364 (N_12364,N_8648,N_9764);
and U12365 (N_12365,N_6013,N_9607);
and U12366 (N_12366,N_8512,N_8162);
and U12367 (N_12367,N_8803,N_9589);
nor U12368 (N_12368,N_8959,N_8748);
nor U12369 (N_12369,N_5994,N_8231);
xnor U12370 (N_12370,N_5601,N_7296);
nand U12371 (N_12371,N_9217,N_9757);
nand U12372 (N_12372,N_7676,N_8337);
or U12373 (N_12373,N_7393,N_6184);
or U12374 (N_12374,N_9763,N_9923);
nand U12375 (N_12375,N_8289,N_9313);
and U12376 (N_12376,N_6693,N_6438);
and U12377 (N_12377,N_8446,N_9994);
nand U12378 (N_12378,N_8116,N_5145);
and U12379 (N_12379,N_9829,N_8626);
nand U12380 (N_12380,N_7863,N_6636);
and U12381 (N_12381,N_9685,N_9079);
and U12382 (N_12382,N_6676,N_8324);
nand U12383 (N_12383,N_7192,N_5858);
or U12384 (N_12384,N_7404,N_8467);
nor U12385 (N_12385,N_5865,N_7003);
nand U12386 (N_12386,N_7846,N_9258);
and U12387 (N_12387,N_6389,N_5214);
and U12388 (N_12388,N_6198,N_9772);
and U12389 (N_12389,N_5871,N_7603);
nand U12390 (N_12390,N_6825,N_6160);
nand U12391 (N_12391,N_5650,N_6652);
or U12392 (N_12392,N_6907,N_6277);
nand U12393 (N_12393,N_5229,N_9789);
nor U12394 (N_12394,N_6841,N_5917);
nand U12395 (N_12395,N_5251,N_5930);
nand U12396 (N_12396,N_7269,N_7492);
and U12397 (N_12397,N_9699,N_9937);
or U12398 (N_12398,N_8272,N_8266);
nor U12399 (N_12399,N_7468,N_8469);
nor U12400 (N_12400,N_6157,N_6234);
nand U12401 (N_12401,N_8714,N_6818);
nor U12402 (N_12402,N_9171,N_5114);
nand U12403 (N_12403,N_5423,N_9930);
nand U12404 (N_12404,N_6597,N_7349);
and U12405 (N_12405,N_7513,N_7125);
nand U12406 (N_12406,N_5537,N_5165);
nand U12407 (N_12407,N_7366,N_7709);
or U12408 (N_12408,N_5271,N_7956);
and U12409 (N_12409,N_5928,N_9181);
or U12410 (N_12410,N_7871,N_6980);
or U12411 (N_12411,N_9955,N_6936);
and U12412 (N_12412,N_8619,N_7782);
nor U12413 (N_12413,N_9363,N_9371);
and U12414 (N_12414,N_5984,N_7224);
nor U12415 (N_12415,N_8486,N_7705);
nand U12416 (N_12416,N_7791,N_5352);
nand U12417 (N_12417,N_5269,N_7844);
or U12418 (N_12418,N_8944,N_7589);
nor U12419 (N_12419,N_7360,N_8416);
or U12420 (N_12420,N_8715,N_7398);
and U12421 (N_12421,N_5598,N_9244);
and U12422 (N_12422,N_7921,N_7976);
nand U12423 (N_12423,N_8129,N_8218);
nand U12424 (N_12424,N_5477,N_9119);
or U12425 (N_12425,N_8970,N_6840);
nor U12426 (N_12426,N_8161,N_8802);
nand U12427 (N_12427,N_8174,N_7190);
nand U12428 (N_12428,N_6820,N_8153);
nor U12429 (N_12429,N_7028,N_7673);
nand U12430 (N_12430,N_8535,N_5717);
xnor U12431 (N_12431,N_5240,N_5369);
nor U12432 (N_12432,N_8010,N_6798);
and U12433 (N_12433,N_5678,N_9060);
nand U12434 (N_12434,N_6682,N_6649);
and U12435 (N_12435,N_7157,N_6190);
nand U12436 (N_12436,N_8428,N_7592);
and U12437 (N_12437,N_9445,N_8933);
or U12438 (N_12438,N_5690,N_5011);
nand U12439 (N_12439,N_6268,N_9051);
xor U12440 (N_12440,N_9883,N_5191);
or U12441 (N_12441,N_6115,N_7121);
or U12442 (N_12442,N_5875,N_5129);
and U12443 (N_12443,N_6617,N_8693);
nor U12444 (N_12444,N_5429,N_6864);
nand U12445 (N_12445,N_8828,N_5413);
or U12446 (N_12446,N_9143,N_5189);
or U12447 (N_12447,N_9620,N_7004);
and U12448 (N_12448,N_8561,N_9877);
nor U12449 (N_12449,N_5393,N_7089);
xor U12450 (N_12450,N_7062,N_8661);
and U12451 (N_12451,N_7800,N_8086);
nand U12452 (N_12452,N_7257,N_6851);
or U12453 (N_12453,N_6195,N_9418);
nand U12454 (N_12454,N_8710,N_8309);
nor U12455 (N_12455,N_8499,N_9900);
and U12456 (N_12456,N_5233,N_7696);
xnor U12457 (N_12457,N_5302,N_7177);
nor U12458 (N_12458,N_7201,N_9164);
nand U12459 (N_12459,N_8422,N_7546);
or U12460 (N_12460,N_9208,N_6379);
nor U12461 (N_12461,N_5769,N_7752);
or U12462 (N_12462,N_8117,N_8188);
and U12463 (N_12463,N_5469,N_6813);
and U12464 (N_12464,N_9781,N_6183);
and U12465 (N_12465,N_9252,N_7901);
or U12466 (N_12466,N_5898,N_5556);
and U12467 (N_12467,N_5805,N_5217);
nand U12468 (N_12468,N_7255,N_9989);
nand U12469 (N_12469,N_6811,N_8044);
or U12470 (N_12470,N_8717,N_7773);
and U12471 (N_12471,N_6092,N_6363);
or U12472 (N_12472,N_7718,N_8424);
or U12473 (N_12473,N_8615,N_5539);
nor U12474 (N_12474,N_5941,N_9215);
nor U12475 (N_12475,N_9961,N_7961);
or U12476 (N_12476,N_7301,N_6414);
and U12477 (N_12477,N_8547,N_6365);
or U12478 (N_12478,N_5409,N_5379);
nor U12479 (N_12479,N_6357,N_7623);
or U12480 (N_12480,N_8220,N_5090);
or U12481 (N_12481,N_6775,N_8019);
and U12482 (N_12482,N_8085,N_9755);
nor U12483 (N_12483,N_6744,N_6328);
xnor U12484 (N_12484,N_5499,N_8219);
nor U12485 (N_12485,N_9431,N_5207);
nor U12486 (N_12486,N_8756,N_5330);
or U12487 (N_12487,N_5181,N_7670);
and U12488 (N_12488,N_9145,N_5112);
nor U12489 (N_12489,N_7755,N_9867);
nand U12490 (N_12490,N_8713,N_9560);
nor U12491 (N_12491,N_9471,N_9966);
and U12492 (N_12492,N_7030,N_5729);
nor U12493 (N_12493,N_5640,N_6444);
nor U12494 (N_12494,N_8700,N_9665);
or U12495 (N_12495,N_6550,N_7197);
and U12496 (N_12496,N_6467,N_7385);
nand U12497 (N_12497,N_6219,N_8537);
nor U12498 (N_12498,N_9765,N_9920);
and U12499 (N_12499,N_6671,N_9187);
nand U12500 (N_12500,N_8678,N_7390);
or U12501 (N_12501,N_5036,N_8346);
and U12502 (N_12502,N_8075,N_7038);
nand U12503 (N_12503,N_9176,N_7082);
and U12504 (N_12504,N_9555,N_8101);
xor U12505 (N_12505,N_8047,N_7367);
nor U12506 (N_12506,N_7967,N_6935);
xor U12507 (N_12507,N_7513,N_8209);
nand U12508 (N_12508,N_9578,N_8369);
or U12509 (N_12509,N_7283,N_9591);
or U12510 (N_12510,N_5263,N_9941);
nand U12511 (N_12511,N_9225,N_8363);
nor U12512 (N_12512,N_9758,N_6036);
nand U12513 (N_12513,N_6373,N_7758);
nor U12514 (N_12514,N_7247,N_9617);
nand U12515 (N_12515,N_8842,N_7244);
nand U12516 (N_12516,N_6032,N_5717);
nor U12517 (N_12517,N_7368,N_5218);
xnor U12518 (N_12518,N_9699,N_6235);
nand U12519 (N_12519,N_9527,N_5055);
nand U12520 (N_12520,N_9950,N_5773);
nor U12521 (N_12521,N_7852,N_8993);
xor U12522 (N_12522,N_8068,N_7814);
xnor U12523 (N_12523,N_8776,N_9429);
nor U12524 (N_12524,N_6903,N_6002);
or U12525 (N_12525,N_9778,N_5425);
nor U12526 (N_12526,N_8427,N_6284);
nand U12527 (N_12527,N_8061,N_9281);
nor U12528 (N_12528,N_9672,N_9777);
or U12529 (N_12529,N_9089,N_9658);
or U12530 (N_12530,N_6704,N_9590);
and U12531 (N_12531,N_6829,N_7267);
and U12532 (N_12532,N_5534,N_8760);
xnor U12533 (N_12533,N_7126,N_8782);
nand U12534 (N_12534,N_5267,N_9304);
nor U12535 (N_12535,N_9650,N_9845);
nor U12536 (N_12536,N_7106,N_9334);
and U12537 (N_12537,N_9072,N_7360);
nor U12538 (N_12538,N_7069,N_7122);
or U12539 (N_12539,N_8750,N_6245);
or U12540 (N_12540,N_7018,N_6769);
nand U12541 (N_12541,N_8955,N_5079);
nor U12542 (N_12542,N_9091,N_5198);
or U12543 (N_12543,N_7947,N_6655);
nand U12544 (N_12544,N_6117,N_7065);
or U12545 (N_12545,N_9651,N_7316);
nand U12546 (N_12546,N_6679,N_7058);
and U12547 (N_12547,N_5267,N_5325);
or U12548 (N_12548,N_8091,N_7113);
and U12549 (N_12549,N_5156,N_9342);
nand U12550 (N_12550,N_6883,N_8763);
nor U12551 (N_12551,N_5658,N_9804);
nand U12552 (N_12552,N_5128,N_6937);
nor U12553 (N_12553,N_7690,N_7045);
nand U12554 (N_12554,N_7503,N_8078);
and U12555 (N_12555,N_5995,N_9033);
nand U12556 (N_12556,N_9938,N_6339);
nand U12557 (N_12557,N_6375,N_8433);
and U12558 (N_12558,N_7468,N_5554);
nor U12559 (N_12559,N_5234,N_9142);
and U12560 (N_12560,N_8678,N_9066);
or U12561 (N_12561,N_9092,N_5669);
or U12562 (N_12562,N_6124,N_7265);
nor U12563 (N_12563,N_7269,N_8941);
nor U12564 (N_12564,N_7769,N_8702);
or U12565 (N_12565,N_5445,N_6345);
or U12566 (N_12566,N_9651,N_5403);
and U12567 (N_12567,N_7334,N_8556);
nand U12568 (N_12568,N_6697,N_7266);
nand U12569 (N_12569,N_8107,N_9460);
xnor U12570 (N_12570,N_6333,N_6776);
and U12571 (N_12571,N_6680,N_5152);
nand U12572 (N_12572,N_5671,N_6902);
xor U12573 (N_12573,N_7037,N_9911);
xnor U12574 (N_12574,N_8628,N_7598);
nand U12575 (N_12575,N_7287,N_9518);
or U12576 (N_12576,N_8263,N_8358);
nor U12577 (N_12577,N_5008,N_6983);
nand U12578 (N_12578,N_6035,N_8463);
and U12579 (N_12579,N_8097,N_5273);
or U12580 (N_12580,N_7916,N_5105);
nand U12581 (N_12581,N_7471,N_5385);
xnor U12582 (N_12582,N_7069,N_8230);
nand U12583 (N_12583,N_7312,N_8001);
and U12584 (N_12584,N_5847,N_9224);
and U12585 (N_12585,N_7632,N_9835);
nor U12586 (N_12586,N_9309,N_8699);
nand U12587 (N_12587,N_9121,N_8464);
xor U12588 (N_12588,N_8677,N_5431);
and U12589 (N_12589,N_6437,N_7335);
nor U12590 (N_12590,N_5368,N_7570);
nand U12591 (N_12591,N_5585,N_5968);
or U12592 (N_12592,N_7448,N_6485);
nand U12593 (N_12593,N_5752,N_6911);
or U12594 (N_12594,N_7814,N_5186);
xnor U12595 (N_12595,N_8341,N_9263);
or U12596 (N_12596,N_7238,N_6718);
and U12597 (N_12597,N_9743,N_9444);
and U12598 (N_12598,N_6945,N_8758);
and U12599 (N_12599,N_7469,N_7156);
nand U12600 (N_12600,N_6302,N_5058);
nand U12601 (N_12601,N_7421,N_8518);
nor U12602 (N_12602,N_8330,N_5954);
or U12603 (N_12603,N_6997,N_5615);
nor U12604 (N_12604,N_5124,N_9943);
nand U12605 (N_12605,N_9317,N_8085);
xnor U12606 (N_12606,N_9668,N_7908);
nand U12607 (N_12607,N_5302,N_9742);
or U12608 (N_12608,N_6553,N_8601);
or U12609 (N_12609,N_9510,N_7749);
xnor U12610 (N_12610,N_7851,N_8484);
or U12611 (N_12611,N_9067,N_8609);
nand U12612 (N_12612,N_5036,N_5196);
nand U12613 (N_12613,N_9827,N_5891);
or U12614 (N_12614,N_8069,N_8197);
or U12615 (N_12615,N_8400,N_7303);
or U12616 (N_12616,N_6349,N_9083);
nor U12617 (N_12617,N_7307,N_7407);
and U12618 (N_12618,N_8870,N_9323);
and U12619 (N_12619,N_7151,N_8465);
and U12620 (N_12620,N_8216,N_6595);
nor U12621 (N_12621,N_7984,N_8439);
nor U12622 (N_12622,N_8083,N_5951);
nor U12623 (N_12623,N_8982,N_9502);
nand U12624 (N_12624,N_6359,N_5550);
nand U12625 (N_12625,N_8630,N_6069);
nor U12626 (N_12626,N_5426,N_6772);
nor U12627 (N_12627,N_8065,N_8932);
nor U12628 (N_12628,N_8188,N_8885);
nand U12629 (N_12629,N_7223,N_8396);
nand U12630 (N_12630,N_9300,N_5563);
nand U12631 (N_12631,N_7881,N_7629);
nor U12632 (N_12632,N_9575,N_6695);
nand U12633 (N_12633,N_5240,N_6691);
nor U12634 (N_12634,N_6166,N_8722);
nor U12635 (N_12635,N_7008,N_9446);
nor U12636 (N_12636,N_6974,N_6060);
and U12637 (N_12637,N_8576,N_9469);
nand U12638 (N_12638,N_5207,N_6593);
or U12639 (N_12639,N_5354,N_5138);
xnor U12640 (N_12640,N_8349,N_6580);
or U12641 (N_12641,N_6127,N_7364);
or U12642 (N_12642,N_8764,N_5851);
and U12643 (N_12643,N_8374,N_6984);
nor U12644 (N_12644,N_7235,N_7174);
nand U12645 (N_12645,N_9552,N_9381);
or U12646 (N_12646,N_7579,N_6343);
or U12647 (N_12647,N_9698,N_9741);
or U12648 (N_12648,N_5024,N_8949);
and U12649 (N_12649,N_5810,N_8067);
xor U12650 (N_12650,N_9420,N_6179);
nand U12651 (N_12651,N_8675,N_6274);
nor U12652 (N_12652,N_8002,N_5014);
nor U12653 (N_12653,N_8793,N_7472);
nand U12654 (N_12654,N_5078,N_5767);
or U12655 (N_12655,N_8523,N_5773);
xor U12656 (N_12656,N_7597,N_5146);
nand U12657 (N_12657,N_6413,N_9704);
and U12658 (N_12658,N_8227,N_5463);
nor U12659 (N_12659,N_5362,N_9218);
and U12660 (N_12660,N_6040,N_5560);
nor U12661 (N_12661,N_8648,N_6719);
nor U12662 (N_12662,N_8752,N_7633);
nand U12663 (N_12663,N_5469,N_9716);
nand U12664 (N_12664,N_5442,N_6768);
or U12665 (N_12665,N_7277,N_6212);
or U12666 (N_12666,N_6483,N_8362);
and U12667 (N_12667,N_7514,N_7245);
or U12668 (N_12668,N_7552,N_7716);
xnor U12669 (N_12669,N_7289,N_5990);
nand U12670 (N_12670,N_8712,N_9331);
or U12671 (N_12671,N_8745,N_6147);
and U12672 (N_12672,N_6391,N_6684);
nor U12673 (N_12673,N_7353,N_9893);
nand U12674 (N_12674,N_6625,N_7165);
nor U12675 (N_12675,N_9848,N_8175);
nor U12676 (N_12676,N_7734,N_6160);
nand U12677 (N_12677,N_9723,N_8164);
nand U12678 (N_12678,N_9368,N_9806);
and U12679 (N_12679,N_5507,N_7532);
xor U12680 (N_12680,N_9327,N_8710);
nand U12681 (N_12681,N_6927,N_8805);
and U12682 (N_12682,N_8630,N_8716);
nand U12683 (N_12683,N_8817,N_8839);
xnor U12684 (N_12684,N_9102,N_7148);
or U12685 (N_12685,N_9705,N_7892);
xnor U12686 (N_12686,N_9371,N_5623);
xor U12687 (N_12687,N_9580,N_5149);
nand U12688 (N_12688,N_9146,N_9199);
nand U12689 (N_12689,N_5576,N_7066);
and U12690 (N_12690,N_7402,N_8185);
xnor U12691 (N_12691,N_5122,N_7428);
or U12692 (N_12692,N_9063,N_6052);
or U12693 (N_12693,N_9849,N_5626);
nor U12694 (N_12694,N_5777,N_6218);
nand U12695 (N_12695,N_9160,N_5479);
and U12696 (N_12696,N_7807,N_6252);
nor U12697 (N_12697,N_9555,N_8651);
nor U12698 (N_12698,N_6844,N_9777);
or U12699 (N_12699,N_6009,N_5707);
nor U12700 (N_12700,N_8033,N_9721);
nand U12701 (N_12701,N_8516,N_7039);
nor U12702 (N_12702,N_8921,N_7151);
xor U12703 (N_12703,N_6988,N_8152);
nor U12704 (N_12704,N_9566,N_5474);
and U12705 (N_12705,N_7532,N_6724);
and U12706 (N_12706,N_6773,N_5396);
nand U12707 (N_12707,N_6846,N_8056);
nor U12708 (N_12708,N_9294,N_6372);
and U12709 (N_12709,N_6630,N_7751);
nand U12710 (N_12710,N_8901,N_9096);
nor U12711 (N_12711,N_6432,N_5878);
nor U12712 (N_12712,N_7420,N_8491);
nor U12713 (N_12713,N_5732,N_7974);
nand U12714 (N_12714,N_7060,N_7303);
and U12715 (N_12715,N_7784,N_9659);
or U12716 (N_12716,N_9892,N_6319);
and U12717 (N_12717,N_9022,N_8365);
nor U12718 (N_12718,N_7306,N_5526);
nand U12719 (N_12719,N_6175,N_8601);
nor U12720 (N_12720,N_8246,N_8068);
nor U12721 (N_12721,N_9915,N_7481);
nand U12722 (N_12722,N_6345,N_9469);
nand U12723 (N_12723,N_6022,N_5842);
or U12724 (N_12724,N_8728,N_7756);
or U12725 (N_12725,N_8914,N_7885);
or U12726 (N_12726,N_5962,N_8984);
and U12727 (N_12727,N_7321,N_8500);
xnor U12728 (N_12728,N_9983,N_8150);
or U12729 (N_12729,N_7508,N_8799);
or U12730 (N_12730,N_7937,N_7832);
nand U12731 (N_12731,N_5216,N_6649);
and U12732 (N_12732,N_5161,N_9485);
or U12733 (N_12733,N_8764,N_9428);
and U12734 (N_12734,N_6080,N_7470);
and U12735 (N_12735,N_8503,N_8630);
or U12736 (N_12736,N_9958,N_7142);
nor U12737 (N_12737,N_9480,N_8484);
and U12738 (N_12738,N_5289,N_9775);
and U12739 (N_12739,N_8127,N_8423);
and U12740 (N_12740,N_6254,N_6968);
and U12741 (N_12741,N_6777,N_8363);
nand U12742 (N_12742,N_8421,N_7737);
and U12743 (N_12743,N_8312,N_5225);
nor U12744 (N_12744,N_5316,N_6117);
nand U12745 (N_12745,N_7961,N_6573);
and U12746 (N_12746,N_6049,N_8949);
nor U12747 (N_12747,N_9109,N_6794);
and U12748 (N_12748,N_5609,N_5831);
nor U12749 (N_12749,N_6614,N_9295);
and U12750 (N_12750,N_6865,N_6582);
or U12751 (N_12751,N_7918,N_8868);
and U12752 (N_12752,N_5849,N_5885);
xor U12753 (N_12753,N_9086,N_7161);
nand U12754 (N_12754,N_7145,N_9107);
and U12755 (N_12755,N_8726,N_8405);
and U12756 (N_12756,N_8441,N_7929);
and U12757 (N_12757,N_7905,N_8875);
nor U12758 (N_12758,N_9625,N_7359);
nor U12759 (N_12759,N_6089,N_8445);
nand U12760 (N_12760,N_7427,N_5326);
or U12761 (N_12761,N_9445,N_7025);
nor U12762 (N_12762,N_6648,N_8815);
nor U12763 (N_12763,N_9266,N_5058);
xnor U12764 (N_12764,N_5867,N_8466);
xnor U12765 (N_12765,N_6083,N_9440);
or U12766 (N_12766,N_5230,N_7965);
and U12767 (N_12767,N_7862,N_5223);
or U12768 (N_12768,N_9139,N_8353);
nand U12769 (N_12769,N_6305,N_9086);
nand U12770 (N_12770,N_8833,N_5870);
or U12771 (N_12771,N_9720,N_6055);
nor U12772 (N_12772,N_9391,N_9933);
and U12773 (N_12773,N_9646,N_5458);
or U12774 (N_12774,N_8069,N_8392);
xnor U12775 (N_12775,N_7138,N_6675);
and U12776 (N_12776,N_5797,N_8937);
and U12777 (N_12777,N_9998,N_5312);
nor U12778 (N_12778,N_5133,N_8552);
or U12779 (N_12779,N_5488,N_7469);
or U12780 (N_12780,N_8453,N_5581);
xor U12781 (N_12781,N_6942,N_7675);
or U12782 (N_12782,N_7330,N_5709);
nor U12783 (N_12783,N_5453,N_6982);
or U12784 (N_12784,N_6062,N_9850);
and U12785 (N_12785,N_5090,N_7388);
or U12786 (N_12786,N_7406,N_9943);
nor U12787 (N_12787,N_6737,N_7562);
and U12788 (N_12788,N_6552,N_7113);
xor U12789 (N_12789,N_9618,N_5895);
and U12790 (N_12790,N_9792,N_8695);
or U12791 (N_12791,N_5973,N_7036);
nor U12792 (N_12792,N_6218,N_8805);
nor U12793 (N_12793,N_6989,N_6962);
nor U12794 (N_12794,N_5276,N_5357);
nor U12795 (N_12795,N_8225,N_7872);
or U12796 (N_12796,N_7964,N_9404);
nor U12797 (N_12797,N_9998,N_9668);
xor U12798 (N_12798,N_5961,N_8402);
and U12799 (N_12799,N_7197,N_5996);
nor U12800 (N_12800,N_7285,N_8087);
or U12801 (N_12801,N_5860,N_9206);
and U12802 (N_12802,N_9852,N_5222);
xor U12803 (N_12803,N_8057,N_5908);
nor U12804 (N_12804,N_7897,N_5395);
and U12805 (N_12805,N_6835,N_9710);
xnor U12806 (N_12806,N_8937,N_5149);
nand U12807 (N_12807,N_5268,N_6162);
or U12808 (N_12808,N_6139,N_7827);
xnor U12809 (N_12809,N_9840,N_5278);
nor U12810 (N_12810,N_6535,N_8899);
nor U12811 (N_12811,N_7953,N_5919);
and U12812 (N_12812,N_9770,N_7175);
nand U12813 (N_12813,N_6774,N_9865);
and U12814 (N_12814,N_6173,N_8296);
nand U12815 (N_12815,N_5839,N_8257);
and U12816 (N_12816,N_6303,N_8904);
nor U12817 (N_12817,N_5615,N_7493);
or U12818 (N_12818,N_7916,N_5761);
or U12819 (N_12819,N_7287,N_7714);
xor U12820 (N_12820,N_9623,N_6217);
nand U12821 (N_12821,N_9589,N_6926);
nor U12822 (N_12822,N_7892,N_6390);
or U12823 (N_12823,N_5433,N_8534);
nand U12824 (N_12824,N_5907,N_6153);
or U12825 (N_12825,N_9254,N_7098);
nand U12826 (N_12826,N_5321,N_5951);
nand U12827 (N_12827,N_8247,N_6107);
xnor U12828 (N_12828,N_9060,N_7127);
and U12829 (N_12829,N_9178,N_7720);
and U12830 (N_12830,N_7030,N_5761);
nor U12831 (N_12831,N_7698,N_7658);
or U12832 (N_12832,N_6603,N_6797);
xor U12833 (N_12833,N_8528,N_7083);
nor U12834 (N_12834,N_6042,N_9828);
nor U12835 (N_12835,N_9646,N_9566);
and U12836 (N_12836,N_5162,N_8874);
nor U12837 (N_12837,N_9789,N_8105);
or U12838 (N_12838,N_8736,N_9890);
or U12839 (N_12839,N_7873,N_9129);
nor U12840 (N_12840,N_7298,N_7088);
nor U12841 (N_12841,N_6452,N_7883);
or U12842 (N_12842,N_9564,N_8263);
nor U12843 (N_12843,N_7431,N_6004);
or U12844 (N_12844,N_5514,N_8563);
and U12845 (N_12845,N_5789,N_9920);
nor U12846 (N_12846,N_6259,N_9865);
or U12847 (N_12847,N_5605,N_7750);
or U12848 (N_12848,N_9805,N_9846);
nor U12849 (N_12849,N_6800,N_6842);
nand U12850 (N_12850,N_6301,N_8828);
xnor U12851 (N_12851,N_6508,N_8731);
or U12852 (N_12852,N_9785,N_6368);
nand U12853 (N_12853,N_8990,N_5458);
and U12854 (N_12854,N_7187,N_6379);
or U12855 (N_12855,N_7522,N_7417);
or U12856 (N_12856,N_9119,N_6802);
nand U12857 (N_12857,N_7219,N_8876);
and U12858 (N_12858,N_6691,N_7143);
nor U12859 (N_12859,N_6584,N_5384);
and U12860 (N_12860,N_6856,N_6308);
or U12861 (N_12861,N_7225,N_8605);
nand U12862 (N_12862,N_6823,N_8574);
nor U12863 (N_12863,N_8007,N_6506);
and U12864 (N_12864,N_7744,N_8579);
xnor U12865 (N_12865,N_7498,N_5617);
nor U12866 (N_12866,N_9349,N_8467);
nor U12867 (N_12867,N_5256,N_8621);
nand U12868 (N_12868,N_9005,N_7545);
nor U12869 (N_12869,N_8013,N_8266);
nand U12870 (N_12870,N_5085,N_9158);
nor U12871 (N_12871,N_6292,N_8327);
nor U12872 (N_12872,N_7859,N_7832);
or U12873 (N_12873,N_8249,N_5082);
nand U12874 (N_12874,N_7389,N_5221);
and U12875 (N_12875,N_9253,N_8016);
nor U12876 (N_12876,N_8749,N_6459);
nand U12877 (N_12877,N_6804,N_6389);
xor U12878 (N_12878,N_8693,N_9524);
nand U12879 (N_12879,N_7177,N_6591);
or U12880 (N_12880,N_5887,N_9434);
and U12881 (N_12881,N_8986,N_9171);
and U12882 (N_12882,N_9461,N_7476);
nor U12883 (N_12883,N_5810,N_7774);
or U12884 (N_12884,N_8661,N_5091);
nand U12885 (N_12885,N_7377,N_8164);
xor U12886 (N_12886,N_6410,N_5919);
or U12887 (N_12887,N_7339,N_6333);
nor U12888 (N_12888,N_7882,N_7154);
and U12889 (N_12889,N_5576,N_5746);
nand U12890 (N_12890,N_6603,N_7651);
or U12891 (N_12891,N_6326,N_5460);
or U12892 (N_12892,N_9059,N_5324);
or U12893 (N_12893,N_9042,N_5618);
nand U12894 (N_12894,N_9197,N_7094);
nor U12895 (N_12895,N_5725,N_7822);
nor U12896 (N_12896,N_7260,N_8497);
or U12897 (N_12897,N_7495,N_7951);
and U12898 (N_12898,N_5305,N_9241);
and U12899 (N_12899,N_5238,N_5738);
nor U12900 (N_12900,N_8665,N_5899);
or U12901 (N_12901,N_7975,N_9077);
nor U12902 (N_12902,N_6720,N_8742);
nor U12903 (N_12903,N_6573,N_8031);
nor U12904 (N_12904,N_7825,N_7404);
or U12905 (N_12905,N_8850,N_5210);
and U12906 (N_12906,N_8360,N_5255);
nor U12907 (N_12907,N_5909,N_5660);
and U12908 (N_12908,N_5846,N_7727);
or U12909 (N_12909,N_6821,N_9681);
or U12910 (N_12910,N_8610,N_5880);
or U12911 (N_12911,N_6553,N_5314);
and U12912 (N_12912,N_7842,N_8689);
or U12913 (N_12913,N_6962,N_8802);
and U12914 (N_12914,N_7968,N_6447);
nand U12915 (N_12915,N_5915,N_7747);
nor U12916 (N_12916,N_8010,N_5245);
xnor U12917 (N_12917,N_5668,N_9874);
nor U12918 (N_12918,N_8609,N_8502);
xor U12919 (N_12919,N_7086,N_8077);
nor U12920 (N_12920,N_9021,N_7215);
nor U12921 (N_12921,N_8182,N_6175);
and U12922 (N_12922,N_9078,N_6211);
or U12923 (N_12923,N_6142,N_5423);
xnor U12924 (N_12924,N_6661,N_8966);
or U12925 (N_12925,N_6563,N_8000);
xnor U12926 (N_12926,N_6033,N_7092);
and U12927 (N_12927,N_8214,N_7202);
or U12928 (N_12928,N_9833,N_9461);
nand U12929 (N_12929,N_5404,N_7819);
and U12930 (N_12930,N_9860,N_7517);
and U12931 (N_12931,N_6195,N_8539);
and U12932 (N_12932,N_7985,N_9442);
or U12933 (N_12933,N_5018,N_6810);
nand U12934 (N_12934,N_6440,N_7162);
nor U12935 (N_12935,N_9457,N_8369);
nand U12936 (N_12936,N_7855,N_8947);
nor U12937 (N_12937,N_5723,N_6200);
or U12938 (N_12938,N_9027,N_5395);
xnor U12939 (N_12939,N_9238,N_9628);
nor U12940 (N_12940,N_9396,N_7934);
nand U12941 (N_12941,N_7922,N_8536);
and U12942 (N_12942,N_7914,N_9962);
or U12943 (N_12943,N_5589,N_6333);
xnor U12944 (N_12944,N_8550,N_6650);
and U12945 (N_12945,N_7719,N_5856);
xor U12946 (N_12946,N_5739,N_6403);
nor U12947 (N_12947,N_9497,N_9378);
xnor U12948 (N_12948,N_9682,N_5677);
nand U12949 (N_12949,N_9919,N_9797);
xnor U12950 (N_12950,N_5093,N_5697);
and U12951 (N_12951,N_6241,N_9168);
and U12952 (N_12952,N_5397,N_5005);
xnor U12953 (N_12953,N_9444,N_6361);
nor U12954 (N_12954,N_6963,N_7686);
and U12955 (N_12955,N_9148,N_7761);
xnor U12956 (N_12956,N_5952,N_6614);
and U12957 (N_12957,N_9469,N_7854);
or U12958 (N_12958,N_7405,N_9601);
or U12959 (N_12959,N_5541,N_8624);
and U12960 (N_12960,N_9633,N_5930);
and U12961 (N_12961,N_9669,N_9302);
xnor U12962 (N_12962,N_8793,N_6412);
nand U12963 (N_12963,N_9727,N_5497);
or U12964 (N_12964,N_6219,N_7696);
or U12965 (N_12965,N_7424,N_7082);
nor U12966 (N_12966,N_9233,N_6723);
nand U12967 (N_12967,N_7399,N_6200);
or U12968 (N_12968,N_9823,N_6621);
and U12969 (N_12969,N_5132,N_8146);
nand U12970 (N_12970,N_5539,N_5474);
nor U12971 (N_12971,N_6233,N_7202);
and U12972 (N_12972,N_7334,N_9442);
nand U12973 (N_12973,N_5438,N_6370);
nand U12974 (N_12974,N_5565,N_7636);
or U12975 (N_12975,N_7964,N_8924);
nor U12976 (N_12976,N_7513,N_5067);
nor U12977 (N_12977,N_6882,N_7958);
nand U12978 (N_12978,N_5714,N_5966);
nand U12979 (N_12979,N_7610,N_9659);
nand U12980 (N_12980,N_8707,N_7391);
nand U12981 (N_12981,N_5568,N_8019);
or U12982 (N_12982,N_6533,N_7896);
or U12983 (N_12983,N_6477,N_9259);
or U12984 (N_12984,N_9162,N_8413);
and U12985 (N_12985,N_5841,N_5696);
and U12986 (N_12986,N_6871,N_6200);
or U12987 (N_12987,N_9477,N_9591);
nor U12988 (N_12988,N_7018,N_7056);
nand U12989 (N_12989,N_9433,N_5219);
nand U12990 (N_12990,N_8098,N_9843);
nor U12991 (N_12991,N_5263,N_9687);
nand U12992 (N_12992,N_7142,N_5901);
and U12993 (N_12993,N_6473,N_7085);
and U12994 (N_12994,N_5747,N_9647);
and U12995 (N_12995,N_5048,N_8676);
and U12996 (N_12996,N_6326,N_7629);
xor U12997 (N_12997,N_6486,N_7190);
or U12998 (N_12998,N_9539,N_5240);
nand U12999 (N_12999,N_9306,N_7249);
nand U13000 (N_13000,N_8494,N_6645);
or U13001 (N_13001,N_5528,N_5083);
and U13002 (N_13002,N_8952,N_9816);
and U13003 (N_13003,N_8939,N_5316);
and U13004 (N_13004,N_8702,N_5186);
nor U13005 (N_13005,N_8048,N_7171);
nand U13006 (N_13006,N_9662,N_7637);
nor U13007 (N_13007,N_8044,N_8640);
or U13008 (N_13008,N_8249,N_9881);
nor U13009 (N_13009,N_5210,N_9492);
nor U13010 (N_13010,N_6176,N_9466);
nand U13011 (N_13011,N_5721,N_8084);
and U13012 (N_13012,N_6722,N_6729);
nor U13013 (N_13013,N_5194,N_8581);
and U13014 (N_13014,N_7559,N_8287);
nand U13015 (N_13015,N_8885,N_6949);
nand U13016 (N_13016,N_7568,N_8105);
nor U13017 (N_13017,N_9325,N_6092);
or U13018 (N_13018,N_9911,N_8973);
and U13019 (N_13019,N_5756,N_5732);
and U13020 (N_13020,N_8082,N_7491);
nor U13021 (N_13021,N_5507,N_8371);
and U13022 (N_13022,N_7193,N_9015);
nor U13023 (N_13023,N_6387,N_9878);
and U13024 (N_13024,N_8163,N_9182);
and U13025 (N_13025,N_8805,N_5441);
nand U13026 (N_13026,N_7505,N_9159);
or U13027 (N_13027,N_7775,N_6030);
or U13028 (N_13028,N_5189,N_8975);
and U13029 (N_13029,N_5376,N_6424);
or U13030 (N_13030,N_9135,N_9311);
and U13031 (N_13031,N_7742,N_8565);
nand U13032 (N_13032,N_9869,N_6800);
or U13033 (N_13033,N_5872,N_9391);
or U13034 (N_13034,N_7047,N_7094);
and U13035 (N_13035,N_9349,N_9034);
nor U13036 (N_13036,N_7919,N_6911);
or U13037 (N_13037,N_9042,N_5906);
nand U13038 (N_13038,N_7949,N_6399);
nor U13039 (N_13039,N_5348,N_9615);
nand U13040 (N_13040,N_9817,N_9745);
nor U13041 (N_13041,N_7650,N_9745);
nor U13042 (N_13042,N_6536,N_6411);
nand U13043 (N_13043,N_8642,N_8080);
nand U13044 (N_13044,N_9580,N_7295);
and U13045 (N_13045,N_5048,N_8354);
nand U13046 (N_13046,N_7767,N_6609);
nor U13047 (N_13047,N_6755,N_8878);
xor U13048 (N_13048,N_8987,N_7753);
nor U13049 (N_13049,N_7435,N_6900);
or U13050 (N_13050,N_7114,N_7154);
and U13051 (N_13051,N_9033,N_7014);
and U13052 (N_13052,N_9710,N_7191);
nand U13053 (N_13053,N_7238,N_5732);
nand U13054 (N_13054,N_8808,N_6107);
nor U13055 (N_13055,N_9908,N_5818);
or U13056 (N_13056,N_8943,N_9670);
and U13057 (N_13057,N_8533,N_8215);
and U13058 (N_13058,N_9212,N_8555);
nor U13059 (N_13059,N_6869,N_9266);
nor U13060 (N_13060,N_8126,N_9018);
nand U13061 (N_13061,N_6802,N_6069);
nand U13062 (N_13062,N_6532,N_9030);
nor U13063 (N_13063,N_6757,N_5828);
and U13064 (N_13064,N_8363,N_9114);
nor U13065 (N_13065,N_6251,N_7174);
nor U13066 (N_13066,N_5282,N_9825);
or U13067 (N_13067,N_8766,N_8251);
nand U13068 (N_13068,N_8338,N_9792);
and U13069 (N_13069,N_7061,N_8815);
and U13070 (N_13070,N_8977,N_6333);
nor U13071 (N_13071,N_9658,N_7040);
or U13072 (N_13072,N_9645,N_7725);
nor U13073 (N_13073,N_8861,N_9424);
and U13074 (N_13074,N_9966,N_5863);
and U13075 (N_13075,N_5046,N_7079);
nor U13076 (N_13076,N_5350,N_9946);
or U13077 (N_13077,N_9970,N_9334);
nand U13078 (N_13078,N_8136,N_5231);
nor U13079 (N_13079,N_6707,N_7051);
or U13080 (N_13080,N_8852,N_8770);
nor U13081 (N_13081,N_8415,N_5891);
nand U13082 (N_13082,N_9866,N_8958);
and U13083 (N_13083,N_7731,N_7651);
xnor U13084 (N_13084,N_9498,N_7733);
or U13085 (N_13085,N_9286,N_6055);
xnor U13086 (N_13086,N_9271,N_8666);
nand U13087 (N_13087,N_7897,N_5473);
or U13088 (N_13088,N_7609,N_7003);
nor U13089 (N_13089,N_8330,N_6908);
and U13090 (N_13090,N_6008,N_7768);
or U13091 (N_13091,N_8612,N_9930);
nand U13092 (N_13092,N_5901,N_8808);
nand U13093 (N_13093,N_6070,N_8566);
nor U13094 (N_13094,N_5233,N_7425);
nand U13095 (N_13095,N_5498,N_8082);
nand U13096 (N_13096,N_8865,N_6751);
or U13097 (N_13097,N_5155,N_6044);
nand U13098 (N_13098,N_6815,N_9615);
nand U13099 (N_13099,N_8410,N_8798);
nand U13100 (N_13100,N_7742,N_9661);
or U13101 (N_13101,N_8963,N_7021);
and U13102 (N_13102,N_5668,N_8213);
and U13103 (N_13103,N_9483,N_7977);
nand U13104 (N_13104,N_5113,N_7456);
or U13105 (N_13105,N_7614,N_7354);
and U13106 (N_13106,N_8185,N_8565);
nand U13107 (N_13107,N_6698,N_7017);
and U13108 (N_13108,N_8100,N_7233);
nor U13109 (N_13109,N_6832,N_6324);
nand U13110 (N_13110,N_9636,N_9670);
nand U13111 (N_13111,N_7963,N_7342);
xor U13112 (N_13112,N_6806,N_5414);
or U13113 (N_13113,N_9119,N_7877);
nand U13114 (N_13114,N_9880,N_6012);
nor U13115 (N_13115,N_8030,N_6232);
xor U13116 (N_13116,N_9634,N_5349);
nor U13117 (N_13117,N_7244,N_6180);
xnor U13118 (N_13118,N_6085,N_5972);
nand U13119 (N_13119,N_6220,N_9651);
nor U13120 (N_13120,N_8363,N_8388);
and U13121 (N_13121,N_5008,N_6954);
nor U13122 (N_13122,N_5217,N_8691);
and U13123 (N_13123,N_8532,N_8049);
nand U13124 (N_13124,N_6381,N_7046);
or U13125 (N_13125,N_7833,N_5062);
or U13126 (N_13126,N_6665,N_6180);
nor U13127 (N_13127,N_6747,N_7759);
or U13128 (N_13128,N_5063,N_9053);
nand U13129 (N_13129,N_8591,N_7271);
nor U13130 (N_13130,N_8191,N_5618);
and U13131 (N_13131,N_6264,N_6938);
nor U13132 (N_13132,N_9682,N_9538);
and U13133 (N_13133,N_9598,N_6008);
and U13134 (N_13134,N_6221,N_5097);
xnor U13135 (N_13135,N_5118,N_7942);
and U13136 (N_13136,N_6317,N_5447);
nor U13137 (N_13137,N_8436,N_7679);
and U13138 (N_13138,N_8942,N_9601);
nor U13139 (N_13139,N_5568,N_6777);
and U13140 (N_13140,N_7522,N_8322);
nand U13141 (N_13141,N_7898,N_6941);
or U13142 (N_13142,N_8301,N_8712);
and U13143 (N_13143,N_7909,N_5919);
and U13144 (N_13144,N_8661,N_6701);
xor U13145 (N_13145,N_6879,N_8103);
nor U13146 (N_13146,N_9446,N_7140);
nand U13147 (N_13147,N_6466,N_7494);
nor U13148 (N_13148,N_5916,N_9643);
and U13149 (N_13149,N_8538,N_5221);
and U13150 (N_13150,N_6030,N_7270);
and U13151 (N_13151,N_6501,N_7075);
nor U13152 (N_13152,N_5171,N_6655);
or U13153 (N_13153,N_5943,N_5305);
or U13154 (N_13154,N_7261,N_6637);
and U13155 (N_13155,N_8364,N_5456);
or U13156 (N_13156,N_7837,N_6861);
and U13157 (N_13157,N_8692,N_8952);
or U13158 (N_13158,N_6113,N_8746);
or U13159 (N_13159,N_6111,N_7867);
and U13160 (N_13160,N_8781,N_9917);
and U13161 (N_13161,N_8269,N_8008);
and U13162 (N_13162,N_6651,N_9652);
or U13163 (N_13163,N_5696,N_5912);
nand U13164 (N_13164,N_9677,N_6637);
or U13165 (N_13165,N_5635,N_9781);
and U13166 (N_13166,N_5249,N_9713);
or U13167 (N_13167,N_9431,N_9698);
or U13168 (N_13168,N_8501,N_9704);
nor U13169 (N_13169,N_5729,N_5798);
xor U13170 (N_13170,N_8713,N_8142);
or U13171 (N_13171,N_9164,N_5653);
nor U13172 (N_13172,N_5737,N_7747);
nor U13173 (N_13173,N_8326,N_9056);
nand U13174 (N_13174,N_6060,N_8182);
xnor U13175 (N_13175,N_9012,N_8288);
and U13176 (N_13176,N_5649,N_8492);
nor U13177 (N_13177,N_8764,N_7096);
nor U13178 (N_13178,N_9161,N_7095);
xnor U13179 (N_13179,N_9823,N_7558);
xor U13180 (N_13180,N_7586,N_7478);
or U13181 (N_13181,N_7709,N_6128);
nor U13182 (N_13182,N_9853,N_5403);
and U13183 (N_13183,N_6505,N_6644);
or U13184 (N_13184,N_7394,N_7401);
xnor U13185 (N_13185,N_5096,N_6831);
xnor U13186 (N_13186,N_9627,N_5685);
or U13187 (N_13187,N_8867,N_8998);
or U13188 (N_13188,N_5223,N_6660);
and U13189 (N_13189,N_6878,N_7703);
nor U13190 (N_13190,N_7902,N_8382);
xnor U13191 (N_13191,N_5635,N_9987);
nor U13192 (N_13192,N_6445,N_5396);
and U13193 (N_13193,N_6573,N_7130);
nor U13194 (N_13194,N_8783,N_8847);
nand U13195 (N_13195,N_9416,N_5710);
nor U13196 (N_13196,N_9505,N_9883);
or U13197 (N_13197,N_5411,N_8411);
and U13198 (N_13198,N_6792,N_7146);
nor U13199 (N_13199,N_5285,N_9209);
nor U13200 (N_13200,N_7282,N_7666);
nand U13201 (N_13201,N_9620,N_6363);
or U13202 (N_13202,N_8326,N_9328);
or U13203 (N_13203,N_9415,N_7782);
nor U13204 (N_13204,N_9509,N_9763);
and U13205 (N_13205,N_8712,N_7023);
nand U13206 (N_13206,N_6566,N_6271);
xor U13207 (N_13207,N_8214,N_6144);
nand U13208 (N_13208,N_8047,N_5451);
nand U13209 (N_13209,N_5027,N_9530);
and U13210 (N_13210,N_7858,N_5133);
nand U13211 (N_13211,N_5224,N_5004);
nor U13212 (N_13212,N_8948,N_9593);
nand U13213 (N_13213,N_9813,N_9188);
nor U13214 (N_13214,N_9923,N_5004);
or U13215 (N_13215,N_9662,N_7686);
nand U13216 (N_13216,N_7226,N_5314);
or U13217 (N_13217,N_9872,N_6404);
nor U13218 (N_13218,N_8564,N_6045);
xor U13219 (N_13219,N_6782,N_5088);
xor U13220 (N_13220,N_7612,N_9538);
and U13221 (N_13221,N_8083,N_7423);
xnor U13222 (N_13222,N_5763,N_7791);
nand U13223 (N_13223,N_5988,N_5060);
nand U13224 (N_13224,N_7087,N_7479);
nor U13225 (N_13225,N_7153,N_7711);
nand U13226 (N_13226,N_5169,N_8345);
xor U13227 (N_13227,N_9115,N_6186);
nand U13228 (N_13228,N_8534,N_7447);
nand U13229 (N_13229,N_9671,N_5793);
or U13230 (N_13230,N_7967,N_5966);
nand U13231 (N_13231,N_6424,N_5668);
and U13232 (N_13232,N_8335,N_8010);
and U13233 (N_13233,N_8688,N_6778);
and U13234 (N_13234,N_7083,N_5326);
nor U13235 (N_13235,N_9994,N_7635);
xor U13236 (N_13236,N_9456,N_5743);
nand U13237 (N_13237,N_6836,N_8515);
xnor U13238 (N_13238,N_6589,N_9973);
nor U13239 (N_13239,N_9029,N_6163);
or U13240 (N_13240,N_9133,N_5929);
nor U13241 (N_13241,N_5081,N_6611);
xor U13242 (N_13242,N_7142,N_6706);
or U13243 (N_13243,N_6049,N_8808);
nand U13244 (N_13244,N_6294,N_5470);
or U13245 (N_13245,N_7921,N_5801);
nor U13246 (N_13246,N_5471,N_9559);
nand U13247 (N_13247,N_6596,N_7235);
xnor U13248 (N_13248,N_9087,N_5313);
nor U13249 (N_13249,N_6065,N_8992);
and U13250 (N_13250,N_6873,N_7159);
and U13251 (N_13251,N_8791,N_9120);
or U13252 (N_13252,N_9369,N_9841);
nand U13253 (N_13253,N_9990,N_8792);
and U13254 (N_13254,N_8110,N_9845);
nor U13255 (N_13255,N_6909,N_9456);
nor U13256 (N_13256,N_8662,N_7874);
or U13257 (N_13257,N_9098,N_5195);
nor U13258 (N_13258,N_9439,N_9052);
nand U13259 (N_13259,N_8826,N_8726);
or U13260 (N_13260,N_7882,N_5225);
nand U13261 (N_13261,N_5641,N_7588);
and U13262 (N_13262,N_8824,N_9505);
and U13263 (N_13263,N_6826,N_8437);
or U13264 (N_13264,N_5926,N_5764);
nor U13265 (N_13265,N_6053,N_9460);
or U13266 (N_13266,N_8391,N_9307);
and U13267 (N_13267,N_7776,N_6450);
or U13268 (N_13268,N_6795,N_6674);
or U13269 (N_13269,N_9158,N_9299);
or U13270 (N_13270,N_7911,N_5338);
nor U13271 (N_13271,N_8671,N_9987);
and U13272 (N_13272,N_8861,N_9065);
xnor U13273 (N_13273,N_5348,N_7430);
nor U13274 (N_13274,N_5958,N_8035);
or U13275 (N_13275,N_7685,N_5288);
xor U13276 (N_13276,N_5929,N_5077);
nor U13277 (N_13277,N_6734,N_8184);
xor U13278 (N_13278,N_5057,N_5649);
nand U13279 (N_13279,N_5734,N_8469);
nand U13280 (N_13280,N_7848,N_6696);
nand U13281 (N_13281,N_5851,N_7320);
nor U13282 (N_13282,N_7226,N_9489);
or U13283 (N_13283,N_7281,N_6409);
and U13284 (N_13284,N_7328,N_7414);
nor U13285 (N_13285,N_5995,N_8513);
nor U13286 (N_13286,N_5431,N_9110);
xor U13287 (N_13287,N_7017,N_8665);
and U13288 (N_13288,N_5360,N_9343);
xor U13289 (N_13289,N_8397,N_7615);
or U13290 (N_13290,N_9529,N_5789);
and U13291 (N_13291,N_9486,N_8264);
or U13292 (N_13292,N_8303,N_8746);
or U13293 (N_13293,N_8381,N_7536);
xnor U13294 (N_13294,N_5183,N_5240);
nand U13295 (N_13295,N_6511,N_5971);
or U13296 (N_13296,N_6223,N_7529);
nor U13297 (N_13297,N_9584,N_5499);
and U13298 (N_13298,N_7115,N_5746);
nand U13299 (N_13299,N_8172,N_7138);
nor U13300 (N_13300,N_8521,N_5387);
xor U13301 (N_13301,N_8565,N_9269);
nand U13302 (N_13302,N_7905,N_7290);
and U13303 (N_13303,N_5656,N_6843);
nand U13304 (N_13304,N_9693,N_8462);
nand U13305 (N_13305,N_8568,N_6272);
nand U13306 (N_13306,N_8202,N_8367);
nor U13307 (N_13307,N_8606,N_6639);
nand U13308 (N_13308,N_6933,N_9002);
nand U13309 (N_13309,N_6751,N_8634);
xor U13310 (N_13310,N_6809,N_9649);
nand U13311 (N_13311,N_7184,N_6777);
nor U13312 (N_13312,N_9174,N_9160);
and U13313 (N_13313,N_8067,N_8428);
nor U13314 (N_13314,N_6793,N_7982);
or U13315 (N_13315,N_7116,N_8635);
nand U13316 (N_13316,N_5341,N_6613);
nor U13317 (N_13317,N_6920,N_9376);
nor U13318 (N_13318,N_9153,N_8100);
or U13319 (N_13319,N_9295,N_7006);
nor U13320 (N_13320,N_5149,N_9881);
or U13321 (N_13321,N_5175,N_6864);
and U13322 (N_13322,N_8297,N_5898);
and U13323 (N_13323,N_9595,N_6218);
and U13324 (N_13324,N_9832,N_5841);
nand U13325 (N_13325,N_7978,N_5079);
xor U13326 (N_13326,N_5778,N_6804);
nand U13327 (N_13327,N_8450,N_5777);
nor U13328 (N_13328,N_8857,N_5967);
nand U13329 (N_13329,N_9781,N_9216);
or U13330 (N_13330,N_9820,N_9263);
nand U13331 (N_13331,N_5215,N_5465);
and U13332 (N_13332,N_9215,N_7750);
xor U13333 (N_13333,N_9491,N_6861);
or U13334 (N_13334,N_8740,N_8069);
nor U13335 (N_13335,N_7819,N_7217);
xor U13336 (N_13336,N_7897,N_5516);
or U13337 (N_13337,N_7337,N_9838);
and U13338 (N_13338,N_9495,N_6550);
or U13339 (N_13339,N_6450,N_9189);
or U13340 (N_13340,N_7547,N_6128);
nor U13341 (N_13341,N_8860,N_6403);
or U13342 (N_13342,N_8417,N_9791);
xor U13343 (N_13343,N_7189,N_6326);
and U13344 (N_13344,N_8594,N_7570);
nor U13345 (N_13345,N_6006,N_8772);
or U13346 (N_13346,N_7780,N_5880);
or U13347 (N_13347,N_8682,N_8721);
nor U13348 (N_13348,N_7050,N_8787);
xnor U13349 (N_13349,N_9569,N_7374);
nor U13350 (N_13350,N_8382,N_8571);
and U13351 (N_13351,N_6753,N_7717);
nor U13352 (N_13352,N_8713,N_6112);
nor U13353 (N_13353,N_6298,N_8700);
or U13354 (N_13354,N_7952,N_6999);
nor U13355 (N_13355,N_6320,N_8840);
or U13356 (N_13356,N_8519,N_8416);
nor U13357 (N_13357,N_7786,N_9598);
or U13358 (N_13358,N_9178,N_5751);
and U13359 (N_13359,N_7323,N_7708);
nor U13360 (N_13360,N_6029,N_5945);
or U13361 (N_13361,N_8016,N_7868);
or U13362 (N_13362,N_6970,N_9868);
or U13363 (N_13363,N_9610,N_7099);
xnor U13364 (N_13364,N_5951,N_5161);
and U13365 (N_13365,N_6563,N_7502);
or U13366 (N_13366,N_5763,N_8910);
or U13367 (N_13367,N_9576,N_5496);
and U13368 (N_13368,N_7853,N_8704);
and U13369 (N_13369,N_6322,N_9667);
nor U13370 (N_13370,N_8595,N_6195);
nand U13371 (N_13371,N_5754,N_9783);
xor U13372 (N_13372,N_5253,N_6985);
and U13373 (N_13373,N_5323,N_9831);
and U13374 (N_13374,N_9200,N_9321);
nand U13375 (N_13375,N_9355,N_5558);
and U13376 (N_13376,N_5493,N_6994);
or U13377 (N_13377,N_5094,N_9737);
and U13378 (N_13378,N_5145,N_8660);
and U13379 (N_13379,N_8042,N_9834);
or U13380 (N_13380,N_6060,N_6747);
xnor U13381 (N_13381,N_9826,N_9838);
nor U13382 (N_13382,N_8704,N_9588);
or U13383 (N_13383,N_6946,N_6520);
or U13384 (N_13384,N_8493,N_7579);
nand U13385 (N_13385,N_8357,N_7077);
or U13386 (N_13386,N_7236,N_6596);
and U13387 (N_13387,N_8472,N_7828);
or U13388 (N_13388,N_7120,N_7140);
nor U13389 (N_13389,N_9776,N_8626);
xor U13390 (N_13390,N_8477,N_9378);
or U13391 (N_13391,N_9080,N_9943);
nor U13392 (N_13392,N_8793,N_9952);
nand U13393 (N_13393,N_6595,N_7777);
nor U13394 (N_13394,N_6099,N_5543);
xnor U13395 (N_13395,N_7513,N_5028);
nor U13396 (N_13396,N_8717,N_6525);
or U13397 (N_13397,N_5908,N_6689);
nor U13398 (N_13398,N_6623,N_8614);
xor U13399 (N_13399,N_9158,N_5586);
nor U13400 (N_13400,N_5411,N_6198);
nor U13401 (N_13401,N_5787,N_7315);
and U13402 (N_13402,N_8952,N_9723);
nand U13403 (N_13403,N_5133,N_7459);
or U13404 (N_13404,N_8432,N_5885);
nor U13405 (N_13405,N_8045,N_5851);
and U13406 (N_13406,N_8818,N_6269);
or U13407 (N_13407,N_5734,N_9181);
or U13408 (N_13408,N_9502,N_6458);
or U13409 (N_13409,N_8337,N_6214);
nand U13410 (N_13410,N_8755,N_6412);
and U13411 (N_13411,N_9987,N_6286);
nor U13412 (N_13412,N_8489,N_6803);
or U13413 (N_13413,N_9854,N_5827);
and U13414 (N_13414,N_7265,N_7594);
or U13415 (N_13415,N_8213,N_9761);
nand U13416 (N_13416,N_7011,N_5467);
nor U13417 (N_13417,N_5509,N_5989);
xnor U13418 (N_13418,N_9275,N_6168);
nor U13419 (N_13419,N_8134,N_6371);
nand U13420 (N_13420,N_9449,N_6470);
nand U13421 (N_13421,N_9673,N_5085);
nand U13422 (N_13422,N_8063,N_9234);
nor U13423 (N_13423,N_5397,N_9963);
nor U13424 (N_13424,N_9932,N_9636);
nor U13425 (N_13425,N_7077,N_9362);
xnor U13426 (N_13426,N_7993,N_8085);
or U13427 (N_13427,N_5711,N_5530);
and U13428 (N_13428,N_6755,N_9412);
nor U13429 (N_13429,N_5604,N_5779);
nor U13430 (N_13430,N_9446,N_7416);
or U13431 (N_13431,N_6948,N_7560);
and U13432 (N_13432,N_8136,N_9174);
and U13433 (N_13433,N_7325,N_5971);
nor U13434 (N_13434,N_6582,N_9262);
nor U13435 (N_13435,N_8130,N_6376);
and U13436 (N_13436,N_9426,N_8129);
or U13437 (N_13437,N_5143,N_5932);
or U13438 (N_13438,N_9218,N_9054);
nand U13439 (N_13439,N_5566,N_6627);
and U13440 (N_13440,N_7867,N_8406);
nor U13441 (N_13441,N_6283,N_6844);
or U13442 (N_13442,N_6309,N_6401);
nand U13443 (N_13443,N_7341,N_6166);
and U13444 (N_13444,N_7379,N_6296);
nand U13445 (N_13445,N_9390,N_6246);
nand U13446 (N_13446,N_7379,N_8388);
xor U13447 (N_13447,N_5958,N_6893);
or U13448 (N_13448,N_5460,N_5355);
nor U13449 (N_13449,N_8506,N_5556);
or U13450 (N_13450,N_9119,N_7933);
xor U13451 (N_13451,N_7671,N_6437);
or U13452 (N_13452,N_6241,N_7773);
and U13453 (N_13453,N_7502,N_7167);
nor U13454 (N_13454,N_7566,N_6697);
nand U13455 (N_13455,N_9006,N_9927);
nand U13456 (N_13456,N_6029,N_6541);
nand U13457 (N_13457,N_9357,N_6759);
nor U13458 (N_13458,N_9146,N_7188);
and U13459 (N_13459,N_6576,N_7819);
nor U13460 (N_13460,N_9018,N_7364);
or U13461 (N_13461,N_6981,N_5205);
nand U13462 (N_13462,N_6866,N_7854);
xor U13463 (N_13463,N_6427,N_6315);
and U13464 (N_13464,N_6313,N_5154);
and U13465 (N_13465,N_8207,N_5928);
and U13466 (N_13466,N_9687,N_7688);
or U13467 (N_13467,N_9545,N_6119);
nand U13468 (N_13468,N_8076,N_6071);
nand U13469 (N_13469,N_8162,N_6470);
and U13470 (N_13470,N_9510,N_7581);
xnor U13471 (N_13471,N_6717,N_6929);
and U13472 (N_13472,N_7861,N_5519);
xor U13473 (N_13473,N_9663,N_9427);
nor U13474 (N_13474,N_9781,N_5789);
nor U13475 (N_13475,N_7644,N_6628);
xor U13476 (N_13476,N_9390,N_7618);
xor U13477 (N_13477,N_8507,N_7351);
or U13478 (N_13478,N_6539,N_5033);
nor U13479 (N_13479,N_6392,N_7817);
nor U13480 (N_13480,N_5554,N_9785);
and U13481 (N_13481,N_6823,N_8605);
nor U13482 (N_13482,N_9552,N_8714);
or U13483 (N_13483,N_6192,N_7055);
and U13484 (N_13484,N_7521,N_9960);
nor U13485 (N_13485,N_7808,N_8962);
xnor U13486 (N_13486,N_9685,N_8080);
and U13487 (N_13487,N_7438,N_7321);
nor U13488 (N_13488,N_9621,N_9973);
nor U13489 (N_13489,N_9526,N_7582);
and U13490 (N_13490,N_7507,N_6558);
xnor U13491 (N_13491,N_8506,N_6657);
nand U13492 (N_13492,N_6601,N_9106);
and U13493 (N_13493,N_8930,N_8121);
nand U13494 (N_13494,N_8995,N_6184);
nor U13495 (N_13495,N_6543,N_5342);
nand U13496 (N_13496,N_5685,N_9286);
nor U13497 (N_13497,N_7401,N_7762);
nor U13498 (N_13498,N_9341,N_6104);
nand U13499 (N_13499,N_9007,N_6248);
nor U13500 (N_13500,N_5445,N_9046);
or U13501 (N_13501,N_5121,N_6234);
and U13502 (N_13502,N_5646,N_5628);
or U13503 (N_13503,N_7603,N_6025);
nand U13504 (N_13504,N_7294,N_8137);
xnor U13505 (N_13505,N_9783,N_6472);
or U13506 (N_13506,N_9187,N_5141);
and U13507 (N_13507,N_7943,N_7773);
xnor U13508 (N_13508,N_8761,N_6108);
nand U13509 (N_13509,N_7423,N_7972);
nand U13510 (N_13510,N_8544,N_5984);
or U13511 (N_13511,N_5899,N_9423);
and U13512 (N_13512,N_6374,N_8442);
and U13513 (N_13513,N_7501,N_9653);
nand U13514 (N_13514,N_9226,N_9944);
nand U13515 (N_13515,N_8547,N_6396);
nor U13516 (N_13516,N_6855,N_9286);
and U13517 (N_13517,N_9247,N_6492);
or U13518 (N_13518,N_8730,N_7882);
or U13519 (N_13519,N_8008,N_7629);
nor U13520 (N_13520,N_9989,N_6029);
and U13521 (N_13521,N_7595,N_7249);
or U13522 (N_13522,N_9267,N_8438);
or U13523 (N_13523,N_8588,N_7830);
and U13524 (N_13524,N_7692,N_8297);
or U13525 (N_13525,N_6452,N_8468);
nor U13526 (N_13526,N_9938,N_5386);
nor U13527 (N_13527,N_9595,N_9912);
or U13528 (N_13528,N_5262,N_7747);
or U13529 (N_13529,N_5812,N_7256);
nand U13530 (N_13530,N_5817,N_9892);
or U13531 (N_13531,N_5137,N_8380);
nor U13532 (N_13532,N_7479,N_8037);
or U13533 (N_13533,N_7866,N_8987);
nand U13534 (N_13534,N_9735,N_7077);
nand U13535 (N_13535,N_9662,N_6325);
nor U13536 (N_13536,N_6582,N_6867);
nor U13537 (N_13537,N_5707,N_5009);
nand U13538 (N_13538,N_5574,N_5169);
nor U13539 (N_13539,N_5397,N_5660);
nand U13540 (N_13540,N_6485,N_6849);
nand U13541 (N_13541,N_8398,N_8132);
or U13542 (N_13542,N_8325,N_9902);
nor U13543 (N_13543,N_6213,N_7191);
and U13544 (N_13544,N_9312,N_5075);
and U13545 (N_13545,N_9968,N_5759);
xor U13546 (N_13546,N_5718,N_8689);
and U13547 (N_13547,N_5819,N_7575);
or U13548 (N_13548,N_5191,N_5351);
and U13549 (N_13549,N_7713,N_6799);
nor U13550 (N_13550,N_7585,N_8946);
nand U13551 (N_13551,N_6594,N_6974);
nand U13552 (N_13552,N_8376,N_6854);
nor U13553 (N_13553,N_8593,N_5699);
xor U13554 (N_13554,N_5343,N_8445);
and U13555 (N_13555,N_7888,N_7420);
or U13556 (N_13556,N_8415,N_6652);
nand U13557 (N_13557,N_8630,N_6922);
or U13558 (N_13558,N_9694,N_6571);
or U13559 (N_13559,N_7570,N_9616);
nand U13560 (N_13560,N_9610,N_6820);
nor U13561 (N_13561,N_9344,N_9517);
or U13562 (N_13562,N_5366,N_8765);
xor U13563 (N_13563,N_6063,N_6369);
nand U13564 (N_13564,N_6635,N_7787);
and U13565 (N_13565,N_5625,N_6902);
or U13566 (N_13566,N_9538,N_6135);
and U13567 (N_13567,N_5772,N_9041);
or U13568 (N_13568,N_8654,N_5607);
nand U13569 (N_13569,N_6460,N_5454);
nand U13570 (N_13570,N_5226,N_6537);
and U13571 (N_13571,N_6268,N_7473);
and U13572 (N_13572,N_9077,N_7123);
and U13573 (N_13573,N_5484,N_6879);
nand U13574 (N_13574,N_6975,N_7330);
or U13575 (N_13575,N_9490,N_9561);
nor U13576 (N_13576,N_6710,N_5992);
xnor U13577 (N_13577,N_6052,N_5920);
or U13578 (N_13578,N_6488,N_6349);
or U13579 (N_13579,N_7056,N_9390);
nand U13580 (N_13580,N_9525,N_6430);
and U13581 (N_13581,N_8272,N_7735);
and U13582 (N_13582,N_8231,N_5959);
nor U13583 (N_13583,N_9299,N_9753);
and U13584 (N_13584,N_6532,N_8110);
nand U13585 (N_13585,N_5080,N_8225);
nor U13586 (N_13586,N_7271,N_8706);
nand U13587 (N_13587,N_9086,N_7271);
nand U13588 (N_13588,N_8892,N_5992);
xnor U13589 (N_13589,N_9086,N_6993);
and U13590 (N_13590,N_6351,N_8836);
xor U13591 (N_13591,N_9579,N_7277);
nor U13592 (N_13592,N_5658,N_5499);
and U13593 (N_13593,N_9782,N_6789);
or U13594 (N_13594,N_7316,N_9040);
xnor U13595 (N_13595,N_6815,N_8891);
nand U13596 (N_13596,N_9421,N_5424);
and U13597 (N_13597,N_9892,N_6910);
nand U13598 (N_13598,N_5928,N_9255);
nand U13599 (N_13599,N_5347,N_5273);
or U13600 (N_13600,N_8557,N_9878);
nand U13601 (N_13601,N_5689,N_6870);
and U13602 (N_13602,N_5797,N_7339);
nor U13603 (N_13603,N_6900,N_9958);
nor U13604 (N_13604,N_7075,N_5370);
xnor U13605 (N_13605,N_8769,N_8442);
or U13606 (N_13606,N_5392,N_9253);
and U13607 (N_13607,N_5996,N_5387);
nor U13608 (N_13608,N_8835,N_8353);
and U13609 (N_13609,N_8591,N_9512);
nor U13610 (N_13610,N_7680,N_5284);
nor U13611 (N_13611,N_9563,N_8629);
and U13612 (N_13612,N_5456,N_8088);
nand U13613 (N_13613,N_5401,N_9206);
and U13614 (N_13614,N_5075,N_9621);
or U13615 (N_13615,N_5350,N_8787);
xnor U13616 (N_13616,N_9619,N_9125);
nand U13617 (N_13617,N_7488,N_7792);
or U13618 (N_13618,N_5688,N_8820);
or U13619 (N_13619,N_5091,N_5462);
and U13620 (N_13620,N_6166,N_5053);
nand U13621 (N_13621,N_5419,N_8791);
nor U13622 (N_13622,N_7608,N_9263);
nand U13623 (N_13623,N_6057,N_9312);
nand U13624 (N_13624,N_5325,N_7436);
nand U13625 (N_13625,N_5551,N_7783);
or U13626 (N_13626,N_5525,N_8165);
nand U13627 (N_13627,N_7300,N_5591);
nand U13628 (N_13628,N_7802,N_8864);
nand U13629 (N_13629,N_7596,N_9780);
nand U13630 (N_13630,N_6805,N_8448);
nand U13631 (N_13631,N_7162,N_6999);
nor U13632 (N_13632,N_5788,N_9128);
nand U13633 (N_13633,N_5256,N_7747);
and U13634 (N_13634,N_6607,N_7603);
nor U13635 (N_13635,N_9735,N_5337);
nor U13636 (N_13636,N_5345,N_8670);
or U13637 (N_13637,N_8149,N_9366);
and U13638 (N_13638,N_8781,N_7232);
nand U13639 (N_13639,N_6242,N_9182);
nand U13640 (N_13640,N_7410,N_9063);
and U13641 (N_13641,N_5498,N_9992);
or U13642 (N_13642,N_8244,N_9209);
nand U13643 (N_13643,N_8041,N_8533);
nor U13644 (N_13644,N_5709,N_6248);
and U13645 (N_13645,N_9462,N_5109);
nor U13646 (N_13646,N_5596,N_5640);
xor U13647 (N_13647,N_6115,N_8918);
and U13648 (N_13648,N_8605,N_5400);
nor U13649 (N_13649,N_6549,N_8091);
xnor U13650 (N_13650,N_9940,N_9774);
and U13651 (N_13651,N_5166,N_7056);
nor U13652 (N_13652,N_5993,N_7163);
nand U13653 (N_13653,N_6250,N_7431);
xnor U13654 (N_13654,N_9818,N_9832);
xor U13655 (N_13655,N_8595,N_5519);
nand U13656 (N_13656,N_7625,N_5253);
and U13657 (N_13657,N_8721,N_7910);
nand U13658 (N_13658,N_7927,N_9564);
nand U13659 (N_13659,N_7241,N_6114);
nor U13660 (N_13660,N_9731,N_9211);
nand U13661 (N_13661,N_7806,N_5907);
and U13662 (N_13662,N_7567,N_5981);
nand U13663 (N_13663,N_8848,N_8423);
nor U13664 (N_13664,N_7064,N_5492);
nor U13665 (N_13665,N_7662,N_6998);
nand U13666 (N_13666,N_5339,N_8768);
nor U13667 (N_13667,N_6299,N_6796);
and U13668 (N_13668,N_6586,N_6720);
or U13669 (N_13669,N_8677,N_8826);
xnor U13670 (N_13670,N_5516,N_5455);
nand U13671 (N_13671,N_6542,N_5113);
and U13672 (N_13672,N_5321,N_5048);
nand U13673 (N_13673,N_6592,N_7595);
and U13674 (N_13674,N_6413,N_8823);
nand U13675 (N_13675,N_5290,N_8079);
nor U13676 (N_13676,N_9173,N_6180);
nand U13677 (N_13677,N_9183,N_6563);
or U13678 (N_13678,N_8752,N_7705);
nor U13679 (N_13679,N_5848,N_6857);
or U13680 (N_13680,N_5115,N_5013);
nand U13681 (N_13681,N_9348,N_5714);
and U13682 (N_13682,N_9464,N_6169);
nor U13683 (N_13683,N_7276,N_8056);
nand U13684 (N_13684,N_6715,N_7425);
and U13685 (N_13685,N_7741,N_8820);
or U13686 (N_13686,N_5462,N_5286);
or U13687 (N_13687,N_6224,N_9244);
nand U13688 (N_13688,N_7047,N_7603);
and U13689 (N_13689,N_9076,N_8507);
and U13690 (N_13690,N_9298,N_9266);
or U13691 (N_13691,N_7144,N_5004);
nand U13692 (N_13692,N_6632,N_5214);
nand U13693 (N_13693,N_5942,N_8496);
nand U13694 (N_13694,N_5311,N_6199);
or U13695 (N_13695,N_9300,N_6293);
xor U13696 (N_13696,N_7385,N_6085);
or U13697 (N_13697,N_9164,N_7533);
nand U13698 (N_13698,N_6149,N_9583);
nand U13699 (N_13699,N_8389,N_6322);
or U13700 (N_13700,N_9500,N_5470);
or U13701 (N_13701,N_7335,N_5664);
and U13702 (N_13702,N_5338,N_8820);
nand U13703 (N_13703,N_7496,N_8114);
nor U13704 (N_13704,N_9921,N_7982);
or U13705 (N_13705,N_5408,N_6476);
nand U13706 (N_13706,N_5435,N_6346);
or U13707 (N_13707,N_7566,N_6129);
xor U13708 (N_13708,N_6816,N_6591);
nand U13709 (N_13709,N_7890,N_6404);
xnor U13710 (N_13710,N_5198,N_5039);
nand U13711 (N_13711,N_7764,N_6081);
nand U13712 (N_13712,N_5549,N_5174);
xor U13713 (N_13713,N_8261,N_9741);
nand U13714 (N_13714,N_5691,N_7884);
and U13715 (N_13715,N_5642,N_9253);
and U13716 (N_13716,N_6667,N_9672);
nor U13717 (N_13717,N_9799,N_6909);
and U13718 (N_13718,N_9014,N_7568);
and U13719 (N_13719,N_6003,N_8802);
xnor U13720 (N_13720,N_9382,N_5869);
nor U13721 (N_13721,N_6042,N_7953);
and U13722 (N_13722,N_5136,N_7479);
nand U13723 (N_13723,N_6570,N_8501);
and U13724 (N_13724,N_7993,N_6191);
nor U13725 (N_13725,N_5920,N_8285);
nand U13726 (N_13726,N_9031,N_8811);
xor U13727 (N_13727,N_6779,N_5923);
or U13728 (N_13728,N_9630,N_8140);
or U13729 (N_13729,N_8101,N_7466);
nand U13730 (N_13730,N_8338,N_8489);
nand U13731 (N_13731,N_9416,N_9639);
nor U13732 (N_13732,N_9718,N_6754);
or U13733 (N_13733,N_9043,N_7310);
nand U13734 (N_13734,N_7018,N_7643);
nand U13735 (N_13735,N_6222,N_7331);
nor U13736 (N_13736,N_8932,N_9081);
or U13737 (N_13737,N_6413,N_7896);
nor U13738 (N_13738,N_7998,N_5956);
nor U13739 (N_13739,N_5164,N_8573);
and U13740 (N_13740,N_7366,N_6689);
or U13741 (N_13741,N_5192,N_6176);
and U13742 (N_13742,N_8442,N_5393);
nand U13743 (N_13743,N_8019,N_9376);
and U13744 (N_13744,N_7745,N_5803);
nor U13745 (N_13745,N_8519,N_6155);
or U13746 (N_13746,N_9218,N_7149);
xor U13747 (N_13747,N_8082,N_7575);
or U13748 (N_13748,N_7406,N_8168);
and U13749 (N_13749,N_9680,N_7952);
nand U13750 (N_13750,N_5754,N_7084);
nand U13751 (N_13751,N_6402,N_9401);
and U13752 (N_13752,N_7469,N_8803);
or U13753 (N_13753,N_7154,N_9959);
nor U13754 (N_13754,N_9676,N_7059);
nor U13755 (N_13755,N_5618,N_6772);
xnor U13756 (N_13756,N_9899,N_8677);
and U13757 (N_13757,N_5305,N_6305);
or U13758 (N_13758,N_5115,N_8577);
nor U13759 (N_13759,N_5737,N_9585);
and U13760 (N_13760,N_7901,N_5689);
nor U13761 (N_13761,N_7528,N_5427);
nor U13762 (N_13762,N_8905,N_9850);
and U13763 (N_13763,N_8609,N_8129);
xor U13764 (N_13764,N_8021,N_5705);
nor U13765 (N_13765,N_8322,N_8347);
and U13766 (N_13766,N_7262,N_5856);
nand U13767 (N_13767,N_5819,N_9558);
xor U13768 (N_13768,N_5763,N_5202);
nand U13769 (N_13769,N_5891,N_6524);
xnor U13770 (N_13770,N_9983,N_7431);
or U13771 (N_13771,N_7760,N_8499);
and U13772 (N_13772,N_8857,N_6500);
or U13773 (N_13773,N_5855,N_9776);
or U13774 (N_13774,N_8943,N_6774);
and U13775 (N_13775,N_8084,N_7638);
and U13776 (N_13776,N_5100,N_6446);
nand U13777 (N_13777,N_5283,N_5753);
or U13778 (N_13778,N_7394,N_7598);
or U13779 (N_13779,N_7125,N_8642);
or U13780 (N_13780,N_9768,N_5894);
nor U13781 (N_13781,N_6599,N_9982);
nor U13782 (N_13782,N_5268,N_8200);
nand U13783 (N_13783,N_7216,N_5817);
and U13784 (N_13784,N_8019,N_9823);
nand U13785 (N_13785,N_5227,N_6897);
nor U13786 (N_13786,N_8250,N_5371);
nand U13787 (N_13787,N_6259,N_5912);
or U13788 (N_13788,N_8747,N_5877);
xor U13789 (N_13789,N_9317,N_9355);
or U13790 (N_13790,N_7730,N_6781);
and U13791 (N_13791,N_5648,N_8747);
or U13792 (N_13792,N_6274,N_9187);
nand U13793 (N_13793,N_7451,N_8658);
nand U13794 (N_13794,N_8336,N_6288);
or U13795 (N_13795,N_5083,N_6698);
or U13796 (N_13796,N_6138,N_5004);
nor U13797 (N_13797,N_8862,N_9278);
or U13798 (N_13798,N_6944,N_9682);
or U13799 (N_13799,N_6168,N_6574);
and U13800 (N_13800,N_5914,N_5246);
xor U13801 (N_13801,N_6132,N_7658);
and U13802 (N_13802,N_7672,N_7401);
and U13803 (N_13803,N_6465,N_9979);
nand U13804 (N_13804,N_9091,N_8898);
or U13805 (N_13805,N_8672,N_5215);
xor U13806 (N_13806,N_5469,N_9646);
or U13807 (N_13807,N_5943,N_8617);
or U13808 (N_13808,N_8655,N_8432);
nor U13809 (N_13809,N_7687,N_5072);
or U13810 (N_13810,N_7709,N_5620);
nand U13811 (N_13811,N_6623,N_6599);
or U13812 (N_13812,N_7217,N_8323);
xnor U13813 (N_13813,N_7644,N_8718);
nor U13814 (N_13814,N_9663,N_5818);
nand U13815 (N_13815,N_5532,N_5614);
nand U13816 (N_13816,N_8502,N_9598);
or U13817 (N_13817,N_8247,N_6828);
nor U13818 (N_13818,N_6684,N_5301);
and U13819 (N_13819,N_6394,N_9019);
nand U13820 (N_13820,N_5317,N_5200);
nand U13821 (N_13821,N_5228,N_9603);
nand U13822 (N_13822,N_8083,N_6367);
or U13823 (N_13823,N_9534,N_8035);
or U13824 (N_13824,N_8243,N_5333);
or U13825 (N_13825,N_7749,N_5171);
or U13826 (N_13826,N_5146,N_9226);
nand U13827 (N_13827,N_9322,N_8393);
and U13828 (N_13828,N_5570,N_7496);
or U13829 (N_13829,N_9752,N_7198);
nor U13830 (N_13830,N_6917,N_9651);
nor U13831 (N_13831,N_8111,N_9690);
nand U13832 (N_13832,N_8881,N_6410);
or U13833 (N_13833,N_5109,N_8645);
nor U13834 (N_13834,N_8402,N_7889);
or U13835 (N_13835,N_8141,N_6043);
nor U13836 (N_13836,N_8307,N_5034);
nand U13837 (N_13837,N_8768,N_6424);
or U13838 (N_13838,N_7101,N_5628);
or U13839 (N_13839,N_8869,N_9147);
and U13840 (N_13840,N_7352,N_9025);
or U13841 (N_13841,N_7619,N_9602);
nor U13842 (N_13842,N_9903,N_8868);
nor U13843 (N_13843,N_7989,N_5832);
nand U13844 (N_13844,N_6967,N_7999);
nor U13845 (N_13845,N_8208,N_9197);
xor U13846 (N_13846,N_9146,N_7627);
and U13847 (N_13847,N_9557,N_8645);
or U13848 (N_13848,N_7990,N_8613);
nand U13849 (N_13849,N_6269,N_6864);
nor U13850 (N_13850,N_8138,N_6707);
nand U13851 (N_13851,N_9675,N_9250);
nor U13852 (N_13852,N_6407,N_9537);
and U13853 (N_13853,N_9494,N_5068);
nand U13854 (N_13854,N_9891,N_7046);
nand U13855 (N_13855,N_8905,N_9320);
nor U13856 (N_13856,N_7212,N_7636);
nand U13857 (N_13857,N_9089,N_6824);
xor U13858 (N_13858,N_5601,N_9788);
or U13859 (N_13859,N_9781,N_9881);
nand U13860 (N_13860,N_7304,N_9157);
or U13861 (N_13861,N_5872,N_5170);
xor U13862 (N_13862,N_6833,N_8662);
and U13863 (N_13863,N_9538,N_5889);
or U13864 (N_13864,N_8787,N_5207);
nor U13865 (N_13865,N_6687,N_6925);
xor U13866 (N_13866,N_5259,N_5467);
nand U13867 (N_13867,N_7303,N_9215);
nor U13868 (N_13868,N_5723,N_5709);
and U13869 (N_13869,N_5596,N_8158);
nand U13870 (N_13870,N_8487,N_8430);
nor U13871 (N_13871,N_9279,N_5720);
nand U13872 (N_13872,N_9448,N_8730);
or U13873 (N_13873,N_6481,N_6955);
or U13874 (N_13874,N_9045,N_7375);
or U13875 (N_13875,N_8841,N_8355);
or U13876 (N_13876,N_7266,N_6563);
or U13877 (N_13877,N_5645,N_7131);
or U13878 (N_13878,N_8044,N_9118);
or U13879 (N_13879,N_5186,N_6960);
and U13880 (N_13880,N_5065,N_7936);
or U13881 (N_13881,N_9389,N_9658);
and U13882 (N_13882,N_8125,N_9335);
xor U13883 (N_13883,N_5977,N_5524);
and U13884 (N_13884,N_8208,N_9855);
and U13885 (N_13885,N_7798,N_8555);
and U13886 (N_13886,N_5075,N_7699);
nor U13887 (N_13887,N_9160,N_8514);
xnor U13888 (N_13888,N_8411,N_9142);
or U13889 (N_13889,N_5778,N_8019);
nand U13890 (N_13890,N_8433,N_9486);
nor U13891 (N_13891,N_5898,N_7948);
xor U13892 (N_13892,N_7752,N_6479);
nand U13893 (N_13893,N_5875,N_7873);
nor U13894 (N_13894,N_8429,N_5192);
and U13895 (N_13895,N_8561,N_9625);
xor U13896 (N_13896,N_9816,N_5363);
or U13897 (N_13897,N_8790,N_6761);
and U13898 (N_13898,N_7706,N_5223);
xor U13899 (N_13899,N_5121,N_8115);
nand U13900 (N_13900,N_9071,N_9817);
or U13901 (N_13901,N_7557,N_5300);
or U13902 (N_13902,N_6295,N_5750);
or U13903 (N_13903,N_5737,N_5037);
nor U13904 (N_13904,N_5795,N_8171);
nand U13905 (N_13905,N_6147,N_9985);
nand U13906 (N_13906,N_5595,N_9735);
nor U13907 (N_13907,N_8352,N_9418);
nand U13908 (N_13908,N_5587,N_5850);
nand U13909 (N_13909,N_9397,N_8617);
or U13910 (N_13910,N_7986,N_9490);
nand U13911 (N_13911,N_6409,N_5759);
xnor U13912 (N_13912,N_9246,N_7647);
or U13913 (N_13913,N_9457,N_9310);
nor U13914 (N_13914,N_8064,N_8137);
xnor U13915 (N_13915,N_9998,N_7164);
nor U13916 (N_13916,N_5860,N_9031);
nor U13917 (N_13917,N_7596,N_6911);
nand U13918 (N_13918,N_6553,N_5620);
xnor U13919 (N_13919,N_6521,N_7356);
nand U13920 (N_13920,N_5602,N_5145);
nor U13921 (N_13921,N_8157,N_7749);
nand U13922 (N_13922,N_9282,N_6381);
and U13923 (N_13923,N_6060,N_9369);
or U13924 (N_13924,N_6261,N_5290);
or U13925 (N_13925,N_6386,N_6580);
or U13926 (N_13926,N_9754,N_7298);
or U13927 (N_13927,N_8512,N_6124);
or U13928 (N_13928,N_8242,N_8944);
nor U13929 (N_13929,N_8305,N_8586);
and U13930 (N_13930,N_7633,N_5659);
and U13931 (N_13931,N_9293,N_9275);
and U13932 (N_13932,N_6365,N_5347);
nand U13933 (N_13933,N_5938,N_6447);
and U13934 (N_13934,N_5972,N_6708);
nor U13935 (N_13935,N_8488,N_8976);
xor U13936 (N_13936,N_5961,N_8236);
and U13937 (N_13937,N_5094,N_5629);
nor U13938 (N_13938,N_7794,N_8518);
and U13939 (N_13939,N_9420,N_6144);
nand U13940 (N_13940,N_5649,N_8543);
nor U13941 (N_13941,N_5469,N_6749);
nand U13942 (N_13942,N_6928,N_6835);
or U13943 (N_13943,N_9863,N_7260);
nand U13944 (N_13944,N_7041,N_5421);
nor U13945 (N_13945,N_8290,N_6003);
or U13946 (N_13946,N_8445,N_9099);
and U13947 (N_13947,N_6428,N_5049);
and U13948 (N_13948,N_5030,N_7355);
and U13949 (N_13949,N_6456,N_6038);
xor U13950 (N_13950,N_5244,N_9412);
nand U13951 (N_13951,N_6551,N_5234);
or U13952 (N_13952,N_7784,N_8903);
or U13953 (N_13953,N_7130,N_8531);
nand U13954 (N_13954,N_6688,N_9575);
nand U13955 (N_13955,N_9778,N_9323);
or U13956 (N_13956,N_6527,N_7550);
nor U13957 (N_13957,N_6756,N_5024);
or U13958 (N_13958,N_5823,N_7473);
or U13959 (N_13959,N_5667,N_7999);
and U13960 (N_13960,N_9955,N_8277);
and U13961 (N_13961,N_5681,N_7583);
nand U13962 (N_13962,N_6187,N_5825);
or U13963 (N_13963,N_7454,N_7145);
nand U13964 (N_13964,N_7820,N_6531);
or U13965 (N_13965,N_5332,N_5330);
or U13966 (N_13966,N_6371,N_7364);
or U13967 (N_13967,N_9065,N_7176);
nand U13968 (N_13968,N_5432,N_8940);
nor U13969 (N_13969,N_6314,N_5987);
nand U13970 (N_13970,N_8467,N_9843);
or U13971 (N_13971,N_9810,N_6876);
xor U13972 (N_13972,N_5531,N_9755);
nor U13973 (N_13973,N_6702,N_6858);
xor U13974 (N_13974,N_5704,N_8246);
or U13975 (N_13975,N_7536,N_9012);
nor U13976 (N_13976,N_6150,N_8621);
and U13977 (N_13977,N_5944,N_7830);
xnor U13978 (N_13978,N_9411,N_6597);
nand U13979 (N_13979,N_8276,N_5761);
or U13980 (N_13980,N_6668,N_9602);
xor U13981 (N_13981,N_9141,N_9892);
nor U13982 (N_13982,N_6437,N_6560);
and U13983 (N_13983,N_6053,N_5271);
nor U13984 (N_13984,N_8229,N_5172);
nand U13985 (N_13985,N_5901,N_8894);
xor U13986 (N_13986,N_6880,N_7657);
and U13987 (N_13987,N_6004,N_5281);
nor U13988 (N_13988,N_8980,N_8605);
and U13989 (N_13989,N_9793,N_5776);
or U13990 (N_13990,N_8488,N_9002);
xnor U13991 (N_13991,N_5851,N_8438);
nand U13992 (N_13992,N_6433,N_5021);
nand U13993 (N_13993,N_8756,N_5052);
and U13994 (N_13994,N_5175,N_9586);
and U13995 (N_13995,N_9646,N_9392);
xor U13996 (N_13996,N_7656,N_7918);
and U13997 (N_13997,N_6447,N_7573);
and U13998 (N_13998,N_9684,N_5279);
nand U13999 (N_13999,N_8525,N_9073);
or U14000 (N_14000,N_7973,N_5247);
or U14001 (N_14001,N_7573,N_8101);
or U14002 (N_14002,N_6008,N_9071);
and U14003 (N_14003,N_7231,N_8726);
nand U14004 (N_14004,N_8830,N_9287);
and U14005 (N_14005,N_5371,N_7508);
or U14006 (N_14006,N_9434,N_9855);
and U14007 (N_14007,N_7243,N_5697);
or U14008 (N_14008,N_7380,N_6710);
nor U14009 (N_14009,N_7399,N_7625);
nor U14010 (N_14010,N_8387,N_8828);
nand U14011 (N_14011,N_8936,N_6048);
nand U14012 (N_14012,N_5953,N_7380);
or U14013 (N_14013,N_7558,N_9358);
nand U14014 (N_14014,N_7392,N_8315);
nor U14015 (N_14015,N_8028,N_8002);
nand U14016 (N_14016,N_9930,N_6403);
nand U14017 (N_14017,N_8147,N_5800);
nand U14018 (N_14018,N_6200,N_6636);
nor U14019 (N_14019,N_5570,N_7891);
nand U14020 (N_14020,N_9341,N_6945);
or U14021 (N_14021,N_6981,N_5471);
nand U14022 (N_14022,N_6661,N_5415);
and U14023 (N_14023,N_9737,N_5857);
nor U14024 (N_14024,N_6230,N_7126);
or U14025 (N_14025,N_8115,N_6597);
nor U14026 (N_14026,N_7270,N_8508);
nor U14027 (N_14027,N_9799,N_8303);
nand U14028 (N_14028,N_5225,N_8828);
nand U14029 (N_14029,N_8731,N_7765);
and U14030 (N_14030,N_5997,N_5814);
or U14031 (N_14031,N_9923,N_8267);
nor U14032 (N_14032,N_6853,N_5957);
xor U14033 (N_14033,N_6767,N_6375);
or U14034 (N_14034,N_5732,N_5928);
nor U14035 (N_14035,N_6803,N_7895);
nand U14036 (N_14036,N_8174,N_5569);
and U14037 (N_14037,N_7727,N_7885);
and U14038 (N_14038,N_6732,N_7217);
nand U14039 (N_14039,N_8134,N_6198);
or U14040 (N_14040,N_8754,N_6487);
nor U14041 (N_14041,N_5394,N_8124);
nand U14042 (N_14042,N_7166,N_9353);
nor U14043 (N_14043,N_7157,N_5802);
or U14044 (N_14044,N_7077,N_8316);
or U14045 (N_14045,N_9367,N_7328);
and U14046 (N_14046,N_6520,N_6841);
nand U14047 (N_14047,N_8928,N_8633);
and U14048 (N_14048,N_5419,N_5032);
nand U14049 (N_14049,N_8257,N_8606);
or U14050 (N_14050,N_6721,N_9671);
nand U14051 (N_14051,N_6222,N_7768);
xnor U14052 (N_14052,N_9684,N_5379);
xnor U14053 (N_14053,N_6381,N_5377);
xnor U14054 (N_14054,N_5843,N_8992);
nor U14055 (N_14055,N_7098,N_5729);
nor U14056 (N_14056,N_9779,N_6806);
nand U14057 (N_14057,N_9261,N_5321);
nor U14058 (N_14058,N_6609,N_7192);
nand U14059 (N_14059,N_8645,N_7928);
xor U14060 (N_14060,N_5939,N_6856);
nor U14061 (N_14061,N_7116,N_6480);
nand U14062 (N_14062,N_6620,N_8678);
nand U14063 (N_14063,N_5673,N_5686);
and U14064 (N_14064,N_7923,N_8308);
and U14065 (N_14065,N_6494,N_6020);
and U14066 (N_14066,N_9512,N_8615);
or U14067 (N_14067,N_6169,N_6497);
and U14068 (N_14068,N_8681,N_7269);
nand U14069 (N_14069,N_6623,N_6422);
or U14070 (N_14070,N_6909,N_6408);
and U14071 (N_14071,N_5266,N_7790);
and U14072 (N_14072,N_6619,N_6766);
or U14073 (N_14073,N_8944,N_5619);
nand U14074 (N_14074,N_8050,N_8043);
nor U14075 (N_14075,N_5523,N_9213);
and U14076 (N_14076,N_8162,N_8501);
and U14077 (N_14077,N_5773,N_7875);
nor U14078 (N_14078,N_5715,N_6245);
and U14079 (N_14079,N_5424,N_7353);
nor U14080 (N_14080,N_8408,N_5296);
nor U14081 (N_14081,N_6920,N_8058);
and U14082 (N_14082,N_6553,N_8615);
nand U14083 (N_14083,N_9043,N_6045);
and U14084 (N_14084,N_9988,N_7243);
nand U14085 (N_14085,N_7247,N_6725);
nand U14086 (N_14086,N_6920,N_6028);
nand U14087 (N_14087,N_5484,N_7341);
nand U14088 (N_14088,N_9040,N_8968);
nand U14089 (N_14089,N_6078,N_5807);
nand U14090 (N_14090,N_8399,N_7315);
xor U14091 (N_14091,N_9140,N_6022);
and U14092 (N_14092,N_8863,N_9277);
nor U14093 (N_14093,N_8489,N_8927);
xor U14094 (N_14094,N_8518,N_5713);
and U14095 (N_14095,N_8616,N_9165);
and U14096 (N_14096,N_5464,N_7848);
xor U14097 (N_14097,N_8605,N_9344);
or U14098 (N_14098,N_7625,N_7077);
and U14099 (N_14099,N_6285,N_6132);
nor U14100 (N_14100,N_7944,N_7629);
xnor U14101 (N_14101,N_6870,N_8485);
nand U14102 (N_14102,N_6990,N_8071);
nand U14103 (N_14103,N_9843,N_8937);
nand U14104 (N_14104,N_7088,N_5387);
nand U14105 (N_14105,N_5237,N_7546);
xnor U14106 (N_14106,N_6546,N_7776);
nand U14107 (N_14107,N_8851,N_5636);
and U14108 (N_14108,N_5597,N_7105);
nor U14109 (N_14109,N_9589,N_5897);
or U14110 (N_14110,N_5319,N_6164);
and U14111 (N_14111,N_5519,N_5436);
or U14112 (N_14112,N_6837,N_6649);
nor U14113 (N_14113,N_5660,N_8717);
nand U14114 (N_14114,N_9868,N_5330);
nor U14115 (N_14115,N_6987,N_8883);
nor U14116 (N_14116,N_8637,N_6923);
nand U14117 (N_14117,N_9346,N_6351);
nand U14118 (N_14118,N_7654,N_7831);
and U14119 (N_14119,N_9276,N_7587);
nor U14120 (N_14120,N_5867,N_9924);
and U14121 (N_14121,N_7097,N_5207);
or U14122 (N_14122,N_7810,N_9029);
and U14123 (N_14123,N_9768,N_9971);
xnor U14124 (N_14124,N_8151,N_5707);
nor U14125 (N_14125,N_7899,N_7512);
nand U14126 (N_14126,N_8625,N_8362);
nand U14127 (N_14127,N_8055,N_6194);
and U14128 (N_14128,N_5670,N_5951);
nor U14129 (N_14129,N_9371,N_9030);
and U14130 (N_14130,N_7516,N_6343);
nand U14131 (N_14131,N_6062,N_9388);
nor U14132 (N_14132,N_5831,N_5684);
nor U14133 (N_14133,N_5018,N_8839);
or U14134 (N_14134,N_9002,N_6562);
nand U14135 (N_14135,N_6053,N_6284);
or U14136 (N_14136,N_5614,N_6976);
xor U14137 (N_14137,N_5333,N_9845);
or U14138 (N_14138,N_6518,N_6143);
and U14139 (N_14139,N_6876,N_5022);
nor U14140 (N_14140,N_9219,N_5495);
and U14141 (N_14141,N_9615,N_8788);
xor U14142 (N_14142,N_6876,N_9911);
and U14143 (N_14143,N_6313,N_8925);
xor U14144 (N_14144,N_7934,N_8186);
or U14145 (N_14145,N_9622,N_6983);
nor U14146 (N_14146,N_6220,N_9194);
nand U14147 (N_14147,N_9390,N_8085);
nand U14148 (N_14148,N_7963,N_9535);
or U14149 (N_14149,N_6913,N_6881);
nand U14150 (N_14150,N_5942,N_6758);
nor U14151 (N_14151,N_5335,N_8099);
xnor U14152 (N_14152,N_6218,N_7786);
and U14153 (N_14153,N_6805,N_7127);
and U14154 (N_14154,N_8832,N_9311);
nand U14155 (N_14155,N_8861,N_7532);
or U14156 (N_14156,N_6462,N_9559);
nand U14157 (N_14157,N_7977,N_7746);
nor U14158 (N_14158,N_8576,N_7945);
and U14159 (N_14159,N_7827,N_6485);
and U14160 (N_14160,N_8959,N_8701);
or U14161 (N_14161,N_7794,N_9684);
nand U14162 (N_14162,N_6182,N_5062);
and U14163 (N_14163,N_5079,N_9495);
xor U14164 (N_14164,N_7028,N_9363);
and U14165 (N_14165,N_5653,N_5850);
xnor U14166 (N_14166,N_9082,N_5412);
nor U14167 (N_14167,N_5672,N_6833);
and U14168 (N_14168,N_8773,N_7668);
nor U14169 (N_14169,N_5142,N_6137);
nor U14170 (N_14170,N_5629,N_8502);
and U14171 (N_14171,N_9121,N_6221);
nand U14172 (N_14172,N_9831,N_8605);
and U14173 (N_14173,N_5587,N_8674);
and U14174 (N_14174,N_9216,N_7618);
or U14175 (N_14175,N_6112,N_6696);
nand U14176 (N_14176,N_5495,N_9737);
nor U14177 (N_14177,N_8482,N_8214);
nor U14178 (N_14178,N_6349,N_7646);
and U14179 (N_14179,N_8854,N_9827);
xor U14180 (N_14180,N_7166,N_5770);
or U14181 (N_14181,N_5016,N_6580);
and U14182 (N_14182,N_5588,N_9815);
and U14183 (N_14183,N_5562,N_6954);
nand U14184 (N_14184,N_9472,N_6676);
and U14185 (N_14185,N_9972,N_9686);
nand U14186 (N_14186,N_6645,N_6498);
nor U14187 (N_14187,N_5530,N_6602);
xor U14188 (N_14188,N_6857,N_8978);
and U14189 (N_14189,N_8306,N_7318);
nor U14190 (N_14190,N_7721,N_6751);
nor U14191 (N_14191,N_7827,N_5972);
xor U14192 (N_14192,N_6376,N_9334);
or U14193 (N_14193,N_7390,N_7315);
or U14194 (N_14194,N_7585,N_9672);
or U14195 (N_14195,N_7130,N_9548);
and U14196 (N_14196,N_6293,N_5980);
xnor U14197 (N_14197,N_9661,N_7130);
or U14198 (N_14198,N_8364,N_9271);
nand U14199 (N_14199,N_7028,N_9641);
nor U14200 (N_14200,N_6924,N_5197);
xor U14201 (N_14201,N_9630,N_5292);
and U14202 (N_14202,N_8692,N_6072);
nor U14203 (N_14203,N_7391,N_8217);
or U14204 (N_14204,N_8951,N_7770);
and U14205 (N_14205,N_6583,N_6214);
nor U14206 (N_14206,N_7034,N_6860);
nor U14207 (N_14207,N_7457,N_5936);
nor U14208 (N_14208,N_5184,N_9590);
nand U14209 (N_14209,N_9874,N_8884);
and U14210 (N_14210,N_6916,N_7494);
nand U14211 (N_14211,N_8554,N_8082);
or U14212 (N_14212,N_7596,N_7122);
nor U14213 (N_14213,N_7183,N_7437);
and U14214 (N_14214,N_6517,N_7037);
nand U14215 (N_14215,N_8967,N_5038);
nand U14216 (N_14216,N_5070,N_6767);
nor U14217 (N_14217,N_7306,N_9413);
or U14218 (N_14218,N_5335,N_5356);
nor U14219 (N_14219,N_9765,N_9154);
nand U14220 (N_14220,N_8602,N_7150);
and U14221 (N_14221,N_7917,N_6050);
nor U14222 (N_14222,N_9369,N_8196);
or U14223 (N_14223,N_8718,N_7378);
nor U14224 (N_14224,N_5570,N_5603);
or U14225 (N_14225,N_6900,N_9749);
or U14226 (N_14226,N_7846,N_5564);
nor U14227 (N_14227,N_6678,N_6892);
xnor U14228 (N_14228,N_5892,N_6085);
nand U14229 (N_14229,N_6638,N_7756);
nor U14230 (N_14230,N_6196,N_7990);
nor U14231 (N_14231,N_7005,N_9616);
nand U14232 (N_14232,N_9511,N_6305);
and U14233 (N_14233,N_7683,N_6284);
nand U14234 (N_14234,N_9631,N_9901);
nand U14235 (N_14235,N_5681,N_5237);
or U14236 (N_14236,N_7367,N_7049);
nor U14237 (N_14237,N_8205,N_6422);
nand U14238 (N_14238,N_7820,N_7536);
nor U14239 (N_14239,N_7965,N_5256);
or U14240 (N_14240,N_5855,N_5510);
nand U14241 (N_14241,N_8186,N_8045);
nand U14242 (N_14242,N_6815,N_6385);
or U14243 (N_14243,N_7014,N_7031);
nand U14244 (N_14244,N_6417,N_6049);
or U14245 (N_14245,N_5192,N_7252);
nand U14246 (N_14246,N_8172,N_8780);
and U14247 (N_14247,N_9833,N_8392);
or U14248 (N_14248,N_5191,N_7746);
or U14249 (N_14249,N_7668,N_9999);
or U14250 (N_14250,N_5640,N_7379);
or U14251 (N_14251,N_7996,N_6057);
nand U14252 (N_14252,N_8622,N_7909);
nor U14253 (N_14253,N_5847,N_9519);
and U14254 (N_14254,N_5398,N_6453);
xnor U14255 (N_14255,N_5578,N_5497);
and U14256 (N_14256,N_5236,N_5475);
nor U14257 (N_14257,N_8324,N_6635);
nor U14258 (N_14258,N_8857,N_7117);
and U14259 (N_14259,N_7767,N_7975);
xnor U14260 (N_14260,N_9021,N_5158);
and U14261 (N_14261,N_8722,N_9315);
and U14262 (N_14262,N_9509,N_5500);
or U14263 (N_14263,N_7204,N_8472);
nor U14264 (N_14264,N_9522,N_9091);
or U14265 (N_14265,N_7401,N_7664);
nand U14266 (N_14266,N_6844,N_5930);
and U14267 (N_14267,N_7869,N_7238);
or U14268 (N_14268,N_7471,N_8081);
nand U14269 (N_14269,N_7429,N_6716);
nand U14270 (N_14270,N_9516,N_9825);
and U14271 (N_14271,N_7055,N_5605);
nand U14272 (N_14272,N_7541,N_7027);
or U14273 (N_14273,N_8337,N_8126);
nand U14274 (N_14274,N_7830,N_6941);
nor U14275 (N_14275,N_5639,N_8794);
or U14276 (N_14276,N_5183,N_5288);
nor U14277 (N_14277,N_5987,N_7322);
nor U14278 (N_14278,N_9930,N_7476);
nor U14279 (N_14279,N_7357,N_7888);
nor U14280 (N_14280,N_8585,N_5475);
nand U14281 (N_14281,N_9232,N_6907);
and U14282 (N_14282,N_7164,N_9322);
or U14283 (N_14283,N_5657,N_6371);
and U14284 (N_14284,N_5637,N_6722);
nor U14285 (N_14285,N_6389,N_6279);
nor U14286 (N_14286,N_6064,N_7967);
nand U14287 (N_14287,N_7641,N_7687);
nor U14288 (N_14288,N_8934,N_5467);
nand U14289 (N_14289,N_6671,N_8911);
or U14290 (N_14290,N_8391,N_6931);
nor U14291 (N_14291,N_5024,N_6140);
or U14292 (N_14292,N_8346,N_5958);
nand U14293 (N_14293,N_7835,N_6296);
and U14294 (N_14294,N_6179,N_8344);
nor U14295 (N_14295,N_8824,N_6995);
and U14296 (N_14296,N_6265,N_5150);
nor U14297 (N_14297,N_5896,N_5679);
and U14298 (N_14298,N_8446,N_9528);
and U14299 (N_14299,N_9350,N_7732);
nor U14300 (N_14300,N_6435,N_6820);
nor U14301 (N_14301,N_9241,N_8914);
or U14302 (N_14302,N_9855,N_5597);
and U14303 (N_14303,N_7709,N_9267);
and U14304 (N_14304,N_5903,N_9698);
or U14305 (N_14305,N_6428,N_9398);
or U14306 (N_14306,N_9277,N_8787);
nand U14307 (N_14307,N_9292,N_5072);
xnor U14308 (N_14308,N_5616,N_6941);
and U14309 (N_14309,N_7999,N_6202);
nor U14310 (N_14310,N_8224,N_6181);
nor U14311 (N_14311,N_5935,N_7422);
or U14312 (N_14312,N_7139,N_6283);
nor U14313 (N_14313,N_5122,N_9492);
nand U14314 (N_14314,N_8823,N_8441);
and U14315 (N_14315,N_6844,N_8727);
xnor U14316 (N_14316,N_5461,N_7438);
nor U14317 (N_14317,N_5488,N_8691);
nand U14318 (N_14318,N_6400,N_5963);
and U14319 (N_14319,N_6789,N_6537);
nor U14320 (N_14320,N_5828,N_9350);
or U14321 (N_14321,N_9777,N_5120);
or U14322 (N_14322,N_9831,N_6186);
or U14323 (N_14323,N_8800,N_8243);
or U14324 (N_14324,N_8106,N_9419);
or U14325 (N_14325,N_5037,N_7732);
and U14326 (N_14326,N_5660,N_9263);
and U14327 (N_14327,N_5877,N_8957);
xor U14328 (N_14328,N_6537,N_7999);
nand U14329 (N_14329,N_5580,N_8235);
or U14330 (N_14330,N_9548,N_9457);
nor U14331 (N_14331,N_7275,N_8114);
and U14332 (N_14332,N_8182,N_9461);
nor U14333 (N_14333,N_7843,N_9158);
nor U14334 (N_14334,N_6175,N_6012);
nand U14335 (N_14335,N_7963,N_7601);
nor U14336 (N_14336,N_7825,N_6748);
nor U14337 (N_14337,N_6128,N_7535);
or U14338 (N_14338,N_8024,N_6074);
nand U14339 (N_14339,N_5621,N_8438);
nor U14340 (N_14340,N_9981,N_5767);
and U14341 (N_14341,N_7202,N_8852);
and U14342 (N_14342,N_6423,N_5598);
or U14343 (N_14343,N_7145,N_8310);
and U14344 (N_14344,N_7118,N_5565);
nand U14345 (N_14345,N_9173,N_5204);
xnor U14346 (N_14346,N_9401,N_9629);
nor U14347 (N_14347,N_6143,N_6311);
nor U14348 (N_14348,N_7872,N_9210);
nor U14349 (N_14349,N_7146,N_7549);
nor U14350 (N_14350,N_7255,N_9863);
and U14351 (N_14351,N_5203,N_6239);
and U14352 (N_14352,N_6950,N_5305);
or U14353 (N_14353,N_6854,N_7319);
nor U14354 (N_14354,N_6895,N_8936);
nand U14355 (N_14355,N_5066,N_7178);
and U14356 (N_14356,N_9205,N_6042);
nand U14357 (N_14357,N_5948,N_8860);
nor U14358 (N_14358,N_6354,N_6520);
or U14359 (N_14359,N_6491,N_7165);
xor U14360 (N_14360,N_6376,N_8419);
and U14361 (N_14361,N_8212,N_8790);
nand U14362 (N_14362,N_9787,N_8457);
and U14363 (N_14363,N_5219,N_8807);
nor U14364 (N_14364,N_9854,N_6194);
nor U14365 (N_14365,N_6633,N_6419);
or U14366 (N_14366,N_9837,N_9304);
nor U14367 (N_14367,N_8663,N_9925);
or U14368 (N_14368,N_8779,N_8801);
nand U14369 (N_14369,N_8956,N_7121);
nor U14370 (N_14370,N_9051,N_5239);
and U14371 (N_14371,N_8982,N_8783);
and U14372 (N_14372,N_5188,N_5448);
nand U14373 (N_14373,N_5959,N_8364);
or U14374 (N_14374,N_7757,N_8219);
nand U14375 (N_14375,N_9669,N_5564);
and U14376 (N_14376,N_6789,N_5294);
nand U14377 (N_14377,N_5615,N_6871);
nor U14378 (N_14378,N_5236,N_5468);
or U14379 (N_14379,N_7868,N_7957);
and U14380 (N_14380,N_5930,N_8058);
nand U14381 (N_14381,N_7473,N_6825);
nor U14382 (N_14382,N_8100,N_8988);
or U14383 (N_14383,N_6720,N_9138);
and U14384 (N_14384,N_9248,N_7866);
nor U14385 (N_14385,N_8813,N_7780);
and U14386 (N_14386,N_6264,N_8213);
nand U14387 (N_14387,N_5431,N_5542);
nand U14388 (N_14388,N_6363,N_9371);
nand U14389 (N_14389,N_9111,N_7300);
and U14390 (N_14390,N_5897,N_5455);
and U14391 (N_14391,N_7277,N_6884);
nand U14392 (N_14392,N_7176,N_8827);
nor U14393 (N_14393,N_7632,N_7194);
and U14394 (N_14394,N_7841,N_5015);
nor U14395 (N_14395,N_5011,N_7175);
nand U14396 (N_14396,N_5321,N_5641);
nor U14397 (N_14397,N_8294,N_8895);
or U14398 (N_14398,N_7548,N_8182);
or U14399 (N_14399,N_5630,N_9878);
nor U14400 (N_14400,N_8332,N_8068);
nor U14401 (N_14401,N_7386,N_9315);
nor U14402 (N_14402,N_6171,N_7907);
nor U14403 (N_14403,N_9257,N_9587);
nand U14404 (N_14404,N_5907,N_8622);
or U14405 (N_14405,N_9686,N_5370);
and U14406 (N_14406,N_9574,N_9536);
nor U14407 (N_14407,N_8248,N_6012);
or U14408 (N_14408,N_5919,N_6312);
xor U14409 (N_14409,N_8533,N_7637);
nor U14410 (N_14410,N_9038,N_6862);
xor U14411 (N_14411,N_7158,N_6860);
nand U14412 (N_14412,N_6627,N_9007);
or U14413 (N_14413,N_5255,N_7078);
or U14414 (N_14414,N_8624,N_9087);
and U14415 (N_14415,N_6330,N_5921);
nand U14416 (N_14416,N_9774,N_5848);
and U14417 (N_14417,N_5041,N_7390);
and U14418 (N_14418,N_7588,N_7534);
nand U14419 (N_14419,N_5794,N_5168);
nor U14420 (N_14420,N_8146,N_6670);
xnor U14421 (N_14421,N_6712,N_7840);
nand U14422 (N_14422,N_7303,N_8794);
or U14423 (N_14423,N_7089,N_8973);
or U14424 (N_14424,N_6257,N_7682);
nand U14425 (N_14425,N_9962,N_7274);
or U14426 (N_14426,N_5530,N_7528);
and U14427 (N_14427,N_6319,N_8298);
nand U14428 (N_14428,N_7399,N_8872);
nand U14429 (N_14429,N_7820,N_8380);
and U14430 (N_14430,N_8159,N_6603);
and U14431 (N_14431,N_8170,N_5769);
nor U14432 (N_14432,N_9467,N_5853);
nand U14433 (N_14433,N_5509,N_5303);
and U14434 (N_14434,N_7629,N_5403);
or U14435 (N_14435,N_5694,N_6263);
nand U14436 (N_14436,N_9594,N_6344);
nand U14437 (N_14437,N_7195,N_9785);
nor U14438 (N_14438,N_7991,N_5711);
nor U14439 (N_14439,N_5570,N_5140);
or U14440 (N_14440,N_5024,N_6628);
and U14441 (N_14441,N_5506,N_7391);
nor U14442 (N_14442,N_7738,N_9796);
or U14443 (N_14443,N_8148,N_7141);
nand U14444 (N_14444,N_6747,N_8305);
nor U14445 (N_14445,N_9608,N_5133);
or U14446 (N_14446,N_9512,N_5799);
and U14447 (N_14447,N_6471,N_8528);
nor U14448 (N_14448,N_5821,N_5484);
nand U14449 (N_14449,N_9896,N_5373);
nor U14450 (N_14450,N_6710,N_6220);
or U14451 (N_14451,N_5539,N_9766);
nor U14452 (N_14452,N_6796,N_5337);
or U14453 (N_14453,N_7851,N_7042);
and U14454 (N_14454,N_5550,N_5824);
or U14455 (N_14455,N_5562,N_9176);
and U14456 (N_14456,N_7645,N_9215);
or U14457 (N_14457,N_7428,N_8842);
xor U14458 (N_14458,N_8841,N_7093);
xor U14459 (N_14459,N_9940,N_5170);
nor U14460 (N_14460,N_6125,N_6207);
or U14461 (N_14461,N_9365,N_8800);
or U14462 (N_14462,N_7960,N_7887);
and U14463 (N_14463,N_8777,N_7145);
or U14464 (N_14464,N_5445,N_8546);
nand U14465 (N_14465,N_6434,N_7249);
or U14466 (N_14466,N_9858,N_9990);
and U14467 (N_14467,N_7505,N_7723);
nand U14468 (N_14468,N_9239,N_9572);
or U14469 (N_14469,N_9484,N_5475);
or U14470 (N_14470,N_9751,N_7812);
nand U14471 (N_14471,N_9242,N_6991);
and U14472 (N_14472,N_5251,N_7723);
nand U14473 (N_14473,N_7808,N_7715);
or U14474 (N_14474,N_6249,N_7621);
nand U14475 (N_14475,N_6433,N_9378);
and U14476 (N_14476,N_6109,N_5579);
nand U14477 (N_14477,N_9660,N_9027);
nand U14478 (N_14478,N_9122,N_6354);
nand U14479 (N_14479,N_8575,N_9915);
xor U14480 (N_14480,N_5150,N_6588);
nor U14481 (N_14481,N_8731,N_7370);
nand U14482 (N_14482,N_5741,N_6590);
and U14483 (N_14483,N_8083,N_7330);
nand U14484 (N_14484,N_9662,N_8872);
nor U14485 (N_14485,N_9690,N_9249);
nand U14486 (N_14486,N_9710,N_7230);
and U14487 (N_14487,N_9459,N_6895);
nand U14488 (N_14488,N_7217,N_6285);
nor U14489 (N_14489,N_7433,N_8092);
nor U14490 (N_14490,N_7188,N_5227);
xor U14491 (N_14491,N_8764,N_5238);
nand U14492 (N_14492,N_7396,N_7595);
nor U14493 (N_14493,N_8360,N_7490);
nor U14494 (N_14494,N_9085,N_8926);
and U14495 (N_14495,N_5479,N_6931);
nand U14496 (N_14496,N_8644,N_6256);
and U14497 (N_14497,N_6083,N_6870);
nor U14498 (N_14498,N_6628,N_5915);
xnor U14499 (N_14499,N_5211,N_7909);
or U14500 (N_14500,N_5084,N_7135);
nand U14501 (N_14501,N_9092,N_5133);
or U14502 (N_14502,N_5916,N_5834);
nand U14503 (N_14503,N_5754,N_9222);
xor U14504 (N_14504,N_5771,N_8499);
nor U14505 (N_14505,N_5149,N_6329);
xnor U14506 (N_14506,N_5507,N_7155);
xor U14507 (N_14507,N_5664,N_6911);
nand U14508 (N_14508,N_7456,N_8673);
nor U14509 (N_14509,N_9311,N_8535);
nor U14510 (N_14510,N_6431,N_6249);
or U14511 (N_14511,N_6301,N_6522);
and U14512 (N_14512,N_9898,N_8195);
nor U14513 (N_14513,N_8316,N_7389);
or U14514 (N_14514,N_5556,N_7394);
and U14515 (N_14515,N_6275,N_5689);
or U14516 (N_14516,N_7897,N_8586);
nand U14517 (N_14517,N_8412,N_5961);
xor U14518 (N_14518,N_5362,N_5882);
or U14519 (N_14519,N_9611,N_8715);
nor U14520 (N_14520,N_9672,N_7362);
and U14521 (N_14521,N_7996,N_5702);
and U14522 (N_14522,N_9700,N_6016);
or U14523 (N_14523,N_7588,N_8096);
nor U14524 (N_14524,N_5071,N_7999);
xor U14525 (N_14525,N_7964,N_9835);
or U14526 (N_14526,N_9132,N_8152);
nand U14527 (N_14527,N_9214,N_8000);
nor U14528 (N_14528,N_5309,N_8794);
nor U14529 (N_14529,N_8152,N_6963);
nor U14530 (N_14530,N_8378,N_8144);
xnor U14531 (N_14531,N_6479,N_7362);
xnor U14532 (N_14532,N_5618,N_6874);
or U14533 (N_14533,N_8104,N_8294);
nor U14534 (N_14534,N_5454,N_5594);
nand U14535 (N_14535,N_7762,N_5079);
nor U14536 (N_14536,N_5434,N_7824);
nand U14537 (N_14537,N_5238,N_9013);
nor U14538 (N_14538,N_5958,N_7517);
nand U14539 (N_14539,N_7300,N_5886);
and U14540 (N_14540,N_8576,N_8975);
nor U14541 (N_14541,N_7516,N_9813);
xor U14542 (N_14542,N_6581,N_6138);
nor U14543 (N_14543,N_5426,N_5343);
nor U14544 (N_14544,N_5512,N_6617);
nand U14545 (N_14545,N_9841,N_6401);
nor U14546 (N_14546,N_6163,N_6898);
and U14547 (N_14547,N_6073,N_6718);
xor U14548 (N_14548,N_5559,N_6251);
xor U14549 (N_14549,N_7918,N_8296);
nand U14550 (N_14550,N_8226,N_9298);
nor U14551 (N_14551,N_7622,N_8198);
nand U14552 (N_14552,N_8324,N_6767);
nor U14553 (N_14553,N_7183,N_6205);
nor U14554 (N_14554,N_8720,N_5746);
nand U14555 (N_14555,N_6287,N_7232);
nor U14556 (N_14556,N_5824,N_7098);
nor U14557 (N_14557,N_9623,N_5229);
or U14558 (N_14558,N_5007,N_5306);
nor U14559 (N_14559,N_6166,N_6035);
and U14560 (N_14560,N_9402,N_6518);
or U14561 (N_14561,N_9093,N_5468);
or U14562 (N_14562,N_7271,N_5224);
or U14563 (N_14563,N_8145,N_8962);
nor U14564 (N_14564,N_5950,N_6316);
nor U14565 (N_14565,N_8568,N_8172);
nor U14566 (N_14566,N_5267,N_9729);
or U14567 (N_14567,N_6486,N_7228);
nor U14568 (N_14568,N_6079,N_5161);
and U14569 (N_14569,N_5562,N_6602);
nor U14570 (N_14570,N_9963,N_6413);
nor U14571 (N_14571,N_8481,N_8019);
or U14572 (N_14572,N_9191,N_6397);
and U14573 (N_14573,N_9052,N_8335);
xnor U14574 (N_14574,N_9845,N_8833);
and U14575 (N_14575,N_9109,N_5558);
nand U14576 (N_14576,N_5237,N_5375);
xor U14577 (N_14577,N_5955,N_7000);
and U14578 (N_14578,N_7435,N_6362);
nor U14579 (N_14579,N_5827,N_7136);
or U14580 (N_14580,N_7300,N_5203);
nand U14581 (N_14581,N_5444,N_6526);
nor U14582 (N_14582,N_8268,N_8725);
or U14583 (N_14583,N_8295,N_6062);
or U14584 (N_14584,N_8404,N_7633);
and U14585 (N_14585,N_6764,N_8522);
nand U14586 (N_14586,N_8000,N_6095);
nor U14587 (N_14587,N_5887,N_7027);
nor U14588 (N_14588,N_6436,N_6263);
and U14589 (N_14589,N_8167,N_6507);
nor U14590 (N_14590,N_9913,N_5780);
and U14591 (N_14591,N_6120,N_5384);
nor U14592 (N_14592,N_9701,N_9503);
nand U14593 (N_14593,N_8732,N_7824);
nor U14594 (N_14594,N_5026,N_5186);
or U14595 (N_14595,N_8448,N_9812);
xnor U14596 (N_14596,N_9337,N_8033);
or U14597 (N_14597,N_5812,N_9536);
or U14598 (N_14598,N_6461,N_6001);
nor U14599 (N_14599,N_9169,N_7437);
nor U14600 (N_14600,N_9304,N_9868);
xor U14601 (N_14601,N_9862,N_9328);
nor U14602 (N_14602,N_5883,N_7460);
and U14603 (N_14603,N_7204,N_6920);
nand U14604 (N_14604,N_7495,N_8347);
or U14605 (N_14605,N_7869,N_7546);
or U14606 (N_14606,N_9479,N_5799);
or U14607 (N_14607,N_6938,N_5697);
xor U14608 (N_14608,N_8354,N_5841);
or U14609 (N_14609,N_9081,N_7311);
and U14610 (N_14610,N_6285,N_6456);
nand U14611 (N_14611,N_8042,N_5509);
and U14612 (N_14612,N_7095,N_8617);
and U14613 (N_14613,N_8655,N_5803);
nor U14614 (N_14614,N_7477,N_6927);
or U14615 (N_14615,N_9336,N_8291);
and U14616 (N_14616,N_9844,N_6044);
or U14617 (N_14617,N_9457,N_8176);
nand U14618 (N_14618,N_7190,N_9207);
or U14619 (N_14619,N_9090,N_6760);
xnor U14620 (N_14620,N_8467,N_9276);
or U14621 (N_14621,N_5753,N_7729);
nor U14622 (N_14622,N_7469,N_9241);
nor U14623 (N_14623,N_8587,N_9214);
nand U14624 (N_14624,N_8915,N_6646);
nor U14625 (N_14625,N_9456,N_5145);
or U14626 (N_14626,N_8208,N_6390);
or U14627 (N_14627,N_9069,N_7656);
or U14628 (N_14628,N_8062,N_6714);
nor U14629 (N_14629,N_6494,N_6433);
nand U14630 (N_14630,N_5891,N_8115);
nor U14631 (N_14631,N_7105,N_5651);
or U14632 (N_14632,N_6435,N_8780);
or U14633 (N_14633,N_8144,N_8223);
nand U14634 (N_14634,N_8212,N_9169);
or U14635 (N_14635,N_8940,N_7487);
and U14636 (N_14636,N_8466,N_7404);
or U14637 (N_14637,N_8035,N_9588);
nand U14638 (N_14638,N_8149,N_9705);
xor U14639 (N_14639,N_7059,N_7601);
nor U14640 (N_14640,N_8127,N_6324);
or U14641 (N_14641,N_9314,N_8377);
or U14642 (N_14642,N_8979,N_6504);
and U14643 (N_14643,N_6163,N_9103);
nor U14644 (N_14644,N_8437,N_5798);
nand U14645 (N_14645,N_8406,N_7402);
and U14646 (N_14646,N_6433,N_7667);
or U14647 (N_14647,N_9071,N_6581);
or U14648 (N_14648,N_6388,N_7077);
nand U14649 (N_14649,N_8126,N_8742);
or U14650 (N_14650,N_9109,N_7631);
xor U14651 (N_14651,N_8275,N_6412);
nand U14652 (N_14652,N_5712,N_6354);
nor U14653 (N_14653,N_9488,N_9063);
or U14654 (N_14654,N_8495,N_6495);
and U14655 (N_14655,N_5693,N_7363);
nor U14656 (N_14656,N_9124,N_9294);
xor U14657 (N_14657,N_6642,N_7007);
nand U14658 (N_14658,N_5132,N_7936);
and U14659 (N_14659,N_8838,N_5143);
nor U14660 (N_14660,N_7838,N_6640);
nand U14661 (N_14661,N_8141,N_9468);
nand U14662 (N_14662,N_8302,N_6129);
and U14663 (N_14663,N_7707,N_8041);
nor U14664 (N_14664,N_5790,N_5005);
or U14665 (N_14665,N_8328,N_7703);
nor U14666 (N_14666,N_6693,N_7551);
nor U14667 (N_14667,N_7666,N_6009);
xor U14668 (N_14668,N_5934,N_6732);
nor U14669 (N_14669,N_7133,N_6038);
nor U14670 (N_14670,N_9568,N_6333);
or U14671 (N_14671,N_7822,N_6731);
and U14672 (N_14672,N_6084,N_6851);
nor U14673 (N_14673,N_5627,N_9224);
nand U14674 (N_14674,N_7707,N_5427);
and U14675 (N_14675,N_5169,N_6872);
nor U14676 (N_14676,N_7981,N_8172);
nand U14677 (N_14677,N_6903,N_6867);
nor U14678 (N_14678,N_8276,N_7830);
and U14679 (N_14679,N_5239,N_7348);
nor U14680 (N_14680,N_8322,N_7375);
nand U14681 (N_14681,N_6572,N_7443);
nand U14682 (N_14682,N_8467,N_6470);
nor U14683 (N_14683,N_6801,N_8314);
or U14684 (N_14684,N_7401,N_8978);
nor U14685 (N_14685,N_9021,N_7781);
nor U14686 (N_14686,N_5410,N_5865);
and U14687 (N_14687,N_6739,N_6173);
or U14688 (N_14688,N_8470,N_8552);
or U14689 (N_14689,N_6897,N_6780);
nor U14690 (N_14690,N_8129,N_6464);
and U14691 (N_14691,N_9998,N_5041);
and U14692 (N_14692,N_7316,N_9558);
and U14693 (N_14693,N_6210,N_9385);
or U14694 (N_14694,N_8018,N_9652);
and U14695 (N_14695,N_6298,N_7235);
nor U14696 (N_14696,N_7411,N_5415);
xor U14697 (N_14697,N_9459,N_5581);
and U14698 (N_14698,N_6751,N_5256);
or U14699 (N_14699,N_8551,N_8913);
nor U14700 (N_14700,N_6911,N_6199);
nor U14701 (N_14701,N_7129,N_6318);
xor U14702 (N_14702,N_5689,N_7028);
nor U14703 (N_14703,N_9189,N_5355);
or U14704 (N_14704,N_8444,N_8057);
and U14705 (N_14705,N_6915,N_8635);
xor U14706 (N_14706,N_9344,N_5137);
nand U14707 (N_14707,N_9653,N_8193);
nand U14708 (N_14708,N_6496,N_6601);
xor U14709 (N_14709,N_9655,N_5660);
nor U14710 (N_14710,N_6338,N_6649);
and U14711 (N_14711,N_8821,N_5046);
xor U14712 (N_14712,N_7888,N_8002);
nor U14713 (N_14713,N_7093,N_8547);
xor U14714 (N_14714,N_6536,N_6432);
nand U14715 (N_14715,N_9421,N_8800);
or U14716 (N_14716,N_6758,N_6648);
nor U14717 (N_14717,N_7649,N_6984);
or U14718 (N_14718,N_6745,N_7490);
xnor U14719 (N_14719,N_6619,N_9950);
nand U14720 (N_14720,N_8698,N_9357);
and U14721 (N_14721,N_9660,N_6637);
or U14722 (N_14722,N_8860,N_6561);
or U14723 (N_14723,N_8044,N_9829);
nor U14724 (N_14724,N_7017,N_5808);
nand U14725 (N_14725,N_9353,N_8730);
nand U14726 (N_14726,N_8640,N_5724);
nand U14727 (N_14727,N_8164,N_5636);
and U14728 (N_14728,N_8493,N_8537);
nand U14729 (N_14729,N_6990,N_9064);
xor U14730 (N_14730,N_9363,N_8339);
and U14731 (N_14731,N_9279,N_8190);
or U14732 (N_14732,N_5963,N_9465);
and U14733 (N_14733,N_8228,N_9942);
nor U14734 (N_14734,N_6274,N_7514);
and U14735 (N_14735,N_7756,N_8436);
and U14736 (N_14736,N_5869,N_7990);
nor U14737 (N_14737,N_5111,N_8378);
or U14738 (N_14738,N_5812,N_9472);
nand U14739 (N_14739,N_6672,N_6858);
xnor U14740 (N_14740,N_5060,N_7432);
or U14741 (N_14741,N_8959,N_7472);
and U14742 (N_14742,N_6132,N_9753);
nand U14743 (N_14743,N_5945,N_9810);
and U14744 (N_14744,N_9006,N_6240);
nand U14745 (N_14745,N_9982,N_6723);
xnor U14746 (N_14746,N_6708,N_6211);
nand U14747 (N_14747,N_7814,N_7990);
xor U14748 (N_14748,N_6898,N_5336);
and U14749 (N_14749,N_9413,N_8128);
or U14750 (N_14750,N_6315,N_5840);
xor U14751 (N_14751,N_8841,N_7802);
nand U14752 (N_14752,N_6770,N_7443);
xor U14753 (N_14753,N_7705,N_9134);
nand U14754 (N_14754,N_8110,N_7295);
or U14755 (N_14755,N_8157,N_5714);
nor U14756 (N_14756,N_7253,N_8761);
or U14757 (N_14757,N_8598,N_6533);
or U14758 (N_14758,N_8088,N_8909);
or U14759 (N_14759,N_6358,N_8462);
xnor U14760 (N_14760,N_7789,N_5051);
or U14761 (N_14761,N_7343,N_7759);
nand U14762 (N_14762,N_9152,N_8231);
and U14763 (N_14763,N_5038,N_8924);
or U14764 (N_14764,N_7472,N_9728);
and U14765 (N_14765,N_5452,N_9791);
and U14766 (N_14766,N_8028,N_7033);
nor U14767 (N_14767,N_9948,N_9373);
nor U14768 (N_14768,N_8540,N_9704);
and U14769 (N_14769,N_6735,N_9217);
nand U14770 (N_14770,N_9566,N_9483);
or U14771 (N_14771,N_8656,N_8126);
and U14772 (N_14772,N_9082,N_9940);
nand U14773 (N_14773,N_9108,N_6583);
nand U14774 (N_14774,N_8329,N_8067);
xor U14775 (N_14775,N_5111,N_8543);
and U14776 (N_14776,N_8748,N_6505);
xor U14777 (N_14777,N_6266,N_8449);
or U14778 (N_14778,N_7818,N_5985);
and U14779 (N_14779,N_8686,N_6556);
nor U14780 (N_14780,N_5255,N_8310);
and U14781 (N_14781,N_9595,N_6596);
xor U14782 (N_14782,N_6692,N_9589);
nor U14783 (N_14783,N_8309,N_7909);
xor U14784 (N_14784,N_5639,N_8647);
or U14785 (N_14785,N_5744,N_9445);
nor U14786 (N_14786,N_6339,N_7736);
nand U14787 (N_14787,N_7265,N_9975);
xor U14788 (N_14788,N_6741,N_9160);
or U14789 (N_14789,N_9607,N_5576);
nor U14790 (N_14790,N_5970,N_9574);
nand U14791 (N_14791,N_5224,N_8703);
nand U14792 (N_14792,N_7014,N_5529);
or U14793 (N_14793,N_9063,N_8806);
or U14794 (N_14794,N_7254,N_9606);
nand U14795 (N_14795,N_7722,N_9272);
nand U14796 (N_14796,N_9626,N_5057);
or U14797 (N_14797,N_9596,N_5837);
nand U14798 (N_14798,N_7385,N_8609);
and U14799 (N_14799,N_7462,N_6590);
and U14800 (N_14800,N_7774,N_5650);
nand U14801 (N_14801,N_6214,N_8611);
and U14802 (N_14802,N_6552,N_5285);
or U14803 (N_14803,N_8720,N_8513);
nor U14804 (N_14804,N_9780,N_7164);
nor U14805 (N_14805,N_8780,N_8654);
or U14806 (N_14806,N_6531,N_7226);
nor U14807 (N_14807,N_7003,N_8807);
nand U14808 (N_14808,N_5083,N_9715);
and U14809 (N_14809,N_7223,N_7447);
and U14810 (N_14810,N_5081,N_6397);
nand U14811 (N_14811,N_6409,N_5325);
nor U14812 (N_14812,N_6560,N_5365);
nand U14813 (N_14813,N_5505,N_8262);
and U14814 (N_14814,N_7263,N_6474);
nand U14815 (N_14815,N_9072,N_9327);
or U14816 (N_14816,N_9488,N_5495);
nor U14817 (N_14817,N_8735,N_6738);
and U14818 (N_14818,N_7579,N_8417);
nand U14819 (N_14819,N_8043,N_8320);
and U14820 (N_14820,N_5731,N_9718);
or U14821 (N_14821,N_9746,N_5940);
nand U14822 (N_14822,N_7545,N_6877);
nand U14823 (N_14823,N_8722,N_9191);
nand U14824 (N_14824,N_9734,N_5763);
or U14825 (N_14825,N_9270,N_7891);
nor U14826 (N_14826,N_6238,N_6261);
and U14827 (N_14827,N_8800,N_5091);
nor U14828 (N_14828,N_8258,N_9813);
nand U14829 (N_14829,N_8496,N_5499);
and U14830 (N_14830,N_6080,N_6645);
nand U14831 (N_14831,N_6887,N_7430);
nand U14832 (N_14832,N_8741,N_7627);
nand U14833 (N_14833,N_9339,N_9495);
or U14834 (N_14834,N_6916,N_7702);
and U14835 (N_14835,N_6550,N_7740);
or U14836 (N_14836,N_9187,N_6450);
nor U14837 (N_14837,N_9040,N_9346);
or U14838 (N_14838,N_6782,N_5842);
nand U14839 (N_14839,N_8735,N_5902);
and U14840 (N_14840,N_7643,N_5102);
or U14841 (N_14841,N_8387,N_7573);
nand U14842 (N_14842,N_9845,N_5786);
nand U14843 (N_14843,N_5694,N_7528);
and U14844 (N_14844,N_8419,N_5229);
nand U14845 (N_14845,N_8412,N_5364);
nand U14846 (N_14846,N_5421,N_6173);
nor U14847 (N_14847,N_8934,N_6364);
nand U14848 (N_14848,N_8284,N_8964);
and U14849 (N_14849,N_8918,N_7187);
or U14850 (N_14850,N_5829,N_6594);
nand U14851 (N_14851,N_9183,N_6686);
nor U14852 (N_14852,N_7093,N_6112);
and U14853 (N_14853,N_9902,N_5821);
and U14854 (N_14854,N_7077,N_8920);
xnor U14855 (N_14855,N_7414,N_8683);
nor U14856 (N_14856,N_7081,N_6624);
and U14857 (N_14857,N_9124,N_6343);
nor U14858 (N_14858,N_5455,N_8946);
and U14859 (N_14859,N_7813,N_9944);
nand U14860 (N_14860,N_7402,N_6641);
xnor U14861 (N_14861,N_7661,N_5240);
xor U14862 (N_14862,N_5668,N_9818);
nor U14863 (N_14863,N_9821,N_9662);
nor U14864 (N_14864,N_8905,N_9532);
or U14865 (N_14865,N_6921,N_7072);
and U14866 (N_14866,N_6545,N_5396);
or U14867 (N_14867,N_5505,N_6457);
xnor U14868 (N_14868,N_8642,N_6879);
nand U14869 (N_14869,N_8549,N_5100);
nand U14870 (N_14870,N_8896,N_9686);
and U14871 (N_14871,N_5154,N_6886);
or U14872 (N_14872,N_9675,N_5523);
nor U14873 (N_14873,N_8409,N_5872);
and U14874 (N_14874,N_8863,N_7014);
nor U14875 (N_14875,N_8863,N_5238);
or U14876 (N_14876,N_5252,N_8675);
or U14877 (N_14877,N_9132,N_8564);
and U14878 (N_14878,N_8824,N_6203);
and U14879 (N_14879,N_8437,N_8495);
and U14880 (N_14880,N_8415,N_7745);
nor U14881 (N_14881,N_9112,N_5904);
nand U14882 (N_14882,N_7159,N_5533);
nand U14883 (N_14883,N_7023,N_9135);
or U14884 (N_14884,N_9420,N_7329);
nand U14885 (N_14885,N_7809,N_6506);
nand U14886 (N_14886,N_9775,N_8743);
xor U14887 (N_14887,N_9137,N_9686);
and U14888 (N_14888,N_7376,N_8680);
xnor U14889 (N_14889,N_5743,N_9257);
xor U14890 (N_14890,N_9054,N_6697);
nor U14891 (N_14891,N_6329,N_5802);
nand U14892 (N_14892,N_9713,N_6882);
nand U14893 (N_14893,N_7502,N_5427);
or U14894 (N_14894,N_5765,N_6444);
or U14895 (N_14895,N_5349,N_5155);
xor U14896 (N_14896,N_8732,N_5141);
and U14897 (N_14897,N_5056,N_9362);
xnor U14898 (N_14898,N_9683,N_9495);
xnor U14899 (N_14899,N_6434,N_9206);
or U14900 (N_14900,N_9097,N_6181);
nor U14901 (N_14901,N_5169,N_5924);
or U14902 (N_14902,N_5313,N_7325);
nor U14903 (N_14903,N_9457,N_6165);
and U14904 (N_14904,N_7270,N_8303);
and U14905 (N_14905,N_5550,N_9672);
nand U14906 (N_14906,N_6091,N_5174);
or U14907 (N_14907,N_6972,N_6663);
or U14908 (N_14908,N_9659,N_7047);
nor U14909 (N_14909,N_7377,N_8793);
nor U14910 (N_14910,N_9075,N_8532);
nor U14911 (N_14911,N_9756,N_8485);
nand U14912 (N_14912,N_6412,N_9905);
nor U14913 (N_14913,N_6667,N_8627);
nor U14914 (N_14914,N_9686,N_8335);
xor U14915 (N_14915,N_5507,N_6273);
and U14916 (N_14916,N_6780,N_5857);
nor U14917 (N_14917,N_8092,N_6485);
xor U14918 (N_14918,N_8984,N_6150);
nor U14919 (N_14919,N_9580,N_7476);
and U14920 (N_14920,N_6778,N_7629);
nand U14921 (N_14921,N_8960,N_6249);
or U14922 (N_14922,N_5674,N_7131);
nor U14923 (N_14923,N_8366,N_9141);
or U14924 (N_14924,N_9543,N_5211);
and U14925 (N_14925,N_6218,N_6132);
nand U14926 (N_14926,N_9630,N_9011);
nand U14927 (N_14927,N_7943,N_5978);
nand U14928 (N_14928,N_9350,N_7572);
nand U14929 (N_14929,N_9575,N_6059);
nor U14930 (N_14930,N_8154,N_5190);
xnor U14931 (N_14931,N_8684,N_5592);
and U14932 (N_14932,N_5945,N_6662);
nor U14933 (N_14933,N_9537,N_9600);
nand U14934 (N_14934,N_6750,N_5138);
and U14935 (N_14935,N_9616,N_5776);
xnor U14936 (N_14936,N_5260,N_8880);
or U14937 (N_14937,N_5791,N_8539);
nand U14938 (N_14938,N_9910,N_6431);
nor U14939 (N_14939,N_8964,N_6934);
or U14940 (N_14940,N_7890,N_7715);
nand U14941 (N_14941,N_9050,N_8327);
or U14942 (N_14942,N_6988,N_8553);
nor U14943 (N_14943,N_6491,N_8032);
nor U14944 (N_14944,N_6824,N_8289);
or U14945 (N_14945,N_8196,N_6143);
and U14946 (N_14946,N_6272,N_8391);
xnor U14947 (N_14947,N_8389,N_9042);
nand U14948 (N_14948,N_9923,N_7468);
and U14949 (N_14949,N_9224,N_7502);
nor U14950 (N_14950,N_8186,N_7079);
xnor U14951 (N_14951,N_9588,N_6339);
and U14952 (N_14952,N_9551,N_9744);
and U14953 (N_14953,N_6984,N_8994);
or U14954 (N_14954,N_9747,N_5576);
or U14955 (N_14955,N_6184,N_8111);
nand U14956 (N_14956,N_8682,N_5620);
or U14957 (N_14957,N_5342,N_5848);
nand U14958 (N_14958,N_8639,N_7632);
and U14959 (N_14959,N_8994,N_8524);
or U14960 (N_14960,N_8672,N_8298);
and U14961 (N_14961,N_6524,N_8591);
xor U14962 (N_14962,N_6905,N_8110);
or U14963 (N_14963,N_8388,N_8161);
and U14964 (N_14964,N_7625,N_6353);
nand U14965 (N_14965,N_5525,N_7477);
or U14966 (N_14966,N_8326,N_5446);
or U14967 (N_14967,N_6944,N_7024);
and U14968 (N_14968,N_7832,N_5083);
and U14969 (N_14969,N_5350,N_7202);
nand U14970 (N_14970,N_6259,N_7492);
nand U14971 (N_14971,N_7622,N_8874);
and U14972 (N_14972,N_6410,N_9236);
nor U14973 (N_14973,N_6372,N_8084);
or U14974 (N_14974,N_7336,N_6189);
or U14975 (N_14975,N_7443,N_7583);
or U14976 (N_14976,N_9779,N_7670);
nor U14977 (N_14977,N_7186,N_5362);
or U14978 (N_14978,N_6592,N_5518);
nor U14979 (N_14979,N_7257,N_9069);
or U14980 (N_14980,N_6590,N_9557);
nand U14981 (N_14981,N_7073,N_6212);
and U14982 (N_14982,N_6298,N_9530);
nand U14983 (N_14983,N_6592,N_7760);
or U14984 (N_14984,N_9234,N_7575);
nor U14985 (N_14985,N_5301,N_5836);
xor U14986 (N_14986,N_5838,N_7253);
nand U14987 (N_14987,N_7456,N_8584);
nand U14988 (N_14988,N_8185,N_7205);
or U14989 (N_14989,N_9822,N_9814);
xnor U14990 (N_14990,N_5967,N_7414);
or U14991 (N_14991,N_5953,N_6735);
nor U14992 (N_14992,N_7154,N_8116);
or U14993 (N_14993,N_7145,N_9393);
nand U14994 (N_14994,N_5452,N_8879);
or U14995 (N_14995,N_7074,N_8208);
nand U14996 (N_14996,N_9511,N_5831);
and U14997 (N_14997,N_5449,N_6108);
nor U14998 (N_14998,N_8224,N_5454);
nor U14999 (N_14999,N_9819,N_9775);
nor U15000 (N_15000,N_10673,N_11199);
or U15001 (N_15001,N_13769,N_12244);
nor U15002 (N_15002,N_10613,N_12710);
or U15003 (N_15003,N_13872,N_13469);
xnor U15004 (N_15004,N_12917,N_14622);
nand U15005 (N_15005,N_14030,N_10454);
nand U15006 (N_15006,N_14756,N_11045);
and U15007 (N_15007,N_10269,N_11367);
nand U15008 (N_15008,N_12181,N_13235);
nor U15009 (N_15009,N_14658,N_12110);
or U15010 (N_15010,N_12236,N_12163);
or U15011 (N_15011,N_10261,N_14791);
and U15012 (N_15012,N_12472,N_11815);
xnor U15013 (N_15013,N_14455,N_14090);
nor U15014 (N_15014,N_13299,N_13520);
or U15015 (N_15015,N_12176,N_13077);
or U15016 (N_15016,N_11703,N_14017);
nor U15017 (N_15017,N_13193,N_13923);
or U15018 (N_15018,N_12873,N_14394);
or U15019 (N_15019,N_13924,N_12752);
and U15020 (N_15020,N_14713,N_14126);
or U15021 (N_15021,N_13699,N_12449);
nand U15022 (N_15022,N_11166,N_13435);
nor U15023 (N_15023,N_13312,N_14200);
nand U15024 (N_15024,N_10243,N_12211);
and U15025 (N_15025,N_11223,N_11531);
xnor U15026 (N_15026,N_11306,N_13362);
or U15027 (N_15027,N_13969,N_14101);
nor U15028 (N_15028,N_13373,N_14241);
nor U15029 (N_15029,N_13115,N_12495);
nor U15030 (N_15030,N_13968,N_10048);
and U15031 (N_15031,N_13619,N_13411);
nor U15032 (N_15032,N_12898,N_13735);
nand U15033 (N_15033,N_10817,N_12773);
nor U15034 (N_15034,N_10918,N_13212);
and U15035 (N_15035,N_10207,N_13948);
or U15036 (N_15036,N_13987,N_10850);
and U15037 (N_15037,N_13484,N_10272);
or U15038 (N_15038,N_13124,N_11101);
nand U15039 (N_15039,N_14240,N_11858);
xnor U15040 (N_15040,N_13117,N_13454);
and U15041 (N_15041,N_12154,N_14239);
nand U15042 (N_15042,N_11609,N_10390);
nor U15043 (N_15043,N_14122,N_12708);
nor U15044 (N_15044,N_14108,N_13204);
nand U15045 (N_15045,N_12237,N_12706);
nor U15046 (N_15046,N_12668,N_13874);
nor U15047 (N_15047,N_10432,N_12200);
or U15048 (N_15048,N_11336,N_11911);
xor U15049 (N_15049,N_13947,N_14326);
and U15050 (N_15050,N_14714,N_10450);
nand U15051 (N_15051,N_13630,N_12278);
nor U15052 (N_15052,N_12908,N_12552);
nand U15053 (N_15053,N_10080,N_10268);
or U15054 (N_15054,N_10433,N_12334);
xnor U15055 (N_15055,N_10139,N_13870);
and U15056 (N_15056,N_13096,N_11125);
or U15057 (N_15057,N_13816,N_14105);
and U15058 (N_15058,N_11744,N_14013);
or U15059 (N_15059,N_13988,N_14439);
nand U15060 (N_15060,N_12796,N_10363);
nor U15061 (N_15061,N_14115,N_11186);
or U15062 (N_15062,N_13094,N_14798);
or U15063 (N_15063,N_13216,N_13171);
and U15064 (N_15064,N_11242,N_11152);
and U15065 (N_15065,N_10977,N_12214);
xnor U15066 (N_15066,N_10019,N_12989);
nand U15067 (N_15067,N_11022,N_14540);
or U15068 (N_15068,N_11096,N_10560);
or U15069 (N_15069,N_13669,N_10287);
nand U15070 (N_15070,N_11277,N_11628);
and U15071 (N_15071,N_14972,N_12024);
xor U15072 (N_15072,N_12604,N_11780);
xor U15073 (N_15073,N_13965,N_12974);
nand U15074 (N_15074,N_12539,N_14515);
or U15075 (N_15075,N_12043,N_13943);
nor U15076 (N_15076,N_10506,N_14176);
nor U15077 (N_15077,N_11740,N_10930);
nand U15078 (N_15078,N_10836,N_11134);
nor U15079 (N_15079,N_13028,N_10769);
nand U15080 (N_15080,N_12153,N_14334);
and U15081 (N_15081,N_11091,N_12367);
nor U15082 (N_15082,N_11322,N_14116);
nand U15083 (N_15083,N_14818,N_13062);
or U15084 (N_15084,N_14372,N_10777);
and U15085 (N_15085,N_12500,N_12084);
nor U15086 (N_15086,N_12112,N_10968);
nand U15087 (N_15087,N_13333,N_11801);
nand U15088 (N_15088,N_11481,N_14926);
or U15089 (N_15089,N_11592,N_10767);
nor U15090 (N_15090,N_12714,N_11455);
and U15091 (N_15091,N_11939,N_11368);
and U15092 (N_15092,N_13175,N_13695);
nand U15093 (N_15093,N_12197,N_10759);
and U15094 (N_15094,N_10205,N_11908);
and U15095 (N_15095,N_11857,N_11817);
nand U15096 (N_15096,N_12879,N_11039);
nand U15097 (N_15097,N_12213,N_14128);
and U15098 (N_15098,N_13169,N_11002);
nor U15099 (N_15099,N_13668,N_11820);
nor U15100 (N_15100,N_11454,N_12527);
nor U15101 (N_15101,N_12355,N_13080);
or U15102 (N_15102,N_11855,N_12032);
nor U15103 (N_15103,N_14891,N_14205);
or U15104 (N_15104,N_11754,N_11494);
xnor U15105 (N_15105,N_14485,N_13319);
and U15106 (N_15106,N_12279,N_13718);
and U15107 (N_15107,N_11221,N_12443);
and U15108 (N_15108,N_14221,N_10928);
and U15109 (N_15109,N_12115,N_12800);
nand U15110 (N_15110,N_10385,N_11729);
and U15111 (N_15111,N_14596,N_10748);
nand U15112 (N_15112,N_12113,N_11109);
nor U15113 (N_15113,N_11582,N_10374);
xnor U15114 (N_15114,N_12673,N_11293);
xnor U15115 (N_15115,N_13102,N_13545);
nor U15116 (N_15116,N_14511,N_13754);
nor U15117 (N_15117,N_13645,N_13772);
or U15118 (N_15118,N_14025,N_13883);
and U15119 (N_15119,N_12344,N_13900);
and U15120 (N_15120,N_10305,N_14007);
nand U15121 (N_15121,N_10805,N_14857);
or U15122 (N_15122,N_13765,N_11225);
and U15123 (N_15123,N_14016,N_10111);
and U15124 (N_15124,N_12466,N_10648);
and U15125 (N_15125,N_11053,N_12223);
nand U15126 (N_15126,N_13258,N_14768);
and U15127 (N_15127,N_12903,N_14933);
or U15128 (N_15128,N_10612,N_10213);
nand U15129 (N_15129,N_11347,N_10940);
and U15130 (N_15130,N_10659,N_11049);
nand U15131 (N_15131,N_13489,N_13250);
and U15132 (N_15132,N_12838,N_14359);
or U15133 (N_15133,N_11499,N_11951);
nand U15134 (N_15134,N_14453,N_13123);
or U15135 (N_15135,N_11844,N_13353);
or U15136 (N_15136,N_13606,N_12654);
nor U15137 (N_15137,N_12476,N_13954);
xor U15138 (N_15138,N_14387,N_11120);
and U15139 (N_15139,N_11567,N_11162);
and U15140 (N_15140,N_10907,N_11493);
and U15141 (N_15141,N_11520,N_14996);
nand U15142 (N_15142,N_14968,N_12304);
nand U15143 (N_15143,N_13082,N_12240);
nor U15144 (N_15144,N_12378,N_14406);
and U15145 (N_15145,N_10933,N_13676);
xor U15146 (N_15146,N_12293,N_14093);
or U15147 (N_15147,N_12263,N_12326);
or U15148 (N_15148,N_12194,N_13902);
and U15149 (N_15149,N_14973,N_14158);
nand U15150 (N_15150,N_11505,N_10253);
nor U15151 (N_15151,N_13823,N_14988);
nand U15152 (N_15152,N_10278,N_12106);
and U15153 (N_15153,N_10566,N_13949);
and U15154 (N_15154,N_10837,N_14276);
nor U15155 (N_15155,N_13329,N_14047);
and U15156 (N_15156,N_13561,N_14644);
nor U15157 (N_15157,N_10472,N_11771);
and U15158 (N_15158,N_10999,N_11661);
nand U15159 (N_15159,N_10168,N_13832);
or U15160 (N_15160,N_13109,N_14464);
and U15161 (N_15161,N_14552,N_11321);
nor U15162 (N_15162,N_13683,N_14048);
nor U15163 (N_15163,N_10224,N_12008);
nor U15164 (N_15164,N_14665,N_13631);
or U15165 (N_15165,N_10250,N_14517);
and U15166 (N_15166,N_12207,N_12645);
nand U15167 (N_15167,N_14398,N_11615);
nand U15168 (N_15168,N_13126,N_10979);
nand U15169 (N_15169,N_13746,N_11249);
and U15170 (N_15170,N_13156,N_14626);
or U15171 (N_15171,N_14340,N_13600);
nor U15172 (N_15172,N_11178,N_13733);
or U15173 (N_15173,N_12306,N_10470);
nor U15174 (N_15174,N_10097,N_13449);
or U15175 (N_15175,N_11102,N_14569);
nor U15176 (N_15176,N_14590,N_10617);
or U15177 (N_15177,N_14365,N_14850);
and U15178 (N_15178,N_12322,N_11851);
nand U15179 (N_15179,N_14646,N_10564);
nand U15180 (N_15180,N_10897,N_10255);
and U15181 (N_15181,N_10707,N_11430);
or U15182 (N_15182,N_14170,N_13195);
nand U15183 (N_15183,N_13448,N_12795);
or U15184 (N_15184,N_11324,N_14703);
nor U15185 (N_15185,N_10187,N_14623);
and U15186 (N_15186,N_12749,N_12486);
or U15187 (N_15187,N_11804,N_11589);
xor U15188 (N_15188,N_10165,N_11822);
xnor U15189 (N_15189,N_11960,N_12740);
or U15190 (N_15190,N_13681,N_10804);
and U15191 (N_15191,N_13432,N_13744);
nand U15192 (N_15192,N_14929,N_14630);
or U15193 (N_15193,N_10592,N_10295);
nand U15194 (N_15194,N_11721,N_14373);
nand U15195 (N_15195,N_14449,N_13912);
nor U15196 (N_15196,N_12190,N_10307);
or U15197 (N_15197,N_13091,N_11876);
nand U15198 (N_15198,N_14556,N_10280);
nor U15199 (N_15199,N_12380,N_11241);
nor U15200 (N_15200,N_14120,N_13065);
and U15201 (N_15201,N_12369,N_14290);
or U15202 (N_15202,N_12191,N_14705);
nor U15203 (N_15203,N_14099,N_12063);
and U15204 (N_15204,N_13950,N_12125);
or U15205 (N_15205,N_10462,N_10012);
nand U15206 (N_15206,N_13566,N_11218);
xnor U15207 (N_15207,N_14846,N_14469);
nor U15208 (N_15208,N_12285,N_14548);
or U15209 (N_15209,N_12597,N_14295);
nor U15210 (N_15210,N_13305,N_11651);
or U15211 (N_15211,N_14306,N_12062);
or U15212 (N_15212,N_11445,N_10246);
xnor U15213 (N_15213,N_11147,N_11196);
nor U15214 (N_15214,N_12399,N_13058);
nand U15215 (N_15215,N_14015,N_12626);
xor U15216 (N_15216,N_11312,N_11233);
xnor U15217 (N_15217,N_12068,N_10885);
or U15218 (N_15218,N_13723,N_14506);
xor U15219 (N_15219,N_12392,N_10082);
nor U15220 (N_15220,N_11818,N_10285);
or U15221 (N_15221,N_10720,N_12571);
nand U15222 (N_15222,N_10591,N_11912);
and U15223 (N_15223,N_10848,N_11366);
and U15224 (N_15224,N_12360,N_10007);
nor U15225 (N_15225,N_12958,N_14881);
nand U15226 (N_15226,N_13188,N_11061);
nor U15227 (N_15227,N_14849,N_11172);
or U15228 (N_15228,N_12672,N_10072);
xor U15229 (N_15229,N_11441,N_10142);
and U15230 (N_15230,N_14234,N_10154);
or U15231 (N_15231,N_13464,N_14650);
or U15232 (N_15232,N_12828,N_10944);
and U15233 (N_15233,N_13575,N_11633);
or U15234 (N_15234,N_14616,N_10294);
nor U15235 (N_15235,N_12761,N_10271);
or U15236 (N_15236,N_10115,N_11301);
or U15237 (N_15237,N_10729,N_11700);
or U15238 (N_15238,N_12577,N_12479);
or U15239 (N_15239,N_11411,N_11971);
and U15240 (N_15240,N_10533,N_13673);
xor U15241 (N_15241,N_14952,N_14530);
xnor U15242 (N_15242,N_12620,N_13849);
nor U15243 (N_15243,N_13989,N_12915);
nor U15244 (N_15244,N_14168,N_12388);
nand U15245 (N_15245,N_12241,N_10137);
or U15246 (N_15246,N_13180,N_12047);
or U15247 (N_15247,N_11214,N_10889);
nand U15248 (N_15248,N_12418,N_10881);
nand U15249 (N_15249,N_14994,N_12333);
and U15250 (N_15250,N_10976,N_10676);
nand U15251 (N_15251,N_11565,N_11252);
nand U15252 (N_15252,N_10449,N_10430);
nand U15253 (N_15253,N_10531,N_11545);
or U15254 (N_15254,N_14056,N_13395);
nor U15255 (N_15255,N_11581,N_11507);
xor U15256 (N_15256,N_13326,N_13045);
nand U15257 (N_15257,N_11590,N_11536);
or U15258 (N_15258,N_12452,N_11970);
and U15259 (N_15259,N_14829,N_13296);
xnor U15260 (N_15260,N_13589,N_10290);
or U15261 (N_15261,N_11638,N_10415);
or U15262 (N_15262,N_11933,N_10672);
or U15263 (N_15263,N_11261,N_12255);
nand U15264 (N_15264,N_13056,N_10909);
nand U15265 (N_15265,N_12807,N_11522);
and U15266 (N_15266,N_11583,N_13907);
or U15267 (N_15267,N_11605,N_10608);
nor U15268 (N_15268,N_14903,N_14139);
nand U15269 (N_15269,N_10380,N_14858);
nor U15270 (N_15270,N_12349,N_12808);
xnor U15271 (N_15271,N_10267,N_13654);
nand U15272 (N_15272,N_12069,N_11396);
and U15273 (N_15273,N_12489,N_10521);
nand U15274 (N_15274,N_10943,N_13026);
nand U15275 (N_15275,N_14539,N_14774);
nand U15276 (N_15276,N_12442,N_11681);
nand U15277 (N_15277,N_13088,N_12018);
nand U15278 (N_15278,N_11268,N_12126);
xnor U15279 (N_15279,N_12957,N_10038);
nand U15280 (N_15280,N_11269,N_13856);
and U15281 (N_15281,N_12187,N_14252);
or U15282 (N_15282,N_13953,N_14213);
and U15283 (N_15283,N_14493,N_10429);
and U15284 (N_15284,N_14243,N_11334);
or U15285 (N_15285,N_14663,N_10320);
or U15286 (N_15286,N_13453,N_10393);
nor U15287 (N_15287,N_11956,N_10838);
or U15288 (N_15288,N_13984,N_12703);
nand U15289 (N_15289,N_13829,N_10279);
and U15290 (N_15290,N_11325,N_14619);
xnor U15291 (N_15291,N_12600,N_13626);
and U15292 (N_15292,N_14327,N_10394);
nor U15293 (N_15293,N_11976,N_10742);
or U15294 (N_15294,N_12079,N_13380);
nand U15295 (N_15295,N_10581,N_13431);
and U15296 (N_15296,N_13703,N_12394);
or U15297 (N_15297,N_13029,N_13404);
or U15298 (N_15298,N_14296,N_10459);
nor U15299 (N_15299,N_13926,N_12912);
xnor U15300 (N_15300,N_12017,N_14987);
nand U15301 (N_15301,N_12423,N_10972);
xor U15302 (N_15302,N_13106,N_14608);
nand U15303 (N_15303,N_10630,N_11916);
nand U15304 (N_15304,N_13410,N_10003);
or U15305 (N_15305,N_11953,N_10806);
nor U15306 (N_15306,N_13551,N_13531);
nand U15307 (N_15307,N_13384,N_10514);
xnor U15308 (N_15308,N_12254,N_11275);
or U15309 (N_15309,N_14341,N_10799);
nand U15310 (N_15310,N_12765,N_12720);
nand U15311 (N_15311,N_11862,N_13491);
nand U15312 (N_15312,N_12872,N_12189);
or U15313 (N_15313,N_10441,N_14046);
nand U15314 (N_15314,N_10411,N_14164);
and U15315 (N_15315,N_10780,N_11436);
or U15316 (N_15316,N_14347,N_12325);
nor U15317 (N_15317,N_11920,N_10391);
and U15318 (N_15318,N_11094,N_14141);
or U15319 (N_15319,N_11263,N_12955);
or U15320 (N_15320,N_14712,N_13402);
nor U15321 (N_15321,N_12104,N_10217);
nand U15322 (N_15322,N_12891,N_14599);
nor U15323 (N_15323,N_12914,N_10347);
and U15324 (N_15324,N_12054,N_10695);
nand U15325 (N_15325,N_10776,N_12789);
nand U15326 (N_15326,N_12031,N_14487);
nor U15327 (N_15327,N_10067,N_12101);
xor U15328 (N_15328,N_10831,N_13934);
nor U15329 (N_15329,N_10008,N_13658);
or U15330 (N_15330,N_10254,N_14148);
and U15331 (N_15331,N_13320,N_12435);
nand U15332 (N_15332,N_13660,N_12586);
nand U15333 (N_15333,N_14825,N_10901);
and U15334 (N_15334,N_13191,N_14757);
or U15335 (N_15335,N_11926,N_11099);
or U15336 (N_15336,N_13539,N_13137);
nor U15337 (N_15337,N_14042,N_12239);
nor U15338 (N_15338,N_10702,N_10632);
xnor U15339 (N_15339,N_12858,N_11563);
xnor U15340 (N_15340,N_14900,N_14685);
xor U15341 (N_15341,N_13141,N_12221);
or U15342 (N_15342,N_14345,N_10016);
xor U15343 (N_15343,N_14331,N_13875);
nand U15344 (N_15344,N_13621,N_14632);
and U15345 (N_15345,N_12338,N_10801);
nor U15346 (N_15346,N_14754,N_10475);
nor U15347 (N_15347,N_11137,N_11831);
nor U15348 (N_15348,N_12158,N_13827);
or U15349 (N_15349,N_11165,N_10884);
nor U15350 (N_15350,N_12471,N_14543);
xnor U15351 (N_15351,N_13293,N_10700);
nand U15352 (N_15352,N_12493,N_10824);
nor U15353 (N_15353,N_14131,N_14109);
nor U15354 (N_15354,N_12432,N_14415);
or U15355 (N_15355,N_12459,N_12738);
xnor U15356 (N_15356,N_11824,N_12837);
nand U15357 (N_15357,N_12389,N_11397);
and U15358 (N_15358,N_13519,N_13921);
or U15359 (N_15359,N_13151,N_12260);
nor U15360 (N_15360,N_12643,N_10021);
nand U15361 (N_15361,N_14209,N_13379);
or U15362 (N_15362,N_10237,N_11755);
nor U15363 (N_15363,N_11897,N_10163);
nor U15364 (N_15364,N_10823,N_10827);
nand U15365 (N_15365,N_14027,N_12948);
nand U15366 (N_15366,N_10456,N_12929);
nor U15367 (N_15367,N_12532,N_12582);
nor U15368 (N_15368,N_10491,N_14005);
or U15369 (N_15369,N_14309,N_13544);
and U15370 (N_15370,N_14708,N_12875);
and U15371 (N_15371,N_14861,N_14593);
and U15372 (N_15372,N_11577,N_11281);
or U15373 (N_15373,N_12270,N_14594);
nand U15374 (N_15374,N_14643,N_10571);
nand U15375 (N_15375,N_11266,N_14664);
and U15376 (N_15376,N_14877,N_12759);
xnor U15377 (N_15377,N_14725,N_14424);
or U15378 (N_15378,N_12843,N_13939);
nand U15379 (N_15379,N_10505,N_13121);
nand U15380 (N_15380,N_11435,N_12557);
and U15381 (N_15381,N_13226,N_12617);
and U15382 (N_15382,N_11018,N_14244);
nor U15383 (N_15383,N_12232,N_11035);
or U15384 (N_15384,N_10228,N_11111);
nand U15385 (N_15385,N_12743,N_14925);
nor U15386 (N_15386,N_10387,N_14481);
nand U15387 (N_15387,N_10525,N_10828);
and U15388 (N_15388,N_12072,N_12767);
and U15389 (N_15389,N_14130,N_10882);
or U15390 (N_15390,N_11059,N_13716);
and U15391 (N_15391,N_12777,N_14161);
or U15392 (N_15392,N_12209,N_11827);
xnor U15393 (N_15393,N_13898,N_12854);
nor U15394 (N_15394,N_11323,N_10225);
xnor U15395 (N_15395,N_11751,N_14367);
xor U15396 (N_15396,N_10716,N_10557);
and U15397 (N_15397,N_13130,N_13807);
nand U15398 (N_15398,N_10910,N_13063);
nor U15399 (N_15399,N_13689,N_10326);
nor U15400 (N_15400,N_13656,N_12004);
or U15401 (N_15401,N_12817,N_13521);
or U15402 (N_15402,N_12461,N_12889);
nor U15403 (N_15403,N_14760,N_14807);
and U15404 (N_15404,N_14173,N_11770);
and U15405 (N_15405,N_14716,N_14982);
and U15406 (N_15406,N_13280,N_10408);
and U15407 (N_15407,N_11087,N_12460);
xor U15408 (N_15408,N_11072,N_13494);
or U15409 (N_15409,N_14719,N_10855);
nand U15410 (N_15410,N_11255,N_14834);
xor U15411 (N_15411,N_11805,N_13433);
and U15412 (N_15412,N_13998,N_14470);
and U15413 (N_15413,N_10196,N_12066);
or U15414 (N_15414,N_13603,N_13976);
or U15415 (N_15415,N_10622,N_10148);
or U15416 (N_15416,N_14856,N_13576);
xnor U15417 (N_15417,N_11062,N_13790);
and U15418 (N_15418,N_13623,N_13777);
nand U15419 (N_15419,N_10350,N_11919);
nor U15420 (N_15420,N_10922,N_10410);
nor U15421 (N_15421,N_14747,N_14274);
or U15422 (N_15422,N_13580,N_14237);
nand U15423 (N_15423,N_13582,N_11787);
or U15424 (N_15424,N_12457,N_12906);
and U15425 (N_15425,N_12121,N_14318);
nand U15426 (N_15426,N_13248,N_10234);
and U15427 (N_15427,N_13496,N_11127);
or U15428 (N_15428,N_14946,N_14136);
nand U15429 (N_15429,N_11378,N_10114);
or U15430 (N_15430,N_13985,N_13006);
or U15431 (N_15431,N_12511,N_13284);
or U15432 (N_15432,N_14041,N_12971);
nor U15433 (N_15433,N_14518,N_11380);
nor U15434 (N_15434,N_10001,N_11341);
nand U15435 (N_15435,N_14202,N_14541);
nand U15436 (N_15436,N_10034,N_10760);
or U15437 (N_15437,N_12206,N_14495);
nor U15438 (N_15438,N_14986,N_10102);
nor U15439 (N_15439,N_14381,N_13766);
nand U15440 (N_15440,N_12734,N_10083);
or U15441 (N_15441,N_14266,N_10685);
xnor U15442 (N_15442,N_11007,N_10956);
xnor U15443 (N_15443,N_10989,N_11727);
or U15444 (N_15444,N_12770,N_12313);
nand U15445 (N_15445,N_12416,N_12936);
nand U15446 (N_15446,N_14098,N_13878);
and U15447 (N_15447,N_10994,N_11264);
and U15448 (N_15448,N_12398,N_10146);
nor U15449 (N_15449,N_11361,N_12138);
nor U15450 (N_15450,N_14782,N_13110);
and U15451 (N_15451,N_14640,N_10407);
nand U15452 (N_15452,N_11044,N_12810);
and U15453 (N_15453,N_13515,N_13279);
nand U15454 (N_15454,N_11027,N_14745);
nand U15455 (N_15455,N_14353,N_12878);
nor U15456 (N_15456,N_12433,N_13750);
and U15457 (N_15457,N_10706,N_11174);
nand U15458 (N_15458,N_13436,N_11946);
nor U15459 (N_15459,N_12947,N_11644);
nor U15460 (N_15460,N_13684,N_10311);
xnor U15461 (N_15461,N_13879,N_10657);
xnor U15462 (N_15462,N_12542,N_14840);
nor U15463 (N_15463,N_14806,N_13225);
nand U15464 (N_15464,N_10084,N_10844);
and U15465 (N_15465,N_10815,N_11071);
and U15466 (N_15466,N_13046,N_11699);
nand U15467 (N_15467,N_12308,N_10852);
nor U15468 (N_15468,N_10569,N_10719);
and U15469 (N_15469,N_14302,N_14003);
xor U15470 (N_15470,N_10949,N_14860);
nor U15471 (N_15471,N_13249,N_12051);
or U15472 (N_15472,N_12099,N_13557);
nor U15473 (N_15473,N_12167,N_11540);
nor U15474 (N_15474,N_10483,N_12847);
or U15475 (N_15475,N_14299,N_10973);
nand U15476 (N_15476,N_10444,N_13134);
or U15477 (N_15477,N_11560,N_13705);
xnor U15478 (N_15478,N_14033,N_10442);
and U15479 (N_15479,N_12377,N_11259);
xor U15480 (N_15480,N_12477,N_10574);
nand U15481 (N_15481,N_12353,N_12140);
nor U15482 (N_15482,N_11429,N_13335);
nor U15483 (N_15483,N_11549,N_13271);
nor U15484 (N_15484,N_14267,N_11154);
and U15485 (N_15485,N_12042,N_14962);
or U15486 (N_15486,N_10174,N_11433);
nand U15487 (N_15487,N_14668,N_13970);
nand U15488 (N_15488,N_14242,N_10666);
and U15489 (N_15489,N_12337,N_11232);
and U15490 (N_15490,N_11200,N_10826);
xnor U15491 (N_15491,N_13955,N_12135);
or U15492 (N_15492,N_14710,N_12548);
and U15493 (N_15493,N_10967,N_10895);
and U15494 (N_15494,N_13559,N_14699);
and U15495 (N_15495,N_11843,N_11904);
or U15496 (N_15496,N_11905,N_11442);
xnor U15497 (N_15497,N_14675,N_12614);
nand U15498 (N_15498,N_12746,N_12856);
or U15499 (N_15499,N_11486,N_11370);
nor U15500 (N_15500,N_11459,N_11997);
or U15501 (N_15501,N_13022,N_12161);
nand U15502 (N_15502,N_10610,N_12390);
or U15503 (N_15503,N_12632,N_11955);
nor U15504 (N_15504,N_13510,N_11273);
nor U15505 (N_15505,N_10351,N_10291);
and U15506 (N_15506,N_10431,N_10919);
or U15507 (N_15507,N_13414,N_13325);
or U15508 (N_15508,N_14826,N_12218);
and U15509 (N_15509,N_12311,N_12453);
and U15510 (N_15510,N_12372,N_14654);
or U15511 (N_15511,N_14859,N_11641);
nor U15512 (N_15512,N_12259,N_10299);
and U15513 (N_15513,N_11769,N_13928);
nor U15514 (N_15514,N_12976,N_10779);
xor U15515 (N_15515,N_12094,N_11034);
nand U15516 (N_15516,N_13524,N_11957);
and U15517 (N_15517,N_12309,N_12677);
xor U15518 (N_15518,N_12913,N_10671);
and U15519 (N_15519,N_13543,N_12327);
and U15520 (N_15520,N_14437,N_11298);
and U15521 (N_15521,N_14395,N_12547);
xnor U15522 (N_15522,N_12258,N_10558);
and U15523 (N_15523,N_12805,N_10405);
xnor U15524 (N_15524,N_10161,N_10770);
nand U15525 (N_15525,N_12001,N_14475);
or U15526 (N_15526,N_14088,N_12646);
nor U15527 (N_15527,N_12177,N_12085);
and U15528 (N_15528,N_13583,N_12899);
nor U15529 (N_15529,N_10732,N_11716);
nor U15530 (N_15530,N_10315,N_11709);
or U15531 (N_15531,N_10133,N_10825);
nor U15532 (N_15532,N_11216,N_10646);
or U15533 (N_15533,N_14023,N_13107);
nor U15534 (N_15534,N_11508,N_11776);
nand U15535 (N_15535,N_14065,N_12690);
and U15536 (N_15536,N_14790,N_13771);
nand U15537 (N_15537,N_13203,N_14927);
nor U15538 (N_15538,N_10588,N_10499);
and U15539 (N_15539,N_11652,N_11379);
xor U15540 (N_15540,N_12490,N_12991);
or U15541 (N_15541,N_12011,N_12419);
nor U15542 (N_15542,N_11236,N_14162);
and U15543 (N_15543,N_13111,N_13644);
nand U15544 (N_15544,N_10413,N_12385);
nand U15545 (N_15545,N_10232,N_10076);
nor U15546 (N_15546,N_12774,N_10236);
nor U15547 (N_15547,N_10175,N_13506);
nor U15548 (N_15548,N_14503,N_14913);
or U15549 (N_15549,N_13680,N_10379);
xor U15550 (N_15550,N_13711,N_13157);
and U15551 (N_15551,N_14468,N_10681);
xor U15552 (N_15552,N_12514,N_11885);
xor U15553 (N_15553,N_11757,N_13906);
nand U15554 (N_15554,N_10763,N_10262);
nor U15555 (N_15555,N_12397,N_12825);
and U15556 (N_15556,N_11662,N_10766);
nand U15557 (N_15557,N_10370,N_13796);
and U15558 (N_15558,N_13336,N_10868);
and U15559 (N_15559,N_12682,N_12470);
nor U15560 (N_15560,N_11313,N_13588);
and U15561 (N_15561,N_13323,N_10155);
nand U15562 (N_15562,N_10414,N_11689);
and U15563 (N_15563,N_14906,N_12363);
nor U15564 (N_15564,N_13895,N_13133);
and U15565 (N_15565,N_12375,N_10573);
nand U15566 (N_15566,N_13294,N_12864);
xor U15567 (N_15567,N_10069,N_11832);
nand U15568 (N_15568,N_11637,N_10814);
nor U15569 (N_15569,N_12533,N_14074);
and U15570 (N_15570,N_14546,N_11934);
or U15571 (N_15571,N_12735,N_14809);
nor U15572 (N_15572,N_13812,N_13382);
or U15573 (N_15573,N_14392,N_11248);
nor U15574 (N_15574,N_14966,N_14905);
nand U15575 (N_15575,N_11654,N_13528);
or U15576 (N_15576,N_14967,N_12117);
nor U15577 (N_15577,N_11555,N_11085);
and U15578 (N_15578,N_11449,N_10210);
or U15579 (N_15579,N_13562,N_11910);
nand U15580 (N_15580,N_11875,N_14547);
and U15581 (N_15581,N_14283,N_10756);
nand U15582 (N_15582,N_13140,N_13143);
xor U15583 (N_15583,N_12077,N_10039);
xnor U15584 (N_15584,N_14414,N_12585);
nand U15585 (N_15585,N_12147,N_14236);
or U15586 (N_15586,N_12426,N_10006);
xor U15587 (N_15587,N_11409,N_11895);
nand U15588 (N_15588,N_12709,N_14814);
and U15589 (N_15589,N_10173,N_14902);
and U15590 (N_15590,N_14978,N_13908);
and U15591 (N_15591,N_10728,N_13000);
nand U15592 (N_15592,N_11686,N_14896);
or U15593 (N_15593,N_10869,N_11081);
and U15594 (N_15594,N_12376,N_13886);
nor U15595 (N_15595,N_12935,N_14736);
nand U15596 (N_15596,N_11251,N_11863);
nand U15597 (N_15597,N_13548,N_13797);
nand U15598 (N_15598,N_14607,N_10835);
xor U15599 (N_15599,N_11142,N_10085);
or U15600 (N_15600,N_11896,N_12998);
nand U15601 (N_15601,N_11639,N_12474);
or U15602 (N_15602,N_11777,N_11672);
nor U15603 (N_15603,N_13670,N_13138);
and U15604 (N_15604,N_10229,N_12904);
nand U15605 (N_15605,N_11033,N_10131);
xnor U15606 (N_15606,N_11140,N_13762);
nor U15607 (N_15607,N_10157,N_13932);
or U15608 (N_15608,N_13956,N_11945);
xnor U15609 (N_15609,N_14634,N_10495);
or U15610 (N_15610,N_14735,N_13227);
xnor U15611 (N_15611,N_10552,N_12166);
or U15612 (N_15612,N_12169,N_12446);
nand U15613 (N_15613,N_13257,N_12421);
nand U15614 (N_15614,N_12465,N_13577);
nor U15615 (N_15615,N_10810,N_12835);
nor U15616 (N_15616,N_12107,N_10747);
or U15617 (N_15617,N_12642,N_10313);
or U15618 (N_15618,N_11538,N_12718);
and U15619 (N_15619,N_14106,N_10458);
or U15620 (N_15620,N_10954,N_12257);
and U15621 (N_15621,N_14508,N_10709);
nand U15622 (N_15622,N_10561,N_14275);
nand U15623 (N_15623,N_14879,N_12216);
and U15624 (N_15624,N_12573,N_13002);
nor U15625 (N_15625,N_12657,N_14971);
nand U15626 (N_15626,N_11962,N_14513);
nor U15627 (N_15627,N_12717,N_12801);
and U15628 (N_15628,N_12782,N_12995);
and U15629 (N_15629,N_12132,N_12314);
or U15630 (N_15630,N_10812,N_13590);
nor U15631 (N_15631,N_10231,N_11778);
nand U15632 (N_15632,N_12275,N_10145);
or U15633 (N_15633,N_13330,N_11393);
or U15634 (N_15634,N_14730,N_14217);
nor U15635 (N_15635,N_12521,N_13666);
nor U15636 (N_15636,N_14738,N_10037);
nor U15637 (N_15637,N_10463,N_10896);
and U15638 (N_15638,N_10266,N_14947);
and U15639 (N_15639,N_14270,N_11124);
nor U15640 (N_15640,N_12702,N_13334);
or U15641 (N_15641,N_10600,N_11270);
nand U15642 (N_15642,N_12243,N_13715);
and U15643 (N_15643,N_13690,N_12316);
xor U15644 (N_15644,N_12950,N_12885);
xor U15645 (N_15645,N_12594,N_11803);
xor U15646 (N_15646,N_12612,N_11463);
or U15647 (N_15647,N_14459,N_10009);
and U15648 (N_15648,N_14399,N_14944);
or U15649 (N_15649,N_12492,N_11523);
and U15650 (N_15650,N_12096,N_11451);
or U15651 (N_15651,N_12984,N_10092);
or U15652 (N_15652,N_12860,N_12053);
or U15653 (N_15653,N_10772,N_14097);
nor U15654 (N_15654,N_10665,N_14951);
xor U15655 (N_15655,N_10138,N_14509);
and U15656 (N_15656,N_12227,N_11052);
xnor U15657 (N_15657,N_12679,N_11276);
nor U15658 (N_15658,N_10615,N_10015);
nor U15659 (N_15659,N_14921,N_11422);
xor U15660 (N_15660,N_11420,N_11892);
and U15661 (N_15661,N_12458,N_12088);
or U15662 (N_15662,N_13087,N_10962);
and U15663 (N_15663,N_14854,N_12622);
nand U15664 (N_15664,N_10579,N_12250);
nand U15665 (N_15665,N_11942,N_13304);
nand U15666 (N_15666,N_13977,N_13833);
nor U15667 (N_15667,N_14995,N_14779);
or U15668 (N_15668,N_10670,N_13122);
nand U15669 (N_15669,N_13911,N_13930);
nand U15670 (N_15670,N_10022,N_12097);
xnor U15671 (N_15671,N_12619,N_13706);
nand U15672 (N_15672,N_12238,N_13393);
nor U15673 (N_15673,N_12319,N_13781);
nor U15674 (N_15674,N_11679,N_13406);
or U15675 (N_15675,N_11929,N_13183);
nand U15676 (N_15676,N_13759,N_11989);
nor U15677 (N_15677,N_10527,N_12226);
and U15678 (N_15678,N_14476,N_14784);
xor U15679 (N_15679,N_12969,N_14303);
xnor U15680 (N_15680,N_11682,N_11917);
xor U15681 (N_15681,N_12134,N_13422);
nand U15682 (N_15682,N_14095,N_10443);
nand U15683 (N_15683,N_11714,N_11217);
and U15684 (N_15684,N_12256,N_13347);
or U15685 (N_15685,N_10186,N_13952);
and U15686 (N_15686,N_11842,N_14885);
nand U15687 (N_15687,N_14498,N_11690);
or U15688 (N_15688,N_14452,N_12882);
or U15689 (N_15689,N_11013,N_13881);
and U15690 (N_15690,N_14839,N_11228);
and U15691 (N_15691,N_11413,N_14742);
xnor U15692 (N_15692,N_13890,N_14410);
nor U15693 (N_15693,N_13846,N_14497);
nand U15694 (N_15694,N_13337,N_12901);
nand U15695 (N_15695,N_14103,N_12498);
and U15696 (N_15696,N_10822,N_14053);
and U15697 (N_15697,N_10843,N_10086);
xor U15698 (N_15698,N_14561,N_11256);
and U15699 (N_15699,N_14195,N_13154);
nor U15700 (N_15700,N_12785,N_13262);
and U15701 (N_15701,N_14659,N_11741);
and U15702 (N_15702,N_12509,N_10589);
nand U15703 (N_15703,N_10093,N_11054);
or U15704 (N_15704,N_14291,N_14936);
and U15705 (N_15705,N_10545,N_11100);
and U15706 (N_15706,N_11834,N_11304);
nand U15707 (N_15707,N_14051,N_13773);
and U15708 (N_15708,N_12328,N_11297);
nand U15709 (N_15709,N_11537,N_13937);
nor U15710 (N_15710,N_12468,N_14637);
nor U15711 (N_15711,N_14955,N_12370);
or U15712 (N_15712,N_11408,N_11491);
or U15713 (N_15713,N_10577,N_10235);
nor U15714 (N_15714,N_10947,N_13256);
and U15715 (N_15715,N_11927,N_12719);
and U15716 (N_15716,N_12436,N_14491);
nand U15717 (N_15717,N_13946,N_13447);
and U15718 (N_15718,N_11728,N_11175);
or U15719 (N_15719,N_11374,N_11031);
and U15720 (N_15720,N_10209,N_14631);
xnor U15721 (N_15721,N_10556,N_14224);
nand U15722 (N_15722,N_11496,N_11462);
nand U15723 (N_15723,N_12420,N_10540);
nand U15724 (N_15724,N_10400,N_14284);
nor U15725 (N_15725,N_13692,N_14778);
and U15726 (N_15726,N_11009,N_13471);
xnor U15727 (N_15727,N_12918,N_11881);
nand U15728 (N_15728,N_14562,N_11395);
or U15729 (N_15729,N_10892,N_10158);
nor U15730 (N_15730,N_11246,N_12507);
or U15731 (N_15731,N_13370,N_12451);
or U15732 (N_15732,N_13542,N_11381);
xor U15733 (N_15733,N_12647,N_10180);
or U15734 (N_15734,N_14125,N_13073);
and U15735 (N_15735,N_13611,N_13052);
or U15736 (N_15736,N_10689,N_10866);
nand U15737 (N_15737,N_14928,N_11114);
nand U15738 (N_15738,N_13150,N_11000);
nor U15739 (N_15739,N_11287,N_14420);
nand U15740 (N_15740,N_11873,N_11731);
nand U15741 (N_15741,N_10360,N_12040);
nand U15742 (N_15742,N_10136,N_10511);
nor U15743 (N_15743,N_10028,N_12407);
nor U15744 (N_15744,N_11572,N_13713);
and U15745 (N_15745,N_14032,N_10105);
or U15746 (N_15746,N_10974,N_12979);
nor U15747 (N_15747,N_14633,N_13776);
or U15748 (N_15748,N_14819,N_13612);
nor U15749 (N_15749,N_12638,N_12545);
nor U15750 (N_15750,N_13255,N_12298);
xor U15751 (N_15751,N_10507,N_13741);
nand U15752 (N_15752,N_11653,N_10597);
or U15753 (N_15753,N_13231,N_11781);
or U15754 (N_15754,N_14034,N_13297);
nor U15755 (N_15755,N_11030,N_10674);
nor U15756 (N_15756,N_12350,N_12525);
nor U15757 (N_15757,N_14157,N_14629);
and U15758 (N_15758,N_14843,N_13570);
nor U15759 (N_15759,N_14525,N_13473);
or U15760 (N_15760,N_11558,N_13498);
nand U15761 (N_15761,N_13245,N_10258);
and U15762 (N_15762,N_13011,N_14134);
and U15763 (N_15763,N_14196,N_10669);
and U15764 (N_15764,N_11475,N_11220);
nand U15765 (N_15765,N_13514,N_11095);
and U15766 (N_15766,N_11850,N_13780);
nor U15767 (N_15767,N_14211,N_11128);
and U15768 (N_15768,N_13477,N_14524);
and U15769 (N_15769,N_10460,N_13529);
nor U15770 (N_15770,N_13345,N_10273);
nor U15771 (N_15771,N_11088,N_11838);
and U15772 (N_15772,N_11510,N_13131);
nor U15773 (N_15773,N_14889,N_12895);
or U15774 (N_15774,N_13821,N_13731);
nor U15775 (N_15775,N_11280,N_13913);
or U15776 (N_15776,N_14815,N_10333);
and U15777 (N_15777,N_11618,N_11513);
and U15778 (N_15778,N_10151,N_11206);
nand U15779 (N_15779,N_13381,N_14389);
nor U15780 (N_15780,N_11743,N_14149);
or U15781 (N_15781,N_12151,N_11438);
nand U15782 (N_15782,N_13556,N_11290);
and U15783 (N_15783,N_10964,N_14649);
nor U15784 (N_15784,N_12529,N_13775);
or U15785 (N_15785,N_14953,N_10398);
nand U15786 (N_15786,N_14432,N_10281);
and U15787 (N_15787,N_13685,N_10886);
nand U15788 (N_15788,N_14336,N_13209);
nand U15789 (N_15789,N_13128,N_14467);
nand U15790 (N_15790,N_13001,N_11415);
and U15791 (N_15791,N_10782,N_13646);
nand U15792 (N_15792,N_11504,N_10796);
and U15793 (N_15793,N_12414,N_13072);
nand U15794 (N_15794,N_12359,N_14273);
and U15795 (N_15795,N_14666,N_12295);
and U15796 (N_15796,N_10289,N_12683);
nand U15797 (N_15797,N_14606,N_12219);
or U15798 (N_15798,N_13343,N_11471);
and U15799 (N_15799,N_13567,N_10058);
and U15800 (N_15800,N_11764,N_14451);
nand U15801 (N_15801,N_12960,N_12114);
or U15802 (N_15802,N_14899,N_14465);
nor U15803 (N_15803,N_12300,N_12804);
nor U15804 (N_15804,N_14915,N_11302);
and U15805 (N_15805,N_12932,N_14679);
nand U15806 (N_15806,N_11474,N_11739);
or U15807 (N_15807,N_10578,N_12540);
nand U15808 (N_15808,N_13704,N_13550);
and U15809 (N_15809,N_11344,N_14067);
nor U15810 (N_15810,N_10355,N_10959);
nand U15811 (N_15811,N_10744,N_10951);
nor U15812 (N_15812,N_10240,N_11527);
xor U15813 (N_15813,N_14144,N_13592);
or U15814 (N_15814,N_11327,N_14479);
or U15815 (N_15815,N_14715,N_11584);
nand U15816 (N_15816,N_10134,N_12431);
and U15817 (N_15817,N_13564,N_12520);
xor U15818 (N_15818,N_14939,N_12776);
nand U15819 (N_15819,N_10502,N_13555);
nor U15820 (N_15820,N_11785,N_10354);
nand U15821 (N_15821,N_11219,N_10265);
xnor U15822 (N_15822,N_10768,N_14797);
nand U15823 (N_15823,N_11038,N_11613);
nor U15824 (N_15824,N_12141,N_12160);
and U15825 (N_15825,N_11423,N_10986);
or U15826 (N_15826,N_13317,N_13709);
nand U15827 (N_15827,N_11333,N_12120);
and U15828 (N_15828,N_11187,N_14300);
and U15829 (N_15829,N_13217,N_11529);
or U15830 (N_15830,N_14227,N_12623);
nor U15831 (N_15831,N_10375,N_10226);
or U15832 (N_15832,N_12265,N_12616);
xnor U15833 (N_15833,N_13119,N_14938);
xor U15834 (N_15834,N_14499,N_11133);
or U15835 (N_15835,N_11867,N_14773);
nand U15836 (N_15836,N_11201,N_11819);
nor U15837 (N_15837,N_13324,N_11469);
and U15838 (N_15838,N_14647,N_14893);
xnor U15839 (N_15839,N_13516,N_14752);
xor U15840 (N_15840,N_14656,N_14618);
nor U15841 (N_15841,N_12822,N_14458);
or U15842 (N_15842,N_14932,N_13120);
nor U15843 (N_15843,N_10629,N_13980);
or U15844 (N_15844,N_14882,N_10089);
nand U15845 (N_15845,N_14305,N_13752);
nor U15846 (N_15846,N_13173,N_14949);
nor U15847 (N_15847,N_14364,N_14132);
and U15848 (N_15848,N_11318,N_12893);
nand U15849 (N_15849,N_12515,N_14189);
nor U15850 (N_15850,N_10975,N_10208);
nor U15851 (N_15851,N_14911,N_10122);
or U15852 (N_15852,N_13758,N_13268);
or U15853 (N_15853,N_10509,N_14294);
nand U15854 (N_15854,N_12644,N_13213);
nand U15855 (N_15855,N_11614,N_11710);
nand U15856 (N_15856,N_14864,N_12754);
and U15857 (N_15857,N_11169,N_13363);
nor U15858 (N_15858,N_14642,N_11573);
and U15859 (N_15859,N_14280,N_10905);
nand U15860 (N_15860,N_10467,N_14639);
nand U15861 (N_15861,N_12384,N_12793);
and U15862 (N_15862,N_14603,N_10296);
xor U15863 (N_15863,N_13184,N_14700);
nor U15864 (N_15864,N_13041,N_14070);
and U15865 (N_15865,N_13272,N_13224);
or U15866 (N_15866,N_14028,N_12425);
xnor U15867 (N_15867,N_11417,N_12182);
and U15868 (N_15868,N_10170,N_10337);
nor U15869 (N_15869,N_12315,N_10125);
or U15870 (N_15870,N_12756,N_13620);
nor U15871 (N_15871,N_10714,N_11680);
nor U15872 (N_15872,N_14887,N_12408);
xor U15873 (N_15873,N_11105,N_11561);
or U15874 (N_15874,N_12144,N_13664);
and U15875 (N_15875,N_12082,N_13700);
and U15876 (N_15876,N_12651,N_11328);
or U15877 (N_15877,N_14442,N_12694);
or U15878 (N_15878,N_13500,N_11427);
nor U15879 (N_15879,N_14072,N_11535);
and U15880 (N_15880,N_14076,N_10535);
or U15881 (N_15881,N_11056,N_11702);
or U15882 (N_15882,N_11258,N_13013);
or U15883 (N_15883,N_10582,N_12233);
and U15884 (N_15884,N_11996,N_12519);
xor U15885 (N_15885,N_13865,N_13694);
nand U15886 (N_15886,N_11267,N_14999);
nor U15887 (N_15887,N_13321,N_10300);
or U15888 (N_15888,N_13308,N_14792);
xnor U15889 (N_15889,N_12676,N_10202);
xor U15890 (N_15890,N_13025,N_14954);
and U15891 (N_15891,N_13513,N_10338);
nand U15892 (N_15892,N_12480,N_12092);
nand U15893 (N_15893,N_11398,N_14535);
nand U15894 (N_15894,N_14904,N_10087);
and U15895 (N_15895,N_14054,N_13597);
nand U15896 (N_15896,N_13152,N_13230);
or U15897 (N_15897,N_12943,N_14684);
and U15898 (N_15898,N_10854,N_11807);
and U15899 (N_15899,N_13147,N_14998);
nor U15900 (N_15900,N_12578,N_14897);
xnor U15901 (N_15901,N_13067,N_11182);
nor U15902 (N_15902,N_11720,N_13434);
or U15903 (N_15903,N_13220,N_14055);
and U15904 (N_15904,N_11426,N_14426);
nand U15905 (N_15905,N_11452,N_12297);
nor U15906 (N_15906,N_12572,N_12444);
nand U15907 (N_15907,N_12745,N_10377);
nand U15908 (N_15908,N_13309,N_13791);
nor U15909 (N_15909,N_10875,N_11608);
nor U15910 (N_15910,N_14147,N_14580);
nor U15911 (N_15911,N_11136,N_12558);
or U15912 (N_15912,N_13896,N_12021);
nand U15913 (N_15913,N_11570,N_14941);
or U15914 (N_15914,N_14869,N_10830);
nor U15915 (N_15915,N_12924,N_12366);
and U15916 (N_15916,N_14040,N_14313);
xnor U15917 (N_15917,N_13457,N_14335);
and U15918 (N_15918,N_12028,N_13468);
or U15919 (N_15919,N_12930,N_13421);
and U15920 (N_15920,N_12168,N_10791);
nand U15921 (N_15921,N_13820,N_12933);
nand U15922 (N_15922,N_12965,N_11840);
or U15923 (N_15923,N_11901,N_10169);
or U15924 (N_15924,N_12173,N_10753);
and U15925 (N_15925,N_13678,N_13824);
and U15926 (N_15926,N_11213,N_13941);
nand U15927 (N_15927,N_14749,N_14124);
nand U15928 (N_15928,N_13661,N_14721);
and U15929 (N_15929,N_13331,N_14011);
and U15930 (N_15930,N_14344,N_13019);
nand U15931 (N_15931,N_12119,N_13116);
nor U15932 (N_15932,N_11148,N_10839);
or U15933 (N_15933,N_12636,N_11197);
and U15934 (N_15934,N_14876,N_13889);
or U15935 (N_15935,N_10184,N_10302);
nor U15936 (N_15936,N_10614,N_12707);
xnor U15937 (N_15937,N_13974,N_11316);
nand U15938 (N_15938,N_12273,N_14259);
nor U15939 (N_15939,N_12787,N_10635);
nand U15940 (N_15940,N_14037,N_12827);
nand U15941 (N_15941,N_12387,N_13635);
nor U15942 (N_15942,N_10953,N_12347);
and U15943 (N_15943,N_10755,N_14624);
and U15944 (N_15944,N_10902,N_12288);
and U15945 (N_15945,N_10249,N_12109);
or U15946 (N_15946,N_11578,N_11358);
nor U15947 (N_15947,N_14177,N_14729);
nor U15948 (N_15948,N_10966,N_13060);
xnor U15949 (N_15949,N_10056,N_12569);
nand U15950 (N_15950,N_13441,N_13467);
or U15951 (N_15951,N_10416,N_13888);
nor U15952 (N_15952,N_11023,N_12386);
xnor U15953 (N_15953,N_11708,N_11534);
or U15954 (N_15954,N_13289,N_11036);
or U15955 (N_15955,N_13472,N_10811);
or U15956 (N_15956,N_12902,N_11410);
or U15957 (N_15957,N_13344,N_14412);
and U15958 (N_15958,N_13069,N_11163);
nor U15959 (N_15959,N_14758,N_12345);
nor U15960 (N_15960,N_11768,N_14375);
or U15961 (N_15961,N_14817,N_11788);
or U15962 (N_15962,N_13021,N_10418);
nand U15963 (N_15963,N_13314,N_10818);
nand U15964 (N_15964,N_12127,N_11181);
or U15965 (N_15965,N_11692,N_14066);
nor U15966 (N_15966,N_14943,N_12985);
nand U15967 (N_15967,N_13160,N_10447);
xor U15968 (N_15968,N_12146,N_14142);
or U15969 (N_15969,N_13501,N_11797);
or U15970 (N_15970,N_14750,N_10113);
and U15971 (N_15971,N_14292,N_11286);
nand U15972 (N_15972,N_10453,N_12274);
or U15973 (N_15973,N_12156,N_13032);
and U15974 (N_15974,N_13729,N_11813);
or U15975 (N_15975,N_11759,N_14184);
and U15976 (N_15976,N_11664,N_12791);
and U15977 (N_15977,N_12402,N_11972);
xnor U15978 (N_15978,N_14462,N_11406);
nor U15979 (N_15979,N_11948,N_11048);
and U15980 (N_15980,N_14358,N_12551);
nor U15981 (N_15981,N_14870,N_12320);
nor U15982 (N_15982,N_10075,N_10649);
or U15983 (N_15983,N_10466,N_12248);
nor U15984 (N_15984,N_13378,N_14199);
nand U15985 (N_15985,N_13266,N_12225);
and U15986 (N_15986,N_11222,N_12071);
nand U15987 (N_15987,N_10650,N_13478);
nor U15988 (N_15988,N_14004,N_12845);
and U15989 (N_15989,N_10050,N_12852);
nor U15990 (N_15990,N_10787,N_14523);
or U15991 (N_15991,N_14583,N_14413);
or U15992 (N_15992,N_11211,N_10183);
nor U15993 (N_15993,N_11464,N_11629);
or U15994 (N_15994,N_11922,N_11084);
nand U15995 (N_15995,N_12036,N_14560);
or U15996 (N_15996,N_10162,N_10746);
xnor U15997 (N_15997,N_10104,N_10764);
and U15998 (N_15998,N_13437,N_13536);
or U15999 (N_15999,N_10199,N_12742);
nor U16000 (N_16000,N_10023,N_13038);
xnor U16001 (N_16001,N_13318,N_10642);
and U16002 (N_16002,N_13672,N_13887);
nand U16003 (N_16003,N_11852,N_11472);
or U16004 (N_16004,N_13269,N_11239);
or U16005 (N_16005,N_10389,N_12661);
or U16006 (N_16006,N_11465,N_11055);
nor U16007 (N_16007,N_10891,N_11821);
nand U16008 (N_16008,N_11458,N_14174);
or U16009 (N_16009,N_10599,N_11234);
nand U16010 (N_16010,N_14963,N_10042);
and U16011 (N_16011,N_11250,N_14255);
and U16012 (N_16012,N_13493,N_10576);
nor U16013 (N_16013,N_14557,N_14123);
and U16014 (N_16014,N_12129,N_12429);
or U16015 (N_16015,N_12262,N_14107);
and U16016 (N_16016,N_12178,N_13282);
or U16017 (N_16017,N_10678,N_12266);
xnor U16018 (N_16018,N_10925,N_10842);
nor U16019 (N_16019,N_14441,N_14969);
xor U16020 (N_16020,N_14592,N_11574);
nand U16021 (N_16021,N_10030,N_12563);
or U16022 (N_16022,N_10699,N_12133);
and U16023 (N_16023,N_13295,N_12462);
and U16024 (N_16024,N_10871,N_14605);
and U16025 (N_16025,N_10103,N_10955);
nor U16026 (N_16026,N_12006,N_11964);
and U16027 (N_16027,N_13938,N_13427);
and U16028 (N_16028,N_11514,N_14528);
or U16029 (N_16029,N_11394,N_11969);
nand U16030 (N_16030,N_14502,N_13005);
or U16031 (N_16031,N_11526,N_13721);
nand U16032 (N_16032,N_12892,N_13640);
nor U16033 (N_16033,N_11037,N_12473);
or U16034 (N_16034,N_12357,N_12130);
nor U16035 (N_16035,N_11603,N_11202);
xor U16036 (N_16036,N_13371,N_10445);
nand U16037 (N_16037,N_14324,N_11882);
and U16038 (N_16038,N_13306,N_14117);
xnor U16039 (N_16039,N_11046,N_10858);
or U16040 (N_16040,N_10304,N_12890);
nand U16041 (N_16041,N_11717,N_10620);
xnor U16042 (N_16042,N_14422,N_10684);
nand U16043 (N_16043,N_11028,N_14489);
and U16044 (N_16044,N_10011,N_14024);
nor U16045 (N_16045,N_12618,N_13356);
nor U16046 (N_16046,N_10775,N_11606);
nand U16047 (N_16047,N_11825,N_10523);
nor U16048 (N_16048,N_13535,N_10754);
nand U16049 (N_16049,N_14002,N_10957);
nand U16050 (N_16050,N_10528,N_10052);
or U16051 (N_16051,N_11802,N_14376);
nor U16052 (N_16052,N_10035,N_10733);
xnor U16053 (N_16053,N_11453,N_14851);
nand U16054 (N_16054,N_11339,N_11693);
xor U16055 (N_16055,N_14214,N_10264);
nor U16056 (N_16056,N_11146,N_12478);
nor U16057 (N_16057,N_11961,N_11938);
or U16058 (N_16058,N_11319,N_10778);
and U16059 (N_16059,N_14482,N_13232);
or U16060 (N_16060,N_11158,N_11765);
and U16061 (N_16061,N_14231,N_12635);
nand U16062 (N_16062,N_10309,N_13298);
nor U16063 (N_16063,N_11164,N_11183);
or U16064 (N_16064,N_11893,N_10563);
and U16065 (N_16065,N_12601,N_11502);
and U16066 (N_16066,N_12276,N_12699);
or U16067 (N_16067,N_10284,N_12982);
and U16068 (N_16068,N_13641,N_11375);
or U16069 (N_16069,N_10140,N_14113);
nand U16070 (N_16070,N_11300,N_11240);
nor U16071 (N_16071,N_10873,N_13290);
or U16072 (N_16072,N_14050,N_13459);
nand U16073 (N_16073,N_10929,N_14118);
and U16074 (N_16074,N_11879,N_13009);
and U16075 (N_16075,N_11029,N_13302);
or U16076 (N_16076,N_14384,N_11224);
nor U16077 (N_16077,N_14759,N_12850);
or U16078 (N_16078,N_14704,N_10306);
or U16079 (N_16079,N_11001,N_12603);
and U16080 (N_16080,N_10725,N_10623);
and U16081 (N_16081,N_11809,N_12396);
xor U16082 (N_16082,N_13397,N_13675);
and U16083 (N_16083,N_13990,N_12588);
nor U16084 (N_16084,N_12391,N_14400);
nand U16085 (N_16085,N_14150,N_14917);
or U16086 (N_16086,N_14681,N_13419);
nor U16087 (N_16087,N_10745,N_12027);
nand U16088 (N_16088,N_10032,N_13919);
or U16089 (N_16089,N_11051,N_11829);
xnor U16090 (N_16090,N_11575,N_14804);
xor U16091 (N_16091,N_12764,N_12832);
nand U16092 (N_16092,N_13742,N_13159);
nor U16093 (N_16093,N_14802,N_13186);
xor U16094 (N_16094,N_13815,N_10223);
nor U16095 (N_16095,N_10440,N_13609);
or U16096 (N_16096,N_10656,N_10476);
and U16097 (N_16097,N_12687,N_14801);
nor U16098 (N_16098,N_14094,N_11847);
or U16099 (N_16099,N_11694,N_13084);
nand U16100 (N_16100,N_13616,N_10963);
nor U16101 (N_16101,N_12354,N_11126);
or U16102 (N_16102,N_12231,N_10212);
and U16103 (N_16103,N_11155,N_12546);
nand U16104 (N_16104,N_13719,N_10639);
xnor U16105 (N_16105,N_11198,N_14614);
or U16106 (N_16106,N_14645,N_14673);
and U16107 (N_16107,N_14388,N_10538);
and U16108 (N_16108,N_11791,N_12732);
or U16109 (N_16109,N_11497,N_11665);
or U16110 (N_16110,N_13552,N_12871);
nor U16111 (N_16111,N_10583,N_11697);
or U16112 (N_16112,N_12152,N_11794);
nor U16113 (N_16113,N_12286,N_14293);
or U16114 (N_16114,N_13986,N_14059);
or U16115 (N_16115,N_11345,N_13412);
nand U16116 (N_16116,N_14609,N_14686);
and U16117 (N_16117,N_10790,N_11748);
nor U16118 (N_16118,N_11446,N_12543);
nand U16119 (N_16119,N_14360,N_11619);
and U16120 (N_16120,N_13627,N_10361);
nand U16121 (N_16121,N_10070,N_10203);
and U16122 (N_16122,N_12896,N_10053);
or U16123 (N_16123,N_10474,N_14667);
xor U16124 (N_16124,N_14155,N_11437);
and U16125 (N_16125,N_13876,N_10197);
or U16126 (N_16126,N_13967,N_14976);
or U16127 (N_16127,N_12078,N_12592);
xor U16128 (N_16128,N_14390,N_11864);
and U16129 (N_16129,N_14404,N_10937);
xor U16130 (N_16130,N_12625,N_10880);
nor U16131 (N_16131,N_11245,N_14253);
xor U16132 (N_16132,N_13207,N_11932);
or U16133 (N_16133,N_10270,N_12639);
xor U16134 (N_16134,N_11974,N_12730);
and U16135 (N_16135,N_14471,N_13853);
nor U16136 (N_16136,N_10033,N_11683);
or U16137 (N_16137,N_10308,N_14753);
nand U16138 (N_16138,N_13757,N_11798);
nor U16139 (N_16139,N_14888,N_10662);
xor U16140 (N_16140,N_11539,N_14216);
nand U16141 (N_16141,N_12271,N_11265);
nor U16142 (N_16142,N_10316,N_10924);
and U16143 (N_16143,N_11386,N_12061);
nand U16144 (N_16144,N_13399,N_10490);
nand U16145 (N_16145,N_11066,N_14997);
nor U16146 (N_16146,N_12034,N_10479);
xor U16147 (N_16147,N_11161,N_13877);
or U16148 (N_16148,N_14733,N_13578);
nand U16149 (N_16149,N_14121,N_11229);
and U16150 (N_16150,N_13918,N_11371);
nand U16151 (N_16151,N_10063,N_11532);
and U16152 (N_16152,N_12050,N_12228);
nand U16153 (N_16153,N_14153,N_11959);
and U16154 (N_16154,N_12652,N_13836);
nand U16155 (N_16155,N_12715,N_11230);
nand U16156 (N_16156,N_12724,N_12887);
or U16157 (N_16157,N_14617,N_14322);
nor U16158 (N_16158,N_13278,N_12931);
or U16159 (N_16159,N_12526,N_12811);
nand U16160 (N_16160,N_14981,N_10029);
and U16161 (N_16161,N_14542,N_13488);
or U16162 (N_16162,N_10073,N_13726);
nand U16163 (N_16163,N_10152,N_14448);
or U16164 (N_16164,N_12550,N_12868);
or U16165 (N_16165,N_14383,N_10041);
nor U16166 (N_16166,N_13935,N_11883);
or U16167 (N_16167,N_13135,N_14408);
or U16168 (N_16168,N_13819,N_10002);
nand U16169 (N_16169,N_14371,N_13774);
nand U16170 (N_16170,N_12684,N_12629);
nor U16171 (N_16171,N_13838,N_13239);
and U16172 (N_16172,N_14852,N_12111);
nor U16173 (N_16173,N_13481,N_13205);
or U16174 (N_16174,N_13261,N_10000);
and U16175 (N_16175,N_14382,N_13413);
or U16176 (N_16176,N_11706,N_10987);
and U16177 (N_16177,N_14545,N_11789);
nor U16178 (N_16178,N_10562,N_12665);
or U16179 (N_16179,N_13931,N_12229);
nor U16180 (N_16180,N_11403,N_13341);
and U16181 (N_16181,N_11026,N_10735);
nand U16182 (N_16182,N_14167,N_14549);
or U16183 (N_16183,N_13192,N_11698);
nand U16184 (N_16184,N_13055,N_14855);
nand U16185 (N_16185,N_10893,N_12090);
nor U16186 (N_16186,N_14058,N_11871);
nor U16187 (N_16187,N_10920,N_13486);
and U16188 (N_16188,N_12523,N_11515);
nor U16189 (N_16189,N_11952,N_13161);
and U16190 (N_16190,N_12401,N_10548);
or U16191 (N_16191,N_13964,N_13179);
and U16192 (N_16192,N_12865,N_10911);
or U16193 (N_16193,N_13178,N_10690);
and U16194 (N_16194,N_11704,N_14958);
nand U16195 (N_16195,N_12867,N_14576);
or U16196 (N_16196,N_12348,N_12812);
nor U16197 (N_16197,N_14942,N_11988);
and U16198 (N_16198,N_10473,N_10227);
nor U16199 (N_16199,N_11767,N_12648);
and U16200 (N_16200,N_13386,N_14538);
or U16201 (N_16201,N_11610,N_10501);
nor U16202 (N_16202,N_13842,N_13653);
and U16203 (N_16203,N_12744,N_12830);
xor U16204 (N_16204,N_14100,N_10068);
or U16205 (N_16205,N_11121,N_13914);
and U16206 (N_16206,N_11746,N_10356);
nand U16207 (N_16207,N_10065,N_10486);
and U16208 (N_16208,N_10856,N_14356);
nand U16209 (N_16209,N_14156,N_11732);
nand U16210 (N_16210,N_11994,N_13376);
nand U16211 (N_16211,N_10900,N_12996);
xor U16212 (N_16212,N_10088,N_13251);
nor U16213 (N_16213,N_11711,N_11799);
and U16214 (N_16214,N_12973,N_12324);
nand U16215 (N_16215,N_14514,N_12691);
or U16216 (N_16216,N_14014,N_13648);
xnor U16217 (N_16217,N_12869,N_14366);
or U16218 (N_16218,N_10541,N_13398);
xnor U16219 (N_16219,N_13407,N_14922);
or U16220 (N_16220,N_11479,N_10883);
xnor U16221 (N_16221,N_11015,N_13502);
and U16222 (N_16222,N_12992,N_10153);
and U16223 (N_16223,N_14289,N_10480);
or U16224 (N_16224,N_14229,N_12196);
nand U16225 (N_16225,N_10248,N_11898);
or U16226 (N_16226,N_14795,N_10821);
nand U16227 (N_16227,N_13442,N_14786);
or U16228 (N_16228,N_14320,N_14707);
and U16229 (N_16229,N_12779,N_12441);
or U16230 (N_16230,N_10329,N_13858);
nand U16231 (N_16231,N_11995,N_10679);
xnor U16232 (N_16232,N_13749,N_10403);
and U16233 (N_16233,N_10833,N_13813);
nor U16234 (N_16234,N_14628,N_12713);
and U16235 (N_16235,N_10349,N_11416);
nand U16236 (N_16236,N_11025,N_13652);
and U16237 (N_16237,N_12282,N_10123);
or U16238 (N_16238,N_11752,N_13340);
and U16239 (N_16239,N_10425,N_12427);
xor U16240 (N_16240,N_10981,N_14391);
nand U16241 (N_16241,N_14964,N_10211);
or U16242 (N_16242,N_14431,N_12670);
and U16243 (N_16243,N_14737,N_13244);
nand U16244 (N_16244,N_13174,N_13390);
nor U16245 (N_16245,N_14775,N_12839);
nand U16246 (N_16246,N_12155,N_13963);
and U16247 (N_16247,N_14082,N_11546);
or U16248 (N_16248,N_11257,N_13920);
or U16249 (N_16249,N_13843,N_13097);
nor U16250 (N_16250,N_12536,N_11305);
and U16251 (N_16251,N_14584,N_12788);
and U16252 (N_16252,N_13034,N_10182);
nand U16253 (N_16253,N_12755,N_13354);
and U16254 (N_16254,N_13808,N_13818);
or U16255 (N_16255,N_11342,N_13463);
nand U16256 (N_16256,N_12590,N_13657);
xnor U16257 (N_16257,N_11688,N_14160);
xor U16258 (N_16258,N_12222,N_11554);
or U16259 (N_16259,N_14377,N_13495);
and U16260 (N_16260,N_10376,N_14762);
nand U16261 (N_16261,N_14661,N_10970);
or U16262 (N_16262,N_14282,N_12002);
nand U16263 (N_16263,N_10036,N_11205);
and U16264 (N_16264,N_11135,N_11977);
nor U16265 (N_16265,N_14361,N_13276);
and U16266 (N_16266,N_11562,N_12919);
nor U16267 (N_16267,N_11089,N_13633);
or U16268 (N_16268,N_13346,N_10298);
xor U16269 (N_16269,N_11833,N_13665);
nor U16270 (N_16270,N_12145,N_14924);
nand U16271 (N_16271,N_10141,N_12438);
or U16272 (N_16272,N_12301,N_12180);
nand U16273 (N_16273,N_12341,N_12859);
and U16274 (N_16274,N_12075,N_14472);
xor U16275 (N_16275,N_11587,N_10539);
nor U16276 (N_16276,N_14651,N_14288);
nor U16277 (N_16277,N_11837,N_11790);
or U16278 (N_16278,N_11082,N_10870);
nor U16279 (N_16279,N_10121,N_13831);
nor U16280 (N_16280,N_12641,N_10950);
nand U16281 (N_16281,N_12076,N_12205);
or U16282 (N_16282,N_10598,N_10172);
or U16283 (N_16283,N_12164,N_10585);
xor U16284 (N_16284,N_10587,N_10619);
and U16285 (N_16285,N_11736,N_13747);
nand U16286 (N_16286,N_12143,N_11530);
nand U16287 (N_16287,N_13994,N_14660);
nand U16288 (N_16288,N_10477,N_14083);
xnor U16289 (N_16289,N_10633,N_10263);
and U16290 (N_16290,N_11670,N_11872);
or U16291 (N_16291,N_11774,N_10820);
or U16292 (N_16292,N_11548,N_13722);
xnor U16293 (N_16293,N_13057,N_12880);
or U16294 (N_16294,N_13639,N_13618);
nand U16295 (N_16295,N_13383,N_13465);
or U16296 (N_16296,N_10636,N_11580);
nand U16297 (N_16297,N_10192,N_14772);
and U16298 (N_16298,N_13415,N_13795);
nand U16299 (N_16299,N_13971,N_14490);
xnor U16300 (N_16300,N_10005,N_11738);
or U16301 (N_16301,N_10640,N_14325);
xor U16302 (N_16302,N_13901,N_10047);
nand U16303 (N_16303,N_12430,N_11060);
nor U16304 (N_16304,N_14796,N_12607);
nand U16305 (N_16305,N_13845,N_14912);
and U16306 (N_16306,N_12508,N_12044);
nor U16307 (N_16307,N_13394,N_11967);
and U16308 (N_16308,N_10879,N_11122);
nand U16309 (N_16309,N_14178,N_10624);
nor U16310 (N_16310,N_11569,N_11750);
nor U16311 (N_16311,N_13051,N_11594);
xnor U16312 (N_16312,N_14577,N_11667);
nor U16313 (N_16313,N_13208,N_14780);
nand U16314 (N_16314,N_13825,N_11511);
nor U16315 (N_16315,N_11559,N_10667);
nor U16316 (N_16316,N_12688,N_13785);
or U16317 (N_16317,N_11192,N_10605);
nor U16318 (N_16318,N_13997,N_11854);
nand U16319 (N_16319,N_13388,N_10596);
or U16320 (N_16320,N_10568,N_12203);
or U16321 (N_16321,N_10049,N_11925);
and U16322 (N_16322,N_14226,N_10200);
nor U16323 (N_16323,N_10345,N_10898);
and U16324 (N_16324,N_14883,N_14680);
nor U16325 (N_16325,N_14555,N_13401);
and U16326 (N_16326,N_14104,N_12704);
or U16327 (N_16327,N_11151,N_14423);
nand U16328 (N_16328,N_10381,N_12598);
and U16329 (N_16329,N_11928,N_10860);
nor U16330 (N_16330,N_11986,N_10946);
nand U16331 (N_16331,N_14690,N_12700);
nand U16332 (N_16332,N_12513,N_13247);
and U16333 (N_16333,N_14337,N_10251);
nand U16334 (N_16334,N_12428,N_12518);
nor U16335 (N_16335,N_13105,N_11991);
or U16336 (N_16336,N_13806,N_13229);
nor U16337 (N_16337,N_14186,N_14683);
or U16338 (N_16338,N_11965,N_13569);
or U16339 (N_16339,N_13264,N_11231);
nor U16340 (N_16340,N_14648,N_11391);
or U16341 (N_16341,N_13839,N_11383);
and U16342 (N_16342,N_13275,N_10857);
nand U16343 (N_16343,N_10680,N_10124);
and U16344 (N_16344,N_13428,N_13525);
and U16345 (N_16345,N_10417,N_13405);
or U16346 (N_16346,N_13558,N_11640);
and U16347 (N_16347,N_13503,N_12990);
nand U16348 (N_16348,N_10851,N_11576);
xnor U16349 (N_16349,N_10980,N_14355);
and U16350 (N_16350,N_11887,N_14036);
xnor U16351 (N_16351,N_12771,N_10520);
and U16352 (N_16352,N_10095,N_10219);
nand U16353 (N_16353,N_12580,N_12159);
or U16354 (N_16354,N_13905,N_13074);
and U16355 (N_16355,N_14636,N_11058);
nor U16356 (N_16356,N_10435,N_13788);
and U16357 (N_16357,N_12975,N_13075);
nor U16358 (N_16358,N_12294,N_12666);
and U16359 (N_16359,N_12123,N_13315);
and U16360 (N_16360,N_12105,N_11707);
nand U16361 (N_16361,N_10366,N_13030);
and U16362 (N_16362,N_13581,N_13579);
nand U16363 (N_16363,N_14363,N_12000);
nand U16364 (N_16364,N_10061,N_12108);
nor U16365 (N_16365,N_12289,N_11006);
or U16366 (N_16366,N_14880,N_10752);
nor U16367 (N_16367,N_12988,N_11207);
nor U16368 (N_16368,N_14402,N_14957);
nor U16369 (N_16369,N_13707,N_11524);
or U16370 (N_16370,N_12060,N_11600);
and U16371 (N_16371,N_11890,N_12023);
xor U16372 (N_16372,N_10797,N_10572);
nor U16373 (N_16373,N_10990,N_12649);
xor U16374 (N_16374,N_14718,N_10025);
and U16375 (N_16375,N_14812,N_11992);
nor U16376 (N_16376,N_13112,N_12234);
or U16377 (N_16377,N_14368,N_14165);
xnor U16378 (N_16378,N_12570,N_11021);
and U16379 (N_16379,N_11443,N_14720);
and U16380 (N_16380,N_12696,N_10654);
nor U16381 (N_16381,N_12920,N_14440);
and U16382 (N_16382,N_12689,N_12821);
nor U16383 (N_16383,N_10693,N_12013);
and U16384 (N_16384,N_12953,N_13098);
or U16385 (N_16385,N_10983,N_10127);
or U16386 (N_16386,N_14039,N_10590);
xnor U16387 (N_16387,N_11176,N_11632);
nand U16388 (N_16388,N_13814,N_12581);
nand U16389 (N_16389,N_10783,N_10185);
nor U16390 (N_16390,N_11737,N_13332);
nor U16391 (N_16391,N_11601,N_12611);
xor U16392 (N_16392,N_14977,N_14793);
nand U16393 (N_16393,N_11646,N_14794);
and U16394 (N_16394,N_10388,N_14245);
nand U16395 (N_16395,N_13717,N_11106);
nand U16396 (N_16396,N_11846,N_10621);
or U16397 (N_16397,N_13328,N_13455);
and U16398 (N_16398,N_13092,N_12760);
or U16399 (N_16399,N_12537,N_10331);
and U16400 (N_16400,N_13238,N_10921);
xnor U16401 (N_16401,N_12491,N_13936);
and U16402 (N_16402,N_14800,N_14728);
and U16403 (N_16403,N_12323,N_14805);
xor U16404 (N_16404,N_10546,N_11019);
nand U16405 (N_16405,N_14063,N_11516);
and U16406 (N_16406,N_14421,N_11884);
xor U16407 (N_16407,N_14898,N_14204);
nor U16408 (N_16408,N_12179,N_11157);
or U16409 (N_16409,N_12549,N_11468);
nand U16410 (N_16410,N_11359,N_14950);
nand U16411 (N_16411,N_12726,N_11117);
and U16412 (N_16412,N_14179,N_14304);
nor U16413 (N_16413,N_11753,N_12628);
nor U16414 (N_16414,N_12100,N_12659);
or U16415 (N_16415,N_10098,N_13095);
and U16416 (N_16416,N_10221,N_12124);
nand U16417 (N_16417,N_14563,N_12015);
or U16418 (N_16418,N_10637,N_11156);
nor U16419 (N_16419,N_14935,N_11356);
and U16420 (N_16420,N_11244,N_12157);
or U16421 (N_16421,N_12098,N_10274);
or U16422 (N_16422,N_11004,N_10758);
nor U16423 (N_16423,N_10064,N_12056);
nand U16424 (N_16424,N_11401,N_13554);
nor U16425 (N_16425,N_12621,N_12693);
or U16426 (N_16426,N_13327,N_11067);
and U16427 (N_16427,N_10813,N_14581);
or U16428 (N_16428,N_11235,N_10859);
and U16429 (N_16429,N_13975,N_11772);
and U16430 (N_16430,N_13607,N_11622);
or U16431 (N_16431,N_11878,N_12281);
nor U16432 (N_16432,N_14001,N_14411);
and U16433 (N_16433,N_11204,N_11761);
nand U16434 (N_16434,N_12711,N_11913);
nand U16435 (N_16435,N_13995,N_10478);
nand U16436 (N_16436,N_10611,N_12658);
xnor U16437 (N_16437,N_10945,N_14092);
or U16438 (N_16438,N_10584,N_14378);
nor U16439 (N_16439,N_13139,N_12959);
nand U16440 (N_16440,N_10634,N_10722);
nand U16441 (N_16441,N_12741,N_10877);
or U16442 (N_16442,N_11816,N_13050);
or U16443 (N_16443,N_14863,N_14206);
and U16444 (N_16444,N_10570,N_11098);
or U16445 (N_16445,N_12561,N_13800);
nand U16446 (N_16446,N_10926,N_10786);
or U16447 (N_16447,N_10079,N_14062);
nor U16448 (N_16448,N_10419,N_13966);
and U16449 (N_16449,N_14457,N_10723);
nor U16450 (N_16450,N_12137,N_12506);
nand U16451 (N_16451,N_13352,N_13085);
nand U16452 (N_16452,N_12048,N_11830);
nand U16453 (N_16453,N_11329,N_13805);
nand U16454 (N_16454,N_13351,N_11254);
or U16455 (N_16455,N_11193,N_12183);
or U16456 (N_16456,N_12674,N_14811);
and U16457 (N_16457,N_13273,N_12284);
and U16458 (N_16458,N_14466,N_11941);
nor U16459 (N_16459,N_14362,N_10691);
or U16460 (N_16460,N_14531,N_10757);
nor U16461 (N_16461,N_13104,N_13756);
nand U16462 (N_16462,N_11509,N_13996);
and U16463 (N_16463,N_11283,N_12806);
or U16464 (N_16464,N_11310,N_13852);
or U16465 (N_16465,N_10252,N_13662);
and U16466 (N_16466,N_13599,N_14401);
nand U16467 (N_16467,N_13828,N_11849);
or U16468 (N_16468,N_14833,N_11541);
nor U16469 (N_16469,N_14379,N_13367);
nor U16470 (N_16470,N_12792,N_12198);
or U16471 (N_16471,N_14271,N_11428);
nand U16472 (N_16472,N_10942,N_12065);
nand U16473 (N_16473,N_12942,N_12212);
nand U16474 (N_16474,N_10867,N_13061);
nand U16475 (N_16475,N_14956,N_10874);
and U16476 (N_16476,N_14615,N_12564);
nor U16477 (N_16477,N_12022,N_12870);
nand U16478 (N_16478,N_11331,N_11024);
or U16479 (N_16479,N_13517,N_11184);
nor U16480 (N_16480,N_14079,N_11364);
and U16481 (N_16481,N_13526,N_10357);
nor U16482 (N_16482,N_14127,N_10054);
or U16483 (N_16483,N_11047,N_12606);
or U16484 (N_16484,N_13739,N_14319);
nor U16485 (N_16485,N_13163,N_10936);
nor U16486 (N_16486,N_12272,N_12046);
or U16487 (N_16487,N_14317,N_10422);
and U16488 (N_16488,N_12352,N_12819);
and U16489 (N_16489,N_14166,N_11466);
nor U16490 (N_16490,N_14694,N_11260);
or U16491 (N_16491,N_12949,N_10721);
and U16492 (N_16492,N_11191,N_11617);
nor U16493 (N_16493,N_10696,N_14077);
and U16494 (N_16494,N_13263,N_13322);
nand U16495 (N_16495,N_13482,N_13044);
and U16496 (N_16496,N_14865,N_13359);
nor U16497 (N_16497,N_13915,N_10147);
or U16498 (N_16498,N_12035,N_13751);
nor U16499 (N_16499,N_13910,N_13687);
nand U16500 (N_16500,N_10863,N_12368);
nand U16501 (N_16501,N_13638,N_13042);
nor U16502 (N_16502,N_10312,N_11800);
and U16503 (N_16503,N_12501,N_14692);
nand U16504 (N_16504,N_14281,N_12317);
or U16505 (N_16505,N_11645,N_10365);
or U16506 (N_16506,N_11810,N_11733);
or U16507 (N_16507,N_12877,N_14456);
nor U16508 (N_16508,N_11503,N_10800);
or U16509 (N_16509,N_14323,N_12267);
and U16510 (N_16510,N_14298,N_10988);
or U16511 (N_16511,N_14612,N_14764);
or U16512 (N_16512,N_13361,N_13162);
nor U16513 (N_16513,N_13099,N_13389);
nand U16514 (N_16514,N_14554,N_13020);
and U16515 (N_16515,N_11108,N_11650);
or U16516 (N_16516,N_14838,N_12667);
xor U16517 (N_16517,N_14678,N_12591);
nand U16518 (N_16518,N_13624,N_12731);
nor U16519 (N_16519,N_10492,N_14767);
nand U16520 (N_16520,N_13586,N_13973);
nand U16521 (N_16521,N_11295,N_12855);
or U16522 (N_16522,N_10436,N_12881);
and U16523 (N_16523,N_11796,N_11907);
nand U16524 (N_16524,N_13466,N_10167);
or U16525 (N_16525,N_11756,N_10626);
or U16526 (N_16526,N_12928,N_10055);
nand U16527 (N_16527,N_11372,N_12829);
xor U16528 (N_16528,N_13940,N_14504);
nor U16529 (N_16529,N_13798,N_11551);
or U16530 (N_16530,N_10534,N_14374);
or U16531 (N_16531,N_10451,N_11238);
and U16532 (N_16532,N_12848,N_14755);
nand U16533 (N_16533,N_13801,N_14597);
and U16534 (N_16534,N_10887,N_14433);
nor U16535 (N_16535,N_14307,N_11547);
nand U16536 (N_16536,N_13206,N_13470);
and U16537 (N_16537,N_14019,N_14578);
and U16538 (N_16538,N_13643,N_11346);
nor U16539 (N_16539,N_10960,N_10471);
nand U16540 (N_16540,N_13512,N_13533);
or U16541 (N_16541,N_12307,N_13445);
and U16542 (N_16542,N_10386,N_14930);
nand U16543 (N_16543,N_10242,N_12172);
nand U16544 (N_16544,N_13530,N_12961);
nand U16545 (N_16545,N_10339,N_10409);
and U16546 (N_16546,N_14010,N_11050);
and U16547 (N_16547,N_11160,N_11377);
or U16548 (N_16548,N_10493,N_10771);
or U16549 (N_16549,N_14689,N_11392);
and U16550 (N_16550,N_12678,N_14185);
nand U16551 (N_16551,N_10784,N_13403);
nand U16552 (N_16552,N_12602,N_11010);
or U16553 (N_16553,N_13629,N_14486);
nor U16554 (N_16554,N_14835,N_13222);
nand U16555 (N_16555,N_12968,N_14585);
nand U16556 (N_16556,N_12833,N_11363);
or U16557 (N_16557,N_10257,N_13426);
nor U16558 (N_16558,N_12945,N_10335);
nand U16559 (N_16559,N_14526,N_10555);
nand U16560 (N_16560,N_11598,N_14496);
nor U16561 (N_16561,N_13090,N_11470);
xor U16562 (N_16562,N_12728,N_12358);
and U16563 (N_16563,N_14197,N_11011);
and U16564 (N_16564,N_12631,N_14769);
nand U16565 (N_16565,N_13882,N_11369);
nand U16566 (N_16566,N_12783,N_10512);
or U16567 (N_16567,N_12925,N_10904);
xnor U16568 (N_16568,N_11210,N_12010);
nor U16569 (N_16569,N_13593,N_12224);
nand U16570 (N_16570,N_11808,N_11712);
nor U16571 (N_16571,N_14693,N_12463);
and U16572 (N_16572,N_10107,N_13929);
xnor U16573 (N_16573,N_11784,N_10508);
nand U16574 (N_16574,N_11150,N_14194);
and U16575 (N_16575,N_14081,N_10201);
and U16576 (N_16576,N_11040,N_14212);
nor U16577 (N_16577,N_11130,N_14061);
and U16578 (N_16578,N_10066,N_10218);
nor U16579 (N_16579,N_10359,N_11131);
and U16580 (N_16580,N_12861,N_14193);
and U16581 (N_16581,N_12874,N_11407);
and U16582 (N_16582,N_10984,N_12029);
and U16583 (N_16583,N_12853,N_12560);
or U16584 (N_16584,N_12434,N_10601);
nand U16585 (N_16585,N_12249,N_13884);
xnor U16586 (N_16586,N_13851,N_12080);
nand U16587 (N_16587,N_13125,N_12242);
nand U16588 (N_16588,N_11431,N_13893);
nand U16589 (N_16589,N_10489,N_10939);
and U16590 (N_16590,N_13037,N_11982);
xnor U16591 (N_16591,N_11978,N_12296);
or U16592 (N_16592,N_14674,N_11141);
and U16593 (N_16593,N_12517,N_12409);
or U16594 (N_16594,N_10692,N_10551);
nand U16595 (N_16595,N_11484,N_12559);
nand U16596 (N_16596,N_14770,N_13181);
nand U16597 (N_16597,N_12876,N_13300);
and U16598 (N_16598,N_13532,N_10727);
nand U16599 (N_16599,N_11591,N_11237);
or U16600 (N_16600,N_14709,N_13927);
or U16601 (N_16601,N_13443,N_11954);
and U16602 (N_16602,N_13651,N_12778);
and U16603 (N_16603,N_11490,N_13804);
nand U16604 (N_16604,N_10602,N_10109);
or U16605 (N_16605,N_12335,N_12381);
and U16606 (N_16606,N_14435,N_11621);
xnor U16607 (N_16607,N_14537,N_10117);
nand U16608 (N_16608,N_10078,N_10465);
and U16609 (N_16609,N_12290,N_11461);
or U16610 (N_16610,N_13523,N_14080);
and U16611 (N_16611,N_10958,N_10378);
and U16612 (N_16612,N_13857,N_12116);
or U16613 (N_16613,N_14676,N_11722);
or U16614 (N_16614,N_13360,N_12966);
or U16615 (N_16615,N_13732,N_12809);
and U16616 (N_16616,N_10160,N_12637);
and U16617 (N_16617,N_12073,N_11705);
nor U16618 (N_16618,N_11695,N_11170);
nor U16619 (N_16619,N_12395,N_11936);
and U16620 (N_16620,N_10734,N_14931);
nand U16621 (N_16621,N_11950,N_10726);
or U16622 (N_16622,N_10004,N_11990);
and U16623 (N_16623,N_10701,N_12762);
nor U16624 (N_16624,N_12610,N_13476);
and U16625 (N_16625,N_14488,N_13342);
or U16626 (N_16626,N_10544,N_13942);
nor U16627 (N_16627,N_12841,N_14571);
nor U16628 (N_16628,N_12857,N_10641);
and U16629 (N_16629,N_12751,N_10675);
and U16630 (N_16630,N_11078,N_10031);
and U16631 (N_16631,N_14894,N_10794);
nand U16632 (N_16632,N_13031,N_12750);
nand U16633 (N_16633,N_11292,N_14342);
or U16634 (N_16634,N_11730,N_13799);
xor U16635 (N_16635,N_14188,N_11439);
or U16636 (N_16636,N_12763,N_11921);
or U16637 (N_16637,N_11180,N_12516);
nand U16638 (N_16638,N_10788,N_10628);
or U16639 (N_16639,N_11636,N_13168);
nor U16640 (N_16640,N_12019,N_12894);
or U16641 (N_16641,N_13054,N_13899);
nand U16642 (N_16642,N_11626,N_14507);
nand U16643 (N_16643,N_11656,N_11284);
and U16644 (N_16644,N_10120,N_14330);
and U16645 (N_16645,N_14143,N_10961);
or U16646 (N_16646,N_12799,N_14872);
and U16647 (N_16647,N_12844,N_11063);
nand U16648 (N_16648,N_12329,N_10643);
nor U16649 (N_16649,N_10713,N_11643);
and U16650 (N_16650,N_12052,N_13189);
nor U16651 (N_16651,N_11860,N_10872);
nor U16652 (N_16652,N_10318,N_12318);
xor U16653 (N_16653,N_11353,N_14519);
xor U16654 (N_16654,N_12727,N_14510);
or U16655 (N_16655,N_13591,N_12944);
or U16656 (N_16656,N_11291,N_10216);
xor U16657 (N_16657,N_11966,N_11724);
or U16658 (N_16658,N_11315,N_13369);
nor U16659 (N_16659,N_12382,N_12510);
or U16660 (N_16660,N_14220,N_12379);
nand U16661 (N_16661,N_14734,N_13803);
xnor U16662 (N_16662,N_11975,N_14570);
nor U16663 (N_16663,N_14018,N_13219);
xor U16664 (N_16664,N_12671,N_14369);
nand U16665 (N_16665,N_12149,N_12277);
or U16666 (N_16666,N_11713,N_11311);
or U16667 (N_16667,N_14343,N_13565);
nor U16668 (N_16668,N_11074,N_14279);
and U16669 (N_16669,N_14960,N_14349);
nor U16670 (N_16670,N_10682,N_10809);
nor U16671 (N_16671,N_13166,N_10993);
nand U16672 (N_16672,N_13897,N_10215);
nor U16673 (N_16673,N_10024,N_10731);
nand U16674 (N_16674,N_13767,N_11841);
or U16675 (N_16675,N_14940,N_14328);
nor U16676 (N_16676,N_14268,N_13423);
nand U16677 (N_16677,N_14853,N_12940);
xor U16678 (N_16678,N_14682,N_14461);
xor U16679 (N_16679,N_13563,N_12102);
and U16680 (N_16680,N_10382,N_11041);
and U16681 (N_16681,N_12014,N_14595);
nor U16682 (N_16682,N_11701,N_13628);
nand U16683 (N_16683,N_11194,N_13145);
or U16684 (N_16684,N_13451,N_10353);
and U16685 (N_16685,N_13199,N_14600);
or U16686 (N_16686,N_11658,N_11620);
nor U16687 (N_16687,N_13078,N_11763);
nor U16688 (N_16688,N_10171,N_12412);
and U16689 (N_16689,N_14203,N_11684);
nor U16690 (N_16690,N_13349,N_13375);
nand U16691 (N_16691,N_11149,N_13835);
nand U16692 (N_16692,N_11602,N_14321);
or U16693 (N_16693,N_10071,N_10014);
or U16694 (N_16694,N_14740,N_13010);
and U16695 (N_16695,N_12650,N_13710);
and U16696 (N_16696,N_14446,N_12826);
and U16697 (N_16697,N_10013,N_14586);
nor U16698 (N_16698,N_12437,N_14572);
nor U16699 (N_16699,N_14260,N_14175);
nor U16700 (N_16700,N_10332,N_10181);
nor U16701 (N_16701,N_11923,N_10017);
nand U16702 (N_16702,N_10932,N_10485);
nand U16703 (N_16703,N_14119,N_14945);
nor U16704 (N_16704,N_10487,N_10803);
and U16705 (N_16705,N_12911,N_11877);
xor U16706 (N_16706,N_14086,N_14278);
or U16707 (N_16707,N_12716,N_12680);
or U16708 (N_16708,N_14723,N_11673);
nor U16709 (N_16709,N_14604,N_12964);
and U16710 (N_16710,N_12721,N_11718);
or U16711 (N_16711,N_10191,N_10244);
or U16712 (N_16712,N_12842,N_12299);
nand U16713 (N_16713,N_10081,N_11533);
nor U16714 (N_16714,N_11209,N_13696);
xor U16715 (N_16715,N_12103,N_10119);
xor U16716 (N_16716,N_10912,N_13108);
nand U16717 (N_16717,N_10406,N_13873);
nor U16718 (N_16718,N_12030,N_14085);
and U16719 (N_16719,N_12009,N_10517);
nor U16720 (N_16720,N_10899,N_11485);
nor U16721 (N_16721,N_11676,N_10323);
nor U16722 (N_16722,N_13534,N_14182);
nor U16723 (N_16723,N_14029,N_14477);
or U16724 (N_16724,N_10908,N_10876);
and U16725 (N_16725,N_13416,N_11869);
nand U16726 (N_16726,N_11303,N_14601);
nor U16727 (N_16727,N_13959,N_14171);
or U16728 (N_16728,N_13003,N_14828);
xnor U16729 (N_16729,N_13708,N_10807);
nand U16730 (N_16730,N_12185,N_11376);
or U16731 (N_16731,N_14348,N_11981);
nor U16732 (N_16732,N_13040,N_11460);
and U16733 (N_16733,N_12439,N_11104);
or U16734 (N_16734,N_13458,N_14985);
or U16735 (N_16735,N_10795,N_13572);
nor U16736 (N_16736,N_13144,N_10849);
or U16737 (N_16737,N_10352,N_10750);
xor U16738 (N_16738,N_11836,N_14980);
and U16739 (N_16739,N_10861,N_11868);
or U16740 (N_16740,N_14909,N_10010);
or U16741 (N_16741,N_10532,N_14038);
nand U16742 (N_16742,N_11564,N_10046);
xor U16743 (N_16743,N_11579,N_11826);
nand U16744 (N_16744,N_10607,N_14638);
or U16745 (N_16745,N_11958,N_11616);
or U16746 (N_16746,N_10130,N_13691);
nand U16747 (N_16747,N_10074,N_13277);
nand U16748 (N_16748,N_11648,N_11092);
and U16749 (N_16749,N_10344,N_11203);
or U16750 (N_16750,N_13540,N_10101);
and U16751 (N_16751,N_14316,N_11865);
xnor U16752 (N_16752,N_10434,N_13854);
nand U16753 (N_16753,N_14022,N_12302);
and U16754 (N_16754,N_10740,N_13642);
nand U16755 (N_16755,N_13485,N_12045);
and U16756 (N_16756,N_12798,N_14761);
or U16757 (N_16757,N_14765,N_13841);
nor U16758 (N_16758,N_12188,N_13610);
and U16759 (N_16759,N_10424,N_14012);
nor U16760 (N_16760,N_10938,N_14908);
and U16761 (N_16761,N_14989,N_11307);
and U16762 (N_16762,N_10724,N_11856);
nor U16763 (N_16763,N_10718,N_13650);
nand U16764 (N_16764,N_12003,N_10934);
or U16765 (N_16765,N_12393,N_13992);
xnor U16766 (N_16766,N_11647,N_14417);
nor U16767 (N_16767,N_12499,N_12884);
and U16768 (N_16768,N_13210,N_14974);
nand U16769 (N_16769,N_10504,N_13659);
nor U16770 (N_16770,N_14527,N_12662);
or U16771 (N_16771,N_12064,N_13507);
or U16772 (N_16772,N_14346,N_10233);
nor U16773 (N_16773,N_13392,N_14397);
nor U16774 (N_16774,N_12900,N_12669);
nand U16775 (N_16775,N_12067,N_14385);
and U16776 (N_16776,N_13136,N_10739);
and U16777 (N_16777,N_13444,N_10116);
nand U16778 (N_16778,N_13348,N_14181);
nand U16779 (N_16779,N_10368,N_13142);
nor U16780 (N_16780,N_13730,N_13270);
nor U16781 (N_16781,N_13826,N_12697);
xor U16782 (N_16782,N_13793,N_10653);
nor U16783 (N_16783,N_14311,N_14803);
and U16784 (N_16784,N_12404,N_11456);
and U16785 (N_16785,N_11008,N_11335);
nand U16786 (N_16786,N_13714,N_10497);
nand U16787 (N_16787,N_12831,N_12775);
nand U16788 (N_16788,N_12584,N_14172);
nor U16789 (N_16789,N_10488,N_14573);
nor U16790 (N_16790,N_14152,N_13260);
nor U16791 (N_16791,N_11389,N_14301);
nand U16792 (N_16792,N_13101,N_13490);
xnor U16793 (N_16793,N_14447,N_14351);
nand U16794 (N_16794,N_10077,N_12362);
nand U16795 (N_16795,N_14396,N_13492);
or U16796 (N_16796,N_14544,N_14529);
nand U16797 (N_16797,N_14308,N_14444);
and U16798 (N_16798,N_12531,N_12148);
or U16799 (N_16799,N_13553,N_13527);
nor U16800 (N_16800,N_12567,N_10917);
or U16801 (N_16801,N_11309,N_11902);
and U16802 (N_16802,N_12923,N_14979);
nor U16803 (N_16803,N_10426,N_10618);
xnor U16804 (N_16804,N_14726,N_13438);
or U16805 (N_16805,N_10247,N_12467);
or U16806 (N_16806,N_14695,N_10687);
nand U16807 (N_16807,N_12093,N_13246);
xor U16808 (N_16808,N_10513,N_13945);
nand U16809 (N_16809,N_12790,N_10845);
and U16810 (N_16810,N_14701,N_12193);
xnor U16811 (N_16811,N_14052,N_14045);
nand U16812 (N_16812,N_10762,N_14031);
or U16813 (N_16813,N_10297,N_10222);
and U16814 (N_16814,N_10586,N_13693);
and U16815 (N_16815,N_12497,N_10062);
nand U16816 (N_16816,N_11110,N_13286);
xnor U16817 (N_16817,N_11918,N_11773);
nand U16818 (N_16818,N_12346,N_13033);
xnor U16819 (N_16819,N_10177,N_14799);
and U16820 (N_16820,N_13933,N_13864);
nor U16821 (N_16821,N_11655,N_11906);
or U16822 (N_16822,N_10688,N_14886);
nand U16823 (N_16823,N_14691,N_11634);
nor U16824 (N_16824,N_11766,N_14233);
nand U16825 (N_16825,N_10457,N_10045);
and U16826 (N_16826,N_14588,N_11057);
nand U16827 (N_16827,N_11177,N_10996);
nand U16828 (N_16828,N_14102,N_13840);
xnor U16829 (N_16829,N_13081,N_10526);
and U16830 (N_16830,N_14816,N_11457);
nand U16831 (N_16831,N_11669,N_11985);
or U16832 (N_16832,N_12356,N_10126);
and U16833 (N_16833,N_13446,N_12165);
nor U16834 (N_16834,N_12544,N_13479);
and U16835 (N_16835,N_10542,N_10841);
xor U16836 (N_16836,N_13048,N_10282);
and U16837 (N_16837,N_13961,N_10214);
nor U16838 (N_16838,N_13417,N_14297);
and U16839 (N_16839,N_12794,N_12633);
xnor U16840 (N_16840,N_12012,N_11402);
nor U16841 (N_16841,N_10238,N_12737);
or U16842 (N_16842,N_12230,N_12217);
and U16843 (N_16843,N_12685,N_11593);
and U16844 (N_16844,N_13608,N_11145);
and U16845 (N_16845,N_12916,N_14965);
or U16846 (N_16846,N_11215,N_12007);
and U16847 (N_16847,N_11385,N_13768);
and U16848 (N_16848,N_11043,N_12692);
nand U16849 (N_16849,N_13810,N_13240);
or U16850 (N_16850,N_13594,N_14427);
nor U16851 (N_16851,N_13962,N_12220);
or U16852 (N_16852,N_13697,N_12291);
and U16853 (N_16853,N_11899,N_12025);
nor U16854 (N_16854,N_13667,N_10283);
and U16855 (N_16855,N_13573,N_10697);
nor U16856 (N_16856,N_10371,N_12951);
nor U16857 (N_16857,N_10894,N_10164);
nand U16858 (N_16858,N_10292,N_14370);
and U16859 (N_16859,N_14078,N_14653);
nor U16860 (N_16860,N_10969,N_13724);
nand U16861 (N_16861,N_12883,N_11139);
xnor U16862 (N_16862,N_14246,N_13237);
xor U16863 (N_16863,N_10683,N_10341);
and U16864 (N_16864,N_12836,N_10395);
nor U16865 (N_16865,N_14873,N_10658);
xnor U16866 (N_16866,N_13316,N_12057);
nand U16867 (N_16867,N_11189,N_12522);
nand U16868 (N_16868,N_10317,N_12342);
nand U16869 (N_16869,N_10923,N_13615);
or U16870 (N_16870,N_10484,N_12340);
or U16871 (N_16871,N_13891,N_10567);
nor U16872 (N_16872,N_13185,N_14722);
and U16873 (N_16873,N_13764,N_10108);
and U16874 (N_16874,N_11171,N_10865);
or U16875 (N_16875,N_10129,N_12907);
and U16876 (N_16876,N_11568,N_10677);
nand U16877 (N_16877,N_13674,N_12210);
and U16878 (N_16878,N_14970,N_13236);
or U16879 (N_16879,N_11498,N_10096);
xnor U16880 (N_16880,N_10468,N_12494);
nor U16881 (N_16881,N_11935,N_14254);
or U16882 (N_16882,N_14277,N_11949);
or U16883 (N_16883,N_13366,N_12246);
nand U16884 (N_16884,N_11839,N_13291);
nand U16885 (N_16885,N_13274,N_10518);
and U16886 (N_16886,N_11501,N_14837);
nand U16887 (N_16887,N_11247,N_11118);
xnor U16888 (N_16888,N_10998,N_11866);
or U16889 (N_16889,N_12983,N_11571);
or U16890 (N_16890,N_11253,N_10455);
and U16891 (N_16891,N_10537,N_14310);
nor U16892 (N_16892,N_13855,N_12383);
nor U16893 (N_16893,N_11012,N_10927);
or U16894 (N_16894,N_10260,N_14823);
and U16895 (N_16895,N_13036,N_12041);
nor U16896 (N_16896,N_12448,N_12780);
and U16897 (N_16897,N_11726,N_11595);
or U16898 (N_16898,N_11489,N_14553);
or U16899 (N_16899,N_11400,N_13164);
nand U16900 (N_16900,N_10159,N_14916);
nor U16901 (N_16901,N_11138,N_12575);
xnor U16902 (N_16902,N_14332,N_14821);
nor U16903 (N_16903,N_14741,N_13241);
nand U16904 (N_16904,N_10789,N_13167);
and U16905 (N_16905,N_10043,N_13365);
nand U16906 (N_16906,N_13254,N_14627);
nor U16907 (N_16907,N_14512,N_10647);
nand U16908 (N_16908,N_14844,N_14706);
nor U16909 (N_16909,N_13999,N_12574);
nand U16910 (N_16910,N_11993,N_12303);
nor U16911 (N_16911,N_14405,N_14429);
or U16912 (N_16912,N_13165,N_10565);
or U16913 (N_16913,N_12977,N_14564);
and U16914 (N_16914,N_11519,N_13787);
or U16915 (N_16915,N_12150,N_14064);
and U16916 (N_16916,N_13460,N_13784);
and U16917 (N_16917,N_14901,N_13909);
and U16918 (N_16918,N_13748,N_11075);
nor U16919 (N_16919,N_11387,N_11775);
or U16920 (N_16920,N_10503,N_11792);
or U16921 (N_16921,N_11940,N_13958);
and U16922 (N_16922,N_11762,N_11859);
nand U16923 (N_16923,N_14961,N_11444);
and U16924 (N_16924,N_14075,N_13571);
and U16925 (N_16925,N_12199,N_10369);
nor U16926 (N_16926,N_13671,N_12609);
xnor U16927 (N_16927,N_11627,N_11874);
nand U16928 (N_16928,N_11404,N_11845);
nand U16929 (N_16929,N_12503,N_14192);
or U16930 (N_16930,N_14403,N_13737);
or U16931 (N_16931,N_12524,N_13802);
and U16932 (N_16932,N_10482,N_12934);
and U16933 (N_16933,N_14820,N_13450);
nand U16934 (N_16934,N_13372,N_11747);
nor U16935 (N_16935,N_11340,N_13522);
nor U16936 (N_16936,N_14711,N_10256);
nor U16937 (N_16937,N_13311,N_11983);
nor U16938 (N_16938,N_12095,N_10627);
and U16939 (N_16939,N_12413,N_12722);
nand U16940 (N_16940,N_14984,N_12447);
nand U16941 (N_16941,N_12660,N_13783);
nor U16942 (N_16942,N_10420,N_11384);
and U16943 (N_16943,N_11179,N_11362);
nor U16944 (N_16944,N_13738,N_12937);
and U16945 (N_16945,N_14521,N_11556);
and U16946 (N_16946,N_12184,N_12235);
nor U16947 (N_16947,N_13039,N_11625);
xor U16948 (N_16948,N_10575,N_11467);
or U16949 (N_16949,N_12475,N_11119);
and U16950 (N_16950,N_11795,N_11278);
or U16951 (N_16951,N_13285,N_14702);
nand U16952 (N_16952,N_13430,N_10106);
or U16953 (N_16953,N_10090,N_13677);
and U16954 (N_16954,N_14848,N_13688);
nand U16955 (N_16955,N_14087,N_10652);
and U16956 (N_16956,N_12405,N_10906);
nand U16957 (N_16957,N_11083,N_13837);
and U16958 (N_16958,N_14641,N_13456);
nor U16959 (N_16959,N_12897,N_10606);
nand U16960 (N_16960,N_12566,N_10397);
nor U16961 (N_16961,N_12201,N_11289);
or U16962 (N_16962,N_14895,N_14073);
nand U16963 (N_16963,N_11272,N_14473);
and U16964 (N_16964,N_14215,N_12723);
xnor U16965 (N_16965,N_11314,N_13850);
nor U16966 (N_16966,N_11032,N_13480);
nor U16967 (N_16967,N_12733,N_10245);
nand U16968 (N_16968,N_12403,N_11909);
nor U16969 (N_16969,N_14262,N_10325);
nand U16970 (N_16970,N_10327,N_10188);
nand U16971 (N_16971,N_14789,N_12343);
nor U16972 (N_16972,N_14140,N_14249);
xor U16973 (N_16973,N_11243,N_14183);
and U16974 (N_16974,N_14871,N_14520);
nand U16975 (N_16975,N_11760,N_12978);
nor U16976 (N_16976,N_11482,N_12701);
nand U16977 (N_16977,N_11132,N_11017);
or U16978 (N_16978,N_13474,N_10773);
xnor U16979 (N_16979,N_10802,N_11903);
and U16980 (N_16980,N_10698,N_10625);
nand U16981 (N_16981,N_11115,N_11914);
nor U16982 (N_16982,N_14918,N_12530);
nand U16983 (N_16983,N_12485,N_11512);
nor U16984 (N_16984,N_10730,N_10846);
nor U16985 (N_16985,N_14558,N_12768);
and U16986 (N_16986,N_14534,N_10198);
nor U16987 (N_16987,N_13972,N_14450);
or U16988 (N_16988,N_10738,N_11793);
nor U16989 (N_16989,N_13701,N_14910);
nand U16990 (N_16990,N_13585,N_12086);
or U16991 (N_16991,N_10519,N_11630);
nand U16992 (N_16992,N_12312,N_11631);
and U16993 (N_16993,N_10091,N_11828);
nor U16994 (N_16994,N_10992,N_14380);
nand U16995 (N_16995,N_13655,N_14591);
xor U16996 (N_16996,N_13066,N_12624);
and U16997 (N_16997,N_12840,N_13632);
xnor U16998 (N_16998,N_13357,N_13602);
and U16999 (N_16999,N_11552,N_10878);
nand U17000 (N_17000,N_10765,N_13211);
or U17001 (N_17001,N_13598,N_13925);
or U17002 (N_17002,N_13396,N_13281);
nor U17003 (N_17003,N_13779,N_12888);
or U17004 (N_17004,N_13511,N_11326);
and U17005 (N_17005,N_10554,N_14842);
nand U17006 (N_17006,N_13649,N_10890);
xor U17007 (N_17007,N_14744,N_10189);
and U17008 (N_17008,N_13595,N_10099);
nand U17009 (N_17009,N_13538,N_14574);
and U17010 (N_17010,N_12851,N_14207);
or U17011 (N_17011,N_10496,N_12886);
and U17012 (N_17012,N_13574,N_12365);
or U17013 (N_17013,N_13770,N_14613);
and U17014 (N_17014,N_14163,N_14008);
nand U17015 (N_17015,N_12963,N_11365);
and U17016 (N_17016,N_10348,N_13387);
nor U17017 (N_17017,N_14522,N_12534);
and U17018 (N_17018,N_10362,N_11597);
nor U17019 (N_17019,N_11557,N_14532);
nor U17020 (N_17020,N_14884,N_12862);
and U17021 (N_17021,N_13093,N_14672);
nand U17022 (N_17022,N_13866,N_13982);
nand U17023 (N_17023,N_11488,N_14265);
nand U17024 (N_17024,N_10286,N_11483);
and U17025 (N_17025,N_12364,N_12321);
or U17026 (N_17026,N_14286,N_14009);
nor U17027 (N_17027,N_10494,N_14434);
or U17028 (N_17028,N_14096,N_13127);
or U17029 (N_17029,N_12846,N_11943);
nor U17030 (N_17030,N_13734,N_13584);
and U17031 (N_17031,N_11317,N_11891);
xor U17032 (N_17032,N_12020,N_14652);
nand U17033 (N_17033,N_11604,N_14919);
or U17034 (N_17034,N_13265,N_14494);
nand U17035 (N_17035,N_12089,N_12596);
and U17036 (N_17036,N_13155,N_13698);
nor U17037 (N_17037,N_13076,N_11678);
nand U17038 (N_17038,N_12287,N_10717);
or U17039 (N_17039,N_10704,N_13338);
or U17040 (N_17040,N_12118,N_13983);
or U17041 (N_17041,N_12556,N_11129);
nand U17042 (N_17042,N_13049,N_14610);
nand U17043 (N_17043,N_11544,N_13863);
nand U17044 (N_17044,N_10997,N_13978);
nand U17045 (N_17045,N_12450,N_12952);
nor U17046 (N_17046,N_11348,N_14354);
nand U17047 (N_17047,N_13234,N_14565);
or U17048 (N_17048,N_10785,N_12456);
nand U17049 (N_17049,N_11998,N_14026);
nor U17050 (N_17050,N_12251,N_10888);
nand U17051 (N_17051,N_13440,N_13068);
nor U17052 (N_17052,N_11889,N_11937);
nor U17053 (N_17053,N_10220,N_10510);
nor U17054 (N_17054,N_11349,N_14287);
nand U17055 (N_17055,N_12481,N_12310);
nor U17056 (N_17056,N_14620,N_14781);
and U17057 (N_17057,N_13614,N_13059);
or U17058 (N_17058,N_11167,N_14579);
nor U17059 (N_17059,N_10301,N_11719);
nand U17060 (N_17060,N_14436,N_14575);
or U17061 (N_17061,N_11550,N_13504);
or U17062 (N_17062,N_12410,N_10373);
and U17063 (N_17063,N_14264,N_12039);
or U17064 (N_17064,N_10018,N_11742);
or U17065 (N_17065,N_10638,N_13197);
nor U17066 (N_17066,N_11079,N_11093);
nor U17067 (N_17067,N_10530,N_12784);
or U17068 (N_17068,N_12136,N_14669);
and U17069 (N_17069,N_11412,N_10660);
and U17070 (N_17070,N_11274,N_12253);
nand U17071 (N_17071,N_13960,N_12215);
xor U17072 (N_17072,N_10798,N_10206);
or U17073 (N_17073,N_12175,N_11432);
nor U17074 (N_17074,N_13303,N_10040);
and U17075 (N_17075,N_13518,N_11623);
nand U17076 (N_17076,N_14044,N_14484);
nand U17077 (N_17077,N_14787,N_10319);
or U17078 (N_17078,N_12736,N_10593);
and U17079 (N_17079,N_10230,N_12162);
or U17080 (N_17080,N_11984,N_13622);
nor U17081 (N_17081,N_11811,N_11390);
and U17082 (N_17082,N_12374,N_12037);
and U17083 (N_17083,N_10971,N_13364);
and U17084 (N_17084,N_10358,N_14920);
or U17085 (N_17085,N_11779,N_10461);
or U17086 (N_17086,N_12781,N_14043);
and U17087 (N_17087,N_10952,N_13221);
nand U17088 (N_17088,N_11332,N_12562);
or U17089 (N_17089,N_14727,N_14000);
and U17090 (N_17090,N_13546,N_13374);
nand U17091 (N_17091,N_12786,N_12922);
nand U17092 (N_17092,N_14129,N_13439);
and U17093 (N_17093,N_13869,N_12997);
and U17094 (N_17094,N_11835,N_14785);
and U17095 (N_17095,N_14890,N_11153);
and U17096 (N_17096,N_14269,N_12820);
xor U17097 (N_17097,N_14831,N_11542);
or U17098 (N_17098,N_12813,N_13267);
nand U17099 (N_17099,N_10193,N_13420);
or U17100 (N_17100,N_10935,N_14743);
nand U17101 (N_17101,N_13118,N_11440);
and U17102 (N_17102,N_10603,N_14146);
nor U17103 (N_17103,N_10259,N_14751);
or U17104 (N_17104,N_12406,N_12748);
nor U17105 (N_17105,N_14258,N_11691);
or U17106 (N_17106,N_14315,N_12797);
and U17107 (N_17107,N_10481,N_11227);
or U17108 (N_17108,N_14671,N_11525);
nand U17109 (N_17109,N_10840,N_12464);
nand U17110 (N_17110,N_14808,N_11758);
nand U17111 (N_17111,N_11848,N_13196);
xnor U17112 (N_17112,N_13070,N_14783);
or U17113 (N_17113,N_14223,N_14724);
nand U17114 (N_17114,N_10594,N_11586);
and U17115 (N_17115,N_13190,N_10324);
xor U17116 (N_17116,N_11861,N_13904);
and U17117 (N_17117,N_13023,N_11612);
and U17118 (N_17118,N_14635,N_12747);
nor U17119 (N_17119,N_13483,N_10781);
xor U17120 (N_17120,N_13158,N_10913);
nor U17121 (N_17121,N_12483,N_13745);
nand U17122 (N_17122,N_11666,N_12576);
or U17123 (N_17123,N_10710,N_14333);
nor U17124 (N_17124,N_10774,N_12816);
nand U17125 (N_17125,N_10498,N_12170);
nor U17126 (N_17126,N_14892,N_12252);
nand U17127 (N_17127,N_10609,N_13596);
nand U17128 (N_17128,N_11900,N_12171);
nand U17129 (N_17129,N_13292,N_13035);
nor U17130 (N_17130,N_13740,N_10144);
nand U17131 (N_17131,N_13015,N_13425);
or U17132 (N_17132,N_12938,N_12993);
xnor U17133 (N_17133,N_13728,N_10178);
or U17134 (N_17134,N_10847,N_12192);
xnor U17135 (N_17135,N_10547,N_11097);
nor U17136 (N_17136,N_13053,N_12339);
and U17137 (N_17137,N_10741,N_13339);
nand U17138 (N_17138,N_10915,N_10328);
nor U17139 (N_17139,N_10132,N_11351);
nor U17140 (N_17140,N_11077,N_13817);
nor U17141 (N_17141,N_12411,N_13957);
or U17142 (N_17142,N_13146,N_12142);
nand U17143 (N_17143,N_12772,N_12579);
or U17144 (N_17144,N_10412,N_13024);
nand U17145 (N_17145,N_14068,N_10421);
or U17146 (N_17146,N_10190,N_13253);
or U17147 (N_17147,N_12505,N_13047);
nand U17148 (N_17148,N_11434,N_12656);
and U17149 (N_17149,N_12729,N_11930);
xor U17150 (N_17150,N_11635,N_14272);
nor U17151 (N_17151,N_11113,N_11607);
nand U17152 (N_17152,N_14135,N_11495);
xnor U17153 (N_17153,N_14225,N_11168);
nand U17154 (N_17154,N_14983,N_14151);
and U17155 (N_17155,N_13587,N_11112);
nand U17156 (N_17156,N_12528,N_10427);
and U17157 (N_17157,N_14285,N_14218);
nand U17158 (N_17158,N_13679,N_14180);
nor U17159 (N_17159,N_11947,N_13288);
nand U17160 (N_17160,N_10664,N_14159);
or U17161 (N_17161,N_12583,N_14049);
nor U17162 (N_17162,N_11350,N_12371);
or U17163 (N_17163,N_13922,N_10276);
or U17164 (N_17164,N_14536,N_10694);
xor U17165 (N_17165,N_10100,N_11492);
nor U17166 (N_17166,N_13310,N_10343);
or U17167 (N_17167,N_14238,N_11806);
nor U17168 (N_17168,N_11735,N_14625);
or U17169 (N_17169,N_10550,N_13541);
and U17170 (N_17170,N_13763,N_12954);
nand U17171 (N_17171,N_13811,N_14830);
and U17172 (N_17172,N_12910,N_11500);
or U17173 (N_17173,N_13830,N_11723);
nor U17174 (N_17174,N_10112,N_12283);
nand U17175 (N_17175,N_14187,N_11963);
nor U17176 (N_17176,N_12599,N_10399);
and U17177 (N_17177,N_14657,N_12361);
nor U17178 (N_17178,N_13004,N_11823);
or U17179 (N_17179,N_14133,N_10686);
nor U17180 (N_17180,N_12400,N_13822);
xnor U17181 (N_17181,N_12675,N_13487);
nand U17182 (N_17182,N_11279,N_13071);
and U17183 (N_17183,N_14232,N_10239);
or U17184 (N_17184,N_14428,N_13917);
nand U17185 (N_17185,N_12417,N_13350);
nand U17186 (N_17186,N_12195,N_10864);
nor U17187 (N_17187,N_12595,N_14089);
or U17188 (N_17188,N_11979,N_10708);
nand U17189 (N_17189,N_13916,N_13867);
or U17190 (N_17190,N_13760,N_14222);
nand U17191 (N_17191,N_10712,N_10834);
nand U17192 (N_17192,N_14992,N_14567);
nor U17193 (N_17193,N_10027,N_11418);
nand U17194 (N_17194,N_13016,N_12681);
or U17195 (N_17195,N_14845,N_12373);
nor U17196 (N_17196,N_12128,N_11814);
nor U17197 (N_17197,N_11663,N_12987);
nor U17198 (N_17198,N_12705,N_10529);
nand U17199 (N_17199,N_14875,N_12967);
nor U17200 (N_17200,N_11330,N_10383);
nor U17201 (N_17201,N_11144,N_13712);
nor U17202 (N_17202,N_11786,N_13743);
and U17203 (N_17203,N_14190,N_10644);
nor U17204 (N_17204,N_11296,N_14352);
nand U17205 (N_17205,N_12245,N_10446);
and U17206 (N_17206,N_14419,N_11517);
nor U17207 (N_17207,N_14698,N_13499);
nor U17208 (N_17208,N_13736,N_11973);
or U17209 (N_17209,N_14696,N_14492);
or U17210 (N_17210,N_11185,N_12487);
or U17211 (N_17211,N_14084,N_12712);
and U17212 (N_17212,N_11288,N_12823);
and U17213 (N_17213,N_11360,N_12081);
or U17214 (N_17214,N_14145,N_10616);
or U17215 (N_17215,N_13761,N_12758);
and U17216 (N_17216,N_13283,N_14201);
nor U17217 (N_17217,N_11068,N_10663);
and U17218 (N_17218,N_12555,N_13218);
and U17219 (N_17219,N_12554,N_11599);
xor U17220 (N_17220,N_11425,N_14060);
nand U17221 (N_17221,N_12496,N_14112);
nand U17222 (N_17222,N_14991,N_12803);
or U17223 (N_17223,N_12655,N_14732);
and U17224 (N_17224,N_12445,N_12070);
nand U17225 (N_17225,N_13177,N_10751);
nor U17226 (N_17226,N_14587,N_14688);
nand U17227 (N_17227,N_14867,N_14091);
or U17228 (N_17228,N_11671,N_13194);
or U17229 (N_17229,N_14256,N_14500);
nand U17230 (N_17230,N_11299,N_11734);
and U17231 (N_17231,N_11480,N_11674);
nor U17232 (N_17232,N_13862,N_13892);
nor U17233 (N_17233,N_14247,N_11308);
nand U17234 (N_17234,N_10330,N_11143);
and U17235 (N_17235,N_14937,N_13885);
and U17236 (N_17236,N_10914,N_12083);
nor U17237 (N_17237,N_10402,N_13233);
nor U17238 (N_17238,N_10991,N_11073);
nor U17239 (N_17239,N_11566,N_11685);
nand U17240 (N_17240,N_14057,N_10195);
and U17241 (N_17241,N_13202,N_12905);
nand U17242 (N_17242,N_10948,N_12469);
nor U17243 (N_17243,N_11696,N_12753);
or U17244 (N_17244,N_13148,N_11659);
nand U17245 (N_17245,N_10808,N_13809);
or U17246 (N_17246,N_12058,N_12766);
and U17247 (N_17247,N_14559,N_13243);
nand U17248 (N_17248,N_11382,N_14771);
nand U17249 (N_17249,N_10340,N_11931);
and U17250 (N_17250,N_13079,N_14934);
xor U17251 (N_17251,N_14035,N_14990);
nand U17252 (N_17252,N_14154,N_13182);
or U17253 (N_17253,N_11399,N_12834);
nand U17254 (N_17254,N_14251,N_13792);
nand U17255 (N_17255,N_11980,N_11107);
nor U17256 (N_17256,N_11065,N_12087);
nand U17257 (N_17257,N_12970,N_13409);
nand U17258 (N_17258,N_13475,N_13176);
or U17259 (N_17259,N_13647,N_14677);
and U17260 (N_17260,N_12698,N_13170);
nor U17261 (N_17261,N_10334,N_10916);
or U17262 (N_17262,N_13894,N_12926);
and U17263 (N_17263,N_11924,N_12016);
nand U17264 (N_17264,N_10604,N_11487);
nor U17265 (N_17265,N_13753,N_12980);
nor U17266 (N_17266,N_14841,N_14438);
nor U17267 (N_17267,N_12455,N_10143);
nor U17268 (N_17268,N_12757,N_13007);
and U17269 (N_17269,N_10428,N_12541);
nor U17270 (N_17270,N_11968,N_14137);
nor U17271 (N_17271,N_10392,N_13017);
nor U17272 (N_17272,N_12502,N_10595);
nand U17273 (N_17273,N_14339,N_14425);
nand U17274 (N_17274,N_13568,N_10703);
or U17275 (N_17275,N_11354,N_14198);
nor U17276 (N_17276,N_14827,N_11782);
nor U17277 (N_17277,N_10156,N_11357);
and U17278 (N_17278,N_10346,N_10396);
nand U17279 (N_17279,N_12634,N_13307);
nand U17280 (N_17280,N_10118,N_14914);
or U17281 (N_17281,N_12247,N_11506);
xor U17282 (N_17282,N_10819,N_14551);
nand U17283 (N_17283,N_14959,N_10384);
xor U17284 (N_17284,N_13301,N_11042);
or U17285 (N_17285,N_13018,N_12921);
nand U17286 (N_17286,N_14219,N_11080);
nor U17287 (N_17287,N_11894,N_10303);
or U17288 (N_17288,N_13418,N_11282);
nand U17289 (N_17289,N_10437,N_10439);
and U17290 (N_17290,N_11687,N_14478);
or U17291 (N_17291,N_10057,N_13089);
nor U17292 (N_17292,N_13377,N_10342);
and U17293 (N_17293,N_13702,N_11388);
nand U17294 (N_17294,N_12488,N_10293);
xnor U17295 (N_17295,N_14350,N_13252);
or U17296 (N_17296,N_13008,N_14566);
nand U17297 (N_17297,N_13313,N_11588);
nor U17298 (N_17298,N_10094,N_11812);
and U17299 (N_17299,N_14868,N_13848);
or U17300 (N_17300,N_12202,N_13198);
or U17301 (N_17301,N_13508,N_12565);
nand U17302 (N_17302,N_12440,N_11725);
nand U17303 (N_17303,N_13452,N_13868);
nand U17304 (N_17304,N_11915,N_11070);
nand U17305 (N_17305,N_13461,N_13634);
nor U17306 (N_17306,N_14611,N_11405);
nor U17307 (N_17307,N_13086,N_14169);
or U17308 (N_17308,N_10438,N_11373);
or U17309 (N_17309,N_10423,N_10816);
and U17310 (N_17310,N_13604,N_11195);
xor U17311 (N_17311,N_13391,N_10965);
nand U17312 (N_17312,N_14975,N_13129);
or U17313 (N_17313,N_13794,N_11473);
and U17314 (N_17314,N_14235,N_12999);
nor U17315 (N_17315,N_10761,N_13149);
and U17316 (N_17316,N_13720,N_14071);
nor U17317 (N_17317,N_10310,N_13981);
nor U17318 (N_17318,N_12292,N_12351);
or U17319 (N_17319,N_10516,N_10668);
nor U17320 (N_17320,N_12593,N_14746);
and U17321 (N_17321,N_12332,N_12640);
and U17322 (N_17322,N_14862,N_13287);
nor U17323 (N_17323,N_11003,N_14516);
nor U17324 (N_17324,N_14589,N_14847);
nor U17325 (N_17325,N_11212,N_10903);
or U17326 (N_17326,N_13993,N_14763);
nor U17327 (N_17327,N_14813,N_10705);
and U17328 (N_17328,N_14460,N_11226);
nor U17329 (N_17329,N_14329,N_12538);
nor U17330 (N_17330,N_14250,N_11090);
and U17331 (N_17331,N_13991,N_11553);
and U17332 (N_17332,N_14550,N_10853);
nor U17333 (N_17333,N_14777,N_14697);
nand U17334 (N_17334,N_11173,N_11450);
or U17335 (N_17335,N_13132,N_12033);
or U17336 (N_17336,N_13625,N_12174);
xor U17337 (N_17337,N_12589,N_12208);
nand U17338 (N_17338,N_14602,N_14474);
and U17339 (N_17339,N_13944,N_10322);
nand U17340 (N_17340,N_11069,N_12122);
nor U17341 (N_17341,N_10176,N_13663);
or U17342 (N_17342,N_13903,N_11208);
and U17343 (N_17343,N_14386,N_14923);
nor U17344 (N_17344,N_13408,N_11870);
and U17345 (N_17345,N_13014,N_12091);
and U17346 (N_17346,N_11987,N_11016);
or U17347 (N_17347,N_13424,N_12484);
nor U17348 (N_17348,N_12956,N_11103);
xor U17349 (N_17349,N_10404,N_11159);
or U17350 (N_17350,N_14505,N_12824);
nand U17351 (N_17351,N_12139,N_11188);
and U17352 (N_17352,N_13537,N_10536);
nor U17353 (N_17353,N_12504,N_10736);
nand U17354 (N_17354,N_14662,N_14582);
nor U17355 (N_17355,N_10314,N_14409);
nor U17356 (N_17356,N_14069,N_11657);
nor U17357 (N_17357,N_11642,N_12802);
nor U17358 (N_17358,N_14208,N_13201);
or U17359 (N_17359,N_11447,N_11285);
and U17360 (N_17360,N_14739,N_13505);
xnor U17361 (N_17361,N_14866,N_12939);
nor U17362 (N_17362,N_12055,N_13228);
nand U17363 (N_17363,N_13200,N_14228);
nor U17364 (N_17364,N_12972,N_13847);
or U17365 (N_17365,N_10931,N_11355);
and U17366 (N_17366,N_10711,N_10452);
and U17367 (N_17367,N_14463,N_13782);
nand U17368 (N_17368,N_11783,N_11521);
and U17369 (N_17369,N_13509,N_13786);
nand U17370 (N_17370,N_11624,N_13215);
nand U17371 (N_17371,N_12568,N_14810);
and U17372 (N_17372,N_12686,N_13755);
nor U17373 (N_17373,N_10655,N_14257);
nor U17374 (N_17374,N_10026,N_12849);
and U17375 (N_17375,N_10372,N_14111);
nand U17376 (N_17376,N_14598,N_14230);
and U17377 (N_17377,N_12059,N_10982);
or U17378 (N_17378,N_13605,N_14006);
or U17379 (N_17379,N_10275,N_10985);
nor U17380 (N_17380,N_11478,N_14430);
or U17381 (N_17381,N_12026,N_12725);
or U17382 (N_17382,N_11880,N_13682);
or U17383 (N_17383,N_10631,N_11294);
or U17384 (N_17384,N_13951,N_14210);
nand U17385 (N_17385,N_12739,N_11476);
nand U17386 (N_17386,N_14874,N_14836);
or U17387 (N_17387,N_14832,N_14445);
nor U17388 (N_17388,N_13979,N_10060);
or U17389 (N_17389,N_12049,N_10321);
nand U17390 (N_17390,N_12131,N_10277);
nor U17391 (N_17391,N_13725,N_14021);
xor U17392 (N_17392,N_13187,N_11421);
nand U17393 (N_17393,N_13637,N_12815);
nor U17394 (N_17394,N_10241,N_11014);
or U17395 (N_17395,N_14907,N_14443);
nand U17396 (N_17396,N_13012,N_10367);
and U17397 (N_17397,N_10135,N_10743);
or U17398 (N_17398,N_13259,N_12615);
nand U17399 (N_17399,N_14687,N_10549);
and U17400 (N_17400,N_11020,N_14824);
nor U17401 (N_17401,N_11123,N_11086);
nand U17402 (N_17402,N_13686,N_10580);
or U17403 (N_17403,N_11448,N_11116);
nand U17404 (N_17404,N_14110,N_12074);
or U17405 (N_17405,N_12605,N_11944);
and U17406 (N_17406,N_10792,N_10149);
nor U17407 (N_17407,N_14533,N_14788);
nor U17408 (N_17408,N_14114,N_12613);
nand U17409 (N_17409,N_10051,N_10469);
nor U17410 (N_17410,N_11745,N_14312);
and U17411 (N_17411,N_10737,N_13617);
or U17412 (N_17412,N_10829,N_10978);
or U17413 (N_17413,N_13083,N_14138);
nor U17414 (N_17414,N_13613,N_10020);
or U17415 (N_17415,N_11424,N_10059);
nand U17416 (N_17416,N_12186,N_10166);
nand U17417 (N_17417,N_14483,N_10150);
or U17418 (N_17418,N_13385,N_14357);
nor U17419 (N_17419,N_11337,N_10524);
nand U17420 (N_17420,N_12863,N_14338);
nand U17421 (N_17421,N_12268,N_14776);
nor U17422 (N_17422,N_14621,N_14261);
nand U17423 (N_17423,N_10128,N_12204);
or U17424 (N_17424,N_14878,N_13880);
or U17425 (N_17425,N_10661,N_12512);
nor U17426 (N_17426,N_14731,N_10464);
nor U17427 (N_17427,N_11715,N_12330);
nor U17428 (N_17428,N_13859,N_14501);
or U17429 (N_17429,N_12962,N_13358);
or U17430 (N_17430,N_14248,N_10543);
xor U17431 (N_17431,N_12627,N_10448);
and U17432 (N_17432,N_14822,N_10179);
nand U17433 (N_17433,N_10522,N_11596);
or U17434 (N_17434,N_12261,N_11352);
nor U17435 (N_17435,N_12269,N_14314);
nor U17436 (N_17436,N_14748,N_14020);
or U17437 (N_17437,N_13153,N_11611);
nand U17438 (N_17438,N_13429,N_14670);
and U17439 (N_17439,N_11668,N_13462);
nand U17440 (N_17440,N_13778,N_12769);
nand U17441 (N_17441,N_13027,N_11543);
nand U17442 (N_17442,N_13727,N_12927);
nor U17443 (N_17443,N_11338,N_13100);
nand U17444 (N_17444,N_12535,N_11419);
nand U17445 (N_17445,N_10336,N_10194);
or U17446 (N_17446,N_13368,N_13355);
and U17447 (N_17447,N_11585,N_11999);
and U17448 (N_17448,N_12994,N_12866);
nor U17449 (N_17449,N_12038,N_11675);
nor U17450 (N_17450,N_13871,N_12415);
nor U17451 (N_17451,N_10553,N_12946);
nor U17452 (N_17452,N_12909,N_11886);
or U17453 (N_17453,N_12422,N_10793);
xor U17454 (N_17454,N_13560,N_12005);
and U17455 (N_17455,N_12264,N_10651);
or U17456 (N_17456,N_11343,N_11749);
nand U17457 (N_17457,N_10364,N_11271);
nand U17458 (N_17458,N_13844,N_14480);
or U17459 (N_17459,N_13547,N_11076);
nand U17460 (N_17460,N_13789,N_13223);
nor U17461 (N_17461,N_13172,N_14717);
nor U17462 (N_17462,N_12482,N_12305);
nand U17463 (N_17463,N_13861,N_13214);
and U17464 (N_17464,N_10288,N_12331);
nand U17465 (N_17465,N_13601,N_13400);
nand U17466 (N_17466,N_12653,N_14407);
nand U17467 (N_17467,N_13043,N_11518);
nor U17468 (N_17468,N_11190,N_12695);
nand U17469 (N_17469,N_11005,N_13834);
and U17470 (N_17470,N_13497,N_12454);
and U17471 (N_17471,N_11528,N_11064);
nor U17472 (N_17472,N_13549,N_12424);
nor U17473 (N_17473,N_12818,N_10110);
nand U17474 (N_17474,N_12941,N_14948);
and U17475 (N_17475,N_10401,N_10645);
or U17476 (N_17476,N_10749,N_11888);
nand U17477 (N_17477,N_10204,N_12814);
nor U17478 (N_17478,N_12663,N_13103);
or U17479 (N_17479,N_13064,N_14393);
nor U17480 (N_17480,N_14568,N_10044);
and U17481 (N_17481,N_13636,N_11320);
or U17482 (N_17482,N_12553,N_10559);
and U17483 (N_17483,N_12981,N_11262);
nand U17484 (N_17484,N_11677,N_13242);
and U17485 (N_17485,N_14418,N_13113);
or U17486 (N_17486,N_14191,N_12986);
nand U17487 (N_17487,N_14454,N_12664);
nand U17488 (N_17488,N_11660,N_10995);
xnor U17489 (N_17489,N_11649,N_12630);
nor U17490 (N_17490,N_13114,N_14416);
and U17491 (N_17491,N_12608,N_10941);
or U17492 (N_17492,N_11414,N_14655);
xnor U17493 (N_17493,N_11477,N_12280);
nor U17494 (N_17494,N_12587,N_11853);
nand U17495 (N_17495,N_10515,N_10715);
nor U17496 (N_17496,N_10862,N_13860);
or U17497 (N_17497,N_14766,N_10500);
xor U17498 (N_17498,N_12336,N_14993);
or U17499 (N_17499,N_10832,N_14263);
or U17500 (N_17500,N_14724,N_14737);
or U17501 (N_17501,N_10487,N_11784);
nand U17502 (N_17502,N_12930,N_10324);
nand U17503 (N_17503,N_14197,N_10739);
and U17504 (N_17504,N_13573,N_12919);
nor U17505 (N_17505,N_12828,N_11232);
and U17506 (N_17506,N_11969,N_11877);
nor U17507 (N_17507,N_12058,N_13152);
and U17508 (N_17508,N_14718,N_11356);
nor U17509 (N_17509,N_11094,N_10636);
and U17510 (N_17510,N_10697,N_11617);
or U17511 (N_17511,N_14496,N_10506);
and U17512 (N_17512,N_10730,N_14775);
nand U17513 (N_17513,N_12114,N_10391);
and U17514 (N_17514,N_11344,N_12067);
xnor U17515 (N_17515,N_14529,N_14628);
or U17516 (N_17516,N_13853,N_14951);
xnor U17517 (N_17517,N_10404,N_10203);
or U17518 (N_17518,N_12328,N_14910);
or U17519 (N_17519,N_14496,N_12178);
nor U17520 (N_17520,N_12543,N_10790);
nor U17521 (N_17521,N_12756,N_12774);
xnor U17522 (N_17522,N_11458,N_10440);
and U17523 (N_17523,N_10343,N_10744);
nor U17524 (N_17524,N_14261,N_12403);
nor U17525 (N_17525,N_11632,N_11566);
xnor U17526 (N_17526,N_13865,N_13204);
nor U17527 (N_17527,N_14345,N_10867);
nor U17528 (N_17528,N_12719,N_14747);
nor U17529 (N_17529,N_13352,N_12808);
and U17530 (N_17530,N_14554,N_10479);
xnor U17531 (N_17531,N_12309,N_10797);
xnor U17532 (N_17532,N_12533,N_11722);
nor U17533 (N_17533,N_14782,N_12646);
nor U17534 (N_17534,N_11427,N_14909);
or U17535 (N_17535,N_12146,N_11354);
nand U17536 (N_17536,N_11643,N_11540);
nor U17537 (N_17537,N_11616,N_13239);
xnor U17538 (N_17538,N_10430,N_10300);
or U17539 (N_17539,N_12969,N_11836);
nand U17540 (N_17540,N_10372,N_11367);
nand U17541 (N_17541,N_11132,N_10312);
or U17542 (N_17542,N_14985,N_11472);
xnor U17543 (N_17543,N_13605,N_11672);
or U17544 (N_17544,N_12098,N_13349);
nand U17545 (N_17545,N_12733,N_10689);
or U17546 (N_17546,N_10260,N_10635);
nand U17547 (N_17547,N_12757,N_12991);
nand U17548 (N_17548,N_12622,N_12539);
xnor U17549 (N_17549,N_12614,N_12807);
nor U17550 (N_17550,N_13648,N_12285);
and U17551 (N_17551,N_13518,N_10808);
or U17552 (N_17552,N_10651,N_11383);
or U17553 (N_17553,N_12008,N_10068);
nand U17554 (N_17554,N_11308,N_13178);
and U17555 (N_17555,N_12879,N_11015);
nor U17556 (N_17556,N_13676,N_14785);
or U17557 (N_17557,N_13562,N_12751);
and U17558 (N_17558,N_14725,N_10445);
nor U17559 (N_17559,N_11074,N_11637);
nor U17560 (N_17560,N_14791,N_10509);
nand U17561 (N_17561,N_10309,N_10260);
nor U17562 (N_17562,N_10228,N_10394);
xnor U17563 (N_17563,N_14015,N_12773);
nor U17564 (N_17564,N_14660,N_12519);
nor U17565 (N_17565,N_14502,N_10743);
or U17566 (N_17566,N_12184,N_14487);
or U17567 (N_17567,N_10056,N_11328);
or U17568 (N_17568,N_12137,N_14171);
and U17569 (N_17569,N_10241,N_13265);
nand U17570 (N_17570,N_10477,N_13682);
nor U17571 (N_17571,N_14179,N_13511);
and U17572 (N_17572,N_14345,N_11759);
or U17573 (N_17573,N_13129,N_14965);
and U17574 (N_17574,N_12535,N_11639);
and U17575 (N_17575,N_13841,N_10200);
nand U17576 (N_17576,N_14797,N_12558);
nor U17577 (N_17577,N_12694,N_12660);
nand U17578 (N_17578,N_14753,N_14462);
and U17579 (N_17579,N_11185,N_13540);
and U17580 (N_17580,N_11282,N_12643);
and U17581 (N_17581,N_10253,N_12103);
nand U17582 (N_17582,N_14077,N_13719);
xnor U17583 (N_17583,N_10717,N_14615);
xor U17584 (N_17584,N_14866,N_13303);
and U17585 (N_17585,N_11383,N_12348);
nor U17586 (N_17586,N_12233,N_14982);
nor U17587 (N_17587,N_10476,N_12667);
nand U17588 (N_17588,N_10890,N_11684);
xor U17589 (N_17589,N_12170,N_10150);
or U17590 (N_17590,N_11976,N_11545);
xnor U17591 (N_17591,N_10865,N_10729);
nand U17592 (N_17592,N_14502,N_10885);
or U17593 (N_17593,N_12808,N_14178);
nand U17594 (N_17594,N_11650,N_12393);
nor U17595 (N_17595,N_14378,N_12108);
xor U17596 (N_17596,N_11578,N_11162);
nand U17597 (N_17597,N_12517,N_10900);
nand U17598 (N_17598,N_10508,N_13756);
nand U17599 (N_17599,N_10699,N_12988);
xor U17600 (N_17600,N_13504,N_13978);
xor U17601 (N_17601,N_10190,N_11739);
nor U17602 (N_17602,N_14571,N_14128);
nor U17603 (N_17603,N_12942,N_10296);
and U17604 (N_17604,N_10156,N_11299);
or U17605 (N_17605,N_12762,N_11427);
nor U17606 (N_17606,N_10003,N_10474);
and U17607 (N_17607,N_10096,N_11979);
and U17608 (N_17608,N_14316,N_10634);
and U17609 (N_17609,N_12450,N_11904);
nand U17610 (N_17610,N_13402,N_12181);
nor U17611 (N_17611,N_11166,N_14621);
or U17612 (N_17612,N_14780,N_13531);
xnor U17613 (N_17613,N_13188,N_11682);
or U17614 (N_17614,N_12032,N_13504);
nor U17615 (N_17615,N_11955,N_12223);
nand U17616 (N_17616,N_14676,N_10258);
nor U17617 (N_17617,N_14564,N_12255);
and U17618 (N_17618,N_10589,N_11767);
nor U17619 (N_17619,N_14523,N_14676);
and U17620 (N_17620,N_13196,N_11493);
xnor U17621 (N_17621,N_13459,N_14144);
or U17622 (N_17622,N_13075,N_12614);
and U17623 (N_17623,N_14736,N_12752);
nor U17624 (N_17624,N_14495,N_14525);
or U17625 (N_17625,N_10605,N_14913);
and U17626 (N_17626,N_13516,N_10085);
and U17627 (N_17627,N_14358,N_10573);
and U17628 (N_17628,N_10800,N_14134);
xor U17629 (N_17629,N_11370,N_10852);
xnor U17630 (N_17630,N_11280,N_13565);
nor U17631 (N_17631,N_14762,N_13968);
and U17632 (N_17632,N_12252,N_13857);
nand U17633 (N_17633,N_13277,N_11483);
and U17634 (N_17634,N_12256,N_14447);
nor U17635 (N_17635,N_14063,N_13855);
xnor U17636 (N_17636,N_12107,N_13380);
nand U17637 (N_17637,N_10619,N_14440);
and U17638 (N_17638,N_13720,N_13284);
nor U17639 (N_17639,N_10366,N_11659);
or U17640 (N_17640,N_14213,N_14346);
or U17641 (N_17641,N_14394,N_14046);
and U17642 (N_17642,N_14702,N_12400);
and U17643 (N_17643,N_10241,N_10315);
or U17644 (N_17644,N_12229,N_13543);
nand U17645 (N_17645,N_14855,N_11730);
xor U17646 (N_17646,N_13976,N_13037);
and U17647 (N_17647,N_12663,N_12809);
nand U17648 (N_17648,N_11209,N_13769);
xnor U17649 (N_17649,N_14358,N_10950);
xnor U17650 (N_17650,N_12714,N_12494);
or U17651 (N_17651,N_13445,N_11024);
nand U17652 (N_17652,N_12504,N_14587);
nor U17653 (N_17653,N_12822,N_13010);
or U17654 (N_17654,N_10576,N_12551);
nand U17655 (N_17655,N_12798,N_13039);
or U17656 (N_17656,N_13162,N_13322);
nand U17657 (N_17657,N_11075,N_14871);
nand U17658 (N_17658,N_13022,N_10249);
nor U17659 (N_17659,N_14984,N_13332);
nand U17660 (N_17660,N_14391,N_14772);
and U17661 (N_17661,N_13556,N_11849);
and U17662 (N_17662,N_14707,N_11796);
and U17663 (N_17663,N_12764,N_14381);
xor U17664 (N_17664,N_11475,N_14168);
nand U17665 (N_17665,N_12286,N_14598);
nor U17666 (N_17666,N_13372,N_12819);
xnor U17667 (N_17667,N_11630,N_12414);
xor U17668 (N_17668,N_12546,N_14295);
or U17669 (N_17669,N_14693,N_14981);
or U17670 (N_17670,N_13887,N_13676);
nor U17671 (N_17671,N_12038,N_10779);
or U17672 (N_17672,N_12212,N_11825);
xnor U17673 (N_17673,N_13174,N_14161);
nor U17674 (N_17674,N_12372,N_10678);
and U17675 (N_17675,N_13643,N_10572);
and U17676 (N_17676,N_13532,N_14180);
and U17677 (N_17677,N_14844,N_13340);
or U17678 (N_17678,N_11716,N_12456);
or U17679 (N_17679,N_12070,N_12656);
nor U17680 (N_17680,N_10809,N_14039);
and U17681 (N_17681,N_14324,N_11859);
and U17682 (N_17682,N_14350,N_14023);
nand U17683 (N_17683,N_13657,N_11390);
and U17684 (N_17684,N_12216,N_12314);
nor U17685 (N_17685,N_14053,N_10888);
nor U17686 (N_17686,N_12399,N_12133);
and U17687 (N_17687,N_11411,N_10938);
and U17688 (N_17688,N_14210,N_14376);
nor U17689 (N_17689,N_12194,N_10759);
nor U17690 (N_17690,N_11902,N_11514);
and U17691 (N_17691,N_13327,N_13606);
nor U17692 (N_17692,N_13529,N_12661);
nor U17693 (N_17693,N_14905,N_10935);
or U17694 (N_17694,N_13896,N_13598);
or U17695 (N_17695,N_12418,N_14335);
nor U17696 (N_17696,N_10470,N_13947);
nand U17697 (N_17697,N_14341,N_13889);
nand U17698 (N_17698,N_12123,N_11635);
nor U17699 (N_17699,N_11537,N_10725);
xnor U17700 (N_17700,N_14477,N_14706);
nand U17701 (N_17701,N_11555,N_10972);
or U17702 (N_17702,N_14305,N_11719);
and U17703 (N_17703,N_12139,N_11644);
xor U17704 (N_17704,N_12052,N_13542);
nor U17705 (N_17705,N_10708,N_12441);
or U17706 (N_17706,N_14639,N_12962);
or U17707 (N_17707,N_12805,N_10541);
or U17708 (N_17708,N_14940,N_12494);
nand U17709 (N_17709,N_12943,N_12724);
nand U17710 (N_17710,N_14752,N_13982);
or U17711 (N_17711,N_12129,N_11066);
or U17712 (N_17712,N_14795,N_14534);
nor U17713 (N_17713,N_13936,N_11426);
or U17714 (N_17714,N_14855,N_12102);
nor U17715 (N_17715,N_11990,N_12617);
or U17716 (N_17716,N_12568,N_11236);
xor U17717 (N_17717,N_11192,N_12476);
xnor U17718 (N_17718,N_12800,N_12174);
or U17719 (N_17719,N_13973,N_11066);
nor U17720 (N_17720,N_11360,N_11705);
or U17721 (N_17721,N_11138,N_12545);
and U17722 (N_17722,N_12356,N_12025);
nor U17723 (N_17723,N_10071,N_13525);
xnor U17724 (N_17724,N_13632,N_11194);
and U17725 (N_17725,N_14516,N_13290);
nor U17726 (N_17726,N_14539,N_11496);
xnor U17727 (N_17727,N_12326,N_10932);
xor U17728 (N_17728,N_10356,N_11694);
and U17729 (N_17729,N_14040,N_10910);
nand U17730 (N_17730,N_10954,N_10159);
or U17731 (N_17731,N_14374,N_11805);
and U17732 (N_17732,N_12038,N_11728);
and U17733 (N_17733,N_11155,N_12265);
and U17734 (N_17734,N_10611,N_11027);
and U17735 (N_17735,N_11892,N_12267);
nand U17736 (N_17736,N_10159,N_14242);
nand U17737 (N_17737,N_12081,N_10970);
nor U17738 (N_17738,N_10345,N_12248);
and U17739 (N_17739,N_12107,N_13148);
xnor U17740 (N_17740,N_11815,N_14908);
nor U17741 (N_17741,N_11924,N_13599);
nor U17742 (N_17742,N_12812,N_14467);
or U17743 (N_17743,N_11342,N_14157);
or U17744 (N_17744,N_10440,N_13924);
nor U17745 (N_17745,N_10421,N_13757);
or U17746 (N_17746,N_10865,N_10443);
or U17747 (N_17747,N_11766,N_12814);
and U17748 (N_17748,N_13993,N_12895);
nand U17749 (N_17749,N_10006,N_12095);
and U17750 (N_17750,N_13757,N_10217);
nand U17751 (N_17751,N_11004,N_13531);
nand U17752 (N_17752,N_10769,N_11392);
nor U17753 (N_17753,N_11408,N_11691);
nand U17754 (N_17754,N_12304,N_11027);
or U17755 (N_17755,N_10021,N_11981);
xnor U17756 (N_17756,N_12484,N_11857);
nor U17757 (N_17757,N_13520,N_13020);
nor U17758 (N_17758,N_12329,N_12448);
or U17759 (N_17759,N_10741,N_11058);
or U17760 (N_17760,N_11894,N_11352);
nor U17761 (N_17761,N_10402,N_12558);
or U17762 (N_17762,N_11853,N_14327);
nand U17763 (N_17763,N_13263,N_12931);
nand U17764 (N_17764,N_11880,N_13233);
or U17765 (N_17765,N_13738,N_14712);
or U17766 (N_17766,N_13527,N_11508);
nor U17767 (N_17767,N_14228,N_13175);
nand U17768 (N_17768,N_12859,N_14299);
and U17769 (N_17769,N_14051,N_14735);
and U17770 (N_17770,N_13671,N_14227);
or U17771 (N_17771,N_11227,N_11689);
xor U17772 (N_17772,N_14333,N_10165);
nor U17773 (N_17773,N_11227,N_13240);
xnor U17774 (N_17774,N_10340,N_11287);
xor U17775 (N_17775,N_13207,N_10232);
and U17776 (N_17776,N_12845,N_10419);
xor U17777 (N_17777,N_11895,N_11659);
and U17778 (N_17778,N_12482,N_10554);
or U17779 (N_17779,N_12110,N_12862);
nor U17780 (N_17780,N_10395,N_12807);
and U17781 (N_17781,N_13452,N_14376);
and U17782 (N_17782,N_11312,N_13854);
or U17783 (N_17783,N_10799,N_10267);
or U17784 (N_17784,N_13336,N_12395);
or U17785 (N_17785,N_12001,N_12595);
nor U17786 (N_17786,N_10602,N_11328);
and U17787 (N_17787,N_12995,N_14676);
or U17788 (N_17788,N_12652,N_14403);
nor U17789 (N_17789,N_10807,N_10848);
and U17790 (N_17790,N_10249,N_14043);
nand U17791 (N_17791,N_12387,N_11856);
and U17792 (N_17792,N_14182,N_12748);
nor U17793 (N_17793,N_11849,N_13398);
or U17794 (N_17794,N_10151,N_12425);
xnor U17795 (N_17795,N_14931,N_12880);
nor U17796 (N_17796,N_11454,N_10382);
and U17797 (N_17797,N_10622,N_12876);
or U17798 (N_17798,N_12534,N_12991);
or U17799 (N_17799,N_11233,N_10396);
nor U17800 (N_17800,N_13390,N_11530);
nor U17801 (N_17801,N_12608,N_12719);
or U17802 (N_17802,N_13682,N_13934);
nor U17803 (N_17803,N_10563,N_10304);
or U17804 (N_17804,N_11380,N_12809);
xnor U17805 (N_17805,N_12935,N_11587);
and U17806 (N_17806,N_10955,N_10735);
nand U17807 (N_17807,N_11435,N_11237);
nor U17808 (N_17808,N_13618,N_13225);
nand U17809 (N_17809,N_14340,N_11468);
xnor U17810 (N_17810,N_12947,N_11974);
nor U17811 (N_17811,N_13104,N_10404);
nor U17812 (N_17812,N_14087,N_13780);
nor U17813 (N_17813,N_14984,N_10703);
nor U17814 (N_17814,N_13558,N_10503);
or U17815 (N_17815,N_13168,N_12215);
nand U17816 (N_17816,N_13679,N_14142);
and U17817 (N_17817,N_11666,N_12789);
and U17818 (N_17818,N_10082,N_10951);
and U17819 (N_17819,N_14662,N_13232);
nor U17820 (N_17820,N_11939,N_14057);
nand U17821 (N_17821,N_13748,N_14728);
or U17822 (N_17822,N_11420,N_10979);
or U17823 (N_17823,N_11043,N_12724);
nand U17824 (N_17824,N_11249,N_14620);
and U17825 (N_17825,N_11930,N_14190);
nor U17826 (N_17826,N_12042,N_11842);
and U17827 (N_17827,N_11690,N_14775);
nand U17828 (N_17828,N_14375,N_12307);
xnor U17829 (N_17829,N_12059,N_14358);
xor U17830 (N_17830,N_13858,N_10893);
or U17831 (N_17831,N_14552,N_10271);
nand U17832 (N_17832,N_10082,N_11780);
nor U17833 (N_17833,N_12124,N_11868);
or U17834 (N_17834,N_10500,N_12868);
nor U17835 (N_17835,N_11483,N_14921);
and U17836 (N_17836,N_11213,N_13424);
or U17837 (N_17837,N_13537,N_14311);
nor U17838 (N_17838,N_14969,N_12210);
xor U17839 (N_17839,N_13453,N_11276);
and U17840 (N_17840,N_10023,N_12323);
and U17841 (N_17841,N_10584,N_12489);
nand U17842 (N_17842,N_12047,N_11109);
xor U17843 (N_17843,N_12807,N_11794);
nand U17844 (N_17844,N_13043,N_12178);
nor U17845 (N_17845,N_13649,N_10985);
nand U17846 (N_17846,N_14614,N_12612);
nand U17847 (N_17847,N_12012,N_10859);
or U17848 (N_17848,N_14157,N_10103);
nand U17849 (N_17849,N_10932,N_12001);
or U17850 (N_17850,N_13377,N_14522);
nor U17851 (N_17851,N_10880,N_13549);
nand U17852 (N_17852,N_14228,N_12716);
and U17853 (N_17853,N_13967,N_14200);
nand U17854 (N_17854,N_11240,N_13010);
nor U17855 (N_17855,N_14208,N_14427);
and U17856 (N_17856,N_14918,N_13693);
and U17857 (N_17857,N_12690,N_10408);
nor U17858 (N_17858,N_12660,N_14971);
or U17859 (N_17859,N_11656,N_14860);
and U17860 (N_17860,N_14643,N_13062);
nand U17861 (N_17861,N_12919,N_11281);
and U17862 (N_17862,N_13448,N_13300);
or U17863 (N_17863,N_12859,N_11163);
or U17864 (N_17864,N_12875,N_10027);
and U17865 (N_17865,N_11463,N_14792);
xnor U17866 (N_17866,N_11037,N_12553);
and U17867 (N_17867,N_13715,N_13259);
nand U17868 (N_17868,N_10304,N_11783);
and U17869 (N_17869,N_14353,N_14971);
nand U17870 (N_17870,N_14868,N_14110);
and U17871 (N_17871,N_13421,N_12056);
nor U17872 (N_17872,N_13313,N_13175);
or U17873 (N_17873,N_11748,N_14814);
or U17874 (N_17874,N_13398,N_10487);
nand U17875 (N_17875,N_14004,N_14717);
and U17876 (N_17876,N_13006,N_11079);
xor U17877 (N_17877,N_11540,N_12046);
nand U17878 (N_17878,N_11715,N_13183);
xor U17879 (N_17879,N_14751,N_12743);
or U17880 (N_17880,N_14073,N_11329);
nor U17881 (N_17881,N_14460,N_11921);
or U17882 (N_17882,N_11015,N_12305);
and U17883 (N_17883,N_10863,N_13673);
or U17884 (N_17884,N_10691,N_11872);
nand U17885 (N_17885,N_13331,N_14740);
nor U17886 (N_17886,N_11525,N_12699);
nand U17887 (N_17887,N_13902,N_11487);
or U17888 (N_17888,N_14519,N_12356);
xor U17889 (N_17889,N_12359,N_14614);
nand U17890 (N_17890,N_14660,N_11013);
xnor U17891 (N_17891,N_11239,N_14496);
and U17892 (N_17892,N_12718,N_13271);
nor U17893 (N_17893,N_12545,N_10786);
and U17894 (N_17894,N_10232,N_12129);
nor U17895 (N_17895,N_13561,N_13027);
nor U17896 (N_17896,N_11040,N_10422);
nor U17897 (N_17897,N_14157,N_14423);
or U17898 (N_17898,N_13855,N_14409);
nor U17899 (N_17899,N_10883,N_14155);
xor U17900 (N_17900,N_14752,N_13966);
xor U17901 (N_17901,N_12175,N_13250);
and U17902 (N_17902,N_13157,N_13515);
xnor U17903 (N_17903,N_10057,N_10609);
xnor U17904 (N_17904,N_12398,N_12357);
nor U17905 (N_17905,N_12099,N_14940);
and U17906 (N_17906,N_11308,N_14441);
and U17907 (N_17907,N_13634,N_10689);
and U17908 (N_17908,N_11604,N_12790);
and U17909 (N_17909,N_13608,N_10105);
nand U17910 (N_17910,N_13081,N_14267);
nor U17911 (N_17911,N_14742,N_11063);
or U17912 (N_17912,N_10102,N_10367);
or U17913 (N_17913,N_14850,N_14685);
nand U17914 (N_17914,N_13990,N_11956);
nand U17915 (N_17915,N_14558,N_11581);
nand U17916 (N_17916,N_14930,N_13566);
nand U17917 (N_17917,N_14993,N_10815);
nand U17918 (N_17918,N_10177,N_13242);
or U17919 (N_17919,N_11000,N_11056);
and U17920 (N_17920,N_10719,N_13055);
and U17921 (N_17921,N_10148,N_10802);
xor U17922 (N_17922,N_13029,N_13405);
nand U17923 (N_17923,N_11982,N_10072);
nor U17924 (N_17924,N_13830,N_13960);
nor U17925 (N_17925,N_13590,N_10644);
nor U17926 (N_17926,N_13874,N_14440);
nand U17927 (N_17927,N_13548,N_11878);
nor U17928 (N_17928,N_14292,N_11759);
nand U17929 (N_17929,N_11817,N_10344);
nand U17930 (N_17930,N_13325,N_12060);
or U17931 (N_17931,N_13174,N_12543);
and U17932 (N_17932,N_11647,N_10308);
and U17933 (N_17933,N_13302,N_14426);
and U17934 (N_17934,N_13473,N_10073);
or U17935 (N_17935,N_13418,N_11148);
or U17936 (N_17936,N_13020,N_14980);
or U17937 (N_17937,N_12882,N_10247);
or U17938 (N_17938,N_10422,N_11581);
and U17939 (N_17939,N_10504,N_11617);
xnor U17940 (N_17940,N_12111,N_13600);
or U17941 (N_17941,N_14477,N_10405);
nand U17942 (N_17942,N_14910,N_10045);
or U17943 (N_17943,N_14998,N_11465);
nand U17944 (N_17944,N_13799,N_14762);
and U17945 (N_17945,N_11581,N_14864);
and U17946 (N_17946,N_10403,N_11610);
or U17947 (N_17947,N_11414,N_12126);
or U17948 (N_17948,N_11946,N_14682);
xnor U17949 (N_17949,N_12305,N_13855);
nor U17950 (N_17950,N_14159,N_11735);
and U17951 (N_17951,N_14436,N_14962);
nand U17952 (N_17952,N_10129,N_10573);
nor U17953 (N_17953,N_13032,N_14223);
nor U17954 (N_17954,N_11934,N_12678);
and U17955 (N_17955,N_14972,N_14401);
nand U17956 (N_17956,N_14117,N_14414);
nand U17957 (N_17957,N_14215,N_10408);
nand U17958 (N_17958,N_13759,N_11789);
or U17959 (N_17959,N_12019,N_11709);
or U17960 (N_17960,N_10297,N_10745);
and U17961 (N_17961,N_10003,N_14528);
nor U17962 (N_17962,N_12026,N_10362);
and U17963 (N_17963,N_11995,N_12203);
nor U17964 (N_17964,N_11490,N_11859);
nand U17965 (N_17965,N_10897,N_11890);
and U17966 (N_17966,N_14500,N_11581);
nor U17967 (N_17967,N_11337,N_13511);
nor U17968 (N_17968,N_14872,N_13813);
nor U17969 (N_17969,N_11685,N_10849);
or U17970 (N_17970,N_14794,N_14004);
nor U17971 (N_17971,N_13761,N_14189);
or U17972 (N_17972,N_11943,N_10214);
and U17973 (N_17973,N_12859,N_14630);
and U17974 (N_17974,N_11380,N_10264);
or U17975 (N_17975,N_11551,N_10354);
nor U17976 (N_17976,N_12829,N_12933);
nand U17977 (N_17977,N_13194,N_10914);
or U17978 (N_17978,N_14625,N_13443);
xnor U17979 (N_17979,N_11939,N_14221);
and U17980 (N_17980,N_12271,N_12742);
and U17981 (N_17981,N_13861,N_11532);
and U17982 (N_17982,N_14162,N_12167);
or U17983 (N_17983,N_11040,N_14951);
and U17984 (N_17984,N_13105,N_11365);
xnor U17985 (N_17985,N_13611,N_13647);
xnor U17986 (N_17986,N_14971,N_11424);
or U17987 (N_17987,N_10646,N_12922);
nand U17988 (N_17988,N_13971,N_12702);
and U17989 (N_17989,N_11003,N_11016);
nor U17990 (N_17990,N_13541,N_12680);
and U17991 (N_17991,N_11566,N_13757);
nand U17992 (N_17992,N_10828,N_14476);
and U17993 (N_17993,N_13083,N_10135);
or U17994 (N_17994,N_11285,N_14263);
nor U17995 (N_17995,N_10550,N_11816);
xor U17996 (N_17996,N_14273,N_10501);
nor U17997 (N_17997,N_13343,N_13883);
and U17998 (N_17998,N_10536,N_12313);
nor U17999 (N_17999,N_11227,N_11602);
nor U18000 (N_18000,N_14961,N_13389);
nand U18001 (N_18001,N_13995,N_13258);
or U18002 (N_18002,N_11317,N_12750);
or U18003 (N_18003,N_14471,N_14201);
and U18004 (N_18004,N_12687,N_13897);
and U18005 (N_18005,N_10007,N_13453);
and U18006 (N_18006,N_10362,N_10485);
and U18007 (N_18007,N_12447,N_11986);
and U18008 (N_18008,N_10884,N_12254);
xor U18009 (N_18009,N_10681,N_12761);
nor U18010 (N_18010,N_11131,N_14844);
or U18011 (N_18011,N_12562,N_11746);
nor U18012 (N_18012,N_14365,N_13758);
nand U18013 (N_18013,N_11806,N_12031);
nand U18014 (N_18014,N_12913,N_10982);
nor U18015 (N_18015,N_13230,N_12521);
or U18016 (N_18016,N_10986,N_13402);
xor U18017 (N_18017,N_13551,N_13423);
and U18018 (N_18018,N_13031,N_11780);
or U18019 (N_18019,N_12999,N_10927);
nor U18020 (N_18020,N_14546,N_12608);
or U18021 (N_18021,N_11205,N_10825);
nor U18022 (N_18022,N_10768,N_14587);
or U18023 (N_18023,N_13928,N_11008);
nor U18024 (N_18024,N_12437,N_11737);
xor U18025 (N_18025,N_11048,N_12234);
nor U18026 (N_18026,N_12813,N_13596);
nor U18027 (N_18027,N_13167,N_14220);
and U18028 (N_18028,N_13146,N_14938);
nand U18029 (N_18029,N_11649,N_12739);
or U18030 (N_18030,N_14457,N_13545);
nor U18031 (N_18031,N_13562,N_14616);
xnor U18032 (N_18032,N_10938,N_13290);
and U18033 (N_18033,N_11627,N_11127);
nand U18034 (N_18034,N_14851,N_12607);
nand U18035 (N_18035,N_14130,N_12583);
or U18036 (N_18036,N_14477,N_10111);
nor U18037 (N_18037,N_13309,N_14154);
xor U18038 (N_18038,N_11551,N_12598);
or U18039 (N_18039,N_10832,N_12994);
nor U18040 (N_18040,N_13802,N_10491);
and U18041 (N_18041,N_13214,N_11412);
or U18042 (N_18042,N_10822,N_11090);
or U18043 (N_18043,N_10171,N_14389);
xor U18044 (N_18044,N_13852,N_10025);
and U18045 (N_18045,N_13056,N_12850);
and U18046 (N_18046,N_11788,N_10483);
or U18047 (N_18047,N_13935,N_13127);
or U18048 (N_18048,N_11360,N_10170);
nand U18049 (N_18049,N_12132,N_10992);
nand U18050 (N_18050,N_11691,N_11181);
nand U18051 (N_18051,N_14938,N_14741);
nor U18052 (N_18052,N_14759,N_12556);
nand U18053 (N_18053,N_11727,N_13607);
nand U18054 (N_18054,N_11378,N_11848);
nand U18055 (N_18055,N_11285,N_13963);
xor U18056 (N_18056,N_10894,N_10033);
or U18057 (N_18057,N_12103,N_13433);
nand U18058 (N_18058,N_10983,N_11778);
nand U18059 (N_18059,N_10115,N_10605);
and U18060 (N_18060,N_13471,N_12888);
or U18061 (N_18061,N_11976,N_10320);
and U18062 (N_18062,N_11367,N_13263);
or U18063 (N_18063,N_14985,N_13886);
or U18064 (N_18064,N_14317,N_13886);
or U18065 (N_18065,N_12889,N_14344);
nand U18066 (N_18066,N_11591,N_10520);
or U18067 (N_18067,N_11563,N_14732);
and U18068 (N_18068,N_14088,N_11351);
and U18069 (N_18069,N_11782,N_13131);
nor U18070 (N_18070,N_11891,N_14790);
xnor U18071 (N_18071,N_12055,N_10081);
and U18072 (N_18072,N_14802,N_14875);
xnor U18073 (N_18073,N_10897,N_10221);
nand U18074 (N_18074,N_11166,N_11351);
or U18075 (N_18075,N_11325,N_11381);
nor U18076 (N_18076,N_14342,N_14058);
or U18077 (N_18077,N_11785,N_11667);
or U18078 (N_18078,N_14284,N_13218);
and U18079 (N_18079,N_10237,N_10573);
nand U18080 (N_18080,N_11317,N_11693);
nand U18081 (N_18081,N_13185,N_13023);
or U18082 (N_18082,N_13223,N_13694);
or U18083 (N_18083,N_11302,N_12666);
nor U18084 (N_18084,N_13485,N_10937);
or U18085 (N_18085,N_14834,N_11466);
nor U18086 (N_18086,N_11062,N_14963);
nor U18087 (N_18087,N_12588,N_11901);
nor U18088 (N_18088,N_13294,N_10738);
and U18089 (N_18089,N_12170,N_11901);
or U18090 (N_18090,N_13503,N_13411);
xor U18091 (N_18091,N_13107,N_11496);
or U18092 (N_18092,N_11647,N_11628);
or U18093 (N_18093,N_14591,N_11117);
nand U18094 (N_18094,N_12845,N_13002);
and U18095 (N_18095,N_10668,N_13361);
nand U18096 (N_18096,N_14396,N_12514);
and U18097 (N_18097,N_11541,N_13259);
nor U18098 (N_18098,N_11114,N_12691);
nor U18099 (N_18099,N_10412,N_13998);
nor U18100 (N_18100,N_12219,N_13781);
or U18101 (N_18101,N_12744,N_11198);
and U18102 (N_18102,N_13269,N_10491);
nand U18103 (N_18103,N_14914,N_13248);
nor U18104 (N_18104,N_14803,N_10640);
xor U18105 (N_18105,N_12147,N_13951);
xor U18106 (N_18106,N_14546,N_10792);
nor U18107 (N_18107,N_10993,N_13379);
or U18108 (N_18108,N_10600,N_12190);
xor U18109 (N_18109,N_11022,N_10348);
or U18110 (N_18110,N_13257,N_12225);
xor U18111 (N_18111,N_10133,N_10733);
nand U18112 (N_18112,N_12703,N_11628);
or U18113 (N_18113,N_14935,N_10442);
xnor U18114 (N_18114,N_13286,N_12549);
and U18115 (N_18115,N_12215,N_10649);
and U18116 (N_18116,N_10996,N_11166);
nor U18117 (N_18117,N_13106,N_14198);
and U18118 (N_18118,N_13491,N_11222);
nor U18119 (N_18119,N_14138,N_14993);
and U18120 (N_18120,N_12371,N_10862);
nor U18121 (N_18121,N_12003,N_13406);
nand U18122 (N_18122,N_13969,N_14589);
and U18123 (N_18123,N_10180,N_10643);
or U18124 (N_18124,N_11922,N_10844);
and U18125 (N_18125,N_12630,N_12866);
xor U18126 (N_18126,N_11626,N_11347);
nor U18127 (N_18127,N_10657,N_11170);
nand U18128 (N_18128,N_14547,N_12738);
and U18129 (N_18129,N_10542,N_10837);
and U18130 (N_18130,N_11978,N_13336);
or U18131 (N_18131,N_10440,N_13034);
nand U18132 (N_18132,N_14919,N_14534);
nor U18133 (N_18133,N_13384,N_13764);
and U18134 (N_18134,N_12351,N_12652);
and U18135 (N_18135,N_14644,N_13772);
or U18136 (N_18136,N_14731,N_13742);
and U18137 (N_18137,N_10511,N_12685);
nand U18138 (N_18138,N_10776,N_11739);
and U18139 (N_18139,N_10884,N_13795);
or U18140 (N_18140,N_13591,N_14032);
and U18141 (N_18141,N_11306,N_13780);
nand U18142 (N_18142,N_11453,N_13694);
nor U18143 (N_18143,N_14320,N_12796);
or U18144 (N_18144,N_13164,N_13817);
and U18145 (N_18145,N_14497,N_14439);
nand U18146 (N_18146,N_10142,N_14083);
nand U18147 (N_18147,N_12417,N_14955);
xor U18148 (N_18148,N_13756,N_11966);
and U18149 (N_18149,N_13130,N_12160);
or U18150 (N_18150,N_13966,N_11578);
and U18151 (N_18151,N_13945,N_13931);
nand U18152 (N_18152,N_14559,N_10449);
nand U18153 (N_18153,N_14970,N_14684);
nor U18154 (N_18154,N_10578,N_10427);
nand U18155 (N_18155,N_14206,N_11878);
nand U18156 (N_18156,N_12956,N_10012);
nor U18157 (N_18157,N_10074,N_14102);
or U18158 (N_18158,N_10341,N_11988);
nand U18159 (N_18159,N_12564,N_10706);
nor U18160 (N_18160,N_14708,N_12229);
or U18161 (N_18161,N_10986,N_10029);
and U18162 (N_18162,N_14692,N_10203);
and U18163 (N_18163,N_12120,N_14576);
nor U18164 (N_18164,N_12123,N_10157);
and U18165 (N_18165,N_12733,N_14238);
or U18166 (N_18166,N_11301,N_14387);
and U18167 (N_18167,N_14243,N_13697);
xor U18168 (N_18168,N_11118,N_14935);
nand U18169 (N_18169,N_11908,N_13524);
or U18170 (N_18170,N_13600,N_10816);
or U18171 (N_18171,N_14343,N_10787);
nor U18172 (N_18172,N_13952,N_14057);
and U18173 (N_18173,N_14683,N_11444);
or U18174 (N_18174,N_10067,N_11541);
nand U18175 (N_18175,N_10156,N_12510);
nand U18176 (N_18176,N_13461,N_11170);
and U18177 (N_18177,N_10161,N_10804);
nand U18178 (N_18178,N_10643,N_11814);
and U18179 (N_18179,N_11999,N_10047);
nor U18180 (N_18180,N_14513,N_14340);
nand U18181 (N_18181,N_10910,N_11035);
nand U18182 (N_18182,N_11332,N_14671);
nor U18183 (N_18183,N_12082,N_14710);
xnor U18184 (N_18184,N_12437,N_12095);
or U18185 (N_18185,N_11942,N_13357);
nor U18186 (N_18186,N_14541,N_10831);
xnor U18187 (N_18187,N_12928,N_12815);
nand U18188 (N_18188,N_11987,N_13972);
nand U18189 (N_18189,N_13422,N_12686);
or U18190 (N_18190,N_14077,N_14310);
and U18191 (N_18191,N_13752,N_11260);
nor U18192 (N_18192,N_13407,N_12539);
xor U18193 (N_18193,N_13182,N_14483);
nor U18194 (N_18194,N_13092,N_10368);
nand U18195 (N_18195,N_14725,N_11342);
nor U18196 (N_18196,N_10973,N_12922);
and U18197 (N_18197,N_13489,N_11091);
or U18198 (N_18198,N_11587,N_14192);
nand U18199 (N_18199,N_13203,N_14215);
nor U18200 (N_18200,N_11657,N_10801);
xor U18201 (N_18201,N_13839,N_10888);
and U18202 (N_18202,N_13470,N_11314);
or U18203 (N_18203,N_13829,N_13168);
nor U18204 (N_18204,N_10362,N_10925);
and U18205 (N_18205,N_10746,N_11715);
and U18206 (N_18206,N_10826,N_13769);
nor U18207 (N_18207,N_11036,N_11766);
nand U18208 (N_18208,N_12515,N_14987);
and U18209 (N_18209,N_13275,N_13476);
or U18210 (N_18210,N_13789,N_10340);
and U18211 (N_18211,N_12427,N_11000);
nor U18212 (N_18212,N_12365,N_12254);
and U18213 (N_18213,N_13756,N_10832);
xor U18214 (N_18214,N_12887,N_13647);
and U18215 (N_18215,N_13121,N_13640);
nor U18216 (N_18216,N_12071,N_12887);
nand U18217 (N_18217,N_13792,N_11395);
nand U18218 (N_18218,N_14901,N_14768);
nor U18219 (N_18219,N_10202,N_12931);
nor U18220 (N_18220,N_12805,N_10653);
nor U18221 (N_18221,N_11787,N_10426);
and U18222 (N_18222,N_11454,N_13068);
nand U18223 (N_18223,N_11205,N_10340);
and U18224 (N_18224,N_12352,N_12242);
nand U18225 (N_18225,N_14190,N_10516);
or U18226 (N_18226,N_12178,N_11676);
and U18227 (N_18227,N_12806,N_11178);
nor U18228 (N_18228,N_10559,N_10810);
and U18229 (N_18229,N_11092,N_14373);
or U18230 (N_18230,N_14817,N_13802);
or U18231 (N_18231,N_13869,N_11553);
or U18232 (N_18232,N_11097,N_10078);
nand U18233 (N_18233,N_11700,N_13126);
nand U18234 (N_18234,N_10137,N_10253);
nor U18235 (N_18235,N_12311,N_11466);
xnor U18236 (N_18236,N_13412,N_11937);
xnor U18237 (N_18237,N_10624,N_14200);
nand U18238 (N_18238,N_11014,N_14769);
or U18239 (N_18239,N_10866,N_12348);
nor U18240 (N_18240,N_13171,N_13757);
and U18241 (N_18241,N_13175,N_12892);
nor U18242 (N_18242,N_12436,N_14294);
nand U18243 (N_18243,N_14212,N_14852);
and U18244 (N_18244,N_14107,N_13113);
nor U18245 (N_18245,N_11380,N_12360);
nor U18246 (N_18246,N_13120,N_12443);
and U18247 (N_18247,N_12955,N_11080);
nand U18248 (N_18248,N_14754,N_11978);
or U18249 (N_18249,N_11380,N_12128);
or U18250 (N_18250,N_12624,N_11911);
xnor U18251 (N_18251,N_11045,N_13800);
nand U18252 (N_18252,N_11486,N_10105);
or U18253 (N_18253,N_13931,N_12180);
nand U18254 (N_18254,N_13904,N_11516);
nor U18255 (N_18255,N_12199,N_12573);
nand U18256 (N_18256,N_14220,N_14040);
and U18257 (N_18257,N_11900,N_14104);
nand U18258 (N_18258,N_11903,N_11277);
or U18259 (N_18259,N_11131,N_12293);
and U18260 (N_18260,N_14880,N_13376);
or U18261 (N_18261,N_12482,N_14608);
and U18262 (N_18262,N_13487,N_10319);
and U18263 (N_18263,N_13443,N_13244);
and U18264 (N_18264,N_11966,N_12071);
xor U18265 (N_18265,N_12479,N_11352);
xor U18266 (N_18266,N_10027,N_11184);
and U18267 (N_18267,N_14376,N_12835);
or U18268 (N_18268,N_13142,N_13712);
nor U18269 (N_18269,N_14598,N_10134);
nand U18270 (N_18270,N_12873,N_12675);
or U18271 (N_18271,N_10945,N_11824);
and U18272 (N_18272,N_12366,N_14155);
xnor U18273 (N_18273,N_14638,N_14153);
nand U18274 (N_18274,N_11144,N_14737);
nand U18275 (N_18275,N_10945,N_10808);
or U18276 (N_18276,N_10011,N_13810);
nand U18277 (N_18277,N_14316,N_14752);
or U18278 (N_18278,N_11181,N_11510);
nand U18279 (N_18279,N_14179,N_11419);
nand U18280 (N_18280,N_12610,N_14767);
or U18281 (N_18281,N_13521,N_12294);
and U18282 (N_18282,N_11212,N_13078);
and U18283 (N_18283,N_12834,N_10645);
or U18284 (N_18284,N_14191,N_14601);
nand U18285 (N_18285,N_11276,N_13299);
and U18286 (N_18286,N_13727,N_10435);
or U18287 (N_18287,N_13198,N_13512);
and U18288 (N_18288,N_10432,N_14500);
or U18289 (N_18289,N_10433,N_11518);
or U18290 (N_18290,N_13779,N_12167);
or U18291 (N_18291,N_10608,N_11411);
nor U18292 (N_18292,N_13008,N_13422);
nand U18293 (N_18293,N_14230,N_11581);
and U18294 (N_18294,N_14223,N_12473);
or U18295 (N_18295,N_12056,N_14271);
or U18296 (N_18296,N_10592,N_12831);
nand U18297 (N_18297,N_10271,N_13874);
xnor U18298 (N_18298,N_13384,N_10357);
nor U18299 (N_18299,N_13769,N_14391);
nand U18300 (N_18300,N_10120,N_14082);
nor U18301 (N_18301,N_10338,N_12303);
nor U18302 (N_18302,N_10069,N_14997);
nand U18303 (N_18303,N_14387,N_12427);
nand U18304 (N_18304,N_14445,N_13184);
and U18305 (N_18305,N_10628,N_12806);
nor U18306 (N_18306,N_12055,N_11421);
nor U18307 (N_18307,N_12401,N_14664);
and U18308 (N_18308,N_11855,N_11819);
and U18309 (N_18309,N_13956,N_12382);
xor U18310 (N_18310,N_11832,N_14023);
xor U18311 (N_18311,N_12279,N_13420);
or U18312 (N_18312,N_11167,N_12081);
and U18313 (N_18313,N_10002,N_11001);
nand U18314 (N_18314,N_14661,N_13277);
and U18315 (N_18315,N_13184,N_10974);
nor U18316 (N_18316,N_14378,N_13988);
or U18317 (N_18317,N_13191,N_14018);
nor U18318 (N_18318,N_12827,N_11584);
and U18319 (N_18319,N_10934,N_13137);
nor U18320 (N_18320,N_12735,N_10808);
and U18321 (N_18321,N_12840,N_14565);
or U18322 (N_18322,N_11436,N_12402);
and U18323 (N_18323,N_14234,N_12292);
xnor U18324 (N_18324,N_13859,N_13761);
and U18325 (N_18325,N_14471,N_12093);
and U18326 (N_18326,N_10626,N_14931);
nand U18327 (N_18327,N_14268,N_11614);
nand U18328 (N_18328,N_14610,N_11453);
nand U18329 (N_18329,N_13732,N_13420);
and U18330 (N_18330,N_13583,N_10602);
nand U18331 (N_18331,N_13961,N_12520);
and U18332 (N_18332,N_13196,N_14004);
xor U18333 (N_18333,N_14557,N_12475);
nor U18334 (N_18334,N_11026,N_13834);
nor U18335 (N_18335,N_14669,N_12188);
or U18336 (N_18336,N_10369,N_12698);
or U18337 (N_18337,N_10646,N_14742);
and U18338 (N_18338,N_10809,N_11536);
nand U18339 (N_18339,N_11929,N_11899);
and U18340 (N_18340,N_13704,N_12392);
nor U18341 (N_18341,N_11572,N_10728);
or U18342 (N_18342,N_14968,N_12110);
nand U18343 (N_18343,N_13551,N_10840);
nor U18344 (N_18344,N_14078,N_13110);
xor U18345 (N_18345,N_14097,N_14066);
and U18346 (N_18346,N_13448,N_10090);
and U18347 (N_18347,N_14115,N_11667);
xor U18348 (N_18348,N_14576,N_12573);
nand U18349 (N_18349,N_13459,N_14884);
nand U18350 (N_18350,N_11998,N_11053);
xor U18351 (N_18351,N_14912,N_11743);
nand U18352 (N_18352,N_14341,N_12942);
nor U18353 (N_18353,N_12694,N_13230);
and U18354 (N_18354,N_12001,N_10465);
nand U18355 (N_18355,N_11304,N_10855);
or U18356 (N_18356,N_11410,N_14089);
and U18357 (N_18357,N_10923,N_13538);
or U18358 (N_18358,N_12776,N_13119);
nand U18359 (N_18359,N_13287,N_12341);
nand U18360 (N_18360,N_12983,N_14470);
and U18361 (N_18361,N_11624,N_14897);
nand U18362 (N_18362,N_11457,N_12535);
and U18363 (N_18363,N_10811,N_11287);
nand U18364 (N_18364,N_13157,N_14662);
nor U18365 (N_18365,N_11503,N_10558);
and U18366 (N_18366,N_13417,N_13785);
nand U18367 (N_18367,N_11972,N_10911);
and U18368 (N_18368,N_10053,N_14807);
nand U18369 (N_18369,N_10712,N_11932);
and U18370 (N_18370,N_10226,N_12585);
nand U18371 (N_18371,N_13506,N_14095);
nor U18372 (N_18372,N_13245,N_12974);
nor U18373 (N_18373,N_13924,N_11294);
nor U18374 (N_18374,N_10620,N_12508);
xor U18375 (N_18375,N_14187,N_12652);
or U18376 (N_18376,N_11731,N_14384);
nand U18377 (N_18377,N_14736,N_14727);
nand U18378 (N_18378,N_10508,N_14611);
or U18379 (N_18379,N_14659,N_12811);
nand U18380 (N_18380,N_11504,N_11851);
nor U18381 (N_18381,N_13074,N_11376);
nor U18382 (N_18382,N_12771,N_13628);
nand U18383 (N_18383,N_11762,N_12218);
and U18384 (N_18384,N_13311,N_11770);
nand U18385 (N_18385,N_13105,N_14540);
nand U18386 (N_18386,N_11270,N_12785);
and U18387 (N_18387,N_11215,N_11432);
nand U18388 (N_18388,N_13303,N_11897);
and U18389 (N_18389,N_14379,N_13726);
nor U18390 (N_18390,N_14648,N_12365);
nand U18391 (N_18391,N_13655,N_10403);
and U18392 (N_18392,N_14967,N_14471);
nand U18393 (N_18393,N_13533,N_11736);
and U18394 (N_18394,N_13586,N_12080);
nand U18395 (N_18395,N_14071,N_12070);
or U18396 (N_18396,N_12125,N_10084);
and U18397 (N_18397,N_10811,N_13928);
and U18398 (N_18398,N_11792,N_14249);
and U18399 (N_18399,N_10476,N_11189);
or U18400 (N_18400,N_12393,N_12197);
or U18401 (N_18401,N_14747,N_14697);
and U18402 (N_18402,N_12469,N_14605);
nor U18403 (N_18403,N_11899,N_14897);
nand U18404 (N_18404,N_10625,N_12144);
nand U18405 (N_18405,N_13732,N_12749);
and U18406 (N_18406,N_11262,N_14248);
and U18407 (N_18407,N_11120,N_12346);
and U18408 (N_18408,N_13495,N_11913);
xnor U18409 (N_18409,N_14024,N_14481);
and U18410 (N_18410,N_11695,N_11317);
nand U18411 (N_18411,N_10868,N_13874);
nand U18412 (N_18412,N_14417,N_11102);
nor U18413 (N_18413,N_12578,N_12516);
or U18414 (N_18414,N_11650,N_14800);
nor U18415 (N_18415,N_14308,N_10749);
or U18416 (N_18416,N_11015,N_11829);
and U18417 (N_18417,N_11718,N_14574);
or U18418 (N_18418,N_12752,N_11046);
xor U18419 (N_18419,N_11373,N_12869);
or U18420 (N_18420,N_11577,N_10745);
nand U18421 (N_18421,N_10457,N_11923);
xnor U18422 (N_18422,N_13022,N_14784);
and U18423 (N_18423,N_10440,N_10986);
and U18424 (N_18424,N_13168,N_12297);
nand U18425 (N_18425,N_13254,N_10410);
and U18426 (N_18426,N_13749,N_13807);
nand U18427 (N_18427,N_11305,N_14490);
nor U18428 (N_18428,N_14887,N_12474);
nor U18429 (N_18429,N_13424,N_11095);
and U18430 (N_18430,N_14881,N_13542);
nor U18431 (N_18431,N_12596,N_13646);
nor U18432 (N_18432,N_13946,N_13318);
nand U18433 (N_18433,N_10328,N_12165);
or U18434 (N_18434,N_14200,N_14915);
or U18435 (N_18435,N_11037,N_13060);
nand U18436 (N_18436,N_14611,N_12668);
nand U18437 (N_18437,N_13725,N_11173);
nor U18438 (N_18438,N_12550,N_14830);
or U18439 (N_18439,N_10819,N_14700);
or U18440 (N_18440,N_10800,N_12509);
or U18441 (N_18441,N_12805,N_12865);
or U18442 (N_18442,N_14027,N_13707);
or U18443 (N_18443,N_12143,N_14072);
nand U18444 (N_18444,N_14433,N_12383);
and U18445 (N_18445,N_10338,N_14993);
nand U18446 (N_18446,N_11090,N_11600);
nor U18447 (N_18447,N_11306,N_10188);
nor U18448 (N_18448,N_11151,N_11730);
nand U18449 (N_18449,N_13668,N_10121);
nand U18450 (N_18450,N_13997,N_11060);
and U18451 (N_18451,N_13206,N_13545);
xnor U18452 (N_18452,N_14290,N_12938);
nand U18453 (N_18453,N_14748,N_13797);
and U18454 (N_18454,N_12828,N_13189);
or U18455 (N_18455,N_13179,N_10570);
nand U18456 (N_18456,N_11293,N_11955);
nor U18457 (N_18457,N_13484,N_14896);
nand U18458 (N_18458,N_12101,N_10283);
or U18459 (N_18459,N_10349,N_13501);
nand U18460 (N_18460,N_14856,N_14063);
or U18461 (N_18461,N_13605,N_10987);
nand U18462 (N_18462,N_13255,N_13097);
and U18463 (N_18463,N_14345,N_14462);
or U18464 (N_18464,N_14880,N_11399);
and U18465 (N_18465,N_11176,N_13955);
nand U18466 (N_18466,N_11707,N_10347);
nor U18467 (N_18467,N_10889,N_11046);
or U18468 (N_18468,N_11553,N_14293);
xor U18469 (N_18469,N_10660,N_10225);
or U18470 (N_18470,N_10390,N_11158);
nor U18471 (N_18471,N_11430,N_11173);
or U18472 (N_18472,N_12971,N_10667);
nor U18473 (N_18473,N_10795,N_14988);
nor U18474 (N_18474,N_12216,N_11223);
and U18475 (N_18475,N_13711,N_14149);
nor U18476 (N_18476,N_11904,N_14760);
xor U18477 (N_18477,N_12156,N_11890);
xor U18478 (N_18478,N_10603,N_12668);
and U18479 (N_18479,N_10668,N_14837);
nor U18480 (N_18480,N_10865,N_13419);
nor U18481 (N_18481,N_11552,N_10936);
nor U18482 (N_18482,N_12816,N_11053);
or U18483 (N_18483,N_12360,N_13521);
or U18484 (N_18484,N_12108,N_11087);
or U18485 (N_18485,N_12855,N_13233);
nor U18486 (N_18486,N_10030,N_13977);
nor U18487 (N_18487,N_14406,N_13319);
nand U18488 (N_18488,N_10991,N_11030);
or U18489 (N_18489,N_10009,N_11355);
nand U18490 (N_18490,N_14985,N_13774);
nand U18491 (N_18491,N_14427,N_14876);
or U18492 (N_18492,N_11433,N_11255);
or U18493 (N_18493,N_14297,N_10826);
and U18494 (N_18494,N_13511,N_13392);
or U18495 (N_18495,N_14564,N_13277);
or U18496 (N_18496,N_13595,N_10525);
nor U18497 (N_18497,N_12630,N_14527);
nand U18498 (N_18498,N_12130,N_13593);
xor U18499 (N_18499,N_13695,N_12744);
nand U18500 (N_18500,N_13065,N_12509);
or U18501 (N_18501,N_13084,N_12139);
or U18502 (N_18502,N_11496,N_12449);
or U18503 (N_18503,N_13443,N_13178);
nand U18504 (N_18504,N_10264,N_13777);
and U18505 (N_18505,N_12451,N_10817);
nor U18506 (N_18506,N_12242,N_10695);
nor U18507 (N_18507,N_11327,N_13640);
or U18508 (N_18508,N_11851,N_12760);
nor U18509 (N_18509,N_11064,N_13894);
nor U18510 (N_18510,N_10642,N_13680);
and U18511 (N_18511,N_12728,N_11511);
nand U18512 (N_18512,N_13993,N_11621);
and U18513 (N_18513,N_13327,N_11057);
or U18514 (N_18514,N_10331,N_12804);
or U18515 (N_18515,N_11848,N_14193);
or U18516 (N_18516,N_11860,N_11429);
xnor U18517 (N_18517,N_11442,N_12745);
or U18518 (N_18518,N_11120,N_12046);
or U18519 (N_18519,N_11640,N_11389);
and U18520 (N_18520,N_13859,N_12223);
or U18521 (N_18521,N_14028,N_14435);
xnor U18522 (N_18522,N_13234,N_13485);
xnor U18523 (N_18523,N_10832,N_12049);
nand U18524 (N_18524,N_10565,N_12598);
nor U18525 (N_18525,N_10700,N_14446);
nor U18526 (N_18526,N_14374,N_14065);
nand U18527 (N_18527,N_10772,N_12036);
nand U18528 (N_18528,N_13882,N_13634);
nor U18529 (N_18529,N_14753,N_13403);
nor U18530 (N_18530,N_12414,N_13192);
nor U18531 (N_18531,N_11232,N_10004);
or U18532 (N_18532,N_11789,N_13098);
nor U18533 (N_18533,N_13424,N_10657);
or U18534 (N_18534,N_11214,N_11654);
xor U18535 (N_18535,N_13151,N_12695);
nand U18536 (N_18536,N_10258,N_12815);
or U18537 (N_18537,N_10905,N_14671);
or U18538 (N_18538,N_10044,N_14045);
and U18539 (N_18539,N_14568,N_13629);
xor U18540 (N_18540,N_10649,N_14271);
nand U18541 (N_18541,N_13440,N_13722);
nor U18542 (N_18542,N_14140,N_12558);
nand U18543 (N_18543,N_13659,N_13518);
xnor U18544 (N_18544,N_13431,N_10188);
or U18545 (N_18545,N_14325,N_12736);
nand U18546 (N_18546,N_14931,N_14529);
nand U18547 (N_18547,N_13750,N_14465);
nand U18548 (N_18548,N_12969,N_14729);
nand U18549 (N_18549,N_12487,N_12630);
and U18550 (N_18550,N_11680,N_11836);
and U18551 (N_18551,N_14728,N_13523);
and U18552 (N_18552,N_13886,N_12158);
or U18553 (N_18553,N_13159,N_11251);
and U18554 (N_18554,N_10558,N_10339);
nand U18555 (N_18555,N_10921,N_10204);
and U18556 (N_18556,N_12529,N_11438);
or U18557 (N_18557,N_10150,N_12250);
or U18558 (N_18558,N_11390,N_12983);
or U18559 (N_18559,N_14695,N_10922);
and U18560 (N_18560,N_11852,N_13567);
nand U18561 (N_18561,N_11645,N_12093);
or U18562 (N_18562,N_12860,N_12027);
or U18563 (N_18563,N_14425,N_11861);
and U18564 (N_18564,N_11611,N_10119);
nor U18565 (N_18565,N_11522,N_13316);
nor U18566 (N_18566,N_12499,N_10639);
or U18567 (N_18567,N_10051,N_14905);
and U18568 (N_18568,N_12145,N_12361);
xor U18569 (N_18569,N_12487,N_10332);
nand U18570 (N_18570,N_11203,N_12414);
and U18571 (N_18571,N_14850,N_13487);
nor U18572 (N_18572,N_13323,N_13215);
nand U18573 (N_18573,N_11617,N_11319);
or U18574 (N_18574,N_11532,N_10474);
nand U18575 (N_18575,N_13050,N_12567);
nor U18576 (N_18576,N_12683,N_13945);
nor U18577 (N_18577,N_11174,N_14423);
and U18578 (N_18578,N_13761,N_13281);
xor U18579 (N_18579,N_13219,N_14218);
and U18580 (N_18580,N_11422,N_11272);
nor U18581 (N_18581,N_14137,N_12655);
nor U18582 (N_18582,N_12443,N_12755);
or U18583 (N_18583,N_10962,N_13691);
nand U18584 (N_18584,N_13423,N_13641);
or U18585 (N_18585,N_11810,N_10073);
or U18586 (N_18586,N_13480,N_11244);
and U18587 (N_18587,N_11595,N_11169);
xnor U18588 (N_18588,N_11822,N_10734);
nand U18589 (N_18589,N_10297,N_12355);
and U18590 (N_18590,N_12599,N_13270);
or U18591 (N_18591,N_14982,N_14896);
nor U18592 (N_18592,N_11686,N_12696);
and U18593 (N_18593,N_10771,N_11957);
xor U18594 (N_18594,N_11227,N_11149);
nor U18595 (N_18595,N_11539,N_10680);
and U18596 (N_18596,N_14413,N_14809);
nand U18597 (N_18597,N_14193,N_12393);
xnor U18598 (N_18598,N_11475,N_11121);
xor U18599 (N_18599,N_12646,N_12191);
nand U18600 (N_18600,N_11275,N_11239);
nor U18601 (N_18601,N_12752,N_14632);
and U18602 (N_18602,N_14208,N_12390);
nor U18603 (N_18603,N_10442,N_14534);
and U18604 (N_18604,N_14161,N_13684);
and U18605 (N_18605,N_11127,N_13030);
nand U18606 (N_18606,N_10169,N_14542);
nor U18607 (N_18607,N_14506,N_13797);
nand U18608 (N_18608,N_13656,N_10447);
nor U18609 (N_18609,N_10890,N_12400);
nand U18610 (N_18610,N_11979,N_11963);
nor U18611 (N_18611,N_12599,N_13570);
or U18612 (N_18612,N_12456,N_14291);
or U18613 (N_18613,N_13845,N_11669);
nor U18614 (N_18614,N_13109,N_13743);
and U18615 (N_18615,N_10578,N_11111);
nor U18616 (N_18616,N_14187,N_13445);
or U18617 (N_18617,N_12426,N_12268);
or U18618 (N_18618,N_10989,N_12227);
nor U18619 (N_18619,N_14917,N_13189);
and U18620 (N_18620,N_12471,N_12551);
nand U18621 (N_18621,N_10396,N_13384);
or U18622 (N_18622,N_12696,N_14060);
or U18623 (N_18623,N_12685,N_12434);
nor U18624 (N_18624,N_14167,N_12006);
nor U18625 (N_18625,N_12042,N_10931);
xnor U18626 (N_18626,N_10379,N_10082);
nor U18627 (N_18627,N_12400,N_11626);
nor U18628 (N_18628,N_14429,N_10993);
and U18629 (N_18629,N_12390,N_14693);
nor U18630 (N_18630,N_13788,N_10719);
nor U18631 (N_18631,N_11922,N_14677);
xnor U18632 (N_18632,N_10650,N_13175);
and U18633 (N_18633,N_10458,N_13032);
or U18634 (N_18634,N_11284,N_12721);
nand U18635 (N_18635,N_14736,N_10293);
or U18636 (N_18636,N_14455,N_11238);
xor U18637 (N_18637,N_14755,N_14319);
nor U18638 (N_18638,N_14757,N_11836);
or U18639 (N_18639,N_12795,N_12602);
and U18640 (N_18640,N_12380,N_14295);
nand U18641 (N_18641,N_13324,N_14735);
nand U18642 (N_18642,N_13624,N_14047);
or U18643 (N_18643,N_12039,N_12897);
or U18644 (N_18644,N_10782,N_12700);
and U18645 (N_18645,N_11873,N_11305);
and U18646 (N_18646,N_14071,N_11396);
nor U18647 (N_18647,N_11278,N_14784);
or U18648 (N_18648,N_11322,N_12190);
xor U18649 (N_18649,N_13046,N_13304);
and U18650 (N_18650,N_14089,N_13066);
nand U18651 (N_18651,N_10058,N_12315);
xor U18652 (N_18652,N_13846,N_12560);
and U18653 (N_18653,N_12546,N_14386);
or U18654 (N_18654,N_11843,N_10899);
xor U18655 (N_18655,N_11915,N_11208);
or U18656 (N_18656,N_14172,N_10350);
xnor U18657 (N_18657,N_10197,N_13583);
or U18658 (N_18658,N_12801,N_10272);
xnor U18659 (N_18659,N_10276,N_14285);
or U18660 (N_18660,N_13109,N_13587);
nor U18661 (N_18661,N_14649,N_14933);
or U18662 (N_18662,N_12036,N_11988);
nor U18663 (N_18663,N_10384,N_10076);
xor U18664 (N_18664,N_10646,N_10295);
nor U18665 (N_18665,N_12916,N_10817);
and U18666 (N_18666,N_13183,N_14815);
nand U18667 (N_18667,N_10895,N_10573);
xor U18668 (N_18668,N_13711,N_13108);
and U18669 (N_18669,N_13903,N_12615);
nor U18670 (N_18670,N_14270,N_13211);
or U18671 (N_18671,N_13784,N_10657);
xor U18672 (N_18672,N_11018,N_10807);
or U18673 (N_18673,N_13718,N_10050);
or U18674 (N_18674,N_10766,N_11451);
nor U18675 (N_18675,N_10815,N_10475);
nor U18676 (N_18676,N_12636,N_11640);
nor U18677 (N_18677,N_11416,N_13583);
or U18678 (N_18678,N_13405,N_12126);
xnor U18679 (N_18679,N_10667,N_11742);
nand U18680 (N_18680,N_11095,N_13597);
xor U18681 (N_18681,N_14749,N_14069);
and U18682 (N_18682,N_11278,N_14801);
xor U18683 (N_18683,N_11476,N_12034);
or U18684 (N_18684,N_14134,N_13196);
and U18685 (N_18685,N_12194,N_14516);
and U18686 (N_18686,N_14076,N_10108);
nand U18687 (N_18687,N_12864,N_12098);
and U18688 (N_18688,N_14466,N_12360);
and U18689 (N_18689,N_13897,N_12587);
or U18690 (N_18690,N_14652,N_13425);
or U18691 (N_18691,N_11696,N_12732);
nand U18692 (N_18692,N_13670,N_12122);
nor U18693 (N_18693,N_13379,N_10455);
or U18694 (N_18694,N_11310,N_12311);
nor U18695 (N_18695,N_14383,N_11505);
or U18696 (N_18696,N_11091,N_10253);
and U18697 (N_18697,N_14063,N_12414);
nand U18698 (N_18698,N_13949,N_13350);
or U18699 (N_18699,N_11995,N_13457);
nand U18700 (N_18700,N_12519,N_12377);
or U18701 (N_18701,N_12756,N_11854);
and U18702 (N_18702,N_12714,N_13073);
nand U18703 (N_18703,N_11501,N_11213);
or U18704 (N_18704,N_14372,N_10038);
nand U18705 (N_18705,N_14244,N_10769);
nand U18706 (N_18706,N_12953,N_11184);
nand U18707 (N_18707,N_12692,N_10055);
nand U18708 (N_18708,N_11307,N_13054);
xnor U18709 (N_18709,N_11783,N_11600);
and U18710 (N_18710,N_11242,N_13588);
nand U18711 (N_18711,N_11343,N_13993);
and U18712 (N_18712,N_10339,N_12745);
nor U18713 (N_18713,N_10753,N_12252);
nor U18714 (N_18714,N_11322,N_13961);
or U18715 (N_18715,N_14696,N_10384);
xor U18716 (N_18716,N_13019,N_10887);
or U18717 (N_18717,N_13008,N_12164);
nand U18718 (N_18718,N_12410,N_14060);
nor U18719 (N_18719,N_10024,N_11517);
nand U18720 (N_18720,N_12873,N_13664);
or U18721 (N_18721,N_10203,N_11680);
xnor U18722 (N_18722,N_14143,N_12785);
nand U18723 (N_18723,N_11903,N_12903);
nand U18724 (N_18724,N_12631,N_12417);
nor U18725 (N_18725,N_13169,N_12165);
or U18726 (N_18726,N_12203,N_14869);
or U18727 (N_18727,N_12126,N_14413);
or U18728 (N_18728,N_10293,N_10151);
and U18729 (N_18729,N_12692,N_12256);
or U18730 (N_18730,N_10478,N_12103);
or U18731 (N_18731,N_14717,N_12952);
nor U18732 (N_18732,N_13410,N_10965);
and U18733 (N_18733,N_13412,N_11945);
and U18734 (N_18734,N_12757,N_11454);
nand U18735 (N_18735,N_13545,N_10637);
or U18736 (N_18736,N_14891,N_11779);
nor U18737 (N_18737,N_10133,N_12825);
xor U18738 (N_18738,N_13031,N_12214);
nor U18739 (N_18739,N_10794,N_11816);
or U18740 (N_18740,N_10377,N_13177);
xnor U18741 (N_18741,N_12983,N_14506);
xor U18742 (N_18742,N_11480,N_14045);
nor U18743 (N_18743,N_12028,N_11717);
nor U18744 (N_18744,N_10771,N_14676);
and U18745 (N_18745,N_12473,N_12825);
nand U18746 (N_18746,N_11267,N_12152);
nand U18747 (N_18747,N_14956,N_11448);
or U18748 (N_18748,N_14606,N_12338);
xnor U18749 (N_18749,N_11599,N_14843);
nand U18750 (N_18750,N_12086,N_14364);
nor U18751 (N_18751,N_14426,N_14695);
nor U18752 (N_18752,N_14021,N_14192);
nand U18753 (N_18753,N_11923,N_10130);
nor U18754 (N_18754,N_12259,N_14627);
or U18755 (N_18755,N_10554,N_13551);
nand U18756 (N_18756,N_13849,N_11246);
or U18757 (N_18757,N_13004,N_14286);
and U18758 (N_18758,N_12338,N_13475);
nor U18759 (N_18759,N_10471,N_14628);
nand U18760 (N_18760,N_11088,N_10917);
or U18761 (N_18761,N_14835,N_11086);
or U18762 (N_18762,N_14777,N_14607);
nand U18763 (N_18763,N_12403,N_12529);
nor U18764 (N_18764,N_12285,N_13429);
nor U18765 (N_18765,N_10862,N_10472);
nor U18766 (N_18766,N_10642,N_12836);
nor U18767 (N_18767,N_14319,N_11728);
nand U18768 (N_18768,N_12532,N_11347);
xnor U18769 (N_18769,N_14840,N_10875);
nand U18770 (N_18770,N_12142,N_11471);
nand U18771 (N_18771,N_13395,N_10934);
nor U18772 (N_18772,N_13312,N_10728);
and U18773 (N_18773,N_10439,N_12700);
nand U18774 (N_18774,N_12882,N_10103);
or U18775 (N_18775,N_12122,N_13964);
nand U18776 (N_18776,N_13055,N_12406);
nand U18777 (N_18777,N_14875,N_14464);
nor U18778 (N_18778,N_12446,N_14855);
xnor U18779 (N_18779,N_11915,N_14164);
nand U18780 (N_18780,N_14684,N_13342);
and U18781 (N_18781,N_10971,N_10838);
and U18782 (N_18782,N_14406,N_13091);
nor U18783 (N_18783,N_10685,N_12759);
nor U18784 (N_18784,N_13733,N_13534);
xnor U18785 (N_18785,N_12194,N_13962);
nor U18786 (N_18786,N_14009,N_11523);
nand U18787 (N_18787,N_14165,N_12041);
nand U18788 (N_18788,N_14344,N_10493);
or U18789 (N_18789,N_13278,N_13330);
nand U18790 (N_18790,N_13313,N_10858);
nor U18791 (N_18791,N_13445,N_14810);
nor U18792 (N_18792,N_13316,N_10708);
or U18793 (N_18793,N_14835,N_12812);
nor U18794 (N_18794,N_11997,N_11371);
nor U18795 (N_18795,N_10345,N_12249);
nor U18796 (N_18796,N_11629,N_11503);
or U18797 (N_18797,N_13860,N_11349);
or U18798 (N_18798,N_12819,N_10944);
or U18799 (N_18799,N_12850,N_14948);
and U18800 (N_18800,N_10690,N_11872);
nand U18801 (N_18801,N_11209,N_13335);
xor U18802 (N_18802,N_13010,N_14285);
and U18803 (N_18803,N_11372,N_10839);
and U18804 (N_18804,N_14832,N_12386);
nand U18805 (N_18805,N_13029,N_11805);
nor U18806 (N_18806,N_12659,N_10098);
and U18807 (N_18807,N_13387,N_10309);
xor U18808 (N_18808,N_14450,N_12916);
and U18809 (N_18809,N_11714,N_13103);
nor U18810 (N_18810,N_11475,N_10132);
and U18811 (N_18811,N_14625,N_11820);
nor U18812 (N_18812,N_14946,N_13964);
nand U18813 (N_18813,N_14861,N_10963);
nor U18814 (N_18814,N_10152,N_12238);
or U18815 (N_18815,N_10613,N_10211);
and U18816 (N_18816,N_14137,N_14895);
nor U18817 (N_18817,N_13165,N_11870);
nor U18818 (N_18818,N_10275,N_14849);
nor U18819 (N_18819,N_14203,N_10096);
xnor U18820 (N_18820,N_11122,N_13492);
nor U18821 (N_18821,N_14650,N_10946);
nand U18822 (N_18822,N_10404,N_11116);
or U18823 (N_18823,N_10463,N_10627);
and U18824 (N_18824,N_14714,N_12872);
xor U18825 (N_18825,N_12191,N_14318);
or U18826 (N_18826,N_13511,N_12651);
nor U18827 (N_18827,N_11819,N_10707);
xnor U18828 (N_18828,N_13057,N_11957);
or U18829 (N_18829,N_10449,N_13332);
nand U18830 (N_18830,N_11060,N_11514);
or U18831 (N_18831,N_12636,N_10654);
nor U18832 (N_18832,N_10895,N_12700);
nor U18833 (N_18833,N_11411,N_12578);
xor U18834 (N_18834,N_11076,N_10538);
and U18835 (N_18835,N_11710,N_13811);
nor U18836 (N_18836,N_12521,N_14918);
nand U18837 (N_18837,N_13926,N_14554);
and U18838 (N_18838,N_13296,N_11351);
or U18839 (N_18839,N_12101,N_14885);
nor U18840 (N_18840,N_14934,N_12710);
nor U18841 (N_18841,N_12205,N_11621);
and U18842 (N_18842,N_10136,N_12619);
or U18843 (N_18843,N_14512,N_11446);
nor U18844 (N_18844,N_13561,N_11393);
nor U18845 (N_18845,N_10114,N_10762);
or U18846 (N_18846,N_14150,N_13916);
or U18847 (N_18847,N_12141,N_12947);
nor U18848 (N_18848,N_11325,N_10123);
and U18849 (N_18849,N_10887,N_12689);
xnor U18850 (N_18850,N_14677,N_14367);
nand U18851 (N_18851,N_10518,N_10682);
or U18852 (N_18852,N_13119,N_10640);
xor U18853 (N_18853,N_12816,N_14800);
or U18854 (N_18854,N_11125,N_12069);
or U18855 (N_18855,N_14736,N_14281);
xor U18856 (N_18856,N_14388,N_12073);
nor U18857 (N_18857,N_10237,N_11000);
nor U18858 (N_18858,N_10422,N_13293);
or U18859 (N_18859,N_14152,N_10449);
nor U18860 (N_18860,N_13054,N_13782);
nor U18861 (N_18861,N_10510,N_13597);
nand U18862 (N_18862,N_11572,N_14004);
or U18863 (N_18863,N_10940,N_12994);
or U18864 (N_18864,N_10931,N_11640);
or U18865 (N_18865,N_14024,N_14184);
or U18866 (N_18866,N_14775,N_12445);
and U18867 (N_18867,N_14337,N_10267);
nand U18868 (N_18868,N_12120,N_13345);
and U18869 (N_18869,N_11240,N_10698);
nand U18870 (N_18870,N_10693,N_13282);
or U18871 (N_18871,N_12838,N_10385);
nand U18872 (N_18872,N_14151,N_14914);
or U18873 (N_18873,N_11130,N_11804);
and U18874 (N_18874,N_13914,N_10216);
nand U18875 (N_18875,N_12659,N_11007);
and U18876 (N_18876,N_14833,N_13790);
and U18877 (N_18877,N_10446,N_10655);
nand U18878 (N_18878,N_11283,N_11876);
xnor U18879 (N_18879,N_14619,N_12378);
and U18880 (N_18880,N_11497,N_12537);
nor U18881 (N_18881,N_13721,N_10509);
xor U18882 (N_18882,N_14745,N_14345);
and U18883 (N_18883,N_10449,N_11706);
nand U18884 (N_18884,N_13396,N_11372);
or U18885 (N_18885,N_14778,N_14717);
nand U18886 (N_18886,N_10057,N_10943);
or U18887 (N_18887,N_12618,N_13674);
and U18888 (N_18888,N_11297,N_14669);
or U18889 (N_18889,N_12796,N_14735);
or U18890 (N_18890,N_14368,N_12611);
and U18891 (N_18891,N_12570,N_14844);
nand U18892 (N_18892,N_11279,N_10574);
or U18893 (N_18893,N_11957,N_14520);
or U18894 (N_18894,N_14752,N_14967);
xor U18895 (N_18895,N_12368,N_13842);
nand U18896 (N_18896,N_13668,N_11949);
nor U18897 (N_18897,N_13677,N_10238);
or U18898 (N_18898,N_10570,N_12663);
xnor U18899 (N_18899,N_14145,N_10841);
or U18900 (N_18900,N_14401,N_12045);
and U18901 (N_18901,N_13486,N_14138);
nor U18902 (N_18902,N_14879,N_13892);
nor U18903 (N_18903,N_11270,N_10223);
or U18904 (N_18904,N_12477,N_12573);
xnor U18905 (N_18905,N_10989,N_11260);
or U18906 (N_18906,N_11819,N_10314);
and U18907 (N_18907,N_14332,N_14747);
or U18908 (N_18908,N_12334,N_14548);
nor U18909 (N_18909,N_11243,N_12603);
and U18910 (N_18910,N_14029,N_14812);
or U18911 (N_18911,N_11537,N_13622);
nand U18912 (N_18912,N_10069,N_13082);
nand U18913 (N_18913,N_11058,N_14992);
or U18914 (N_18914,N_14088,N_11585);
and U18915 (N_18915,N_14665,N_11749);
nor U18916 (N_18916,N_14591,N_14811);
nor U18917 (N_18917,N_14006,N_12923);
or U18918 (N_18918,N_11774,N_12885);
nand U18919 (N_18919,N_11467,N_14959);
nand U18920 (N_18920,N_13452,N_12393);
nor U18921 (N_18921,N_14007,N_12573);
nand U18922 (N_18922,N_12875,N_13071);
and U18923 (N_18923,N_14354,N_12183);
or U18924 (N_18924,N_11052,N_11688);
and U18925 (N_18925,N_11751,N_14787);
nand U18926 (N_18926,N_12408,N_10060);
nand U18927 (N_18927,N_12457,N_13816);
and U18928 (N_18928,N_14194,N_10478);
nand U18929 (N_18929,N_12697,N_12505);
or U18930 (N_18930,N_10921,N_11795);
nor U18931 (N_18931,N_12568,N_14270);
nor U18932 (N_18932,N_14964,N_13974);
nand U18933 (N_18933,N_10669,N_13804);
or U18934 (N_18934,N_12795,N_14541);
xnor U18935 (N_18935,N_12750,N_14014);
and U18936 (N_18936,N_12396,N_12111);
nand U18937 (N_18937,N_11589,N_11221);
nand U18938 (N_18938,N_10705,N_12576);
or U18939 (N_18939,N_10890,N_10126);
nand U18940 (N_18940,N_11634,N_12712);
nor U18941 (N_18941,N_11646,N_12316);
or U18942 (N_18942,N_14022,N_12410);
nor U18943 (N_18943,N_13484,N_13004);
nand U18944 (N_18944,N_13368,N_10814);
nor U18945 (N_18945,N_11632,N_12130);
and U18946 (N_18946,N_10432,N_14348);
nand U18947 (N_18947,N_12828,N_13093);
nor U18948 (N_18948,N_13090,N_11769);
or U18949 (N_18949,N_14140,N_12177);
nor U18950 (N_18950,N_14584,N_13466);
nand U18951 (N_18951,N_11288,N_12992);
nor U18952 (N_18952,N_13718,N_10358);
nor U18953 (N_18953,N_10378,N_13135);
or U18954 (N_18954,N_10862,N_13396);
or U18955 (N_18955,N_14200,N_13016);
nor U18956 (N_18956,N_13593,N_14138);
and U18957 (N_18957,N_11480,N_14278);
or U18958 (N_18958,N_12838,N_12768);
or U18959 (N_18959,N_14816,N_10013);
or U18960 (N_18960,N_13724,N_11918);
and U18961 (N_18961,N_13495,N_10457);
xor U18962 (N_18962,N_13807,N_12268);
and U18963 (N_18963,N_13006,N_14279);
and U18964 (N_18964,N_13350,N_13875);
xor U18965 (N_18965,N_14540,N_12768);
nand U18966 (N_18966,N_14380,N_13358);
nor U18967 (N_18967,N_14295,N_10787);
and U18968 (N_18968,N_14618,N_11869);
nand U18969 (N_18969,N_14798,N_12436);
nor U18970 (N_18970,N_13977,N_12262);
or U18971 (N_18971,N_12070,N_12078);
and U18972 (N_18972,N_10296,N_13623);
xnor U18973 (N_18973,N_13270,N_12566);
nand U18974 (N_18974,N_12805,N_11283);
nand U18975 (N_18975,N_10355,N_10020);
or U18976 (N_18976,N_13768,N_13001);
or U18977 (N_18977,N_11981,N_13328);
nand U18978 (N_18978,N_10597,N_12838);
nor U18979 (N_18979,N_11659,N_10695);
or U18980 (N_18980,N_12544,N_14996);
nor U18981 (N_18981,N_14617,N_13299);
nand U18982 (N_18982,N_13705,N_10924);
and U18983 (N_18983,N_12278,N_12756);
nand U18984 (N_18984,N_13984,N_10367);
nor U18985 (N_18985,N_14038,N_13198);
nor U18986 (N_18986,N_14551,N_11178);
nor U18987 (N_18987,N_11915,N_13820);
nand U18988 (N_18988,N_10054,N_14060);
or U18989 (N_18989,N_11606,N_11917);
nand U18990 (N_18990,N_12146,N_13940);
nand U18991 (N_18991,N_14037,N_11159);
xnor U18992 (N_18992,N_11626,N_14906);
nor U18993 (N_18993,N_10242,N_14642);
or U18994 (N_18994,N_10603,N_13751);
and U18995 (N_18995,N_14126,N_11279);
nor U18996 (N_18996,N_11339,N_10565);
or U18997 (N_18997,N_10010,N_10879);
nor U18998 (N_18998,N_13991,N_14438);
or U18999 (N_18999,N_10569,N_12955);
or U19000 (N_19000,N_13460,N_12186);
and U19001 (N_19001,N_10770,N_10926);
nor U19002 (N_19002,N_12397,N_14663);
nand U19003 (N_19003,N_12719,N_13208);
nor U19004 (N_19004,N_14364,N_11592);
nor U19005 (N_19005,N_13497,N_11816);
and U19006 (N_19006,N_10950,N_14522);
or U19007 (N_19007,N_14621,N_12047);
and U19008 (N_19008,N_12982,N_13448);
nand U19009 (N_19009,N_14664,N_14412);
nor U19010 (N_19010,N_14286,N_13405);
nand U19011 (N_19011,N_11676,N_11857);
xnor U19012 (N_19012,N_10890,N_11267);
nand U19013 (N_19013,N_10365,N_14709);
nand U19014 (N_19014,N_11730,N_10174);
nand U19015 (N_19015,N_13953,N_12554);
nor U19016 (N_19016,N_11394,N_14264);
and U19017 (N_19017,N_12903,N_14719);
nor U19018 (N_19018,N_11502,N_14185);
and U19019 (N_19019,N_10676,N_10340);
or U19020 (N_19020,N_14881,N_13362);
or U19021 (N_19021,N_14836,N_13669);
nand U19022 (N_19022,N_14787,N_12519);
xor U19023 (N_19023,N_13615,N_12361);
or U19024 (N_19024,N_11286,N_13906);
or U19025 (N_19025,N_10498,N_14602);
nand U19026 (N_19026,N_11694,N_11407);
nor U19027 (N_19027,N_11080,N_10921);
nor U19028 (N_19028,N_11792,N_14979);
nand U19029 (N_19029,N_10971,N_11463);
nor U19030 (N_19030,N_10303,N_13874);
or U19031 (N_19031,N_14220,N_12845);
xnor U19032 (N_19032,N_14965,N_13600);
nand U19033 (N_19033,N_11315,N_10020);
and U19034 (N_19034,N_12028,N_14209);
nand U19035 (N_19035,N_14438,N_14643);
nand U19036 (N_19036,N_13033,N_12803);
nand U19037 (N_19037,N_10358,N_10566);
xor U19038 (N_19038,N_13683,N_13439);
or U19039 (N_19039,N_14131,N_10534);
nor U19040 (N_19040,N_13963,N_11195);
and U19041 (N_19041,N_11223,N_10487);
xor U19042 (N_19042,N_12616,N_13560);
and U19043 (N_19043,N_13351,N_10855);
and U19044 (N_19044,N_12808,N_14727);
or U19045 (N_19045,N_13872,N_14905);
nand U19046 (N_19046,N_11713,N_13926);
nand U19047 (N_19047,N_10677,N_11604);
and U19048 (N_19048,N_11945,N_11062);
or U19049 (N_19049,N_13923,N_13932);
nor U19050 (N_19050,N_13222,N_10904);
nor U19051 (N_19051,N_14125,N_10072);
and U19052 (N_19052,N_13943,N_11265);
or U19053 (N_19053,N_10415,N_10672);
or U19054 (N_19054,N_10206,N_11569);
nor U19055 (N_19055,N_14671,N_13803);
nor U19056 (N_19056,N_14752,N_13761);
or U19057 (N_19057,N_10469,N_14018);
nor U19058 (N_19058,N_11099,N_14557);
or U19059 (N_19059,N_13979,N_14400);
nor U19060 (N_19060,N_10928,N_10289);
nand U19061 (N_19061,N_14969,N_12878);
and U19062 (N_19062,N_14582,N_10239);
and U19063 (N_19063,N_11398,N_11441);
or U19064 (N_19064,N_14095,N_12721);
xnor U19065 (N_19065,N_11185,N_13073);
xor U19066 (N_19066,N_12126,N_14686);
or U19067 (N_19067,N_13194,N_12710);
nand U19068 (N_19068,N_10158,N_12952);
nor U19069 (N_19069,N_11597,N_13571);
or U19070 (N_19070,N_10193,N_13435);
and U19071 (N_19071,N_13225,N_10816);
or U19072 (N_19072,N_14101,N_13116);
nand U19073 (N_19073,N_14579,N_14222);
or U19074 (N_19074,N_14702,N_13575);
or U19075 (N_19075,N_10512,N_13945);
and U19076 (N_19076,N_14467,N_11544);
nor U19077 (N_19077,N_10124,N_13195);
or U19078 (N_19078,N_11940,N_13922);
nor U19079 (N_19079,N_14533,N_13187);
and U19080 (N_19080,N_14901,N_13607);
nor U19081 (N_19081,N_11810,N_12260);
or U19082 (N_19082,N_10236,N_12158);
nor U19083 (N_19083,N_12362,N_10705);
or U19084 (N_19084,N_11277,N_10166);
nor U19085 (N_19085,N_13492,N_11612);
or U19086 (N_19086,N_14122,N_13652);
or U19087 (N_19087,N_10861,N_11235);
nand U19088 (N_19088,N_11899,N_14929);
or U19089 (N_19089,N_14358,N_10243);
and U19090 (N_19090,N_10584,N_12345);
nor U19091 (N_19091,N_13353,N_14452);
nand U19092 (N_19092,N_14175,N_11638);
nor U19093 (N_19093,N_10354,N_11942);
xor U19094 (N_19094,N_10260,N_13931);
and U19095 (N_19095,N_14791,N_13180);
nand U19096 (N_19096,N_11855,N_14627);
and U19097 (N_19097,N_14074,N_13537);
and U19098 (N_19098,N_10710,N_13525);
nor U19099 (N_19099,N_14844,N_11965);
nor U19100 (N_19100,N_10865,N_10090);
or U19101 (N_19101,N_12685,N_13182);
or U19102 (N_19102,N_12951,N_13963);
or U19103 (N_19103,N_11576,N_12939);
xnor U19104 (N_19104,N_14162,N_14081);
or U19105 (N_19105,N_11016,N_11169);
nand U19106 (N_19106,N_10323,N_10370);
or U19107 (N_19107,N_12455,N_10188);
and U19108 (N_19108,N_13244,N_12569);
nor U19109 (N_19109,N_14386,N_11494);
nor U19110 (N_19110,N_10863,N_12809);
and U19111 (N_19111,N_11777,N_12643);
nor U19112 (N_19112,N_13986,N_11343);
xor U19113 (N_19113,N_10302,N_14014);
nand U19114 (N_19114,N_14782,N_10701);
and U19115 (N_19115,N_12401,N_10919);
or U19116 (N_19116,N_12612,N_10627);
nor U19117 (N_19117,N_13139,N_10694);
and U19118 (N_19118,N_12915,N_10296);
nand U19119 (N_19119,N_11414,N_11291);
nand U19120 (N_19120,N_14962,N_14801);
nand U19121 (N_19121,N_10203,N_13561);
nor U19122 (N_19122,N_12832,N_12969);
nand U19123 (N_19123,N_10197,N_14144);
or U19124 (N_19124,N_12096,N_12330);
nor U19125 (N_19125,N_10082,N_14788);
or U19126 (N_19126,N_11821,N_13369);
or U19127 (N_19127,N_14643,N_12702);
or U19128 (N_19128,N_12700,N_10507);
and U19129 (N_19129,N_12812,N_12319);
or U19130 (N_19130,N_14166,N_11079);
or U19131 (N_19131,N_12854,N_12301);
xnor U19132 (N_19132,N_12247,N_12582);
nor U19133 (N_19133,N_11086,N_12232);
or U19134 (N_19134,N_11730,N_12151);
xor U19135 (N_19135,N_12627,N_11673);
or U19136 (N_19136,N_14154,N_13256);
and U19137 (N_19137,N_13249,N_11691);
and U19138 (N_19138,N_10077,N_13891);
and U19139 (N_19139,N_13540,N_13480);
or U19140 (N_19140,N_14422,N_12957);
and U19141 (N_19141,N_10083,N_11050);
and U19142 (N_19142,N_14222,N_14626);
nor U19143 (N_19143,N_12148,N_11965);
nand U19144 (N_19144,N_12682,N_12224);
nor U19145 (N_19145,N_12219,N_12105);
and U19146 (N_19146,N_14022,N_10935);
and U19147 (N_19147,N_12706,N_10159);
nor U19148 (N_19148,N_14354,N_12939);
nand U19149 (N_19149,N_13021,N_14792);
nand U19150 (N_19150,N_10219,N_10253);
and U19151 (N_19151,N_10819,N_10882);
xor U19152 (N_19152,N_14021,N_12132);
nor U19153 (N_19153,N_11516,N_12299);
xnor U19154 (N_19154,N_12930,N_13922);
nand U19155 (N_19155,N_13792,N_12613);
nor U19156 (N_19156,N_11234,N_13434);
or U19157 (N_19157,N_10834,N_10314);
nor U19158 (N_19158,N_12018,N_11046);
nor U19159 (N_19159,N_11548,N_10316);
or U19160 (N_19160,N_14391,N_10895);
nand U19161 (N_19161,N_13159,N_11594);
or U19162 (N_19162,N_12032,N_12491);
nor U19163 (N_19163,N_14784,N_13153);
nor U19164 (N_19164,N_13446,N_13664);
and U19165 (N_19165,N_12716,N_14925);
nor U19166 (N_19166,N_13127,N_12028);
xnor U19167 (N_19167,N_11985,N_11710);
nor U19168 (N_19168,N_11941,N_14971);
nor U19169 (N_19169,N_14268,N_14555);
and U19170 (N_19170,N_13460,N_14568);
or U19171 (N_19171,N_13343,N_11519);
and U19172 (N_19172,N_12912,N_14180);
nand U19173 (N_19173,N_12758,N_11298);
xor U19174 (N_19174,N_10765,N_10801);
and U19175 (N_19175,N_14446,N_13222);
and U19176 (N_19176,N_14518,N_11253);
xor U19177 (N_19177,N_10718,N_12728);
nor U19178 (N_19178,N_10269,N_11992);
and U19179 (N_19179,N_14702,N_11430);
nor U19180 (N_19180,N_11308,N_14105);
nand U19181 (N_19181,N_12670,N_10072);
or U19182 (N_19182,N_12447,N_11084);
nor U19183 (N_19183,N_14722,N_11396);
nand U19184 (N_19184,N_14298,N_11256);
nor U19185 (N_19185,N_11249,N_10412);
nor U19186 (N_19186,N_11733,N_11589);
nand U19187 (N_19187,N_12716,N_11297);
nand U19188 (N_19188,N_11062,N_14428);
or U19189 (N_19189,N_11157,N_11030);
or U19190 (N_19190,N_10190,N_13294);
xor U19191 (N_19191,N_11341,N_10746);
and U19192 (N_19192,N_10251,N_12646);
nor U19193 (N_19193,N_10074,N_13723);
and U19194 (N_19194,N_10250,N_12481);
xor U19195 (N_19195,N_11165,N_14186);
nor U19196 (N_19196,N_12607,N_12754);
and U19197 (N_19197,N_14030,N_11501);
and U19198 (N_19198,N_14950,N_11849);
nand U19199 (N_19199,N_13859,N_14330);
and U19200 (N_19200,N_10638,N_11812);
nand U19201 (N_19201,N_13924,N_11454);
and U19202 (N_19202,N_11463,N_10416);
nor U19203 (N_19203,N_10448,N_12816);
nand U19204 (N_19204,N_10563,N_10646);
xor U19205 (N_19205,N_13818,N_13554);
nand U19206 (N_19206,N_12616,N_10820);
xnor U19207 (N_19207,N_14892,N_10683);
or U19208 (N_19208,N_10322,N_13549);
and U19209 (N_19209,N_12309,N_13379);
xnor U19210 (N_19210,N_10711,N_10540);
xor U19211 (N_19211,N_12469,N_13630);
nand U19212 (N_19212,N_10847,N_11214);
xor U19213 (N_19213,N_14243,N_11857);
and U19214 (N_19214,N_14407,N_13151);
and U19215 (N_19215,N_12779,N_10326);
nor U19216 (N_19216,N_13568,N_13622);
nand U19217 (N_19217,N_12772,N_12722);
and U19218 (N_19218,N_12545,N_14059);
and U19219 (N_19219,N_13436,N_11209);
and U19220 (N_19220,N_12074,N_14907);
and U19221 (N_19221,N_14004,N_10608);
and U19222 (N_19222,N_13493,N_13534);
and U19223 (N_19223,N_12925,N_10558);
and U19224 (N_19224,N_12942,N_14990);
nor U19225 (N_19225,N_11767,N_11348);
xor U19226 (N_19226,N_13622,N_12562);
nor U19227 (N_19227,N_10287,N_10236);
nand U19228 (N_19228,N_14402,N_13462);
or U19229 (N_19229,N_14410,N_13595);
or U19230 (N_19230,N_14851,N_12421);
nand U19231 (N_19231,N_13914,N_11790);
or U19232 (N_19232,N_11748,N_14255);
and U19233 (N_19233,N_14381,N_12750);
or U19234 (N_19234,N_10939,N_14557);
nand U19235 (N_19235,N_10167,N_11886);
and U19236 (N_19236,N_13713,N_12413);
or U19237 (N_19237,N_13859,N_12917);
xor U19238 (N_19238,N_11013,N_11730);
and U19239 (N_19239,N_10442,N_12299);
and U19240 (N_19240,N_11093,N_14582);
and U19241 (N_19241,N_11948,N_14834);
and U19242 (N_19242,N_12840,N_14244);
nor U19243 (N_19243,N_10494,N_14690);
xor U19244 (N_19244,N_12059,N_14110);
nor U19245 (N_19245,N_12289,N_14108);
nor U19246 (N_19246,N_12221,N_13402);
or U19247 (N_19247,N_11051,N_14663);
nor U19248 (N_19248,N_10163,N_12441);
nor U19249 (N_19249,N_12220,N_14222);
and U19250 (N_19250,N_14365,N_13466);
nor U19251 (N_19251,N_11673,N_12919);
or U19252 (N_19252,N_12647,N_11446);
nand U19253 (N_19253,N_10871,N_13358);
nand U19254 (N_19254,N_11641,N_11142);
and U19255 (N_19255,N_12260,N_14925);
or U19256 (N_19256,N_10539,N_11786);
nor U19257 (N_19257,N_10970,N_11599);
and U19258 (N_19258,N_11408,N_13486);
nor U19259 (N_19259,N_13404,N_14774);
or U19260 (N_19260,N_10590,N_13051);
or U19261 (N_19261,N_10071,N_14352);
xor U19262 (N_19262,N_11344,N_13727);
and U19263 (N_19263,N_14223,N_11023);
or U19264 (N_19264,N_11582,N_13007);
nor U19265 (N_19265,N_13870,N_13565);
nor U19266 (N_19266,N_12975,N_10598);
nor U19267 (N_19267,N_11775,N_11617);
nor U19268 (N_19268,N_12450,N_13986);
and U19269 (N_19269,N_14500,N_14776);
nor U19270 (N_19270,N_11847,N_10953);
nor U19271 (N_19271,N_14973,N_12133);
nand U19272 (N_19272,N_13789,N_14442);
nor U19273 (N_19273,N_11660,N_12695);
nand U19274 (N_19274,N_14998,N_11340);
nor U19275 (N_19275,N_11335,N_11487);
and U19276 (N_19276,N_10588,N_11495);
nor U19277 (N_19277,N_13000,N_11640);
or U19278 (N_19278,N_13321,N_11263);
nand U19279 (N_19279,N_12618,N_14366);
or U19280 (N_19280,N_12043,N_10582);
xor U19281 (N_19281,N_11602,N_11059);
or U19282 (N_19282,N_12748,N_10711);
and U19283 (N_19283,N_13209,N_13173);
nand U19284 (N_19284,N_12188,N_14856);
and U19285 (N_19285,N_12647,N_11810);
or U19286 (N_19286,N_11239,N_12254);
and U19287 (N_19287,N_12459,N_11943);
or U19288 (N_19288,N_12294,N_10644);
and U19289 (N_19289,N_10839,N_11434);
or U19290 (N_19290,N_10042,N_13971);
or U19291 (N_19291,N_13358,N_14021);
nand U19292 (N_19292,N_11555,N_14072);
nand U19293 (N_19293,N_11023,N_12583);
and U19294 (N_19294,N_14678,N_14997);
or U19295 (N_19295,N_13822,N_14851);
xnor U19296 (N_19296,N_13479,N_10340);
nor U19297 (N_19297,N_11022,N_10838);
nand U19298 (N_19298,N_11995,N_10843);
or U19299 (N_19299,N_13518,N_12062);
nor U19300 (N_19300,N_13399,N_14529);
and U19301 (N_19301,N_14906,N_12686);
nor U19302 (N_19302,N_10284,N_13253);
nor U19303 (N_19303,N_12864,N_12412);
and U19304 (N_19304,N_14996,N_12518);
nor U19305 (N_19305,N_11551,N_11067);
or U19306 (N_19306,N_14857,N_11911);
xnor U19307 (N_19307,N_14183,N_12239);
and U19308 (N_19308,N_10097,N_10176);
nand U19309 (N_19309,N_10870,N_10873);
or U19310 (N_19310,N_10921,N_10391);
nor U19311 (N_19311,N_11052,N_12252);
nand U19312 (N_19312,N_11369,N_10851);
and U19313 (N_19313,N_11898,N_12961);
nor U19314 (N_19314,N_10399,N_13762);
nand U19315 (N_19315,N_14088,N_12585);
nand U19316 (N_19316,N_10440,N_12332);
and U19317 (N_19317,N_11564,N_10983);
nand U19318 (N_19318,N_14999,N_14361);
nor U19319 (N_19319,N_13540,N_14861);
or U19320 (N_19320,N_10594,N_11675);
nor U19321 (N_19321,N_11338,N_11990);
nand U19322 (N_19322,N_11148,N_11758);
nand U19323 (N_19323,N_11998,N_11842);
nand U19324 (N_19324,N_13325,N_10366);
nand U19325 (N_19325,N_10790,N_12467);
or U19326 (N_19326,N_14117,N_10181);
xor U19327 (N_19327,N_10818,N_13779);
or U19328 (N_19328,N_10389,N_12001);
and U19329 (N_19329,N_13038,N_12523);
and U19330 (N_19330,N_14509,N_10074);
nor U19331 (N_19331,N_13645,N_14775);
or U19332 (N_19332,N_11108,N_13516);
nor U19333 (N_19333,N_10988,N_10778);
and U19334 (N_19334,N_14929,N_10150);
nand U19335 (N_19335,N_12929,N_14043);
xnor U19336 (N_19336,N_11541,N_12496);
nand U19337 (N_19337,N_13401,N_12613);
and U19338 (N_19338,N_11940,N_10422);
nand U19339 (N_19339,N_13515,N_12276);
nor U19340 (N_19340,N_12396,N_13393);
nand U19341 (N_19341,N_12234,N_14091);
or U19342 (N_19342,N_10782,N_11980);
nand U19343 (N_19343,N_11046,N_13312);
or U19344 (N_19344,N_10441,N_12083);
nand U19345 (N_19345,N_14961,N_14372);
xnor U19346 (N_19346,N_10005,N_12668);
nand U19347 (N_19347,N_14804,N_10370);
and U19348 (N_19348,N_13747,N_11722);
or U19349 (N_19349,N_11351,N_11532);
nor U19350 (N_19350,N_10801,N_10907);
xor U19351 (N_19351,N_14440,N_11035);
nor U19352 (N_19352,N_13982,N_12945);
and U19353 (N_19353,N_12998,N_13473);
and U19354 (N_19354,N_11379,N_14582);
and U19355 (N_19355,N_14530,N_10652);
and U19356 (N_19356,N_11031,N_13494);
and U19357 (N_19357,N_10390,N_10437);
or U19358 (N_19358,N_13723,N_12916);
nand U19359 (N_19359,N_13141,N_12938);
xnor U19360 (N_19360,N_10767,N_10121);
nor U19361 (N_19361,N_10695,N_10889);
nand U19362 (N_19362,N_14543,N_14516);
nor U19363 (N_19363,N_10233,N_14508);
nor U19364 (N_19364,N_13702,N_13233);
nand U19365 (N_19365,N_12327,N_14388);
xor U19366 (N_19366,N_11835,N_13296);
and U19367 (N_19367,N_10166,N_10185);
nand U19368 (N_19368,N_10830,N_13664);
nor U19369 (N_19369,N_14673,N_10380);
nand U19370 (N_19370,N_11398,N_14287);
nor U19371 (N_19371,N_14413,N_10434);
and U19372 (N_19372,N_13381,N_14557);
or U19373 (N_19373,N_11149,N_11260);
nand U19374 (N_19374,N_13538,N_13140);
nor U19375 (N_19375,N_14719,N_14865);
nand U19376 (N_19376,N_10115,N_12378);
nand U19377 (N_19377,N_13819,N_13003);
nor U19378 (N_19378,N_10518,N_11021);
xor U19379 (N_19379,N_10509,N_10555);
nor U19380 (N_19380,N_10508,N_11726);
nand U19381 (N_19381,N_10219,N_13567);
nor U19382 (N_19382,N_12746,N_10454);
and U19383 (N_19383,N_10646,N_14950);
xnor U19384 (N_19384,N_11900,N_10676);
xnor U19385 (N_19385,N_11372,N_13667);
or U19386 (N_19386,N_12805,N_11855);
and U19387 (N_19387,N_11738,N_10334);
or U19388 (N_19388,N_13026,N_11461);
nor U19389 (N_19389,N_10475,N_13758);
nand U19390 (N_19390,N_13467,N_10499);
xnor U19391 (N_19391,N_10371,N_12255);
or U19392 (N_19392,N_10784,N_14733);
xor U19393 (N_19393,N_12710,N_14133);
and U19394 (N_19394,N_12477,N_12681);
xnor U19395 (N_19395,N_10443,N_14035);
or U19396 (N_19396,N_11713,N_13402);
xnor U19397 (N_19397,N_11143,N_10937);
and U19398 (N_19398,N_14065,N_14105);
and U19399 (N_19399,N_14278,N_14408);
nor U19400 (N_19400,N_14108,N_12606);
nor U19401 (N_19401,N_12905,N_11411);
xnor U19402 (N_19402,N_13569,N_13268);
or U19403 (N_19403,N_13209,N_12953);
xor U19404 (N_19404,N_13157,N_10181);
nand U19405 (N_19405,N_13436,N_12720);
and U19406 (N_19406,N_10468,N_10840);
and U19407 (N_19407,N_10156,N_13210);
nand U19408 (N_19408,N_12750,N_12763);
or U19409 (N_19409,N_12901,N_11455);
xor U19410 (N_19410,N_10789,N_11671);
xor U19411 (N_19411,N_13782,N_13398);
xor U19412 (N_19412,N_10559,N_11641);
nor U19413 (N_19413,N_11645,N_14837);
or U19414 (N_19414,N_14565,N_10637);
or U19415 (N_19415,N_13753,N_10100);
nand U19416 (N_19416,N_13469,N_12853);
nor U19417 (N_19417,N_14931,N_14837);
nor U19418 (N_19418,N_10991,N_14581);
or U19419 (N_19419,N_13720,N_13610);
nor U19420 (N_19420,N_14347,N_11316);
or U19421 (N_19421,N_11776,N_13976);
nor U19422 (N_19422,N_11024,N_11464);
nand U19423 (N_19423,N_13804,N_11408);
nand U19424 (N_19424,N_12183,N_10313);
xor U19425 (N_19425,N_13967,N_13487);
nand U19426 (N_19426,N_13864,N_13322);
or U19427 (N_19427,N_12636,N_13396);
nand U19428 (N_19428,N_13471,N_14891);
xnor U19429 (N_19429,N_10144,N_14399);
and U19430 (N_19430,N_10245,N_12353);
nand U19431 (N_19431,N_14198,N_10780);
xnor U19432 (N_19432,N_11661,N_10843);
nand U19433 (N_19433,N_10029,N_10589);
nand U19434 (N_19434,N_10538,N_13853);
nand U19435 (N_19435,N_14502,N_11727);
xor U19436 (N_19436,N_11761,N_11123);
and U19437 (N_19437,N_12156,N_12115);
and U19438 (N_19438,N_14872,N_14523);
nor U19439 (N_19439,N_12873,N_13419);
nand U19440 (N_19440,N_13008,N_14444);
or U19441 (N_19441,N_11698,N_11020);
nand U19442 (N_19442,N_14867,N_13974);
or U19443 (N_19443,N_14439,N_11291);
nand U19444 (N_19444,N_11000,N_12059);
and U19445 (N_19445,N_11819,N_12073);
nand U19446 (N_19446,N_14788,N_13724);
nor U19447 (N_19447,N_13305,N_14024);
and U19448 (N_19448,N_12134,N_14592);
or U19449 (N_19449,N_12553,N_11460);
or U19450 (N_19450,N_10393,N_12551);
or U19451 (N_19451,N_14942,N_13090);
or U19452 (N_19452,N_11074,N_13291);
nor U19453 (N_19453,N_12669,N_14251);
and U19454 (N_19454,N_12467,N_10847);
or U19455 (N_19455,N_10626,N_13330);
and U19456 (N_19456,N_13630,N_12880);
nor U19457 (N_19457,N_14173,N_11594);
nor U19458 (N_19458,N_11727,N_10957);
xnor U19459 (N_19459,N_11911,N_14475);
nor U19460 (N_19460,N_13765,N_13037);
nand U19461 (N_19461,N_11151,N_10125);
nor U19462 (N_19462,N_13981,N_12532);
and U19463 (N_19463,N_12486,N_10072);
or U19464 (N_19464,N_10808,N_10794);
nand U19465 (N_19465,N_11093,N_12110);
or U19466 (N_19466,N_14929,N_14900);
or U19467 (N_19467,N_10043,N_12519);
or U19468 (N_19468,N_12832,N_10405);
nand U19469 (N_19469,N_11605,N_12724);
or U19470 (N_19470,N_11828,N_10291);
and U19471 (N_19471,N_13115,N_11540);
nand U19472 (N_19472,N_10980,N_12202);
nand U19473 (N_19473,N_14140,N_12332);
nand U19474 (N_19474,N_11340,N_12529);
nor U19475 (N_19475,N_10982,N_14361);
and U19476 (N_19476,N_11350,N_12895);
nor U19477 (N_19477,N_14985,N_12783);
and U19478 (N_19478,N_10940,N_12178);
or U19479 (N_19479,N_11538,N_12814);
and U19480 (N_19480,N_14158,N_13423);
xor U19481 (N_19481,N_11988,N_11091);
xor U19482 (N_19482,N_11198,N_13784);
and U19483 (N_19483,N_14226,N_11558);
nand U19484 (N_19484,N_10469,N_14830);
nor U19485 (N_19485,N_10300,N_14716);
or U19486 (N_19486,N_13828,N_13234);
nand U19487 (N_19487,N_14423,N_11035);
and U19488 (N_19488,N_12546,N_12737);
nand U19489 (N_19489,N_11698,N_12406);
nor U19490 (N_19490,N_13038,N_14661);
and U19491 (N_19491,N_13338,N_13199);
or U19492 (N_19492,N_12691,N_14209);
and U19493 (N_19493,N_12036,N_12799);
and U19494 (N_19494,N_10701,N_12518);
and U19495 (N_19495,N_10539,N_14491);
nand U19496 (N_19496,N_12710,N_10480);
xnor U19497 (N_19497,N_10728,N_14934);
nand U19498 (N_19498,N_12702,N_13339);
or U19499 (N_19499,N_13895,N_14643);
xor U19500 (N_19500,N_13140,N_11582);
xor U19501 (N_19501,N_14248,N_12320);
and U19502 (N_19502,N_11133,N_11975);
and U19503 (N_19503,N_10173,N_10139);
nor U19504 (N_19504,N_11769,N_11739);
nand U19505 (N_19505,N_10315,N_12737);
and U19506 (N_19506,N_14381,N_13789);
nand U19507 (N_19507,N_12351,N_11114);
or U19508 (N_19508,N_14112,N_11734);
and U19509 (N_19509,N_14242,N_10846);
nand U19510 (N_19510,N_11387,N_10430);
nor U19511 (N_19511,N_14690,N_13077);
nor U19512 (N_19512,N_10735,N_12557);
and U19513 (N_19513,N_12548,N_11511);
and U19514 (N_19514,N_11295,N_10088);
xor U19515 (N_19515,N_11522,N_11023);
or U19516 (N_19516,N_13424,N_14863);
nand U19517 (N_19517,N_12334,N_12040);
nor U19518 (N_19518,N_12074,N_10941);
nor U19519 (N_19519,N_11311,N_11894);
xor U19520 (N_19520,N_12974,N_10194);
or U19521 (N_19521,N_10698,N_14050);
nor U19522 (N_19522,N_11856,N_11022);
and U19523 (N_19523,N_10350,N_10629);
xor U19524 (N_19524,N_10676,N_13567);
or U19525 (N_19525,N_14898,N_14509);
nand U19526 (N_19526,N_12988,N_13733);
nor U19527 (N_19527,N_11564,N_14260);
nand U19528 (N_19528,N_11184,N_12004);
and U19529 (N_19529,N_14085,N_14043);
nand U19530 (N_19530,N_13177,N_13618);
and U19531 (N_19531,N_13691,N_14316);
or U19532 (N_19532,N_10076,N_10950);
xor U19533 (N_19533,N_11530,N_11950);
and U19534 (N_19534,N_13251,N_10480);
xor U19535 (N_19535,N_11692,N_10244);
nand U19536 (N_19536,N_10456,N_14525);
xor U19537 (N_19537,N_10836,N_13886);
nor U19538 (N_19538,N_12071,N_11469);
xnor U19539 (N_19539,N_10798,N_10812);
nand U19540 (N_19540,N_10601,N_13093);
nor U19541 (N_19541,N_14322,N_14933);
or U19542 (N_19542,N_13040,N_12568);
or U19543 (N_19543,N_11283,N_12188);
nand U19544 (N_19544,N_10894,N_14989);
xnor U19545 (N_19545,N_14661,N_13163);
and U19546 (N_19546,N_11605,N_13971);
or U19547 (N_19547,N_13185,N_12768);
nand U19548 (N_19548,N_11046,N_10519);
and U19549 (N_19549,N_14674,N_14105);
nor U19550 (N_19550,N_13423,N_13364);
nor U19551 (N_19551,N_13255,N_11710);
nor U19552 (N_19552,N_14377,N_11066);
or U19553 (N_19553,N_14595,N_11893);
nand U19554 (N_19554,N_13519,N_10007);
or U19555 (N_19555,N_12199,N_10629);
or U19556 (N_19556,N_14569,N_11484);
nand U19557 (N_19557,N_12708,N_14136);
xor U19558 (N_19558,N_14486,N_11113);
nand U19559 (N_19559,N_13912,N_14744);
and U19560 (N_19560,N_10816,N_14116);
or U19561 (N_19561,N_12243,N_11284);
and U19562 (N_19562,N_13574,N_13679);
nand U19563 (N_19563,N_14675,N_13440);
nor U19564 (N_19564,N_11316,N_14780);
nand U19565 (N_19565,N_13786,N_10855);
or U19566 (N_19566,N_10320,N_14858);
and U19567 (N_19567,N_13113,N_12767);
nand U19568 (N_19568,N_13000,N_14785);
and U19569 (N_19569,N_11363,N_11748);
and U19570 (N_19570,N_13666,N_12590);
or U19571 (N_19571,N_10764,N_10459);
nand U19572 (N_19572,N_13948,N_10737);
xnor U19573 (N_19573,N_12234,N_10597);
nand U19574 (N_19574,N_14909,N_13359);
or U19575 (N_19575,N_13960,N_12893);
xnor U19576 (N_19576,N_12817,N_10755);
and U19577 (N_19577,N_12509,N_11894);
nand U19578 (N_19578,N_11642,N_11388);
or U19579 (N_19579,N_13282,N_14187);
nor U19580 (N_19580,N_12892,N_13972);
nand U19581 (N_19581,N_10659,N_11813);
and U19582 (N_19582,N_10458,N_13551);
or U19583 (N_19583,N_12109,N_13664);
or U19584 (N_19584,N_13139,N_12047);
nor U19585 (N_19585,N_13034,N_13434);
and U19586 (N_19586,N_11096,N_12686);
nor U19587 (N_19587,N_10671,N_13698);
nor U19588 (N_19588,N_13986,N_12720);
and U19589 (N_19589,N_10514,N_14665);
nand U19590 (N_19590,N_10597,N_11866);
and U19591 (N_19591,N_12102,N_13428);
and U19592 (N_19592,N_11708,N_11019);
and U19593 (N_19593,N_14554,N_14510);
nand U19594 (N_19594,N_13333,N_13528);
xnor U19595 (N_19595,N_11899,N_11936);
and U19596 (N_19596,N_13970,N_14083);
nand U19597 (N_19597,N_14328,N_14832);
nor U19598 (N_19598,N_14138,N_12108);
and U19599 (N_19599,N_11110,N_11934);
nand U19600 (N_19600,N_14284,N_14618);
xor U19601 (N_19601,N_12989,N_11188);
nand U19602 (N_19602,N_12046,N_13496);
nand U19603 (N_19603,N_14507,N_12399);
and U19604 (N_19604,N_10409,N_12864);
nor U19605 (N_19605,N_10453,N_10675);
or U19606 (N_19606,N_10560,N_14310);
nor U19607 (N_19607,N_11147,N_14118);
and U19608 (N_19608,N_14583,N_14188);
nand U19609 (N_19609,N_12310,N_11025);
nand U19610 (N_19610,N_13852,N_11913);
nand U19611 (N_19611,N_13455,N_10084);
nand U19612 (N_19612,N_13975,N_14710);
nand U19613 (N_19613,N_10352,N_14916);
nand U19614 (N_19614,N_12756,N_11492);
and U19615 (N_19615,N_11470,N_14529);
nand U19616 (N_19616,N_11053,N_11713);
nor U19617 (N_19617,N_13559,N_11226);
nor U19618 (N_19618,N_14179,N_11562);
nand U19619 (N_19619,N_14529,N_13759);
and U19620 (N_19620,N_10103,N_12719);
nand U19621 (N_19621,N_14577,N_11723);
and U19622 (N_19622,N_14740,N_12880);
or U19623 (N_19623,N_14733,N_13457);
or U19624 (N_19624,N_14888,N_10219);
and U19625 (N_19625,N_10942,N_11190);
nand U19626 (N_19626,N_11107,N_14781);
and U19627 (N_19627,N_12134,N_10008);
or U19628 (N_19628,N_12257,N_10457);
nor U19629 (N_19629,N_13025,N_12395);
nor U19630 (N_19630,N_13631,N_12944);
nor U19631 (N_19631,N_13810,N_12412);
and U19632 (N_19632,N_12161,N_11229);
nand U19633 (N_19633,N_12570,N_10661);
or U19634 (N_19634,N_12964,N_14644);
nor U19635 (N_19635,N_11259,N_14672);
xnor U19636 (N_19636,N_14724,N_11280);
or U19637 (N_19637,N_11603,N_10168);
and U19638 (N_19638,N_12324,N_12823);
nor U19639 (N_19639,N_11549,N_14055);
and U19640 (N_19640,N_12846,N_12066);
or U19641 (N_19641,N_10685,N_11141);
and U19642 (N_19642,N_14663,N_11945);
nand U19643 (N_19643,N_13194,N_13048);
nor U19644 (N_19644,N_13029,N_12696);
xor U19645 (N_19645,N_10367,N_13376);
nor U19646 (N_19646,N_13688,N_13209);
nor U19647 (N_19647,N_10057,N_12068);
and U19648 (N_19648,N_12916,N_14936);
or U19649 (N_19649,N_12521,N_14749);
nand U19650 (N_19650,N_12680,N_13134);
nand U19651 (N_19651,N_12395,N_11839);
and U19652 (N_19652,N_10258,N_12298);
nor U19653 (N_19653,N_12682,N_14020);
nand U19654 (N_19654,N_13881,N_10288);
or U19655 (N_19655,N_14465,N_13861);
nand U19656 (N_19656,N_13349,N_11385);
nand U19657 (N_19657,N_10976,N_14434);
nor U19658 (N_19658,N_12903,N_13317);
or U19659 (N_19659,N_11170,N_11163);
nand U19660 (N_19660,N_12367,N_14486);
nand U19661 (N_19661,N_12519,N_10287);
nand U19662 (N_19662,N_12592,N_12470);
xor U19663 (N_19663,N_11004,N_13921);
or U19664 (N_19664,N_10247,N_14520);
nand U19665 (N_19665,N_11892,N_11733);
nor U19666 (N_19666,N_10536,N_12372);
or U19667 (N_19667,N_13369,N_13320);
or U19668 (N_19668,N_11435,N_13106);
nor U19669 (N_19669,N_10515,N_13965);
nand U19670 (N_19670,N_13709,N_12024);
nor U19671 (N_19671,N_11370,N_13535);
nand U19672 (N_19672,N_14565,N_14249);
nand U19673 (N_19673,N_12380,N_14030);
and U19674 (N_19674,N_12400,N_10733);
nand U19675 (N_19675,N_12945,N_14125);
and U19676 (N_19676,N_10924,N_11808);
nand U19677 (N_19677,N_14818,N_10703);
nand U19678 (N_19678,N_11116,N_14787);
nand U19679 (N_19679,N_10555,N_13916);
nor U19680 (N_19680,N_14900,N_12377);
nor U19681 (N_19681,N_14216,N_14882);
nand U19682 (N_19682,N_10701,N_12154);
or U19683 (N_19683,N_10959,N_11821);
nor U19684 (N_19684,N_11452,N_12592);
nand U19685 (N_19685,N_12549,N_11269);
or U19686 (N_19686,N_10760,N_10399);
nor U19687 (N_19687,N_12083,N_13016);
nand U19688 (N_19688,N_13682,N_11090);
nand U19689 (N_19689,N_12863,N_13717);
nand U19690 (N_19690,N_13644,N_12512);
nor U19691 (N_19691,N_14149,N_13598);
and U19692 (N_19692,N_11145,N_12197);
and U19693 (N_19693,N_14132,N_12120);
or U19694 (N_19694,N_14904,N_12476);
and U19695 (N_19695,N_10805,N_13933);
nor U19696 (N_19696,N_14040,N_10268);
and U19697 (N_19697,N_12724,N_13797);
xor U19698 (N_19698,N_11915,N_11206);
nor U19699 (N_19699,N_10029,N_10711);
nand U19700 (N_19700,N_12155,N_10820);
xnor U19701 (N_19701,N_13424,N_13382);
or U19702 (N_19702,N_10357,N_14598);
and U19703 (N_19703,N_12912,N_12648);
nand U19704 (N_19704,N_14794,N_13127);
nand U19705 (N_19705,N_14229,N_11400);
or U19706 (N_19706,N_14675,N_12389);
nor U19707 (N_19707,N_14330,N_11110);
or U19708 (N_19708,N_11447,N_12532);
or U19709 (N_19709,N_13832,N_14184);
nor U19710 (N_19710,N_14317,N_13810);
nor U19711 (N_19711,N_13414,N_11534);
xor U19712 (N_19712,N_11257,N_13624);
and U19713 (N_19713,N_11225,N_13851);
or U19714 (N_19714,N_12085,N_14392);
or U19715 (N_19715,N_12835,N_11529);
nand U19716 (N_19716,N_14325,N_14730);
or U19717 (N_19717,N_11385,N_13260);
and U19718 (N_19718,N_13101,N_13389);
and U19719 (N_19719,N_12855,N_10190);
or U19720 (N_19720,N_12833,N_13522);
and U19721 (N_19721,N_14656,N_14162);
and U19722 (N_19722,N_11536,N_10097);
or U19723 (N_19723,N_12985,N_14944);
nand U19724 (N_19724,N_14636,N_11945);
or U19725 (N_19725,N_13872,N_10849);
or U19726 (N_19726,N_10550,N_13324);
and U19727 (N_19727,N_11417,N_10838);
nand U19728 (N_19728,N_14403,N_11700);
and U19729 (N_19729,N_12259,N_13557);
nand U19730 (N_19730,N_11415,N_13951);
xnor U19731 (N_19731,N_10615,N_13385);
nor U19732 (N_19732,N_12079,N_13151);
or U19733 (N_19733,N_14303,N_14876);
or U19734 (N_19734,N_14134,N_13282);
xor U19735 (N_19735,N_13455,N_11015);
xnor U19736 (N_19736,N_14309,N_10133);
nor U19737 (N_19737,N_12235,N_12063);
nand U19738 (N_19738,N_14909,N_11932);
nand U19739 (N_19739,N_13195,N_11279);
and U19740 (N_19740,N_14540,N_12624);
or U19741 (N_19741,N_13447,N_11097);
nand U19742 (N_19742,N_13028,N_14809);
and U19743 (N_19743,N_13001,N_14778);
nand U19744 (N_19744,N_10485,N_11666);
and U19745 (N_19745,N_10599,N_12178);
xnor U19746 (N_19746,N_11766,N_13069);
nor U19747 (N_19747,N_14823,N_12997);
or U19748 (N_19748,N_12935,N_10757);
or U19749 (N_19749,N_11881,N_12702);
and U19750 (N_19750,N_10846,N_14575);
nor U19751 (N_19751,N_13961,N_12082);
nand U19752 (N_19752,N_11891,N_12302);
and U19753 (N_19753,N_13469,N_14890);
nor U19754 (N_19754,N_13852,N_13808);
or U19755 (N_19755,N_14659,N_11449);
nor U19756 (N_19756,N_14945,N_10538);
nor U19757 (N_19757,N_11620,N_11264);
nor U19758 (N_19758,N_12722,N_11872);
or U19759 (N_19759,N_13057,N_12717);
nand U19760 (N_19760,N_14937,N_12383);
nor U19761 (N_19761,N_10453,N_12550);
xnor U19762 (N_19762,N_11639,N_13337);
nand U19763 (N_19763,N_14950,N_12548);
or U19764 (N_19764,N_10790,N_12621);
or U19765 (N_19765,N_14130,N_13791);
nor U19766 (N_19766,N_11625,N_10414);
nand U19767 (N_19767,N_13277,N_11705);
or U19768 (N_19768,N_10188,N_14688);
nand U19769 (N_19769,N_11036,N_13379);
nor U19770 (N_19770,N_13745,N_14775);
nor U19771 (N_19771,N_13535,N_13709);
nor U19772 (N_19772,N_14841,N_13439);
and U19773 (N_19773,N_11205,N_10748);
nor U19774 (N_19774,N_12026,N_13527);
and U19775 (N_19775,N_14918,N_13589);
nor U19776 (N_19776,N_10907,N_12762);
nand U19777 (N_19777,N_14084,N_10524);
or U19778 (N_19778,N_14509,N_11468);
and U19779 (N_19779,N_12795,N_12687);
nand U19780 (N_19780,N_13887,N_11287);
and U19781 (N_19781,N_13386,N_10857);
and U19782 (N_19782,N_11581,N_11422);
and U19783 (N_19783,N_11391,N_11643);
nor U19784 (N_19784,N_12171,N_12997);
nor U19785 (N_19785,N_12075,N_10529);
or U19786 (N_19786,N_11313,N_11012);
xor U19787 (N_19787,N_14443,N_12131);
nor U19788 (N_19788,N_12902,N_13532);
xnor U19789 (N_19789,N_10608,N_14179);
and U19790 (N_19790,N_11537,N_14039);
or U19791 (N_19791,N_10856,N_11936);
nor U19792 (N_19792,N_14815,N_12580);
nand U19793 (N_19793,N_11471,N_13046);
or U19794 (N_19794,N_13854,N_12893);
or U19795 (N_19795,N_13509,N_11768);
and U19796 (N_19796,N_10323,N_13425);
nor U19797 (N_19797,N_10762,N_14941);
xnor U19798 (N_19798,N_11994,N_11806);
nand U19799 (N_19799,N_13138,N_12938);
and U19800 (N_19800,N_11533,N_13667);
nor U19801 (N_19801,N_11985,N_10070);
xor U19802 (N_19802,N_14558,N_10492);
and U19803 (N_19803,N_13172,N_13419);
nand U19804 (N_19804,N_10520,N_10206);
xnor U19805 (N_19805,N_10842,N_10596);
nor U19806 (N_19806,N_13438,N_10832);
or U19807 (N_19807,N_11191,N_14984);
or U19808 (N_19808,N_11839,N_14574);
and U19809 (N_19809,N_14313,N_11478);
nand U19810 (N_19810,N_10126,N_11954);
or U19811 (N_19811,N_12499,N_14643);
nor U19812 (N_19812,N_11643,N_10910);
nand U19813 (N_19813,N_14534,N_11532);
nand U19814 (N_19814,N_14238,N_13015);
or U19815 (N_19815,N_12849,N_10992);
nand U19816 (N_19816,N_11814,N_11401);
nand U19817 (N_19817,N_13148,N_12332);
xnor U19818 (N_19818,N_11908,N_12678);
nand U19819 (N_19819,N_13480,N_10868);
and U19820 (N_19820,N_14585,N_11711);
nand U19821 (N_19821,N_12551,N_14163);
nor U19822 (N_19822,N_12400,N_13952);
and U19823 (N_19823,N_14050,N_10004);
nand U19824 (N_19824,N_14023,N_14327);
nor U19825 (N_19825,N_14136,N_11173);
and U19826 (N_19826,N_13453,N_12760);
nor U19827 (N_19827,N_11896,N_14531);
nor U19828 (N_19828,N_10515,N_14142);
nand U19829 (N_19829,N_11382,N_14042);
nand U19830 (N_19830,N_12268,N_13126);
nand U19831 (N_19831,N_11879,N_10127);
or U19832 (N_19832,N_13689,N_11958);
nand U19833 (N_19833,N_14377,N_10608);
and U19834 (N_19834,N_10815,N_14104);
nor U19835 (N_19835,N_13497,N_13735);
nand U19836 (N_19836,N_13831,N_11905);
nor U19837 (N_19837,N_10173,N_14422);
nand U19838 (N_19838,N_13961,N_12009);
or U19839 (N_19839,N_14217,N_11299);
or U19840 (N_19840,N_13209,N_10535);
nand U19841 (N_19841,N_10643,N_12014);
or U19842 (N_19842,N_10089,N_10137);
and U19843 (N_19843,N_12291,N_13703);
nor U19844 (N_19844,N_12759,N_10714);
or U19845 (N_19845,N_14158,N_12704);
or U19846 (N_19846,N_10913,N_13649);
nor U19847 (N_19847,N_10905,N_12193);
nor U19848 (N_19848,N_12166,N_14354);
or U19849 (N_19849,N_11736,N_14286);
nand U19850 (N_19850,N_10039,N_12815);
and U19851 (N_19851,N_12282,N_14019);
or U19852 (N_19852,N_11411,N_10888);
nand U19853 (N_19853,N_14061,N_14819);
and U19854 (N_19854,N_10945,N_13171);
nand U19855 (N_19855,N_12460,N_11403);
and U19856 (N_19856,N_11942,N_12770);
nor U19857 (N_19857,N_12485,N_11310);
nor U19858 (N_19858,N_11862,N_10291);
nand U19859 (N_19859,N_13513,N_13509);
nand U19860 (N_19860,N_12482,N_11372);
xor U19861 (N_19861,N_13280,N_13014);
and U19862 (N_19862,N_11653,N_13653);
nor U19863 (N_19863,N_14209,N_10263);
xor U19864 (N_19864,N_14735,N_13775);
and U19865 (N_19865,N_11810,N_12485);
nor U19866 (N_19866,N_12694,N_13913);
and U19867 (N_19867,N_13053,N_14148);
and U19868 (N_19868,N_13264,N_14069);
nand U19869 (N_19869,N_12684,N_12048);
and U19870 (N_19870,N_10447,N_10022);
and U19871 (N_19871,N_11468,N_14148);
and U19872 (N_19872,N_12911,N_10071);
nor U19873 (N_19873,N_10667,N_13145);
or U19874 (N_19874,N_10452,N_10896);
or U19875 (N_19875,N_12714,N_12177);
nand U19876 (N_19876,N_13625,N_12677);
nor U19877 (N_19877,N_13772,N_10593);
nor U19878 (N_19878,N_12621,N_13768);
nor U19879 (N_19879,N_11122,N_13829);
xor U19880 (N_19880,N_11013,N_10637);
nor U19881 (N_19881,N_10019,N_11808);
and U19882 (N_19882,N_10433,N_11295);
nor U19883 (N_19883,N_14104,N_13539);
nor U19884 (N_19884,N_14185,N_12436);
and U19885 (N_19885,N_11984,N_13417);
nor U19886 (N_19886,N_12403,N_14573);
nor U19887 (N_19887,N_11851,N_11146);
xnor U19888 (N_19888,N_11638,N_10856);
or U19889 (N_19889,N_12934,N_13505);
or U19890 (N_19890,N_10320,N_14782);
and U19891 (N_19891,N_10127,N_12127);
and U19892 (N_19892,N_13437,N_12491);
nor U19893 (N_19893,N_10680,N_10734);
or U19894 (N_19894,N_12656,N_13639);
or U19895 (N_19895,N_12765,N_13835);
or U19896 (N_19896,N_11956,N_10240);
and U19897 (N_19897,N_10279,N_12736);
nand U19898 (N_19898,N_12265,N_13131);
xor U19899 (N_19899,N_12917,N_12465);
or U19900 (N_19900,N_14101,N_14097);
nor U19901 (N_19901,N_12727,N_12505);
and U19902 (N_19902,N_12508,N_14803);
and U19903 (N_19903,N_10742,N_10021);
or U19904 (N_19904,N_11937,N_11504);
nand U19905 (N_19905,N_11248,N_11576);
nor U19906 (N_19906,N_12766,N_13167);
or U19907 (N_19907,N_14380,N_10683);
or U19908 (N_19908,N_10828,N_11778);
xor U19909 (N_19909,N_13230,N_13635);
and U19910 (N_19910,N_10117,N_14850);
or U19911 (N_19911,N_12334,N_13903);
nand U19912 (N_19912,N_14190,N_13240);
or U19913 (N_19913,N_13750,N_12278);
xor U19914 (N_19914,N_11842,N_13486);
nand U19915 (N_19915,N_11312,N_10106);
or U19916 (N_19916,N_11615,N_11336);
nor U19917 (N_19917,N_14953,N_10779);
xnor U19918 (N_19918,N_12445,N_11712);
or U19919 (N_19919,N_13928,N_10501);
nand U19920 (N_19920,N_14181,N_12344);
nand U19921 (N_19921,N_10273,N_14795);
or U19922 (N_19922,N_12108,N_14800);
and U19923 (N_19923,N_13042,N_10055);
or U19924 (N_19924,N_10442,N_14478);
nor U19925 (N_19925,N_12726,N_12429);
or U19926 (N_19926,N_12929,N_14768);
nand U19927 (N_19927,N_10986,N_13135);
nor U19928 (N_19928,N_12650,N_10299);
and U19929 (N_19929,N_14329,N_14374);
nand U19930 (N_19930,N_14982,N_10444);
nand U19931 (N_19931,N_13764,N_13133);
xnor U19932 (N_19932,N_13261,N_10641);
xnor U19933 (N_19933,N_13159,N_12970);
or U19934 (N_19934,N_10674,N_14368);
xnor U19935 (N_19935,N_12775,N_14512);
and U19936 (N_19936,N_11581,N_11505);
nand U19937 (N_19937,N_11963,N_13045);
and U19938 (N_19938,N_11495,N_11785);
nor U19939 (N_19939,N_13326,N_10573);
nor U19940 (N_19940,N_11218,N_11160);
or U19941 (N_19941,N_13018,N_11171);
and U19942 (N_19942,N_10504,N_14017);
and U19943 (N_19943,N_12018,N_12365);
xnor U19944 (N_19944,N_12932,N_13776);
or U19945 (N_19945,N_10921,N_10896);
nor U19946 (N_19946,N_10198,N_11376);
or U19947 (N_19947,N_13628,N_13296);
nand U19948 (N_19948,N_12647,N_13666);
or U19949 (N_19949,N_12966,N_11318);
nor U19950 (N_19950,N_14067,N_14515);
nand U19951 (N_19951,N_11651,N_11130);
and U19952 (N_19952,N_13907,N_14225);
nor U19953 (N_19953,N_13933,N_10395);
nor U19954 (N_19954,N_10573,N_12425);
nor U19955 (N_19955,N_14751,N_11571);
or U19956 (N_19956,N_10028,N_13889);
and U19957 (N_19957,N_13503,N_14018);
nand U19958 (N_19958,N_10821,N_13161);
nor U19959 (N_19959,N_13441,N_10603);
xor U19960 (N_19960,N_12102,N_12106);
nand U19961 (N_19961,N_14816,N_12484);
nor U19962 (N_19962,N_11525,N_10751);
and U19963 (N_19963,N_12371,N_12801);
and U19964 (N_19964,N_11385,N_13273);
xor U19965 (N_19965,N_11564,N_14320);
nor U19966 (N_19966,N_12520,N_14764);
and U19967 (N_19967,N_14936,N_14028);
xnor U19968 (N_19968,N_11255,N_11041);
and U19969 (N_19969,N_12432,N_10410);
and U19970 (N_19970,N_14641,N_12145);
nand U19971 (N_19971,N_11534,N_11952);
nand U19972 (N_19972,N_13906,N_10414);
or U19973 (N_19973,N_13205,N_12744);
or U19974 (N_19974,N_11482,N_11228);
or U19975 (N_19975,N_11920,N_13331);
nor U19976 (N_19976,N_12235,N_10504);
nor U19977 (N_19977,N_12551,N_11754);
nand U19978 (N_19978,N_11982,N_11612);
nor U19979 (N_19979,N_13716,N_12022);
or U19980 (N_19980,N_10104,N_14295);
and U19981 (N_19981,N_10417,N_11774);
nor U19982 (N_19982,N_12165,N_13574);
xor U19983 (N_19983,N_12321,N_14399);
nand U19984 (N_19984,N_14487,N_13361);
nor U19985 (N_19985,N_14553,N_11349);
and U19986 (N_19986,N_14087,N_11797);
nand U19987 (N_19987,N_11399,N_12066);
nand U19988 (N_19988,N_14338,N_12359);
or U19989 (N_19989,N_11069,N_12271);
xor U19990 (N_19990,N_10390,N_10839);
nand U19991 (N_19991,N_11761,N_11051);
and U19992 (N_19992,N_11102,N_10780);
nor U19993 (N_19993,N_13910,N_11925);
and U19994 (N_19994,N_11353,N_12211);
xnor U19995 (N_19995,N_14517,N_14198);
nand U19996 (N_19996,N_10301,N_13316);
and U19997 (N_19997,N_13869,N_10223);
and U19998 (N_19998,N_11256,N_10502);
and U19999 (N_19999,N_11673,N_13770);
and UO_0 (O_0,N_17940,N_17616);
and UO_1 (O_1,N_19334,N_16981);
xnor UO_2 (O_2,N_19883,N_17517);
or UO_3 (O_3,N_16469,N_15311);
and UO_4 (O_4,N_19267,N_18382);
or UO_5 (O_5,N_18089,N_19551);
nand UO_6 (O_6,N_19656,N_19878);
nand UO_7 (O_7,N_15068,N_16008);
xnor UO_8 (O_8,N_17835,N_18341);
nor UO_9 (O_9,N_16644,N_19349);
nand UO_10 (O_10,N_17992,N_16078);
nor UO_11 (O_11,N_18779,N_15574);
nor UO_12 (O_12,N_16444,N_19830);
or UO_13 (O_13,N_16255,N_19645);
nand UO_14 (O_14,N_19232,N_16794);
nand UO_15 (O_15,N_19062,N_16711);
or UO_16 (O_16,N_16997,N_16335);
and UO_17 (O_17,N_17243,N_15290);
nor UO_18 (O_18,N_18570,N_17503);
xnor UO_19 (O_19,N_18688,N_18032);
and UO_20 (O_20,N_17312,N_16562);
or UO_21 (O_21,N_16724,N_15751);
nand UO_22 (O_22,N_18073,N_15828);
xor UO_23 (O_23,N_19189,N_15930);
or UO_24 (O_24,N_15050,N_17552);
nor UO_25 (O_25,N_16945,N_18223);
nor UO_26 (O_26,N_16486,N_18886);
nand UO_27 (O_27,N_18762,N_15743);
nand UO_28 (O_28,N_15782,N_17620);
and UO_29 (O_29,N_18707,N_15062);
nor UO_30 (O_30,N_19407,N_16654);
nor UO_31 (O_31,N_15647,N_17608);
nand UO_32 (O_32,N_16870,N_18631);
and UO_33 (O_33,N_15665,N_18623);
or UO_34 (O_34,N_17177,N_19723);
or UO_35 (O_35,N_15307,N_17640);
and UO_36 (O_36,N_19041,N_17626);
nand UO_37 (O_37,N_18397,N_17295);
and UO_38 (O_38,N_17353,N_18460);
or UO_39 (O_39,N_16509,N_15882);
and UO_40 (O_40,N_15366,N_17642);
and UO_41 (O_41,N_18479,N_19499);
and UO_42 (O_42,N_18435,N_17595);
nor UO_43 (O_43,N_16854,N_18617);
xor UO_44 (O_44,N_16390,N_18517);
nand UO_45 (O_45,N_16754,N_15224);
or UO_46 (O_46,N_16225,N_18437);
nor UO_47 (O_47,N_19184,N_18713);
nor UO_48 (O_48,N_19691,N_18967);
or UO_49 (O_49,N_19966,N_17046);
nand UO_50 (O_50,N_15429,N_19084);
xnor UO_51 (O_51,N_18134,N_15187);
or UO_52 (O_52,N_15523,N_17514);
nand UO_53 (O_53,N_15262,N_18512);
nand UO_54 (O_54,N_16044,N_17559);
and UO_55 (O_55,N_18219,N_19101);
or UO_56 (O_56,N_18061,N_19209);
nand UO_57 (O_57,N_18399,N_17403);
and UO_58 (O_58,N_19763,N_18589);
xnor UO_59 (O_59,N_15084,N_19671);
nand UO_60 (O_60,N_15735,N_18645);
and UO_61 (O_61,N_17737,N_15291);
or UO_62 (O_62,N_15431,N_19177);
nand UO_63 (O_63,N_18354,N_15915);
nand UO_64 (O_64,N_17275,N_18173);
nor UO_65 (O_65,N_16687,N_16529);
nand UO_66 (O_66,N_19976,N_16580);
nor UO_67 (O_67,N_18567,N_17605);
nor UO_68 (O_68,N_19556,N_17763);
and UO_69 (O_69,N_18454,N_18198);
nor UO_70 (O_70,N_17561,N_18402);
and UO_71 (O_71,N_16143,N_19716);
nor UO_72 (O_72,N_19555,N_19153);
nor UO_73 (O_73,N_15544,N_15428);
nand UO_74 (O_74,N_18192,N_15340);
and UO_75 (O_75,N_18357,N_16114);
nor UO_76 (O_76,N_18318,N_16670);
or UO_77 (O_77,N_19954,N_17250);
nand UO_78 (O_78,N_17369,N_18823);
xnor UO_79 (O_79,N_17970,N_19051);
nor UO_80 (O_80,N_19438,N_19481);
xnor UO_81 (O_81,N_19767,N_19627);
and UO_82 (O_82,N_15280,N_16310);
nand UO_83 (O_83,N_17844,N_16136);
nor UO_84 (O_84,N_16911,N_15095);
or UO_85 (O_85,N_15259,N_18736);
or UO_86 (O_86,N_17804,N_15323);
or UO_87 (O_87,N_15245,N_19038);
nand UO_88 (O_88,N_17743,N_18153);
nand UO_89 (O_89,N_15957,N_16278);
and UO_90 (O_90,N_16680,N_15802);
and UO_91 (O_91,N_16744,N_15070);
or UO_92 (O_92,N_15912,N_17210);
nand UO_93 (O_93,N_16702,N_15637);
and UO_94 (O_94,N_18747,N_16435);
nand UO_95 (O_95,N_17102,N_15922);
and UO_96 (O_96,N_15473,N_17478);
nor UO_97 (O_97,N_15391,N_15766);
nand UO_98 (O_98,N_15266,N_15639);
nor UO_99 (O_99,N_19251,N_15174);
or UO_100 (O_100,N_16084,N_15347);
or UO_101 (O_101,N_17493,N_18102);
or UO_102 (O_102,N_15142,N_18822);
and UO_103 (O_103,N_16919,N_16589);
nor UO_104 (O_104,N_16466,N_18758);
or UO_105 (O_105,N_15332,N_16100);
and UO_106 (O_106,N_18473,N_15125);
or UO_107 (O_107,N_18542,N_17044);
nand UO_108 (O_108,N_19922,N_19310);
nand UO_109 (O_109,N_19701,N_18244);
nand UO_110 (O_110,N_17445,N_19930);
or UO_111 (O_111,N_17920,N_15555);
or UO_112 (O_112,N_18915,N_17239);
xor UO_113 (O_113,N_19414,N_15533);
xnor UO_114 (O_114,N_18983,N_19936);
nor UO_115 (O_115,N_18828,N_17834);
nand UO_116 (O_116,N_16260,N_19539);
nand UO_117 (O_117,N_16208,N_19875);
and UO_118 (O_118,N_18656,N_17346);
nand UO_119 (O_119,N_18597,N_15459);
or UO_120 (O_120,N_16629,N_19468);
or UO_121 (O_121,N_18576,N_18651);
nand UO_122 (O_122,N_16398,N_18378);
or UO_123 (O_123,N_18522,N_15680);
or UO_124 (O_124,N_18520,N_19149);
nor UO_125 (O_125,N_17717,N_17810);
nand UO_126 (O_126,N_18844,N_19262);
nor UO_127 (O_127,N_19650,N_17913);
or UO_128 (O_128,N_18963,N_16844);
xor UO_129 (O_129,N_15385,N_19092);
or UO_130 (O_130,N_17814,N_16986);
and UO_131 (O_131,N_18529,N_16798);
and UO_132 (O_132,N_19117,N_18921);
nor UO_133 (O_133,N_15622,N_15502);
nor UO_134 (O_134,N_17785,N_19751);
nand UO_135 (O_135,N_19429,N_16358);
and UO_136 (O_136,N_16170,N_17340);
and UO_137 (O_137,N_19885,N_17683);
or UO_138 (O_138,N_18776,N_19367);
nor UO_139 (O_139,N_18857,N_15662);
and UO_140 (O_140,N_15993,N_19781);
nor UO_141 (O_141,N_19896,N_15052);
and UO_142 (O_142,N_15963,N_19582);
xnor UO_143 (O_143,N_18184,N_18824);
or UO_144 (O_144,N_17002,N_15832);
and UO_145 (O_145,N_16635,N_19554);
xnor UO_146 (O_146,N_19055,N_17131);
nor UO_147 (O_147,N_19252,N_18128);
and UO_148 (O_148,N_18701,N_16004);
and UO_149 (O_149,N_18429,N_19379);
nand UO_150 (O_150,N_18668,N_16735);
nand UO_151 (O_151,N_19508,N_17342);
nor UO_152 (O_152,N_15001,N_17427);
or UO_153 (O_153,N_18025,N_16683);
nor UO_154 (O_154,N_17741,N_17720);
nand UO_155 (O_155,N_16340,N_19743);
nand UO_156 (O_156,N_19591,N_15975);
or UO_157 (O_157,N_17057,N_17454);
nor UO_158 (O_158,N_19257,N_15867);
and UO_159 (O_159,N_16734,N_18260);
nor UO_160 (O_160,N_17974,N_19151);
or UO_161 (O_161,N_15506,N_16952);
xnor UO_162 (O_162,N_18271,N_18005);
or UO_163 (O_163,N_16209,N_15475);
nor UO_164 (O_164,N_16576,N_17227);
nand UO_165 (O_165,N_15976,N_18481);
nand UO_166 (O_166,N_18505,N_17512);
xor UO_167 (O_167,N_17196,N_18979);
or UO_168 (O_168,N_16824,N_17412);
nor UO_169 (O_169,N_17022,N_19576);
and UO_170 (O_170,N_17927,N_17672);
or UO_171 (O_171,N_15615,N_16662);
nor UO_172 (O_172,N_15518,N_18948);
or UO_173 (O_173,N_17694,N_15586);
nand UO_174 (O_174,N_19984,N_18974);
nand UO_175 (O_175,N_15282,N_16324);
nor UO_176 (O_176,N_19827,N_16174);
nor UO_177 (O_177,N_17055,N_18328);
and UO_178 (O_178,N_15914,N_18230);
or UO_179 (O_179,N_16941,N_15191);
nor UO_180 (O_180,N_19791,N_19190);
or UO_181 (O_181,N_15626,N_16133);
and UO_182 (O_182,N_16611,N_18735);
and UO_183 (O_183,N_18262,N_19597);
or UO_184 (O_184,N_16508,N_19406);
nand UO_185 (O_185,N_19297,N_15893);
and UO_186 (O_186,N_18106,N_15447);
nor UO_187 (O_187,N_18289,N_16428);
nor UO_188 (O_188,N_18063,N_18780);
nor UO_189 (O_189,N_18482,N_15433);
nand UO_190 (O_190,N_16312,N_18165);
and UO_191 (O_191,N_18581,N_16989);
nand UO_192 (O_192,N_18761,N_19536);
nand UO_193 (O_193,N_18075,N_17398);
or UO_194 (O_194,N_15685,N_15595);
or UO_195 (O_195,N_18253,N_15945);
nor UO_196 (O_196,N_19320,N_15166);
nor UO_197 (O_197,N_16139,N_19534);
nor UO_198 (O_198,N_15772,N_15926);
nor UO_199 (O_199,N_18453,N_19321);
nor UO_200 (O_200,N_19660,N_16007);
or UO_201 (O_201,N_16916,N_19123);
or UO_202 (O_202,N_16883,N_15721);
nor UO_203 (O_203,N_16606,N_15997);
or UO_204 (O_204,N_17719,N_15846);
or UO_205 (O_205,N_16054,N_18124);
nor UO_206 (O_206,N_15939,N_17952);
nor UO_207 (O_207,N_19887,N_16763);
or UO_208 (O_208,N_19509,N_17891);
and UO_209 (O_209,N_15512,N_17021);
and UO_210 (O_210,N_17315,N_16453);
nor UO_211 (O_211,N_15919,N_15033);
nor UO_212 (O_212,N_18784,N_17726);
and UO_213 (O_213,N_19754,N_19129);
nand UO_214 (O_214,N_17484,N_16210);
and UO_215 (O_215,N_18572,N_19090);
nand UO_216 (O_216,N_19580,N_15493);
nor UO_217 (O_217,N_15702,N_18026);
or UO_218 (O_218,N_18640,N_18555);
or UO_219 (O_219,N_19500,N_19135);
and UO_220 (O_220,N_18694,N_19083);
nor UO_221 (O_221,N_16727,N_19156);
and UO_222 (O_222,N_18282,N_17482);
or UO_223 (O_223,N_17975,N_18462);
and UO_224 (O_224,N_16481,N_17266);
and UO_225 (O_225,N_16692,N_17795);
nand UO_226 (O_226,N_17467,N_16715);
nand UO_227 (O_227,N_15202,N_16623);
nand UO_228 (O_228,N_17531,N_16033);
and UO_229 (O_229,N_15749,N_17040);
xnor UO_230 (O_230,N_15289,N_15906);
xor UO_231 (O_231,N_19002,N_16161);
or UO_232 (O_232,N_16781,N_15139);
nor UO_233 (O_233,N_16013,N_18418);
and UO_234 (O_234,N_19000,N_16056);
and UO_235 (O_235,N_17453,N_17845);
nand UO_236 (O_236,N_16974,N_19547);
nand UO_237 (O_237,N_19617,N_16821);
and UO_238 (O_238,N_16516,N_16112);
or UO_239 (O_239,N_15313,N_17762);
or UO_240 (O_240,N_17780,N_18962);
and UO_241 (O_241,N_19787,N_16863);
nor UO_242 (O_242,N_17915,N_15235);
or UO_243 (O_243,N_15596,N_17732);
nand UO_244 (O_244,N_16321,N_17392);
nand UO_245 (O_245,N_16944,N_16395);
and UO_246 (O_246,N_18486,N_16757);
or UO_247 (O_247,N_18647,N_18493);
nor UO_248 (O_248,N_19488,N_19994);
and UO_249 (O_249,N_19828,N_19684);
nor UO_250 (O_250,N_19946,N_18087);
nor UO_251 (O_251,N_19565,N_17233);
xnor UO_252 (O_252,N_19586,N_15520);
nor UO_253 (O_253,N_16904,N_17166);
or UO_254 (O_254,N_17964,N_18883);
or UO_255 (O_255,N_18930,N_18286);
nor UO_256 (O_256,N_16837,N_16705);
nand UO_257 (O_257,N_19250,N_15481);
nand UO_258 (O_258,N_15031,N_19624);
or UO_259 (O_259,N_17284,N_15826);
xor UO_260 (O_260,N_18444,N_17337);
or UO_261 (O_261,N_19440,N_15989);
and UO_262 (O_262,N_15781,N_15465);
nor UO_263 (O_263,N_19360,N_17142);
or UO_264 (O_264,N_17201,N_17064);
nor UO_265 (O_265,N_19799,N_15264);
xor UO_266 (O_266,N_15342,N_16593);
and UO_267 (O_267,N_15184,N_19464);
nand UO_268 (O_268,N_17189,N_19545);
or UO_269 (O_269,N_17259,N_15793);
and UO_270 (O_270,N_15078,N_19940);
nand UO_271 (O_271,N_19019,N_17494);
nand UO_272 (O_272,N_19643,N_16094);
xor UO_273 (O_273,N_19694,N_16771);
or UO_274 (O_274,N_19079,N_18778);
nand UO_275 (O_275,N_17747,N_18122);
nand UO_276 (O_276,N_17045,N_16261);
nor UO_277 (O_277,N_16559,N_15617);
nor UO_278 (O_278,N_19958,N_19895);
nor UO_279 (O_279,N_15953,N_18491);
nand UO_280 (O_280,N_17148,N_17215);
and UO_281 (O_281,N_18600,N_17322);
nand UO_282 (O_282,N_15729,N_16686);
nand UO_283 (O_283,N_19371,N_16828);
nor UO_284 (O_284,N_17410,N_16567);
or UO_285 (O_285,N_19093,N_19127);
nor UO_286 (O_286,N_15122,N_16943);
nor UO_287 (O_287,N_16990,N_15408);
nand UO_288 (O_288,N_17678,N_16785);
or UO_289 (O_289,N_18239,N_17837);
nand UO_290 (O_290,N_19696,N_19498);
and UO_291 (O_291,N_17367,N_15686);
nor UO_292 (O_292,N_15949,N_17422);
and UO_293 (O_293,N_15208,N_18312);
xnor UO_294 (O_294,N_15761,N_17783);
or UO_295 (O_295,N_19526,N_17397);
xnor UO_296 (O_296,N_17596,N_19630);
nor UO_297 (O_297,N_19221,N_17130);
xnor UO_298 (O_298,N_17649,N_18194);
and UO_299 (O_299,N_19034,N_18228);
and UO_300 (O_300,N_17223,N_17697);
xor UO_301 (O_301,N_17869,N_17666);
or UO_302 (O_302,N_18249,N_16353);
nand UO_303 (O_303,N_19622,N_16368);
nand UO_304 (O_304,N_19842,N_19215);
or UO_305 (O_305,N_15434,N_18841);
or UO_306 (O_306,N_19663,N_16582);
or UO_307 (O_307,N_15209,N_15500);
xnor UO_308 (O_308,N_19013,N_17555);
xor UO_309 (O_309,N_19385,N_17262);
and UO_310 (O_310,N_17008,N_17286);
nor UO_311 (O_311,N_18415,N_16632);
xnor UO_312 (O_312,N_16924,N_16167);
nor UO_313 (O_313,N_18665,N_18675);
xor UO_314 (O_314,N_16826,N_18654);
nor UO_315 (O_315,N_17860,N_15581);
and UO_316 (O_316,N_19255,N_16528);
or UO_317 (O_317,N_16247,N_15795);
nand UO_318 (O_318,N_18234,N_18995);
nand UO_319 (O_319,N_17129,N_15551);
nand UO_320 (O_320,N_17742,N_18528);
xor UO_321 (O_321,N_15442,N_15328);
or UO_322 (O_322,N_19537,N_18786);
nand UO_323 (O_323,N_19324,N_15886);
or UO_324 (O_324,N_18386,N_19131);
nor UO_325 (O_325,N_15946,N_19424);
and UO_326 (O_326,N_15638,N_19581);
and UO_327 (O_327,N_17598,N_15252);
or UO_328 (O_328,N_19693,N_17734);
and UO_329 (O_329,N_18033,N_19672);
and UO_330 (O_330,N_19141,N_16245);
xnor UO_331 (O_331,N_16690,N_16908);
and UO_332 (O_332,N_17281,N_19943);
nand UO_333 (O_333,N_19686,N_16476);
and UO_334 (O_334,N_15578,N_18568);
and UO_335 (O_335,N_16688,N_19095);
nor UO_336 (O_336,N_15348,N_16577);
nor UO_337 (O_337,N_15297,N_19318);
nand UO_338 (O_338,N_18850,N_17409);
nor UO_339 (O_339,N_18970,N_19520);
nand UO_340 (O_340,N_18351,N_19031);
nand UO_341 (O_341,N_19336,N_18052);
or UO_342 (O_342,N_19486,N_19973);
and UO_343 (O_343,N_15267,N_17871);
or UO_344 (O_344,N_18989,N_19241);
or UO_345 (O_345,N_17787,N_18206);
and UO_346 (O_346,N_16759,N_16263);
nor UO_347 (O_347,N_19351,N_19768);
xor UO_348 (O_348,N_16953,N_15404);
and UO_349 (O_349,N_15199,N_18584);
and UO_350 (O_350,N_19978,N_15416);
and UO_351 (O_351,N_19546,N_19821);
or UO_352 (O_352,N_16901,N_17520);
xor UO_353 (O_353,N_19575,N_15361);
nand UO_354 (O_354,N_17232,N_16274);
nor UO_355 (O_355,N_15383,N_16907);
nor UO_356 (O_356,N_15146,N_17961);
nand UO_357 (O_357,N_16909,N_17693);
or UO_358 (O_358,N_16572,N_15195);
and UO_359 (O_359,N_17160,N_18416);
or UO_360 (O_360,N_18202,N_19201);
nand UO_361 (O_361,N_16959,N_16218);
or UO_362 (O_362,N_18464,N_15315);
nor UO_363 (O_363,N_16352,N_19569);
and UO_364 (O_364,N_19989,N_15986);
nor UO_365 (O_365,N_15709,N_18916);
and UO_366 (O_366,N_16465,N_19086);
or UO_367 (O_367,N_17765,N_17803);
nor UO_368 (O_368,N_19132,N_16511);
nand UO_369 (O_369,N_18035,N_18250);
nor UO_370 (O_370,N_19303,N_17067);
and UO_371 (O_371,N_16490,N_18123);
or UO_372 (O_372,N_15938,N_17931);
nand UO_373 (O_373,N_19441,N_16602);
nor UO_374 (O_374,N_19606,N_15454);
nand UO_375 (O_375,N_15263,N_16085);
nand UO_376 (O_376,N_17035,N_16362);
nand UO_377 (O_377,N_18363,N_15403);
nand UO_378 (O_378,N_18489,N_19834);
or UO_379 (O_379,N_19449,N_18737);
nand UO_380 (O_380,N_15696,N_18468);
nor UO_381 (O_381,N_15030,N_19502);
or UO_382 (O_382,N_15367,N_15856);
nor UO_383 (O_383,N_19926,N_15636);
nor UO_384 (O_384,N_16720,N_17754);
nand UO_385 (O_385,N_18217,N_17428);
or UO_386 (O_386,N_17466,N_16969);
and UO_387 (O_387,N_17908,N_19489);
nand UO_388 (O_388,N_16913,N_15994);
or UO_389 (O_389,N_19792,N_17526);
and UO_390 (O_390,N_17336,N_18405);
xor UO_391 (O_391,N_15731,N_18065);
xor UO_392 (O_392,N_16808,N_16429);
and UO_393 (O_393,N_15104,N_15422);
nand UO_394 (O_394,N_17856,N_15837);
or UO_395 (O_395,N_15251,N_18596);
and UO_396 (O_396,N_18527,N_18703);
or UO_397 (O_397,N_15387,N_17280);
and UO_398 (O_398,N_19841,N_15485);
nor UO_399 (O_399,N_18296,N_18047);
nand UO_400 (O_400,N_19463,N_15546);
nor UO_401 (O_401,N_15974,N_17193);
nor UO_402 (O_402,N_18885,N_19124);
nand UO_403 (O_403,N_18254,N_18067);
nand UO_404 (O_404,N_18988,N_15655);
nor UO_405 (O_405,N_17135,N_18679);
or UO_406 (O_406,N_19292,N_16115);
nor UO_407 (O_407,N_15777,N_16823);
nand UO_408 (O_408,N_19274,N_19317);
nor UO_409 (O_409,N_18678,N_18972);
nand UO_410 (O_410,N_15679,N_17098);
nor UO_411 (O_411,N_19725,N_15330);
nor UO_412 (O_412,N_19746,N_19413);
nand UO_413 (O_413,N_17247,N_17735);
or UO_414 (O_414,N_15003,N_17388);
and UO_415 (O_415,N_17440,N_18705);
or UO_416 (O_416,N_16045,N_15634);
nand UO_417 (O_417,N_16416,N_18251);
or UO_418 (O_418,N_19507,N_18059);
or UO_419 (O_419,N_17536,N_17060);
nor UO_420 (O_420,N_15232,N_17585);
nor UO_421 (O_421,N_19572,N_19923);
and UO_422 (O_422,N_19742,N_16202);
and UO_423 (O_423,N_18307,N_16503);
or UO_424 (O_424,N_18634,N_17211);
nor UO_425 (O_425,N_15650,N_19103);
or UO_426 (O_426,N_18370,N_18212);
and UO_427 (O_427,N_19295,N_16548);
nand UO_428 (O_428,N_15868,N_18537);
nor UO_429 (O_429,N_17544,N_18441);
or UO_430 (O_430,N_19246,N_15354);
or UO_431 (O_431,N_19036,N_16081);
nand UO_432 (O_432,N_18361,N_16608);
or UO_433 (O_433,N_18672,N_16520);
nand UO_434 (O_434,N_15539,N_18827);
or UO_435 (O_435,N_17190,N_17857);
or UO_436 (O_436,N_19296,N_17907);
and UO_437 (O_437,N_15640,N_16439);
or UO_438 (O_438,N_18721,N_18870);
or UO_439 (O_439,N_19427,N_18507);
nor UO_440 (O_440,N_18290,N_17725);
or UO_441 (O_441,N_15833,N_18193);
and UO_442 (O_442,N_16873,N_17411);
or UO_443 (O_443,N_18743,N_15942);
xor UO_444 (O_444,N_16935,N_17235);
or UO_445 (O_445,N_17662,N_18613);
xor UO_446 (O_446,N_16965,N_16016);
and UO_447 (O_447,N_16841,N_18265);
and UO_448 (O_448,N_15630,N_17446);
nand UO_449 (O_449,N_16474,N_15362);
or UO_450 (O_450,N_16545,N_16658);
nor UO_451 (O_451,N_19106,N_16915);
nand UO_452 (O_452,N_17968,N_19788);
and UO_453 (O_453,N_18037,N_15478);
or UO_454 (O_454,N_15241,N_16751);
and UO_455 (O_455,N_16265,N_19155);
or UO_456 (O_456,N_16665,N_18904);
nand UO_457 (O_457,N_18174,N_16641);
and UO_458 (O_458,N_18582,N_16614);
xor UO_459 (O_459,N_18657,N_17489);
or UO_460 (O_460,N_19361,N_18845);
or UO_461 (O_461,N_19260,N_18285);
nand UO_462 (O_462,N_19247,N_19237);
nor UO_463 (O_463,N_19453,N_19941);
or UO_464 (O_464,N_18179,N_17248);
nor UO_465 (O_465,N_17444,N_17056);
or UO_466 (O_466,N_15716,N_16048);
nand UO_467 (O_467,N_16153,N_15300);
nand UO_468 (O_468,N_18946,N_16375);
nand UO_469 (O_469,N_16049,N_19717);
and UO_470 (O_470,N_19678,N_18105);
nor UO_471 (O_471,N_17301,N_16296);
nor UO_472 (O_472,N_18628,N_16027);
nor UO_473 (O_473,N_15979,N_16615);
and UO_474 (O_474,N_15453,N_16541);
or UO_475 (O_475,N_15444,N_19212);
nor UO_476 (O_476,N_18986,N_19474);
or UO_477 (O_477,N_15746,N_15564);
nor UO_478 (O_478,N_19187,N_17958);
nor UO_479 (O_479,N_15498,N_16640);
nand UO_480 (O_480,N_19170,N_16728);
nor UO_481 (O_481,N_19897,N_16515);
or UO_482 (O_482,N_17178,N_19955);
nor UO_483 (O_483,N_15722,N_17217);
or UO_484 (O_484,N_15689,N_15148);
and UO_485 (O_485,N_17420,N_18711);
xnor UO_486 (O_486,N_17938,N_18120);
nand UO_487 (O_487,N_17425,N_16458);
nor UO_488 (O_488,N_16918,N_16594);
or UO_489 (O_489,N_18064,N_19601);
nor UO_490 (O_490,N_16586,N_17847);
nor UO_491 (O_491,N_15284,N_19409);
xor UO_492 (O_492,N_15043,N_16792);
nor UO_493 (O_493,N_17206,N_16832);
nand UO_494 (O_494,N_17898,N_17457);
nor UO_495 (O_495,N_15278,N_19710);
or UO_496 (O_496,N_18697,N_16464);
xor UO_497 (O_497,N_16988,N_19739);
xnor UO_498 (O_498,N_19396,N_18578);
and UO_499 (O_499,N_16427,N_19181);
nor UO_500 (O_500,N_17221,N_17358);
nand UO_501 (O_501,N_17363,N_18150);
or UO_502 (O_502,N_16730,N_15014);
nand UO_503 (O_503,N_15071,N_15847);
nor UO_504 (O_504,N_18203,N_15244);
nand UO_505 (O_505,N_19053,N_19313);
nor UO_506 (O_506,N_18573,N_17488);
nor UO_507 (O_507,N_18792,N_16180);
nand UO_508 (O_508,N_19425,N_17667);
or UO_509 (O_509,N_15302,N_19762);
or UO_510 (O_510,N_16955,N_16206);
or UO_511 (O_511,N_16886,N_16342);
or UO_512 (O_512,N_19431,N_19049);
nor UO_513 (O_513,N_18958,N_15247);
or UO_514 (O_514,N_15150,N_19148);
nor UO_515 (O_515,N_19910,N_17459);
or UO_516 (O_516,N_18204,N_17876);
nand UO_517 (O_517,N_19230,N_15704);
or UO_518 (O_518,N_19778,N_16479);
nand UO_519 (O_519,N_19992,N_15117);
and UO_520 (O_520,N_19348,N_17923);
nand UO_521 (O_521,N_16963,N_17897);
and UO_522 (O_522,N_17853,N_18896);
or UO_523 (O_523,N_15389,N_18135);
nor UO_524 (O_524,N_19609,N_15301);
or UO_525 (O_525,N_16329,N_17539);
or UO_526 (O_526,N_16169,N_16159);
or UO_527 (O_527,N_19902,N_17759);
xnor UO_528 (O_528,N_15299,N_17345);
xnor UO_529 (O_529,N_17019,N_16491);
nor UO_530 (O_530,N_16099,N_17945);
nand UO_531 (O_531,N_16147,N_18220);
and UO_532 (O_532,N_15272,N_16304);
or UO_533 (O_533,N_15483,N_15576);
xnor UO_534 (O_534,N_17347,N_16947);
nor UO_535 (O_535,N_17740,N_15896);
and UO_536 (O_536,N_19515,N_18984);
or UO_537 (O_537,N_15320,N_16299);
nor UO_538 (O_538,N_17807,N_16175);
nand UO_539 (O_539,N_19557,N_19948);
xnor UO_540 (O_540,N_15494,N_17338);
and UO_541 (O_541,N_15980,N_19404);
nor UO_542 (O_542,N_18041,N_17812);
nand UO_543 (O_543,N_17123,N_15103);
nor UO_544 (O_544,N_19692,N_15841);
nand UO_545 (O_545,N_16418,N_15931);
or UO_546 (O_546,N_15859,N_17387);
nand UO_547 (O_547,N_19319,N_16122);
and UO_548 (O_548,N_15457,N_18147);
and UO_549 (O_549,N_19718,N_19015);
or UO_550 (O_550,N_15530,N_15618);
nand UO_551 (O_551,N_19583,N_16790);
and UO_552 (O_552,N_15339,N_16659);
nor UO_553 (O_553,N_16812,N_15789);
or UO_554 (O_554,N_19552,N_16315);
nand UO_555 (O_555,N_18066,N_18773);
nand UO_556 (O_556,N_15132,N_15042);
and UO_557 (O_557,N_15250,N_18076);
and UO_558 (O_558,N_15983,N_19702);
and UO_559 (O_559,N_15124,N_19094);
and UO_560 (O_560,N_19072,N_17850);
xnor UO_561 (O_561,N_16618,N_17645);
nand UO_562 (O_562,N_16307,N_17679);
xor UO_563 (O_563,N_18820,N_17165);
or UO_564 (O_564,N_15764,N_16135);
nor UO_565 (O_565,N_17508,N_19568);
nor UO_566 (O_566,N_19766,N_17150);
and UO_567 (O_567,N_16457,N_17639);
nor UO_568 (O_568,N_17097,N_19598);
nor UO_569 (O_569,N_15409,N_18012);
and UO_570 (O_570,N_16319,N_17326);
or UO_571 (O_571,N_15817,N_15402);
nand UO_572 (O_572,N_18801,N_16925);
xnor UO_573 (O_573,N_16647,N_17458);
nor UO_574 (O_574,N_17134,N_15780);
nand UO_575 (O_575,N_17269,N_15065);
or UO_576 (O_576,N_18478,N_15559);
or UO_577 (O_577,N_19140,N_15869);
nand UO_578 (O_578,N_18907,N_17511);
nor UO_579 (O_579,N_15898,N_15611);
or UO_580 (O_580,N_17702,N_15643);
and UO_581 (O_581,N_16130,N_15435);
and UO_582 (O_582,N_18716,N_15258);
or UO_583 (O_583,N_19437,N_17048);
or UO_584 (O_584,N_19909,N_15159);
nor UO_585 (O_585,N_17532,N_18509);
nand UO_586 (O_586,N_18882,N_18376);
or UO_587 (O_587,N_16207,N_18750);
nand UO_588 (O_588,N_16475,N_19258);
xor UO_589 (O_589,N_19745,N_18058);
nand UO_590 (O_590,N_19159,N_18616);
or UO_591 (O_591,N_16738,N_18353);
nand UO_592 (O_592,N_17157,N_15438);
or UO_593 (O_593,N_19443,N_19730);
or UO_594 (O_594,N_18164,N_17820);
nor UO_595 (O_595,N_16872,N_19654);
nor UO_596 (O_596,N_15991,N_15904);
nand UO_597 (O_597,N_16243,N_18659);
xnor UO_598 (O_598,N_15327,N_17788);
nand UO_599 (O_599,N_15645,N_18935);
nand UO_600 (O_600,N_15985,N_16778);
and UO_601 (O_601,N_15852,N_16018);
nand UO_602 (O_602,N_19272,N_17128);
nand UO_603 (O_603,N_15853,N_16928);
or UO_604 (O_604,N_19293,N_15120);
or UO_605 (O_605,N_18932,N_16813);
nor UO_606 (O_606,N_19428,N_16718);
nand UO_607 (O_607,N_19061,N_15376);
nor UO_608 (O_608,N_19199,N_15140);
or UO_609 (O_609,N_18011,N_15053);
xnor UO_610 (O_610,N_17724,N_17175);
nand UO_611 (O_611,N_18829,N_17730);
and UO_612 (O_612,N_15691,N_19338);
xnor UO_613 (O_613,N_16468,N_19146);
xor UO_614 (O_614,N_17287,N_16379);
xnor UO_615 (O_615,N_18877,N_15306);
and UO_616 (O_616,N_18890,N_17306);
nand UO_617 (O_617,N_17256,N_17966);
or UO_618 (O_618,N_19231,N_19229);
nand UO_619 (O_619,N_17591,N_17758);
nand UO_620 (O_620,N_15916,N_19477);
or UO_621 (O_621,N_15675,N_18018);
nor UO_622 (O_622,N_16978,N_16816);
and UO_623 (O_623,N_18867,N_15216);
nor UO_624 (O_624,N_17382,N_16063);
and UO_625 (O_625,N_18472,N_18113);
and UO_626 (O_626,N_18412,N_17863);
nor UO_627 (O_627,N_16148,N_16306);
nor UO_628 (O_628,N_17969,N_16746);
and UO_629 (O_629,N_16859,N_17562);
nand UO_630 (O_630,N_16184,N_15038);
and UO_631 (O_631,N_16704,N_17418);
and UO_632 (O_632,N_19233,N_16628);
nor UO_633 (O_633,N_18619,N_16729);
and UO_634 (O_634,N_17716,N_16150);
or UO_635 (O_635,N_18817,N_17443);
and UO_636 (O_636,N_18215,N_16768);
nand UO_637 (O_637,N_15190,N_16074);
xor UO_638 (O_638,N_17558,N_18839);
xnor UO_639 (O_639,N_19023,N_19600);
nand UO_640 (O_640,N_17074,N_17162);
and UO_641 (O_641,N_19816,N_18344);
and UO_642 (O_642,N_18030,N_16185);
and UO_643 (O_643,N_19843,N_17028);
nand UO_644 (O_644,N_19793,N_17084);
nor UO_645 (O_645,N_18917,N_15600);
nand UO_646 (O_646,N_17864,N_17132);
or UO_647 (O_647,N_18818,N_19111);
xnor UO_648 (O_648,N_18502,N_18458);
or UO_649 (O_649,N_17049,N_17513);
or UO_650 (O_650,N_17404,N_16852);
or UO_651 (O_651,N_17840,N_16361);
and UO_652 (O_652,N_18717,N_15305);
or UO_653 (O_653,N_18676,N_15542);
nor UO_654 (O_654,N_18633,N_19687);
nor UO_655 (O_655,N_16320,N_15717);
and UO_656 (O_656,N_17357,N_16561);
nand UO_657 (O_657,N_17188,N_19253);
nand UO_658 (O_658,N_15791,N_19291);
or UO_659 (O_659,N_15000,N_16966);
nand UO_660 (O_660,N_18710,N_16424);
nand UO_661 (O_661,N_17808,N_16583);
nor UO_662 (O_662,N_15669,N_17545);
or UO_663 (O_663,N_19983,N_15295);
and UO_664 (O_664,N_16693,N_19063);
nor UO_665 (O_665,N_16097,N_18888);
xor UO_666 (O_666,N_19454,N_16282);
xor UO_667 (O_667,N_18101,N_18340);
nor UO_668 (O_668,N_19020,N_15954);
nand UO_669 (O_669,N_16755,N_16082);
or UO_670 (O_670,N_17089,N_19375);
nor UO_671 (O_671,N_17971,N_18232);
and UO_672 (O_672,N_17297,N_19029);
nand UO_673 (O_673,N_15028,N_19612);
nand UO_674 (O_674,N_18936,N_19301);
and UO_675 (O_675,N_15745,N_19851);
or UO_676 (O_676,N_16403,N_15959);
nor UO_677 (O_677,N_15138,N_18293);
nand UO_678 (O_678,N_17203,N_17784);
or UO_679 (O_679,N_19543,N_18796);
or UO_680 (O_680,N_16737,N_16786);
or UO_681 (O_681,N_19548,N_18793);
nor UO_682 (O_682,N_17439,N_16083);
nand UO_683 (O_683,N_15943,N_18236);
or UO_684 (O_684,N_18630,N_19771);
nor UO_685 (O_685,N_15466,N_17090);
nor UO_686 (O_686,N_18027,N_18819);
and UO_687 (O_687,N_15621,N_15670);
and UO_688 (O_688,N_17078,N_19623);
or UO_689 (O_689,N_17229,N_18926);
xnor UO_690 (O_690,N_17929,N_19125);
and UO_691 (O_691,N_16750,N_16145);
nand UO_692 (O_692,N_17321,N_19191);
and UO_693 (O_693,N_15567,N_17528);
nor UO_694 (O_694,N_16268,N_19286);
and UO_695 (O_695,N_19307,N_18139);
and UO_696 (O_696,N_15510,N_17075);
or UO_697 (O_697,N_18432,N_19950);
and UO_698 (O_698,N_16188,N_19939);
nor UO_699 (O_699,N_17768,N_18039);
and UO_700 (O_700,N_18496,N_15182);
or UO_701 (O_701,N_18862,N_15531);
nand UO_702 (O_702,N_19857,N_18261);
xnor UO_703 (O_703,N_18375,N_17505);
and UO_704 (O_704,N_16810,N_17435);
and UO_705 (O_705,N_18534,N_16797);
and UO_706 (O_706,N_18199,N_19849);
or UO_707 (O_707,N_19986,N_19920);
and UO_708 (O_708,N_18138,N_18111);
nor UO_709 (O_709,N_18965,N_18015);
xnor UO_710 (O_710,N_15157,N_18557);
and UO_711 (O_711,N_17077,N_17607);
xor UO_712 (O_712,N_18902,N_18794);
or UO_713 (O_713,N_18308,N_15334);
and UO_714 (O_714,N_16722,N_16271);
nand UO_715 (O_715,N_17490,N_15580);
or UO_716 (O_716,N_19605,N_19363);
nor UO_717 (O_717,N_17416,N_19480);
or UO_718 (O_718,N_16111,N_15589);
and UO_719 (O_719,N_17476,N_19120);
nand UO_720 (O_720,N_19944,N_18615);
xnor UO_721 (O_721,N_15720,N_17584);
and UO_722 (O_722,N_16987,N_17220);
or UO_723 (O_723,N_17507,N_17731);
xor UO_724 (O_724,N_18431,N_16436);
or UO_725 (O_725,N_16241,N_16326);
or UO_726 (O_726,N_15412,N_17877);
nor UO_727 (O_727,N_19942,N_18814);
or UO_728 (O_728,N_17942,N_15754);
nor UO_729 (O_729,N_15631,N_16240);
and UO_730 (O_730,N_15968,N_15144);
and UO_731 (O_731,N_19423,N_15197);
and UO_732 (O_732,N_17380,N_19087);
nand UO_733 (O_733,N_15785,N_15992);
or UO_734 (O_734,N_15273,N_15681);
nand UO_735 (O_735,N_18729,N_16667);
nand UO_736 (O_736,N_15948,N_17995);
xor UO_737 (O_737,N_17030,N_18783);
nor UO_738 (O_738,N_15077,N_19122);
and UO_739 (O_739,N_17487,N_15489);
nor UO_740 (O_740,N_19091,N_16244);
nand UO_741 (O_741,N_15911,N_17689);
nor UO_742 (O_742,N_16940,N_17283);
xnor UO_743 (O_743,N_16221,N_18214);
or UO_744 (O_744,N_19753,N_19214);
xor UO_745 (O_745,N_17238,N_16172);
nand UO_746 (O_746,N_19081,N_16592);
and UO_747 (O_747,N_15063,N_19491);
or UO_748 (O_748,N_16330,N_16009);
nand UO_749 (O_749,N_16473,N_17582);
or UO_750 (O_750,N_18944,N_16295);
nand UO_751 (O_751,N_18990,N_17948);
nor UO_752 (O_752,N_16634,N_15786);
nor UO_753 (O_753,N_18566,N_19854);
and UO_754 (O_754,N_19903,N_19138);
nor UO_755 (O_755,N_19179,N_16780);
or UO_756 (O_756,N_19369,N_19677);
and UO_757 (O_757,N_16887,N_16364);
nor UO_758 (O_758,N_15213,N_15797);
nor UO_759 (O_759,N_15857,N_16926);
nor UO_760 (O_760,N_19608,N_19003);
nand UO_761 (O_761,N_17174,N_16789);
or UO_762 (O_762,N_17936,N_15056);
or UO_763 (O_763,N_19271,N_15861);
nand UO_764 (O_764,N_16417,N_17652);
and UO_765 (O_765,N_19243,N_17712);
and UO_766 (O_766,N_19137,N_16573);
or UO_767 (O_767,N_15039,N_17323);
xor UO_768 (O_768,N_16382,N_18144);
nor UO_769 (O_769,N_16420,N_16752);
or UO_770 (O_770,N_17925,N_18853);
or UO_771 (O_771,N_15460,N_19890);
xnor UO_772 (O_772,N_19662,N_17234);
nand UO_773 (O_773,N_18414,N_15325);
or UO_774 (O_774,N_15088,N_15810);
xnor UO_775 (O_775,N_17967,N_17677);
or UO_776 (O_776,N_16827,N_18274);
or UO_777 (O_777,N_16770,N_18727);
nor UO_778 (O_778,N_17996,N_15776);
and UO_779 (O_779,N_15073,N_17624);
nor UO_780 (O_780,N_18755,N_15541);
nor UO_781 (O_781,N_17351,N_19864);
or UO_782 (O_782,N_15894,N_18372);
nor UO_783 (O_783,N_17415,N_17769);
nor UO_784 (O_784,N_19947,N_15952);
nand UO_785 (O_785,N_16656,N_15324);
nand UO_786 (O_786,N_16347,N_18802);
xnor UO_787 (O_787,N_15288,N_18669);
xnor UO_788 (O_788,N_16957,N_18954);
or UO_789 (O_789,N_17983,N_15015);
or UO_790 (O_790,N_16889,N_16782);
nor UO_791 (O_791,N_18586,N_18369);
and UO_792 (O_792,N_19618,N_16625);
xor UO_793 (O_793,N_17900,N_15338);
nand UO_794 (O_794,N_15160,N_17935);
or UO_795 (O_795,N_17991,N_19863);
xnor UO_796 (O_796,N_16079,N_17500);
nor UO_797 (O_797,N_17125,N_17276);
nand UO_798 (O_798,N_17273,N_15393);
nand UO_799 (O_799,N_18510,N_15246);
and UO_800 (O_800,N_16843,N_18959);
and UO_801 (O_801,N_15750,N_17866);
nand UO_802 (O_802,N_18746,N_17091);
or UO_803 (O_803,N_19800,N_17705);
and UO_804 (O_804,N_19553,N_19050);
nand UO_805 (O_805,N_16552,N_19056);
nand UO_806 (O_806,N_15855,N_17263);
nand UO_807 (O_807,N_15491,N_18789);
nand UO_808 (O_808,N_18547,N_17575);
nand UO_809 (O_809,N_18413,N_18343);
xor UO_810 (O_810,N_19244,N_18393);
or UO_811 (O_811,N_19485,N_19567);
nor UO_812 (O_812,N_16386,N_15480);
or UO_813 (O_813,N_17862,N_15309);
or UO_814 (O_814,N_19471,N_17352);
and UO_815 (O_815,N_16305,N_18699);
or UO_816 (O_816,N_16946,N_17550);
xnor UO_817 (O_817,N_18884,N_18785);
nand UO_818 (O_818,N_16958,N_16651);
and UO_819 (O_819,N_16617,N_18927);
or UO_820 (O_820,N_18531,N_18258);
nor UO_821 (O_821,N_18210,N_16222);
or UO_822 (O_822,N_16703,N_18324);
nand UO_823 (O_823,N_16214,N_15106);
and UO_824 (O_824,N_16001,N_15835);
nor UO_825 (O_825,N_17790,N_18110);
nand UO_826 (O_826,N_17471,N_19194);
nor UO_827 (O_827,N_15446,N_18533);
and UO_828 (O_828,N_19426,N_15175);
nand UO_829 (O_829,N_15854,N_15411);
or UO_830 (O_830,N_15575,N_18821);
and UO_831 (O_831,N_18718,N_19649);
or UO_832 (O_832,N_19410,N_15374);
nand UO_833 (O_833,N_15771,N_16726);
nor UO_834 (O_834,N_15069,N_17771);
xnor UO_835 (O_835,N_18176,N_18595);
nand UO_836 (O_836,N_15599,N_16587);
nor UO_837 (O_837,N_15887,N_18433);
nor UO_838 (O_838,N_18169,N_16230);
nand UO_839 (O_839,N_16448,N_16971);
xnor UO_840 (O_840,N_19064,N_18088);
nor UO_841 (O_841,N_16213,N_19196);
nor UO_842 (O_842,N_15521,N_15096);
nand UO_843 (O_843,N_16566,N_19579);
nand UO_844 (O_844,N_19972,N_18901);
nor UO_845 (O_845,N_15194,N_18057);
xor UO_846 (O_846,N_15418,N_19985);
nand UO_847 (O_847,N_15901,N_15864);
and UO_848 (O_848,N_16930,N_16401);
and UO_849 (O_849,N_18757,N_19245);
and UO_850 (O_850,N_16570,N_17518);
or UO_851 (O_851,N_16809,N_15787);
nand UO_852 (O_852,N_17005,N_16098);
or UO_853 (O_853,N_16894,N_15998);
nor UO_854 (O_854,N_17739,N_15895);
nor UO_855 (O_855,N_17556,N_18554);
nor UO_856 (O_856,N_17291,N_15632);
nor UO_857 (O_857,N_17278,N_15227);
and UO_858 (O_858,N_17309,N_18722);
nor UO_859 (O_859,N_15188,N_18996);
or UO_860 (O_860,N_18731,N_19493);
nand UO_861 (O_861,N_17314,N_19925);
nand UO_862 (O_862,N_19699,N_17065);
nand UO_863 (O_863,N_18103,N_17299);
xnor UO_864 (O_864,N_17377,N_19929);
nand UO_865 (O_865,N_19840,N_18342);
or UO_866 (O_866,N_19697,N_15741);
and UO_867 (O_867,N_15726,N_19820);
and UO_868 (O_868,N_19285,N_15059);
or UO_869 (O_869,N_18653,N_15331);
nor UO_870 (O_870,N_18366,N_17917);
or UO_871 (O_871,N_15885,N_15814);
nand UO_872 (O_872,N_15970,N_15359);
or UO_873 (O_873,N_17146,N_16162);
and UO_874 (O_874,N_18606,N_18408);
or UO_875 (O_875,N_18514,N_19143);
and UO_876 (O_876,N_17288,N_18908);
and UO_877 (O_877,N_19335,N_16354);
nor UO_878 (O_878,N_17052,N_15767);
or UO_879 (O_879,N_17053,N_15379);
nand UO_880 (O_880,N_16487,N_17636);
and UO_881 (O_881,N_15875,N_17887);
nand UO_882 (O_882,N_15243,N_19796);
xor UO_883 (O_883,N_17599,N_19373);
or UO_884 (O_884,N_18992,N_17230);
nor UO_885 (O_885,N_15816,N_15221);
nand UO_886 (O_886,N_17141,N_17156);
nand UO_887 (O_887,N_18427,N_15584);
or UO_888 (O_888,N_18749,N_17973);
nand UO_889 (O_889,N_18480,N_15110);
nor UO_890 (O_890,N_15094,N_17169);
nand UO_891 (O_891,N_18092,N_18269);
and UO_892 (O_892,N_15891,N_16571);
and UO_893 (O_893,N_15497,N_15355);
nor UO_894 (O_894,N_18866,N_18513);
and UO_895 (O_895,N_15740,N_19099);
and UO_896 (O_896,N_15881,N_16507);
nand UO_897 (O_897,N_18190,N_15844);
nand UO_898 (O_898,N_15283,N_16591);
xnor UO_899 (O_899,N_16998,N_16179);
nand UO_900 (O_900,N_19719,N_16660);
nor UO_901 (O_901,N_15228,N_18301);
nand UO_902 (O_902,N_18085,N_19542);
nor UO_903 (O_903,N_17939,N_18790);
nor UO_904 (O_904,N_19030,N_16146);
or UO_905 (O_905,N_15628,N_18145);
or UO_906 (O_906,N_16898,N_18574);
nor UO_907 (O_907,N_17551,N_15413);
nand UO_908 (O_908,N_17643,N_18130);
or UO_909 (O_909,N_19901,N_16236);
nor UO_910 (O_910,N_15192,N_19304);
and UO_911 (O_911,N_19161,N_16496);
and UO_912 (O_912,N_16706,N_15370);
nand UO_913 (O_913,N_18224,N_15233);
nand UO_914 (O_914,N_18070,N_16663);
or UO_915 (O_915,N_19987,N_17986);
xor UO_916 (O_916,N_16695,N_18002);
or UO_917 (O_917,N_17903,N_19430);
nor UO_918 (O_918,N_18279,N_17122);
or UO_919 (O_919,N_19621,N_17680);
nor UO_920 (O_920,N_18730,N_15607);
xnor UO_921 (O_921,N_18808,N_18769);
and UO_922 (O_922,N_16251,N_16962);
nor UO_923 (O_923,N_18356,N_17821);
nor UO_924 (O_924,N_15514,N_18299);
nand UO_925 (O_925,N_16830,N_18938);
nand UO_926 (O_926,N_19530,N_15661);
nor UO_927 (O_927,N_19035,N_17629);
or UO_928 (O_928,N_19860,N_19465);
nand UO_929 (O_929,N_17147,N_18622);
xnor UO_930 (O_930,N_18799,N_19651);
nor UO_931 (O_931,N_16598,N_15236);
nand UO_932 (O_932,N_17729,N_15486);
or UO_933 (O_933,N_18446,N_17658);
or UO_934 (O_934,N_16199,N_19825);
nor UO_935 (O_935,N_15688,N_15445);
or UO_936 (O_936,N_15198,N_19640);
nand UO_937 (O_937,N_17896,N_19846);
and UO_938 (O_938,N_18609,N_17910);
nor UO_939 (O_939,N_17112,N_17846);
nand UO_940 (O_940,N_16105,N_17121);
and UO_941 (O_941,N_18390,N_15845);
nand UO_942 (O_942,N_19398,N_16975);
nor UO_943 (O_943,N_19822,N_17414);
and UO_944 (O_944,N_18587,N_18837);
nand UO_945 (O_945,N_15515,N_15292);
and UO_946 (O_946,N_17542,N_16776);
and UO_947 (O_947,N_17786,N_15788);
nor UO_948 (O_948,N_16183,N_16039);
xor UO_949 (O_949,N_18398,N_18129);
or UO_950 (O_950,N_15779,N_17469);
nor UO_951 (O_951,N_18754,N_16421);
nand UO_952 (O_952,N_17127,N_16309);
xor UO_953 (O_953,N_17710,N_19283);
xor UO_954 (O_954,N_18119,N_18038);
or UO_955 (O_955,N_16743,N_18698);
and UO_956 (O_956,N_15322,N_15577);
nor UO_957 (O_957,N_19747,N_19574);
nand UO_958 (O_958,N_16638,N_17774);
and UO_959 (O_959,N_18465,N_15201);
and UO_960 (O_960,N_15656,N_18781);
and UO_961 (O_961,N_18807,N_19610);
or UO_962 (O_962,N_17191,N_16532);
or UO_963 (O_963,N_15601,N_16211);
or UO_964 (O_964,N_16325,N_15254);
and UO_965 (O_965,N_16020,N_15579);
or UO_966 (O_966,N_19472,N_16661);
nand UO_967 (O_967,N_15345,N_16973);
or UO_968 (O_968,N_15526,N_16252);
nor UO_969 (O_969,N_17473,N_19964);
or UO_970 (O_970,N_16867,N_18334);
or UO_971 (O_971,N_19773,N_18770);
or UO_972 (O_972,N_15999,N_19403);
or UO_973 (O_973,N_18125,N_17257);
nand UO_974 (O_974,N_18162,N_16800);
xor UO_975 (O_975,N_15827,N_17058);
nor UO_976 (O_976,N_16341,N_15128);
nand UO_977 (O_977,N_15200,N_17692);
or UO_978 (O_978,N_18660,N_16749);
or UO_979 (O_979,N_19535,N_17187);
and UO_980 (O_980,N_17576,N_15049);
nand UO_981 (O_981,N_18691,N_19528);
and UO_982 (O_982,N_16086,N_15303);
nor UO_983 (O_983,N_19238,N_16613);
and UO_984 (O_984,N_19970,N_19374);
or UO_985 (O_985,N_17711,N_16012);
or UO_986 (O_986,N_19075,N_15727);
and UO_987 (O_987,N_18976,N_17254);
nor UO_988 (O_988,N_19222,N_17685);
nand UO_989 (O_989,N_19005,N_18626);
nor UO_990 (O_990,N_16254,N_19511);
and UO_991 (O_991,N_18813,N_15009);
and UO_992 (O_992,N_17797,N_15654);
and UO_993 (O_993,N_17167,N_16596);
or UO_994 (O_994,N_16229,N_16525);
and UO_995 (O_995,N_19891,N_19876);
nor UO_996 (O_996,N_19206,N_17465);
nor UO_997 (O_997,N_18627,N_19531);
or UO_998 (O_998,N_15134,N_18281);
nor UO_999 (O_999,N_18314,N_16544);
nand UO_1000 (O_1000,N_17874,N_15400);
nand UO_1001 (O_1001,N_16639,N_18272);
nand UO_1002 (O_1002,N_18255,N_15929);
nand UO_1003 (O_1003,N_18728,N_15658);
xnor UO_1004 (O_1004,N_17686,N_16607);
nand UO_1005 (O_1005,N_17109,N_19467);
or UO_1006 (O_1006,N_15988,N_19996);
and UO_1007 (O_1007,N_16801,N_19900);
nor UO_1008 (O_1008,N_17901,N_15739);
and UO_1009 (O_1009,N_15260,N_17883);
nand UO_1010 (O_1010,N_19659,N_15973);
and UO_1011 (O_1011,N_19482,N_18734);
xnor UO_1012 (O_1012,N_16906,N_15425);
or UO_1013 (O_1013,N_17186,N_19256);
nand UO_1014 (O_1014,N_16494,N_15603);
and UO_1015 (O_1015,N_16877,N_17859);
nor UO_1016 (O_1016,N_15229,N_18098);
or UO_1017 (O_1017,N_17653,N_18148);
or UO_1018 (O_1018,N_18387,N_19236);
xnor UO_1019 (O_1019,N_16288,N_17260);
and UO_1020 (O_1020,N_18404,N_15863);
and UO_1021 (O_1021,N_15153,N_15395);
and UO_1022 (O_1022,N_16192,N_18292);
and UO_1023 (O_1023,N_17329,N_15090);
nor UO_1024 (O_1024,N_17095,N_17375);
and UO_1025 (O_1025,N_19390,N_19707);
and UO_1026 (O_1026,N_15455,N_19868);
and UO_1027 (O_1027,N_19647,N_18291);
nand UO_1028 (O_1028,N_15108,N_16445);
or UO_1029 (O_1029,N_17782,N_16825);
or UO_1030 (O_1030,N_18006,N_19496);
nand UO_1031 (O_1031,N_19735,N_18816);
nand UO_1032 (O_1032,N_18603,N_18487);
xnor UO_1033 (O_1033,N_15386,N_18358);
xor UO_1034 (O_1034,N_18858,N_16302);
and UO_1035 (O_1035,N_16351,N_18023);
and UO_1036 (O_1036,N_17580,N_18010);
nand UO_1037 (O_1037,N_15588,N_15378);
nor UO_1038 (O_1038,N_16875,N_19366);
and UO_1039 (O_1039,N_17799,N_18900);
nor UO_1040 (O_1040,N_15808,N_18003);
xnor UO_1041 (O_1041,N_16929,N_18379);
nand UO_1042 (O_1042,N_18024,N_15960);
or UO_1043 (O_1043,N_17612,N_17713);
nor UO_1044 (O_1044,N_16204,N_19752);
nand UO_1045 (O_1045,N_18685,N_19541);
xnor UO_1046 (O_1046,N_17192,N_19756);
nand UO_1047 (O_1047,N_18664,N_19171);
or UO_1048 (O_1048,N_19492,N_17222);
or UO_1049 (O_1049,N_19275,N_16736);
nand UO_1050 (O_1050,N_18501,N_15773);
or UO_1051 (O_1051,N_16374,N_15424);
or UO_1052 (O_1052,N_19033,N_17714);
nand UO_1053 (O_1053,N_18337,N_15874);
or UO_1054 (O_1054,N_16725,N_17143);
and UO_1055 (O_1055,N_15705,N_16698);
xnor UO_1056 (O_1056,N_17477,N_16380);
and UO_1057 (O_1057,N_15932,N_18714);
or UO_1058 (O_1058,N_17087,N_18744);
nand UO_1059 (O_1059,N_18787,N_17848);
nand UO_1060 (O_1060,N_19802,N_19100);
nand UO_1061 (O_1061,N_16627,N_18044);
and UO_1062 (O_1062,N_17164,N_19921);
and UO_1063 (O_1063,N_15113,N_16140);
nand UO_1064 (O_1064,N_17564,N_19782);
or UO_1065 (O_1065,N_17603,N_16697);
or UO_1066 (O_1066,N_17588,N_16488);
nand UO_1067 (O_1067,N_17696,N_15562);
nor UO_1068 (O_1068,N_16173,N_16538);
nor UO_1069 (O_1069,N_19705,N_17566);
nand UO_1070 (O_1070,N_18577,N_16581);
nor UO_1071 (O_1071,N_18692,N_16710);
xor UO_1072 (O_1072,N_17704,N_17311);
and UO_1073 (O_1073,N_19726,N_16317);
or UO_1074 (O_1074,N_18997,N_16195);
or UO_1075 (O_1075,N_19277,N_18719);
nor UO_1076 (O_1076,N_19912,N_16066);
nor UO_1077 (O_1077,N_15364,N_18524);
nor UO_1078 (O_1078,N_15760,N_16419);
and UO_1079 (O_1079,N_16449,N_16979);
and UO_1080 (O_1080,N_19419,N_15956);
or UO_1081 (O_1081,N_18894,N_15573);
nand UO_1082 (O_1082,N_15451,N_17569);
nand UO_1083 (O_1083,N_15087,N_18593);
nor UO_1084 (O_1084,N_15405,N_18371);
and UO_1085 (O_1085,N_15525,N_17140);
nor UO_1086 (O_1086,N_15536,N_15382);
xnor UO_1087 (O_1087,N_16077,N_19870);
nand UO_1088 (O_1088,N_17255,N_15186);
nor UO_1089 (O_1089,N_19774,N_16447);
nor UO_1090 (O_1090,N_18635,N_19073);
nor UO_1091 (O_1091,N_18835,N_17698);
and UO_1092 (O_1092,N_15940,N_16643);
and UO_1093 (O_1093,N_19866,N_17872);
or UO_1094 (O_1094,N_19340,N_19590);
nor UO_1095 (O_1095,N_19447,N_19115);
xor UO_1096 (O_1096,N_18569,N_15145);
nor UO_1097 (O_1097,N_19126,N_17016);
or UO_1098 (O_1098,N_18693,N_15831);
nand UO_1099 (O_1099,N_15337,N_19180);
and UO_1100 (O_1100,N_15692,N_17510);
nand UO_1101 (O_1101,N_16126,N_16674);
or UO_1102 (O_1102,N_16408,N_19715);
and UO_1103 (O_1103,N_17423,N_18084);
and UO_1104 (O_1104,N_18708,N_15560);
and UO_1105 (O_1105,N_16095,N_15482);
and UO_1106 (O_1106,N_17426,N_19856);
and UO_1107 (O_1107,N_16791,N_16861);
nand UO_1108 (O_1108,N_18086,N_16092);
nor UO_1109 (O_1109,N_16530,N_18461);
nand UO_1110 (O_1110,N_16937,N_19737);
nand UO_1111 (O_1111,N_15176,N_17076);
or UO_1112 (O_1112,N_19845,N_19631);
nor UO_1113 (O_1113,N_15100,N_15155);
nand UO_1114 (O_1114,N_16936,N_16502);
nand UO_1115 (O_1115,N_19638,N_18854);
nand UO_1116 (O_1116,N_17623,N_16762);
nor UO_1117 (O_1117,N_16177,N_16719);
or UO_1118 (O_1118,N_17522,N_18470);
xor UO_1119 (O_1119,N_18594,N_19877);
and UO_1120 (O_1120,N_16684,N_15982);
nor UO_1121 (O_1121,N_17391,N_18211);
and UO_1122 (O_1122,N_16266,N_19052);
or UO_1123 (O_1123,N_18897,N_16477);
and UO_1124 (O_1124,N_16158,N_16227);
nor UO_1125 (O_1125,N_18686,N_16980);
xor UO_1126 (O_1126,N_19469,N_18702);
and UO_1127 (O_1127,N_19932,N_19951);
nor UO_1128 (O_1128,N_19018,N_15093);
nor UO_1129 (O_1129,N_19069,N_16334);
or UO_1130 (O_1130,N_16539,N_18919);
or UO_1131 (O_1131,N_18999,N_19178);
nor UO_1132 (O_1132,N_17622,N_17161);
or UO_1133 (O_1133,N_19004,N_19422);
xnor UO_1134 (O_1134,N_16992,N_15918);
or UO_1135 (O_1135,N_17755,N_17827);
nand UO_1136 (O_1136,N_19637,N_15167);
nor UO_1137 (O_1137,N_16673,N_19239);
and UO_1138 (O_1138,N_19562,N_18966);
nand UO_1139 (O_1139,N_18518,N_19370);
nor UO_1140 (O_1140,N_17749,N_19070);
nand UO_1141 (O_1141,N_16910,N_17389);
nor UO_1142 (O_1142,N_18095,N_19312);
nand UO_1143 (O_1143,N_17024,N_15585);
or UO_1144 (O_1144,N_15265,N_17557);
or UO_1145 (O_1145,N_17746,N_16280);
and UO_1146 (O_1146,N_15477,N_16238);
or UO_1147 (O_1147,N_18498,N_15329);
nand UO_1148 (O_1148,N_16489,N_17099);
xnor UO_1149 (O_1149,N_18078,N_17789);
nor UO_1150 (O_1150,N_19894,N_16461);
nand UO_1151 (O_1151,N_17395,N_15044);
nand UO_1152 (O_1152,N_15928,N_16732);
or UO_1153 (O_1153,N_15971,N_19008);
nor UO_1154 (O_1154,N_17947,N_18977);
nor UO_1155 (O_1155,N_18419,N_17882);
xnor UO_1156 (O_1156,N_16125,N_15333);
nand UO_1157 (O_1157,N_17852,N_18874);
nor UO_1158 (O_1158,N_16691,N_18004);
or UO_1159 (O_1159,N_16977,N_16168);
nor UO_1160 (O_1160,N_18715,N_15005);
nor UO_1161 (O_1161,N_19198,N_19700);
nand UO_1162 (O_1162,N_17316,N_17906);
nor UO_1163 (O_1163,N_17198,N_17145);
and UO_1164 (O_1164,N_17956,N_16774);
or UO_1165 (O_1165,N_15604,N_16677);
or UO_1166 (O_1166,N_17138,N_16262);
nand UO_1167 (O_1167,N_16405,N_16524);
and UO_1168 (O_1168,N_16181,N_15488);
nand UO_1169 (O_1169,N_17111,N_18864);
and UO_1170 (O_1170,N_16694,N_16438);
and UO_1171 (O_1171,N_19648,N_15839);
and UO_1172 (O_1172,N_15862,N_19154);
and UO_1173 (O_1173,N_19065,N_19208);
nor UO_1174 (O_1174,N_19327,N_15693);
or UO_1175 (O_1175,N_19818,N_16002);
or UO_1176 (O_1176,N_15616,N_18083);
nand UO_1177 (O_1177,N_17168,N_16434);
and UO_1178 (O_1178,N_18511,N_16556);
and UO_1179 (O_1179,N_15414,N_19833);
and UO_1180 (O_1180,N_15678,N_15592);
or UO_1181 (O_1181,N_19517,N_15261);
nor UO_1182 (O_1182,N_17051,N_16372);
nor UO_1183 (O_1183,N_15476,N_19175);
and UO_1184 (O_1184,N_15427,N_17646);
nor UO_1185 (O_1185,N_16716,N_18591);
and UO_1186 (O_1186,N_19372,N_19869);
or UO_1187 (O_1187,N_16383,N_15824);
or UO_1188 (O_1188,N_18127,N_18742);
nor UO_1189 (O_1189,N_15045,N_17750);
and UO_1190 (O_1190,N_16531,N_18068);
nor UO_1191 (O_1191,N_17688,N_18367);
nand UO_1192 (O_1192,N_17955,N_17826);
and UO_1193 (O_1193,N_18322,N_19119);
and UO_1194 (O_1194,N_16970,N_15203);
nand UO_1195 (O_1195,N_19886,N_17092);
or UO_1196 (O_1196,N_15156,N_17386);
or UO_1197 (O_1197,N_17951,N_16505);
nor UO_1198 (O_1198,N_15116,N_16912);
nand UO_1199 (O_1199,N_16542,N_16713);
nor UO_1200 (O_1200,N_18759,N_19619);
nor UO_1201 (O_1201,N_17354,N_15392);
nand UO_1202 (O_1202,N_15664,N_17082);
nand UO_1203 (O_1203,N_18525,N_17665);
or UO_1204 (O_1204,N_18474,N_17932);
nor UO_1205 (O_1205,N_16856,N_16788);
xor UO_1206 (O_1206,N_18968,N_18218);
and UO_1207 (O_1207,N_18519,N_16584);
xnor UO_1208 (O_1208,N_18443,N_19803);
nor UO_1209 (O_1209,N_16504,N_17006);
xor UO_1210 (O_1210,N_17924,N_17833);
xnor UO_1211 (O_1211,N_19323,N_19658);
and UO_1212 (O_1212,N_16557,N_17452);
nand UO_1213 (O_1213,N_16851,N_18081);
nor UO_1214 (O_1214,N_18149,N_18925);
xor UO_1215 (O_1215,N_18532,N_19724);
or UO_1216 (O_1216,N_16197,N_15057);
nand UO_1217 (O_1217,N_19365,N_17370);
nand UO_1218 (O_1218,N_19824,N_18226);
or UO_1219 (O_1219,N_15220,N_19977);
or UO_1220 (O_1220,N_18283,N_15350);
nand UO_1221 (O_1221,N_17880,N_16028);
nand UO_1222 (O_1222,N_15660,N_16772);
or UO_1223 (O_1223,N_18280,N_17101);
nand UO_1224 (O_1224,N_19933,N_18998);
and UO_1225 (O_1225,N_16523,N_19988);
nor UO_1226 (O_1226,N_15181,N_17043);
nor UO_1227 (O_1227,N_17776,N_19908);
or UO_1228 (O_1228,N_16938,N_19888);
and UO_1229 (O_1229,N_18942,N_19733);
nand UO_1230 (O_1230,N_19585,N_19057);
and UO_1231 (O_1231,N_17800,N_18439);
or UO_1232 (O_1232,N_15870,N_17225);
and UO_1233 (O_1233,N_18007,N_19789);
nand UO_1234 (O_1234,N_16951,N_15369);
nor UO_1235 (O_1235,N_19969,N_15007);
and UO_1236 (O_1236,N_16072,N_15419);
nor UO_1237 (O_1237,N_18971,N_18810);
xnor UO_1238 (O_1238,N_15185,N_19593);
nand UO_1239 (O_1239,N_19599,N_17502);
nor UO_1240 (O_1240,N_15529,N_15211);
nor UO_1241 (O_1241,N_15602,N_19917);
or UO_1242 (O_1242,N_19408,N_19478);
and UO_1243 (O_1243,N_16060,N_16154);
and UO_1244 (O_1244,N_19136,N_17265);
and UO_1245 (O_1245,N_19355,N_16818);
xnor UO_1246 (O_1246,N_18021,N_18766);
and UO_1247 (O_1247,N_19487,N_19172);
and UO_1248 (O_1248,N_17832,N_15897);
nand UO_1249 (O_1249,N_18492,N_18381);
or UO_1250 (O_1250,N_18544,N_18663);
or UO_1251 (O_1251,N_17200,N_18550);
xor UO_1252 (O_1252,N_15011,N_17475);
or UO_1253 (O_1253,N_15509,N_19968);
and UO_1254 (O_1254,N_19871,N_18652);
or UO_1255 (O_1255,N_16601,N_17606);
or UO_1256 (O_1256,N_18695,N_17104);
nand UO_1257 (O_1257,N_16270,N_15080);
and UO_1258 (O_1258,N_18937,N_19089);
or UO_1259 (O_1259,N_15294,N_17208);
xnor UO_1260 (O_1260,N_15268,N_16517);
or UO_1261 (O_1261,N_16549,N_19708);
nand UO_1262 (O_1262,N_17778,N_19402);
or UO_1263 (O_1263,N_19769,N_16356);
and UO_1264 (O_1264,N_16679,N_17020);
and UO_1265 (O_1265,N_17794,N_18910);
nand UO_1266 (O_1266,N_16483,N_17634);
or UO_1267 (O_1267,N_17251,N_15067);
nor UO_1268 (O_1268,N_18561,N_16413);
or UO_1269 (O_1269,N_19721,N_17365);
and UO_1270 (O_1270,N_19931,N_17535);
nor UO_1271 (O_1271,N_15426,N_18564);
and UO_1272 (O_1272,N_17029,N_15449);
and UO_1273 (O_1273,N_16533,N_19009);
nand UO_1274 (O_1274,N_15620,N_15210);
nand UO_1275 (O_1275,N_17890,N_16893);
nand UO_1276 (O_1276,N_18471,N_18182);
nor UO_1277 (O_1277,N_19734,N_16462);
xor UO_1278 (O_1278,N_18726,N_15219);
nor UO_1279 (O_1279,N_19027,N_18898);
and UO_1280 (O_1280,N_19071,N_19259);
or UO_1281 (O_1281,N_17861,N_15223);
nor UO_1282 (O_1282,N_17691,N_16275);
or UO_1283 (O_1283,N_16059,N_19963);
or UO_1284 (O_1284,N_16960,N_17185);
nand UO_1285 (O_1285,N_18267,N_15770);
nand UO_1286 (O_1286,N_15344,N_17093);
nor UO_1287 (O_1287,N_17170,N_19999);
nor UO_1288 (O_1288,N_17965,N_19330);
xor UO_1289 (O_1289,N_16124,N_17801);
nor UO_1290 (O_1290,N_16119,N_17240);
and UO_1291 (O_1291,N_15635,N_18000);
xnor UO_1292 (O_1292,N_17436,N_18945);
nand UO_1293 (O_1293,N_17361,N_15029);
or UO_1294 (O_1294,N_15778,N_17023);
xor UO_1295 (O_1295,N_17027,N_16328);
and UO_1296 (O_1296,N_19613,N_18712);
or UO_1297 (O_1297,N_18104,N_17615);
nand UO_1298 (O_1298,N_19356,N_18800);
nand UO_1299 (O_1299,N_17954,N_19806);
or UO_1300 (O_1300,N_16338,N_19192);
and UO_1301 (O_1301,N_19607,N_18767);
nor UO_1302 (O_1302,N_17663,N_16237);
nor UO_1303 (O_1303,N_16051,N_18306);
or UO_1304 (O_1304,N_16360,N_17313);
nor UO_1305 (O_1305,N_19104,N_16905);
or UO_1306 (O_1306,N_19434,N_15105);
xor UO_1307 (O_1307,N_18931,N_18947);
xor UO_1308 (O_1308,N_16857,N_19611);
nand UO_1309 (O_1309,N_18658,N_19168);
nor UO_1310 (O_1310,N_18317,N_19879);
or UO_1311 (O_1311,N_19698,N_16739);
or UO_1312 (O_1312,N_16822,N_17204);
nand UO_1313 (O_1313,N_18560,N_19078);
nand UO_1314 (O_1314,N_19653,N_17474);
xor UO_1315 (O_1315,N_17611,N_19838);
or UO_1316 (O_1316,N_17767,N_18409);
nor UO_1317 (O_1317,N_17930,N_19169);
nor UO_1318 (O_1318,N_15674,N_16766);
nand UO_1319 (O_1319,N_16537,N_16630);
xor UO_1320 (O_1320,N_15842,N_17902);
nand UO_1321 (O_1321,N_15214,N_16290);
or UO_1322 (O_1322,N_18795,N_15752);
and UO_1323 (O_1323,N_17638,N_17547);
nand UO_1324 (O_1324,N_15212,N_19043);
or UO_1325 (O_1325,N_17979,N_19039);
and UO_1326 (O_1326,N_17656,N_19346);
nand UO_1327 (O_1327,N_16149,N_18978);
nor UO_1328 (O_1328,N_18191,N_19704);
and UO_1329 (O_1329,N_15627,N_17884);
nand UO_1330 (O_1330,N_16452,N_17682);
or UO_1331 (O_1331,N_19709,N_17424);
nand UO_1332 (O_1332,N_19060,N_16783);
or UO_1333 (O_1333,N_15137,N_16814);
or UO_1334 (O_1334,N_17870,N_16235);
nand UO_1335 (O_1335,N_16407,N_16376);
and UO_1336 (O_1336,N_18546,N_16285);
nand UO_1337 (O_1337,N_16291,N_16522);
or UO_1338 (O_1338,N_19810,N_17271);
and UO_1339 (O_1339,N_15838,N_17000);
or UO_1340 (O_1340,N_18868,N_18612);
nor UO_1341 (O_1341,N_18760,N_16855);
xor UO_1342 (O_1342,N_15724,N_18929);
nand UO_1343 (O_1343,N_16769,N_19387);
nor UO_1344 (O_1344,N_15849,N_18848);
nand UO_1345 (O_1345,N_16993,N_17980);
nor UO_1346 (O_1346,N_18475,N_18171);
and UO_1347 (O_1347,N_19288,N_18503);
and UO_1348 (O_1348,N_18536,N_19971);
nor UO_1349 (O_1349,N_19350,N_18108);
nand UO_1350 (O_1350,N_18928,N_19420);
and UO_1351 (O_1351,N_16480,N_19642);
nand UO_1352 (O_1352,N_16519,N_16547);
xnor UO_1353 (O_1353,N_17707,N_19938);
nand UO_1354 (O_1354,N_16067,N_16521);
xnor UO_1355 (O_1355,N_17671,N_18046);
and UO_1356 (O_1356,N_17501,N_15377);
nor UO_1357 (O_1357,N_19512,N_19603);
or UO_1358 (O_1358,N_15417,N_19490);
xnor UO_1359 (O_1359,N_18457,N_17943);
nand UO_1360 (O_1360,N_19096,N_15089);
or UO_1361 (O_1361,N_15461,N_19024);
nor UO_1362 (O_1362,N_19054,N_19142);
or UO_1363 (O_1363,N_15571,N_19620);
nand UO_1364 (O_1364,N_16499,N_16976);
nand UO_1365 (O_1365,N_15910,N_17149);
or UO_1366 (O_1366,N_16619,N_19067);
or UO_1367 (O_1367,N_15484,N_19889);
nor UO_1368 (O_1368,N_19690,N_19501);
nand UO_1369 (O_1369,N_16422,N_19195);
nand UO_1370 (O_1370,N_16484,N_16267);
nor UO_1371 (O_1371,N_15668,N_16191);
and UO_1372 (O_1372,N_19048,N_16040);
nand UO_1373 (O_1373,N_15927,N_16701);
nand UO_1374 (O_1374,N_17911,N_15256);
or UO_1375 (O_1375,N_17703,N_17982);
nand UO_1376 (O_1376,N_15730,N_17587);
nand UO_1377 (O_1377,N_17070,N_16764);
nand UO_1378 (O_1378,N_15713,N_16279);
or UO_1379 (O_1379,N_16182,N_18670);
or UO_1380 (O_1380,N_17792,N_15703);
nor UO_1381 (O_1381,N_15708,N_16534);
or UO_1382 (O_1382,N_18256,N_15594);
or UO_1383 (O_1383,N_18009,N_15114);
and UO_1384 (O_1384,N_18605,N_18360);
nor UO_1385 (O_1385,N_18060,N_16171);
nand UO_1386 (O_1386,N_19533,N_15308);
or UO_1387 (O_1387,N_17383,N_19294);
and UO_1388 (O_1388,N_16096,N_19046);
nand UO_1389 (O_1389,N_18490,N_15276);
nor UO_1390 (O_1390,N_17630,N_16336);
nor UO_1391 (O_1391,N_19278,N_16250);
or UO_1392 (O_1392,N_15225,N_16337);
nand UO_1393 (O_1393,N_18768,N_17368);
and UO_1394 (O_1394,N_17307,N_17687);
or UO_1395 (O_1395,N_15765,N_15748);
nand UO_1396 (O_1396,N_19473,N_18825);
xnor UO_1397 (O_1397,N_15889,N_16298);
or UO_1398 (O_1398,N_18763,N_17757);
or UO_1399 (O_1399,N_17464,N_18923);
and UO_1400 (O_1400,N_18319,N_16820);
and UO_1401 (O_1401,N_18565,N_17199);
or UO_1402 (O_1402,N_16273,N_16506);
or UO_1403 (O_1403,N_18304,N_16840);
nor UO_1404 (O_1404,N_19240,N_15102);
or UO_1405 (O_1405,N_16920,N_19741);
or UO_1406 (O_1406,N_15646,N_16914);
and UO_1407 (O_1407,N_16160,N_15699);
nand UO_1408 (O_1408,N_18116,N_17292);
and UO_1409 (O_1409,N_19670,N_15572);
and UO_1410 (O_1410,N_16316,N_15456);
or UO_1411 (O_1411,N_15381,N_17324);
nor UO_1412 (O_1412,N_19483,N_17236);
or UO_1413 (O_1413,N_18477,N_17258);
or UO_1414 (O_1414,N_16866,N_17836);
nand UO_1415 (O_1415,N_18644,N_15723);
nand UO_1416 (O_1416,N_18774,N_17495);
and UO_1417 (O_1417,N_18241,N_15170);
nor UO_1418 (O_1418,N_17977,N_16367);
nand UO_1419 (O_1419,N_17727,N_16107);
or UO_1420 (O_1420,N_19695,N_19918);
nor UO_1421 (O_1421,N_18056,N_19577);
or UO_1422 (O_1422,N_19633,N_15061);
and UO_1423 (O_1423,N_15744,N_15649);
nor UO_1424 (O_1424,N_17339,N_17442);
and UO_1425 (O_1425,N_15834,N_17873);
nand UO_1426 (O_1426,N_18552,N_18911);
and UO_1427 (O_1427,N_15492,N_19566);
nand UO_1428 (O_1428,N_15274,N_19967);
nor UO_1429 (O_1429,N_19105,N_16300);
nand UO_1430 (O_1430,N_16717,N_19808);
nor UO_1431 (O_1431,N_19722,N_19333);
nand UO_1432 (O_1432,N_19220,N_19380);
nor UO_1433 (O_1433,N_16890,N_16075);
or UO_1434 (O_1434,N_15738,N_17069);
or UO_1435 (O_1435,N_15995,N_19466);
and UO_1436 (O_1436,N_15131,N_18614);
or UO_1437 (O_1437,N_19911,N_15257);
and UO_1438 (O_1438,N_16308,N_17455);
nor UO_1439 (O_1439,N_16707,N_16672);
nor UO_1440 (O_1440,N_16152,N_15947);
and UO_1441 (O_1441,N_16865,N_15519);
or UO_1442 (O_1442,N_19904,N_19026);
and UO_1443 (O_1443,N_18403,N_15147);
nor UO_1444 (O_1444,N_17176,N_17990);
nor UO_1445 (O_1445,N_18036,N_19794);
nor UO_1446 (O_1446,N_17209,N_18001);
and UO_1447 (O_1447,N_18826,N_15516);
xnor UO_1448 (O_1448,N_15673,N_18463);
or UO_1449 (O_1449,N_18842,N_19919);
xor UO_1450 (O_1450,N_19513,N_15353);
xnor UO_1451 (O_1451,N_18051,N_18684);
nor UO_1452 (O_1452,N_18806,N_16565);
nor UO_1453 (O_1453,N_19082,N_16653);
nand UO_1454 (O_1454,N_17277,N_18158);
or UO_1455 (O_1455,N_16385,N_19185);
xnor UO_1456 (O_1456,N_19162,N_19345);
and UO_1457 (O_1457,N_16014,N_18709);
nand UO_1458 (O_1458,N_15800,N_17120);
or UO_1459 (O_1459,N_17390,N_16631);
nor UO_1460 (O_1460,N_18838,N_17798);
and UO_1461 (O_1461,N_17441,N_16536);
nor UO_1462 (O_1462,N_19270,N_15432);
and UO_1463 (O_1463,N_16015,N_16010);
and UO_1464 (O_1464,N_17304,N_15753);
nor UO_1465 (O_1465,N_19088,N_19042);
or UO_1466 (O_1466,N_17497,N_17842);
and UO_1467 (O_1467,N_16120,N_18836);
or UO_1468 (O_1468,N_18674,N_15304);
nor UO_1469 (O_1469,N_16495,N_19265);
nor UO_1470 (O_1470,N_18167,N_18287);
xnor UO_1471 (O_1471,N_15177,N_19629);
nor UO_1472 (O_1472,N_15164,N_18756);
xnor UO_1473 (O_1473,N_17637,N_17635);
and UO_1474 (O_1474,N_17268,N_18683);
and UO_1475 (O_1475,N_19974,N_19205);
nor UO_1476 (O_1476,N_18545,N_18920);
nand UO_1477 (O_1477,N_16689,N_17483);
nor UO_1478 (O_1478,N_17319,N_16685);
nor UO_1479 (O_1479,N_16482,N_17197);
and UO_1480 (O_1480,N_16731,N_18495);
nor UO_1481 (O_1481,N_16668,N_19202);
and UO_1482 (O_1482,N_17617,N_15755);
nand UO_1483 (O_1483,N_17537,N_17350);
or UO_1484 (O_1484,N_18034,N_18231);
xor UO_1485 (O_1485,N_19519,N_17079);
or UO_1486 (O_1486,N_17379,N_19216);
nor UO_1487 (O_1487,N_15672,N_15207);
or UO_1488 (O_1488,N_16106,N_15081);
and UO_1489 (O_1489,N_15129,N_18863);
nor UO_1490 (O_1490,N_16259,N_17867);
and UO_1491 (O_1491,N_18303,N_16819);
xor UO_1492 (O_1492,N_19785,N_18374);
or UO_1493 (O_1493,N_17515,N_15180);
nand UO_1494 (O_1494,N_16470,N_18924);
nand UO_1495 (O_1495,N_18329,N_17738);
nor UO_1496 (O_1496,N_19446,N_15908);
nand UO_1497 (O_1497,N_18019,N_16311);
nor UO_1498 (O_1498,N_17107,N_15172);
nor UO_1499 (O_1499,N_18467,N_16301);
xnor UO_1500 (O_1500,N_18535,N_15154);
nor UO_1501 (O_1501,N_18137,N_15934);
and UO_1502 (O_1502,N_17302,N_17328);
and UO_1503 (O_1503,N_16642,N_18384);
xor UO_1504 (O_1504,N_16070,N_19571);
nand UO_1505 (O_1505,N_16043,N_16620);
nor UO_1506 (O_1506,N_18891,N_16610);
nand UO_1507 (O_1507,N_19795,N_16032);
and UO_1508 (O_1508,N_19188,N_16612);
xor UO_1509 (O_1509,N_17570,N_19852);
or UO_1510 (O_1510,N_17761,N_18655);
nand UO_1511 (O_1511,N_15130,N_19786);
nand UO_1512 (O_1512,N_16555,N_16068);
nor UO_1513 (O_1513,N_16817,N_19436);
or UO_1514 (O_1514,N_19770,N_17491);
or UO_1515 (O_1515,N_18650,N_19399);
or UO_1516 (O_1516,N_15495,N_15179);
nor UO_1517 (O_1517,N_15286,N_17376);
nor UO_1518 (O_1518,N_15371,N_18943);
xnor UO_1519 (O_1519,N_18880,N_15504);
xnor UO_1520 (O_1520,N_17802,N_16131);
nand UO_1521 (O_1521,N_16165,N_16127);
nand UO_1522 (O_1522,N_15848,N_17950);
nor UO_1523 (O_1523,N_19836,N_18732);
nand UO_1524 (O_1524,N_19758,N_17879);
nand UO_1525 (O_1525,N_17657,N_19905);
nor UO_1526 (O_1526,N_17809,N_16864);
nand UO_1527 (O_1527,N_18327,N_19524);
or UO_1528 (O_1528,N_18263,N_16363);
xor UO_1529 (O_1529,N_18861,N_19391);
or UO_1530 (O_1530,N_17928,N_18311);
and UO_1531 (O_1531,N_18689,N_15285);
and UO_1532 (O_1532,N_19397,N_16036);
or UO_1533 (O_1533,N_16568,N_15725);
nor UO_1534 (O_1534,N_18448,N_15490);
and UO_1535 (O_1535,N_18248,N_16795);
nor UO_1536 (O_1536,N_16708,N_15806);
nor UO_1537 (O_1537,N_18682,N_16000);
nand UO_1538 (O_1538,N_16269,N_18424);
nor UO_1539 (O_1539,N_19711,N_19433);
nand UO_1540 (O_1540,N_16318,N_17356);
and UO_1541 (O_1541,N_19614,N_17791);
nand UO_1542 (O_1542,N_16017,N_16093);
or UO_1543 (O_1543,N_16888,N_16626);
or UO_1544 (O_1544,N_18551,N_19990);
nor UO_1545 (O_1545,N_19744,N_15158);
nand UO_1546 (O_1546,N_15168,N_15064);
nor UO_1547 (O_1547,N_17062,N_16600);
or UO_1548 (O_1548,N_18391,N_18610);
or UO_1549 (O_1549,N_15768,N_15240);
nor UO_1550 (O_1550,N_17267,N_18417);
xnor UO_1551 (O_1551,N_16103,N_15550);
or UO_1552 (O_1552,N_19872,N_19306);
or UO_1553 (O_1553,N_15851,N_18161);
nand UO_1554 (O_1554,N_18834,N_16805);
and UO_1555 (O_1555,N_18054,N_17480);
or UO_1556 (O_1556,N_17012,N_15255);
or UO_1557 (O_1557,N_19316,N_15326);
nand UO_1558 (O_1558,N_19204,N_15091);
and UO_1559 (O_1559,N_18960,N_15024);
xor UO_1560 (O_1560,N_17981,N_18300);
or UO_1561 (O_1561,N_15231,N_17538);
nand UO_1562 (O_1562,N_15441,N_17534);
or UO_1563 (O_1563,N_16132,N_18080);
or UO_1564 (O_1564,N_17310,N_17499);
and UO_1565 (O_1565,N_19281,N_17066);
or UO_1566 (O_1566,N_17895,N_15955);
nand UO_1567 (O_1567,N_16189,N_17242);
or UO_1568 (O_1568,N_18345,N_17274);
and UO_1569 (O_1569,N_15614,N_15663);
nand UO_1570 (O_1570,N_19044,N_16377);
and UO_1571 (O_1571,N_16595,N_15532);
nor UO_1572 (O_1572,N_16994,N_19280);
or UO_1573 (O_1573,N_18590,N_18497);
or UO_1574 (O_1574,N_19276,N_17325);
nor UO_1575 (O_1575,N_17270,N_19217);
nor UO_1576 (O_1576,N_19328,N_15135);
nor UO_1577 (O_1577,N_16836,N_18278);
or UO_1578 (O_1578,N_19261,N_15563);
and UO_1579 (O_1579,N_19962,N_16779);
and UO_1580 (O_1580,N_18830,N_15763);
nand UO_1581 (O_1581,N_17899,N_17760);
nand UO_1582 (O_1582,N_19848,N_17825);
nand UO_1583 (O_1583,N_19353,N_18229);
xnor UO_1584 (O_1584,N_19442,N_16394);
nor UO_1585 (O_1585,N_15035,N_15464);
nor UO_1586 (O_1586,N_16510,N_17937);
nand UO_1587 (O_1587,N_16108,N_15756);
xor UO_1588 (O_1588,N_15813,N_19314);
or UO_1589 (O_1589,N_17332,N_15511);
nand UO_1590 (O_1590,N_15978,N_15684);
or UO_1591 (O_1591,N_19326,N_18090);
nand UO_1592 (O_1592,N_19311,N_18964);
and UO_1593 (O_1593,N_15420,N_17641);
or UO_1594 (O_1594,N_16882,N_15872);
or UO_1595 (O_1595,N_17660,N_17450);
xnor UO_1596 (O_1596,N_17934,N_16761);
and UO_1597 (O_1597,N_18832,N_17038);
and UO_1598 (O_1598,N_16849,N_16286);
and UO_1599 (O_1599,N_17408,N_19881);
nor UO_1600 (O_1600,N_19479,N_19646);
nor UO_1601 (O_1601,N_17581,N_16289);
xnor UO_1602 (O_1602,N_18235,N_17583);
or UO_1603 (O_1603,N_16297,N_18879);
or UO_1604 (O_1604,N_19874,N_18642);
nor UO_1605 (O_1605,N_16842,N_19378);
and UO_1606 (O_1606,N_19166,N_18530);
nor UO_1607 (O_1607,N_19934,N_16917);
nor UO_1608 (O_1608,N_16283,N_19415);
nand UO_1609 (O_1609,N_18053,N_17701);
nand UO_1610 (O_1610,N_17133,N_19615);
nor UO_1611 (O_1611,N_17261,N_15981);
nor UO_1612 (O_1612,N_15336,N_16102);
nand UO_1613 (O_1613,N_19076,N_19772);
and UO_1614 (O_1614,N_16949,N_17878);
nor UO_1615 (O_1615,N_16806,N_15136);
or UO_1616 (O_1616,N_17086,N_18071);
or UO_1617 (O_1617,N_16272,N_17601);
or UO_1618 (O_1618,N_15287,N_16669);
nand UO_1619 (O_1619,N_15363,N_15319);
and UO_1620 (O_1620,N_16389,N_18107);
xor UO_1621 (O_1621,N_19655,N_19405);
nor UO_1622 (O_1622,N_19602,N_15178);
xnor UO_1623 (O_1623,N_19173,N_16038);
nand UO_1624 (O_1624,N_17858,N_15905);
or UO_1625 (O_1625,N_19210,N_15697);
xnor UO_1626 (O_1626,N_17009,N_18049);
nand UO_1627 (O_1627,N_18455,N_15591);
nor UO_1628 (O_1628,N_18666,N_19470);
nand UO_1629 (O_1629,N_19343,N_16991);
nand UO_1630 (O_1630,N_16441,N_15443);
xnor UO_1631 (O_1631,N_17811,N_18620);
nor UO_1632 (O_1632,N_17627,N_15372);
nor UO_1633 (O_1633,N_17226,N_17881);
nor UO_1634 (O_1634,N_19344,N_18476);
nor UO_1635 (O_1635,N_15553,N_15878);
nand UO_1636 (O_1636,N_18575,N_19290);
nor UO_1637 (O_1637,N_18205,N_17059);
nand UO_1638 (O_1638,N_18733,N_16564);
nand UO_1639 (O_1639,N_18208,N_16034);
nand UO_1640 (O_1640,N_16574,N_18117);
nor UO_1641 (O_1641,N_18969,N_18320);
or UO_1642 (O_1642,N_19299,N_18131);
nor UO_1643 (O_1643,N_19302,N_15984);
or UO_1644 (O_1644,N_18175,N_18132);
and UO_1645 (O_1645,N_16142,N_16323);
nor UO_1646 (O_1646,N_16956,N_16676);
and UO_1647 (O_1647,N_16569,N_16035);
or UO_1648 (O_1648,N_17690,N_15141);
or UO_1649 (O_1649,N_15690,N_18295);
nand UO_1650 (O_1650,N_15625,N_18905);
and UO_1651 (O_1651,N_17068,N_15152);
or UO_1652 (O_1652,N_19037,N_17618);
xor UO_1653 (O_1653,N_16554,N_19961);
and UO_1654 (O_1654,N_15742,N_17429);
nand UO_1655 (O_1655,N_15121,N_16765);
or UO_1656 (O_1656,N_15714,N_18913);
nor UO_1657 (O_1657,N_18141,N_19213);
or UO_1658 (O_1658,N_19757,N_19644);
xor UO_1659 (O_1659,N_19981,N_15659);
nand UO_1660 (O_1660,N_15351,N_19207);
and UO_1661 (O_1661,N_15218,N_15570);
xnor UO_1662 (O_1662,N_17224,N_18893);
and UO_1663 (O_1663,N_19855,N_16055);
or UO_1664 (O_1664,N_15840,N_17137);
and UO_1665 (O_1665,N_16402,N_18425);
nand UO_1666 (O_1666,N_19714,N_15903);
nand UO_1667 (O_1667,N_19906,N_15314);
and UO_1668 (O_1668,N_16426,N_19584);
nor UO_1669 (O_1669,N_19544,N_18499);
or UO_1670 (O_1670,N_17994,N_18991);
or UO_1671 (O_1671,N_15458,N_16514);
xor UO_1672 (O_1672,N_15118,N_19632);
nand UO_1673 (O_1673,N_18483,N_16187);
or UO_1674 (O_1674,N_18865,N_16741);
and UO_1675 (O_1675,N_19882,N_19570);
nand UO_1676 (O_1676,N_15036,N_16597);
nand UO_1677 (O_1677,N_18266,N_19504);
nand UO_1678 (O_1678,N_15843,N_19826);
and UO_1679 (O_1679,N_18268,N_17506);
or UO_1680 (O_1680,N_17407,N_15335);
nand UO_1681 (O_1681,N_18434,N_15312);
nor UO_1682 (O_1682,N_18860,N_16500);
and UO_1683 (O_1683,N_17675,N_16384);
nand UO_1684 (O_1684,N_16455,N_16983);
nand UO_1685 (O_1685,N_16603,N_18571);
and UO_1686 (O_1686,N_15368,N_17944);
and UO_1687 (O_1687,N_18608,N_18876);
or UO_1688 (O_1688,N_19765,N_18775);
nand UO_1689 (O_1689,N_17647,N_17525);
nand UO_1690 (O_1690,N_17673,N_15467);
xor UO_1691 (O_1691,N_16560,N_18452);
nand UO_1692 (O_1692,N_17014,N_18934);
or UO_1693 (O_1693,N_16031,N_17816);
nor UO_1694 (O_1694,N_16343,N_16365);
nor UO_1695 (O_1695,N_19266,N_17003);
and UO_1696 (O_1696,N_16025,N_16220);
nand UO_1697 (O_1697,N_15734,N_17333);
or UO_1698 (O_1698,N_15508,N_17371);
nand UO_1699 (O_1699,N_18906,N_18771);
nand UO_1700 (O_1700,N_15522,N_19858);
and UO_1701 (O_1701,N_15825,N_19592);
nand UO_1702 (O_1702,N_16526,N_17025);
nor UO_1703 (O_1703,N_17723,N_15902);
and UO_1704 (O_1704,N_15360,N_17613);
xor UO_1705 (O_1705,N_18856,N_17300);
nor UO_1706 (O_1706,N_17289,N_16391);
nand UO_1707 (O_1707,N_17434,N_17349);
nor UO_1708 (O_1708,N_17843,N_19777);
nor UO_1709 (O_1709,N_16090,N_16633);
nand UO_1710 (O_1710,N_19616,N_18753);
nand UO_1711 (O_1711,N_18373,N_16942);
nor UO_1712 (O_1712,N_15107,N_19130);
xor UO_1713 (O_1713,N_15358,N_19121);
or UO_1714 (O_1714,N_18407,N_16412);
nand UO_1715 (O_1715,N_19032,N_18539);
nor UO_1716 (O_1716,N_17854,N_19675);
nor UO_1717 (O_1717,N_15695,N_15866);
nand UO_1718 (O_1718,N_16666,N_16223);
nand UO_1719 (O_1719,N_17745,N_19914);
or UO_1720 (O_1720,N_17886,N_18350);
and UO_1721 (O_1721,N_19817,N_15549);
nor UO_1722 (O_1722,N_17541,N_19025);
and UO_1723 (O_1723,N_16723,N_18611);
or UO_1724 (O_1724,N_17063,N_17171);
or UO_1725 (O_1725,N_17781,N_19811);
xnor UO_1726 (O_1726,N_19559,N_16249);
and UO_1727 (O_1727,N_19993,N_17237);
nor UO_1728 (O_1728,N_16089,N_18163);
nand UO_1729 (O_1729,N_16069,N_19998);
nor UO_1730 (O_1730,N_19193,N_16091);
or UO_1731 (O_1731,N_18484,N_16513);
and UO_1732 (O_1732,N_19952,N_18298);
nand UO_1733 (O_1733,N_15037,N_17628);
nand UO_1734 (O_1734,N_19144,N_17721);
and UO_1735 (O_1735,N_18121,N_16881);
nor UO_1736 (O_1736,N_16294,N_17571);
nor UO_1737 (O_1737,N_17530,N_19727);
nand UO_1738 (O_1738,N_15468,N_19688);
nand UO_1739 (O_1739,N_19525,N_15921);
or UO_1740 (O_1740,N_15925,N_16802);
xnor UO_1741 (O_1741,N_17579,N_18852);
nand UO_1742 (O_1742,N_16493,N_18671);
nand UO_1743 (O_1743,N_18872,N_18336);
nand UO_1744 (O_1744,N_15747,N_16234);
or UO_1745 (O_1745,N_16585,N_18955);
nor UO_1746 (O_1746,N_17567,N_19807);
nor UO_1747 (O_1747,N_17394,N_17709);
nor UO_1748 (O_1748,N_17824,N_19028);
or UO_1749 (O_1749,N_15648,N_17037);
and UO_1750 (O_1750,N_19505,N_17460);
or UO_1751 (O_1751,N_17609,N_17718);
nand UO_1752 (O_1752,N_17524,N_18661);
nand UO_1753 (O_1753,N_15269,N_16371);
and UO_1754 (O_1754,N_19014,N_16157);
or UO_1755 (O_1755,N_16876,N_16884);
or UO_1756 (O_1756,N_16277,N_16388);
and UO_1757 (O_1757,N_17061,N_15557);
nand UO_1758 (O_1758,N_17228,N_15682);
or UO_1759 (O_1759,N_17831,N_16931);
and UO_1760 (O_1760,N_19497,N_17527);
or UO_1761 (O_1761,N_17610,N_16021);
or UO_1762 (O_1762,N_16896,N_19045);
and UO_1763 (O_1763,N_17914,N_18451);
nand UO_1764 (O_1764,N_19315,N_15021);
nor UO_1765 (O_1765,N_18426,N_18288);
or UO_1766 (O_1766,N_15499,N_17540);
and UO_1767 (O_1767,N_17600,N_16355);
nand UO_1768 (O_1768,N_15552,N_17343);
nand UO_1769 (O_1769,N_19837,N_19401);
nand UO_1770 (O_1770,N_15082,N_15913);
xor UO_1771 (O_1771,N_17578,N_15920);
nand UO_1772 (O_1772,N_19110,N_19832);
and UO_1773 (O_1773,N_15098,N_19560);
nand UO_1774 (O_1774,N_18245,N_19867);
nand UO_1775 (O_1775,N_17017,N_16232);
nand UO_1776 (O_1776,N_18745,N_15054);
or UO_1777 (O_1777,N_16121,N_19113);
xnor UO_1778 (O_1778,N_15079,N_19937);
and UO_1779 (O_1779,N_19017,N_18851);
and UO_1780 (O_1780,N_18791,N_16276);
and UO_1781 (O_1781,N_16287,N_17572);
nand UO_1782 (O_1782,N_18352,N_15888);
and UO_1783 (O_1783,N_16964,N_16950);
nor UO_1784 (O_1784,N_17793,N_15222);
and UO_1785 (O_1785,N_16923,N_18765);
or UO_1786 (O_1786,N_18168,N_18013);
nand UO_1787 (O_1787,N_19595,N_17359);
and UO_1788 (O_1788,N_16982,N_19728);
nand UO_1789 (O_1789,N_17770,N_16700);
and UO_1790 (O_1790,N_15907,N_18411);
or UO_1791 (O_1791,N_19850,N_19098);
nand UO_1792 (O_1792,N_15871,N_19384);
xor UO_1793 (O_1793,N_17777,N_17892);
nor UO_1794 (O_1794,N_15215,N_17402);
or UO_1795 (O_1795,N_15900,N_17946);
and UO_1796 (O_1796,N_16057,N_17838);
or UO_1797 (O_1797,N_19254,N_18136);
xor UO_1798 (O_1798,N_17153,N_18213);
or UO_1799 (O_1799,N_16787,N_18442);
nand UO_1800 (O_1800,N_15365,N_16164);
nor UO_1801 (O_1801,N_19047,N_17661);
xnor UO_1802 (O_1802,N_15624,N_15017);
or UO_1803 (O_1803,N_16345,N_19884);
nand UO_1804 (O_1804,N_17385,N_17373);
and UO_1805 (O_1805,N_16699,N_18079);
nand UO_1806 (O_1806,N_18649,N_17496);
or UO_1807 (O_1807,N_15242,N_18748);
nor UO_1808 (O_1808,N_18237,N_18346);
nor UO_1809 (O_1809,N_17912,N_15248);
or UO_1810 (O_1810,N_19109,N_18017);
xnor UO_1811 (O_1811,N_18094,N_18833);
and UO_1812 (O_1812,N_19183,N_17100);
nor UO_1813 (O_1813,N_19561,N_19669);
nand UO_1814 (O_1814,N_18887,N_16463);
nand UO_1815 (O_1815,N_15352,N_17219);
and UO_1816 (O_1816,N_18994,N_19128);
nor UO_1817 (O_1817,N_19475,N_19518);
or UO_1818 (O_1818,N_16339,N_16922);
and UO_1819 (O_1819,N_15321,N_15633);
nor UO_1820 (O_1820,N_16932,N_18450);
or UO_1821 (O_1821,N_17963,N_18154);
and UO_1822 (O_1822,N_18912,N_19685);
nand UO_1823 (O_1823,N_18957,N_16155);
or UO_1824 (O_1824,N_18869,N_15877);
nor UO_1825 (O_1825,N_17103,N_19626);
and UO_1826 (O_1826,N_18980,N_15641);
nand UO_1827 (O_1827,N_18680,N_19400);
nand UO_1828 (O_1828,N_16138,N_17305);
xnor UO_1829 (O_1829,N_19451,N_19147);
or UO_1830 (O_1830,N_17565,N_18632);
nor UO_1831 (O_1831,N_18724,N_17519);
and UO_1832 (O_1832,N_16314,N_19814);
nor UO_1833 (O_1833,N_18406,N_17885);
nor UO_1834 (O_1834,N_15858,N_15619);
nand UO_1835 (O_1835,N_17116,N_15025);
or UO_1836 (O_1836,N_17205,N_16053);
or UO_1837 (O_1837,N_17384,N_18580);
xor UO_1838 (O_1838,N_19445,N_16331);
or UO_1839 (O_1839,N_15972,N_15074);
or UO_1840 (O_1840,N_15967,N_17202);
and UO_1841 (O_1841,N_18155,N_16551);
nand UO_1842 (O_1842,N_17485,N_19516);
and UO_1843 (O_1843,N_16041,N_17406);
nor UO_1844 (O_1844,N_17334,N_16459);
nor UO_1845 (O_1845,N_17988,N_19859);
nand UO_1846 (O_1846,N_19523,N_17543);
or UO_1847 (O_1847,N_17081,N_17007);
and UO_1848 (O_1848,N_16073,N_19713);
or UO_1849 (O_1849,N_15020,N_19264);
nand UO_1850 (O_1850,N_19731,N_15644);
or UO_1851 (O_1851,N_18197,N_19022);
xnor UO_1852 (O_1852,N_15653,N_18521);
nand UO_1853 (O_1853,N_15775,N_19749);
xnor UO_1854 (O_1854,N_17364,N_16709);
xnor UO_1855 (O_1855,N_17308,N_19012);
nand UO_1856 (O_1856,N_16239,N_19657);
nand UO_1857 (O_1857,N_16024,N_19635);
nor UO_1858 (O_1858,N_19589,N_19667);
nand UO_1859 (O_1859,N_17144,N_18042);
nor UO_1860 (O_1860,N_18195,N_16733);
nand UO_1861 (O_1861,N_18681,N_17419);
xor UO_1862 (O_1862,N_16869,N_15083);
or UO_1863 (O_1863,N_18677,N_19813);
nor UO_1864 (O_1864,N_17126,N_16871);
nor UO_1865 (O_1865,N_16433,N_18395);
nand UO_1866 (O_1866,N_19282,N_17036);
xor UO_1867 (O_1867,N_16621,N_18764);
nor UO_1868 (O_1868,N_19596,N_17381);
and UO_1869 (O_1869,N_18200,N_18072);
and UO_1870 (O_1870,N_17405,N_19529);
nor UO_1871 (O_1871,N_19991,N_17417);
nand UO_1872 (O_1872,N_19831,N_16646);
or UO_1873 (O_1873,N_15401,N_17401);
and UO_1874 (O_1874,N_17533,N_15430);
or UO_1875 (O_1875,N_16415,N_18873);
or UO_1876 (O_1876,N_18918,N_19329);
and UO_1877 (O_1877,N_17073,N_18892);
and UO_1878 (O_1878,N_16558,N_17775);
nor UO_1879 (O_1879,N_18096,N_17604);
nor UO_1880 (O_1880,N_16128,N_19134);
or UO_1881 (O_1881,N_16369,N_17563);
and UO_1882 (O_1882,N_19750,N_18183);
or UO_1883 (O_1883,N_17684,N_15173);
xor UO_1884 (O_1884,N_15590,N_19995);
and UO_1885 (O_1885,N_16756,N_15318);
and UO_1886 (O_1886,N_18720,N_18325);
and UO_1887 (O_1887,N_16231,N_18196);
or UO_1888 (O_1888,N_18939,N_16151);
and UO_1889 (O_1889,N_19325,N_15732);
nand UO_1890 (O_1890,N_15032,N_19898);
and UO_1891 (O_1891,N_16163,N_18321);
nor UO_1892 (O_1892,N_17212,N_17909);
nand UO_1893 (O_1893,N_15239,N_17010);
nor UO_1894 (O_1894,N_17463,N_18048);
nor UO_1895 (O_1895,N_17796,N_16440);
or UO_1896 (O_1896,N_17400,N_18275);
or UO_1897 (O_1897,N_17449,N_15718);
or UO_1898 (O_1898,N_19844,N_15018);
nor UO_1899 (O_1899,N_16399,N_19460);
or UO_1900 (O_1900,N_19755,N_18188);
or UO_1901 (O_1901,N_17026,N_18430);
xnor UO_1902 (O_1902,N_19823,N_18456);
and UO_1903 (O_1903,N_15527,N_15317);
and UO_1904 (O_1904,N_16885,N_17753);
nor UO_1905 (O_1905,N_15569,N_16550);
nor UO_1906 (O_1906,N_16967,N_15503);
and UO_1907 (O_1907,N_17631,N_16934);
or UO_1908 (O_1908,N_18246,N_17018);
or UO_1909 (O_1909,N_16212,N_15933);
nor UO_1910 (O_1910,N_15161,N_18798);
and UO_1911 (O_1911,N_18751,N_18172);
nor UO_1912 (O_1912,N_15436,N_18952);
nor UO_1913 (O_1913,N_16903,N_17290);
nor UO_1914 (O_1914,N_18178,N_18146);
and UO_1915 (O_1915,N_17393,N_19218);
nor UO_1916 (O_1916,N_18362,N_17593);
nor UO_1917 (O_1917,N_15879,N_18400);
nor UO_1918 (O_1918,N_15439,N_18114);
or UO_1919 (O_1919,N_16201,N_16224);
or UO_1920 (O_1920,N_18601,N_18333);
or UO_1921 (O_1921,N_19269,N_15085);
or UO_1922 (O_1922,N_15316,N_18704);
and UO_1923 (O_1923,N_18809,N_16176);
nand UO_1924 (O_1924,N_15410,N_18585);
nor UO_1925 (O_1925,N_19068,N_15010);
nor UO_1926 (O_1926,N_17592,N_15384);
nand UO_1927 (O_1927,N_18624,N_18159);
or UO_1928 (O_1928,N_18142,N_17119);
and UO_1929 (O_1929,N_18029,N_17047);
xor UO_1930 (O_1930,N_17715,N_19118);
nand UO_1931 (O_1931,N_18359,N_17674);
nand UO_1932 (O_1932,N_15058,N_17154);
and UO_1933 (O_1933,N_16217,N_19107);
nor UO_1934 (O_1934,N_17184,N_15666);
nor UO_1935 (O_1935,N_15701,N_15119);
nand UO_1936 (O_1936,N_16046,N_17348);
or UO_1937 (O_1937,N_15076,N_17396);
or UO_1938 (O_1938,N_18050,N_17241);
and UO_1939 (O_1939,N_17004,N_15964);
or UO_1940 (O_1940,N_18667,N_17676);
nor UO_1941 (O_1941,N_17096,N_16860);
and UO_1942 (O_1942,N_15792,N_16414);
xor UO_1943 (O_1943,N_16858,N_15924);
nor UO_1944 (O_1944,N_15162,N_19861);
or UO_1945 (O_1945,N_15528,N_18553);
or UO_1946 (O_1946,N_16357,N_17456);
xnor UO_1947 (O_1947,N_16156,N_15026);
and UO_1948 (O_1948,N_15479,N_17461);
and UO_1949 (O_1949,N_19873,N_16378);
or UO_1950 (O_1950,N_19133,N_17855);
nand UO_1951 (O_1951,N_16590,N_15609);
and UO_1952 (O_1952,N_19298,N_19279);
nand UO_1953 (O_1953,N_19676,N_19703);
xnor UO_1954 (O_1954,N_19563,N_17207);
and UO_1955 (O_1955,N_17320,N_19639);
and UO_1956 (O_1956,N_19892,N_18160);
xnor UO_1957 (O_1957,N_17648,N_19975);
xor UO_1958 (O_1958,N_18741,N_17372);
xnor UO_1959 (O_1959,N_16712,N_16456);
and UO_1960 (O_1960,N_17670,N_16799);
xor UO_1961 (O_1961,N_16984,N_17516);
or UO_1962 (O_1962,N_16471,N_18297);
xnor UO_1963 (O_1963,N_15189,N_17894);
xor UO_1964 (O_1964,N_16467,N_15513);
and UO_1965 (O_1965,N_18392,N_19853);
nand UO_1966 (O_1966,N_18466,N_18673);
nor UO_1967 (O_1967,N_15123,N_19628);
nor UO_1968 (O_1968,N_16831,N_18899);
nand UO_1969 (O_1969,N_15899,N_17865);
and UO_1970 (O_1970,N_16332,N_15558);
xor UO_1971 (O_1971,N_15126,N_19927);
nor UO_1972 (O_1972,N_16773,N_19495);
nor UO_1973 (O_1973,N_19010,N_16745);
or UO_1974 (O_1974,N_18339,N_18788);
or UO_1975 (O_1975,N_15606,N_17115);
and UO_1976 (O_1976,N_16359,N_17953);
xnor UO_1977 (O_1977,N_19411,N_17819);
nor UO_1978 (O_1978,N_17751,N_19219);
or UO_1979 (O_1979,N_15554,N_16897);
xnor UO_1980 (O_1980,N_18240,N_16472);
nor UO_1981 (O_1981,N_15206,N_15398);
and UO_1982 (O_1982,N_19783,N_19359);
nand UO_1983 (O_1983,N_15496,N_15271);
nor UO_1984 (O_1984,N_18739,N_16742);
nor UO_1985 (O_1985,N_15819,N_16604);
or UO_1986 (O_1986,N_15099,N_19661);
nor UO_1987 (O_1987,N_17011,N_19145);
nor UO_1988 (O_1988,N_19332,N_17828);
nor UO_1989 (O_1989,N_15873,N_18118);
or UO_1990 (O_1990,N_19957,N_19953);
nand UO_1991 (O_1991,N_15587,N_17094);
or UO_1992 (O_1992,N_17817,N_15950);
nand UO_1993 (O_1993,N_15115,N_19636);
nand UO_1994 (O_1994,N_17054,N_18216);
or UO_1995 (O_1995,N_15537,N_16753);
nand UO_1996 (O_1996,N_16215,N_18243);
nor UO_1997 (O_1997,N_17772,N_18469);
or UO_1998 (O_1998,N_15296,N_18388);
nor UO_1999 (O_1999,N_16784,N_16313);
nand UO_2000 (O_2000,N_17344,N_18940);
nor UO_2001 (O_2001,N_15798,N_15448);
or UO_2002 (O_2002,N_16134,N_19289);
nand UO_2003 (O_2003,N_15375,N_15341);
nand UO_2004 (O_2004,N_15965,N_19362);
and UO_2005 (O_2005,N_19594,N_18903);
and UO_2006 (O_2006,N_18592,N_18562);
and UO_2007 (O_2007,N_17015,N_17546);
or UO_2008 (O_2008,N_15876,N_15774);
and UO_2009 (O_2009,N_17479,N_19347);
or UO_2010 (O_2010,N_19573,N_16518);
or UO_2011 (O_2011,N_19228,N_17264);
nand UO_2012 (O_2012,N_19748,N_19227);
nor UO_2013 (O_2013,N_15004,N_18014);
nand UO_2014 (O_2014,N_18326,N_15923);
nand UO_2015 (O_2015,N_17594,N_18941);
or UO_2016 (O_2016,N_19444,N_19273);
and UO_2017 (O_2017,N_16834,N_19223);
nand UO_2018 (O_2018,N_18895,N_17218);
xor UO_2019 (O_2019,N_17619,N_16264);
or UO_2020 (O_2020,N_19706,N_15540);
nor UO_2021 (O_2021,N_17589,N_15112);
nand UO_2022 (O_2022,N_19225,N_17331);
xnor UO_2023 (O_2023,N_17355,N_18305);
nor UO_2024 (O_2024,N_16019,N_19862);
nand UO_2025 (O_2025,N_16933,N_17904);
nand UO_2026 (O_2026,N_18270,N_15237);
nand UO_2027 (O_2027,N_19680,N_19382);
xnor UO_2028 (O_2028,N_18364,N_16397);
and UO_2029 (O_2029,N_17560,N_15583);
or UO_2030 (O_2030,N_19165,N_18602);
and UO_2031 (O_2031,N_15047,N_19880);
and UO_2032 (O_2032,N_16804,N_16186);
nand UO_2033 (O_2033,N_19200,N_18100);
and UO_2034 (O_2034,N_18914,N_15548);
nor UO_2035 (O_2035,N_16835,N_19959);
nand UO_2036 (O_2036,N_15450,N_19455);
xor UO_2037 (O_2037,N_19158,N_18421);
nand UO_2038 (O_2038,N_19322,N_18276);
or UO_2039 (O_2039,N_18112,N_17748);
nand UO_2040 (O_2040,N_16622,N_17072);
and UO_2041 (O_2041,N_16006,N_15683);
and UO_2042 (O_2042,N_17681,N_19235);
or UO_2043 (O_2043,N_16058,N_18782);
or UO_2044 (O_2044,N_15357,N_16113);
and UO_2045 (O_2045,N_16437,N_16026);
and UO_2046 (O_2046,N_16874,N_16605);
nand UO_2047 (O_2047,N_17549,N_18273);
nand UO_2048 (O_2048,N_18091,N_16575);
or UO_2049 (O_2049,N_19764,N_17318);
and UO_2050 (O_2050,N_18045,N_18723);
nor UO_2051 (O_2051,N_18982,N_15698);
or UO_2052 (O_2052,N_19416,N_17421);
nand UO_2053 (O_2053,N_16588,N_19540);
nand UO_2054 (O_2054,N_18302,N_15711);
and UO_2055 (O_2055,N_19736,N_16748);
nor UO_2056 (O_2056,N_16381,N_16985);
nand UO_2057 (O_2057,N_18259,N_18459);
and UO_2058 (O_2058,N_19666,N_18348);
and UO_2059 (O_2059,N_16370,N_16030);
and UO_2060 (O_2060,N_19641,N_18074);
and UO_2061 (O_2061,N_19893,N_16637);
nand UO_2062 (O_2062,N_19683,N_18209);
nand UO_2063 (O_2063,N_18093,N_18700);
nor UO_2064 (O_2064,N_16485,N_16322);
or UO_2065 (O_2065,N_18156,N_19484);
nor UO_2066 (O_2066,N_18447,N_18170);
xor UO_2067 (O_2067,N_19980,N_18909);
and UO_2068 (O_2068,N_19388,N_16927);
nor UO_2069 (O_2069,N_15610,N_15275);
nand UO_2070 (O_2070,N_17194,N_16141);
and UO_2071 (O_2071,N_18383,N_16432);
or UO_2072 (O_2072,N_15373,N_17231);
nand UO_2073 (O_2073,N_16853,N_18973);
and UO_2074 (O_2074,N_15270,N_17105);
nand UO_2075 (O_2075,N_15534,N_17163);
nor UO_2076 (O_2076,N_15238,N_17034);
nor UO_2077 (O_2077,N_15700,N_16425);
nand UO_2078 (O_2078,N_15469,N_15006);
and UO_2079 (O_2079,N_15829,N_18618);
nand UO_2080 (O_2080,N_15757,N_15388);
nand UO_2081 (O_2081,N_18815,N_15969);
xor UO_2082 (O_2082,N_17272,N_15958);
and UO_2083 (O_2083,N_15892,N_15796);
and UO_2084 (O_2084,N_17001,N_19389);
nand UO_2085 (O_2085,N_15470,N_19421);
nor UO_2086 (O_2086,N_15783,N_19459);
and UO_2087 (O_2087,N_18040,N_19835);
nor UO_2088 (O_2088,N_16393,N_15818);
nand UO_2089 (O_2089,N_17472,N_15715);
nor UO_2090 (O_2090,N_19341,N_19776);
and UO_2091 (O_2091,N_19339,N_16721);
nand UO_2092 (O_2092,N_18368,N_18062);
or UO_2093 (O_2093,N_18331,N_19432);
nand UO_2094 (O_2094,N_16137,N_16166);
nand UO_2095 (O_2095,N_19532,N_17253);
xnor UO_2096 (O_2096,N_15865,N_16087);
nor UO_2097 (O_2097,N_15710,N_18636);
or UO_2098 (O_2098,N_15230,N_15657);
nand UO_2099 (O_2099,N_18186,N_18638);
and UO_2100 (O_2100,N_15462,N_19674);
nand UO_2101 (O_2101,N_15545,N_15013);
and UO_2102 (O_2102,N_15092,N_18227);
nand UO_2103 (O_2103,N_18201,N_18396);
or UO_2104 (O_2104,N_19907,N_18881);
nor UO_2105 (O_2105,N_19805,N_19819);
nor UO_2106 (O_2106,N_18538,N_19720);
or UO_2107 (O_2107,N_18871,N_19458);
and UO_2108 (O_2108,N_18855,N_15407);
nor UO_2109 (O_2109,N_17959,N_15226);
and UO_2110 (O_2110,N_17088,N_17216);
or UO_2111 (O_2111,N_17159,N_16062);
and UO_2112 (O_2112,N_17341,N_19865);
nand UO_2113 (O_2113,N_17989,N_15253);
or UO_2114 (O_2114,N_16064,N_18389);
or UO_2115 (O_2115,N_16011,N_15561);
or UO_2116 (O_2116,N_15719,N_16902);
or UO_2117 (O_2117,N_17113,N_17779);
and UO_2118 (O_2118,N_18277,N_15440);
nand UO_2119 (O_2119,N_15343,N_15890);
nor UO_2120 (O_2120,N_15880,N_19249);
xnor UO_2121 (O_2121,N_16431,N_17978);
nor UO_2122 (O_2122,N_15293,N_16747);
nand UO_2123 (O_2123,N_18950,N_15505);
or UO_2124 (O_2124,N_19522,N_16682);
nor UO_2125 (O_2125,N_15805,N_17997);
and UO_2126 (O_2126,N_16845,N_16410);
nor UO_2127 (O_2127,N_18309,N_15707);
nor UO_2128 (O_2128,N_19761,N_16110);
nand UO_2129 (O_2129,N_15823,N_16579);
and UO_2130 (O_2130,N_17632,N_17554);
or UO_2131 (O_2131,N_17590,N_17293);
xor UO_2132 (O_2132,N_16193,N_15582);
or UO_2133 (O_2133,N_15996,N_18811);
and UO_2134 (O_2134,N_16648,N_16190);
nand UO_2135 (O_2135,N_16348,N_18022);
nand UO_2136 (O_2136,N_16442,N_15075);
and UO_2137 (O_2137,N_15676,N_15961);
and UO_2138 (O_2138,N_15016,N_18187);
nand UO_2139 (O_2139,N_17083,N_19521);
and UO_2140 (O_2140,N_17985,N_18242);
or UO_2141 (O_2141,N_19007,N_19448);
nor UO_2142 (O_2142,N_19790,N_16144);
nor UO_2143 (O_2143,N_15452,N_18598);
xnor UO_2144 (O_2144,N_17195,N_19462);
xnor UO_2145 (O_2145,N_16775,N_18740);
nor UO_2146 (O_2146,N_18055,N_16205);
and UO_2147 (O_2147,N_15543,N_19673);
nor UO_2148 (O_2148,N_15836,N_18420);
and UO_2149 (O_2149,N_16117,N_16430);
nand UO_2150 (O_2150,N_15380,N_18772);
nand UO_2151 (O_2151,N_18508,N_17708);
nand UO_2152 (O_2152,N_19732,N_19625);
nand UO_2153 (O_2153,N_17999,N_18804);
or UO_2154 (O_2154,N_19364,N_18380);
nand UO_2155 (O_2155,N_19587,N_18385);
nor UO_2156 (O_2156,N_15944,N_16868);
xor UO_2157 (O_2157,N_17303,N_18365);
nand UO_2158 (O_2158,N_19224,N_18878);
nor UO_2159 (O_2159,N_16846,N_19804);
nor UO_2160 (O_2160,N_18846,N_19809);
nor UO_2161 (O_2161,N_15667,N_16226);
nand UO_2162 (O_2162,N_16948,N_19248);
nand UO_2163 (O_2163,N_19956,N_18177);
or UO_2164 (O_2164,N_18332,N_17602);
nor UO_2165 (O_2165,N_18151,N_17118);
and UO_2166 (O_2166,N_15860,N_15193);
nand UO_2167 (O_2167,N_18097,N_18706);
nand UO_2168 (O_2168,N_18840,N_16616);
nand UO_2169 (O_2169,N_19284,N_16451);
and UO_2170 (O_2170,N_15171,N_18077);
nor UO_2171 (O_2171,N_19108,N_16200);
xnor UO_2172 (O_2172,N_15556,N_17245);
nor UO_2173 (O_2173,N_18987,N_15809);
or UO_2174 (O_2174,N_15002,N_19263);
or UO_2175 (O_2175,N_16767,N_18540);
nand UO_2176 (O_2176,N_16047,N_16815);
or UO_2177 (O_2177,N_18330,N_16023);
nand UO_2178 (O_2178,N_17625,N_15951);
xor UO_2179 (O_2179,N_17815,N_17431);
and UO_2180 (O_2180,N_16253,N_19357);
nor UO_2181 (O_2181,N_18687,N_16061);
nor UO_2182 (O_2182,N_16650,N_16878);
or UO_2183 (O_2183,N_19377,N_16454);
nand UO_2184 (O_2184,N_19394,N_18185);
nor UO_2185 (O_2185,N_18812,N_16999);
or UO_2186 (O_2186,N_17362,N_19461);
or UO_2187 (O_2187,N_15390,N_16609);
nor UO_2188 (O_2188,N_19139,N_16535);
and UO_2189 (O_2189,N_19549,N_17597);
nor UO_2190 (O_2190,N_16599,N_17032);
nor UO_2191 (O_2191,N_16303,N_19059);
and UO_2192 (O_2192,N_15736,N_16681);
xor UO_2193 (O_2193,N_19331,N_19066);
or UO_2194 (O_2194,N_17700,N_17889);
and UO_2195 (O_2195,N_18752,N_15109);
and UO_2196 (O_2196,N_16333,N_15111);
nand UO_2197 (O_2197,N_16293,N_16492);
and UO_2198 (O_2198,N_17773,N_19494);
or UO_2199 (O_2199,N_15086,N_17179);
and UO_2200 (O_2200,N_19665,N_15612);
or UO_2201 (O_2201,N_19829,N_19182);
or UO_2202 (O_2202,N_19797,N_16065);
nand UO_2203 (O_2203,N_19506,N_16396);
and UO_2204 (O_2204,N_18933,N_16829);
nor UO_2205 (O_2205,N_19913,N_17659);
or UO_2206 (O_2206,N_19203,N_16400);
xor UO_2207 (O_2207,N_15041,N_16042);
nand UO_2208 (O_2208,N_16921,N_18335);
and UO_2209 (O_2209,N_16995,N_18629);
xor UO_2210 (O_2210,N_17285,N_17413);
nor UO_2211 (O_2211,N_15623,N_19456);
xnor UO_2212 (O_2212,N_19916,N_19588);
nor UO_2213 (O_2213,N_17972,N_16005);
nor UO_2214 (O_2214,N_17039,N_17654);
or UO_2215 (O_2215,N_19077,N_17568);
and UO_2216 (O_2216,N_19114,N_16071);
xor UO_2217 (O_2217,N_17823,N_18140);
and UO_2218 (O_2218,N_19839,N_15917);
and UO_2219 (O_2219,N_17110,N_18847);
and UO_2220 (O_2220,N_15990,N_15524);
nor UO_2221 (O_2221,N_15397,N_17919);
xnor UO_2222 (O_2222,N_16972,N_17432);
or UO_2223 (O_2223,N_15217,N_19358);
or UO_2224 (O_2224,N_18643,N_18849);
nand UO_2225 (O_2225,N_17553,N_17136);
nor UO_2226 (O_2226,N_19779,N_18428);
and UO_2227 (O_2227,N_15812,N_15101);
nand UO_2228 (O_2228,N_19234,N_16198);
and UO_2229 (O_2229,N_18313,N_17577);
and UO_2230 (O_2230,N_16242,N_19503);
nor UO_2231 (O_2231,N_19058,N_15762);
or UO_2232 (O_2232,N_16109,N_15356);
xnor UO_2233 (O_2233,N_19738,N_16664);
or UO_2234 (O_2234,N_17621,N_15807);
and UO_2235 (O_2235,N_15023,N_16652);
nor UO_2236 (O_2236,N_16327,N_18394);
nand UO_2237 (O_2237,N_15613,N_17987);
nor UO_2238 (O_2238,N_16655,N_15784);
and UO_2239 (O_2239,N_15794,N_16954);
or UO_2240 (O_2240,N_15883,N_17916);
and UO_2241 (O_2241,N_18152,N_16796);
or UO_2242 (O_2242,N_15463,N_19242);
or UO_2243 (O_2243,N_19268,N_16649);
nor UO_2244 (O_2244,N_17918,N_15629);
or UO_2245 (O_2245,N_15651,N_16645);
and UO_2246 (O_2246,N_15962,N_18579);
or UO_2247 (O_2247,N_18583,N_16807);
or UO_2248 (O_2248,N_19417,N_19211);
or UO_2249 (O_2249,N_18115,N_17246);
and UO_2250 (O_2250,N_18981,N_17905);
nor UO_2251 (O_2251,N_19928,N_16373);
nand UO_2252 (O_2252,N_19342,N_16968);
nor UO_2253 (O_2253,N_15277,N_16675);
or UO_2254 (O_2254,N_19157,N_18257);
xnor UO_2255 (O_2255,N_16961,N_17976);
nor UO_2256 (O_2256,N_18993,N_15937);
nor UO_2257 (O_2257,N_19354,N_19412);
and UO_2258 (O_2258,N_18445,N_15566);
nor UO_2259 (O_2259,N_15535,N_18264);
or UO_2260 (O_2260,N_17296,N_17031);
nand UO_2261 (O_2261,N_17669,N_15298);
nand UO_2262 (O_2262,N_19915,N_19538);
and UO_2263 (O_2263,N_18020,N_18559);
and UO_2264 (O_2264,N_15349,N_16228);
xor UO_2265 (O_2265,N_17481,N_16839);
nand UO_2266 (O_2266,N_16478,N_16196);
nand UO_2267 (O_2267,N_18423,N_17080);
and UO_2268 (O_2268,N_17875,N_19682);
or UO_2269 (O_2269,N_18181,N_15046);
or UO_2270 (O_2270,N_19300,N_19305);
and UO_2271 (O_2271,N_15935,N_18247);
nand UO_2272 (O_2272,N_17181,N_16501);
or UO_2273 (O_2273,N_15677,N_17252);
nor UO_2274 (O_2274,N_17733,N_19681);
nor UO_2275 (O_2275,N_15605,N_17851);
and UO_2276 (O_2276,N_15538,N_19564);
and UO_2277 (O_2277,N_18777,N_16246);
or UO_2278 (O_2278,N_18541,N_16216);
nand UO_2279 (O_2279,N_19510,N_16446);
nand UO_2280 (O_2280,N_19935,N_17071);
or UO_2281 (O_2281,N_18875,N_17139);
or UO_2282 (O_2282,N_19016,N_16498);
xor UO_2283 (O_2283,N_19815,N_18797);
and UO_2284 (O_2284,N_16838,N_18238);
nor UO_2285 (O_2285,N_19740,N_16497);
or UO_2286 (O_2286,N_16284,N_17152);
nor UO_2287 (O_2287,N_17706,N_17279);
xnor UO_2288 (O_2288,N_17651,N_19945);
or UO_2289 (O_2289,N_17374,N_17574);
or UO_2290 (O_2290,N_16129,N_16350);
nor UO_2291 (O_2291,N_17614,N_19006);
and UO_2292 (O_2292,N_15060,N_17941);
and UO_2293 (O_2293,N_16460,N_16076);
or UO_2294 (O_2294,N_17183,N_19979);
nor UO_2295 (O_2295,N_18985,N_17335);
nor UO_2296 (O_2296,N_16406,N_18157);
nand UO_2297 (O_2297,N_19965,N_17399);
xnor UO_2298 (O_2298,N_16423,N_17805);
and UO_2299 (O_2299,N_15471,N_16387);
or UO_2300 (O_2300,N_18831,N_18889);
xnor UO_2301 (O_2301,N_15712,N_19001);
nand UO_2302 (O_2302,N_19418,N_17013);
or UO_2303 (O_2303,N_15281,N_19167);
and UO_2304 (O_2304,N_15820,N_15143);
or UO_2305 (O_2305,N_15758,N_17330);
nand UO_2306 (O_2306,N_19226,N_15051);
nand UO_2307 (O_2307,N_19160,N_16050);
xnor UO_2308 (O_2308,N_15706,N_15936);
nand UO_2309 (O_2309,N_15804,N_17993);
nor UO_2310 (O_2310,N_15234,N_15149);
and UO_2311 (O_2311,N_15884,N_15204);
or UO_2312 (O_2312,N_17926,N_19550);
xnor UO_2313 (O_2313,N_18549,N_18516);
nand UO_2314 (O_2314,N_18607,N_16740);
nor UO_2315 (O_2315,N_15769,N_17922);
and UO_2316 (O_2316,N_17829,N_17151);
or UO_2317 (O_2317,N_15568,N_16443);
nand UO_2318 (O_2318,N_17650,N_16895);
nor UO_2319 (O_2319,N_18843,N_17764);
nor UO_2320 (O_2320,N_16777,N_17158);
or UO_2321 (O_2321,N_18082,N_17521);
nor UO_2322 (O_2322,N_19309,N_16546);
nand UO_2323 (O_2323,N_15421,N_18338);
and UO_2324 (O_2324,N_16392,N_18548);
nand UO_2325 (O_2325,N_18316,N_19308);
nor UO_2326 (O_2326,N_16118,N_16678);
and UO_2327 (O_2327,N_17699,N_16899);
and UO_2328 (O_2328,N_17124,N_16080);
nand UO_2329 (O_2329,N_18621,N_18252);
or UO_2330 (O_2330,N_15346,N_15909);
and UO_2331 (O_2331,N_19775,N_17633);
or UO_2332 (O_2332,N_16578,N_15987);
nand UO_2333 (O_2333,N_16258,N_18422);
and UO_2334 (O_2334,N_15671,N_18449);
nand UO_2335 (O_2335,N_19604,N_19712);
or UO_2336 (O_2336,N_18410,N_19527);
xnor UO_2337 (O_2337,N_15396,N_17957);
nor UO_2338 (O_2338,N_17366,N_15012);
and UO_2339 (O_2339,N_17447,N_16409);
nand UO_2340 (O_2340,N_15055,N_16450);
or UO_2341 (O_2341,N_18662,N_16256);
and UO_2342 (O_2342,N_19011,N_16527);
or UO_2343 (O_2343,N_15048,N_16543);
xnor UO_2344 (O_2344,N_15165,N_16714);
or UO_2345 (O_2345,N_15811,N_16203);
nor UO_2346 (O_2346,N_17214,N_15127);
and UO_2347 (O_2347,N_16553,N_18805);
nor UO_2348 (O_2348,N_17041,N_18803);
or UO_2349 (O_2349,N_19578,N_17462);
or UO_2350 (O_2350,N_16257,N_18109);
nand UO_2351 (O_2351,N_18028,N_16411);
nand UO_2352 (O_2352,N_17813,N_17438);
nor UO_2353 (O_2353,N_17155,N_17042);
nand UO_2354 (O_2354,N_17664,N_19476);
nor UO_2355 (O_2355,N_19383,N_15966);
nand UO_2356 (O_2356,N_15163,N_16512);
or UO_2357 (O_2357,N_18043,N_17960);
and UO_2358 (O_2358,N_18975,N_19392);
or UO_2359 (O_2359,N_19097,N_18588);
nand UO_2360 (O_2360,N_18504,N_17984);
nand UO_2361 (O_2361,N_17470,N_16292);
nor UO_2362 (O_2362,N_17893,N_19393);
xnor UO_2363 (O_2363,N_19924,N_15598);
and UO_2364 (O_2364,N_19899,N_16178);
nand UO_2365 (O_2365,N_18859,N_18207);
nand UO_2366 (O_2366,N_18953,N_16833);
and UO_2367 (O_2367,N_18949,N_17722);
nor UO_2368 (O_2368,N_18438,N_18222);
or UO_2369 (O_2369,N_18133,N_18725);
xor UO_2370 (O_2370,N_17172,N_15830);
nor UO_2371 (O_2371,N_16900,N_18506);
or UO_2372 (O_2372,N_18523,N_19664);
nor UO_2373 (O_2373,N_15593,N_18315);
nand UO_2374 (O_2374,N_18436,N_17668);
nand UO_2375 (O_2375,N_15406,N_16563);
nor UO_2376 (O_2376,N_16366,N_19558);
nand UO_2377 (O_2377,N_19040,N_18526);
nor UO_2378 (O_2378,N_15737,N_17213);
xnor UO_2379 (O_2379,N_15799,N_16022);
nor UO_2380 (O_2380,N_17492,N_17839);
nand UO_2381 (O_2381,N_19780,N_17360);
nand UO_2382 (O_2382,N_17806,N_19174);
nand UO_2383 (O_2383,N_18310,N_16803);
and UO_2384 (O_2384,N_18738,N_15815);
nand UO_2385 (O_2385,N_15196,N_19074);
nand UO_2386 (O_2386,N_18143,N_15803);
and UO_2387 (O_2387,N_19381,N_19080);
nand UO_2388 (O_2388,N_17050,N_16123);
or UO_2389 (O_2389,N_19085,N_18599);
or UO_2390 (O_2390,N_16879,N_18558);
nor UO_2391 (O_2391,N_19798,N_17744);
nand UO_2392 (O_2392,N_15394,N_15022);
xor UO_2393 (O_2393,N_17509,N_15652);
nand UO_2394 (O_2394,N_15040,N_17586);
nor UO_2395 (O_2395,N_19176,N_15565);
nor UO_2396 (O_2396,N_16003,N_18233);
nand UO_2397 (O_2397,N_16793,N_18180);
xor UO_2398 (O_2398,N_15133,N_19352);
nand UO_2399 (O_2399,N_17114,N_18401);
and UO_2400 (O_2400,N_17486,N_18556);
nor UO_2401 (O_2401,N_15507,N_15977);
nor UO_2402 (O_2402,N_17433,N_19514);
nor UO_2403 (O_2403,N_17294,N_17327);
and UO_2404 (O_2404,N_18494,N_19949);
or UO_2405 (O_2405,N_17117,N_19439);
nor UO_2406 (O_2406,N_17430,N_19197);
nor UO_2407 (O_2407,N_18031,N_19450);
or UO_2408 (O_2408,N_16850,N_18696);
nor UO_2409 (O_2409,N_17106,N_15687);
nand UO_2410 (O_2410,N_16344,N_17849);
nor UO_2411 (O_2411,N_17736,N_15474);
or UO_2412 (O_2412,N_17752,N_19847);
or UO_2413 (O_2413,N_16696,N_18488);
nand UO_2414 (O_2414,N_16219,N_18625);
nor UO_2415 (O_2415,N_15694,N_18225);
nand UO_2416 (O_2416,N_19729,N_17504);
nor UO_2417 (O_2417,N_17468,N_17548);
nand UO_2418 (O_2418,N_18069,N_16636);
or UO_2419 (O_2419,N_15027,N_19452);
or UO_2420 (O_2420,N_15501,N_18355);
and UO_2421 (O_2421,N_19812,N_16540);
nand UO_2422 (O_2422,N_17822,N_16891);
nand UO_2423 (O_2423,N_15850,N_15790);
nor UO_2424 (O_2424,N_16939,N_15205);
and UO_2425 (O_2425,N_18016,N_15801);
and UO_2426 (O_2426,N_19457,N_15008);
nor UO_2427 (O_2427,N_15608,N_18500);
or UO_2428 (O_2428,N_15019,N_17249);
nor UO_2429 (O_2429,N_18166,N_18347);
nor UO_2430 (O_2430,N_16847,N_17888);
and UO_2431 (O_2431,N_17033,N_15941);
or UO_2432 (O_2432,N_15487,N_18323);
nand UO_2433 (O_2433,N_15249,N_19435);
or UO_2434 (O_2434,N_18922,N_19652);
nor UO_2435 (O_2435,N_17573,N_16088);
nor UO_2436 (O_2436,N_17298,N_17998);
xnor UO_2437 (O_2437,N_19760,N_19021);
nor UO_2438 (O_2438,N_19150,N_19395);
nand UO_2439 (O_2439,N_18637,N_18961);
or UO_2440 (O_2440,N_19164,N_19112);
nand UO_2441 (O_2441,N_18221,N_15279);
xor UO_2442 (O_2442,N_15759,N_17921);
and UO_2443 (O_2443,N_16862,N_19102);
and UO_2444 (O_2444,N_18648,N_16101);
and UO_2445 (O_2445,N_18126,N_15034);
nor UO_2446 (O_2446,N_17949,N_16104);
xor UO_2447 (O_2447,N_16404,N_17378);
xor UO_2448 (O_2448,N_18099,N_17437);
or UO_2449 (O_2449,N_17766,N_17282);
and UO_2450 (O_2450,N_17830,N_15728);
nor UO_2451 (O_2451,N_16760,N_16892);
or UO_2452 (O_2452,N_16811,N_17868);
xor UO_2453 (O_2453,N_19186,N_18690);
nor UO_2454 (O_2454,N_18284,N_15151);
nor UO_2455 (O_2455,N_15642,N_18189);
nor UO_2456 (O_2456,N_19679,N_18563);
and UO_2457 (O_2457,N_19163,N_18951);
nor UO_2458 (O_2458,N_15733,N_17244);
or UO_2459 (O_2459,N_17529,N_17085);
or UO_2460 (O_2460,N_15822,N_15597);
nand UO_2461 (O_2461,N_18646,N_15310);
nand UO_2462 (O_2462,N_15517,N_18377);
nor UO_2463 (O_2463,N_18604,N_17173);
and UO_2464 (O_2464,N_18008,N_17655);
xor UO_2465 (O_2465,N_17644,N_19337);
and UO_2466 (O_2466,N_15072,N_17498);
nand UO_2467 (O_2467,N_16233,N_16281);
and UO_2468 (O_2468,N_19152,N_15169);
or UO_2469 (O_2469,N_18440,N_19689);
nor UO_2470 (O_2470,N_19982,N_19997);
xnor UO_2471 (O_2471,N_15399,N_16029);
or UO_2472 (O_2472,N_17451,N_16248);
or UO_2473 (O_2473,N_17180,N_17108);
xor UO_2474 (O_2474,N_17523,N_15097);
nor UO_2475 (O_2475,N_17818,N_17448);
and UO_2476 (O_2476,N_16657,N_19759);
and UO_2477 (O_2477,N_17182,N_19668);
nor UO_2478 (O_2478,N_17841,N_15415);
nor UO_2479 (O_2479,N_16349,N_18485);
nand UO_2480 (O_2480,N_16624,N_18294);
xnor UO_2481 (O_2481,N_17695,N_17728);
and UO_2482 (O_2482,N_18543,N_15183);
nor UO_2483 (O_2483,N_17933,N_16194);
nor UO_2484 (O_2484,N_18956,N_19287);
or UO_2485 (O_2485,N_16037,N_19386);
or UO_2486 (O_2486,N_16346,N_15066);
or UO_2487 (O_2487,N_18515,N_16848);
and UO_2488 (O_2488,N_16052,N_19801);
or UO_2489 (O_2489,N_16758,N_19960);
xnor UO_2490 (O_2490,N_15472,N_19634);
nor UO_2491 (O_2491,N_17962,N_16996);
and UO_2492 (O_2492,N_16116,N_16880);
nor UO_2493 (O_2493,N_16671,N_19784);
nor UO_2494 (O_2494,N_15821,N_19116);
or UO_2495 (O_2495,N_18349,N_19376);
and UO_2496 (O_2496,N_15437,N_19368);
nand UO_2497 (O_2497,N_18641,N_17317);
and UO_2498 (O_2498,N_17756,N_15547);
nor UO_2499 (O_2499,N_18639,N_15423);
endmodule