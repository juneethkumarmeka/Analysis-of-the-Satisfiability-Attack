module basic_1000_10000_1500_10_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
and U0 (N_0,In_195,In_490);
xor U1 (N_1,In_831,In_101);
nor U2 (N_2,In_224,In_638);
nor U3 (N_3,In_604,In_268);
nand U4 (N_4,In_353,In_299);
nor U5 (N_5,In_547,In_303);
nor U6 (N_6,In_730,In_568);
and U7 (N_7,In_612,In_354);
and U8 (N_8,In_566,In_881);
nand U9 (N_9,In_617,In_986);
xnor U10 (N_10,In_713,In_40);
nor U11 (N_11,In_912,In_697);
nor U12 (N_12,In_652,In_773);
and U13 (N_13,In_699,In_808);
or U14 (N_14,In_736,In_732);
xor U15 (N_15,In_508,In_650);
nand U16 (N_16,In_579,In_138);
or U17 (N_17,In_246,In_1);
and U18 (N_18,In_830,In_92);
nor U19 (N_19,In_464,In_918);
and U20 (N_20,In_476,In_387);
nand U21 (N_21,In_893,In_882);
and U22 (N_22,In_645,In_729);
nor U23 (N_23,In_160,In_189);
nand U24 (N_24,In_456,In_781);
nor U25 (N_25,In_647,In_156);
or U26 (N_26,In_479,In_174);
xor U27 (N_27,In_153,In_328);
xor U28 (N_28,In_110,In_149);
and U29 (N_29,In_178,In_368);
or U30 (N_30,In_176,In_289);
nand U31 (N_31,In_544,In_70);
or U32 (N_32,In_217,In_596);
or U33 (N_33,In_471,In_292);
or U34 (N_34,In_747,In_10);
and U35 (N_35,In_534,In_28);
nand U36 (N_36,In_784,In_513);
nand U37 (N_37,In_553,In_839);
xnor U38 (N_38,In_469,In_585);
nor U39 (N_39,In_897,In_120);
xor U40 (N_40,In_477,In_127);
nor U41 (N_41,In_648,In_284);
xor U42 (N_42,In_663,In_459);
or U43 (N_43,In_431,In_678);
or U44 (N_44,In_518,In_852);
and U45 (N_45,In_18,In_61);
xnor U46 (N_46,In_443,In_14);
nor U47 (N_47,In_792,In_54);
nand U48 (N_48,In_623,In_777);
and U49 (N_49,In_653,In_631);
nor U50 (N_50,In_819,In_436);
nand U51 (N_51,In_822,In_901);
and U52 (N_52,In_228,In_398);
nand U53 (N_53,In_415,In_25);
nand U54 (N_54,In_786,In_0);
nor U55 (N_55,In_975,In_362);
nor U56 (N_56,In_472,In_187);
and U57 (N_57,In_506,In_993);
or U58 (N_58,In_129,In_32);
or U59 (N_59,In_919,In_49);
and U60 (N_60,In_821,In_649);
nand U61 (N_61,In_332,In_619);
xor U62 (N_62,In_846,In_673);
nand U63 (N_63,In_595,In_221);
nand U64 (N_64,In_709,In_529);
or U65 (N_65,In_628,In_770);
xnor U66 (N_66,In_744,In_403);
xnor U67 (N_67,In_820,In_378);
xnor U68 (N_68,In_832,In_861);
or U69 (N_69,In_266,In_416);
and U70 (N_70,In_757,In_389);
or U71 (N_71,In_966,In_945);
and U72 (N_72,In_36,In_778);
xnor U73 (N_73,In_43,In_935);
xor U74 (N_74,In_760,In_150);
and U75 (N_75,In_449,In_375);
or U76 (N_76,In_31,In_970);
or U77 (N_77,In_504,In_636);
xor U78 (N_78,In_72,In_698);
nand U79 (N_79,In_510,In_4);
nand U80 (N_80,In_835,In_34);
nand U81 (N_81,In_583,In_637);
or U82 (N_82,In_580,In_38);
xnor U83 (N_83,In_458,In_564);
and U84 (N_84,In_420,In_626);
nand U85 (N_85,In_344,In_202);
xnor U86 (N_86,In_588,In_322);
and U87 (N_87,In_664,In_498);
or U88 (N_88,In_275,In_853);
or U89 (N_89,In_6,In_294);
nor U90 (N_90,In_184,In_512);
xor U91 (N_91,In_335,In_85);
nand U92 (N_92,In_842,In_738);
nand U93 (N_93,In_116,In_291);
nor U94 (N_94,In_843,In_687);
nor U95 (N_95,In_179,In_593);
and U96 (N_96,In_305,In_561);
nor U97 (N_97,In_502,In_983);
nand U98 (N_98,In_88,In_761);
or U99 (N_99,In_943,In_39);
nor U100 (N_100,In_177,In_310);
or U101 (N_101,In_142,In_696);
xnor U102 (N_102,In_348,In_962);
nand U103 (N_103,In_355,In_263);
or U104 (N_104,In_418,In_557);
nand U105 (N_105,In_2,In_98);
nand U106 (N_106,In_454,In_349);
or U107 (N_107,In_183,In_740);
and U108 (N_108,In_260,In_682);
nand U109 (N_109,In_857,In_237);
nor U110 (N_110,In_47,In_190);
nor U111 (N_111,In_324,In_312);
nor U112 (N_112,In_735,In_837);
or U113 (N_113,In_694,In_392);
xor U114 (N_114,In_944,In_51);
nor U115 (N_115,In_692,In_317);
and U116 (N_116,In_685,In_491);
or U117 (N_117,In_269,In_277);
nand U118 (N_118,In_474,In_231);
and U119 (N_119,In_505,In_841);
and U120 (N_120,In_932,In_122);
nand U121 (N_121,In_995,In_118);
nand U122 (N_122,In_394,In_964);
or U123 (N_123,In_62,In_391);
nor U124 (N_124,In_703,In_300);
nor U125 (N_125,In_91,In_106);
nor U126 (N_126,In_531,In_571);
nand U127 (N_127,In_429,In_136);
or U128 (N_128,In_79,In_655);
xor U129 (N_129,In_186,In_802);
and U130 (N_130,In_771,In_968);
and U131 (N_131,In_370,In_511);
xnor U132 (N_132,In_680,In_222);
or U133 (N_133,In_996,In_427);
nand U134 (N_134,In_325,In_811);
nand U135 (N_135,In_577,In_295);
or U136 (N_136,In_223,In_849);
nand U137 (N_137,In_515,In_794);
or U138 (N_138,In_871,In_807);
or U139 (N_139,In_360,In_621);
nor U140 (N_140,In_446,In_766);
and U141 (N_141,In_691,In_939);
nand U142 (N_142,In_969,In_565);
nand U143 (N_143,In_288,In_878);
or U144 (N_144,In_957,In_574);
or U145 (N_145,In_308,In_599);
nor U146 (N_146,In_862,In_319);
and U147 (N_147,In_985,In_722);
xor U148 (N_148,In_542,In_94);
nand U149 (N_149,In_592,In_608);
nor U150 (N_150,In_941,In_590);
or U151 (N_151,In_175,In_734);
nand U152 (N_152,In_441,In_748);
nand U153 (N_153,In_311,In_892);
nand U154 (N_154,In_530,In_203);
and U155 (N_155,In_690,In_789);
xnor U156 (N_156,In_782,In_232);
or U157 (N_157,In_211,In_358);
xor U158 (N_158,In_89,In_976);
nand U159 (N_159,In_992,In_793);
nor U160 (N_160,In_80,In_439);
nor U161 (N_161,In_972,In_618);
xor U162 (N_162,In_874,In_890);
and U163 (N_163,In_676,In_147);
xnor U164 (N_164,In_487,In_933);
nor U165 (N_165,In_280,In_208);
or U166 (N_166,In_250,In_629);
or U167 (N_167,In_408,In_213);
or U168 (N_168,In_661,In_902);
or U169 (N_169,In_154,In_644);
or U170 (N_170,In_710,In_484);
nor U171 (N_171,In_405,In_594);
and U172 (N_172,In_109,In_172);
or U173 (N_173,In_538,In_486);
or U174 (N_174,In_905,In_753);
or U175 (N_175,In_244,In_768);
and U176 (N_176,In_410,In_111);
and U177 (N_177,In_15,In_666);
nand U178 (N_178,In_705,In_642);
xor U179 (N_179,In_276,In_380);
and U180 (N_180,In_982,In_974);
and U181 (N_181,In_501,In_146);
nand U182 (N_182,In_739,In_795);
and U183 (N_183,In_297,In_78);
or U184 (N_184,In_827,In_435);
or U185 (N_185,In_906,In_242);
nand U186 (N_186,In_990,In_714);
or U187 (N_187,In_550,In_340);
nand U188 (N_188,In_475,In_314);
or U189 (N_189,In_913,In_724);
xnor U190 (N_190,In_489,In_667);
nor U191 (N_191,In_763,In_342);
nor U192 (N_192,In_745,In_401);
nor U193 (N_193,In_455,In_81);
and U194 (N_194,In_826,In_979);
nor U195 (N_195,In_818,In_41);
and U196 (N_196,In_910,In_977);
and U197 (N_197,In_96,In_824);
nor U198 (N_198,In_468,In_866);
nand U199 (N_199,In_876,In_921);
and U200 (N_200,In_614,In_914);
nand U201 (N_201,In_315,In_980);
or U202 (N_202,In_677,In_602);
nor U203 (N_203,In_872,In_115);
or U204 (N_204,In_404,In_955);
nor U205 (N_205,In_74,In_445);
nor U206 (N_206,In_265,In_702);
and U207 (N_207,In_665,In_848);
xor U208 (N_208,In_407,In_584);
nor U209 (N_209,In_790,In_293);
xnor U210 (N_210,In_836,In_157);
and U211 (N_211,In_825,In_365);
nand U212 (N_212,In_956,In_591);
or U213 (N_213,In_53,In_400);
nand U214 (N_214,In_382,In_50);
nor U215 (N_215,In_715,In_77);
and U216 (N_216,In_999,In_625);
nand U217 (N_217,In_69,In_113);
nand U218 (N_218,In_520,In_723);
nor U219 (N_219,In_804,In_488);
and U220 (N_220,In_681,In_218);
xor U221 (N_221,In_797,In_788);
xor U222 (N_222,In_803,In_357);
xnor U223 (N_223,In_562,In_60);
xor U224 (N_224,In_143,In_546);
and U225 (N_225,In_952,In_169);
xnor U226 (N_226,In_963,In_75);
or U227 (N_227,In_199,In_316);
and U228 (N_228,In_726,In_423);
and U229 (N_229,In_984,In_904);
nor U230 (N_230,In_785,In_167);
nor U231 (N_231,In_27,In_519);
or U232 (N_232,In_121,In_103);
and U233 (N_233,In_670,In_227);
and U234 (N_234,In_573,In_385);
and U235 (N_235,In_13,In_847);
and U236 (N_236,In_216,In_76);
xor U237 (N_237,In_219,In_397);
xor U238 (N_238,In_194,In_895);
nor U239 (N_239,In_799,In_589);
nand U240 (N_240,In_522,In_298);
nand U241 (N_241,In_376,In_381);
and U242 (N_242,In_615,In_9);
and U243 (N_243,In_279,In_609);
nor U244 (N_244,In_998,In_256);
or U245 (N_245,In_662,In_442);
nand U246 (N_246,In_386,In_128);
or U247 (N_247,In_537,In_500);
and U248 (N_248,In_457,In_988);
or U249 (N_249,In_450,In_336);
or U250 (N_250,In_16,In_758);
xnor U251 (N_251,In_497,In_273);
xnor U252 (N_252,In_624,In_880);
or U253 (N_253,In_11,In_411);
or U254 (N_254,In_885,In_728);
xor U255 (N_255,In_52,In_927);
and U256 (N_256,In_815,In_460);
nor U257 (N_257,In_750,In_278);
or U258 (N_258,In_865,In_930);
xor U259 (N_259,In_946,In_509);
and U260 (N_260,In_163,In_331);
and U261 (N_261,In_801,In_413);
xnor U262 (N_262,In_12,In_967);
or U263 (N_263,In_139,In_341);
or U264 (N_264,In_249,In_828);
nor U265 (N_265,In_214,In_225);
xor U266 (N_266,In_524,In_124);
nor U267 (N_267,In_971,In_669);
nor U268 (N_268,In_923,In_719);
xor U269 (N_269,In_347,In_704);
and U270 (N_270,In_675,In_434);
and U271 (N_271,In_108,In_137);
xor U272 (N_272,In_168,In_869);
nand U273 (N_273,In_119,In_236);
or U274 (N_274,In_55,In_285);
nor U275 (N_275,In_605,In_64);
nor U276 (N_276,In_388,In_164);
nand U277 (N_277,In_99,In_720);
nand U278 (N_278,In_422,In_873);
and U279 (N_279,In_751,In_492);
or U280 (N_280,In_377,In_356);
xor U281 (N_281,In_533,In_679);
nand U282 (N_282,In_166,In_688);
or U283 (N_283,In_953,In_598);
nor U284 (N_284,In_516,In_258);
and U285 (N_285,In_706,In_390);
nor U286 (N_286,In_743,In_911);
and U287 (N_287,In_616,In_654);
or U288 (N_288,In_527,In_428);
or U289 (N_289,In_960,In_765);
nor U290 (N_290,In_112,In_65);
nor U291 (N_291,In_507,In_417);
nor U292 (N_292,In_68,In_659);
xnor U293 (N_293,In_406,In_627);
nand U294 (N_294,In_950,In_686);
nand U295 (N_295,In_635,In_367);
nor U296 (N_296,In_205,In_29);
nand U297 (N_297,In_270,In_586);
or U298 (N_298,In_948,In_241);
and U299 (N_299,In_155,In_525);
or U300 (N_300,In_57,In_97);
nand U301 (N_301,In_20,In_233);
nand U302 (N_302,In_742,In_235);
and U303 (N_303,In_909,In_264);
or U304 (N_304,In_622,In_535);
or U305 (N_305,In_132,In_338);
nand U306 (N_306,In_282,In_483);
xor U307 (N_307,In_95,In_152);
nor U308 (N_308,In_526,In_783);
nand U309 (N_309,In_672,In_741);
xor U310 (N_310,In_949,In_46);
and U311 (N_311,In_306,In_674);
nand U312 (N_312,In_894,In_452);
and U313 (N_313,In_366,In_554);
and U314 (N_314,In_318,In_274);
and U315 (N_315,In_363,In_188);
nor U316 (N_316,In_937,In_93);
nand U317 (N_317,In_643,In_145);
and U318 (N_318,In_117,In_220);
xor U319 (N_319,In_125,In_234);
nor U320 (N_320,In_259,In_240);
and U321 (N_321,In_467,In_560);
xnor U322 (N_322,In_343,In_817);
nand U323 (N_323,In_684,In_806);
or U324 (N_324,In_576,In_131);
and U325 (N_325,In_453,In_767);
or U326 (N_326,In_620,In_425);
and U327 (N_327,In_100,In_958);
and U328 (N_328,In_915,In_182);
xor U329 (N_329,In_339,In_517);
nor U330 (N_330,In_201,In_931);
nand U331 (N_331,In_942,In_495);
nand U332 (N_332,In_731,In_272);
nor U333 (N_333,In_359,In_695);
or U334 (N_334,In_920,In_973);
nor U335 (N_335,In_860,In_287);
nand U336 (N_336,In_180,In_606);
xor U337 (N_337,In_481,In_896);
xor U338 (N_338,In_572,In_746);
xnor U339 (N_339,In_267,In_255);
nor U340 (N_340,In_463,In_45);
or U341 (N_341,In_523,In_198);
or U342 (N_342,In_430,In_286);
nor U343 (N_343,In_104,In_708);
nand U344 (N_344,In_290,In_42);
nand U345 (N_345,In_374,In_987);
and U346 (N_346,In_929,In_823);
and U347 (N_347,In_426,In_321);
xnor U348 (N_348,In_536,In_140);
xnor U349 (N_349,In_875,In_462);
and U350 (N_350,In_334,In_800);
or U351 (N_351,In_361,In_409);
and U352 (N_352,In_337,In_610);
or U353 (N_353,In_780,In_485);
nand U354 (N_354,In_204,In_888);
xor U355 (N_355,In_759,In_668);
xnor U356 (N_356,In_296,In_600);
or U357 (N_357,In_587,In_257);
nand U358 (N_358,In_283,In_539);
and U359 (N_359,In_226,In_133);
nor U360 (N_360,In_123,In_575);
and U361 (N_361,In_925,In_165);
or U362 (N_362,In_922,In_215);
nor U363 (N_363,In_916,In_991);
or U364 (N_364,In_640,In_549);
and U365 (N_365,In_989,In_981);
xor U366 (N_366,In_601,In_805);
or U367 (N_367,In_86,In_717);
xnor U368 (N_368,In_58,In_954);
nor U369 (N_369,In_711,In_83);
and U370 (N_370,In_752,In_755);
and U371 (N_371,In_301,In_603);
xnor U372 (N_372,In_421,In_859);
and U373 (N_373,In_33,In_552);
nand U374 (N_374,In_364,In_87);
and U375 (N_375,In_521,In_440);
xnor U376 (N_376,In_170,In_307);
nor U377 (N_377,In_309,In_940);
nor U378 (N_378,In_934,In_7);
nor U379 (N_379,In_480,In_633);
nand U380 (N_380,In_660,In_281);
xnor U381 (N_381,In_372,In_8);
nor U382 (N_382,In_809,In_883);
nor U383 (N_383,In_854,In_891);
or U384 (N_384,In_864,In_813);
nand U385 (N_385,In_56,In_230);
nand U386 (N_386,In_938,In_856);
nor U387 (N_387,In_448,In_229);
or U388 (N_388,In_302,In_494);
and U389 (N_389,In_994,In_84);
or U390 (N_390,In_251,In_917);
xnor U391 (N_391,In_151,In_689);
and U392 (N_392,In_559,In_238);
xor U393 (N_393,In_383,In_438);
and U394 (N_394,In_181,In_67);
or U395 (N_395,In_30,In_838);
nand U396 (N_396,In_262,In_725);
xor U397 (N_397,In_886,In_162);
or U398 (N_398,In_173,In_158);
and U399 (N_399,In_191,In_114);
nand U400 (N_400,In_210,In_769);
nor U401 (N_401,In_197,In_141);
and U402 (N_402,In_570,In_253);
nor U403 (N_403,In_727,In_721);
or U404 (N_404,In_997,In_834);
xnor U405 (N_405,In_558,In_639);
and U406 (N_406,In_582,In_693);
or U407 (N_407,In_884,In_936);
xnor U408 (N_408,In_323,In_701);
and U409 (N_409,In_379,In_393);
nor U410 (N_410,In_466,In_924);
xor U411 (N_411,In_541,In_22);
nand U412 (N_412,In_499,In_764);
nand U413 (N_413,In_271,In_247);
or U414 (N_414,In_3,In_17);
or U415 (N_415,In_716,In_451);
xor U416 (N_416,In_185,In_59);
nor U417 (N_417,In_641,In_19);
nand U418 (N_418,In_514,In_461);
xnor U419 (N_419,In_396,In_73);
nand U420 (N_420,In_556,In_209);
and U421 (N_421,In_63,In_329);
or U422 (N_422,In_754,In_850);
nand U423 (N_423,In_555,In_35);
and U424 (N_424,In_24,In_212);
nand U425 (N_425,In_718,In_243);
and U426 (N_426,In_569,In_908);
nor U427 (N_427,In_898,In_196);
xnor U428 (N_428,In_630,In_252);
nor U429 (N_429,In_432,In_102);
and U430 (N_430,In_611,In_814);
and U431 (N_431,In_798,In_134);
nor U432 (N_432,In_352,In_207);
or U433 (N_433,In_350,In_161);
nand U434 (N_434,In_887,In_193);
or U435 (N_435,In_829,In_419);
xnor U436 (N_436,In_23,In_656);
xor U437 (N_437,In_470,In_5);
xnor U438 (N_438,In_737,In_482);
nor U439 (N_439,In_791,In_749);
or U440 (N_440,In_840,In_369);
nor U441 (N_441,In_532,In_496);
xnor U442 (N_442,In_683,In_581);
nand U443 (N_443,In_774,In_159);
xnor U444 (N_444,In_206,In_130);
xnor U445 (N_445,In_528,In_414);
or U446 (N_446,In_907,In_26);
and U447 (N_447,In_346,In_444);
or U448 (N_448,In_543,In_597);
nand U449 (N_449,In_607,In_578);
nor U450 (N_450,In_867,In_44);
or U451 (N_451,In_700,In_926);
nand U452 (N_452,In_961,In_254);
nand U453 (N_453,In_870,In_493);
or U454 (N_454,In_816,In_632);
and U455 (N_455,In_473,In_812);
nor U456 (N_456,In_567,In_775);
xnor U457 (N_457,In_978,In_135);
and U458 (N_458,In_21,In_399);
and U459 (N_459,In_779,In_37);
and U460 (N_460,In_563,In_863);
and U461 (N_461,In_503,In_877);
and U462 (N_462,In_796,In_551);
nand U463 (N_463,In_657,In_373);
nor U464 (N_464,In_424,In_144);
and U465 (N_465,In_326,In_402);
or U466 (N_466,In_879,In_951);
nand U467 (N_467,In_192,In_646);
and U468 (N_468,In_707,In_671);
or U469 (N_469,In_903,In_787);
xor U470 (N_470,In_959,In_756);
nand U471 (N_471,In_900,In_545);
nand U472 (N_472,In_107,In_855);
or U473 (N_473,In_658,In_651);
nor U474 (N_474,In_947,In_447);
nand U475 (N_475,In_437,In_851);
xnor U476 (N_476,In_548,In_845);
xor U477 (N_477,In_148,In_540);
xnor U478 (N_478,In_858,In_762);
nand U479 (N_479,In_327,In_333);
and U480 (N_480,In_261,In_90);
and U481 (N_481,In_200,In_899);
nand U482 (N_482,In_810,In_345);
or U483 (N_483,In_48,In_965);
nor U484 (N_484,In_772,In_330);
nor U485 (N_485,In_126,In_239);
nand U486 (N_486,In_351,In_248);
and U487 (N_487,In_868,In_712);
nor U488 (N_488,In_833,In_478);
or U489 (N_489,In_82,In_844);
and U490 (N_490,In_384,In_245);
xnor U491 (N_491,In_733,In_171);
xnor U492 (N_492,In_776,In_412);
nand U493 (N_493,In_465,In_395);
xor U494 (N_494,In_433,In_613);
xor U495 (N_495,In_371,In_320);
nor U496 (N_496,In_928,In_313);
and U497 (N_497,In_66,In_304);
or U498 (N_498,In_105,In_889);
and U499 (N_499,In_71,In_634);
and U500 (N_500,In_775,In_168);
or U501 (N_501,In_135,In_891);
or U502 (N_502,In_691,In_147);
and U503 (N_503,In_267,In_290);
nor U504 (N_504,In_353,In_467);
and U505 (N_505,In_123,In_139);
and U506 (N_506,In_97,In_112);
or U507 (N_507,In_518,In_67);
or U508 (N_508,In_899,In_357);
nand U509 (N_509,In_210,In_509);
and U510 (N_510,In_903,In_95);
and U511 (N_511,In_866,In_108);
or U512 (N_512,In_868,In_296);
or U513 (N_513,In_19,In_501);
nor U514 (N_514,In_21,In_898);
and U515 (N_515,In_159,In_592);
xnor U516 (N_516,In_75,In_45);
xor U517 (N_517,In_7,In_48);
or U518 (N_518,In_481,In_381);
nor U519 (N_519,In_159,In_289);
nand U520 (N_520,In_322,In_865);
or U521 (N_521,In_380,In_864);
xor U522 (N_522,In_531,In_871);
nand U523 (N_523,In_342,In_348);
xnor U524 (N_524,In_404,In_54);
or U525 (N_525,In_226,In_807);
and U526 (N_526,In_361,In_108);
xor U527 (N_527,In_975,In_677);
nor U528 (N_528,In_961,In_319);
and U529 (N_529,In_766,In_132);
or U530 (N_530,In_695,In_105);
and U531 (N_531,In_285,In_780);
and U532 (N_532,In_686,In_847);
xnor U533 (N_533,In_703,In_316);
nor U534 (N_534,In_720,In_518);
or U535 (N_535,In_371,In_526);
or U536 (N_536,In_170,In_89);
xnor U537 (N_537,In_696,In_222);
nor U538 (N_538,In_964,In_19);
nor U539 (N_539,In_967,In_283);
nand U540 (N_540,In_308,In_675);
xor U541 (N_541,In_533,In_23);
nor U542 (N_542,In_928,In_282);
nand U543 (N_543,In_375,In_464);
nand U544 (N_544,In_859,In_141);
xor U545 (N_545,In_591,In_580);
nor U546 (N_546,In_485,In_644);
or U547 (N_547,In_153,In_545);
xnor U548 (N_548,In_362,In_373);
or U549 (N_549,In_349,In_657);
or U550 (N_550,In_765,In_102);
xor U551 (N_551,In_891,In_675);
nand U552 (N_552,In_98,In_414);
xnor U553 (N_553,In_527,In_544);
and U554 (N_554,In_586,In_494);
nand U555 (N_555,In_743,In_438);
and U556 (N_556,In_433,In_120);
nand U557 (N_557,In_714,In_424);
xor U558 (N_558,In_582,In_90);
nor U559 (N_559,In_207,In_42);
nand U560 (N_560,In_240,In_292);
and U561 (N_561,In_406,In_871);
or U562 (N_562,In_425,In_649);
nor U563 (N_563,In_43,In_3);
nand U564 (N_564,In_616,In_278);
xnor U565 (N_565,In_495,In_910);
and U566 (N_566,In_717,In_685);
and U567 (N_567,In_61,In_441);
and U568 (N_568,In_840,In_577);
nand U569 (N_569,In_507,In_171);
nor U570 (N_570,In_797,In_852);
nand U571 (N_571,In_917,In_397);
nor U572 (N_572,In_486,In_303);
or U573 (N_573,In_463,In_974);
nor U574 (N_574,In_202,In_980);
nor U575 (N_575,In_465,In_241);
xnor U576 (N_576,In_899,In_300);
nor U577 (N_577,In_911,In_217);
nor U578 (N_578,In_17,In_854);
nand U579 (N_579,In_339,In_252);
xnor U580 (N_580,In_464,In_270);
or U581 (N_581,In_537,In_3);
and U582 (N_582,In_254,In_521);
nand U583 (N_583,In_26,In_541);
xnor U584 (N_584,In_541,In_409);
nand U585 (N_585,In_815,In_161);
or U586 (N_586,In_584,In_314);
nor U587 (N_587,In_991,In_580);
nor U588 (N_588,In_612,In_109);
or U589 (N_589,In_627,In_879);
and U590 (N_590,In_530,In_233);
nor U591 (N_591,In_623,In_402);
nor U592 (N_592,In_884,In_859);
nor U593 (N_593,In_175,In_631);
nor U594 (N_594,In_222,In_985);
xnor U595 (N_595,In_581,In_134);
nand U596 (N_596,In_737,In_513);
xor U597 (N_597,In_598,In_440);
nand U598 (N_598,In_444,In_540);
and U599 (N_599,In_875,In_749);
nor U600 (N_600,In_214,In_245);
xor U601 (N_601,In_182,In_686);
or U602 (N_602,In_536,In_27);
or U603 (N_603,In_97,In_82);
nor U604 (N_604,In_265,In_856);
xor U605 (N_605,In_750,In_221);
and U606 (N_606,In_644,In_144);
nor U607 (N_607,In_525,In_724);
nor U608 (N_608,In_132,In_744);
nand U609 (N_609,In_300,In_473);
xnor U610 (N_610,In_113,In_730);
or U611 (N_611,In_190,In_448);
or U612 (N_612,In_767,In_488);
nor U613 (N_613,In_778,In_412);
nor U614 (N_614,In_360,In_619);
and U615 (N_615,In_140,In_211);
nor U616 (N_616,In_330,In_847);
xor U617 (N_617,In_355,In_815);
xor U618 (N_618,In_893,In_703);
or U619 (N_619,In_578,In_312);
and U620 (N_620,In_934,In_39);
or U621 (N_621,In_810,In_309);
nand U622 (N_622,In_454,In_399);
nand U623 (N_623,In_63,In_668);
and U624 (N_624,In_441,In_407);
xnor U625 (N_625,In_566,In_382);
xor U626 (N_626,In_166,In_900);
nand U627 (N_627,In_828,In_81);
nor U628 (N_628,In_895,In_119);
or U629 (N_629,In_555,In_321);
nor U630 (N_630,In_82,In_214);
xnor U631 (N_631,In_594,In_662);
nand U632 (N_632,In_49,In_217);
or U633 (N_633,In_146,In_773);
or U634 (N_634,In_80,In_120);
nand U635 (N_635,In_377,In_3);
nor U636 (N_636,In_481,In_78);
xnor U637 (N_637,In_678,In_425);
xor U638 (N_638,In_390,In_931);
and U639 (N_639,In_636,In_241);
nor U640 (N_640,In_789,In_398);
and U641 (N_641,In_44,In_940);
nor U642 (N_642,In_454,In_987);
nand U643 (N_643,In_779,In_277);
or U644 (N_644,In_102,In_762);
nor U645 (N_645,In_251,In_102);
nand U646 (N_646,In_937,In_135);
nand U647 (N_647,In_156,In_637);
and U648 (N_648,In_410,In_739);
nor U649 (N_649,In_250,In_298);
or U650 (N_650,In_992,In_738);
and U651 (N_651,In_621,In_928);
and U652 (N_652,In_579,In_824);
and U653 (N_653,In_402,In_152);
xnor U654 (N_654,In_142,In_748);
and U655 (N_655,In_349,In_754);
xnor U656 (N_656,In_918,In_236);
nand U657 (N_657,In_397,In_517);
or U658 (N_658,In_955,In_496);
nor U659 (N_659,In_587,In_197);
or U660 (N_660,In_878,In_101);
nor U661 (N_661,In_895,In_361);
nor U662 (N_662,In_233,In_337);
nor U663 (N_663,In_923,In_836);
xor U664 (N_664,In_147,In_960);
xnor U665 (N_665,In_367,In_362);
nand U666 (N_666,In_128,In_282);
xnor U667 (N_667,In_146,In_509);
or U668 (N_668,In_783,In_875);
and U669 (N_669,In_71,In_606);
nor U670 (N_670,In_93,In_62);
xor U671 (N_671,In_886,In_800);
nand U672 (N_672,In_204,In_746);
nor U673 (N_673,In_921,In_160);
xnor U674 (N_674,In_309,In_589);
and U675 (N_675,In_24,In_325);
and U676 (N_676,In_457,In_864);
nand U677 (N_677,In_982,In_262);
and U678 (N_678,In_782,In_825);
nor U679 (N_679,In_313,In_63);
xnor U680 (N_680,In_910,In_473);
nor U681 (N_681,In_910,In_591);
nor U682 (N_682,In_65,In_102);
or U683 (N_683,In_404,In_628);
nor U684 (N_684,In_970,In_408);
and U685 (N_685,In_734,In_22);
nand U686 (N_686,In_107,In_348);
nor U687 (N_687,In_312,In_978);
or U688 (N_688,In_31,In_704);
nand U689 (N_689,In_971,In_779);
and U690 (N_690,In_250,In_609);
nor U691 (N_691,In_75,In_819);
nor U692 (N_692,In_450,In_967);
nor U693 (N_693,In_525,In_888);
nand U694 (N_694,In_977,In_165);
and U695 (N_695,In_377,In_733);
or U696 (N_696,In_723,In_978);
xnor U697 (N_697,In_983,In_722);
nand U698 (N_698,In_111,In_705);
xor U699 (N_699,In_629,In_519);
or U700 (N_700,In_852,In_127);
nand U701 (N_701,In_661,In_557);
nand U702 (N_702,In_854,In_615);
nand U703 (N_703,In_399,In_361);
and U704 (N_704,In_207,In_322);
xor U705 (N_705,In_411,In_602);
nor U706 (N_706,In_938,In_436);
nand U707 (N_707,In_450,In_836);
xor U708 (N_708,In_921,In_308);
xor U709 (N_709,In_1,In_410);
or U710 (N_710,In_524,In_23);
nor U711 (N_711,In_630,In_951);
xor U712 (N_712,In_73,In_86);
nor U713 (N_713,In_333,In_660);
or U714 (N_714,In_373,In_491);
or U715 (N_715,In_926,In_833);
or U716 (N_716,In_582,In_32);
or U717 (N_717,In_472,In_387);
nor U718 (N_718,In_994,In_969);
nor U719 (N_719,In_503,In_631);
or U720 (N_720,In_371,In_348);
or U721 (N_721,In_785,In_573);
nand U722 (N_722,In_394,In_348);
xor U723 (N_723,In_736,In_989);
or U724 (N_724,In_263,In_831);
xnor U725 (N_725,In_763,In_360);
or U726 (N_726,In_349,In_453);
or U727 (N_727,In_248,In_299);
and U728 (N_728,In_84,In_488);
xor U729 (N_729,In_687,In_143);
xor U730 (N_730,In_17,In_847);
nor U731 (N_731,In_364,In_685);
nor U732 (N_732,In_900,In_751);
and U733 (N_733,In_740,In_509);
or U734 (N_734,In_41,In_501);
nand U735 (N_735,In_628,In_435);
and U736 (N_736,In_6,In_857);
xnor U737 (N_737,In_199,In_775);
and U738 (N_738,In_40,In_615);
nor U739 (N_739,In_750,In_797);
and U740 (N_740,In_60,In_778);
or U741 (N_741,In_161,In_649);
and U742 (N_742,In_359,In_384);
nor U743 (N_743,In_946,In_165);
and U744 (N_744,In_373,In_134);
or U745 (N_745,In_673,In_753);
xor U746 (N_746,In_16,In_45);
nand U747 (N_747,In_952,In_561);
nor U748 (N_748,In_714,In_360);
xor U749 (N_749,In_721,In_797);
nand U750 (N_750,In_79,In_633);
and U751 (N_751,In_781,In_138);
nor U752 (N_752,In_783,In_151);
xnor U753 (N_753,In_842,In_766);
and U754 (N_754,In_889,In_820);
xnor U755 (N_755,In_160,In_844);
xnor U756 (N_756,In_849,In_329);
or U757 (N_757,In_166,In_490);
xnor U758 (N_758,In_716,In_45);
nor U759 (N_759,In_20,In_199);
nand U760 (N_760,In_792,In_603);
nor U761 (N_761,In_292,In_823);
nand U762 (N_762,In_418,In_467);
or U763 (N_763,In_133,In_996);
or U764 (N_764,In_58,In_635);
nor U765 (N_765,In_0,In_932);
nor U766 (N_766,In_298,In_740);
or U767 (N_767,In_648,In_507);
nor U768 (N_768,In_39,In_154);
and U769 (N_769,In_793,In_92);
and U770 (N_770,In_732,In_415);
and U771 (N_771,In_337,In_102);
nand U772 (N_772,In_362,In_407);
nor U773 (N_773,In_664,In_366);
or U774 (N_774,In_79,In_402);
nand U775 (N_775,In_302,In_449);
or U776 (N_776,In_312,In_251);
xnor U777 (N_777,In_800,In_119);
nor U778 (N_778,In_35,In_848);
nor U779 (N_779,In_672,In_884);
or U780 (N_780,In_267,In_402);
nor U781 (N_781,In_668,In_552);
nand U782 (N_782,In_565,In_96);
nor U783 (N_783,In_147,In_192);
and U784 (N_784,In_169,In_839);
or U785 (N_785,In_995,In_489);
and U786 (N_786,In_158,In_705);
nand U787 (N_787,In_203,In_822);
nor U788 (N_788,In_108,In_402);
or U789 (N_789,In_948,In_364);
or U790 (N_790,In_781,In_660);
nand U791 (N_791,In_139,In_728);
or U792 (N_792,In_470,In_71);
xor U793 (N_793,In_185,In_141);
nand U794 (N_794,In_759,In_333);
nand U795 (N_795,In_118,In_78);
nand U796 (N_796,In_399,In_321);
or U797 (N_797,In_688,In_859);
nor U798 (N_798,In_622,In_904);
nor U799 (N_799,In_516,In_46);
or U800 (N_800,In_552,In_772);
xnor U801 (N_801,In_319,In_731);
and U802 (N_802,In_582,In_465);
or U803 (N_803,In_166,In_764);
xnor U804 (N_804,In_651,In_763);
and U805 (N_805,In_372,In_285);
nor U806 (N_806,In_815,In_664);
nand U807 (N_807,In_995,In_864);
nand U808 (N_808,In_233,In_288);
nand U809 (N_809,In_969,In_996);
and U810 (N_810,In_751,In_190);
nor U811 (N_811,In_720,In_750);
nor U812 (N_812,In_684,In_604);
and U813 (N_813,In_180,In_843);
nand U814 (N_814,In_534,In_749);
and U815 (N_815,In_812,In_639);
and U816 (N_816,In_333,In_814);
and U817 (N_817,In_280,In_8);
nor U818 (N_818,In_516,In_162);
or U819 (N_819,In_742,In_99);
xnor U820 (N_820,In_205,In_869);
or U821 (N_821,In_9,In_236);
nand U822 (N_822,In_262,In_891);
nor U823 (N_823,In_321,In_933);
and U824 (N_824,In_938,In_388);
nand U825 (N_825,In_873,In_759);
nor U826 (N_826,In_833,In_325);
xnor U827 (N_827,In_143,In_879);
xnor U828 (N_828,In_860,In_567);
or U829 (N_829,In_166,In_651);
and U830 (N_830,In_695,In_183);
xor U831 (N_831,In_726,In_634);
or U832 (N_832,In_337,In_780);
and U833 (N_833,In_148,In_669);
xor U834 (N_834,In_830,In_366);
xnor U835 (N_835,In_983,In_39);
and U836 (N_836,In_266,In_450);
xor U837 (N_837,In_444,In_796);
nand U838 (N_838,In_113,In_205);
or U839 (N_839,In_311,In_375);
xnor U840 (N_840,In_271,In_380);
nand U841 (N_841,In_216,In_283);
and U842 (N_842,In_402,In_154);
and U843 (N_843,In_246,In_486);
xnor U844 (N_844,In_523,In_357);
xor U845 (N_845,In_233,In_697);
nor U846 (N_846,In_327,In_989);
nor U847 (N_847,In_432,In_475);
and U848 (N_848,In_231,In_316);
nor U849 (N_849,In_729,In_777);
and U850 (N_850,In_878,In_638);
nor U851 (N_851,In_683,In_42);
nand U852 (N_852,In_605,In_299);
nor U853 (N_853,In_279,In_25);
or U854 (N_854,In_263,In_576);
nand U855 (N_855,In_836,In_582);
and U856 (N_856,In_594,In_623);
and U857 (N_857,In_636,In_677);
or U858 (N_858,In_589,In_350);
xnor U859 (N_859,In_954,In_521);
nand U860 (N_860,In_122,In_676);
or U861 (N_861,In_686,In_536);
nand U862 (N_862,In_645,In_464);
nand U863 (N_863,In_683,In_644);
or U864 (N_864,In_834,In_465);
and U865 (N_865,In_413,In_24);
nor U866 (N_866,In_332,In_715);
nor U867 (N_867,In_567,In_48);
and U868 (N_868,In_570,In_284);
nor U869 (N_869,In_926,In_475);
nand U870 (N_870,In_767,In_875);
and U871 (N_871,In_660,In_124);
and U872 (N_872,In_192,In_69);
xnor U873 (N_873,In_17,In_134);
or U874 (N_874,In_422,In_542);
and U875 (N_875,In_916,In_14);
nor U876 (N_876,In_590,In_734);
or U877 (N_877,In_478,In_781);
nand U878 (N_878,In_317,In_925);
xor U879 (N_879,In_247,In_815);
xor U880 (N_880,In_592,In_419);
nor U881 (N_881,In_627,In_971);
or U882 (N_882,In_737,In_622);
xnor U883 (N_883,In_570,In_821);
or U884 (N_884,In_545,In_429);
xnor U885 (N_885,In_753,In_884);
xnor U886 (N_886,In_910,In_924);
nor U887 (N_887,In_181,In_705);
xor U888 (N_888,In_236,In_333);
nand U889 (N_889,In_140,In_836);
nand U890 (N_890,In_568,In_31);
nand U891 (N_891,In_571,In_970);
nor U892 (N_892,In_649,In_701);
nand U893 (N_893,In_448,In_443);
nand U894 (N_894,In_479,In_136);
and U895 (N_895,In_686,In_292);
or U896 (N_896,In_650,In_324);
xor U897 (N_897,In_125,In_982);
or U898 (N_898,In_60,In_555);
nand U899 (N_899,In_773,In_713);
and U900 (N_900,In_520,In_364);
or U901 (N_901,In_748,In_105);
and U902 (N_902,In_19,In_588);
and U903 (N_903,In_705,In_68);
nor U904 (N_904,In_625,In_483);
nand U905 (N_905,In_20,In_931);
and U906 (N_906,In_893,In_313);
and U907 (N_907,In_748,In_213);
nand U908 (N_908,In_697,In_230);
nor U909 (N_909,In_171,In_57);
nand U910 (N_910,In_62,In_297);
xor U911 (N_911,In_328,In_300);
xnor U912 (N_912,In_142,In_787);
nand U913 (N_913,In_525,In_158);
nand U914 (N_914,In_24,In_520);
nor U915 (N_915,In_151,In_649);
and U916 (N_916,In_33,In_503);
or U917 (N_917,In_136,In_130);
or U918 (N_918,In_305,In_393);
and U919 (N_919,In_169,In_939);
nand U920 (N_920,In_318,In_943);
xor U921 (N_921,In_418,In_532);
or U922 (N_922,In_881,In_239);
xnor U923 (N_923,In_703,In_429);
nand U924 (N_924,In_569,In_492);
xor U925 (N_925,In_315,In_299);
xnor U926 (N_926,In_734,In_687);
nor U927 (N_927,In_611,In_973);
xnor U928 (N_928,In_517,In_790);
and U929 (N_929,In_619,In_374);
and U930 (N_930,In_491,In_854);
and U931 (N_931,In_994,In_654);
xnor U932 (N_932,In_107,In_78);
and U933 (N_933,In_963,In_950);
and U934 (N_934,In_555,In_478);
xnor U935 (N_935,In_645,In_446);
and U936 (N_936,In_716,In_370);
nand U937 (N_937,In_945,In_965);
or U938 (N_938,In_41,In_737);
or U939 (N_939,In_49,In_243);
nand U940 (N_940,In_84,In_839);
nand U941 (N_941,In_942,In_980);
xnor U942 (N_942,In_293,In_349);
xor U943 (N_943,In_515,In_298);
and U944 (N_944,In_942,In_281);
xor U945 (N_945,In_97,In_402);
and U946 (N_946,In_769,In_120);
and U947 (N_947,In_357,In_246);
nor U948 (N_948,In_163,In_792);
nor U949 (N_949,In_88,In_634);
nor U950 (N_950,In_238,In_177);
xor U951 (N_951,In_496,In_746);
or U952 (N_952,In_605,In_461);
xnor U953 (N_953,In_837,In_289);
or U954 (N_954,In_309,In_690);
or U955 (N_955,In_661,In_938);
nand U956 (N_956,In_252,In_354);
or U957 (N_957,In_549,In_703);
or U958 (N_958,In_845,In_839);
and U959 (N_959,In_642,In_834);
nor U960 (N_960,In_465,In_649);
or U961 (N_961,In_571,In_454);
or U962 (N_962,In_349,In_683);
or U963 (N_963,In_489,In_606);
and U964 (N_964,In_965,In_750);
xnor U965 (N_965,In_753,In_984);
or U966 (N_966,In_946,In_320);
xor U967 (N_967,In_259,In_716);
nand U968 (N_968,In_3,In_738);
nor U969 (N_969,In_391,In_592);
or U970 (N_970,In_79,In_32);
and U971 (N_971,In_902,In_119);
or U972 (N_972,In_362,In_833);
or U973 (N_973,In_898,In_438);
and U974 (N_974,In_418,In_653);
or U975 (N_975,In_219,In_638);
nor U976 (N_976,In_839,In_490);
or U977 (N_977,In_80,In_399);
and U978 (N_978,In_330,In_482);
and U979 (N_979,In_749,In_295);
and U980 (N_980,In_969,In_330);
nor U981 (N_981,In_506,In_839);
xor U982 (N_982,In_113,In_39);
nand U983 (N_983,In_189,In_284);
or U984 (N_984,In_412,In_148);
nand U985 (N_985,In_316,In_295);
nor U986 (N_986,In_416,In_511);
or U987 (N_987,In_962,In_968);
xnor U988 (N_988,In_571,In_190);
nor U989 (N_989,In_49,In_694);
and U990 (N_990,In_678,In_705);
nor U991 (N_991,In_930,In_850);
or U992 (N_992,In_724,In_640);
and U993 (N_993,In_806,In_831);
and U994 (N_994,In_142,In_560);
nand U995 (N_995,In_294,In_715);
or U996 (N_996,In_581,In_329);
nand U997 (N_997,In_710,In_252);
and U998 (N_998,In_746,In_222);
nor U999 (N_999,In_844,In_274);
nand U1000 (N_1000,N_163,N_18);
or U1001 (N_1001,N_0,N_588);
nand U1002 (N_1002,N_221,N_944);
or U1003 (N_1003,N_204,N_336);
nand U1004 (N_1004,N_430,N_520);
and U1005 (N_1005,N_749,N_586);
and U1006 (N_1006,N_122,N_15);
nor U1007 (N_1007,N_128,N_503);
nand U1008 (N_1008,N_864,N_264);
xor U1009 (N_1009,N_350,N_528);
and U1010 (N_1010,N_142,N_306);
nor U1011 (N_1011,N_370,N_120);
nand U1012 (N_1012,N_810,N_705);
and U1013 (N_1013,N_923,N_470);
nor U1014 (N_1014,N_140,N_73);
and U1015 (N_1015,N_80,N_595);
xor U1016 (N_1016,N_486,N_517);
nor U1017 (N_1017,N_628,N_364);
nand U1018 (N_1018,N_970,N_507);
and U1019 (N_1019,N_324,N_622);
nand U1020 (N_1020,N_19,N_937);
nand U1021 (N_1021,N_183,N_434);
nand U1022 (N_1022,N_375,N_292);
or U1023 (N_1023,N_687,N_621);
nor U1024 (N_1024,N_669,N_405);
nand U1025 (N_1025,N_900,N_935);
nor U1026 (N_1026,N_360,N_514);
or U1027 (N_1027,N_872,N_524);
nand U1028 (N_1028,N_270,N_545);
and U1029 (N_1029,N_881,N_340);
xor U1030 (N_1030,N_368,N_388);
or U1031 (N_1031,N_485,N_400);
nor U1032 (N_1032,N_309,N_831);
xor U1033 (N_1033,N_420,N_167);
nor U1034 (N_1034,N_195,N_521);
xnor U1035 (N_1035,N_487,N_263);
and U1036 (N_1036,N_236,N_266);
or U1037 (N_1037,N_206,N_158);
or U1038 (N_1038,N_9,N_982);
or U1039 (N_1039,N_413,N_700);
nor U1040 (N_1040,N_753,N_801);
nand U1041 (N_1041,N_65,N_876);
and U1042 (N_1042,N_768,N_216);
nor U1043 (N_1043,N_180,N_160);
and U1044 (N_1044,N_22,N_869);
and U1045 (N_1045,N_693,N_76);
or U1046 (N_1046,N_792,N_232);
and U1047 (N_1047,N_566,N_969);
nand U1048 (N_1048,N_543,N_882);
or U1049 (N_1049,N_387,N_680);
or U1050 (N_1050,N_722,N_793);
xnor U1051 (N_1051,N_251,N_157);
and U1052 (N_1052,N_377,N_534);
xnor U1053 (N_1053,N_150,N_636);
and U1054 (N_1054,N_352,N_629);
nor U1055 (N_1055,N_562,N_772);
xor U1056 (N_1056,N_980,N_96);
nor U1057 (N_1057,N_519,N_525);
and U1058 (N_1058,N_369,N_974);
xor U1059 (N_1059,N_919,N_593);
or U1060 (N_1060,N_94,N_452);
nor U1061 (N_1061,N_690,N_911);
nor U1062 (N_1062,N_408,N_963);
nor U1063 (N_1063,N_590,N_613);
xor U1064 (N_1064,N_939,N_426);
xnor U1065 (N_1065,N_783,N_604);
or U1066 (N_1066,N_657,N_927);
or U1067 (N_1067,N_274,N_343);
nor U1068 (N_1068,N_776,N_45);
nand U1069 (N_1069,N_741,N_995);
and U1070 (N_1070,N_798,N_223);
or U1071 (N_1071,N_956,N_288);
nand U1072 (N_1072,N_345,N_24);
and U1073 (N_1073,N_91,N_5);
nor U1074 (N_1074,N_250,N_746);
nand U1075 (N_1075,N_111,N_536);
nor U1076 (N_1076,N_500,N_946);
nand U1077 (N_1077,N_666,N_63);
nand U1078 (N_1078,N_713,N_284);
and U1079 (N_1079,N_589,N_255);
xnor U1080 (N_1080,N_422,N_253);
nor U1081 (N_1081,N_269,N_162);
nand U1082 (N_1082,N_126,N_668);
nor U1083 (N_1083,N_925,N_121);
nor U1084 (N_1084,N_461,N_124);
and U1085 (N_1085,N_763,N_349);
nand U1086 (N_1086,N_540,N_197);
and U1087 (N_1087,N_610,N_782);
nand U1088 (N_1088,N_698,N_809);
or U1089 (N_1089,N_551,N_703);
xnor U1090 (N_1090,N_196,N_720);
nor U1091 (N_1091,N_397,N_751);
and U1092 (N_1092,N_61,N_362);
and U1093 (N_1093,N_609,N_648);
or U1094 (N_1094,N_878,N_243);
xor U1095 (N_1095,N_635,N_846);
or U1096 (N_1096,N_338,N_228);
xor U1097 (N_1097,N_608,N_215);
nor U1098 (N_1098,N_110,N_897);
or U1099 (N_1099,N_415,N_737);
xor U1100 (N_1100,N_605,N_538);
nor U1101 (N_1101,N_407,N_456);
and U1102 (N_1102,N_78,N_978);
or U1103 (N_1103,N_219,N_52);
or U1104 (N_1104,N_342,N_254);
nor U1105 (N_1105,N_842,N_325);
or U1106 (N_1106,N_488,N_570);
nor U1107 (N_1107,N_615,N_733);
and U1108 (N_1108,N_748,N_957);
nand U1109 (N_1109,N_665,N_479);
or U1110 (N_1110,N_36,N_193);
xor U1111 (N_1111,N_619,N_135);
nand U1112 (N_1112,N_533,N_492);
or U1113 (N_1113,N_379,N_177);
nand U1114 (N_1114,N_996,N_976);
nor U1115 (N_1115,N_711,N_478);
or U1116 (N_1116,N_750,N_888);
nor U1117 (N_1117,N_164,N_468);
xnor U1118 (N_1118,N_189,N_473);
or U1119 (N_1119,N_752,N_27);
and U1120 (N_1120,N_743,N_355);
nor U1121 (N_1121,N_823,N_10);
and U1122 (N_1122,N_942,N_312);
or U1123 (N_1123,N_499,N_290);
nand U1124 (N_1124,N_912,N_418);
nor U1125 (N_1125,N_109,N_301);
and U1126 (N_1126,N_261,N_824);
or U1127 (N_1127,N_686,N_43);
xor U1128 (N_1128,N_267,N_887);
or U1129 (N_1129,N_639,N_244);
nor U1130 (N_1130,N_42,N_32);
xor U1131 (N_1131,N_527,N_439);
or U1132 (N_1132,N_116,N_159);
nor U1133 (N_1133,N_885,N_674);
nand U1134 (N_1134,N_424,N_522);
and U1135 (N_1135,N_363,N_186);
and U1136 (N_1136,N_715,N_175);
or U1137 (N_1137,N_248,N_154);
and U1138 (N_1138,N_392,N_817);
nor U1139 (N_1139,N_231,N_453);
and U1140 (N_1140,N_697,N_68);
and U1141 (N_1141,N_191,N_217);
and U1142 (N_1142,N_161,N_311);
nand U1143 (N_1143,N_575,N_282);
nand U1144 (N_1144,N_318,N_950);
or U1145 (N_1145,N_867,N_441);
nand U1146 (N_1146,N_74,N_707);
xor U1147 (N_1147,N_670,N_103);
nor U1148 (N_1148,N_786,N_239);
xor U1149 (N_1149,N_472,N_139);
xnor U1150 (N_1150,N_865,N_893);
nor U1151 (N_1151,N_509,N_726);
nand U1152 (N_1152,N_638,N_565);
nor U1153 (N_1153,N_483,N_184);
nand U1154 (N_1154,N_322,N_240);
nand U1155 (N_1155,N_378,N_922);
nor U1156 (N_1156,N_144,N_423);
and U1157 (N_1157,N_832,N_155);
or U1158 (N_1158,N_491,N_993);
xor U1159 (N_1159,N_417,N_141);
nor U1160 (N_1160,N_427,N_357);
and U1161 (N_1161,N_932,N_297);
xor U1162 (N_1162,N_553,N_779);
xor U1163 (N_1163,N_41,N_211);
nor U1164 (N_1164,N_884,N_818);
nand U1165 (N_1165,N_626,N_961);
nand U1166 (N_1166,N_904,N_469);
and U1167 (N_1167,N_11,N_403);
xnor U1168 (N_1168,N_745,N_477);
xnor U1169 (N_1169,N_300,N_170);
xor U1170 (N_1170,N_747,N_108);
nand U1171 (N_1171,N_834,N_572);
nor U1172 (N_1172,N_187,N_953);
nor U1173 (N_1173,N_774,N_257);
nand U1174 (N_1174,N_598,N_870);
nand U1175 (N_1175,N_755,N_879);
and U1176 (N_1176,N_765,N_383);
xor U1177 (N_1177,N_165,N_856);
or U1178 (N_1178,N_358,N_564);
nor U1179 (N_1179,N_637,N_596);
and U1180 (N_1180,N_280,N_848);
nand U1181 (N_1181,N_512,N_830);
nor U1182 (N_1182,N_172,N_718);
or U1183 (N_1183,N_356,N_857);
or U1184 (N_1184,N_808,N_148);
and U1185 (N_1185,N_716,N_320);
nor U1186 (N_1186,N_571,N_833);
xor U1187 (N_1187,N_394,N_855);
nor U1188 (N_1188,N_29,N_490);
xnor U1189 (N_1189,N_295,N_127);
and U1190 (N_1190,N_34,N_348);
and U1191 (N_1191,N_663,N_951);
and U1192 (N_1192,N_815,N_734);
and U1193 (N_1193,N_133,N_984);
or U1194 (N_1194,N_592,N_51);
nand U1195 (N_1195,N_178,N_278);
nand U1196 (N_1196,N_156,N_273);
nor U1197 (N_1197,N_652,N_436);
nand U1198 (N_1198,N_455,N_476);
nand U1199 (N_1199,N_134,N_729);
xor U1200 (N_1200,N_285,N_660);
xnor U1201 (N_1201,N_814,N_526);
nand U1202 (N_1202,N_676,N_242);
xor U1203 (N_1203,N_860,N_740);
or U1204 (N_1204,N_761,N_582);
xor U1205 (N_1205,N_497,N_560);
and U1206 (N_1206,N_992,N_84);
nor U1207 (N_1207,N_3,N_844);
and U1208 (N_1208,N_620,N_840);
and U1209 (N_1209,N_841,N_839);
xor U1210 (N_1210,N_849,N_907);
xor U1211 (N_1211,N_209,N_784);
or U1212 (N_1212,N_958,N_702);
or U1213 (N_1213,N_862,N_87);
and U1214 (N_1214,N_70,N_739);
xnor U1215 (N_1215,N_940,N_296);
nand U1216 (N_1216,N_112,N_401);
nand U1217 (N_1217,N_616,N_502);
nor U1218 (N_1218,N_853,N_495);
xor U1219 (N_1219,N_289,N_431);
or U1220 (N_1220,N_518,N_224);
nor U1221 (N_1221,N_307,N_442);
nor U1222 (N_1222,N_95,N_85);
nor U1223 (N_1223,N_113,N_554);
nand U1224 (N_1224,N_845,N_706);
or U1225 (N_1225,N_13,N_645);
xor U1226 (N_1226,N_218,N_308);
nor U1227 (N_1227,N_75,N_820);
nand U1228 (N_1228,N_901,N_825);
nand U1229 (N_1229,N_412,N_672);
or U1230 (N_1230,N_281,N_791);
nand U1231 (N_1231,N_460,N_339);
and U1232 (N_1232,N_353,N_769);
and U1233 (N_1233,N_396,N_754);
nand U1234 (N_1234,N_171,N_283);
nand U1235 (N_1235,N_760,N_544);
nand U1236 (N_1236,N_235,N_530);
nand U1237 (N_1237,N_37,N_130);
and U1238 (N_1238,N_771,N_123);
xnor U1239 (N_1239,N_661,N_125);
nor U1240 (N_1240,N_173,N_2);
and U1241 (N_1241,N_188,N_354);
nand U1242 (N_1242,N_410,N_515);
and U1243 (N_1243,N_268,N_416);
nand U1244 (N_1244,N_12,N_316);
nand U1245 (N_1245,N_458,N_971);
nand U1246 (N_1246,N_973,N_484);
nand U1247 (N_1247,N_438,N_989);
xnor U1248 (N_1248,N_105,N_730);
or U1249 (N_1249,N_249,N_678);
xnor U1250 (N_1250,N_229,N_291);
or U1251 (N_1251,N_185,N_265);
nand U1252 (N_1252,N_151,N_641);
xnor U1253 (N_1253,N_714,N_828);
nor U1254 (N_1254,N_975,N_895);
nor U1255 (N_1255,N_398,N_909);
and U1256 (N_1256,N_153,N_797);
nor U1257 (N_1257,N_738,N_618);
and U1258 (N_1258,N_914,N_463);
and U1259 (N_1259,N_933,N_928);
nor U1260 (N_1260,N_480,N_640);
or U1261 (N_1261,N_505,N_335);
nor U1262 (N_1262,N_573,N_181);
and U1263 (N_1263,N_179,N_894);
nand U1264 (N_1264,N_321,N_756);
nor U1265 (N_1265,N_938,N_25);
and U1266 (N_1266,N_998,N_777);
or U1267 (N_1267,N_220,N_552);
nor U1268 (N_1268,N_843,N_959);
or U1269 (N_1269,N_835,N_137);
nand U1270 (N_1270,N_145,N_651);
nand U1271 (N_1271,N_685,N_174);
nor U1272 (N_1272,N_117,N_532);
xor U1273 (N_1273,N_81,N_952);
nor U1274 (N_1274,N_39,N_599);
nand U1275 (N_1275,N_447,N_802);
or U1276 (N_1276,N_868,N_448);
xor U1277 (N_1277,N_40,N_631);
and U1278 (N_1278,N_16,N_908);
nor U1279 (N_1279,N_333,N_395);
and U1280 (N_1280,N_459,N_723);
nor U1281 (N_1281,N_892,N_205);
nor U1282 (N_1282,N_757,N_446);
and U1283 (N_1283,N_207,N_812);
nand U1284 (N_1284,N_365,N_851);
xnor U1285 (N_1285,N_227,N_617);
nand U1286 (N_1286,N_773,N_539);
xnor U1287 (N_1287,N_82,N_129);
nand U1288 (N_1288,N_688,N_577);
and U1289 (N_1289,N_567,N_866);
xor U1290 (N_1290,N_531,N_132);
and U1291 (N_1291,N_918,N_385);
nand U1292 (N_1292,N_762,N_708);
xor U1293 (N_1293,N_930,N_276);
or U1294 (N_1294,N_667,N_508);
nand U1295 (N_1295,N_147,N_390);
xnor U1296 (N_1296,N_489,N_838);
nor U1297 (N_1297,N_1,N_404);
or U1298 (N_1298,N_241,N_71);
or U1299 (N_1299,N_38,N_656);
nand U1300 (N_1300,N_948,N_168);
nor U1301 (N_1301,N_587,N_766);
nand U1302 (N_1302,N_896,N_556);
xnor U1303 (N_1303,N_684,N_921);
xor U1304 (N_1304,N_778,N_591);
and U1305 (N_1305,N_481,N_561);
nand U1306 (N_1306,N_329,N_985);
xor U1307 (N_1307,N_262,N_361);
and U1308 (N_1308,N_433,N_298);
or U1309 (N_1309,N_934,N_977);
and U1310 (N_1310,N_585,N_854);
nand U1311 (N_1311,N_941,N_192);
or U1312 (N_1312,N_601,N_863);
nor U1313 (N_1313,N_60,N_633);
nand U1314 (N_1314,N_880,N_146);
xor U1315 (N_1315,N_376,N_107);
nor U1316 (N_1316,N_787,N_719);
nand U1317 (N_1317,N_813,N_47);
xor U1318 (N_1318,N_114,N_28);
and U1319 (N_1319,N_317,N_612);
or U1320 (N_1320,N_198,N_683);
xnor U1321 (N_1321,N_381,N_821);
or U1322 (N_1322,N_371,N_859);
nor U1323 (N_1323,N_873,N_917);
nor U1324 (N_1324,N_359,N_366);
xor U1325 (N_1325,N_482,N_64);
or U1326 (N_1326,N_576,N_981);
xor U1327 (N_1327,N_389,N_910);
or U1328 (N_1328,N_331,N_245);
and U1329 (N_1329,N_54,N_315);
xnor U1330 (N_1330,N_557,N_546);
and U1331 (N_1331,N_658,N_537);
nor U1332 (N_1332,N_454,N_351);
or U1333 (N_1333,N_600,N_102);
nor U1334 (N_1334,N_194,N_451);
and U1335 (N_1335,N_563,N_891);
xnor U1336 (N_1336,N_97,N_962);
nand U1337 (N_1337,N_704,N_319);
or U1338 (N_1338,N_955,N_341);
or U1339 (N_1339,N_614,N_805);
nor U1340 (N_1340,N_504,N_31);
or U1341 (N_1341,N_474,N_653);
xor U1342 (N_1342,N_679,N_875);
nand U1343 (N_1343,N_393,N_735);
xnor U1344 (N_1344,N_682,N_304);
and U1345 (N_1345,N_437,N_926);
xnor U1346 (N_1346,N_212,N_541);
and U1347 (N_1347,N_166,N_579);
or U1348 (N_1348,N_201,N_428);
or U1349 (N_1349,N_644,N_799);
or U1350 (N_1350,N_69,N_230);
or U1351 (N_1351,N_380,N_202);
nor U1352 (N_1352,N_347,N_374);
xnor U1353 (N_1353,N_569,N_681);
nor U1354 (N_1354,N_496,N_991);
or U1355 (N_1355,N_529,N_924);
xor U1356 (N_1356,N_983,N_581);
and U1357 (N_1357,N_988,N_252);
nor U1358 (N_1358,N_929,N_247);
or U1359 (N_1359,N_513,N_190);
xor U1360 (N_1360,N_886,N_21);
or U1361 (N_1361,N_964,N_997);
nor U1362 (N_1362,N_829,N_293);
nand U1363 (N_1363,N_344,N_501);
or U1364 (N_1364,N_429,N_119);
xor U1365 (N_1365,N_313,N_987);
xor U1366 (N_1366,N_234,N_465);
xor U1367 (N_1367,N_66,N_449);
or U1368 (N_1368,N_664,N_643);
xor U1369 (N_1369,N_79,N_99);
nand U1370 (N_1370,N_258,N_182);
nor U1371 (N_1371,N_717,N_852);
or U1372 (N_1372,N_889,N_804);
nand U1373 (N_1373,N_33,N_920);
xnor U1374 (N_1374,N_386,N_35);
xor U1375 (N_1375,N_56,N_999);
or U1376 (N_1376,N_673,N_90);
and U1377 (N_1377,N_506,N_542);
xnor U1378 (N_1378,N_568,N_816);
or U1379 (N_1379,N_945,N_7);
xor U1380 (N_1380,N_384,N_583);
and U1381 (N_1381,N_334,N_26);
xor U1382 (N_1382,N_770,N_642);
or U1383 (N_1383,N_811,N_203);
nand U1384 (N_1384,N_523,N_535);
nor U1385 (N_1385,N_106,N_943);
and U1386 (N_1386,N_607,N_548);
nor U1387 (N_1387,N_256,N_822);
xnor U1388 (N_1388,N_314,N_837);
and U1389 (N_1389,N_781,N_382);
nor U1390 (N_1390,N_819,N_391);
xor U1391 (N_1391,N_649,N_493);
nor U1392 (N_1392,N_800,N_287);
nand U1393 (N_1393,N_86,N_712);
xnor U1394 (N_1394,N_225,N_406);
or U1395 (N_1395,N_55,N_93);
nand U1396 (N_1396,N_602,N_915);
nor U1397 (N_1397,N_411,N_467);
xor U1398 (N_1398,N_214,N_694);
and U1399 (N_1399,N_623,N_659);
or U1400 (N_1400,N_584,N_871);
and U1401 (N_1401,N_947,N_731);
nor U1402 (N_1402,N_850,N_440);
nand U1403 (N_1403,N_104,N_625);
nand U1404 (N_1404,N_302,N_580);
or U1405 (N_1405,N_632,N_421);
or U1406 (N_1406,N_803,N_332);
nor U1407 (N_1407,N_775,N_858);
xor U1408 (N_1408,N_30,N_990);
nand U1409 (N_1409,N_624,N_699);
nand U1410 (N_1410,N_445,N_960);
nand U1411 (N_1411,N_100,N_200);
or U1412 (N_1412,N_138,N_20);
and U1413 (N_1413,N_701,N_728);
or U1414 (N_1414,N_899,N_710);
or U1415 (N_1415,N_330,N_603);
and U1416 (N_1416,N_905,N_326);
or U1417 (N_1417,N_471,N_443);
nand U1418 (N_1418,N_827,N_727);
and U1419 (N_1419,N_795,N_965);
nand U1420 (N_1420,N_611,N_550);
nand U1421 (N_1421,N_402,N_210);
xor U1422 (N_1422,N_14,N_758);
or U1423 (N_1423,N_709,N_294);
and U1424 (N_1424,N_464,N_372);
and U1425 (N_1425,N_647,N_780);
or U1426 (N_1426,N_689,N_399);
or U1427 (N_1427,N_597,N_494);
xor U1428 (N_1428,N_305,N_246);
nor U1429 (N_1429,N_6,N_986);
nand U1430 (N_1430,N_936,N_691);
nor U1431 (N_1431,N_498,N_675);
nor U1432 (N_1432,N_725,N_898);
or U1433 (N_1433,N_655,N_692);
and U1434 (N_1434,N_627,N_271);
nand U1435 (N_1435,N_732,N_303);
xor U1436 (N_1436,N_299,N_83);
nand U1437 (N_1437,N_67,N_574);
nand U1438 (N_1438,N_346,N_475);
and U1439 (N_1439,N_58,N_367);
nor U1440 (N_1440,N_511,N_260);
xnor U1441 (N_1441,N_890,N_199);
nor U1442 (N_1442,N_606,N_444);
nor U1443 (N_1443,N_466,N_373);
or U1444 (N_1444,N_759,N_213);
nor U1445 (N_1445,N_59,N_883);
nand U1446 (N_1446,N_435,N_238);
or U1447 (N_1447,N_237,N_419);
xnor U1448 (N_1448,N_549,N_4);
and U1449 (N_1449,N_861,N_796);
xnor U1450 (N_1450,N_8,N_516);
xnor U1451 (N_1451,N_662,N_337);
xnor U1452 (N_1452,N_874,N_323);
nand U1453 (N_1453,N_695,N_457);
or U1454 (N_1454,N_902,N_630);
or U1455 (N_1455,N_877,N_767);
and U1456 (N_1456,N_88,N_559);
and U1457 (N_1457,N_115,N_57);
nor U1458 (N_1458,N_696,N_98);
or U1459 (N_1459,N_510,N_806);
nor U1460 (N_1460,N_222,N_259);
xor U1461 (N_1461,N_48,N_46);
and U1462 (N_1462,N_555,N_450);
nor U1463 (N_1463,N_736,N_966);
nand U1464 (N_1464,N_578,N_328);
xnor U1465 (N_1465,N_547,N_594);
nand U1466 (N_1466,N_788,N_903);
or U1467 (N_1467,N_906,N_931);
xor U1468 (N_1468,N_916,N_176);
nand U1469 (N_1469,N_77,N_826);
xor U1470 (N_1470,N_101,N_967);
nor U1471 (N_1471,N_310,N_789);
and U1472 (N_1472,N_994,N_272);
nor U1473 (N_1473,N_462,N_275);
or U1474 (N_1474,N_72,N_89);
nor U1475 (N_1475,N_979,N_62);
xor U1476 (N_1476,N_169,N_646);
nor U1477 (N_1477,N_954,N_277);
and U1478 (N_1478,N_949,N_742);
and U1479 (N_1479,N_634,N_847);
xor U1480 (N_1480,N_136,N_409);
or U1481 (N_1481,N_233,N_744);
and U1482 (N_1482,N_44,N_53);
nand U1483 (N_1483,N_968,N_50);
nor U1484 (N_1484,N_226,N_721);
or U1485 (N_1485,N_414,N_92);
xor U1486 (N_1486,N_671,N_432);
or U1487 (N_1487,N_208,N_558);
or U1488 (N_1488,N_764,N_913);
xor U1489 (N_1489,N_327,N_972);
and U1490 (N_1490,N_118,N_425);
and U1491 (N_1491,N_149,N_49);
and U1492 (N_1492,N_677,N_836);
nor U1493 (N_1493,N_279,N_152);
nand U1494 (N_1494,N_724,N_286);
xnor U1495 (N_1495,N_807,N_23);
and U1496 (N_1496,N_794,N_131);
nor U1497 (N_1497,N_650,N_654);
and U1498 (N_1498,N_143,N_790);
xor U1499 (N_1499,N_785,N_17);
nand U1500 (N_1500,N_780,N_577);
and U1501 (N_1501,N_997,N_310);
nand U1502 (N_1502,N_483,N_284);
nor U1503 (N_1503,N_843,N_616);
xor U1504 (N_1504,N_586,N_15);
and U1505 (N_1505,N_246,N_70);
or U1506 (N_1506,N_598,N_922);
nand U1507 (N_1507,N_645,N_682);
and U1508 (N_1508,N_252,N_265);
nand U1509 (N_1509,N_299,N_880);
nor U1510 (N_1510,N_318,N_656);
or U1511 (N_1511,N_980,N_997);
nor U1512 (N_1512,N_752,N_878);
or U1513 (N_1513,N_341,N_772);
nand U1514 (N_1514,N_465,N_644);
nor U1515 (N_1515,N_897,N_458);
xor U1516 (N_1516,N_476,N_379);
nand U1517 (N_1517,N_104,N_282);
nand U1518 (N_1518,N_663,N_308);
nand U1519 (N_1519,N_683,N_102);
xor U1520 (N_1520,N_157,N_396);
nand U1521 (N_1521,N_830,N_672);
xor U1522 (N_1522,N_224,N_39);
and U1523 (N_1523,N_903,N_386);
nand U1524 (N_1524,N_96,N_249);
and U1525 (N_1525,N_115,N_445);
or U1526 (N_1526,N_874,N_970);
and U1527 (N_1527,N_283,N_395);
and U1528 (N_1528,N_968,N_12);
and U1529 (N_1529,N_872,N_468);
nand U1530 (N_1530,N_76,N_340);
nand U1531 (N_1531,N_467,N_67);
and U1532 (N_1532,N_956,N_265);
and U1533 (N_1533,N_86,N_106);
xnor U1534 (N_1534,N_855,N_684);
nand U1535 (N_1535,N_846,N_842);
xnor U1536 (N_1536,N_948,N_774);
xnor U1537 (N_1537,N_257,N_360);
nor U1538 (N_1538,N_687,N_823);
or U1539 (N_1539,N_593,N_100);
and U1540 (N_1540,N_291,N_523);
nand U1541 (N_1541,N_798,N_276);
and U1542 (N_1542,N_597,N_537);
nor U1543 (N_1543,N_122,N_575);
and U1544 (N_1544,N_475,N_642);
and U1545 (N_1545,N_433,N_135);
nor U1546 (N_1546,N_551,N_106);
nor U1547 (N_1547,N_291,N_801);
and U1548 (N_1548,N_283,N_995);
xnor U1549 (N_1549,N_186,N_69);
nor U1550 (N_1550,N_109,N_154);
and U1551 (N_1551,N_190,N_903);
nor U1552 (N_1552,N_594,N_337);
and U1553 (N_1553,N_521,N_442);
and U1554 (N_1554,N_630,N_934);
or U1555 (N_1555,N_945,N_585);
and U1556 (N_1556,N_668,N_343);
xor U1557 (N_1557,N_533,N_777);
nand U1558 (N_1558,N_334,N_624);
nor U1559 (N_1559,N_898,N_635);
and U1560 (N_1560,N_97,N_777);
xnor U1561 (N_1561,N_388,N_226);
and U1562 (N_1562,N_626,N_867);
nor U1563 (N_1563,N_255,N_415);
nand U1564 (N_1564,N_544,N_107);
and U1565 (N_1565,N_64,N_919);
or U1566 (N_1566,N_849,N_479);
nand U1567 (N_1567,N_198,N_477);
nor U1568 (N_1568,N_784,N_739);
or U1569 (N_1569,N_679,N_409);
or U1570 (N_1570,N_559,N_658);
nor U1571 (N_1571,N_276,N_555);
and U1572 (N_1572,N_916,N_741);
nor U1573 (N_1573,N_417,N_525);
nor U1574 (N_1574,N_504,N_636);
nor U1575 (N_1575,N_704,N_1);
xnor U1576 (N_1576,N_581,N_984);
and U1577 (N_1577,N_935,N_429);
nor U1578 (N_1578,N_330,N_323);
and U1579 (N_1579,N_108,N_421);
or U1580 (N_1580,N_493,N_168);
xnor U1581 (N_1581,N_155,N_703);
xor U1582 (N_1582,N_901,N_584);
or U1583 (N_1583,N_135,N_570);
and U1584 (N_1584,N_898,N_57);
and U1585 (N_1585,N_607,N_596);
xor U1586 (N_1586,N_908,N_718);
nor U1587 (N_1587,N_433,N_512);
xnor U1588 (N_1588,N_431,N_9);
or U1589 (N_1589,N_481,N_928);
and U1590 (N_1590,N_600,N_367);
or U1591 (N_1591,N_515,N_572);
or U1592 (N_1592,N_844,N_695);
nand U1593 (N_1593,N_790,N_461);
nor U1594 (N_1594,N_451,N_174);
nor U1595 (N_1595,N_437,N_607);
and U1596 (N_1596,N_942,N_365);
or U1597 (N_1597,N_470,N_319);
and U1598 (N_1598,N_896,N_595);
nand U1599 (N_1599,N_122,N_907);
nor U1600 (N_1600,N_622,N_341);
nand U1601 (N_1601,N_809,N_625);
nor U1602 (N_1602,N_777,N_188);
or U1603 (N_1603,N_939,N_788);
and U1604 (N_1604,N_179,N_544);
or U1605 (N_1605,N_237,N_856);
nor U1606 (N_1606,N_532,N_119);
xnor U1607 (N_1607,N_857,N_353);
nand U1608 (N_1608,N_722,N_19);
nand U1609 (N_1609,N_723,N_440);
or U1610 (N_1610,N_758,N_590);
or U1611 (N_1611,N_392,N_717);
and U1612 (N_1612,N_408,N_589);
nand U1613 (N_1613,N_467,N_136);
and U1614 (N_1614,N_313,N_40);
nor U1615 (N_1615,N_950,N_725);
and U1616 (N_1616,N_16,N_830);
xor U1617 (N_1617,N_671,N_687);
nand U1618 (N_1618,N_696,N_438);
or U1619 (N_1619,N_298,N_631);
nor U1620 (N_1620,N_95,N_590);
xnor U1621 (N_1621,N_664,N_736);
nand U1622 (N_1622,N_215,N_601);
nor U1623 (N_1623,N_610,N_943);
nand U1624 (N_1624,N_827,N_533);
and U1625 (N_1625,N_421,N_500);
and U1626 (N_1626,N_574,N_14);
xor U1627 (N_1627,N_335,N_869);
nor U1628 (N_1628,N_359,N_188);
xor U1629 (N_1629,N_246,N_315);
nor U1630 (N_1630,N_304,N_780);
and U1631 (N_1631,N_776,N_26);
xnor U1632 (N_1632,N_777,N_604);
xor U1633 (N_1633,N_270,N_442);
or U1634 (N_1634,N_160,N_805);
and U1635 (N_1635,N_444,N_81);
nor U1636 (N_1636,N_975,N_287);
or U1637 (N_1637,N_963,N_956);
nand U1638 (N_1638,N_776,N_181);
nand U1639 (N_1639,N_17,N_885);
nor U1640 (N_1640,N_74,N_688);
nor U1641 (N_1641,N_108,N_324);
nor U1642 (N_1642,N_924,N_741);
nor U1643 (N_1643,N_111,N_0);
xnor U1644 (N_1644,N_243,N_40);
or U1645 (N_1645,N_288,N_525);
and U1646 (N_1646,N_530,N_37);
and U1647 (N_1647,N_558,N_319);
or U1648 (N_1648,N_149,N_779);
and U1649 (N_1649,N_671,N_179);
xor U1650 (N_1650,N_124,N_480);
or U1651 (N_1651,N_980,N_85);
nand U1652 (N_1652,N_119,N_283);
or U1653 (N_1653,N_649,N_989);
nand U1654 (N_1654,N_297,N_567);
or U1655 (N_1655,N_141,N_689);
or U1656 (N_1656,N_459,N_113);
nand U1657 (N_1657,N_308,N_512);
or U1658 (N_1658,N_839,N_297);
and U1659 (N_1659,N_268,N_448);
or U1660 (N_1660,N_466,N_23);
and U1661 (N_1661,N_319,N_200);
or U1662 (N_1662,N_255,N_128);
and U1663 (N_1663,N_971,N_846);
nand U1664 (N_1664,N_377,N_853);
nor U1665 (N_1665,N_934,N_695);
nand U1666 (N_1666,N_469,N_645);
nand U1667 (N_1667,N_573,N_419);
nand U1668 (N_1668,N_95,N_914);
nand U1669 (N_1669,N_211,N_833);
nor U1670 (N_1670,N_998,N_989);
xor U1671 (N_1671,N_603,N_379);
nand U1672 (N_1672,N_77,N_307);
and U1673 (N_1673,N_80,N_189);
or U1674 (N_1674,N_243,N_244);
xor U1675 (N_1675,N_641,N_400);
or U1676 (N_1676,N_142,N_97);
nor U1677 (N_1677,N_972,N_588);
xnor U1678 (N_1678,N_635,N_413);
or U1679 (N_1679,N_44,N_539);
or U1680 (N_1680,N_505,N_663);
nor U1681 (N_1681,N_76,N_575);
or U1682 (N_1682,N_715,N_268);
nand U1683 (N_1683,N_166,N_789);
or U1684 (N_1684,N_371,N_405);
xor U1685 (N_1685,N_731,N_467);
and U1686 (N_1686,N_944,N_347);
xnor U1687 (N_1687,N_569,N_42);
or U1688 (N_1688,N_234,N_499);
nor U1689 (N_1689,N_9,N_51);
nand U1690 (N_1690,N_714,N_521);
or U1691 (N_1691,N_731,N_350);
nand U1692 (N_1692,N_525,N_550);
xor U1693 (N_1693,N_459,N_429);
or U1694 (N_1694,N_168,N_880);
and U1695 (N_1695,N_752,N_743);
and U1696 (N_1696,N_663,N_561);
xnor U1697 (N_1697,N_576,N_915);
nand U1698 (N_1698,N_160,N_111);
and U1699 (N_1699,N_770,N_72);
or U1700 (N_1700,N_114,N_922);
nand U1701 (N_1701,N_991,N_239);
xor U1702 (N_1702,N_156,N_936);
nand U1703 (N_1703,N_89,N_560);
and U1704 (N_1704,N_209,N_819);
or U1705 (N_1705,N_405,N_59);
nand U1706 (N_1706,N_918,N_664);
or U1707 (N_1707,N_409,N_757);
xnor U1708 (N_1708,N_126,N_915);
or U1709 (N_1709,N_949,N_339);
xnor U1710 (N_1710,N_234,N_949);
and U1711 (N_1711,N_515,N_283);
nor U1712 (N_1712,N_882,N_3);
or U1713 (N_1713,N_118,N_98);
or U1714 (N_1714,N_503,N_409);
xor U1715 (N_1715,N_591,N_696);
nand U1716 (N_1716,N_882,N_490);
nand U1717 (N_1717,N_188,N_723);
or U1718 (N_1718,N_474,N_441);
nand U1719 (N_1719,N_603,N_163);
nand U1720 (N_1720,N_802,N_548);
nand U1721 (N_1721,N_267,N_425);
or U1722 (N_1722,N_958,N_566);
nor U1723 (N_1723,N_524,N_945);
or U1724 (N_1724,N_913,N_993);
xor U1725 (N_1725,N_461,N_44);
nand U1726 (N_1726,N_55,N_596);
or U1727 (N_1727,N_457,N_150);
nor U1728 (N_1728,N_128,N_292);
xor U1729 (N_1729,N_740,N_741);
or U1730 (N_1730,N_721,N_686);
xor U1731 (N_1731,N_679,N_933);
xor U1732 (N_1732,N_350,N_946);
xor U1733 (N_1733,N_335,N_543);
and U1734 (N_1734,N_168,N_110);
or U1735 (N_1735,N_953,N_160);
or U1736 (N_1736,N_397,N_745);
nand U1737 (N_1737,N_894,N_912);
and U1738 (N_1738,N_484,N_171);
or U1739 (N_1739,N_746,N_989);
nand U1740 (N_1740,N_822,N_55);
or U1741 (N_1741,N_876,N_913);
xor U1742 (N_1742,N_507,N_169);
xnor U1743 (N_1743,N_389,N_671);
nor U1744 (N_1744,N_431,N_428);
nand U1745 (N_1745,N_886,N_668);
nor U1746 (N_1746,N_877,N_992);
nand U1747 (N_1747,N_580,N_989);
or U1748 (N_1748,N_783,N_955);
or U1749 (N_1749,N_75,N_410);
xnor U1750 (N_1750,N_693,N_467);
and U1751 (N_1751,N_0,N_105);
or U1752 (N_1752,N_941,N_277);
nand U1753 (N_1753,N_388,N_547);
or U1754 (N_1754,N_776,N_194);
nor U1755 (N_1755,N_899,N_494);
nand U1756 (N_1756,N_883,N_127);
nor U1757 (N_1757,N_610,N_406);
nand U1758 (N_1758,N_33,N_646);
nand U1759 (N_1759,N_511,N_422);
or U1760 (N_1760,N_62,N_875);
or U1761 (N_1761,N_509,N_202);
xnor U1762 (N_1762,N_223,N_655);
or U1763 (N_1763,N_762,N_105);
and U1764 (N_1764,N_462,N_463);
and U1765 (N_1765,N_46,N_683);
and U1766 (N_1766,N_31,N_160);
xnor U1767 (N_1767,N_678,N_465);
xnor U1768 (N_1768,N_781,N_480);
xor U1769 (N_1769,N_323,N_536);
and U1770 (N_1770,N_149,N_575);
nand U1771 (N_1771,N_336,N_976);
or U1772 (N_1772,N_327,N_21);
nor U1773 (N_1773,N_454,N_743);
nor U1774 (N_1774,N_411,N_802);
or U1775 (N_1775,N_58,N_830);
nor U1776 (N_1776,N_249,N_431);
nand U1777 (N_1777,N_510,N_284);
or U1778 (N_1778,N_981,N_432);
and U1779 (N_1779,N_433,N_422);
xor U1780 (N_1780,N_360,N_187);
and U1781 (N_1781,N_136,N_371);
nand U1782 (N_1782,N_52,N_359);
nor U1783 (N_1783,N_70,N_244);
nand U1784 (N_1784,N_982,N_556);
and U1785 (N_1785,N_972,N_119);
or U1786 (N_1786,N_7,N_405);
nand U1787 (N_1787,N_267,N_256);
and U1788 (N_1788,N_42,N_187);
nor U1789 (N_1789,N_463,N_955);
or U1790 (N_1790,N_650,N_900);
or U1791 (N_1791,N_685,N_544);
or U1792 (N_1792,N_898,N_143);
or U1793 (N_1793,N_972,N_536);
nand U1794 (N_1794,N_898,N_296);
and U1795 (N_1795,N_219,N_475);
and U1796 (N_1796,N_984,N_609);
nand U1797 (N_1797,N_369,N_229);
nand U1798 (N_1798,N_87,N_855);
or U1799 (N_1799,N_465,N_25);
xor U1800 (N_1800,N_928,N_181);
nor U1801 (N_1801,N_48,N_649);
nand U1802 (N_1802,N_797,N_947);
and U1803 (N_1803,N_110,N_991);
nand U1804 (N_1804,N_23,N_626);
and U1805 (N_1805,N_190,N_411);
nand U1806 (N_1806,N_538,N_145);
xnor U1807 (N_1807,N_400,N_637);
nor U1808 (N_1808,N_322,N_458);
nand U1809 (N_1809,N_587,N_839);
nor U1810 (N_1810,N_552,N_313);
or U1811 (N_1811,N_524,N_471);
nand U1812 (N_1812,N_902,N_228);
nand U1813 (N_1813,N_170,N_289);
and U1814 (N_1814,N_585,N_136);
and U1815 (N_1815,N_395,N_865);
or U1816 (N_1816,N_363,N_11);
nand U1817 (N_1817,N_251,N_521);
xor U1818 (N_1818,N_416,N_936);
or U1819 (N_1819,N_656,N_301);
nand U1820 (N_1820,N_158,N_255);
nor U1821 (N_1821,N_104,N_868);
and U1822 (N_1822,N_745,N_450);
nor U1823 (N_1823,N_741,N_445);
nand U1824 (N_1824,N_314,N_942);
nor U1825 (N_1825,N_74,N_718);
and U1826 (N_1826,N_558,N_496);
xor U1827 (N_1827,N_705,N_645);
and U1828 (N_1828,N_670,N_22);
nor U1829 (N_1829,N_428,N_725);
and U1830 (N_1830,N_577,N_73);
xnor U1831 (N_1831,N_880,N_827);
nor U1832 (N_1832,N_943,N_315);
or U1833 (N_1833,N_135,N_605);
and U1834 (N_1834,N_658,N_294);
and U1835 (N_1835,N_387,N_711);
nand U1836 (N_1836,N_545,N_144);
xor U1837 (N_1837,N_926,N_824);
or U1838 (N_1838,N_48,N_610);
and U1839 (N_1839,N_156,N_958);
nor U1840 (N_1840,N_562,N_442);
nand U1841 (N_1841,N_435,N_613);
or U1842 (N_1842,N_374,N_317);
and U1843 (N_1843,N_24,N_500);
or U1844 (N_1844,N_848,N_25);
xor U1845 (N_1845,N_39,N_153);
and U1846 (N_1846,N_101,N_219);
or U1847 (N_1847,N_684,N_828);
or U1848 (N_1848,N_616,N_359);
xnor U1849 (N_1849,N_79,N_977);
and U1850 (N_1850,N_937,N_712);
and U1851 (N_1851,N_528,N_778);
and U1852 (N_1852,N_399,N_605);
xnor U1853 (N_1853,N_0,N_763);
and U1854 (N_1854,N_70,N_468);
nand U1855 (N_1855,N_345,N_854);
or U1856 (N_1856,N_592,N_525);
or U1857 (N_1857,N_555,N_69);
or U1858 (N_1858,N_833,N_332);
xnor U1859 (N_1859,N_151,N_275);
and U1860 (N_1860,N_911,N_597);
nand U1861 (N_1861,N_360,N_865);
or U1862 (N_1862,N_101,N_461);
nor U1863 (N_1863,N_119,N_298);
nand U1864 (N_1864,N_939,N_34);
nand U1865 (N_1865,N_991,N_977);
xor U1866 (N_1866,N_93,N_355);
and U1867 (N_1867,N_343,N_643);
or U1868 (N_1868,N_40,N_800);
nor U1869 (N_1869,N_841,N_306);
xor U1870 (N_1870,N_973,N_815);
or U1871 (N_1871,N_238,N_280);
nor U1872 (N_1872,N_263,N_15);
or U1873 (N_1873,N_178,N_133);
xnor U1874 (N_1874,N_20,N_783);
and U1875 (N_1875,N_644,N_540);
xor U1876 (N_1876,N_495,N_531);
nand U1877 (N_1877,N_112,N_749);
and U1878 (N_1878,N_197,N_585);
xor U1879 (N_1879,N_15,N_328);
xnor U1880 (N_1880,N_789,N_467);
xnor U1881 (N_1881,N_85,N_852);
or U1882 (N_1882,N_636,N_794);
xor U1883 (N_1883,N_990,N_502);
xor U1884 (N_1884,N_753,N_339);
xor U1885 (N_1885,N_876,N_286);
nor U1886 (N_1886,N_493,N_571);
and U1887 (N_1887,N_165,N_503);
nand U1888 (N_1888,N_136,N_534);
and U1889 (N_1889,N_193,N_889);
nor U1890 (N_1890,N_301,N_22);
or U1891 (N_1891,N_256,N_924);
or U1892 (N_1892,N_793,N_884);
xor U1893 (N_1893,N_282,N_948);
nor U1894 (N_1894,N_649,N_664);
xor U1895 (N_1895,N_943,N_22);
nor U1896 (N_1896,N_950,N_877);
or U1897 (N_1897,N_78,N_498);
nand U1898 (N_1898,N_317,N_152);
xor U1899 (N_1899,N_713,N_7);
nor U1900 (N_1900,N_274,N_561);
and U1901 (N_1901,N_37,N_937);
and U1902 (N_1902,N_682,N_660);
xor U1903 (N_1903,N_211,N_807);
nand U1904 (N_1904,N_499,N_990);
nand U1905 (N_1905,N_81,N_238);
or U1906 (N_1906,N_762,N_12);
nand U1907 (N_1907,N_191,N_465);
nor U1908 (N_1908,N_74,N_734);
nor U1909 (N_1909,N_334,N_215);
nor U1910 (N_1910,N_510,N_209);
or U1911 (N_1911,N_272,N_876);
nand U1912 (N_1912,N_558,N_950);
and U1913 (N_1913,N_785,N_817);
or U1914 (N_1914,N_453,N_376);
nor U1915 (N_1915,N_119,N_422);
or U1916 (N_1916,N_382,N_777);
and U1917 (N_1917,N_14,N_603);
and U1918 (N_1918,N_420,N_403);
xnor U1919 (N_1919,N_943,N_577);
nand U1920 (N_1920,N_255,N_354);
nor U1921 (N_1921,N_413,N_757);
or U1922 (N_1922,N_947,N_971);
nand U1923 (N_1923,N_962,N_976);
and U1924 (N_1924,N_703,N_578);
nand U1925 (N_1925,N_911,N_991);
xnor U1926 (N_1926,N_27,N_670);
nor U1927 (N_1927,N_921,N_8);
and U1928 (N_1928,N_939,N_601);
xnor U1929 (N_1929,N_990,N_626);
and U1930 (N_1930,N_888,N_18);
or U1931 (N_1931,N_455,N_277);
xnor U1932 (N_1932,N_793,N_674);
nand U1933 (N_1933,N_678,N_814);
xnor U1934 (N_1934,N_413,N_599);
xor U1935 (N_1935,N_348,N_766);
and U1936 (N_1936,N_829,N_189);
or U1937 (N_1937,N_648,N_540);
or U1938 (N_1938,N_372,N_240);
nor U1939 (N_1939,N_239,N_43);
and U1940 (N_1940,N_126,N_8);
xor U1941 (N_1941,N_769,N_802);
xnor U1942 (N_1942,N_920,N_580);
or U1943 (N_1943,N_538,N_713);
xor U1944 (N_1944,N_742,N_741);
nor U1945 (N_1945,N_359,N_999);
xor U1946 (N_1946,N_426,N_31);
nor U1947 (N_1947,N_369,N_177);
or U1948 (N_1948,N_764,N_983);
and U1949 (N_1949,N_734,N_482);
nor U1950 (N_1950,N_576,N_369);
nand U1951 (N_1951,N_212,N_882);
nand U1952 (N_1952,N_660,N_523);
xor U1953 (N_1953,N_470,N_620);
xor U1954 (N_1954,N_358,N_436);
nand U1955 (N_1955,N_801,N_604);
xnor U1956 (N_1956,N_47,N_133);
or U1957 (N_1957,N_515,N_911);
nor U1958 (N_1958,N_884,N_736);
xnor U1959 (N_1959,N_385,N_301);
nand U1960 (N_1960,N_206,N_940);
or U1961 (N_1961,N_297,N_246);
nor U1962 (N_1962,N_40,N_773);
nand U1963 (N_1963,N_8,N_322);
nand U1964 (N_1964,N_313,N_558);
xnor U1965 (N_1965,N_4,N_962);
or U1966 (N_1966,N_128,N_171);
nor U1967 (N_1967,N_67,N_206);
or U1968 (N_1968,N_828,N_213);
nand U1969 (N_1969,N_14,N_479);
and U1970 (N_1970,N_622,N_204);
nor U1971 (N_1971,N_602,N_568);
and U1972 (N_1972,N_403,N_556);
xnor U1973 (N_1973,N_893,N_183);
xnor U1974 (N_1974,N_83,N_961);
and U1975 (N_1975,N_420,N_364);
xor U1976 (N_1976,N_677,N_670);
nand U1977 (N_1977,N_161,N_377);
or U1978 (N_1978,N_812,N_673);
and U1979 (N_1979,N_628,N_636);
nor U1980 (N_1980,N_215,N_258);
xor U1981 (N_1981,N_798,N_43);
nor U1982 (N_1982,N_580,N_538);
or U1983 (N_1983,N_452,N_187);
nand U1984 (N_1984,N_598,N_209);
nor U1985 (N_1985,N_70,N_970);
nor U1986 (N_1986,N_125,N_805);
and U1987 (N_1987,N_88,N_715);
nand U1988 (N_1988,N_252,N_390);
or U1989 (N_1989,N_831,N_42);
and U1990 (N_1990,N_601,N_947);
nor U1991 (N_1991,N_824,N_559);
and U1992 (N_1992,N_20,N_877);
or U1993 (N_1993,N_22,N_336);
and U1994 (N_1994,N_299,N_907);
xor U1995 (N_1995,N_60,N_346);
and U1996 (N_1996,N_386,N_895);
nand U1997 (N_1997,N_504,N_240);
or U1998 (N_1998,N_705,N_286);
xnor U1999 (N_1999,N_372,N_274);
xnor U2000 (N_2000,N_1536,N_1555);
nand U2001 (N_2001,N_1092,N_1308);
nor U2002 (N_2002,N_1813,N_1313);
nor U2003 (N_2003,N_1862,N_1278);
and U2004 (N_2004,N_1766,N_1131);
nor U2005 (N_2005,N_1192,N_1783);
xnor U2006 (N_2006,N_1366,N_1093);
or U2007 (N_2007,N_1724,N_1275);
and U2008 (N_2008,N_1334,N_1424);
nand U2009 (N_2009,N_1902,N_1455);
nand U2010 (N_2010,N_1452,N_1500);
nor U2011 (N_2011,N_1437,N_1472);
nor U2012 (N_2012,N_1045,N_1518);
and U2013 (N_2013,N_1411,N_1979);
nand U2014 (N_2014,N_1262,N_1319);
nand U2015 (N_2015,N_1527,N_1935);
or U2016 (N_2016,N_1499,N_1342);
xor U2017 (N_2017,N_1198,N_1463);
and U2018 (N_2018,N_1660,N_1205);
or U2019 (N_2019,N_1774,N_1032);
nor U2020 (N_2020,N_1004,N_1807);
xnor U2021 (N_2021,N_1059,N_1804);
and U2022 (N_2022,N_1776,N_1683);
and U2023 (N_2023,N_1893,N_1709);
xor U2024 (N_2024,N_1841,N_1036);
xnor U2025 (N_2025,N_1641,N_1690);
and U2026 (N_2026,N_1579,N_1016);
or U2027 (N_2027,N_1648,N_1870);
or U2028 (N_2028,N_1451,N_1447);
and U2029 (N_2029,N_1480,N_1118);
or U2030 (N_2030,N_1276,N_1446);
nor U2031 (N_2031,N_1537,N_1915);
nor U2032 (N_2032,N_1869,N_1340);
xor U2033 (N_2033,N_1985,N_1269);
and U2034 (N_2034,N_1458,N_1948);
or U2035 (N_2035,N_1691,N_1227);
xor U2036 (N_2036,N_1558,N_1207);
nand U2037 (N_2037,N_1530,N_1578);
nand U2038 (N_2038,N_1692,N_1063);
nor U2039 (N_2039,N_1675,N_1569);
nor U2040 (N_2040,N_1064,N_1021);
nor U2041 (N_2041,N_1324,N_1875);
xor U2042 (N_2042,N_1298,N_1353);
nand U2043 (N_2043,N_1738,N_1779);
nor U2044 (N_2044,N_1356,N_1442);
and U2045 (N_2045,N_1300,N_1461);
or U2046 (N_2046,N_1323,N_1772);
or U2047 (N_2047,N_1819,N_1614);
nand U2048 (N_2048,N_1068,N_1851);
xor U2049 (N_2049,N_1445,N_1834);
or U2050 (N_2050,N_1554,N_1512);
xnor U2051 (N_2051,N_1787,N_1390);
nor U2052 (N_2052,N_1760,N_1011);
xor U2053 (N_2053,N_1155,N_1229);
nand U2054 (N_2054,N_1401,N_1386);
nand U2055 (N_2055,N_1788,N_1933);
nor U2056 (N_2056,N_1650,N_1913);
or U2057 (N_2057,N_1749,N_1894);
xnor U2058 (N_2058,N_1168,N_1291);
and U2059 (N_2059,N_1793,N_1642);
nand U2060 (N_2060,N_1336,N_1397);
nand U2061 (N_2061,N_1995,N_1343);
and U2062 (N_2062,N_1244,N_1528);
nor U2063 (N_2063,N_1423,N_1140);
and U2064 (N_2064,N_1887,N_1221);
nor U2065 (N_2065,N_1364,N_1532);
nor U2066 (N_2066,N_1634,N_1865);
nand U2067 (N_2067,N_1633,N_1620);
or U2068 (N_2068,N_1975,N_1282);
nor U2069 (N_2069,N_1711,N_1402);
or U2070 (N_2070,N_1674,N_1419);
and U2071 (N_2071,N_1273,N_1846);
nand U2072 (N_2072,N_1061,N_1702);
xor U2073 (N_2073,N_1752,N_1242);
or U2074 (N_2074,N_1185,N_1549);
and U2075 (N_2075,N_1514,N_1584);
and U2076 (N_2076,N_1983,N_1111);
xnor U2077 (N_2077,N_1843,N_1701);
and U2078 (N_2078,N_1687,N_1058);
or U2079 (N_2079,N_1450,N_1984);
and U2080 (N_2080,N_1132,N_1492);
xnor U2081 (N_2081,N_1233,N_1861);
or U2082 (N_2082,N_1707,N_1070);
or U2083 (N_2083,N_1076,N_1713);
xnor U2084 (N_2084,N_1164,N_1930);
and U2085 (N_2085,N_1931,N_1741);
and U2086 (N_2086,N_1226,N_1398);
nand U2087 (N_2087,N_1830,N_1812);
nor U2088 (N_2088,N_1968,N_1252);
nor U2089 (N_2089,N_1287,N_1585);
xnor U2090 (N_2090,N_1355,N_1266);
nor U2091 (N_2091,N_1130,N_1265);
nand U2092 (N_2092,N_1062,N_1407);
nor U2093 (N_2093,N_1860,N_1859);
nand U2094 (N_2094,N_1523,N_1609);
xnor U2095 (N_2095,N_1326,N_1435);
and U2096 (N_2096,N_1958,N_1478);
nand U2097 (N_2097,N_1358,N_1110);
and U2098 (N_2098,N_1534,N_1563);
and U2099 (N_2099,N_1806,N_1494);
xor U2100 (N_2100,N_1717,N_1239);
xor U2101 (N_2101,N_1720,N_1393);
and U2102 (N_2102,N_1337,N_1805);
and U2103 (N_2103,N_1941,N_1715);
xor U2104 (N_2104,N_1588,N_1257);
and U2105 (N_2105,N_1947,N_1377);
or U2106 (N_2106,N_1232,N_1214);
nor U2107 (N_2107,N_1989,N_1224);
xor U2108 (N_2108,N_1255,N_1267);
and U2109 (N_2109,N_1350,N_1874);
nand U2110 (N_2110,N_1414,N_1637);
nand U2111 (N_2111,N_1531,N_1876);
and U2112 (N_2112,N_1270,N_1009);
xnor U2113 (N_2113,N_1256,N_1969);
nor U2114 (N_2114,N_1464,N_1284);
xnor U2115 (N_2115,N_1676,N_1910);
or U2116 (N_2116,N_1504,N_1665);
nor U2117 (N_2117,N_1944,N_1114);
xor U2118 (N_2118,N_1029,N_1627);
and U2119 (N_2119,N_1526,N_1200);
xor U2120 (N_2120,N_1848,N_1574);
nor U2121 (N_2121,N_1980,N_1485);
and U2122 (N_2122,N_1066,N_1891);
xnor U2123 (N_2123,N_1959,N_1926);
xnor U2124 (N_2124,N_1375,N_1961);
xnor U2125 (N_2125,N_1421,N_1509);
and U2126 (N_2126,N_1433,N_1780);
nand U2127 (N_2127,N_1814,N_1801);
nand U2128 (N_2128,N_1657,N_1015);
xor U2129 (N_2129,N_1013,N_1039);
nand U2130 (N_2130,N_1123,N_1428);
xnor U2131 (N_2131,N_1133,N_1965);
nor U2132 (N_2132,N_1576,N_1757);
or U2133 (N_2133,N_1231,N_1880);
and U2134 (N_2134,N_1184,N_1924);
and U2135 (N_2135,N_1671,N_1072);
xor U2136 (N_2136,N_1610,N_1593);
and U2137 (N_2137,N_1723,N_1839);
nor U2138 (N_2138,N_1900,N_1371);
xor U2139 (N_2139,N_1999,N_1234);
xnor U2140 (N_2140,N_1466,N_1177);
nor U2141 (N_2141,N_1595,N_1885);
or U2142 (N_2142,N_1580,N_1301);
nand U2143 (N_2143,N_1213,N_1754);
nand U2144 (N_2144,N_1144,N_1069);
xor U2145 (N_2145,N_1479,N_1543);
xnor U2146 (N_2146,N_1653,N_1084);
or U2147 (N_2147,N_1429,N_1604);
or U2148 (N_2148,N_1142,N_1684);
xor U2149 (N_2149,N_1856,N_1338);
or U2150 (N_2150,N_1467,N_1601);
nor U2151 (N_2151,N_1700,N_1572);
or U2152 (N_2152,N_1113,N_1399);
nand U2153 (N_2153,N_1048,N_1903);
and U2154 (N_2154,N_1764,N_1605);
and U2155 (N_2155,N_1628,N_1249);
and U2156 (N_2156,N_1718,N_1139);
and U2157 (N_2157,N_1762,N_1034);
xnor U2158 (N_2158,N_1348,N_1937);
and U2159 (N_2159,N_1594,N_1483);
nand U2160 (N_2160,N_1341,N_1669);
or U2161 (N_2161,N_1368,N_1607);
nand U2162 (N_2162,N_1420,N_1600);
nand U2163 (N_2163,N_1733,N_1954);
or U2164 (N_2164,N_1208,N_1044);
or U2165 (N_2165,N_1497,N_1219);
or U2166 (N_2166,N_1056,N_1295);
nor U2167 (N_2167,N_1310,N_1272);
nand U2168 (N_2168,N_1074,N_1586);
xnor U2169 (N_2169,N_1680,N_1018);
and U2170 (N_2170,N_1649,N_1264);
nor U2171 (N_2171,N_1163,N_1129);
xnor U2172 (N_2172,N_1564,N_1740);
nor U2173 (N_2173,N_1247,N_1087);
and U2174 (N_2174,N_1977,N_1904);
nor U2175 (N_2175,N_1292,N_1288);
and U2176 (N_2176,N_1135,N_1925);
nand U2177 (N_2177,N_1112,N_1384);
nor U2178 (N_2178,N_1837,N_1573);
nor U2179 (N_2179,N_1559,N_1784);
and U2180 (N_2180,N_1756,N_1519);
xor U2181 (N_2181,N_1745,N_1613);
nand U2182 (N_2182,N_1457,N_1729);
nand U2183 (N_2183,N_1259,N_1491);
nand U2184 (N_2184,N_1615,N_1847);
nor U2185 (N_2185,N_1071,N_1042);
nand U2186 (N_2186,N_1545,N_1951);
and U2187 (N_2187,N_1612,N_1410);
nand U2188 (N_2188,N_1845,N_1566);
nand U2189 (N_2189,N_1544,N_1522);
and U2190 (N_2190,N_1912,N_1117);
nor U2191 (N_2191,N_1597,N_1722);
xor U2192 (N_2192,N_1666,N_1978);
nor U2193 (N_2193,N_1879,N_1309);
nor U2194 (N_2194,N_1529,N_1746);
nor U2195 (N_2195,N_1629,N_1141);
nand U2196 (N_2196,N_1484,N_1197);
nand U2197 (N_2197,N_1031,N_1206);
xor U2198 (N_2198,N_1202,N_1037);
nand U2199 (N_2199,N_1817,N_1525);
and U2200 (N_2200,N_1728,N_1007);
or U2201 (N_2201,N_1169,N_1006);
nor U2202 (N_2202,N_1081,N_1165);
nor U2203 (N_2203,N_1489,N_1695);
nor U2204 (N_2204,N_1183,N_1898);
xnor U2205 (N_2205,N_1515,N_1901);
nand U2206 (N_2206,N_1149,N_1770);
nor U2207 (N_2207,N_1750,N_1907);
nor U2208 (N_2208,N_1465,N_1000);
nand U2209 (N_2209,N_1473,N_1359);
or U2210 (N_2210,N_1955,N_1581);
xnor U2211 (N_2211,N_1427,N_1236);
xnor U2212 (N_2212,N_1686,N_1619);
or U2213 (N_2213,N_1743,N_1626);
nor U2214 (N_2214,N_1381,N_1872);
or U2215 (N_2215,N_1100,N_1710);
nand U2216 (N_2216,N_1172,N_1993);
or U2217 (N_2217,N_1120,N_1547);
nand U2218 (N_2218,N_1339,N_1507);
nor U2219 (N_2219,N_1280,N_1922);
nand U2220 (N_2220,N_1990,N_1406);
nand U2221 (N_2221,N_1694,N_1550);
nand U2222 (N_2222,N_1453,N_1173);
and U2223 (N_2223,N_1744,N_1181);
nand U2224 (N_2224,N_1047,N_1060);
and U2225 (N_2225,N_1726,N_1436);
and U2226 (N_2226,N_1542,N_1328);
or U2227 (N_2227,N_1538,N_1682);
or U2228 (N_2228,N_1625,N_1932);
and U2229 (N_2229,N_1121,N_1739);
or U2230 (N_2230,N_1617,N_1430);
or U2231 (N_2231,N_1160,N_1082);
nand U2232 (N_2232,N_1195,N_1191);
nand U2233 (N_2233,N_1373,N_1331);
or U2234 (N_2234,N_1546,N_1260);
xor U2235 (N_2235,N_1152,N_1828);
and U2236 (N_2236,N_1151,N_1474);
and U2237 (N_2237,N_1444,N_1689);
or U2238 (N_2238,N_1618,N_1513);
xnor U2239 (N_2239,N_1575,N_1622);
or U2240 (N_2240,N_1592,N_1055);
or U2241 (N_2241,N_1871,N_1327);
nand U2242 (N_2242,N_1281,N_1970);
and U2243 (N_2243,N_1175,N_1418);
or U2244 (N_2244,N_1046,N_1187);
nand U2245 (N_2245,N_1090,N_1973);
and U2246 (N_2246,N_1128,N_1345);
xor U2247 (N_2247,N_1655,N_1696);
and U2248 (N_2248,N_1391,N_1963);
nor U2249 (N_2249,N_1939,N_1976);
or U2250 (N_2250,N_1404,N_1106);
and U2251 (N_2251,N_1699,N_1318);
nand U2252 (N_2252,N_1456,N_1038);
nand U2253 (N_2253,N_1277,N_1667);
xnor U2254 (N_2254,N_1568,N_1241);
nor U2255 (N_2255,N_1996,N_1520);
nor U2256 (N_2256,N_1054,N_1982);
and U2257 (N_2257,N_1664,N_1225);
and U2258 (N_2258,N_1946,N_1878);
xnor U2259 (N_2259,N_1119,N_1864);
nand U2260 (N_2260,N_1840,N_1816);
and U2261 (N_2261,N_1178,N_1646);
xor U2262 (N_2262,N_1636,N_1987);
and U2263 (N_2263,N_1844,N_1335);
and U2264 (N_2264,N_1268,N_1639);
nand U2265 (N_2265,N_1086,N_1681);
or U2266 (N_2266,N_1981,N_1734);
or U2267 (N_2267,N_1432,N_1583);
nand U2268 (N_2268,N_1223,N_1422);
nor U2269 (N_2269,N_1166,N_1498);
xor U2270 (N_2270,N_1833,N_1917);
or U2271 (N_2271,N_1104,N_1796);
nand U2272 (N_2272,N_1263,N_1017);
nand U2273 (N_2273,N_1590,N_1412);
and U2274 (N_2274,N_1789,N_1890);
and U2275 (N_2275,N_1477,N_1797);
xor U2276 (N_2276,N_1591,N_1376);
nand U2277 (N_2277,N_1773,N_1621);
nand U2278 (N_2278,N_1174,N_1556);
nand U2279 (N_2279,N_1330,N_1886);
or U2280 (N_2280,N_1911,N_1493);
nor U2281 (N_2281,N_1005,N_1798);
xnor U2282 (N_2282,N_1125,N_1988);
xnor U2283 (N_2283,N_1956,N_1321);
and U2284 (N_2284,N_1877,N_1928);
and U2285 (N_2285,N_1103,N_1873);
nand U2286 (N_2286,N_1361,N_1810);
and U2287 (N_2287,N_1352,N_1517);
nand U2288 (N_2288,N_1799,N_1020);
nand U2289 (N_2289,N_1882,N_1194);
xor U2290 (N_2290,N_1261,N_1153);
or U2291 (N_2291,N_1967,N_1842);
or U2292 (N_2292,N_1363,N_1829);
and U2293 (N_2293,N_1325,N_1438);
and U2294 (N_2294,N_1154,N_1077);
nand U2295 (N_2295,N_1240,N_1656);
nand U2296 (N_2296,N_1822,N_1099);
nor U2297 (N_2297,N_1663,N_1654);
nor U2298 (N_2298,N_1630,N_1116);
nor U2299 (N_2299,N_1314,N_1540);
xor U2300 (N_2300,N_1631,N_1026);
nor U2301 (N_2301,N_1571,N_1551);
or U2302 (N_2302,N_1199,N_1274);
or U2303 (N_2303,N_1302,N_1245);
and U2304 (N_2304,N_1992,N_1818);
xor U2305 (N_2305,N_1897,N_1957);
nand U2306 (N_2306,N_1449,N_1821);
nand U2307 (N_2307,N_1248,N_1258);
nand U2308 (N_2308,N_1162,N_1075);
xor U2309 (N_2309,N_1067,N_1329);
or U2310 (N_2310,N_1644,N_1736);
nand U2311 (N_2311,N_1714,N_1124);
and U2312 (N_2312,N_1632,N_1672);
or U2313 (N_2313,N_1027,N_1201);
nand U2314 (N_2314,N_1790,N_1719);
nand U2315 (N_2315,N_1785,N_1468);
and U2316 (N_2316,N_1170,N_1052);
xor U2317 (N_2317,N_1541,N_1596);
and U2318 (N_2318,N_1997,N_1367);
and U2319 (N_2319,N_1297,N_1721);
nor U2320 (N_2320,N_1293,N_1161);
nor U2321 (N_2321,N_1475,N_1439);
or U2322 (N_2322,N_1105,N_1156);
nand U2323 (N_2323,N_1725,N_1881);
or U2324 (N_2324,N_1986,N_1394);
or U2325 (N_2325,N_1598,N_1028);
nor U2326 (N_2326,N_1508,N_1608);
xnor U2327 (N_2327,N_1511,N_1868);
and U2328 (N_2328,N_1496,N_1703);
nand U2329 (N_2329,N_1565,N_1415);
and U2330 (N_2330,N_1688,N_1697);
nand U2331 (N_2331,N_1552,N_1661);
and U2332 (N_2332,N_1487,N_1974);
nor U2333 (N_2333,N_1835,N_1008);
and U2334 (N_2334,N_1285,N_1126);
nand U2335 (N_2335,N_1251,N_1101);
or U2336 (N_2336,N_1747,N_1849);
xor U2337 (N_2337,N_1408,N_1417);
xor U2338 (N_2338,N_1771,N_1148);
nor U2339 (N_2339,N_1186,N_1403);
xor U2340 (N_2340,N_1949,N_1127);
and U2341 (N_2341,N_1501,N_1346);
or U2342 (N_2342,N_1022,N_1651);
nand U2343 (N_2343,N_1378,N_1182);
nor U2344 (N_2344,N_1150,N_1434);
nand U2345 (N_2345,N_1296,N_1180);
nand U2346 (N_2346,N_1677,N_1372);
xor U2347 (N_2347,N_1994,N_1279);
nor U2348 (N_2348,N_1137,N_1866);
or U2349 (N_2349,N_1317,N_1243);
and U2350 (N_2350,N_1362,N_1204);
and U2351 (N_2351,N_1742,N_1158);
or U2352 (N_2352,N_1624,N_1089);
xnor U2353 (N_2353,N_1827,N_1290);
xor U2354 (N_2354,N_1892,N_1557);
xnor U2355 (N_2355,N_1919,N_1838);
and U2356 (N_2356,N_1409,N_1025);
and U2357 (N_2357,N_1109,N_1815);
xor U2358 (N_2358,N_1775,N_1091);
nor U2359 (N_2359,N_1896,N_1502);
or U2360 (N_2360,N_1767,N_1950);
nor U2361 (N_2361,N_1673,N_1476);
nor U2362 (N_2362,N_1030,N_1735);
xnor U2363 (N_2363,N_1670,N_1769);
nand U2364 (N_2364,N_1803,N_1395);
nor U2365 (N_2365,N_1041,N_1826);
nor U2366 (N_2366,N_1645,N_1303);
nor U2367 (N_2367,N_1108,N_1332);
nor U2368 (N_2368,N_1920,N_1899);
nand U2369 (N_2369,N_1010,N_1238);
xnor U2370 (N_2370,N_1972,N_1603);
or U2371 (N_2371,N_1057,N_1209);
and U2372 (N_2372,N_1960,N_1146);
xnor U2373 (N_2373,N_1587,N_1889);
xnor U2374 (N_2374,N_1716,N_1962);
nor U2375 (N_2375,N_1053,N_1831);
nand U2376 (N_2376,N_1351,N_1431);
nor U2377 (N_2377,N_1385,N_1383);
or U2378 (N_2378,N_1003,N_1212);
xor U2379 (N_2379,N_1964,N_1049);
xor U2380 (N_2380,N_1481,N_1811);
and U2381 (N_2381,N_1758,N_1905);
xor U2382 (N_2382,N_1380,N_1854);
nor U2383 (N_2383,N_1616,N_1379);
and U2384 (N_2384,N_1294,N_1416);
or U2385 (N_2385,N_1782,N_1867);
nand U2386 (N_2386,N_1506,N_1283);
and U2387 (N_2387,N_1441,N_1107);
or U2388 (N_2388,N_1159,N_1211);
xnor U2389 (N_2389,N_1708,N_1940);
and U2390 (N_2390,N_1753,N_1495);
or U2391 (N_2391,N_1759,N_1535);
nor U2392 (N_2392,N_1102,N_1024);
nor U2393 (N_2393,N_1157,N_1188);
xnor U2394 (N_2394,N_1704,N_1357);
and U2395 (N_2395,N_1638,N_1971);
xnor U2396 (N_2396,N_1705,N_1658);
nand U2397 (N_2397,N_1085,N_1635);
and U2398 (N_2398,N_1454,N_1577);
and U2399 (N_2399,N_1369,N_1289);
and U2400 (N_2400,N_1425,N_1599);
or U2401 (N_2401,N_1088,N_1800);
xor U2402 (N_2402,N_1909,N_1659);
and U2403 (N_2403,N_1203,N_1755);
or U2404 (N_2404,N_1895,N_1299);
xnor U2405 (N_2405,N_1490,N_1035);
xor U2406 (N_2406,N_1765,N_1448);
xnor U2407 (N_2407,N_1923,N_1179);
and U2408 (N_2408,N_1322,N_1823);
xnor U2409 (N_2409,N_1073,N_1623);
xor U2410 (N_2410,N_1304,N_1908);
and U2411 (N_2411,N_1777,N_1888);
and U2412 (N_2412,N_1853,N_1136);
xnor U2413 (N_2413,N_1080,N_1218);
xor U2414 (N_2414,N_1078,N_1065);
and U2415 (N_2415,N_1014,N_1778);
or U2416 (N_2416,N_1143,N_1712);
nand U2417 (N_2417,N_1333,N_1921);
and U2418 (N_2418,N_1471,N_1392);
nand U2419 (N_2419,N_1706,N_1370);
xnor U2420 (N_2420,N_1365,N_1469);
xor U2421 (N_2421,N_1190,N_1043);
and U2422 (N_2422,N_1679,N_1095);
nand U2423 (N_2423,N_1459,N_1316);
nor U2424 (N_2424,N_1918,N_1751);
nand U2425 (N_2425,N_1791,N_1562);
nand U2426 (N_2426,N_1040,N_1389);
and U2427 (N_2427,N_1311,N_1561);
or U2428 (N_2428,N_1832,N_1320);
xor U2429 (N_2429,N_1503,N_1210);
and U2430 (N_2430,N_1852,N_1914);
and U2431 (N_2431,N_1001,N_1235);
xor U2432 (N_2432,N_1567,N_1548);
and U2433 (N_2433,N_1938,N_1820);
and U2434 (N_2434,N_1470,N_1460);
nor U2435 (N_2435,N_1050,N_1482);
xor U2436 (N_2436,N_1945,N_1929);
nand U2437 (N_2437,N_1189,N_1727);
nand U2438 (N_2438,N_1138,N_1647);
xor U2439 (N_2439,N_1222,N_1606);
xor U2440 (N_2440,N_1906,N_1934);
and U2441 (N_2441,N_1462,N_1134);
nand U2442 (N_2442,N_1307,N_1079);
or U2443 (N_2443,N_1413,N_1443);
xor U2444 (N_2444,N_1405,N_1196);
nor U2445 (N_2445,N_1668,N_1560);
nand U2446 (N_2446,N_1230,N_1685);
nor U2447 (N_2447,N_1786,N_1884);
and U2448 (N_2448,N_1737,N_1510);
nor U2449 (N_2449,N_1652,N_1486);
and U2450 (N_2450,N_1312,N_1936);
xnor U2451 (N_2451,N_1347,N_1516);
nand U2452 (N_2452,N_1349,N_1344);
nand U2453 (N_2453,N_1122,N_1193);
nand U2454 (N_2454,N_1374,N_1693);
nand U2455 (N_2455,N_1228,N_1858);
xnor U2456 (N_2456,N_1387,N_1570);
or U2457 (N_2457,N_1794,N_1602);
nor U2458 (N_2458,N_1857,N_1927);
xnor U2459 (N_2459,N_1253,N_1115);
and U2460 (N_2460,N_1216,N_1094);
or U2461 (N_2461,N_1589,N_1640);
or U2462 (N_2462,N_1098,N_1698);
nor U2463 (N_2463,N_1254,N_1855);
and U2464 (N_2464,N_1792,N_1539);
nand U2465 (N_2465,N_1083,N_1802);
or U2466 (N_2466,N_1217,N_1662);
nand U2467 (N_2467,N_1748,N_1315);
and U2468 (N_2468,N_1271,N_1916);
nand U2469 (N_2469,N_1145,N_1824);
xor U2470 (N_2470,N_1643,N_1360);
or U2471 (N_2471,N_1220,N_1306);
xor U2472 (N_2472,N_1382,N_1250);
and U2473 (N_2473,N_1533,N_1002);
xor U2474 (N_2474,N_1850,N_1400);
nand U2475 (N_2475,N_1763,N_1582);
and U2476 (N_2476,N_1553,N_1440);
nor U2477 (N_2477,N_1998,N_1731);
nand U2478 (N_2478,N_1761,N_1426);
or U2479 (N_2479,N_1396,N_1863);
xor U2480 (N_2480,N_1883,N_1809);
and U2481 (N_2481,N_1521,N_1781);
and U2482 (N_2482,N_1952,N_1678);
xor U2483 (N_2483,N_1611,N_1942);
xor U2484 (N_2484,N_1167,N_1051);
xor U2485 (N_2485,N_1730,N_1953);
and U2486 (N_2486,N_1354,N_1147);
or U2487 (N_2487,N_1305,N_1023);
xor U2488 (N_2488,N_1215,N_1808);
or U2489 (N_2489,N_1825,N_1732);
and U2490 (N_2490,N_1019,N_1286);
nand U2491 (N_2491,N_1795,N_1768);
nor U2492 (N_2492,N_1388,N_1096);
xor U2493 (N_2493,N_1991,N_1836);
nor U2494 (N_2494,N_1966,N_1012);
nand U2495 (N_2495,N_1246,N_1488);
nor U2496 (N_2496,N_1505,N_1171);
nor U2497 (N_2497,N_1176,N_1097);
and U2498 (N_2498,N_1033,N_1943);
nor U2499 (N_2499,N_1524,N_1237);
nand U2500 (N_2500,N_1105,N_1279);
xor U2501 (N_2501,N_1704,N_1555);
nor U2502 (N_2502,N_1343,N_1415);
xor U2503 (N_2503,N_1143,N_1402);
or U2504 (N_2504,N_1128,N_1301);
nor U2505 (N_2505,N_1948,N_1409);
nand U2506 (N_2506,N_1665,N_1271);
and U2507 (N_2507,N_1185,N_1003);
nand U2508 (N_2508,N_1206,N_1377);
and U2509 (N_2509,N_1899,N_1034);
and U2510 (N_2510,N_1932,N_1804);
xnor U2511 (N_2511,N_1639,N_1890);
nand U2512 (N_2512,N_1671,N_1704);
xor U2513 (N_2513,N_1466,N_1549);
and U2514 (N_2514,N_1217,N_1873);
or U2515 (N_2515,N_1222,N_1130);
xor U2516 (N_2516,N_1077,N_1752);
and U2517 (N_2517,N_1052,N_1930);
nand U2518 (N_2518,N_1903,N_1462);
nand U2519 (N_2519,N_1478,N_1247);
xnor U2520 (N_2520,N_1115,N_1029);
nand U2521 (N_2521,N_1969,N_1533);
or U2522 (N_2522,N_1714,N_1253);
and U2523 (N_2523,N_1445,N_1713);
nand U2524 (N_2524,N_1076,N_1510);
nor U2525 (N_2525,N_1917,N_1260);
or U2526 (N_2526,N_1213,N_1666);
and U2527 (N_2527,N_1554,N_1396);
nor U2528 (N_2528,N_1231,N_1912);
and U2529 (N_2529,N_1849,N_1960);
nand U2530 (N_2530,N_1310,N_1164);
nand U2531 (N_2531,N_1958,N_1985);
and U2532 (N_2532,N_1303,N_1870);
nand U2533 (N_2533,N_1993,N_1474);
nor U2534 (N_2534,N_1134,N_1049);
nand U2535 (N_2535,N_1630,N_1130);
xnor U2536 (N_2536,N_1475,N_1363);
or U2537 (N_2537,N_1088,N_1219);
nand U2538 (N_2538,N_1988,N_1622);
nor U2539 (N_2539,N_1821,N_1085);
xor U2540 (N_2540,N_1895,N_1006);
xnor U2541 (N_2541,N_1536,N_1511);
and U2542 (N_2542,N_1716,N_1722);
xor U2543 (N_2543,N_1682,N_1186);
nand U2544 (N_2544,N_1764,N_1530);
nor U2545 (N_2545,N_1904,N_1729);
xor U2546 (N_2546,N_1734,N_1926);
or U2547 (N_2547,N_1377,N_1784);
and U2548 (N_2548,N_1306,N_1677);
xor U2549 (N_2549,N_1651,N_1492);
and U2550 (N_2550,N_1150,N_1753);
nor U2551 (N_2551,N_1404,N_1008);
or U2552 (N_2552,N_1479,N_1850);
xnor U2553 (N_2553,N_1966,N_1363);
nor U2554 (N_2554,N_1157,N_1990);
nand U2555 (N_2555,N_1403,N_1231);
nand U2556 (N_2556,N_1855,N_1657);
xor U2557 (N_2557,N_1660,N_1566);
or U2558 (N_2558,N_1009,N_1980);
nand U2559 (N_2559,N_1574,N_1222);
nor U2560 (N_2560,N_1364,N_1675);
nor U2561 (N_2561,N_1634,N_1597);
and U2562 (N_2562,N_1778,N_1105);
or U2563 (N_2563,N_1440,N_1313);
nor U2564 (N_2564,N_1263,N_1923);
xor U2565 (N_2565,N_1269,N_1161);
or U2566 (N_2566,N_1646,N_1045);
and U2567 (N_2567,N_1823,N_1802);
nand U2568 (N_2568,N_1128,N_1474);
nor U2569 (N_2569,N_1045,N_1318);
and U2570 (N_2570,N_1777,N_1365);
xor U2571 (N_2571,N_1032,N_1520);
nor U2572 (N_2572,N_1267,N_1032);
xnor U2573 (N_2573,N_1913,N_1718);
and U2574 (N_2574,N_1050,N_1750);
and U2575 (N_2575,N_1984,N_1488);
or U2576 (N_2576,N_1855,N_1335);
nand U2577 (N_2577,N_1478,N_1885);
xnor U2578 (N_2578,N_1077,N_1888);
nor U2579 (N_2579,N_1268,N_1929);
nor U2580 (N_2580,N_1183,N_1615);
nor U2581 (N_2581,N_1549,N_1966);
nand U2582 (N_2582,N_1968,N_1425);
or U2583 (N_2583,N_1783,N_1925);
nor U2584 (N_2584,N_1671,N_1550);
xor U2585 (N_2585,N_1962,N_1543);
nor U2586 (N_2586,N_1641,N_1663);
xor U2587 (N_2587,N_1730,N_1769);
nand U2588 (N_2588,N_1672,N_1664);
or U2589 (N_2589,N_1106,N_1204);
nor U2590 (N_2590,N_1181,N_1581);
nand U2591 (N_2591,N_1266,N_1698);
nand U2592 (N_2592,N_1136,N_1846);
xnor U2593 (N_2593,N_1121,N_1520);
xor U2594 (N_2594,N_1800,N_1638);
nor U2595 (N_2595,N_1013,N_1584);
nand U2596 (N_2596,N_1324,N_1857);
or U2597 (N_2597,N_1013,N_1050);
and U2598 (N_2598,N_1199,N_1443);
or U2599 (N_2599,N_1062,N_1479);
xor U2600 (N_2600,N_1975,N_1952);
or U2601 (N_2601,N_1060,N_1660);
nand U2602 (N_2602,N_1423,N_1494);
nand U2603 (N_2603,N_1263,N_1473);
nor U2604 (N_2604,N_1696,N_1327);
and U2605 (N_2605,N_1660,N_1292);
nor U2606 (N_2606,N_1828,N_1437);
nand U2607 (N_2607,N_1044,N_1684);
nor U2608 (N_2608,N_1144,N_1498);
xor U2609 (N_2609,N_1022,N_1115);
nor U2610 (N_2610,N_1024,N_1207);
or U2611 (N_2611,N_1373,N_1388);
and U2612 (N_2612,N_1762,N_1129);
xnor U2613 (N_2613,N_1084,N_1679);
nand U2614 (N_2614,N_1492,N_1334);
nand U2615 (N_2615,N_1964,N_1037);
or U2616 (N_2616,N_1401,N_1389);
and U2617 (N_2617,N_1732,N_1826);
and U2618 (N_2618,N_1459,N_1494);
nand U2619 (N_2619,N_1990,N_1343);
or U2620 (N_2620,N_1084,N_1237);
and U2621 (N_2621,N_1526,N_1350);
xnor U2622 (N_2622,N_1876,N_1297);
nor U2623 (N_2623,N_1447,N_1676);
and U2624 (N_2624,N_1001,N_1226);
and U2625 (N_2625,N_1829,N_1126);
or U2626 (N_2626,N_1342,N_1346);
xnor U2627 (N_2627,N_1566,N_1239);
and U2628 (N_2628,N_1692,N_1358);
or U2629 (N_2629,N_1315,N_1282);
or U2630 (N_2630,N_1526,N_1730);
xor U2631 (N_2631,N_1436,N_1801);
and U2632 (N_2632,N_1143,N_1283);
and U2633 (N_2633,N_1315,N_1514);
nand U2634 (N_2634,N_1614,N_1731);
nand U2635 (N_2635,N_1457,N_1847);
xnor U2636 (N_2636,N_1418,N_1871);
nor U2637 (N_2637,N_1501,N_1224);
nor U2638 (N_2638,N_1562,N_1590);
nor U2639 (N_2639,N_1395,N_1431);
or U2640 (N_2640,N_1872,N_1710);
xnor U2641 (N_2641,N_1975,N_1030);
nor U2642 (N_2642,N_1446,N_1547);
nand U2643 (N_2643,N_1241,N_1251);
or U2644 (N_2644,N_1520,N_1971);
nor U2645 (N_2645,N_1667,N_1998);
nor U2646 (N_2646,N_1892,N_1334);
nand U2647 (N_2647,N_1079,N_1231);
or U2648 (N_2648,N_1826,N_1903);
or U2649 (N_2649,N_1955,N_1720);
or U2650 (N_2650,N_1933,N_1054);
xor U2651 (N_2651,N_1717,N_1952);
and U2652 (N_2652,N_1250,N_1254);
nor U2653 (N_2653,N_1367,N_1547);
xor U2654 (N_2654,N_1392,N_1667);
and U2655 (N_2655,N_1466,N_1181);
and U2656 (N_2656,N_1305,N_1258);
nand U2657 (N_2657,N_1126,N_1756);
and U2658 (N_2658,N_1024,N_1614);
xnor U2659 (N_2659,N_1577,N_1540);
nand U2660 (N_2660,N_1667,N_1794);
or U2661 (N_2661,N_1635,N_1178);
xor U2662 (N_2662,N_1677,N_1300);
nor U2663 (N_2663,N_1530,N_1882);
and U2664 (N_2664,N_1692,N_1288);
nand U2665 (N_2665,N_1346,N_1901);
or U2666 (N_2666,N_1296,N_1713);
xor U2667 (N_2667,N_1304,N_1923);
xor U2668 (N_2668,N_1756,N_1842);
nor U2669 (N_2669,N_1180,N_1016);
xor U2670 (N_2670,N_1390,N_1096);
and U2671 (N_2671,N_1919,N_1896);
xor U2672 (N_2672,N_1811,N_1376);
xor U2673 (N_2673,N_1205,N_1134);
or U2674 (N_2674,N_1573,N_1097);
or U2675 (N_2675,N_1517,N_1572);
or U2676 (N_2676,N_1912,N_1695);
xor U2677 (N_2677,N_1136,N_1726);
xor U2678 (N_2678,N_1909,N_1785);
xnor U2679 (N_2679,N_1884,N_1937);
or U2680 (N_2680,N_1610,N_1851);
nand U2681 (N_2681,N_1748,N_1827);
nor U2682 (N_2682,N_1884,N_1137);
nor U2683 (N_2683,N_1875,N_1676);
and U2684 (N_2684,N_1382,N_1109);
xnor U2685 (N_2685,N_1982,N_1970);
nand U2686 (N_2686,N_1343,N_1204);
and U2687 (N_2687,N_1691,N_1548);
and U2688 (N_2688,N_1056,N_1687);
and U2689 (N_2689,N_1905,N_1706);
nand U2690 (N_2690,N_1011,N_1424);
nand U2691 (N_2691,N_1833,N_1310);
nor U2692 (N_2692,N_1978,N_1833);
xor U2693 (N_2693,N_1758,N_1995);
xor U2694 (N_2694,N_1747,N_1613);
or U2695 (N_2695,N_1352,N_1046);
and U2696 (N_2696,N_1953,N_1003);
xnor U2697 (N_2697,N_1602,N_1042);
xnor U2698 (N_2698,N_1438,N_1265);
nor U2699 (N_2699,N_1557,N_1526);
xor U2700 (N_2700,N_1074,N_1582);
and U2701 (N_2701,N_1438,N_1244);
and U2702 (N_2702,N_1515,N_1918);
and U2703 (N_2703,N_1958,N_1753);
and U2704 (N_2704,N_1821,N_1795);
nor U2705 (N_2705,N_1151,N_1449);
xnor U2706 (N_2706,N_1929,N_1844);
or U2707 (N_2707,N_1807,N_1731);
or U2708 (N_2708,N_1739,N_1217);
nand U2709 (N_2709,N_1513,N_1063);
xnor U2710 (N_2710,N_1101,N_1558);
nor U2711 (N_2711,N_1752,N_1663);
nor U2712 (N_2712,N_1739,N_1170);
and U2713 (N_2713,N_1065,N_1785);
nand U2714 (N_2714,N_1957,N_1222);
and U2715 (N_2715,N_1062,N_1822);
and U2716 (N_2716,N_1713,N_1819);
and U2717 (N_2717,N_1592,N_1206);
nand U2718 (N_2718,N_1540,N_1213);
and U2719 (N_2719,N_1189,N_1933);
nand U2720 (N_2720,N_1562,N_1928);
nor U2721 (N_2721,N_1447,N_1891);
and U2722 (N_2722,N_1500,N_1676);
or U2723 (N_2723,N_1318,N_1325);
nand U2724 (N_2724,N_1508,N_1958);
xor U2725 (N_2725,N_1730,N_1268);
nor U2726 (N_2726,N_1348,N_1072);
or U2727 (N_2727,N_1371,N_1120);
and U2728 (N_2728,N_1873,N_1087);
or U2729 (N_2729,N_1922,N_1526);
nor U2730 (N_2730,N_1658,N_1223);
or U2731 (N_2731,N_1851,N_1246);
xor U2732 (N_2732,N_1082,N_1440);
xnor U2733 (N_2733,N_1953,N_1666);
or U2734 (N_2734,N_1895,N_1937);
and U2735 (N_2735,N_1334,N_1073);
nor U2736 (N_2736,N_1008,N_1238);
and U2737 (N_2737,N_1449,N_1228);
or U2738 (N_2738,N_1777,N_1940);
nand U2739 (N_2739,N_1248,N_1781);
or U2740 (N_2740,N_1769,N_1760);
nor U2741 (N_2741,N_1725,N_1029);
or U2742 (N_2742,N_1207,N_1532);
or U2743 (N_2743,N_1185,N_1027);
or U2744 (N_2744,N_1887,N_1550);
nor U2745 (N_2745,N_1929,N_1018);
or U2746 (N_2746,N_1697,N_1722);
xnor U2747 (N_2747,N_1141,N_1577);
xnor U2748 (N_2748,N_1682,N_1743);
nor U2749 (N_2749,N_1046,N_1614);
nor U2750 (N_2750,N_1777,N_1057);
xnor U2751 (N_2751,N_1176,N_1414);
or U2752 (N_2752,N_1452,N_1928);
nor U2753 (N_2753,N_1569,N_1951);
nor U2754 (N_2754,N_1540,N_1734);
nand U2755 (N_2755,N_1435,N_1181);
and U2756 (N_2756,N_1874,N_1630);
or U2757 (N_2757,N_1534,N_1939);
xnor U2758 (N_2758,N_1696,N_1954);
and U2759 (N_2759,N_1240,N_1040);
nor U2760 (N_2760,N_1931,N_1164);
and U2761 (N_2761,N_1644,N_1740);
nand U2762 (N_2762,N_1442,N_1529);
nand U2763 (N_2763,N_1797,N_1642);
or U2764 (N_2764,N_1996,N_1245);
or U2765 (N_2765,N_1303,N_1147);
nand U2766 (N_2766,N_1660,N_1049);
nor U2767 (N_2767,N_1605,N_1881);
nand U2768 (N_2768,N_1260,N_1831);
and U2769 (N_2769,N_1407,N_1155);
and U2770 (N_2770,N_1269,N_1437);
and U2771 (N_2771,N_1339,N_1937);
nor U2772 (N_2772,N_1475,N_1669);
and U2773 (N_2773,N_1304,N_1901);
or U2774 (N_2774,N_1451,N_1935);
or U2775 (N_2775,N_1137,N_1094);
xor U2776 (N_2776,N_1871,N_1561);
or U2777 (N_2777,N_1269,N_1511);
nor U2778 (N_2778,N_1779,N_1844);
or U2779 (N_2779,N_1300,N_1574);
or U2780 (N_2780,N_1122,N_1640);
nand U2781 (N_2781,N_1059,N_1307);
nor U2782 (N_2782,N_1530,N_1338);
nand U2783 (N_2783,N_1666,N_1699);
xnor U2784 (N_2784,N_1238,N_1556);
nor U2785 (N_2785,N_1323,N_1241);
nand U2786 (N_2786,N_1513,N_1581);
xor U2787 (N_2787,N_1148,N_1490);
nor U2788 (N_2788,N_1215,N_1592);
xor U2789 (N_2789,N_1251,N_1366);
and U2790 (N_2790,N_1374,N_1892);
nor U2791 (N_2791,N_1645,N_1668);
nor U2792 (N_2792,N_1788,N_1685);
nor U2793 (N_2793,N_1524,N_1730);
and U2794 (N_2794,N_1835,N_1528);
nor U2795 (N_2795,N_1712,N_1031);
nand U2796 (N_2796,N_1635,N_1782);
and U2797 (N_2797,N_1225,N_1609);
nor U2798 (N_2798,N_1048,N_1550);
nor U2799 (N_2799,N_1515,N_1759);
nand U2800 (N_2800,N_1040,N_1769);
nor U2801 (N_2801,N_1302,N_1385);
nand U2802 (N_2802,N_1732,N_1338);
and U2803 (N_2803,N_1667,N_1896);
or U2804 (N_2804,N_1258,N_1013);
nor U2805 (N_2805,N_1186,N_1049);
and U2806 (N_2806,N_1489,N_1696);
or U2807 (N_2807,N_1000,N_1280);
or U2808 (N_2808,N_1240,N_1235);
xor U2809 (N_2809,N_1257,N_1126);
xnor U2810 (N_2810,N_1702,N_1263);
nor U2811 (N_2811,N_1231,N_1726);
nand U2812 (N_2812,N_1907,N_1811);
nand U2813 (N_2813,N_1173,N_1497);
or U2814 (N_2814,N_1677,N_1844);
nor U2815 (N_2815,N_1702,N_1660);
and U2816 (N_2816,N_1274,N_1493);
xor U2817 (N_2817,N_1434,N_1818);
nand U2818 (N_2818,N_1015,N_1993);
nand U2819 (N_2819,N_1237,N_1850);
and U2820 (N_2820,N_1331,N_1386);
xor U2821 (N_2821,N_1972,N_1052);
nand U2822 (N_2822,N_1432,N_1974);
nor U2823 (N_2823,N_1727,N_1260);
and U2824 (N_2824,N_1801,N_1225);
and U2825 (N_2825,N_1420,N_1766);
or U2826 (N_2826,N_1944,N_1369);
and U2827 (N_2827,N_1284,N_1967);
or U2828 (N_2828,N_1240,N_1060);
xnor U2829 (N_2829,N_1140,N_1279);
nor U2830 (N_2830,N_1456,N_1290);
nand U2831 (N_2831,N_1201,N_1490);
and U2832 (N_2832,N_1047,N_1039);
or U2833 (N_2833,N_1021,N_1380);
and U2834 (N_2834,N_1649,N_1320);
nor U2835 (N_2835,N_1190,N_1401);
xor U2836 (N_2836,N_1455,N_1132);
or U2837 (N_2837,N_1134,N_1785);
nor U2838 (N_2838,N_1881,N_1441);
xnor U2839 (N_2839,N_1373,N_1522);
and U2840 (N_2840,N_1692,N_1289);
or U2841 (N_2841,N_1349,N_1047);
or U2842 (N_2842,N_1101,N_1824);
and U2843 (N_2843,N_1338,N_1305);
xnor U2844 (N_2844,N_1883,N_1923);
xnor U2845 (N_2845,N_1297,N_1294);
nor U2846 (N_2846,N_1532,N_1620);
or U2847 (N_2847,N_1423,N_1208);
and U2848 (N_2848,N_1240,N_1899);
nor U2849 (N_2849,N_1347,N_1812);
nand U2850 (N_2850,N_1440,N_1433);
nor U2851 (N_2851,N_1824,N_1829);
or U2852 (N_2852,N_1251,N_1942);
xor U2853 (N_2853,N_1797,N_1625);
xnor U2854 (N_2854,N_1281,N_1714);
nand U2855 (N_2855,N_1925,N_1933);
or U2856 (N_2856,N_1421,N_1173);
nor U2857 (N_2857,N_1899,N_1449);
nand U2858 (N_2858,N_1485,N_1897);
nand U2859 (N_2859,N_1759,N_1427);
nand U2860 (N_2860,N_1574,N_1523);
nor U2861 (N_2861,N_1168,N_1448);
nor U2862 (N_2862,N_1048,N_1039);
nor U2863 (N_2863,N_1633,N_1735);
or U2864 (N_2864,N_1935,N_1111);
xnor U2865 (N_2865,N_1761,N_1309);
nand U2866 (N_2866,N_1797,N_1518);
or U2867 (N_2867,N_1361,N_1166);
or U2868 (N_2868,N_1957,N_1755);
or U2869 (N_2869,N_1409,N_1829);
nand U2870 (N_2870,N_1958,N_1400);
nor U2871 (N_2871,N_1490,N_1996);
and U2872 (N_2872,N_1808,N_1160);
or U2873 (N_2873,N_1530,N_1603);
nand U2874 (N_2874,N_1211,N_1678);
xnor U2875 (N_2875,N_1634,N_1686);
or U2876 (N_2876,N_1773,N_1080);
and U2877 (N_2877,N_1693,N_1265);
or U2878 (N_2878,N_1881,N_1664);
xnor U2879 (N_2879,N_1863,N_1730);
or U2880 (N_2880,N_1290,N_1968);
nand U2881 (N_2881,N_1286,N_1465);
or U2882 (N_2882,N_1252,N_1021);
nor U2883 (N_2883,N_1113,N_1178);
xnor U2884 (N_2884,N_1544,N_1193);
or U2885 (N_2885,N_1911,N_1097);
xnor U2886 (N_2886,N_1371,N_1785);
and U2887 (N_2887,N_1623,N_1087);
xnor U2888 (N_2888,N_1790,N_1201);
nor U2889 (N_2889,N_1667,N_1975);
nand U2890 (N_2890,N_1128,N_1901);
xnor U2891 (N_2891,N_1985,N_1710);
nor U2892 (N_2892,N_1331,N_1085);
nand U2893 (N_2893,N_1135,N_1619);
nand U2894 (N_2894,N_1408,N_1135);
nand U2895 (N_2895,N_1842,N_1298);
nor U2896 (N_2896,N_1668,N_1894);
nand U2897 (N_2897,N_1652,N_1715);
nor U2898 (N_2898,N_1913,N_1881);
and U2899 (N_2899,N_1182,N_1099);
or U2900 (N_2900,N_1167,N_1959);
nor U2901 (N_2901,N_1201,N_1313);
nor U2902 (N_2902,N_1454,N_1508);
and U2903 (N_2903,N_1622,N_1182);
nand U2904 (N_2904,N_1089,N_1561);
xor U2905 (N_2905,N_1775,N_1637);
or U2906 (N_2906,N_1885,N_1187);
nand U2907 (N_2907,N_1739,N_1490);
xor U2908 (N_2908,N_1483,N_1554);
or U2909 (N_2909,N_1377,N_1858);
nor U2910 (N_2910,N_1714,N_1522);
and U2911 (N_2911,N_1956,N_1577);
or U2912 (N_2912,N_1255,N_1258);
nor U2913 (N_2913,N_1653,N_1842);
nor U2914 (N_2914,N_1348,N_1290);
xnor U2915 (N_2915,N_1922,N_1897);
xnor U2916 (N_2916,N_1363,N_1118);
xnor U2917 (N_2917,N_1662,N_1709);
and U2918 (N_2918,N_1112,N_1410);
or U2919 (N_2919,N_1972,N_1475);
xnor U2920 (N_2920,N_1696,N_1141);
xnor U2921 (N_2921,N_1449,N_1687);
nor U2922 (N_2922,N_1190,N_1643);
or U2923 (N_2923,N_1700,N_1862);
xor U2924 (N_2924,N_1855,N_1188);
nand U2925 (N_2925,N_1924,N_1934);
xor U2926 (N_2926,N_1271,N_1927);
or U2927 (N_2927,N_1659,N_1295);
or U2928 (N_2928,N_1761,N_1657);
nor U2929 (N_2929,N_1552,N_1226);
nor U2930 (N_2930,N_1711,N_1782);
or U2931 (N_2931,N_1542,N_1985);
and U2932 (N_2932,N_1289,N_1337);
or U2933 (N_2933,N_1271,N_1191);
nand U2934 (N_2934,N_1244,N_1846);
xnor U2935 (N_2935,N_1988,N_1093);
nand U2936 (N_2936,N_1438,N_1698);
nand U2937 (N_2937,N_1085,N_1598);
nand U2938 (N_2938,N_1637,N_1087);
nand U2939 (N_2939,N_1329,N_1509);
or U2940 (N_2940,N_1529,N_1130);
or U2941 (N_2941,N_1443,N_1841);
or U2942 (N_2942,N_1177,N_1112);
or U2943 (N_2943,N_1641,N_1038);
nor U2944 (N_2944,N_1794,N_1939);
nor U2945 (N_2945,N_1279,N_1111);
xor U2946 (N_2946,N_1981,N_1572);
nand U2947 (N_2947,N_1326,N_1424);
xor U2948 (N_2948,N_1520,N_1791);
nor U2949 (N_2949,N_1305,N_1172);
nand U2950 (N_2950,N_1503,N_1098);
nor U2951 (N_2951,N_1317,N_1219);
and U2952 (N_2952,N_1202,N_1960);
nand U2953 (N_2953,N_1359,N_1617);
nor U2954 (N_2954,N_1927,N_1258);
nor U2955 (N_2955,N_1050,N_1525);
and U2956 (N_2956,N_1692,N_1443);
nand U2957 (N_2957,N_1782,N_1411);
or U2958 (N_2958,N_1750,N_1714);
and U2959 (N_2959,N_1262,N_1081);
nor U2960 (N_2960,N_1469,N_1814);
nor U2961 (N_2961,N_1884,N_1486);
or U2962 (N_2962,N_1995,N_1976);
or U2963 (N_2963,N_1717,N_1324);
nor U2964 (N_2964,N_1460,N_1047);
xnor U2965 (N_2965,N_1436,N_1906);
xnor U2966 (N_2966,N_1106,N_1006);
and U2967 (N_2967,N_1747,N_1621);
or U2968 (N_2968,N_1085,N_1178);
and U2969 (N_2969,N_1234,N_1042);
nor U2970 (N_2970,N_1135,N_1725);
xnor U2971 (N_2971,N_1305,N_1295);
nand U2972 (N_2972,N_1558,N_1552);
and U2973 (N_2973,N_1932,N_1976);
nor U2974 (N_2974,N_1454,N_1729);
and U2975 (N_2975,N_1034,N_1098);
xor U2976 (N_2976,N_1142,N_1760);
nor U2977 (N_2977,N_1641,N_1908);
xnor U2978 (N_2978,N_1157,N_1889);
nor U2979 (N_2979,N_1318,N_1327);
or U2980 (N_2980,N_1759,N_1348);
xnor U2981 (N_2981,N_1990,N_1869);
or U2982 (N_2982,N_1218,N_1963);
or U2983 (N_2983,N_1061,N_1318);
and U2984 (N_2984,N_1008,N_1825);
or U2985 (N_2985,N_1745,N_1099);
nand U2986 (N_2986,N_1672,N_1111);
nand U2987 (N_2987,N_1861,N_1340);
or U2988 (N_2988,N_1214,N_1143);
xnor U2989 (N_2989,N_1202,N_1609);
or U2990 (N_2990,N_1310,N_1936);
and U2991 (N_2991,N_1115,N_1419);
nand U2992 (N_2992,N_1937,N_1605);
xnor U2993 (N_2993,N_1270,N_1345);
xor U2994 (N_2994,N_1506,N_1841);
nor U2995 (N_2995,N_1158,N_1673);
and U2996 (N_2996,N_1653,N_1080);
nand U2997 (N_2997,N_1699,N_1818);
nand U2998 (N_2998,N_1051,N_1090);
and U2999 (N_2999,N_1743,N_1008);
and U3000 (N_3000,N_2320,N_2575);
nand U3001 (N_3001,N_2249,N_2263);
xor U3002 (N_3002,N_2574,N_2980);
nand U3003 (N_3003,N_2146,N_2487);
or U3004 (N_3004,N_2592,N_2940);
xor U3005 (N_3005,N_2906,N_2224);
and U3006 (N_3006,N_2774,N_2846);
nand U3007 (N_3007,N_2864,N_2298);
and U3008 (N_3008,N_2710,N_2450);
nor U3009 (N_3009,N_2326,N_2213);
nor U3010 (N_3010,N_2888,N_2470);
and U3011 (N_3011,N_2546,N_2393);
and U3012 (N_3012,N_2388,N_2511);
and U3013 (N_3013,N_2581,N_2957);
or U3014 (N_3014,N_2629,N_2438);
nor U3015 (N_3015,N_2795,N_2212);
or U3016 (N_3016,N_2893,N_2221);
and U3017 (N_3017,N_2429,N_2069);
nand U3018 (N_3018,N_2641,N_2382);
nor U3019 (N_3019,N_2262,N_2228);
nand U3020 (N_3020,N_2352,N_2242);
nand U3021 (N_3021,N_2348,N_2480);
xor U3022 (N_3022,N_2192,N_2937);
and U3023 (N_3023,N_2226,N_2189);
xor U3024 (N_3024,N_2457,N_2391);
nand U3025 (N_3025,N_2589,N_2597);
nor U3026 (N_3026,N_2593,N_2934);
xor U3027 (N_3027,N_2410,N_2079);
and U3028 (N_3028,N_2800,N_2271);
nand U3029 (N_3029,N_2977,N_2880);
nor U3030 (N_3030,N_2144,N_2314);
xor U3031 (N_3031,N_2067,N_2665);
nand U3032 (N_3032,N_2060,N_2055);
nor U3033 (N_3033,N_2380,N_2684);
nand U3034 (N_3034,N_2129,N_2993);
nand U3035 (N_3035,N_2538,N_2149);
and U3036 (N_3036,N_2343,N_2724);
nor U3037 (N_3037,N_2639,N_2720);
xor U3038 (N_3038,N_2825,N_2305);
nand U3039 (N_3039,N_2260,N_2034);
nor U3040 (N_3040,N_2117,N_2790);
nor U3041 (N_3041,N_2572,N_2495);
nor U3042 (N_3042,N_2090,N_2557);
nor U3043 (N_3043,N_2643,N_2194);
xnor U3044 (N_3044,N_2707,N_2103);
nor U3045 (N_3045,N_2679,N_2947);
nor U3046 (N_3046,N_2218,N_2231);
or U3047 (N_3047,N_2872,N_2176);
nor U3048 (N_3048,N_2038,N_2187);
xor U3049 (N_3049,N_2744,N_2281);
xor U3050 (N_3050,N_2664,N_2527);
or U3051 (N_3051,N_2373,N_2808);
nand U3052 (N_3052,N_2162,N_2489);
xor U3053 (N_3053,N_2716,N_2555);
nand U3054 (N_3054,N_2351,N_2497);
nand U3055 (N_3055,N_2304,N_2234);
nand U3056 (N_3056,N_2227,N_2919);
xor U3057 (N_3057,N_2950,N_2381);
xnor U3058 (N_3058,N_2119,N_2163);
nand U3059 (N_3059,N_2990,N_2016);
xor U3060 (N_3060,N_2726,N_2195);
and U3061 (N_3061,N_2412,N_2843);
and U3062 (N_3062,N_2731,N_2289);
and U3063 (N_3063,N_2703,N_2496);
nor U3064 (N_3064,N_2803,N_2600);
or U3065 (N_3065,N_2396,N_2237);
or U3066 (N_3066,N_2723,N_2165);
nor U3067 (N_3067,N_2591,N_2233);
or U3068 (N_3068,N_2246,N_2157);
nand U3069 (N_3069,N_2930,N_2668);
or U3070 (N_3070,N_2503,N_2653);
or U3071 (N_3071,N_2960,N_2137);
or U3072 (N_3072,N_2788,N_2899);
xor U3073 (N_3073,N_2634,N_2911);
and U3074 (N_3074,N_2462,N_2344);
and U3075 (N_3075,N_2984,N_2595);
xnor U3076 (N_3076,N_2070,N_2755);
and U3077 (N_3077,N_2920,N_2091);
and U3078 (N_3078,N_2644,N_2026);
nand U3079 (N_3079,N_2471,N_2245);
xnor U3080 (N_3080,N_2037,N_2540);
and U3081 (N_3081,N_2501,N_2717);
nand U3082 (N_3082,N_2126,N_2883);
nor U3083 (N_3083,N_2513,N_2436);
or U3084 (N_3084,N_2338,N_2833);
and U3085 (N_3085,N_2901,N_2686);
and U3086 (N_3086,N_2324,N_2764);
or U3087 (N_3087,N_2309,N_2181);
or U3088 (N_3088,N_2287,N_2905);
and U3089 (N_3089,N_2140,N_2075);
or U3090 (N_3090,N_2523,N_2935);
xnor U3091 (N_3091,N_2064,N_2578);
nor U3092 (N_3092,N_2619,N_2273);
nand U3093 (N_3093,N_2904,N_2448);
xor U3094 (N_3094,N_2669,N_2625);
xnor U3095 (N_3095,N_2371,N_2473);
nor U3096 (N_3096,N_2204,N_2709);
nor U3097 (N_3097,N_2863,N_2355);
nand U3098 (N_3098,N_2422,N_2778);
nand U3099 (N_3099,N_2995,N_2131);
nand U3100 (N_3100,N_2536,N_2301);
nor U3101 (N_3101,N_2399,N_2022);
nand U3102 (N_3102,N_2549,N_2004);
and U3103 (N_3103,N_2706,N_2111);
and U3104 (N_3104,N_2292,N_2431);
nand U3105 (N_3105,N_2084,N_2678);
or U3106 (N_3106,N_2005,N_2188);
nand U3107 (N_3107,N_2965,N_2838);
nand U3108 (N_3108,N_2630,N_2942);
nor U3109 (N_3109,N_2890,N_2282);
nand U3110 (N_3110,N_2518,N_2214);
or U3111 (N_3111,N_2868,N_2076);
nand U3112 (N_3112,N_2676,N_2582);
xnor U3113 (N_3113,N_2742,N_2831);
or U3114 (N_3114,N_2924,N_2252);
or U3115 (N_3115,N_2345,N_2244);
or U3116 (N_3116,N_2319,N_2491);
nor U3117 (N_3117,N_2584,N_2257);
and U3118 (N_3118,N_2847,N_2000);
xnor U3119 (N_3119,N_2730,N_2892);
or U3120 (N_3120,N_2693,N_2078);
nand U3121 (N_3121,N_2248,N_2692);
nand U3122 (N_3122,N_2398,N_2297);
nand U3123 (N_3123,N_2108,N_2419);
and U3124 (N_3124,N_2095,N_2804);
nand U3125 (N_3125,N_2832,N_2138);
and U3126 (N_3126,N_2830,N_2941);
nor U3127 (N_3127,N_2492,N_2982);
nor U3128 (N_3128,N_2606,N_2670);
nor U3129 (N_3129,N_2981,N_2970);
nand U3130 (N_3130,N_2082,N_2943);
or U3131 (N_3131,N_2631,N_2923);
nor U3132 (N_3132,N_2506,N_2465);
and U3133 (N_3133,N_2087,N_2862);
nor U3134 (N_3134,N_2402,N_2397);
nand U3135 (N_3135,N_2010,N_2921);
or U3136 (N_3136,N_2636,N_2418);
or U3137 (N_3137,N_2505,N_2784);
nand U3138 (N_3138,N_2395,N_2116);
nand U3139 (N_3139,N_2598,N_2529);
and U3140 (N_3140,N_2913,N_2931);
xor U3141 (N_3141,N_2469,N_2533);
nor U3142 (N_3142,N_2541,N_2528);
or U3143 (N_3143,N_2858,N_2269);
nor U3144 (N_3144,N_2929,N_2295);
xor U3145 (N_3145,N_2135,N_2059);
and U3146 (N_3146,N_2002,N_2561);
xnor U3147 (N_3147,N_2551,N_2699);
or U3148 (N_3148,N_2334,N_2829);
and U3149 (N_3149,N_2142,N_2948);
or U3150 (N_3150,N_2805,N_2253);
and U3151 (N_3151,N_2250,N_2278);
nor U3152 (N_3152,N_2855,N_2413);
xnor U3153 (N_3153,N_2183,N_2277);
and U3154 (N_3154,N_2918,N_2682);
or U3155 (N_3155,N_2276,N_2816);
xor U3156 (N_3156,N_2001,N_2737);
nand U3157 (N_3157,N_2308,N_2484);
nor U3158 (N_3158,N_2270,N_2877);
or U3159 (N_3159,N_2360,N_2514);
xnor U3160 (N_3160,N_2907,N_2322);
nand U3161 (N_3161,N_2640,N_2766);
nand U3162 (N_3162,N_2488,N_2346);
or U3163 (N_3163,N_2675,N_2017);
and U3164 (N_3164,N_2882,N_2066);
xor U3165 (N_3165,N_2086,N_2792);
and U3166 (N_3166,N_2186,N_2903);
or U3167 (N_3167,N_2379,N_2417);
nor U3168 (N_3168,N_2736,N_2364);
nor U3169 (N_3169,N_2733,N_2425);
and U3170 (N_3170,N_2121,N_2871);
nand U3171 (N_3171,N_2207,N_2687);
and U3172 (N_3172,N_2439,N_2433);
and U3173 (N_3173,N_2894,N_2875);
and U3174 (N_3174,N_2392,N_2077);
xor U3175 (N_3175,N_2559,N_2172);
nand U3176 (N_3176,N_2945,N_2167);
xnor U3177 (N_3177,N_2760,N_2812);
nor U3178 (N_3178,N_2601,N_2842);
or U3179 (N_3179,N_2377,N_2032);
or U3180 (N_3180,N_2756,N_2255);
or U3181 (N_3181,N_2718,N_2081);
and U3182 (N_3182,N_2562,N_2548);
and U3183 (N_3183,N_2021,N_2220);
or U3184 (N_3184,N_2337,N_2407);
nor U3185 (N_3185,N_2007,N_2696);
and U3186 (N_3186,N_2867,N_2586);
nand U3187 (N_3187,N_2467,N_2190);
and U3188 (N_3188,N_2300,N_2012);
xor U3189 (N_3189,N_2746,N_2761);
and U3190 (N_3190,N_2938,N_2383);
or U3191 (N_3191,N_2106,N_2910);
nand U3192 (N_3192,N_2147,N_2169);
xor U3193 (N_3193,N_2599,N_2751);
or U3194 (N_3194,N_2876,N_2748);
xor U3195 (N_3195,N_2041,N_2112);
nand U3196 (N_3196,N_2652,N_2018);
nand U3197 (N_3197,N_2850,N_2596);
or U3198 (N_3198,N_2762,N_2908);
nand U3199 (N_3199,N_2099,N_2810);
or U3200 (N_3200,N_2254,N_2118);
or U3201 (N_3201,N_2400,N_2158);
and U3202 (N_3202,N_2535,N_2783);
nand U3203 (N_3203,N_2912,N_2564);
nor U3204 (N_3204,N_2992,N_2288);
or U3205 (N_3205,N_2148,N_2628);
nand U3206 (N_3206,N_2421,N_2133);
nand U3207 (N_3207,N_2658,N_2689);
nand U3208 (N_3208,N_2524,N_2985);
nand U3209 (N_3209,N_2240,N_2885);
and U3210 (N_3210,N_2753,N_2083);
nor U3211 (N_3211,N_2044,N_2585);
or U3212 (N_3212,N_2280,N_2811);
or U3213 (N_3213,N_2655,N_2747);
nand U3214 (N_3214,N_2014,N_2145);
and U3215 (N_3215,N_2602,N_2519);
nand U3216 (N_3216,N_2650,N_2657);
or U3217 (N_3217,N_2437,N_2114);
nor U3218 (N_3218,N_2312,N_2268);
nand U3219 (N_3219,N_2442,N_2779);
nand U3220 (N_3220,N_2427,N_2366);
nand U3221 (N_3221,N_2008,N_2335);
xor U3222 (N_3222,N_2780,N_2915);
or U3223 (N_3223,N_2897,N_2443);
nand U3224 (N_3224,N_2841,N_2532);
or U3225 (N_3225,N_2386,N_2860);
or U3226 (N_3226,N_2362,N_2035);
or U3227 (N_3227,N_2754,N_2475);
nand U3228 (N_3228,N_2196,N_2180);
nor U3229 (N_3229,N_2356,N_2460);
nor U3230 (N_3230,N_2136,N_2485);
nand U3231 (N_3231,N_2411,N_2109);
xor U3232 (N_3232,N_2807,N_2115);
xor U3233 (N_3233,N_2886,N_2306);
and U3234 (N_3234,N_2547,N_2879);
and U3235 (N_3235,N_2458,N_2818);
nor U3236 (N_3236,N_2614,N_2656);
xor U3237 (N_3237,N_2205,N_2329);
xor U3238 (N_3238,N_2284,N_2235);
and U3239 (N_3239,N_2568,N_2758);
xor U3240 (N_3240,N_2030,N_2347);
nor U3241 (N_3241,N_2100,N_2521);
nor U3242 (N_3242,N_2368,N_2113);
xor U3243 (N_3243,N_2236,N_2019);
or U3244 (N_3244,N_2516,N_2836);
nor U3245 (N_3245,N_2517,N_2033);
or U3246 (N_3246,N_2522,N_2123);
and U3247 (N_3247,N_2952,N_2445);
nand U3248 (N_3248,N_2608,N_2698);
nor U3249 (N_3249,N_2768,N_2098);
or U3250 (N_3250,N_2702,N_2542);
xnor U3251 (N_3251,N_2478,N_2615);
and U3252 (N_3252,N_2962,N_2241);
xnor U3253 (N_3253,N_2721,N_2325);
xor U3254 (N_3254,N_2525,N_2928);
xnor U3255 (N_3255,N_2141,N_2949);
nand U3256 (N_3256,N_2387,N_2056);
and U3257 (N_3257,N_2006,N_2375);
and U3258 (N_3258,N_2331,N_2683);
nor U3259 (N_3259,N_2127,N_2040);
nor U3260 (N_3260,N_2865,N_2174);
or U3261 (N_3261,N_2197,N_2624);
xnor U3262 (N_3262,N_2583,N_2428);
and U3263 (N_3263,N_2384,N_2027);
nand U3264 (N_3264,N_2358,N_2594);
xnor U3265 (N_3265,N_2185,N_2844);
and U3266 (N_3266,N_2376,N_2617);
or U3267 (N_3267,N_2560,N_2936);
nand U3268 (N_3268,N_2565,N_2739);
or U3269 (N_3269,N_2456,N_2062);
nand U3270 (N_3270,N_2861,N_2944);
nand U3271 (N_3271,N_2130,N_2459);
or U3272 (N_3272,N_2453,N_2217);
nand U3273 (N_3273,N_2092,N_2983);
nor U3274 (N_3274,N_2434,N_2061);
xor U3275 (N_3275,N_2787,N_2323);
and U3276 (N_3276,N_2691,N_2677);
and U3277 (N_3277,N_2203,N_2449);
and U3278 (N_3278,N_2216,N_2215);
and U3279 (N_3279,N_2821,N_2685);
xor U3280 (N_3280,N_2406,N_2620);
nor U3281 (N_3281,N_2011,N_2094);
or U3282 (N_3282,N_2202,N_2315);
nand U3283 (N_3283,N_2953,N_2638);
nor U3284 (N_3284,N_2283,N_2390);
and U3285 (N_3285,N_2068,N_2156);
xor U3286 (N_3286,N_2420,N_2660);
nand U3287 (N_3287,N_2151,N_2740);
nor U3288 (N_3288,N_2802,N_2961);
and U3289 (N_3289,N_2814,N_2490);
nand U3290 (N_3290,N_2729,N_2463);
or U3291 (N_3291,N_2285,N_2697);
nor U3292 (N_3292,N_2430,N_2925);
xor U3293 (N_3293,N_2279,N_2175);
and U3294 (N_3294,N_2367,N_2058);
xor U3295 (N_3295,N_2531,N_2666);
or U3296 (N_3296,N_2963,N_2946);
nor U3297 (N_3297,N_2013,N_2290);
or U3298 (N_3298,N_2820,N_2073);
nand U3299 (N_3299,N_2193,N_2835);
and U3300 (N_3300,N_2849,N_2991);
nand U3301 (N_3301,N_2712,N_2354);
or U3302 (N_3302,N_2303,N_2155);
nor U3303 (N_3303,N_2772,N_2570);
nor U3304 (N_3304,N_2239,N_2072);
nand U3305 (N_3305,N_2797,N_2662);
and U3306 (N_3306,N_2622,N_2286);
xor U3307 (N_3307,N_2461,N_2139);
and U3308 (N_3308,N_2435,N_2455);
and U3309 (N_3309,N_2317,N_2201);
nand U3310 (N_3310,N_2837,N_2318);
nor U3311 (N_3311,N_2799,N_2667);
nand U3312 (N_3312,N_2102,N_2752);
nand U3313 (N_3313,N_2566,N_2369);
nor U3314 (N_3314,N_2869,N_2472);
xor U3315 (N_3315,N_2122,N_2745);
and U3316 (N_3316,N_2793,N_2681);
nand U3317 (N_3317,N_2482,N_2047);
nand U3318 (N_3318,N_2050,N_2827);
xnor U3319 (N_3319,N_2230,N_2432);
or U3320 (N_3320,N_2646,N_2579);
or U3321 (N_3321,N_2711,N_2974);
or U3322 (N_3322,N_2336,N_2967);
nand U3323 (N_3323,N_2857,N_2782);
nor U3324 (N_3324,N_2705,N_2603);
or U3325 (N_3325,N_2848,N_2101);
nand U3326 (N_3326,N_2968,N_2749);
or U3327 (N_3327,N_2637,N_2840);
nand U3328 (N_3328,N_2713,N_2986);
and U3329 (N_3329,N_2958,N_2852);
xnor U3330 (N_3330,N_2039,N_2553);
nor U3331 (N_3331,N_2372,N_2895);
nand U3332 (N_3332,N_2266,N_2854);
nand U3333 (N_3333,N_2604,N_2153);
and U3334 (N_3334,N_2571,N_2370);
or U3335 (N_3335,N_2020,N_2642);
nor U3336 (N_3336,N_2510,N_2889);
and U3337 (N_3337,N_2105,N_2357);
nand U3338 (N_3338,N_2817,N_2870);
xnor U3339 (N_3339,N_2446,N_2359);
nor U3340 (N_3340,N_2587,N_2161);
nor U3341 (N_3341,N_2259,N_2704);
and U3342 (N_3342,N_2024,N_2588);
nand U3343 (N_3343,N_2509,N_2333);
xor U3344 (N_3344,N_2184,N_2451);
xnor U3345 (N_3345,N_2576,N_2632);
or U3346 (N_3346,N_2046,N_2023);
or U3347 (N_3347,N_2232,N_2859);
nand U3348 (N_3348,N_2577,N_2361);
nor U3349 (N_3349,N_2623,N_2671);
and U3350 (N_3350,N_2499,N_2914);
or U3351 (N_3351,N_2539,N_2464);
or U3352 (N_3352,N_2441,N_2403);
or U3353 (N_3353,N_2826,N_2672);
xor U3354 (N_3354,N_2074,N_2563);
xnor U3355 (N_3355,N_2674,N_2654);
xnor U3356 (N_3356,N_2211,N_2688);
xnor U3357 (N_3357,N_2989,N_2474);
and U3358 (N_3358,N_2734,N_2612);
nor U3359 (N_3359,N_2311,N_2182);
nor U3360 (N_3360,N_2468,N_2649);
and U3361 (N_3361,N_2727,N_2627);
nand U3362 (N_3362,N_2975,N_2477);
nor U3363 (N_3363,N_2349,N_2498);
or U3364 (N_3364,N_2104,N_2537);
and U3365 (N_3365,N_2902,N_2964);
nor U3366 (N_3366,N_2222,N_2916);
or U3367 (N_3367,N_2243,N_2447);
nand U3368 (N_3368,N_2313,N_2408);
nor U3369 (N_3369,N_2385,N_2770);
nand U3370 (N_3370,N_2168,N_2159);
and U3371 (N_3371,N_2927,N_2229);
nor U3372 (N_3372,N_2049,N_2444);
or U3373 (N_3373,N_2776,N_2272);
nor U3374 (N_3374,N_2680,N_2173);
xor U3375 (N_3375,N_2789,N_2741);
nor U3376 (N_3376,N_2694,N_2796);
xor U3377 (N_3377,N_2881,N_2342);
and U3378 (N_3378,N_2426,N_2951);
nand U3379 (N_3379,N_2558,N_2609);
nand U3380 (N_3380,N_2423,N_2708);
and U3381 (N_3381,N_2900,N_2618);
and U3382 (N_3382,N_2926,N_2164);
nor U3383 (N_3383,N_2258,N_2878);
xor U3384 (N_3384,N_2663,N_2891);
nand U3385 (N_3385,N_2120,N_2052);
or U3386 (N_3386,N_2813,N_2512);
xnor U3387 (N_3387,N_2898,N_2610);
xnor U3388 (N_3388,N_2028,N_2648);
or U3389 (N_3389,N_2715,N_2097);
or U3390 (N_3390,N_2401,N_2917);
nor U3391 (N_3391,N_2554,N_2966);
or U3392 (N_3392,N_2996,N_2569);
or U3393 (N_3393,N_2978,N_2722);
nor U3394 (N_3394,N_2363,N_2015);
or U3395 (N_3395,N_2500,N_2340);
nor U3396 (N_3396,N_2633,N_2042);
nand U3397 (N_3397,N_2590,N_2170);
nor U3398 (N_3398,N_2743,N_2088);
nor U3399 (N_3399,N_2209,N_2152);
and U3400 (N_3400,N_2988,N_2294);
or U3401 (N_3401,N_2063,N_2607);
or U3402 (N_3402,N_2543,N_2414);
xor U3403 (N_3403,N_2773,N_2972);
nor U3404 (N_3404,N_2009,N_2208);
nand U3405 (N_3405,N_2275,N_2695);
nor U3406 (N_3406,N_2053,N_2611);
nor U3407 (N_3407,N_2775,N_2806);
nor U3408 (N_3408,N_2124,N_2051);
and U3409 (N_3409,N_2732,N_2238);
nor U3410 (N_3410,N_2223,N_2483);
xor U3411 (N_3411,N_2302,N_2520);
xor U3412 (N_3412,N_2274,N_2219);
nand U3413 (N_3413,N_2556,N_2374);
nor U3414 (N_3414,N_2405,N_2031);
nand U3415 (N_3415,N_2828,N_2476);
xnor U3416 (N_3416,N_2178,N_2866);
nand U3417 (N_3417,N_2404,N_2544);
nand U3418 (N_3418,N_2316,N_2494);
xnor U3419 (N_3419,N_2251,N_2763);
or U3420 (N_3420,N_2552,N_2132);
and U3421 (N_3421,N_2339,N_2873);
nor U3422 (N_3422,N_2341,N_2296);
nor U3423 (N_3423,N_2481,N_2029);
xor U3424 (N_3424,N_2690,N_2166);
nand U3425 (N_3425,N_2987,N_2466);
nand U3426 (N_3426,N_2959,N_2191);
or U3427 (N_3427,N_2834,N_2424);
xor U3428 (N_3428,N_2791,N_2080);
nor U3429 (N_3429,N_2997,N_2714);
nand U3430 (N_3430,N_2054,N_2939);
nor U3431 (N_3431,N_2332,N_2976);
or U3432 (N_3432,N_2110,N_2365);
xnor U3433 (N_3433,N_2310,N_2291);
or U3434 (N_3434,N_2125,N_2932);
xnor U3435 (N_3435,N_2307,N_2267);
nand U3436 (N_3436,N_2096,N_2526);
nor U3437 (N_3437,N_2179,N_2065);
nand U3438 (N_3438,N_2328,N_2819);
nand U3439 (N_3439,N_2200,N_2093);
xnor U3440 (N_3440,N_2378,N_2839);
nor U3441 (N_3441,N_2973,N_2621);
nor U3442 (N_3442,N_2801,N_2504);
nor U3443 (N_3443,N_2160,N_2394);
nand U3444 (N_3444,N_2545,N_2824);
nand U3445 (N_3445,N_2651,N_2735);
nor U3446 (N_3446,N_2700,N_2673);
xnor U3447 (N_3447,N_2922,N_2409);
xnor U3448 (N_3448,N_2043,N_2823);
and U3449 (N_3449,N_2321,N_2036);
xor U3450 (N_3450,N_2719,N_2225);
and U3451 (N_3451,N_2171,N_2210);
xor U3452 (N_3452,N_2389,N_2003);
nand U3453 (N_3453,N_2661,N_2057);
xor U3454 (N_3454,N_2261,N_2567);
nor U3455 (N_3455,N_2786,N_2955);
xor U3456 (N_3456,N_2605,N_2198);
nand U3457 (N_3457,N_2256,N_2851);
xnor U3458 (N_3458,N_2769,N_2502);
nor U3459 (N_3459,N_2933,N_2896);
or U3460 (N_3460,N_2454,N_2750);
nand U3461 (N_3461,N_2767,N_2853);
or U3462 (N_3462,N_2822,N_2327);
nor U3463 (N_3463,N_2777,N_2330);
xor U3464 (N_3464,N_2508,N_2645);
xor U3465 (N_3465,N_2994,N_2728);
nor U3466 (N_3466,N_2534,N_2515);
nor U3467 (N_3467,N_2264,N_2048);
and U3468 (N_3468,N_2150,N_2247);
xor U3469 (N_3469,N_2299,N_2440);
xnor U3470 (N_3470,N_2025,N_2350);
or U3471 (N_3471,N_2635,N_2486);
nor U3472 (N_3472,N_2479,N_2507);
xor U3473 (N_3473,N_2909,N_2969);
nand U3474 (N_3474,N_2573,N_2659);
xor U3475 (N_3475,N_2845,N_2998);
xnor U3476 (N_3476,N_2452,N_2874);
and U3477 (N_3477,N_2971,N_2206);
xnor U3478 (N_3478,N_2085,N_2415);
nor U3479 (N_3479,N_2798,N_2979);
and U3480 (N_3480,N_2134,N_2416);
or U3481 (N_3481,N_2626,N_2701);
nor U3482 (N_3482,N_2154,N_2765);
nand U3483 (N_3483,N_2071,N_2884);
and U3484 (N_3484,N_2954,N_2887);
nand U3485 (N_3485,N_2293,N_2530);
nor U3486 (N_3486,N_2045,N_2771);
or U3487 (N_3487,N_2616,N_2738);
and U3488 (N_3488,N_2493,N_2759);
and U3489 (N_3489,N_2550,N_2353);
and U3490 (N_3490,N_2781,N_2856);
nand U3491 (N_3491,N_2128,N_2143);
xor U3492 (N_3492,N_2613,N_2089);
xnor U3493 (N_3493,N_2647,N_2815);
or U3494 (N_3494,N_2107,N_2757);
nand U3495 (N_3495,N_2265,N_2999);
xnor U3496 (N_3496,N_2580,N_2199);
nor U3497 (N_3497,N_2794,N_2956);
xnor U3498 (N_3498,N_2177,N_2785);
and U3499 (N_3499,N_2725,N_2809);
and U3500 (N_3500,N_2928,N_2640);
and U3501 (N_3501,N_2261,N_2347);
xnor U3502 (N_3502,N_2780,N_2965);
nand U3503 (N_3503,N_2535,N_2391);
nand U3504 (N_3504,N_2034,N_2007);
nor U3505 (N_3505,N_2956,N_2674);
nor U3506 (N_3506,N_2388,N_2767);
nor U3507 (N_3507,N_2395,N_2118);
or U3508 (N_3508,N_2147,N_2270);
nor U3509 (N_3509,N_2584,N_2004);
and U3510 (N_3510,N_2193,N_2405);
nor U3511 (N_3511,N_2360,N_2347);
and U3512 (N_3512,N_2251,N_2070);
nand U3513 (N_3513,N_2858,N_2802);
nor U3514 (N_3514,N_2587,N_2016);
or U3515 (N_3515,N_2097,N_2507);
xnor U3516 (N_3516,N_2673,N_2166);
nand U3517 (N_3517,N_2240,N_2190);
or U3518 (N_3518,N_2011,N_2417);
xor U3519 (N_3519,N_2782,N_2855);
or U3520 (N_3520,N_2635,N_2569);
and U3521 (N_3521,N_2160,N_2609);
or U3522 (N_3522,N_2545,N_2102);
xnor U3523 (N_3523,N_2554,N_2704);
or U3524 (N_3524,N_2965,N_2920);
and U3525 (N_3525,N_2747,N_2101);
nand U3526 (N_3526,N_2942,N_2441);
nand U3527 (N_3527,N_2169,N_2199);
xnor U3528 (N_3528,N_2428,N_2196);
nor U3529 (N_3529,N_2647,N_2438);
nor U3530 (N_3530,N_2034,N_2370);
and U3531 (N_3531,N_2645,N_2110);
nor U3532 (N_3532,N_2040,N_2594);
and U3533 (N_3533,N_2882,N_2661);
nand U3534 (N_3534,N_2451,N_2519);
and U3535 (N_3535,N_2239,N_2196);
or U3536 (N_3536,N_2469,N_2547);
or U3537 (N_3537,N_2364,N_2978);
and U3538 (N_3538,N_2080,N_2753);
and U3539 (N_3539,N_2640,N_2734);
nand U3540 (N_3540,N_2934,N_2070);
xnor U3541 (N_3541,N_2327,N_2859);
nand U3542 (N_3542,N_2534,N_2622);
nand U3543 (N_3543,N_2992,N_2936);
nand U3544 (N_3544,N_2147,N_2027);
xnor U3545 (N_3545,N_2333,N_2554);
xnor U3546 (N_3546,N_2065,N_2411);
nand U3547 (N_3547,N_2363,N_2859);
or U3548 (N_3548,N_2719,N_2358);
nor U3549 (N_3549,N_2118,N_2857);
and U3550 (N_3550,N_2945,N_2070);
or U3551 (N_3551,N_2167,N_2695);
or U3552 (N_3552,N_2943,N_2090);
nand U3553 (N_3553,N_2783,N_2962);
nand U3554 (N_3554,N_2975,N_2932);
or U3555 (N_3555,N_2040,N_2737);
nor U3556 (N_3556,N_2408,N_2803);
nand U3557 (N_3557,N_2485,N_2372);
xnor U3558 (N_3558,N_2304,N_2543);
and U3559 (N_3559,N_2513,N_2025);
nand U3560 (N_3560,N_2268,N_2845);
and U3561 (N_3561,N_2944,N_2494);
and U3562 (N_3562,N_2836,N_2231);
and U3563 (N_3563,N_2638,N_2486);
nor U3564 (N_3564,N_2752,N_2384);
nand U3565 (N_3565,N_2229,N_2417);
nor U3566 (N_3566,N_2675,N_2784);
and U3567 (N_3567,N_2728,N_2762);
xor U3568 (N_3568,N_2061,N_2181);
nand U3569 (N_3569,N_2387,N_2680);
nand U3570 (N_3570,N_2389,N_2189);
xnor U3571 (N_3571,N_2960,N_2065);
nor U3572 (N_3572,N_2329,N_2235);
nand U3573 (N_3573,N_2590,N_2482);
and U3574 (N_3574,N_2810,N_2700);
nor U3575 (N_3575,N_2795,N_2735);
xor U3576 (N_3576,N_2963,N_2108);
xor U3577 (N_3577,N_2301,N_2483);
or U3578 (N_3578,N_2841,N_2013);
or U3579 (N_3579,N_2735,N_2144);
and U3580 (N_3580,N_2480,N_2562);
or U3581 (N_3581,N_2247,N_2198);
xor U3582 (N_3582,N_2582,N_2793);
xor U3583 (N_3583,N_2395,N_2946);
nor U3584 (N_3584,N_2865,N_2389);
nor U3585 (N_3585,N_2723,N_2226);
and U3586 (N_3586,N_2940,N_2032);
or U3587 (N_3587,N_2975,N_2228);
or U3588 (N_3588,N_2113,N_2690);
nor U3589 (N_3589,N_2504,N_2922);
xor U3590 (N_3590,N_2669,N_2016);
nand U3591 (N_3591,N_2075,N_2907);
xor U3592 (N_3592,N_2768,N_2360);
xor U3593 (N_3593,N_2062,N_2247);
nand U3594 (N_3594,N_2722,N_2303);
or U3595 (N_3595,N_2599,N_2008);
nand U3596 (N_3596,N_2276,N_2801);
nand U3597 (N_3597,N_2013,N_2516);
nor U3598 (N_3598,N_2702,N_2966);
nand U3599 (N_3599,N_2878,N_2449);
nor U3600 (N_3600,N_2322,N_2277);
or U3601 (N_3601,N_2294,N_2544);
or U3602 (N_3602,N_2646,N_2344);
xor U3603 (N_3603,N_2041,N_2191);
xnor U3604 (N_3604,N_2444,N_2398);
nand U3605 (N_3605,N_2100,N_2614);
xor U3606 (N_3606,N_2861,N_2544);
xnor U3607 (N_3607,N_2143,N_2194);
or U3608 (N_3608,N_2147,N_2315);
and U3609 (N_3609,N_2163,N_2619);
nand U3610 (N_3610,N_2947,N_2498);
xnor U3611 (N_3611,N_2952,N_2448);
and U3612 (N_3612,N_2670,N_2376);
xor U3613 (N_3613,N_2835,N_2336);
nor U3614 (N_3614,N_2850,N_2502);
or U3615 (N_3615,N_2592,N_2097);
nor U3616 (N_3616,N_2880,N_2112);
and U3617 (N_3617,N_2126,N_2038);
and U3618 (N_3618,N_2837,N_2617);
nor U3619 (N_3619,N_2031,N_2019);
xnor U3620 (N_3620,N_2393,N_2291);
nor U3621 (N_3621,N_2995,N_2436);
nor U3622 (N_3622,N_2431,N_2410);
xor U3623 (N_3623,N_2941,N_2947);
xnor U3624 (N_3624,N_2560,N_2801);
nor U3625 (N_3625,N_2432,N_2868);
nand U3626 (N_3626,N_2056,N_2798);
nor U3627 (N_3627,N_2214,N_2172);
nor U3628 (N_3628,N_2480,N_2389);
xnor U3629 (N_3629,N_2649,N_2889);
xor U3630 (N_3630,N_2893,N_2645);
or U3631 (N_3631,N_2627,N_2535);
and U3632 (N_3632,N_2126,N_2930);
nor U3633 (N_3633,N_2683,N_2392);
xor U3634 (N_3634,N_2080,N_2521);
xor U3635 (N_3635,N_2766,N_2006);
xnor U3636 (N_3636,N_2472,N_2809);
and U3637 (N_3637,N_2628,N_2566);
nor U3638 (N_3638,N_2447,N_2290);
nor U3639 (N_3639,N_2940,N_2559);
xor U3640 (N_3640,N_2411,N_2099);
and U3641 (N_3641,N_2059,N_2989);
xnor U3642 (N_3642,N_2770,N_2107);
and U3643 (N_3643,N_2631,N_2736);
xor U3644 (N_3644,N_2146,N_2840);
or U3645 (N_3645,N_2578,N_2374);
nor U3646 (N_3646,N_2076,N_2355);
nor U3647 (N_3647,N_2849,N_2012);
or U3648 (N_3648,N_2564,N_2157);
or U3649 (N_3649,N_2931,N_2001);
or U3650 (N_3650,N_2767,N_2158);
or U3651 (N_3651,N_2971,N_2335);
nor U3652 (N_3652,N_2376,N_2789);
xnor U3653 (N_3653,N_2689,N_2562);
or U3654 (N_3654,N_2042,N_2413);
and U3655 (N_3655,N_2818,N_2493);
or U3656 (N_3656,N_2250,N_2917);
xor U3657 (N_3657,N_2271,N_2740);
nor U3658 (N_3658,N_2196,N_2638);
xnor U3659 (N_3659,N_2296,N_2003);
or U3660 (N_3660,N_2883,N_2020);
xor U3661 (N_3661,N_2917,N_2877);
or U3662 (N_3662,N_2045,N_2175);
nor U3663 (N_3663,N_2925,N_2567);
and U3664 (N_3664,N_2604,N_2944);
or U3665 (N_3665,N_2719,N_2252);
or U3666 (N_3666,N_2299,N_2974);
xor U3667 (N_3667,N_2971,N_2226);
nor U3668 (N_3668,N_2106,N_2809);
xnor U3669 (N_3669,N_2682,N_2033);
nor U3670 (N_3670,N_2671,N_2095);
nand U3671 (N_3671,N_2008,N_2899);
nand U3672 (N_3672,N_2982,N_2990);
or U3673 (N_3673,N_2195,N_2224);
nand U3674 (N_3674,N_2439,N_2541);
nor U3675 (N_3675,N_2719,N_2220);
or U3676 (N_3676,N_2281,N_2376);
or U3677 (N_3677,N_2433,N_2956);
or U3678 (N_3678,N_2766,N_2960);
and U3679 (N_3679,N_2335,N_2932);
nor U3680 (N_3680,N_2909,N_2529);
nand U3681 (N_3681,N_2145,N_2036);
xnor U3682 (N_3682,N_2097,N_2559);
and U3683 (N_3683,N_2644,N_2754);
or U3684 (N_3684,N_2646,N_2536);
and U3685 (N_3685,N_2659,N_2892);
and U3686 (N_3686,N_2115,N_2849);
nor U3687 (N_3687,N_2030,N_2857);
and U3688 (N_3688,N_2223,N_2395);
xor U3689 (N_3689,N_2664,N_2110);
and U3690 (N_3690,N_2309,N_2335);
xnor U3691 (N_3691,N_2794,N_2249);
nand U3692 (N_3692,N_2685,N_2192);
nor U3693 (N_3693,N_2365,N_2621);
and U3694 (N_3694,N_2090,N_2455);
xor U3695 (N_3695,N_2510,N_2387);
nand U3696 (N_3696,N_2257,N_2971);
nand U3697 (N_3697,N_2693,N_2046);
and U3698 (N_3698,N_2723,N_2216);
nand U3699 (N_3699,N_2328,N_2511);
or U3700 (N_3700,N_2114,N_2337);
nor U3701 (N_3701,N_2435,N_2487);
and U3702 (N_3702,N_2499,N_2712);
and U3703 (N_3703,N_2379,N_2969);
xnor U3704 (N_3704,N_2505,N_2005);
nand U3705 (N_3705,N_2809,N_2397);
nand U3706 (N_3706,N_2842,N_2360);
and U3707 (N_3707,N_2915,N_2245);
nand U3708 (N_3708,N_2115,N_2639);
nand U3709 (N_3709,N_2956,N_2176);
and U3710 (N_3710,N_2602,N_2671);
xnor U3711 (N_3711,N_2460,N_2104);
nor U3712 (N_3712,N_2053,N_2464);
or U3713 (N_3713,N_2325,N_2281);
and U3714 (N_3714,N_2229,N_2832);
nor U3715 (N_3715,N_2765,N_2849);
or U3716 (N_3716,N_2457,N_2331);
xor U3717 (N_3717,N_2468,N_2310);
xnor U3718 (N_3718,N_2629,N_2642);
nor U3719 (N_3719,N_2713,N_2706);
nand U3720 (N_3720,N_2163,N_2846);
or U3721 (N_3721,N_2446,N_2658);
or U3722 (N_3722,N_2319,N_2794);
or U3723 (N_3723,N_2990,N_2950);
and U3724 (N_3724,N_2011,N_2870);
nor U3725 (N_3725,N_2393,N_2838);
xnor U3726 (N_3726,N_2129,N_2310);
nor U3727 (N_3727,N_2812,N_2608);
and U3728 (N_3728,N_2622,N_2554);
and U3729 (N_3729,N_2931,N_2373);
nor U3730 (N_3730,N_2219,N_2735);
and U3731 (N_3731,N_2003,N_2360);
or U3732 (N_3732,N_2277,N_2290);
or U3733 (N_3733,N_2447,N_2334);
and U3734 (N_3734,N_2256,N_2815);
nor U3735 (N_3735,N_2273,N_2264);
or U3736 (N_3736,N_2420,N_2433);
xor U3737 (N_3737,N_2084,N_2513);
xor U3738 (N_3738,N_2484,N_2215);
and U3739 (N_3739,N_2960,N_2932);
nor U3740 (N_3740,N_2636,N_2505);
nor U3741 (N_3741,N_2864,N_2009);
nor U3742 (N_3742,N_2486,N_2423);
nor U3743 (N_3743,N_2320,N_2773);
nand U3744 (N_3744,N_2901,N_2733);
xnor U3745 (N_3745,N_2067,N_2632);
or U3746 (N_3746,N_2098,N_2491);
nor U3747 (N_3747,N_2348,N_2612);
xor U3748 (N_3748,N_2338,N_2890);
or U3749 (N_3749,N_2999,N_2239);
nor U3750 (N_3750,N_2329,N_2981);
nor U3751 (N_3751,N_2105,N_2080);
nor U3752 (N_3752,N_2903,N_2662);
and U3753 (N_3753,N_2654,N_2644);
and U3754 (N_3754,N_2975,N_2884);
nand U3755 (N_3755,N_2226,N_2133);
nand U3756 (N_3756,N_2850,N_2562);
and U3757 (N_3757,N_2683,N_2944);
nor U3758 (N_3758,N_2530,N_2410);
or U3759 (N_3759,N_2509,N_2212);
xor U3760 (N_3760,N_2284,N_2964);
nor U3761 (N_3761,N_2733,N_2913);
or U3762 (N_3762,N_2462,N_2972);
xnor U3763 (N_3763,N_2224,N_2234);
and U3764 (N_3764,N_2984,N_2056);
and U3765 (N_3765,N_2411,N_2899);
nor U3766 (N_3766,N_2624,N_2451);
xnor U3767 (N_3767,N_2339,N_2551);
and U3768 (N_3768,N_2448,N_2181);
nand U3769 (N_3769,N_2596,N_2560);
xor U3770 (N_3770,N_2857,N_2850);
nor U3771 (N_3771,N_2693,N_2443);
nor U3772 (N_3772,N_2604,N_2793);
or U3773 (N_3773,N_2650,N_2609);
and U3774 (N_3774,N_2212,N_2938);
nor U3775 (N_3775,N_2151,N_2962);
or U3776 (N_3776,N_2410,N_2516);
and U3777 (N_3777,N_2701,N_2109);
and U3778 (N_3778,N_2710,N_2515);
and U3779 (N_3779,N_2301,N_2684);
or U3780 (N_3780,N_2929,N_2618);
nor U3781 (N_3781,N_2043,N_2689);
nor U3782 (N_3782,N_2491,N_2749);
xnor U3783 (N_3783,N_2786,N_2920);
or U3784 (N_3784,N_2576,N_2667);
nand U3785 (N_3785,N_2953,N_2494);
nor U3786 (N_3786,N_2672,N_2539);
or U3787 (N_3787,N_2590,N_2595);
nor U3788 (N_3788,N_2402,N_2975);
or U3789 (N_3789,N_2807,N_2184);
nand U3790 (N_3790,N_2502,N_2120);
xnor U3791 (N_3791,N_2026,N_2524);
and U3792 (N_3792,N_2473,N_2626);
nor U3793 (N_3793,N_2146,N_2298);
and U3794 (N_3794,N_2151,N_2704);
nor U3795 (N_3795,N_2965,N_2535);
or U3796 (N_3796,N_2783,N_2353);
xor U3797 (N_3797,N_2935,N_2642);
nand U3798 (N_3798,N_2759,N_2588);
and U3799 (N_3799,N_2785,N_2885);
xor U3800 (N_3800,N_2480,N_2185);
nand U3801 (N_3801,N_2820,N_2612);
and U3802 (N_3802,N_2684,N_2319);
or U3803 (N_3803,N_2508,N_2494);
or U3804 (N_3804,N_2477,N_2491);
and U3805 (N_3805,N_2374,N_2575);
nor U3806 (N_3806,N_2694,N_2703);
nor U3807 (N_3807,N_2408,N_2319);
or U3808 (N_3808,N_2060,N_2698);
and U3809 (N_3809,N_2341,N_2645);
nor U3810 (N_3810,N_2789,N_2475);
nor U3811 (N_3811,N_2225,N_2535);
nor U3812 (N_3812,N_2336,N_2104);
or U3813 (N_3813,N_2544,N_2364);
nor U3814 (N_3814,N_2588,N_2921);
xor U3815 (N_3815,N_2131,N_2496);
and U3816 (N_3816,N_2214,N_2267);
xor U3817 (N_3817,N_2831,N_2089);
and U3818 (N_3818,N_2119,N_2315);
or U3819 (N_3819,N_2463,N_2596);
nor U3820 (N_3820,N_2438,N_2631);
nor U3821 (N_3821,N_2149,N_2921);
and U3822 (N_3822,N_2493,N_2137);
nor U3823 (N_3823,N_2703,N_2205);
and U3824 (N_3824,N_2117,N_2650);
nand U3825 (N_3825,N_2735,N_2776);
nand U3826 (N_3826,N_2574,N_2379);
xnor U3827 (N_3827,N_2998,N_2842);
nor U3828 (N_3828,N_2101,N_2187);
xnor U3829 (N_3829,N_2187,N_2029);
and U3830 (N_3830,N_2510,N_2434);
xor U3831 (N_3831,N_2935,N_2646);
nand U3832 (N_3832,N_2735,N_2842);
nand U3833 (N_3833,N_2800,N_2456);
and U3834 (N_3834,N_2192,N_2445);
and U3835 (N_3835,N_2825,N_2083);
nor U3836 (N_3836,N_2408,N_2789);
nand U3837 (N_3837,N_2488,N_2535);
and U3838 (N_3838,N_2515,N_2690);
nand U3839 (N_3839,N_2394,N_2787);
nor U3840 (N_3840,N_2078,N_2517);
nand U3841 (N_3841,N_2347,N_2720);
nand U3842 (N_3842,N_2485,N_2509);
nand U3843 (N_3843,N_2440,N_2013);
xnor U3844 (N_3844,N_2467,N_2260);
nor U3845 (N_3845,N_2605,N_2704);
nor U3846 (N_3846,N_2258,N_2273);
nand U3847 (N_3847,N_2917,N_2315);
and U3848 (N_3848,N_2605,N_2471);
xor U3849 (N_3849,N_2331,N_2456);
xor U3850 (N_3850,N_2730,N_2452);
nand U3851 (N_3851,N_2281,N_2024);
nand U3852 (N_3852,N_2407,N_2703);
or U3853 (N_3853,N_2931,N_2834);
xor U3854 (N_3854,N_2511,N_2808);
nand U3855 (N_3855,N_2399,N_2930);
nor U3856 (N_3856,N_2330,N_2661);
or U3857 (N_3857,N_2590,N_2334);
nand U3858 (N_3858,N_2809,N_2477);
or U3859 (N_3859,N_2564,N_2872);
nand U3860 (N_3860,N_2403,N_2547);
xor U3861 (N_3861,N_2370,N_2952);
nor U3862 (N_3862,N_2047,N_2929);
and U3863 (N_3863,N_2905,N_2375);
or U3864 (N_3864,N_2547,N_2394);
nand U3865 (N_3865,N_2321,N_2772);
nor U3866 (N_3866,N_2070,N_2164);
and U3867 (N_3867,N_2033,N_2858);
xor U3868 (N_3868,N_2738,N_2613);
nand U3869 (N_3869,N_2854,N_2276);
xnor U3870 (N_3870,N_2785,N_2182);
nor U3871 (N_3871,N_2119,N_2890);
xor U3872 (N_3872,N_2694,N_2200);
nor U3873 (N_3873,N_2670,N_2807);
xnor U3874 (N_3874,N_2107,N_2326);
or U3875 (N_3875,N_2227,N_2576);
nand U3876 (N_3876,N_2814,N_2656);
or U3877 (N_3877,N_2840,N_2387);
nor U3878 (N_3878,N_2621,N_2389);
or U3879 (N_3879,N_2851,N_2182);
nor U3880 (N_3880,N_2152,N_2313);
xor U3881 (N_3881,N_2902,N_2039);
and U3882 (N_3882,N_2068,N_2193);
nor U3883 (N_3883,N_2652,N_2351);
and U3884 (N_3884,N_2539,N_2330);
or U3885 (N_3885,N_2344,N_2935);
nor U3886 (N_3886,N_2898,N_2113);
nor U3887 (N_3887,N_2917,N_2641);
nand U3888 (N_3888,N_2618,N_2751);
nor U3889 (N_3889,N_2377,N_2966);
xor U3890 (N_3890,N_2712,N_2273);
or U3891 (N_3891,N_2941,N_2887);
and U3892 (N_3892,N_2388,N_2800);
and U3893 (N_3893,N_2947,N_2885);
or U3894 (N_3894,N_2324,N_2956);
or U3895 (N_3895,N_2811,N_2581);
xnor U3896 (N_3896,N_2551,N_2269);
and U3897 (N_3897,N_2996,N_2397);
xnor U3898 (N_3898,N_2954,N_2392);
or U3899 (N_3899,N_2357,N_2831);
nand U3900 (N_3900,N_2379,N_2651);
nor U3901 (N_3901,N_2592,N_2199);
nand U3902 (N_3902,N_2603,N_2938);
xor U3903 (N_3903,N_2151,N_2414);
or U3904 (N_3904,N_2419,N_2477);
or U3905 (N_3905,N_2267,N_2422);
or U3906 (N_3906,N_2598,N_2410);
nand U3907 (N_3907,N_2878,N_2979);
and U3908 (N_3908,N_2314,N_2176);
nor U3909 (N_3909,N_2487,N_2339);
and U3910 (N_3910,N_2838,N_2270);
nor U3911 (N_3911,N_2459,N_2794);
or U3912 (N_3912,N_2564,N_2429);
or U3913 (N_3913,N_2498,N_2121);
xnor U3914 (N_3914,N_2637,N_2182);
xor U3915 (N_3915,N_2938,N_2805);
xor U3916 (N_3916,N_2304,N_2644);
nand U3917 (N_3917,N_2788,N_2327);
or U3918 (N_3918,N_2893,N_2027);
and U3919 (N_3919,N_2219,N_2473);
and U3920 (N_3920,N_2487,N_2130);
nand U3921 (N_3921,N_2420,N_2657);
nand U3922 (N_3922,N_2904,N_2964);
nand U3923 (N_3923,N_2030,N_2706);
nor U3924 (N_3924,N_2995,N_2641);
or U3925 (N_3925,N_2004,N_2220);
or U3926 (N_3926,N_2539,N_2212);
and U3927 (N_3927,N_2562,N_2396);
nand U3928 (N_3928,N_2717,N_2839);
nand U3929 (N_3929,N_2783,N_2411);
nor U3930 (N_3930,N_2156,N_2650);
nor U3931 (N_3931,N_2607,N_2513);
or U3932 (N_3932,N_2522,N_2150);
and U3933 (N_3933,N_2467,N_2985);
nor U3934 (N_3934,N_2430,N_2188);
nor U3935 (N_3935,N_2477,N_2711);
nand U3936 (N_3936,N_2755,N_2474);
nand U3937 (N_3937,N_2374,N_2842);
and U3938 (N_3938,N_2109,N_2374);
nand U3939 (N_3939,N_2521,N_2330);
nand U3940 (N_3940,N_2421,N_2186);
xnor U3941 (N_3941,N_2511,N_2853);
or U3942 (N_3942,N_2904,N_2379);
nand U3943 (N_3943,N_2562,N_2752);
xnor U3944 (N_3944,N_2266,N_2061);
nand U3945 (N_3945,N_2695,N_2410);
nor U3946 (N_3946,N_2552,N_2380);
and U3947 (N_3947,N_2921,N_2267);
nor U3948 (N_3948,N_2781,N_2097);
and U3949 (N_3949,N_2410,N_2800);
or U3950 (N_3950,N_2168,N_2895);
or U3951 (N_3951,N_2643,N_2219);
xor U3952 (N_3952,N_2261,N_2164);
nand U3953 (N_3953,N_2737,N_2974);
or U3954 (N_3954,N_2117,N_2640);
nand U3955 (N_3955,N_2423,N_2608);
xnor U3956 (N_3956,N_2240,N_2967);
xor U3957 (N_3957,N_2211,N_2743);
nor U3958 (N_3958,N_2751,N_2606);
xor U3959 (N_3959,N_2951,N_2975);
or U3960 (N_3960,N_2193,N_2314);
xor U3961 (N_3961,N_2600,N_2879);
or U3962 (N_3962,N_2126,N_2522);
or U3963 (N_3963,N_2849,N_2476);
or U3964 (N_3964,N_2996,N_2441);
xor U3965 (N_3965,N_2689,N_2655);
or U3966 (N_3966,N_2274,N_2127);
nor U3967 (N_3967,N_2439,N_2859);
nand U3968 (N_3968,N_2808,N_2524);
nor U3969 (N_3969,N_2236,N_2292);
nor U3970 (N_3970,N_2620,N_2787);
nand U3971 (N_3971,N_2524,N_2357);
or U3972 (N_3972,N_2766,N_2316);
or U3973 (N_3973,N_2897,N_2400);
or U3974 (N_3974,N_2092,N_2283);
or U3975 (N_3975,N_2199,N_2604);
and U3976 (N_3976,N_2061,N_2724);
and U3977 (N_3977,N_2462,N_2463);
xor U3978 (N_3978,N_2480,N_2542);
and U3979 (N_3979,N_2450,N_2194);
nand U3980 (N_3980,N_2127,N_2355);
or U3981 (N_3981,N_2255,N_2572);
nor U3982 (N_3982,N_2150,N_2853);
nor U3983 (N_3983,N_2249,N_2088);
xor U3984 (N_3984,N_2493,N_2649);
or U3985 (N_3985,N_2559,N_2944);
xnor U3986 (N_3986,N_2438,N_2123);
nor U3987 (N_3987,N_2154,N_2661);
and U3988 (N_3988,N_2348,N_2656);
or U3989 (N_3989,N_2514,N_2147);
and U3990 (N_3990,N_2687,N_2043);
nor U3991 (N_3991,N_2538,N_2350);
nand U3992 (N_3992,N_2497,N_2600);
and U3993 (N_3993,N_2663,N_2966);
xor U3994 (N_3994,N_2335,N_2051);
nor U3995 (N_3995,N_2540,N_2038);
and U3996 (N_3996,N_2655,N_2032);
or U3997 (N_3997,N_2277,N_2164);
xnor U3998 (N_3998,N_2698,N_2228);
and U3999 (N_3999,N_2479,N_2632);
nand U4000 (N_4000,N_3350,N_3845);
or U4001 (N_4001,N_3843,N_3818);
xor U4002 (N_4002,N_3157,N_3971);
nor U4003 (N_4003,N_3673,N_3007);
nor U4004 (N_4004,N_3160,N_3332);
nand U4005 (N_4005,N_3513,N_3055);
or U4006 (N_4006,N_3531,N_3143);
or U4007 (N_4007,N_3771,N_3993);
nand U4008 (N_4008,N_3838,N_3273);
and U4009 (N_4009,N_3260,N_3276);
nor U4010 (N_4010,N_3465,N_3825);
xnor U4011 (N_4011,N_3967,N_3446);
nor U4012 (N_4012,N_3431,N_3250);
and U4013 (N_4013,N_3682,N_3360);
and U4014 (N_4014,N_3256,N_3867);
nor U4015 (N_4015,N_3476,N_3297);
or U4016 (N_4016,N_3604,N_3738);
and U4017 (N_4017,N_3346,N_3268);
or U4018 (N_4018,N_3568,N_3100);
or U4019 (N_4019,N_3588,N_3869);
nand U4020 (N_4020,N_3364,N_3329);
nor U4021 (N_4021,N_3404,N_3596);
or U4022 (N_4022,N_3603,N_3048);
and U4023 (N_4023,N_3271,N_3621);
nand U4024 (N_4024,N_3963,N_3804);
or U4025 (N_4025,N_3930,N_3846);
xor U4026 (N_4026,N_3285,N_3123);
nand U4027 (N_4027,N_3079,N_3650);
nand U4028 (N_4028,N_3239,N_3909);
nand U4029 (N_4029,N_3395,N_3812);
nand U4030 (N_4030,N_3023,N_3317);
nand U4031 (N_4031,N_3799,N_3502);
nor U4032 (N_4032,N_3393,N_3154);
xnor U4033 (N_4033,N_3547,N_3454);
and U4034 (N_4034,N_3987,N_3555);
xor U4035 (N_4035,N_3684,N_3940);
xnor U4036 (N_4036,N_3182,N_3990);
or U4037 (N_4037,N_3607,N_3891);
and U4038 (N_4038,N_3169,N_3099);
xor U4039 (N_4039,N_3475,N_3235);
xnor U4040 (N_4040,N_3246,N_3075);
and U4041 (N_4041,N_3339,N_3102);
nand U4042 (N_4042,N_3559,N_3678);
or U4043 (N_4043,N_3549,N_3692);
or U4044 (N_4044,N_3952,N_3356);
nand U4045 (N_4045,N_3964,N_3690);
nand U4046 (N_4046,N_3462,N_3253);
nand U4047 (N_4047,N_3808,N_3855);
or U4048 (N_4048,N_3866,N_3649);
nor U4049 (N_4049,N_3831,N_3740);
nor U4050 (N_4050,N_3116,N_3674);
or U4051 (N_4051,N_3227,N_3355);
xnor U4052 (N_4052,N_3929,N_3449);
nor U4053 (N_4053,N_3716,N_3922);
nand U4054 (N_4054,N_3331,N_3597);
and U4055 (N_4055,N_3516,N_3626);
xnor U4056 (N_4056,N_3068,N_3892);
xnor U4057 (N_4057,N_3248,N_3191);
and U4058 (N_4058,N_3022,N_3354);
nor U4059 (N_4059,N_3464,N_3011);
nor U4060 (N_4060,N_3084,N_3905);
xnor U4061 (N_4061,N_3426,N_3608);
xor U4062 (N_4062,N_3323,N_3968);
and U4063 (N_4063,N_3830,N_3748);
nor U4064 (N_4064,N_3312,N_3732);
xnor U4065 (N_4065,N_3257,N_3915);
or U4066 (N_4066,N_3442,N_3082);
xnor U4067 (N_4067,N_3762,N_3036);
or U4068 (N_4068,N_3904,N_3910);
nor U4069 (N_4069,N_3844,N_3753);
and U4070 (N_4070,N_3814,N_3472);
nor U4071 (N_4071,N_3985,N_3939);
nand U4072 (N_4072,N_3936,N_3481);
and U4073 (N_4073,N_3816,N_3189);
nor U4074 (N_4074,N_3121,N_3719);
nor U4075 (N_4075,N_3410,N_3850);
nand U4076 (N_4076,N_3572,N_3875);
xor U4077 (N_4077,N_3744,N_3616);
nand U4078 (N_4078,N_3761,N_3721);
or U4079 (N_4079,N_3303,N_3292);
and U4080 (N_4080,N_3630,N_3113);
or U4081 (N_4081,N_3717,N_3293);
nand U4082 (N_4082,N_3645,N_3118);
and U4083 (N_4083,N_3252,N_3015);
nor U4084 (N_4084,N_3872,N_3402);
xnor U4085 (N_4085,N_3815,N_3708);
nor U4086 (N_4086,N_3991,N_3548);
nand U4087 (N_4087,N_3806,N_3210);
xor U4088 (N_4088,N_3745,N_3772);
nor U4089 (N_4089,N_3700,N_3515);
or U4090 (N_4090,N_3633,N_3265);
or U4091 (N_4091,N_3255,N_3617);
and U4092 (N_4092,N_3856,N_3853);
xor U4093 (N_4093,N_3437,N_3978);
xnor U4094 (N_4094,N_3860,N_3406);
or U4095 (N_4095,N_3918,N_3374);
and U4096 (N_4096,N_3385,N_3032);
nand U4097 (N_4097,N_3409,N_3724);
xor U4098 (N_4098,N_3507,N_3834);
xnor U4099 (N_4099,N_3709,N_3027);
nor U4100 (N_4100,N_3262,N_3398);
or U4101 (N_4101,N_3600,N_3270);
or U4102 (N_4102,N_3605,N_3370);
nand U4103 (N_4103,N_3319,N_3695);
xnor U4104 (N_4104,N_3399,N_3006);
nor U4105 (N_4105,N_3040,N_3474);
xnor U4106 (N_4106,N_3186,N_3888);
nand U4107 (N_4107,N_3284,N_3203);
or U4108 (N_4108,N_3612,N_3024);
or U4109 (N_4109,N_3640,N_3200);
nand U4110 (N_4110,N_3400,N_3304);
xnor U4111 (N_4111,N_3657,N_3897);
nor U4112 (N_4112,N_3881,N_3236);
nor U4113 (N_4113,N_3525,N_3050);
xnor U4114 (N_4114,N_3280,N_3141);
nor U4115 (N_4115,N_3619,N_3705);
nor U4116 (N_4116,N_3039,N_3688);
xor U4117 (N_4117,N_3057,N_3132);
nor U4118 (N_4118,N_3508,N_3676);
or U4119 (N_4119,N_3168,N_3587);
nand U4120 (N_4120,N_3278,N_3667);
nor U4121 (N_4121,N_3106,N_3517);
xor U4122 (N_4122,N_3539,N_3109);
nand U4123 (N_4123,N_3563,N_3043);
or U4124 (N_4124,N_3176,N_3908);
xnor U4125 (N_4125,N_3453,N_3025);
nor U4126 (N_4126,N_3163,N_3658);
nor U4127 (N_4127,N_3177,N_3927);
and U4128 (N_4128,N_3028,N_3122);
xor U4129 (N_4129,N_3158,N_3187);
xor U4130 (N_4130,N_3347,N_3571);
nand U4131 (N_4131,N_3198,N_3183);
xnor U4132 (N_4132,N_3433,N_3215);
nand U4133 (N_4133,N_3552,N_3672);
or U4134 (N_4134,N_3931,N_3219);
nand U4135 (N_4135,N_3598,N_3093);
and U4136 (N_4136,N_3359,N_3272);
or U4137 (N_4137,N_3396,N_3353);
xnor U4138 (N_4138,N_3903,N_3349);
or U4139 (N_4139,N_3880,N_3722);
or U4140 (N_4140,N_3958,N_3501);
nor U4141 (N_4141,N_3368,N_3311);
or U4142 (N_4142,N_3358,N_3938);
xor U4143 (N_4143,N_3144,N_3060);
nand U4144 (N_4144,N_3142,N_3697);
nor U4145 (N_4145,N_3989,N_3451);
or U4146 (N_4146,N_3702,N_3214);
or U4147 (N_4147,N_3521,N_3975);
or U4148 (N_4148,N_3233,N_3301);
or U4149 (N_4149,N_3240,N_3567);
and U4150 (N_4150,N_3403,N_3520);
xnor U4151 (N_4151,N_3792,N_3530);
nand U4152 (N_4152,N_3195,N_3833);
or U4153 (N_4153,N_3035,N_3333);
xor U4154 (N_4154,N_3627,N_3746);
or U4155 (N_4155,N_3942,N_3505);
nand U4156 (N_4156,N_3245,N_3727);
or U4157 (N_4157,N_3140,N_3582);
nor U4158 (N_4158,N_3147,N_3669);
nand U4159 (N_4159,N_3309,N_3886);
or U4160 (N_4160,N_3826,N_3718);
nor U4161 (N_4161,N_3483,N_3857);
nor U4162 (N_4162,N_3809,N_3149);
nor U4163 (N_4163,N_3120,N_3128);
or U4164 (N_4164,N_3326,N_3469);
or U4165 (N_4165,N_3794,N_3421);
xor U4166 (N_4166,N_3047,N_3486);
and U4167 (N_4167,N_3452,N_3334);
or U4168 (N_4168,N_3302,N_3456);
xnor U4169 (N_4169,N_3443,N_3973);
and U4170 (N_4170,N_3473,N_3221);
xnor U4171 (N_4171,N_3174,N_3523);
or U4172 (N_4172,N_3340,N_3008);
nand U4173 (N_4173,N_3294,N_3595);
nand U4174 (N_4174,N_3251,N_3184);
nand U4175 (N_4175,N_3490,N_3212);
and U4176 (N_4176,N_3434,N_3037);
nor U4177 (N_4177,N_3636,N_3056);
xnor U4178 (N_4178,N_3832,N_3254);
xor U4179 (N_4179,N_3824,N_3005);
or U4180 (N_4180,N_3119,N_3088);
and U4181 (N_4181,N_3228,N_3361);
nor U4182 (N_4182,N_3907,N_3108);
xor U4183 (N_4183,N_3059,N_3482);
or U4184 (N_4184,N_3192,N_3497);
nor U4185 (N_4185,N_3861,N_3033);
xor U4186 (N_4186,N_3208,N_3504);
nor U4187 (N_4187,N_3151,N_3923);
and U4188 (N_4188,N_3267,N_3041);
or U4189 (N_4189,N_3391,N_3749);
nor U4190 (N_4190,N_3207,N_3071);
and U4191 (N_4191,N_3901,N_3401);
or U4192 (N_4192,N_3247,N_3864);
xor U4193 (N_4193,N_3898,N_3540);
or U4194 (N_4194,N_3327,N_3791);
nand U4195 (N_4195,N_3310,N_3584);
or U4196 (N_4196,N_3185,N_3775);
or U4197 (N_4197,N_3817,N_3822);
and U4198 (N_4198,N_3703,N_3496);
nor U4199 (N_4199,N_3115,N_3444);
or U4200 (N_4200,N_3849,N_3668);
xnor U4201 (N_4201,N_3110,N_3069);
nor U4202 (N_4202,N_3042,N_3689);
xnor U4203 (N_4203,N_3639,N_3737);
or U4204 (N_4204,N_3381,N_3803);
xor U4205 (N_4205,N_3743,N_3495);
xnor U4206 (N_4206,N_3511,N_3801);
xor U4207 (N_4207,N_3769,N_3710);
nand U4208 (N_4208,N_3884,N_3053);
or U4209 (N_4209,N_3135,N_3786);
nor U4210 (N_4210,N_3983,N_3382);
or U4211 (N_4211,N_3599,N_3882);
and U4212 (N_4212,N_3887,N_3701);
or U4213 (N_4213,N_3779,N_3984);
or U4214 (N_4214,N_3463,N_3706);
or U4215 (N_4215,N_3279,N_3264);
or U4216 (N_4216,N_3492,N_3680);
nor U4217 (N_4217,N_3117,N_3004);
xnor U4218 (N_4218,N_3758,N_3150);
and U4219 (N_4219,N_3220,N_3405);
nor U4220 (N_4220,N_3181,N_3498);
nand U4221 (N_4221,N_3526,N_3167);
xor U4222 (N_4222,N_3031,N_3580);
nand U4223 (N_4223,N_3694,N_3629);
or U4224 (N_4224,N_3466,N_3556);
and U4225 (N_4225,N_3226,N_3029);
xnor U4226 (N_4226,N_3805,N_3665);
nor U4227 (N_4227,N_3238,N_3201);
or U4228 (N_4228,N_3981,N_3739);
nand U4229 (N_4229,N_3720,N_3655);
nor U4230 (N_4230,N_3757,N_3479);
xnor U4231 (N_4231,N_3911,N_3074);
and U4232 (N_4232,N_3581,N_3324);
and U4233 (N_4233,N_3105,N_3336);
nand U4234 (N_4234,N_3954,N_3367);
xor U4235 (N_4235,N_3087,N_3773);
nand U4236 (N_4236,N_3206,N_3145);
and U4237 (N_4237,N_3625,N_3615);
nor U4238 (N_4238,N_3107,N_3551);
nor U4239 (N_4239,N_3928,N_3419);
and U4240 (N_4240,N_3953,N_3286);
nor U4241 (N_4241,N_3766,N_3447);
nor U4242 (N_4242,N_3643,N_3190);
or U4243 (N_4243,N_3959,N_3133);
or U4244 (N_4244,N_3178,N_3995);
nand U4245 (N_4245,N_3536,N_3728);
nand U4246 (N_4246,N_3575,N_3593);
xor U4247 (N_4247,N_3261,N_3561);
nor U4248 (N_4248,N_3759,N_3211);
and U4249 (N_4249,N_3328,N_3380);
xnor U4250 (N_4250,N_3782,N_3545);
or U4251 (N_4251,N_3266,N_3979);
xor U4252 (N_4252,N_3179,N_3698);
or U4253 (N_4253,N_3237,N_3681);
nand U4254 (N_4254,N_3660,N_3944);
and U4255 (N_4255,N_3578,N_3124);
xor U4256 (N_4256,N_3675,N_3934);
nor U4257 (N_4257,N_3223,N_3620);
xnor U4258 (N_4258,N_3155,N_3742);
or U4259 (N_4259,N_3019,N_3982);
nand U4260 (N_4260,N_3683,N_3635);
nand U4261 (N_4261,N_3003,N_3914);
nand U4262 (N_4262,N_3977,N_3017);
nand U4263 (N_4263,N_3933,N_3275);
nor U4264 (N_4264,N_3893,N_3712);
and U4265 (N_4265,N_3009,N_3097);
nor U4266 (N_4266,N_3900,N_3366);
or U4267 (N_4267,N_3876,N_3654);
nand U4268 (N_4268,N_3529,N_3089);
or U4269 (N_4269,N_3579,N_3858);
nor U4270 (N_4270,N_3389,N_3172);
nand U4271 (N_4271,N_3244,N_3499);
nor U4272 (N_4272,N_3471,N_3429);
nor U4273 (N_4273,N_3081,N_3997);
or U4274 (N_4274,N_3819,N_3467);
and U4275 (N_4275,N_3685,N_3577);
and U4276 (N_4276,N_3095,N_3755);
nand U4277 (N_4277,N_3161,N_3715);
or U4278 (N_4278,N_3589,N_3585);
nor U4279 (N_4279,N_3802,N_3080);
nand U4280 (N_4280,N_3330,N_3197);
nor U4281 (N_4281,N_3734,N_3229);
nand U4282 (N_4282,N_3532,N_3662);
xnor U4283 (N_4283,N_3460,N_3136);
and U4284 (N_4284,N_3777,N_3554);
xnor U4285 (N_4285,N_3550,N_3687);
and U4286 (N_4286,N_3793,N_3624);
and U4287 (N_4287,N_3175,N_3798);
nor U4288 (N_4288,N_3926,N_3066);
and U4289 (N_4289,N_3205,N_3946);
nand U4290 (N_4290,N_3352,N_3980);
or U4291 (N_4291,N_3965,N_3859);
or U4292 (N_4292,N_3902,N_3064);
and U4293 (N_4293,N_3781,N_3455);
or U4294 (N_4294,N_3010,N_3423);
nand U4295 (N_4295,N_3194,N_3321);
nand U4296 (N_4296,N_3383,N_3494);
nand U4297 (N_4297,N_3924,N_3371);
and U4298 (N_4298,N_3836,N_3751);
nor U4299 (N_4299,N_3416,N_3125);
nor U4300 (N_4300,N_3774,N_3362);
or U4301 (N_4301,N_3341,N_3750);
nand U4302 (N_4302,N_3837,N_3566);
xnor U4303 (N_4303,N_3077,N_3765);
and U4304 (N_4304,N_3670,N_3527);
nand U4305 (N_4305,N_3591,N_3970);
nand U4306 (N_4306,N_3363,N_3188);
xnor U4307 (N_4307,N_3535,N_3012);
xnor U4308 (N_4308,N_3948,N_3691);
nand U4309 (N_4309,N_3756,N_3874);
nand U4310 (N_4310,N_3955,N_3112);
and U4311 (N_4311,N_3797,N_3659);
and U4312 (N_4312,N_3851,N_3972);
nand U4313 (N_4313,N_3537,N_3103);
nand U4314 (N_4314,N_3435,N_3001);
nand U4315 (N_4315,N_3351,N_3648);
xnor U4316 (N_4316,N_3308,N_3209);
nor U4317 (N_4317,N_3896,N_3384);
nand U4318 (N_4318,N_3863,N_3714);
and U4319 (N_4319,N_3146,N_3813);
nand U4320 (N_4320,N_3842,N_3916);
or U4321 (N_4321,N_3541,N_3852);
xor U4322 (N_4322,N_3974,N_3696);
and U4323 (N_4323,N_3484,N_3947);
and U4324 (N_4324,N_3518,N_3524);
or U4325 (N_4325,N_3018,N_3422);
xor U4326 (N_4326,N_3173,N_3038);
nand U4327 (N_4327,N_3570,N_3428);
xor U4328 (N_4328,N_3729,N_3795);
xnor U4329 (N_4329,N_3320,N_3436);
nand U4330 (N_4330,N_3956,N_3438);
nand U4331 (N_4331,N_3061,N_3470);
nor U4332 (N_4332,N_3306,N_3386);
or U4333 (N_4333,N_3165,N_3638);
nand U4334 (N_4334,N_3686,N_3148);
xor U4335 (N_4335,N_3586,N_3314);
nor U4336 (N_4336,N_3736,N_3249);
nand U4337 (N_4337,N_3564,N_3810);
nand U4338 (N_4338,N_3606,N_3919);
nand U4339 (N_4339,N_3894,N_3046);
xnor U4340 (N_4340,N_3768,N_3424);
and U4341 (N_4341,N_3634,N_3258);
and U4342 (N_4342,N_3637,N_3558);
nor U4343 (N_4343,N_3741,N_3534);
or U4344 (N_4344,N_3020,N_3218);
nor U4345 (N_4345,N_3234,N_3723);
xor U4346 (N_4346,N_3338,N_3425);
xor U4347 (N_4347,N_3274,N_3369);
nor U4348 (N_4348,N_3445,N_3661);
or U4349 (N_4349,N_3512,N_3828);
and U4350 (N_4350,N_3623,N_3785);
nor U4351 (N_4351,N_3085,N_3111);
nor U4352 (N_4352,N_3656,N_3514);
nand U4353 (N_4353,N_3092,N_3949);
xnor U4354 (N_4354,N_3733,N_3912);
or U4355 (N_4355,N_3839,N_3199);
and U4356 (N_4356,N_3357,N_3509);
or U4357 (N_4357,N_3315,N_3013);
or U4358 (N_4358,N_3291,N_3752);
and U4359 (N_4359,N_3413,N_3058);
and U4360 (N_4360,N_3171,N_3459);
and U4361 (N_4361,N_3754,N_3506);
and U4362 (N_4362,N_3618,N_3747);
nand U4363 (N_4363,N_3213,N_3461);
nand U4364 (N_4364,N_3217,N_3962);
and U4365 (N_4365,N_3560,N_3788);
nand U4366 (N_4366,N_3412,N_3835);
nand U4367 (N_4367,N_3131,N_3906);
and U4368 (N_4368,N_3296,N_3644);
xnor U4369 (N_4369,N_3034,N_3313);
xor U4370 (N_4370,N_3780,N_3969);
and U4371 (N_4371,N_3487,N_3241);
nor U4372 (N_4372,N_3281,N_3873);
xnor U4373 (N_4373,N_3420,N_3062);
nand U4374 (N_4374,N_3337,N_3827);
nand U4375 (N_4375,N_3784,N_3544);
and U4376 (N_4376,N_3295,N_3072);
nand U4377 (N_4377,N_3316,N_3493);
xor U4378 (N_4378,N_3992,N_3288);
xnor U4379 (N_4379,N_3343,N_3299);
xnor U4380 (N_4380,N_3538,N_3448);
and U4381 (N_4381,N_3298,N_3601);
xor U4382 (N_4382,N_3427,N_3565);
nand U4383 (N_4383,N_3522,N_3988);
nor U4384 (N_4384,N_3485,N_3305);
nor U4385 (N_4385,N_3647,N_3408);
nand U4386 (N_4386,N_3014,N_3129);
xor U4387 (N_4387,N_3044,N_3653);
xor U4388 (N_4388,N_3943,N_3488);
xor U4389 (N_4389,N_3546,N_3130);
xnor U4390 (N_4390,N_3932,N_3065);
nand U4391 (N_4391,N_3289,N_3776);
and U4392 (N_4392,N_3731,N_3713);
xnor U4393 (N_4393,N_3342,N_3372);
or U4394 (N_4394,N_3170,N_3913);
xor U4395 (N_4395,N_3821,N_3883);
and U4396 (N_4396,N_3344,N_3533);
nor U4397 (N_4397,N_3998,N_3016);
and U4398 (N_4398,N_3263,N_3994);
nor U4399 (N_4399,N_3628,N_3677);
nand U4400 (N_4400,N_3783,N_3999);
nor U4401 (N_4401,N_3073,N_3440);
and U4402 (N_4402,N_3478,N_3760);
nor U4403 (N_4403,N_3789,N_3083);
nand U4404 (N_4404,N_3457,N_3152);
nand U4405 (N_4405,N_3663,N_3283);
nand U4406 (N_4406,N_3300,N_3063);
and U4407 (N_4407,N_3373,N_3840);
and U4408 (N_4408,N_3242,N_3417);
or U4409 (N_4409,N_3439,N_3277);
nor U4410 (N_4410,N_3704,N_3138);
nor U4411 (N_4411,N_3823,N_3937);
nor U4412 (N_4412,N_3961,N_3622);
nand U4413 (N_4413,N_3807,N_3671);
nor U4414 (N_4414,N_3976,N_3432);
or U4415 (N_4415,N_3726,N_3491);
nor U4416 (N_4416,N_3614,N_3067);
and U4417 (N_4417,N_3921,N_3862);
or U4418 (N_4418,N_3945,N_3917);
nand U4419 (N_4419,N_3870,N_3847);
and U4420 (N_4420,N_3162,N_3193);
or U4421 (N_4421,N_3848,N_3335);
nor U4422 (N_4422,N_3202,N_3613);
xor U4423 (N_4423,N_3519,N_3725);
nor U4424 (N_4424,N_3811,N_3450);
xor U4425 (N_4425,N_3259,N_3414);
nand U4426 (N_4426,N_3610,N_3885);
nand U4427 (N_4427,N_3224,N_3957);
and U4428 (N_4428,N_3602,N_3026);
and U4429 (N_4429,N_3592,N_3376);
and U4430 (N_4430,N_3216,N_3679);
and U4431 (N_4431,N_3086,N_3841);
nor U4432 (N_4432,N_3574,N_3800);
nor U4433 (N_4433,N_3699,N_3418);
and U4434 (N_4434,N_3590,N_3282);
xor U4435 (N_4435,N_3094,N_3126);
or U4436 (N_4436,N_3707,N_3583);
or U4437 (N_4437,N_3764,N_3510);
nor U4438 (N_4438,N_3230,N_3153);
xnor U4439 (N_4439,N_3778,N_3269);
or U4440 (N_4440,N_3651,N_3854);
and U4441 (N_4441,N_3090,N_3325);
xor U4442 (N_4442,N_3387,N_3441);
and U4443 (N_4443,N_3407,N_3114);
nand U4444 (N_4444,N_3796,N_3002);
xnor U4445 (N_4445,N_3477,N_3225);
nor U4446 (N_4446,N_3646,N_3390);
nand U4447 (N_4447,N_3569,N_3950);
or U4448 (N_4448,N_3711,N_3134);
xnor U4449 (N_4449,N_3730,N_3735);
nand U4450 (N_4450,N_3632,N_3562);
nand U4451 (N_4451,N_3899,N_3345);
nand U4452 (N_4452,N_3127,N_3767);
xnor U4453 (N_4453,N_3895,N_3960);
nand U4454 (N_4454,N_3693,N_3049);
and U4455 (N_4455,N_3322,N_3166);
xor U4456 (N_4456,N_3232,N_3890);
nand U4457 (N_4457,N_3664,N_3091);
xnor U4458 (N_4458,N_3879,N_3489);
or U4459 (N_4459,N_3573,N_3480);
nor U4460 (N_4460,N_3652,N_3889);
or U4461 (N_4461,N_3503,N_3051);
nor U4462 (N_4462,N_3021,N_3379);
xnor U4463 (N_4463,N_3986,N_3318);
nand U4464 (N_4464,N_3770,N_3528);
and U4465 (N_4465,N_3243,N_3594);
and U4466 (N_4466,N_3156,N_3666);
nand U4467 (N_4467,N_3231,N_3392);
and U4468 (N_4468,N_3631,N_3164);
xor U4469 (N_4469,N_3951,N_3790);
and U4470 (N_4470,N_3641,N_3576);
or U4471 (N_4471,N_3543,N_3611);
nand U4472 (N_4472,N_3307,N_3137);
or U4473 (N_4473,N_3096,N_3553);
and U4474 (N_4474,N_3365,N_3500);
xor U4475 (N_4475,N_3101,N_3925);
nor U4476 (N_4476,N_3820,N_3871);
and U4477 (N_4477,N_3935,N_3098);
xnor U4478 (N_4478,N_3877,N_3787);
nor U4479 (N_4479,N_3868,N_3196);
nor U4480 (N_4480,N_3104,N_3394);
or U4481 (N_4481,N_3763,N_3458);
or U4482 (N_4482,N_3996,N_3378);
or U4483 (N_4483,N_3468,N_3030);
and U4484 (N_4484,N_3430,N_3878);
or U4485 (N_4485,N_3557,N_3941);
xnor U4486 (N_4486,N_3829,N_3070);
xnor U4487 (N_4487,N_3076,N_3222);
nand U4488 (N_4488,N_3078,N_3139);
and U4489 (N_4489,N_3045,N_3287);
xor U4490 (N_4490,N_3290,N_3966);
nand U4491 (N_4491,N_3865,N_3542);
and U4492 (N_4492,N_3052,N_3375);
and U4493 (N_4493,N_3415,N_3411);
and U4494 (N_4494,N_3348,N_3204);
xnor U4495 (N_4495,N_3180,N_3397);
xor U4496 (N_4496,N_3000,N_3609);
and U4497 (N_4497,N_3159,N_3388);
nand U4498 (N_4498,N_3920,N_3054);
nand U4499 (N_4499,N_3642,N_3377);
or U4500 (N_4500,N_3419,N_3173);
nand U4501 (N_4501,N_3626,N_3524);
or U4502 (N_4502,N_3364,N_3804);
nor U4503 (N_4503,N_3499,N_3283);
nand U4504 (N_4504,N_3890,N_3799);
and U4505 (N_4505,N_3362,N_3592);
xor U4506 (N_4506,N_3745,N_3771);
or U4507 (N_4507,N_3396,N_3126);
nor U4508 (N_4508,N_3352,N_3811);
nor U4509 (N_4509,N_3592,N_3282);
nor U4510 (N_4510,N_3154,N_3746);
and U4511 (N_4511,N_3907,N_3243);
nor U4512 (N_4512,N_3233,N_3261);
xnor U4513 (N_4513,N_3686,N_3316);
nor U4514 (N_4514,N_3890,N_3623);
nand U4515 (N_4515,N_3433,N_3744);
nand U4516 (N_4516,N_3588,N_3986);
and U4517 (N_4517,N_3400,N_3018);
and U4518 (N_4518,N_3600,N_3543);
nand U4519 (N_4519,N_3989,N_3199);
xor U4520 (N_4520,N_3300,N_3274);
nor U4521 (N_4521,N_3817,N_3162);
nor U4522 (N_4522,N_3609,N_3576);
or U4523 (N_4523,N_3593,N_3202);
and U4524 (N_4524,N_3351,N_3854);
or U4525 (N_4525,N_3605,N_3066);
xnor U4526 (N_4526,N_3038,N_3072);
nand U4527 (N_4527,N_3712,N_3981);
or U4528 (N_4528,N_3588,N_3675);
and U4529 (N_4529,N_3677,N_3939);
or U4530 (N_4530,N_3187,N_3661);
or U4531 (N_4531,N_3596,N_3623);
nor U4532 (N_4532,N_3403,N_3837);
xnor U4533 (N_4533,N_3305,N_3978);
or U4534 (N_4534,N_3176,N_3608);
and U4535 (N_4535,N_3117,N_3893);
nor U4536 (N_4536,N_3883,N_3890);
nand U4537 (N_4537,N_3217,N_3950);
nand U4538 (N_4538,N_3454,N_3415);
or U4539 (N_4539,N_3383,N_3515);
or U4540 (N_4540,N_3775,N_3424);
and U4541 (N_4541,N_3141,N_3386);
or U4542 (N_4542,N_3214,N_3785);
nor U4543 (N_4543,N_3553,N_3428);
nand U4544 (N_4544,N_3838,N_3545);
and U4545 (N_4545,N_3978,N_3431);
xor U4546 (N_4546,N_3419,N_3978);
nand U4547 (N_4547,N_3186,N_3562);
and U4548 (N_4548,N_3699,N_3271);
xnor U4549 (N_4549,N_3560,N_3927);
and U4550 (N_4550,N_3240,N_3925);
nor U4551 (N_4551,N_3640,N_3274);
xor U4552 (N_4552,N_3712,N_3163);
xor U4553 (N_4553,N_3495,N_3665);
nand U4554 (N_4554,N_3601,N_3732);
xor U4555 (N_4555,N_3166,N_3707);
and U4556 (N_4556,N_3435,N_3289);
and U4557 (N_4557,N_3266,N_3869);
xor U4558 (N_4558,N_3076,N_3915);
or U4559 (N_4559,N_3349,N_3182);
nor U4560 (N_4560,N_3200,N_3002);
or U4561 (N_4561,N_3842,N_3598);
nor U4562 (N_4562,N_3656,N_3599);
or U4563 (N_4563,N_3452,N_3521);
xor U4564 (N_4564,N_3596,N_3423);
and U4565 (N_4565,N_3699,N_3247);
xnor U4566 (N_4566,N_3435,N_3773);
and U4567 (N_4567,N_3441,N_3199);
xnor U4568 (N_4568,N_3275,N_3817);
nand U4569 (N_4569,N_3550,N_3190);
nand U4570 (N_4570,N_3619,N_3514);
xnor U4571 (N_4571,N_3531,N_3311);
or U4572 (N_4572,N_3364,N_3234);
nand U4573 (N_4573,N_3134,N_3213);
xor U4574 (N_4574,N_3502,N_3383);
nand U4575 (N_4575,N_3267,N_3746);
xor U4576 (N_4576,N_3638,N_3835);
xor U4577 (N_4577,N_3578,N_3378);
nor U4578 (N_4578,N_3168,N_3422);
nor U4579 (N_4579,N_3521,N_3691);
or U4580 (N_4580,N_3442,N_3755);
nor U4581 (N_4581,N_3826,N_3722);
nor U4582 (N_4582,N_3978,N_3485);
nand U4583 (N_4583,N_3928,N_3453);
or U4584 (N_4584,N_3129,N_3107);
and U4585 (N_4585,N_3476,N_3434);
and U4586 (N_4586,N_3990,N_3429);
xnor U4587 (N_4587,N_3779,N_3045);
nor U4588 (N_4588,N_3703,N_3569);
nand U4589 (N_4589,N_3250,N_3174);
nand U4590 (N_4590,N_3861,N_3678);
nand U4591 (N_4591,N_3084,N_3093);
nand U4592 (N_4592,N_3455,N_3637);
xnor U4593 (N_4593,N_3552,N_3549);
nand U4594 (N_4594,N_3218,N_3767);
nand U4595 (N_4595,N_3347,N_3436);
nor U4596 (N_4596,N_3193,N_3936);
nor U4597 (N_4597,N_3794,N_3994);
xor U4598 (N_4598,N_3812,N_3910);
or U4599 (N_4599,N_3485,N_3514);
xnor U4600 (N_4600,N_3782,N_3850);
nand U4601 (N_4601,N_3412,N_3391);
nand U4602 (N_4602,N_3349,N_3542);
nor U4603 (N_4603,N_3647,N_3989);
nor U4604 (N_4604,N_3569,N_3786);
nand U4605 (N_4605,N_3541,N_3933);
xnor U4606 (N_4606,N_3558,N_3557);
nand U4607 (N_4607,N_3108,N_3431);
nand U4608 (N_4608,N_3084,N_3087);
nand U4609 (N_4609,N_3965,N_3014);
nand U4610 (N_4610,N_3279,N_3276);
xor U4611 (N_4611,N_3243,N_3597);
nor U4612 (N_4612,N_3229,N_3629);
and U4613 (N_4613,N_3864,N_3414);
nor U4614 (N_4614,N_3996,N_3473);
nor U4615 (N_4615,N_3822,N_3410);
and U4616 (N_4616,N_3718,N_3487);
xor U4617 (N_4617,N_3505,N_3097);
or U4618 (N_4618,N_3502,N_3401);
xor U4619 (N_4619,N_3089,N_3903);
xor U4620 (N_4620,N_3734,N_3576);
nor U4621 (N_4621,N_3940,N_3730);
or U4622 (N_4622,N_3611,N_3667);
nor U4623 (N_4623,N_3656,N_3975);
and U4624 (N_4624,N_3129,N_3855);
nand U4625 (N_4625,N_3003,N_3464);
nand U4626 (N_4626,N_3864,N_3854);
nor U4627 (N_4627,N_3761,N_3906);
nor U4628 (N_4628,N_3844,N_3268);
xnor U4629 (N_4629,N_3381,N_3918);
or U4630 (N_4630,N_3969,N_3994);
nor U4631 (N_4631,N_3175,N_3067);
or U4632 (N_4632,N_3132,N_3427);
nand U4633 (N_4633,N_3794,N_3583);
or U4634 (N_4634,N_3791,N_3773);
xor U4635 (N_4635,N_3046,N_3140);
and U4636 (N_4636,N_3128,N_3357);
and U4637 (N_4637,N_3557,N_3829);
nor U4638 (N_4638,N_3444,N_3772);
nor U4639 (N_4639,N_3739,N_3523);
and U4640 (N_4640,N_3463,N_3782);
and U4641 (N_4641,N_3828,N_3935);
nand U4642 (N_4642,N_3341,N_3928);
or U4643 (N_4643,N_3959,N_3477);
nor U4644 (N_4644,N_3582,N_3481);
or U4645 (N_4645,N_3107,N_3750);
or U4646 (N_4646,N_3440,N_3782);
nand U4647 (N_4647,N_3173,N_3911);
and U4648 (N_4648,N_3998,N_3340);
and U4649 (N_4649,N_3755,N_3082);
nand U4650 (N_4650,N_3999,N_3746);
nor U4651 (N_4651,N_3526,N_3034);
xor U4652 (N_4652,N_3755,N_3187);
nand U4653 (N_4653,N_3820,N_3560);
nor U4654 (N_4654,N_3889,N_3113);
or U4655 (N_4655,N_3682,N_3708);
nor U4656 (N_4656,N_3176,N_3989);
nor U4657 (N_4657,N_3078,N_3754);
or U4658 (N_4658,N_3760,N_3985);
xor U4659 (N_4659,N_3551,N_3459);
xnor U4660 (N_4660,N_3402,N_3083);
and U4661 (N_4661,N_3662,N_3293);
nor U4662 (N_4662,N_3117,N_3734);
nand U4663 (N_4663,N_3877,N_3892);
nand U4664 (N_4664,N_3901,N_3057);
nand U4665 (N_4665,N_3155,N_3994);
and U4666 (N_4666,N_3395,N_3608);
xnor U4667 (N_4667,N_3962,N_3337);
or U4668 (N_4668,N_3877,N_3830);
xor U4669 (N_4669,N_3386,N_3401);
nand U4670 (N_4670,N_3609,N_3906);
nand U4671 (N_4671,N_3484,N_3724);
and U4672 (N_4672,N_3428,N_3730);
or U4673 (N_4673,N_3219,N_3418);
or U4674 (N_4674,N_3436,N_3293);
xor U4675 (N_4675,N_3116,N_3460);
nand U4676 (N_4676,N_3697,N_3522);
nand U4677 (N_4677,N_3543,N_3385);
nand U4678 (N_4678,N_3759,N_3085);
nor U4679 (N_4679,N_3952,N_3274);
xnor U4680 (N_4680,N_3393,N_3818);
and U4681 (N_4681,N_3415,N_3488);
and U4682 (N_4682,N_3129,N_3706);
or U4683 (N_4683,N_3765,N_3721);
and U4684 (N_4684,N_3793,N_3387);
and U4685 (N_4685,N_3376,N_3367);
xnor U4686 (N_4686,N_3091,N_3373);
or U4687 (N_4687,N_3753,N_3443);
xnor U4688 (N_4688,N_3846,N_3576);
nor U4689 (N_4689,N_3075,N_3146);
and U4690 (N_4690,N_3181,N_3782);
or U4691 (N_4691,N_3472,N_3618);
xor U4692 (N_4692,N_3969,N_3225);
xor U4693 (N_4693,N_3654,N_3413);
nand U4694 (N_4694,N_3441,N_3886);
xor U4695 (N_4695,N_3878,N_3106);
nor U4696 (N_4696,N_3004,N_3508);
or U4697 (N_4697,N_3755,N_3961);
nor U4698 (N_4698,N_3568,N_3416);
nand U4699 (N_4699,N_3309,N_3061);
xnor U4700 (N_4700,N_3958,N_3575);
nand U4701 (N_4701,N_3690,N_3465);
nand U4702 (N_4702,N_3787,N_3166);
or U4703 (N_4703,N_3187,N_3326);
xnor U4704 (N_4704,N_3701,N_3648);
xor U4705 (N_4705,N_3100,N_3501);
xor U4706 (N_4706,N_3923,N_3124);
and U4707 (N_4707,N_3302,N_3814);
and U4708 (N_4708,N_3440,N_3909);
nor U4709 (N_4709,N_3609,N_3061);
or U4710 (N_4710,N_3821,N_3919);
and U4711 (N_4711,N_3902,N_3614);
and U4712 (N_4712,N_3766,N_3676);
or U4713 (N_4713,N_3372,N_3509);
or U4714 (N_4714,N_3383,N_3550);
nand U4715 (N_4715,N_3181,N_3299);
nand U4716 (N_4716,N_3939,N_3785);
and U4717 (N_4717,N_3607,N_3430);
nor U4718 (N_4718,N_3697,N_3994);
and U4719 (N_4719,N_3443,N_3463);
nor U4720 (N_4720,N_3616,N_3032);
xor U4721 (N_4721,N_3094,N_3043);
nand U4722 (N_4722,N_3148,N_3228);
nor U4723 (N_4723,N_3522,N_3673);
nor U4724 (N_4724,N_3529,N_3869);
xnor U4725 (N_4725,N_3176,N_3090);
xnor U4726 (N_4726,N_3958,N_3176);
or U4727 (N_4727,N_3387,N_3010);
nand U4728 (N_4728,N_3616,N_3177);
or U4729 (N_4729,N_3436,N_3068);
and U4730 (N_4730,N_3978,N_3663);
nor U4731 (N_4731,N_3062,N_3592);
nor U4732 (N_4732,N_3411,N_3118);
and U4733 (N_4733,N_3871,N_3375);
or U4734 (N_4734,N_3229,N_3952);
xor U4735 (N_4735,N_3287,N_3042);
or U4736 (N_4736,N_3177,N_3715);
or U4737 (N_4737,N_3072,N_3009);
or U4738 (N_4738,N_3144,N_3749);
and U4739 (N_4739,N_3434,N_3439);
xnor U4740 (N_4740,N_3927,N_3497);
nor U4741 (N_4741,N_3266,N_3709);
or U4742 (N_4742,N_3986,N_3620);
and U4743 (N_4743,N_3401,N_3813);
or U4744 (N_4744,N_3852,N_3099);
nand U4745 (N_4745,N_3487,N_3943);
nor U4746 (N_4746,N_3986,N_3837);
xor U4747 (N_4747,N_3692,N_3834);
nand U4748 (N_4748,N_3979,N_3571);
nor U4749 (N_4749,N_3049,N_3531);
or U4750 (N_4750,N_3989,N_3007);
nand U4751 (N_4751,N_3305,N_3017);
nor U4752 (N_4752,N_3057,N_3941);
nand U4753 (N_4753,N_3153,N_3354);
xor U4754 (N_4754,N_3739,N_3750);
nor U4755 (N_4755,N_3145,N_3882);
nand U4756 (N_4756,N_3076,N_3075);
nand U4757 (N_4757,N_3921,N_3464);
and U4758 (N_4758,N_3085,N_3152);
xnor U4759 (N_4759,N_3429,N_3353);
nor U4760 (N_4760,N_3554,N_3905);
xor U4761 (N_4761,N_3063,N_3087);
or U4762 (N_4762,N_3718,N_3202);
nor U4763 (N_4763,N_3098,N_3324);
xnor U4764 (N_4764,N_3458,N_3399);
xor U4765 (N_4765,N_3466,N_3958);
xnor U4766 (N_4766,N_3060,N_3485);
nand U4767 (N_4767,N_3181,N_3491);
nor U4768 (N_4768,N_3968,N_3630);
nand U4769 (N_4769,N_3450,N_3391);
nor U4770 (N_4770,N_3787,N_3066);
nand U4771 (N_4771,N_3147,N_3601);
nor U4772 (N_4772,N_3374,N_3427);
xor U4773 (N_4773,N_3927,N_3309);
nand U4774 (N_4774,N_3431,N_3723);
nand U4775 (N_4775,N_3218,N_3936);
nor U4776 (N_4776,N_3756,N_3819);
xor U4777 (N_4777,N_3362,N_3404);
and U4778 (N_4778,N_3683,N_3724);
or U4779 (N_4779,N_3837,N_3654);
and U4780 (N_4780,N_3394,N_3222);
nor U4781 (N_4781,N_3032,N_3111);
xnor U4782 (N_4782,N_3810,N_3212);
and U4783 (N_4783,N_3750,N_3509);
xnor U4784 (N_4784,N_3637,N_3950);
and U4785 (N_4785,N_3255,N_3011);
nand U4786 (N_4786,N_3033,N_3645);
and U4787 (N_4787,N_3612,N_3267);
nor U4788 (N_4788,N_3814,N_3098);
nand U4789 (N_4789,N_3943,N_3084);
nor U4790 (N_4790,N_3900,N_3422);
xor U4791 (N_4791,N_3139,N_3485);
nand U4792 (N_4792,N_3499,N_3411);
and U4793 (N_4793,N_3044,N_3205);
and U4794 (N_4794,N_3030,N_3284);
nor U4795 (N_4795,N_3144,N_3960);
and U4796 (N_4796,N_3124,N_3518);
nand U4797 (N_4797,N_3807,N_3049);
nor U4798 (N_4798,N_3595,N_3256);
and U4799 (N_4799,N_3653,N_3104);
and U4800 (N_4800,N_3267,N_3422);
nand U4801 (N_4801,N_3719,N_3631);
and U4802 (N_4802,N_3276,N_3685);
and U4803 (N_4803,N_3892,N_3893);
xnor U4804 (N_4804,N_3134,N_3964);
or U4805 (N_4805,N_3902,N_3576);
nor U4806 (N_4806,N_3067,N_3286);
and U4807 (N_4807,N_3284,N_3956);
xnor U4808 (N_4808,N_3561,N_3588);
or U4809 (N_4809,N_3421,N_3704);
or U4810 (N_4810,N_3376,N_3761);
xor U4811 (N_4811,N_3933,N_3364);
xnor U4812 (N_4812,N_3888,N_3753);
nor U4813 (N_4813,N_3649,N_3439);
and U4814 (N_4814,N_3641,N_3509);
xnor U4815 (N_4815,N_3323,N_3422);
nor U4816 (N_4816,N_3538,N_3752);
nor U4817 (N_4817,N_3378,N_3414);
nand U4818 (N_4818,N_3684,N_3448);
or U4819 (N_4819,N_3160,N_3742);
xor U4820 (N_4820,N_3199,N_3194);
and U4821 (N_4821,N_3013,N_3503);
nor U4822 (N_4822,N_3617,N_3471);
and U4823 (N_4823,N_3489,N_3247);
nand U4824 (N_4824,N_3809,N_3182);
or U4825 (N_4825,N_3634,N_3645);
or U4826 (N_4826,N_3632,N_3373);
nor U4827 (N_4827,N_3346,N_3453);
or U4828 (N_4828,N_3647,N_3776);
xnor U4829 (N_4829,N_3418,N_3712);
or U4830 (N_4830,N_3088,N_3859);
xnor U4831 (N_4831,N_3854,N_3311);
xor U4832 (N_4832,N_3080,N_3113);
nor U4833 (N_4833,N_3840,N_3396);
or U4834 (N_4834,N_3807,N_3544);
or U4835 (N_4835,N_3465,N_3049);
nand U4836 (N_4836,N_3560,N_3846);
and U4837 (N_4837,N_3467,N_3673);
and U4838 (N_4838,N_3537,N_3691);
xnor U4839 (N_4839,N_3147,N_3607);
and U4840 (N_4840,N_3028,N_3334);
nand U4841 (N_4841,N_3797,N_3079);
xor U4842 (N_4842,N_3242,N_3490);
xor U4843 (N_4843,N_3529,N_3854);
nand U4844 (N_4844,N_3837,N_3684);
xor U4845 (N_4845,N_3259,N_3409);
nand U4846 (N_4846,N_3499,N_3562);
xnor U4847 (N_4847,N_3177,N_3856);
nor U4848 (N_4848,N_3210,N_3215);
nor U4849 (N_4849,N_3127,N_3421);
and U4850 (N_4850,N_3678,N_3668);
and U4851 (N_4851,N_3104,N_3033);
or U4852 (N_4852,N_3906,N_3794);
or U4853 (N_4853,N_3913,N_3606);
or U4854 (N_4854,N_3518,N_3889);
or U4855 (N_4855,N_3844,N_3576);
and U4856 (N_4856,N_3008,N_3139);
or U4857 (N_4857,N_3685,N_3768);
and U4858 (N_4858,N_3173,N_3708);
and U4859 (N_4859,N_3743,N_3263);
nand U4860 (N_4860,N_3867,N_3599);
xnor U4861 (N_4861,N_3125,N_3624);
xor U4862 (N_4862,N_3752,N_3113);
or U4863 (N_4863,N_3165,N_3865);
xor U4864 (N_4864,N_3216,N_3282);
or U4865 (N_4865,N_3815,N_3739);
and U4866 (N_4866,N_3899,N_3966);
and U4867 (N_4867,N_3567,N_3368);
nand U4868 (N_4868,N_3304,N_3162);
xor U4869 (N_4869,N_3714,N_3165);
and U4870 (N_4870,N_3501,N_3420);
xnor U4871 (N_4871,N_3142,N_3177);
xor U4872 (N_4872,N_3019,N_3942);
nand U4873 (N_4873,N_3686,N_3272);
and U4874 (N_4874,N_3036,N_3065);
and U4875 (N_4875,N_3834,N_3191);
or U4876 (N_4876,N_3445,N_3984);
nor U4877 (N_4877,N_3806,N_3643);
xor U4878 (N_4878,N_3099,N_3661);
nor U4879 (N_4879,N_3042,N_3792);
nor U4880 (N_4880,N_3807,N_3064);
nand U4881 (N_4881,N_3756,N_3080);
nor U4882 (N_4882,N_3948,N_3123);
nor U4883 (N_4883,N_3156,N_3092);
nor U4884 (N_4884,N_3496,N_3608);
or U4885 (N_4885,N_3508,N_3974);
nor U4886 (N_4886,N_3941,N_3114);
and U4887 (N_4887,N_3978,N_3075);
nand U4888 (N_4888,N_3919,N_3120);
and U4889 (N_4889,N_3557,N_3427);
xor U4890 (N_4890,N_3131,N_3494);
and U4891 (N_4891,N_3612,N_3346);
or U4892 (N_4892,N_3547,N_3754);
xnor U4893 (N_4893,N_3547,N_3823);
and U4894 (N_4894,N_3757,N_3685);
xnor U4895 (N_4895,N_3143,N_3450);
xor U4896 (N_4896,N_3341,N_3112);
nand U4897 (N_4897,N_3889,N_3296);
nand U4898 (N_4898,N_3240,N_3868);
nor U4899 (N_4899,N_3619,N_3693);
and U4900 (N_4900,N_3102,N_3730);
or U4901 (N_4901,N_3168,N_3467);
nand U4902 (N_4902,N_3164,N_3445);
or U4903 (N_4903,N_3006,N_3859);
and U4904 (N_4904,N_3454,N_3255);
nor U4905 (N_4905,N_3395,N_3877);
and U4906 (N_4906,N_3059,N_3428);
nor U4907 (N_4907,N_3036,N_3972);
and U4908 (N_4908,N_3976,N_3862);
or U4909 (N_4909,N_3333,N_3191);
nand U4910 (N_4910,N_3555,N_3203);
and U4911 (N_4911,N_3028,N_3281);
or U4912 (N_4912,N_3710,N_3180);
xor U4913 (N_4913,N_3083,N_3032);
nand U4914 (N_4914,N_3406,N_3239);
or U4915 (N_4915,N_3358,N_3260);
nand U4916 (N_4916,N_3692,N_3299);
nor U4917 (N_4917,N_3210,N_3252);
and U4918 (N_4918,N_3107,N_3201);
xor U4919 (N_4919,N_3940,N_3075);
nor U4920 (N_4920,N_3438,N_3172);
and U4921 (N_4921,N_3748,N_3409);
or U4922 (N_4922,N_3506,N_3785);
nand U4923 (N_4923,N_3584,N_3191);
nand U4924 (N_4924,N_3701,N_3903);
and U4925 (N_4925,N_3110,N_3121);
nor U4926 (N_4926,N_3850,N_3234);
and U4927 (N_4927,N_3658,N_3056);
and U4928 (N_4928,N_3301,N_3568);
nor U4929 (N_4929,N_3995,N_3347);
nand U4930 (N_4930,N_3910,N_3863);
or U4931 (N_4931,N_3523,N_3587);
and U4932 (N_4932,N_3373,N_3297);
or U4933 (N_4933,N_3672,N_3427);
and U4934 (N_4934,N_3722,N_3588);
xnor U4935 (N_4935,N_3521,N_3634);
and U4936 (N_4936,N_3291,N_3620);
nand U4937 (N_4937,N_3432,N_3567);
and U4938 (N_4938,N_3009,N_3451);
xor U4939 (N_4939,N_3629,N_3802);
nor U4940 (N_4940,N_3821,N_3790);
nand U4941 (N_4941,N_3323,N_3132);
nand U4942 (N_4942,N_3283,N_3605);
or U4943 (N_4943,N_3068,N_3128);
xnor U4944 (N_4944,N_3375,N_3213);
xnor U4945 (N_4945,N_3034,N_3226);
and U4946 (N_4946,N_3012,N_3524);
and U4947 (N_4947,N_3777,N_3269);
nor U4948 (N_4948,N_3385,N_3133);
nor U4949 (N_4949,N_3756,N_3570);
xor U4950 (N_4950,N_3363,N_3021);
nand U4951 (N_4951,N_3576,N_3044);
nand U4952 (N_4952,N_3329,N_3113);
and U4953 (N_4953,N_3641,N_3979);
nand U4954 (N_4954,N_3522,N_3019);
or U4955 (N_4955,N_3669,N_3486);
and U4956 (N_4956,N_3309,N_3145);
xnor U4957 (N_4957,N_3141,N_3810);
and U4958 (N_4958,N_3686,N_3925);
and U4959 (N_4959,N_3092,N_3344);
and U4960 (N_4960,N_3546,N_3502);
nand U4961 (N_4961,N_3354,N_3404);
xnor U4962 (N_4962,N_3030,N_3298);
or U4963 (N_4963,N_3201,N_3389);
nor U4964 (N_4964,N_3017,N_3672);
or U4965 (N_4965,N_3229,N_3651);
nand U4966 (N_4966,N_3776,N_3746);
nand U4967 (N_4967,N_3309,N_3605);
xor U4968 (N_4968,N_3648,N_3352);
nor U4969 (N_4969,N_3305,N_3449);
xor U4970 (N_4970,N_3027,N_3376);
or U4971 (N_4971,N_3860,N_3122);
nand U4972 (N_4972,N_3581,N_3325);
nor U4973 (N_4973,N_3737,N_3674);
xor U4974 (N_4974,N_3065,N_3395);
or U4975 (N_4975,N_3969,N_3491);
xor U4976 (N_4976,N_3928,N_3757);
nand U4977 (N_4977,N_3512,N_3957);
xor U4978 (N_4978,N_3408,N_3082);
xnor U4979 (N_4979,N_3333,N_3061);
and U4980 (N_4980,N_3542,N_3705);
and U4981 (N_4981,N_3107,N_3920);
xnor U4982 (N_4982,N_3863,N_3582);
or U4983 (N_4983,N_3000,N_3492);
xnor U4984 (N_4984,N_3161,N_3877);
nand U4985 (N_4985,N_3643,N_3891);
and U4986 (N_4986,N_3603,N_3470);
or U4987 (N_4987,N_3187,N_3541);
nor U4988 (N_4988,N_3525,N_3510);
and U4989 (N_4989,N_3501,N_3494);
or U4990 (N_4990,N_3597,N_3662);
or U4991 (N_4991,N_3543,N_3112);
or U4992 (N_4992,N_3066,N_3945);
or U4993 (N_4993,N_3205,N_3896);
and U4994 (N_4994,N_3403,N_3875);
or U4995 (N_4995,N_3132,N_3530);
or U4996 (N_4996,N_3813,N_3825);
and U4997 (N_4997,N_3719,N_3253);
and U4998 (N_4998,N_3517,N_3320);
or U4999 (N_4999,N_3070,N_3045);
or U5000 (N_5000,N_4960,N_4972);
nor U5001 (N_5001,N_4649,N_4629);
or U5002 (N_5002,N_4591,N_4970);
or U5003 (N_5003,N_4148,N_4560);
nor U5004 (N_5004,N_4146,N_4570);
and U5005 (N_5005,N_4187,N_4584);
or U5006 (N_5006,N_4879,N_4380);
nor U5007 (N_5007,N_4093,N_4160);
nand U5008 (N_5008,N_4742,N_4012);
nor U5009 (N_5009,N_4661,N_4441);
nor U5010 (N_5010,N_4278,N_4201);
nor U5011 (N_5011,N_4912,N_4887);
xnor U5012 (N_5012,N_4299,N_4308);
nor U5013 (N_5013,N_4287,N_4491);
nor U5014 (N_5014,N_4151,N_4843);
or U5015 (N_5015,N_4736,N_4870);
xor U5016 (N_5016,N_4783,N_4452);
nand U5017 (N_5017,N_4758,N_4685);
xnor U5018 (N_5018,N_4227,N_4821);
or U5019 (N_5019,N_4237,N_4643);
nor U5020 (N_5020,N_4066,N_4167);
nor U5021 (N_5021,N_4175,N_4875);
nor U5022 (N_5022,N_4181,N_4330);
or U5023 (N_5023,N_4371,N_4717);
and U5024 (N_5024,N_4317,N_4703);
or U5025 (N_5025,N_4674,N_4247);
or U5026 (N_5026,N_4092,N_4898);
and U5027 (N_5027,N_4041,N_4057);
nor U5028 (N_5028,N_4817,N_4506);
nor U5029 (N_5029,N_4851,N_4046);
or U5030 (N_5030,N_4716,N_4630);
or U5031 (N_5031,N_4611,N_4588);
or U5032 (N_5032,N_4221,N_4274);
nor U5033 (N_5033,N_4079,N_4313);
nor U5034 (N_5034,N_4054,N_4044);
nor U5035 (N_5035,N_4375,N_4271);
or U5036 (N_5036,N_4966,N_4383);
xor U5037 (N_5037,N_4862,N_4035);
or U5038 (N_5038,N_4533,N_4848);
xnor U5039 (N_5039,N_4502,N_4082);
nor U5040 (N_5040,N_4714,N_4106);
or U5041 (N_5041,N_4463,N_4314);
nor U5042 (N_5042,N_4615,N_4521);
xor U5043 (N_5043,N_4026,N_4178);
and U5044 (N_5044,N_4216,N_4280);
and U5045 (N_5045,N_4766,N_4258);
nand U5046 (N_5046,N_4888,N_4297);
xnor U5047 (N_5047,N_4285,N_4599);
and U5048 (N_5048,N_4977,N_4908);
nor U5049 (N_5049,N_4042,N_4222);
nand U5050 (N_5050,N_4507,N_4085);
nand U5051 (N_5051,N_4782,N_4874);
nand U5052 (N_5052,N_4865,N_4911);
and U5053 (N_5053,N_4562,N_4087);
and U5054 (N_5054,N_4332,N_4168);
or U5055 (N_5055,N_4186,N_4976);
xor U5056 (N_5056,N_4128,N_4542);
nand U5057 (N_5057,N_4559,N_4544);
nand U5058 (N_5058,N_4637,N_4126);
nor U5059 (N_5059,N_4534,N_4607);
and U5060 (N_5060,N_4586,N_4640);
and U5061 (N_5061,N_4368,N_4407);
or U5062 (N_5062,N_4645,N_4210);
nor U5063 (N_5063,N_4658,N_4757);
nand U5064 (N_5064,N_4249,N_4922);
xor U5065 (N_5065,N_4923,N_4635);
and U5066 (N_5066,N_4055,N_4132);
xor U5067 (N_5067,N_4381,N_4997);
xnor U5068 (N_5068,N_4244,N_4239);
xnor U5069 (N_5069,N_4465,N_4699);
and U5070 (N_5070,N_4854,N_4856);
and U5071 (N_5071,N_4430,N_4633);
or U5072 (N_5072,N_4924,N_4372);
or U5073 (N_5073,N_4162,N_4188);
or U5074 (N_5074,N_4142,N_4283);
nor U5075 (N_5075,N_4303,N_4989);
xnor U5076 (N_5076,N_4695,N_4822);
and U5077 (N_5077,N_4844,N_4479);
or U5078 (N_5078,N_4690,N_4827);
xor U5079 (N_5079,N_4362,N_4841);
and U5080 (N_5080,N_4784,N_4715);
nand U5081 (N_5081,N_4760,N_4726);
and U5082 (N_5082,N_4946,N_4021);
nor U5083 (N_5083,N_4165,N_4941);
or U5084 (N_5084,N_4067,N_4415);
and U5085 (N_5085,N_4064,N_4094);
or U5086 (N_5086,N_4706,N_4652);
or U5087 (N_5087,N_4032,N_4583);
or U5088 (N_5088,N_4979,N_4031);
and U5089 (N_5089,N_4047,N_4945);
xor U5090 (N_5090,N_4537,N_4644);
or U5091 (N_5091,N_4260,N_4340);
or U5092 (N_5092,N_4449,N_4212);
xnor U5093 (N_5093,N_4219,N_4401);
nor U5094 (N_5094,N_4425,N_4356);
nor U5095 (N_5095,N_4855,N_4872);
nand U5096 (N_5096,N_4137,N_4984);
or U5097 (N_5097,N_4820,N_4708);
xor U5098 (N_5098,N_4166,N_4127);
and U5099 (N_5099,N_4907,N_4058);
or U5100 (N_5100,N_4687,N_4824);
or U5101 (N_5101,N_4701,N_4061);
and U5102 (N_5102,N_4204,N_4433);
nor U5103 (N_5103,N_4207,N_4180);
and U5104 (N_5104,N_4097,N_4868);
nor U5105 (N_5105,N_4641,N_4427);
xnor U5106 (N_5106,N_4962,N_4574);
xnor U5107 (N_5107,N_4692,N_4622);
and U5108 (N_5108,N_4581,N_4919);
nand U5109 (N_5109,N_4494,N_4030);
nor U5110 (N_5110,N_4947,N_4014);
or U5111 (N_5111,N_4727,N_4531);
or U5112 (N_5112,N_4763,N_4466);
and U5113 (N_5113,N_4256,N_4255);
nand U5114 (N_5114,N_4655,N_4288);
nand U5115 (N_5115,N_4639,N_4359);
or U5116 (N_5116,N_4298,N_4254);
nor U5117 (N_5117,N_4492,N_4602);
xnor U5118 (N_5118,N_4871,N_4445);
nor U5119 (N_5119,N_4442,N_4469);
nand U5120 (N_5120,N_4199,N_4547);
or U5121 (N_5121,N_4027,N_4744);
and U5122 (N_5122,N_4546,N_4113);
and U5123 (N_5123,N_4322,N_4265);
or U5124 (N_5124,N_4628,N_4704);
nand U5125 (N_5125,N_4662,N_4018);
nand U5126 (N_5126,N_4203,N_4548);
or U5127 (N_5127,N_4225,N_4853);
and U5128 (N_5128,N_4440,N_4954);
and U5129 (N_5129,N_4847,N_4631);
nor U5130 (N_5130,N_4852,N_4096);
xnor U5131 (N_5131,N_4024,N_4198);
nor U5132 (N_5132,N_4156,N_4053);
or U5133 (N_5133,N_4831,N_4567);
nor U5134 (N_5134,N_4917,N_4536);
and U5135 (N_5135,N_4719,N_4001);
and U5136 (N_5136,N_4095,N_4845);
xor U5137 (N_5137,N_4409,N_4850);
or U5138 (N_5138,N_4416,N_4417);
and U5139 (N_5139,N_4377,N_4858);
and U5140 (N_5140,N_4335,N_4691);
nor U5141 (N_5141,N_4517,N_4769);
or U5142 (N_5142,N_4310,N_4264);
xor U5143 (N_5143,N_4139,N_4765);
and U5144 (N_5144,N_4798,N_4569);
and U5145 (N_5145,N_4551,N_4355);
or U5146 (N_5146,N_4712,N_4458);
and U5147 (N_5147,N_4140,N_4177);
and U5148 (N_5148,N_4485,N_4921);
or U5149 (N_5149,N_4208,N_4503);
xnor U5150 (N_5150,N_4321,N_4125);
and U5151 (N_5151,N_4394,N_4194);
or U5152 (N_5152,N_4801,N_4686);
and U5153 (N_5153,N_4185,N_4900);
xnor U5154 (N_5154,N_4353,N_4748);
and U5155 (N_5155,N_4325,N_4245);
xor U5156 (N_5156,N_4124,N_4455);
nand U5157 (N_5157,N_4894,N_4776);
or U5158 (N_5158,N_4789,N_4881);
nand U5159 (N_5159,N_4391,N_4205);
nand U5160 (N_5160,N_4364,N_4558);
xor U5161 (N_5161,N_4050,N_4473);
and U5162 (N_5162,N_4561,N_4345);
xor U5163 (N_5163,N_4971,N_4730);
and U5164 (N_5164,N_4762,N_4481);
nor U5165 (N_5165,N_4963,N_4745);
nor U5166 (N_5166,N_4550,N_4935);
and U5167 (N_5167,N_4286,N_4090);
xor U5168 (N_5168,N_4513,N_4500);
and U5169 (N_5169,N_4796,N_4978);
nand U5170 (N_5170,N_4694,N_4400);
and U5171 (N_5171,N_4150,N_4184);
and U5172 (N_5172,N_4749,N_4179);
and U5173 (N_5173,N_4804,N_4505);
xnor U5174 (N_5174,N_4992,N_4767);
nand U5175 (N_5175,N_4472,N_4882);
or U5176 (N_5176,N_4434,N_4200);
xnor U5177 (N_5177,N_4435,N_4343);
nand U5178 (N_5178,N_4575,N_4829);
xor U5179 (N_5179,N_4968,N_4277);
or U5180 (N_5180,N_4683,N_4610);
nand U5181 (N_5181,N_4376,N_4275);
nor U5182 (N_5182,N_4261,N_4627);
nor U5183 (N_5183,N_4483,N_4008);
and U5184 (N_5184,N_4873,N_4306);
nor U5185 (N_5185,N_4259,N_4597);
nor U5186 (N_5186,N_4251,N_4422);
nor U5187 (N_5187,N_4587,N_4555);
nor U5188 (N_5188,N_4309,N_4461);
xor U5189 (N_5189,N_4689,N_4220);
xnor U5190 (N_5190,N_4944,N_4170);
and U5191 (N_5191,N_4338,N_4609);
or U5192 (N_5192,N_4752,N_4451);
or U5193 (N_5193,N_4423,N_4272);
nand U5194 (N_5194,N_4999,N_4290);
xor U5195 (N_5195,N_4818,N_4616);
or U5196 (N_5196,N_4604,N_4793);
xor U5197 (N_5197,N_4301,N_4957);
and U5198 (N_5198,N_4154,N_4467);
or U5199 (N_5199,N_4480,N_4016);
nor U5200 (N_5200,N_4880,N_4190);
xor U5201 (N_5201,N_4387,N_4747);
nand U5202 (N_5202,N_4861,N_4475);
xor U5203 (N_5203,N_4228,N_4369);
or U5204 (N_5204,N_4753,N_4367);
nand U5205 (N_5205,N_4341,N_4048);
or U5206 (N_5206,N_4476,N_4993);
nand U5207 (N_5207,N_4756,N_4918);
or U5208 (N_5208,N_4007,N_4939);
nand U5209 (N_5209,N_4171,N_4524);
xor U5210 (N_5210,N_4903,N_4135);
nand U5211 (N_5211,N_4884,N_4081);
nor U5212 (N_5212,N_4361,N_4642);
nor U5213 (N_5213,N_4083,N_4432);
xnor U5214 (N_5214,N_4660,N_4266);
nand U5215 (N_5215,N_4996,N_4292);
or U5216 (N_5216,N_4777,N_4234);
and U5217 (N_5217,N_4846,N_4196);
nor U5218 (N_5218,N_4665,N_4075);
nor U5219 (N_5219,N_4837,N_4395);
xnor U5220 (N_5220,N_4823,N_4621);
nand U5221 (N_5221,N_4833,N_4931);
xor U5222 (N_5222,N_4589,N_4020);
xor U5223 (N_5223,N_4183,N_4696);
nand U5224 (N_5224,N_4519,N_4810);
nand U5225 (N_5225,N_4250,N_4498);
xor U5226 (N_5226,N_4596,N_4226);
nor U5227 (N_5227,N_4318,N_4352);
nand U5228 (N_5228,N_4213,N_4350);
nor U5229 (N_5229,N_4487,N_4663);
nor U5230 (N_5230,N_4986,N_4102);
and U5231 (N_5231,N_4114,N_4606);
nand U5232 (N_5232,N_4474,N_4164);
xnor U5233 (N_5233,N_4626,N_4173);
nand U5234 (N_5234,N_4991,N_4059);
xnor U5235 (N_5235,N_4086,N_4681);
xor U5236 (N_5236,N_4541,N_4029);
xor U5237 (N_5237,N_4988,N_4664);
nor U5238 (N_5238,N_4439,N_4932);
xor U5239 (N_5239,N_4682,N_4974);
xnor U5240 (N_5240,N_4952,N_4578);
or U5241 (N_5241,N_4496,N_4182);
or U5242 (N_5242,N_4077,N_4365);
or U5243 (N_5243,N_4866,N_4484);
or U5244 (N_5244,N_4169,N_4650);
nand U5245 (N_5245,N_4806,N_4454);
xor U5246 (N_5246,N_4107,N_4323);
or U5247 (N_5247,N_4478,N_4462);
and U5248 (N_5248,N_4373,N_4477);
or U5249 (N_5249,N_4192,N_4659);
or U5250 (N_5250,N_4925,N_4514);
or U5251 (N_5251,N_4098,N_4358);
xor U5252 (N_5252,N_4828,N_4724);
and U5253 (N_5253,N_4869,N_4241);
and U5254 (N_5254,N_4790,N_4965);
nor U5255 (N_5255,N_4421,N_4316);
xnor U5256 (N_5256,N_4950,N_4403);
or U5257 (N_5257,N_4612,N_4063);
nor U5258 (N_5258,N_4110,N_4311);
nor U5259 (N_5259,N_4839,N_4815);
nand U5260 (N_5260,N_4799,N_4211);
or U5261 (N_5261,N_4928,N_4520);
xor U5262 (N_5262,N_4370,N_4218);
nand U5263 (N_5263,N_4980,N_4257);
xnor U5264 (N_5264,N_4867,N_4565);
nor U5265 (N_5265,N_4552,N_4711);
nand U5266 (N_5266,N_4545,N_4593);
nand U5267 (N_5267,N_4910,N_4038);
xor U5268 (N_5268,N_4624,N_4885);
xor U5269 (N_5269,N_4620,N_4675);
xor U5270 (N_5270,N_4224,N_4319);
or U5271 (N_5271,N_4223,N_4450);
nor U5272 (N_5272,N_4859,N_4797);
nand U5273 (N_5273,N_4671,N_4295);
xnor U5274 (N_5274,N_4312,N_4914);
nor U5275 (N_5275,N_4420,N_4525);
and U5276 (N_5276,N_4805,N_4739);
or U5277 (N_5277,N_4159,N_4133);
and U5278 (N_5278,N_4327,N_4594);
nor U5279 (N_5279,N_4131,N_4120);
nor U5280 (N_5280,N_4056,N_4613);
nor U5281 (N_5281,N_4155,N_4735);
xnor U5282 (N_5282,N_4540,N_4397);
nor U5283 (N_5283,N_4893,N_4291);
xnor U5284 (N_5284,N_4108,N_4229);
and U5285 (N_5285,N_4405,N_4418);
xor U5286 (N_5286,N_4938,N_4625);
and U5287 (N_5287,N_4100,N_4331);
nor U5288 (N_5288,N_4539,N_4927);
xnor U5289 (N_5289,N_4006,N_4145);
nor U5290 (N_5290,N_4413,N_4959);
and U5291 (N_5291,N_4143,N_4411);
or U5292 (N_5292,N_4337,N_4740);
and U5293 (N_5293,N_4289,N_4037);
and U5294 (N_5294,N_4543,N_4608);
or U5295 (N_5295,N_4398,N_4281);
nor U5296 (N_5296,N_4838,N_4571);
or U5297 (N_5297,N_4897,N_4015);
nor U5298 (N_5298,N_4489,N_4961);
and U5299 (N_5299,N_4117,N_4532);
or U5300 (N_5300,N_4022,N_4080);
nor U5301 (N_5301,N_4951,N_4497);
or U5302 (N_5302,N_4495,N_4527);
xor U5303 (N_5303,N_4028,N_4705);
nand U5304 (N_5304,N_4443,N_4779);
nand U5305 (N_5305,N_4891,N_4564);
or U5306 (N_5306,N_4825,N_4122);
or U5307 (N_5307,N_4771,N_4130);
nand U5308 (N_5308,N_4728,N_4913);
or U5309 (N_5309,N_4942,N_4328);
or U5310 (N_5310,N_4429,N_4074);
or U5311 (N_5311,N_4348,N_4388);
and U5312 (N_5312,N_4005,N_4501);
or U5313 (N_5313,N_4515,N_4812);
or U5314 (N_5314,N_4902,N_4538);
xnor U5315 (N_5315,N_4091,N_4654);
or U5316 (N_5316,N_4830,N_4504);
or U5317 (N_5317,N_4590,N_4268);
nand U5318 (N_5318,N_4656,N_4385);
or U5319 (N_5319,N_4457,N_4153);
nand U5320 (N_5320,N_4262,N_4379);
and U5321 (N_5321,N_4955,N_4916);
and U5322 (N_5322,N_4857,N_4573);
or U5323 (N_5323,N_4197,N_4598);
nor U5324 (N_5324,N_4152,N_4176);
nor U5325 (N_5325,N_4780,N_4638);
xor U5326 (N_5326,N_4231,N_4720);
nor U5327 (N_5327,N_4101,N_4576);
xnor U5328 (N_5328,N_4787,N_4040);
xnor U5329 (N_5329,N_4568,N_4103);
xnor U5330 (N_5330,N_4553,N_4099);
or U5331 (N_5331,N_4676,N_4940);
nor U5332 (N_5332,N_4878,N_4267);
nor U5333 (N_5333,N_4956,N_4953);
xnor U5334 (N_5334,N_4428,N_4305);
nand U5335 (N_5335,N_4781,N_4069);
or U5336 (N_5336,N_4808,N_4710);
xor U5337 (N_5337,N_4049,N_4794);
nor U5338 (N_5338,N_4144,N_4967);
xnor U5339 (N_5339,N_4279,N_4490);
nor U5340 (N_5340,N_4349,N_4722);
nand U5341 (N_5341,N_4088,N_4835);
nand U5342 (N_5342,N_4618,N_4214);
nor U5343 (N_5343,N_4723,N_4800);
xor U5344 (N_5344,N_4890,N_4294);
or U5345 (N_5345,N_4304,N_4149);
and U5346 (N_5346,N_4161,N_4713);
and U5347 (N_5347,N_4667,N_4464);
and U5348 (N_5348,N_4382,N_4526);
xnor U5349 (N_5349,N_4410,N_4775);
or U5350 (N_5350,N_4601,N_4399);
nand U5351 (N_5351,N_4393,N_4592);
or U5352 (N_5352,N_4003,N_4406);
and U5353 (N_5353,N_4339,N_4195);
nor U5354 (N_5354,N_4121,N_4981);
and U5355 (N_5355,N_4684,N_4582);
nor U5356 (N_5356,N_4975,N_4414);
xnor U5357 (N_5357,N_4307,N_4269);
xnor U5358 (N_5358,N_4013,N_4347);
or U5359 (N_5359,N_4809,N_4482);
xor U5360 (N_5360,N_4926,N_4886);
nor U5361 (N_5361,N_4774,N_4819);
and U5362 (N_5362,N_4530,N_4202);
nand U5363 (N_5363,N_4426,N_4813);
nand U5364 (N_5364,N_4045,N_4761);
or U5365 (N_5365,N_4437,N_4468);
or U5366 (N_5366,N_4302,N_4746);
nor U5367 (N_5367,N_4390,N_4764);
nor U5368 (N_5368,N_4189,N_4614);
and U5369 (N_5369,N_4019,N_4802);
or U5370 (N_5370,N_4404,N_4732);
nand U5371 (N_5371,N_4253,N_4109);
xnor U5372 (N_5372,N_4904,N_4235);
or U5373 (N_5373,N_4901,N_4721);
xor U5374 (N_5374,N_4209,N_4930);
xnor U5375 (N_5375,N_4899,N_4315);
or U5376 (N_5376,N_4002,N_4915);
nor U5377 (N_5377,N_4105,N_4709);
nand U5378 (N_5378,N_4158,N_4273);
xnor U5379 (N_5379,N_4698,N_4688);
or U5380 (N_5380,N_4572,N_4025);
and U5381 (N_5381,N_4116,N_4985);
xor U5382 (N_5382,N_4792,N_4448);
or U5383 (N_5383,N_4697,N_4248);
or U5384 (N_5384,N_4934,N_4043);
nor U5385 (N_5385,N_4329,N_4943);
nor U5386 (N_5386,N_4786,N_4342);
or U5387 (N_5387,N_4788,N_4778);
nand U5388 (N_5388,N_4010,N_4670);
xnor U5389 (N_5389,N_4004,N_4354);
or U5390 (N_5390,N_4326,N_4270);
nor U5391 (N_5391,N_4104,N_4488);
and U5392 (N_5392,N_4470,N_4679);
nand U5393 (N_5393,N_4785,N_4499);
xnor U5394 (N_5394,N_4123,N_4791);
nand U5395 (N_5395,N_4636,N_4111);
xnor U5396 (N_5396,N_4840,N_4734);
nor U5397 (N_5397,N_4076,N_4282);
nand U5398 (N_5398,N_4528,N_4990);
nand U5399 (N_5399,N_4617,N_4363);
and U5400 (N_5400,N_4755,N_4284);
and U5401 (N_5401,N_4246,N_4754);
nand U5402 (N_5402,N_4619,N_4486);
and U5403 (N_5403,N_4510,N_4346);
and U5404 (N_5404,N_4232,N_4535);
nand U5405 (N_5405,N_4680,N_4073);
or U5406 (N_5406,N_4446,N_4129);
nor U5407 (N_5407,N_4230,N_4163);
xnor U5408 (N_5408,N_4816,N_4238);
xor U5409 (N_5409,N_4549,N_4896);
nor U5410 (N_5410,N_4193,N_4141);
or U5411 (N_5411,N_4933,N_4459);
nand U5412 (N_5412,N_4033,N_4453);
and U5413 (N_5413,N_4677,N_4134);
xnor U5414 (N_5414,N_4419,N_4444);
or U5415 (N_5415,N_4668,N_4000);
and U5416 (N_5416,N_4929,N_4657);
and U5417 (N_5417,N_4072,N_4036);
nor U5418 (N_5418,N_4052,N_4344);
nand U5419 (N_5419,N_4595,N_4741);
xor U5420 (N_5420,N_4849,N_4836);
or U5421 (N_5421,N_4065,N_4673);
xor U5422 (N_5422,N_4949,N_4580);
nor U5423 (N_5423,N_4973,N_4995);
nand U5424 (N_5424,N_4707,N_4554);
nand U5425 (N_5425,N_4136,N_4729);
xnor U5426 (N_5426,N_4773,N_4743);
and U5427 (N_5427,N_4119,N_4039);
nand U5428 (N_5428,N_4623,N_4366);
nor U5429 (N_5429,N_4895,N_4378);
nor U5430 (N_5430,N_4892,N_4060);
nor U5431 (N_5431,N_4669,N_4795);
nor U5432 (N_5432,N_4115,N_4215);
nor U5433 (N_5433,N_4905,N_4509);
or U5434 (N_5434,N_4522,N_4603);
nor U5435 (N_5435,N_4772,N_4860);
or U5436 (N_5436,N_4412,N_4252);
nand U5437 (N_5437,N_4523,N_4678);
nor U5438 (N_5438,N_4217,N_4078);
nand U5439 (N_5439,N_4969,N_4982);
or U5440 (N_5440,N_4994,N_4436);
nor U5441 (N_5441,N_4814,N_4750);
and U5442 (N_5442,N_4936,N_4557);
nor U5443 (N_5443,N_4389,N_4518);
nand U5444 (N_5444,N_4408,N_4998);
xnor U5445 (N_5445,N_4357,N_4648);
xor U5446 (N_5446,N_4438,N_4842);
nor U5447 (N_5447,N_4089,N_4700);
nor U5448 (N_5448,N_4512,N_4242);
nor U5449 (N_5449,N_4062,N_4243);
xor U5450 (N_5450,N_4605,N_4493);
and U5451 (N_5451,N_4646,N_4579);
nand U5452 (N_5452,N_4738,N_4651);
xor U5453 (N_5453,N_4864,N_4112);
nand U5454 (N_5454,N_4334,N_4811);
xor U5455 (N_5455,N_4384,N_4566);
nor U5456 (N_5456,N_4863,N_4751);
and U5457 (N_5457,N_4529,N_4632);
and U5458 (N_5458,N_4834,N_4718);
nand U5459 (N_5459,N_4296,N_4424);
and U5460 (N_5460,N_4877,N_4832);
xnor U5461 (N_5461,N_4351,N_4563);
and U5462 (N_5462,N_4071,N_4770);
or U5463 (N_5463,N_4937,N_4174);
nor U5464 (N_5464,N_4206,N_4759);
nand U5465 (N_5465,N_4768,N_4889);
nor U5466 (N_5466,N_4402,N_4147);
nor U5467 (N_5467,N_4964,N_4647);
or U5468 (N_5468,N_4023,N_4263);
and U5469 (N_5469,N_4807,N_4826);
xnor U5470 (N_5470,N_4693,N_4702);
nand U5471 (N_5471,N_4011,N_4240);
or U5472 (N_5472,N_4374,N_4883);
nand U5473 (N_5473,N_4051,N_4191);
xnor U5474 (N_5474,N_4233,N_4293);
and U5475 (N_5475,N_4084,N_4987);
or U5476 (N_5476,N_4672,N_4138);
nand U5477 (N_5477,N_4600,N_4447);
and U5478 (N_5478,N_4118,N_4017);
xor U5479 (N_5479,N_4431,N_4511);
or U5480 (N_5480,N_4392,N_4360);
and U5481 (N_5481,N_4471,N_4958);
xor U5482 (N_5482,N_4034,N_4333);
xnor U5483 (N_5483,N_4737,N_4324);
nand U5484 (N_5484,N_4920,N_4983);
nor U5485 (N_5485,N_4909,N_4336);
and U5486 (N_5486,N_4666,N_4577);
or U5487 (N_5487,N_4172,N_4725);
nand U5488 (N_5488,N_4300,N_4906);
or U5489 (N_5489,N_4731,N_4236);
and U5490 (N_5490,N_4396,N_4634);
nand U5491 (N_5491,N_4386,N_4460);
and U5492 (N_5492,N_4320,N_4070);
and U5493 (N_5493,N_4516,N_4508);
nor U5494 (N_5494,N_4948,N_4157);
or U5495 (N_5495,N_4876,N_4276);
nand U5496 (N_5496,N_4733,N_4803);
nor U5497 (N_5497,N_4585,N_4653);
and U5498 (N_5498,N_4556,N_4456);
or U5499 (N_5499,N_4009,N_4068);
or U5500 (N_5500,N_4722,N_4783);
nand U5501 (N_5501,N_4510,N_4345);
and U5502 (N_5502,N_4143,N_4691);
xor U5503 (N_5503,N_4263,N_4111);
xor U5504 (N_5504,N_4763,N_4963);
or U5505 (N_5505,N_4703,N_4605);
or U5506 (N_5506,N_4008,N_4050);
xnor U5507 (N_5507,N_4906,N_4576);
and U5508 (N_5508,N_4568,N_4693);
or U5509 (N_5509,N_4624,N_4730);
nor U5510 (N_5510,N_4187,N_4976);
xnor U5511 (N_5511,N_4830,N_4997);
or U5512 (N_5512,N_4122,N_4213);
xor U5513 (N_5513,N_4601,N_4468);
and U5514 (N_5514,N_4779,N_4805);
and U5515 (N_5515,N_4103,N_4944);
or U5516 (N_5516,N_4728,N_4496);
nand U5517 (N_5517,N_4244,N_4770);
and U5518 (N_5518,N_4764,N_4556);
nor U5519 (N_5519,N_4415,N_4235);
or U5520 (N_5520,N_4847,N_4935);
nor U5521 (N_5521,N_4059,N_4217);
or U5522 (N_5522,N_4127,N_4198);
or U5523 (N_5523,N_4893,N_4946);
nor U5524 (N_5524,N_4489,N_4030);
nand U5525 (N_5525,N_4366,N_4634);
or U5526 (N_5526,N_4067,N_4184);
nor U5527 (N_5527,N_4960,N_4325);
nand U5528 (N_5528,N_4244,N_4074);
nor U5529 (N_5529,N_4828,N_4594);
and U5530 (N_5530,N_4622,N_4319);
or U5531 (N_5531,N_4184,N_4530);
or U5532 (N_5532,N_4429,N_4810);
or U5533 (N_5533,N_4771,N_4358);
and U5534 (N_5534,N_4934,N_4130);
or U5535 (N_5535,N_4794,N_4828);
nor U5536 (N_5536,N_4521,N_4486);
and U5537 (N_5537,N_4971,N_4934);
nor U5538 (N_5538,N_4410,N_4651);
and U5539 (N_5539,N_4406,N_4079);
and U5540 (N_5540,N_4503,N_4808);
and U5541 (N_5541,N_4651,N_4320);
and U5542 (N_5542,N_4142,N_4655);
xnor U5543 (N_5543,N_4325,N_4726);
nor U5544 (N_5544,N_4231,N_4520);
nor U5545 (N_5545,N_4640,N_4450);
xor U5546 (N_5546,N_4374,N_4587);
nor U5547 (N_5547,N_4744,N_4650);
nand U5548 (N_5548,N_4574,N_4028);
nand U5549 (N_5549,N_4923,N_4175);
and U5550 (N_5550,N_4174,N_4297);
or U5551 (N_5551,N_4356,N_4517);
nand U5552 (N_5552,N_4393,N_4652);
nand U5553 (N_5553,N_4191,N_4323);
and U5554 (N_5554,N_4617,N_4058);
or U5555 (N_5555,N_4479,N_4551);
nor U5556 (N_5556,N_4530,N_4611);
xnor U5557 (N_5557,N_4808,N_4436);
nor U5558 (N_5558,N_4553,N_4698);
nand U5559 (N_5559,N_4867,N_4251);
nand U5560 (N_5560,N_4217,N_4377);
and U5561 (N_5561,N_4315,N_4981);
nor U5562 (N_5562,N_4749,N_4058);
xnor U5563 (N_5563,N_4523,N_4170);
or U5564 (N_5564,N_4880,N_4683);
nand U5565 (N_5565,N_4957,N_4755);
nor U5566 (N_5566,N_4073,N_4561);
xor U5567 (N_5567,N_4376,N_4434);
and U5568 (N_5568,N_4798,N_4333);
nor U5569 (N_5569,N_4668,N_4958);
nand U5570 (N_5570,N_4255,N_4826);
nor U5571 (N_5571,N_4387,N_4720);
nor U5572 (N_5572,N_4067,N_4267);
and U5573 (N_5573,N_4861,N_4125);
and U5574 (N_5574,N_4610,N_4432);
or U5575 (N_5575,N_4456,N_4987);
xnor U5576 (N_5576,N_4506,N_4350);
nand U5577 (N_5577,N_4834,N_4242);
and U5578 (N_5578,N_4518,N_4795);
and U5579 (N_5579,N_4825,N_4017);
xnor U5580 (N_5580,N_4065,N_4180);
xor U5581 (N_5581,N_4256,N_4988);
or U5582 (N_5582,N_4513,N_4787);
nand U5583 (N_5583,N_4809,N_4290);
nor U5584 (N_5584,N_4652,N_4005);
and U5585 (N_5585,N_4245,N_4914);
xnor U5586 (N_5586,N_4412,N_4486);
nor U5587 (N_5587,N_4386,N_4547);
nor U5588 (N_5588,N_4528,N_4275);
nor U5589 (N_5589,N_4134,N_4528);
xor U5590 (N_5590,N_4054,N_4507);
and U5591 (N_5591,N_4163,N_4419);
and U5592 (N_5592,N_4454,N_4684);
or U5593 (N_5593,N_4747,N_4489);
nor U5594 (N_5594,N_4123,N_4911);
nand U5595 (N_5595,N_4323,N_4438);
and U5596 (N_5596,N_4799,N_4958);
xor U5597 (N_5597,N_4131,N_4710);
nand U5598 (N_5598,N_4680,N_4383);
or U5599 (N_5599,N_4442,N_4386);
nand U5600 (N_5600,N_4225,N_4944);
and U5601 (N_5601,N_4061,N_4940);
nand U5602 (N_5602,N_4119,N_4019);
xor U5603 (N_5603,N_4569,N_4912);
and U5604 (N_5604,N_4209,N_4150);
and U5605 (N_5605,N_4057,N_4383);
or U5606 (N_5606,N_4583,N_4177);
nor U5607 (N_5607,N_4926,N_4983);
xor U5608 (N_5608,N_4006,N_4949);
or U5609 (N_5609,N_4376,N_4653);
nor U5610 (N_5610,N_4563,N_4666);
xnor U5611 (N_5611,N_4359,N_4066);
xnor U5612 (N_5612,N_4964,N_4642);
nor U5613 (N_5613,N_4360,N_4424);
nand U5614 (N_5614,N_4936,N_4010);
and U5615 (N_5615,N_4649,N_4651);
nand U5616 (N_5616,N_4763,N_4026);
xnor U5617 (N_5617,N_4901,N_4498);
and U5618 (N_5618,N_4616,N_4413);
and U5619 (N_5619,N_4782,N_4139);
or U5620 (N_5620,N_4197,N_4472);
nor U5621 (N_5621,N_4717,N_4664);
nor U5622 (N_5622,N_4504,N_4725);
xnor U5623 (N_5623,N_4132,N_4124);
xor U5624 (N_5624,N_4538,N_4665);
xor U5625 (N_5625,N_4887,N_4400);
xnor U5626 (N_5626,N_4574,N_4377);
nor U5627 (N_5627,N_4335,N_4080);
or U5628 (N_5628,N_4232,N_4643);
or U5629 (N_5629,N_4131,N_4123);
or U5630 (N_5630,N_4085,N_4683);
or U5631 (N_5631,N_4707,N_4279);
nand U5632 (N_5632,N_4879,N_4342);
xor U5633 (N_5633,N_4376,N_4352);
nor U5634 (N_5634,N_4587,N_4561);
nor U5635 (N_5635,N_4543,N_4862);
or U5636 (N_5636,N_4159,N_4544);
nand U5637 (N_5637,N_4320,N_4304);
xor U5638 (N_5638,N_4515,N_4672);
and U5639 (N_5639,N_4704,N_4050);
nand U5640 (N_5640,N_4323,N_4946);
or U5641 (N_5641,N_4543,N_4520);
and U5642 (N_5642,N_4581,N_4769);
nand U5643 (N_5643,N_4322,N_4408);
and U5644 (N_5644,N_4782,N_4363);
xor U5645 (N_5645,N_4854,N_4211);
and U5646 (N_5646,N_4718,N_4956);
xor U5647 (N_5647,N_4381,N_4256);
nand U5648 (N_5648,N_4570,N_4108);
or U5649 (N_5649,N_4890,N_4322);
or U5650 (N_5650,N_4920,N_4438);
xnor U5651 (N_5651,N_4747,N_4797);
or U5652 (N_5652,N_4027,N_4610);
or U5653 (N_5653,N_4148,N_4258);
nand U5654 (N_5654,N_4027,N_4547);
nor U5655 (N_5655,N_4619,N_4970);
and U5656 (N_5656,N_4096,N_4962);
xor U5657 (N_5657,N_4042,N_4968);
or U5658 (N_5658,N_4580,N_4674);
nor U5659 (N_5659,N_4176,N_4679);
or U5660 (N_5660,N_4395,N_4590);
nor U5661 (N_5661,N_4998,N_4844);
nand U5662 (N_5662,N_4321,N_4075);
or U5663 (N_5663,N_4232,N_4806);
nand U5664 (N_5664,N_4505,N_4158);
and U5665 (N_5665,N_4969,N_4303);
nor U5666 (N_5666,N_4344,N_4794);
xor U5667 (N_5667,N_4644,N_4187);
or U5668 (N_5668,N_4814,N_4501);
nor U5669 (N_5669,N_4685,N_4708);
or U5670 (N_5670,N_4573,N_4145);
nand U5671 (N_5671,N_4684,N_4359);
nand U5672 (N_5672,N_4253,N_4731);
or U5673 (N_5673,N_4364,N_4726);
or U5674 (N_5674,N_4861,N_4880);
and U5675 (N_5675,N_4880,N_4278);
xor U5676 (N_5676,N_4164,N_4544);
nor U5677 (N_5677,N_4156,N_4004);
or U5678 (N_5678,N_4335,N_4612);
nand U5679 (N_5679,N_4077,N_4063);
or U5680 (N_5680,N_4903,N_4119);
nor U5681 (N_5681,N_4457,N_4711);
or U5682 (N_5682,N_4606,N_4242);
xnor U5683 (N_5683,N_4825,N_4170);
xor U5684 (N_5684,N_4855,N_4886);
nor U5685 (N_5685,N_4095,N_4336);
nand U5686 (N_5686,N_4701,N_4480);
and U5687 (N_5687,N_4718,N_4179);
xnor U5688 (N_5688,N_4876,N_4090);
xnor U5689 (N_5689,N_4276,N_4676);
and U5690 (N_5690,N_4458,N_4438);
nor U5691 (N_5691,N_4404,N_4780);
nor U5692 (N_5692,N_4638,N_4281);
nor U5693 (N_5693,N_4895,N_4421);
xnor U5694 (N_5694,N_4014,N_4952);
xnor U5695 (N_5695,N_4338,N_4702);
xor U5696 (N_5696,N_4544,N_4249);
nand U5697 (N_5697,N_4507,N_4300);
xnor U5698 (N_5698,N_4532,N_4089);
nand U5699 (N_5699,N_4773,N_4610);
and U5700 (N_5700,N_4220,N_4653);
nor U5701 (N_5701,N_4498,N_4814);
nand U5702 (N_5702,N_4711,N_4728);
xnor U5703 (N_5703,N_4329,N_4445);
nand U5704 (N_5704,N_4357,N_4926);
nor U5705 (N_5705,N_4308,N_4449);
nand U5706 (N_5706,N_4944,N_4367);
and U5707 (N_5707,N_4826,N_4336);
nand U5708 (N_5708,N_4888,N_4710);
nor U5709 (N_5709,N_4811,N_4530);
xor U5710 (N_5710,N_4442,N_4413);
nand U5711 (N_5711,N_4929,N_4245);
xnor U5712 (N_5712,N_4474,N_4140);
or U5713 (N_5713,N_4753,N_4911);
nand U5714 (N_5714,N_4848,N_4562);
nor U5715 (N_5715,N_4820,N_4938);
xor U5716 (N_5716,N_4778,N_4161);
nor U5717 (N_5717,N_4401,N_4412);
or U5718 (N_5718,N_4989,N_4006);
nor U5719 (N_5719,N_4560,N_4515);
xor U5720 (N_5720,N_4436,N_4617);
xnor U5721 (N_5721,N_4860,N_4425);
and U5722 (N_5722,N_4550,N_4855);
xnor U5723 (N_5723,N_4275,N_4935);
and U5724 (N_5724,N_4956,N_4141);
or U5725 (N_5725,N_4262,N_4120);
nand U5726 (N_5726,N_4069,N_4494);
or U5727 (N_5727,N_4554,N_4615);
and U5728 (N_5728,N_4201,N_4076);
nand U5729 (N_5729,N_4012,N_4461);
or U5730 (N_5730,N_4005,N_4140);
and U5731 (N_5731,N_4674,N_4626);
and U5732 (N_5732,N_4733,N_4860);
nand U5733 (N_5733,N_4476,N_4999);
nor U5734 (N_5734,N_4558,N_4087);
nor U5735 (N_5735,N_4862,N_4727);
nor U5736 (N_5736,N_4387,N_4415);
xnor U5737 (N_5737,N_4310,N_4030);
and U5738 (N_5738,N_4851,N_4477);
nand U5739 (N_5739,N_4459,N_4611);
xor U5740 (N_5740,N_4799,N_4425);
and U5741 (N_5741,N_4256,N_4648);
nand U5742 (N_5742,N_4736,N_4720);
xnor U5743 (N_5743,N_4531,N_4048);
xnor U5744 (N_5744,N_4420,N_4891);
or U5745 (N_5745,N_4190,N_4527);
xor U5746 (N_5746,N_4235,N_4088);
xor U5747 (N_5747,N_4954,N_4757);
nand U5748 (N_5748,N_4536,N_4767);
nor U5749 (N_5749,N_4128,N_4969);
nand U5750 (N_5750,N_4783,N_4558);
xor U5751 (N_5751,N_4411,N_4632);
and U5752 (N_5752,N_4267,N_4317);
nor U5753 (N_5753,N_4631,N_4444);
or U5754 (N_5754,N_4207,N_4065);
nand U5755 (N_5755,N_4235,N_4625);
or U5756 (N_5756,N_4116,N_4038);
and U5757 (N_5757,N_4601,N_4163);
nor U5758 (N_5758,N_4155,N_4099);
nand U5759 (N_5759,N_4492,N_4812);
or U5760 (N_5760,N_4105,N_4246);
xor U5761 (N_5761,N_4003,N_4226);
nor U5762 (N_5762,N_4774,N_4884);
and U5763 (N_5763,N_4538,N_4107);
nor U5764 (N_5764,N_4683,N_4623);
or U5765 (N_5765,N_4852,N_4505);
xnor U5766 (N_5766,N_4639,N_4248);
and U5767 (N_5767,N_4906,N_4872);
and U5768 (N_5768,N_4693,N_4830);
and U5769 (N_5769,N_4756,N_4401);
xor U5770 (N_5770,N_4781,N_4791);
and U5771 (N_5771,N_4072,N_4756);
xnor U5772 (N_5772,N_4537,N_4619);
nand U5773 (N_5773,N_4217,N_4489);
or U5774 (N_5774,N_4731,N_4368);
nand U5775 (N_5775,N_4851,N_4058);
nor U5776 (N_5776,N_4118,N_4024);
nor U5777 (N_5777,N_4944,N_4505);
and U5778 (N_5778,N_4360,N_4839);
or U5779 (N_5779,N_4327,N_4931);
xnor U5780 (N_5780,N_4310,N_4245);
and U5781 (N_5781,N_4126,N_4759);
and U5782 (N_5782,N_4845,N_4393);
nor U5783 (N_5783,N_4904,N_4157);
nor U5784 (N_5784,N_4507,N_4938);
xor U5785 (N_5785,N_4956,N_4167);
xnor U5786 (N_5786,N_4638,N_4690);
and U5787 (N_5787,N_4046,N_4187);
xor U5788 (N_5788,N_4903,N_4146);
nor U5789 (N_5789,N_4590,N_4986);
nor U5790 (N_5790,N_4712,N_4123);
nor U5791 (N_5791,N_4930,N_4172);
or U5792 (N_5792,N_4232,N_4969);
nor U5793 (N_5793,N_4551,N_4465);
xor U5794 (N_5794,N_4555,N_4529);
nor U5795 (N_5795,N_4357,N_4505);
xnor U5796 (N_5796,N_4534,N_4769);
or U5797 (N_5797,N_4274,N_4666);
xnor U5798 (N_5798,N_4725,N_4270);
nor U5799 (N_5799,N_4178,N_4288);
or U5800 (N_5800,N_4313,N_4924);
nor U5801 (N_5801,N_4382,N_4368);
nand U5802 (N_5802,N_4602,N_4130);
xor U5803 (N_5803,N_4608,N_4369);
nor U5804 (N_5804,N_4045,N_4246);
nor U5805 (N_5805,N_4982,N_4245);
or U5806 (N_5806,N_4298,N_4950);
xor U5807 (N_5807,N_4724,N_4018);
or U5808 (N_5808,N_4149,N_4560);
nand U5809 (N_5809,N_4465,N_4137);
xor U5810 (N_5810,N_4075,N_4816);
nand U5811 (N_5811,N_4652,N_4999);
or U5812 (N_5812,N_4566,N_4429);
nor U5813 (N_5813,N_4273,N_4382);
nand U5814 (N_5814,N_4072,N_4969);
nor U5815 (N_5815,N_4738,N_4982);
or U5816 (N_5816,N_4089,N_4873);
or U5817 (N_5817,N_4799,N_4186);
or U5818 (N_5818,N_4811,N_4852);
or U5819 (N_5819,N_4364,N_4359);
and U5820 (N_5820,N_4415,N_4176);
nand U5821 (N_5821,N_4173,N_4766);
nand U5822 (N_5822,N_4342,N_4338);
nor U5823 (N_5823,N_4841,N_4645);
nand U5824 (N_5824,N_4902,N_4630);
or U5825 (N_5825,N_4994,N_4014);
nand U5826 (N_5826,N_4030,N_4333);
nor U5827 (N_5827,N_4121,N_4568);
nor U5828 (N_5828,N_4381,N_4466);
nand U5829 (N_5829,N_4181,N_4280);
or U5830 (N_5830,N_4322,N_4012);
and U5831 (N_5831,N_4752,N_4786);
nand U5832 (N_5832,N_4417,N_4254);
xnor U5833 (N_5833,N_4646,N_4245);
nand U5834 (N_5834,N_4124,N_4678);
nor U5835 (N_5835,N_4626,N_4105);
or U5836 (N_5836,N_4368,N_4103);
xor U5837 (N_5837,N_4704,N_4312);
nand U5838 (N_5838,N_4768,N_4036);
and U5839 (N_5839,N_4448,N_4298);
nor U5840 (N_5840,N_4737,N_4067);
xor U5841 (N_5841,N_4260,N_4900);
and U5842 (N_5842,N_4771,N_4925);
or U5843 (N_5843,N_4949,N_4991);
or U5844 (N_5844,N_4838,N_4856);
or U5845 (N_5845,N_4363,N_4180);
and U5846 (N_5846,N_4016,N_4454);
nor U5847 (N_5847,N_4743,N_4488);
nand U5848 (N_5848,N_4642,N_4956);
xnor U5849 (N_5849,N_4860,N_4919);
and U5850 (N_5850,N_4647,N_4136);
and U5851 (N_5851,N_4333,N_4651);
or U5852 (N_5852,N_4924,N_4467);
xor U5853 (N_5853,N_4663,N_4736);
nor U5854 (N_5854,N_4620,N_4541);
and U5855 (N_5855,N_4255,N_4742);
nor U5856 (N_5856,N_4419,N_4883);
xor U5857 (N_5857,N_4193,N_4213);
or U5858 (N_5858,N_4185,N_4622);
nor U5859 (N_5859,N_4249,N_4537);
or U5860 (N_5860,N_4535,N_4403);
nand U5861 (N_5861,N_4433,N_4688);
nor U5862 (N_5862,N_4661,N_4004);
xnor U5863 (N_5863,N_4191,N_4532);
nand U5864 (N_5864,N_4221,N_4692);
xor U5865 (N_5865,N_4340,N_4910);
xor U5866 (N_5866,N_4597,N_4170);
or U5867 (N_5867,N_4655,N_4461);
nor U5868 (N_5868,N_4499,N_4953);
nand U5869 (N_5869,N_4767,N_4221);
nor U5870 (N_5870,N_4056,N_4289);
nand U5871 (N_5871,N_4637,N_4736);
or U5872 (N_5872,N_4390,N_4895);
xor U5873 (N_5873,N_4841,N_4695);
xor U5874 (N_5874,N_4018,N_4987);
and U5875 (N_5875,N_4064,N_4939);
and U5876 (N_5876,N_4086,N_4067);
nand U5877 (N_5877,N_4127,N_4544);
nand U5878 (N_5878,N_4779,N_4286);
and U5879 (N_5879,N_4704,N_4673);
and U5880 (N_5880,N_4252,N_4976);
or U5881 (N_5881,N_4974,N_4558);
nand U5882 (N_5882,N_4879,N_4206);
or U5883 (N_5883,N_4834,N_4339);
and U5884 (N_5884,N_4554,N_4401);
xor U5885 (N_5885,N_4691,N_4302);
or U5886 (N_5886,N_4314,N_4283);
nand U5887 (N_5887,N_4743,N_4593);
or U5888 (N_5888,N_4629,N_4554);
and U5889 (N_5889,N_4387,N_4321);
or U5890 (N_5890,N_4513,N_4060);
nor U5891 (N_5891,N_4936,N_4764);
xnor U5892 (N_5892,N_4148,N_4982);
nor U5893 (N_5893,N_4693,N_4234);
nor U5894 (N_5894,N_4506,N_4661);
or U5895 (N_5895,N_4632,N_4132);
nand U5896 (N_5896,N_4003,N_4626);
nor U5897 (N_5897,N_4776,N_4550);
nand U5898 (N_5898,N_4384,N_4489);
nor U5899 (N_5899,N_4627,N_4196);
xor U5900 (N_5900,N_4958,N_4297);
nor U5901 (N_5901,N_4651,N_4621);
nor U5902 (N_5902,N_4401,N_4626);
nor U5903 (N_5903,N_4935,N_4990);
and U5904 (N_5904,N_4373,N_4508);
nor U5905 (N_5905,N_4433,N_4613);
nor U5906 (N_5906,N_4425,N_4157);
nand U5907 (N_5907,N_4189,N_4965);
xnor U5908 (N_5908,N_4339,N_4992);
or U5909 (N_5909,N_4772,N_4913);
and U5910 (N_5910,N_4544,N_4711);
xor U5911 (N_5911,N_4387,N_4890);
nor U5912 (N_5912,N_4309,N_4043);
and U5913 (N_5913,N_4701,N_4094);
xnor U5914 (N_5914,N_4317,N_4701);
and U5915 (N_5915,N_4495,N_4566);
nand U5916 (N_5916,N_4175,N_4840);
xnor U5917 (N_5917,N_4354,N_4077);
or U5918 (N_5918,N_4882,N_4363);
nor U5919 (N_5919,N_4541,N_4235);
or U5920 (N_5920,N_4868,N_4808);
and U5921 (N_5921,N_4219,N_4442);
nor U5922 (N_5922,N_4575,N_4427);
xnor U5923 (N_5923,N_4929,N_4038);
nand U5924 (N_5924,N_4855,N_4966);
or U5925 (N_5925,N_4887,N_4761);
xor U5926 (N_5926,N_4601,N_4288);
nand U5927 (N_5927,N_4055,N_4539);
nor U5928 (N_5928,N_4554,N_4995);
nor U5929 (N_5929,N_4453,N_4644);
or U5930 (N_5930,N_4773,N_4311);
or U5931 (N_5931,N_4966,N_4345);
or U5932 (N_5932,N_4800,N_4006);
or U5933 (N_5933,N_4316,N_4578);
nor U5934 (N_5934,N_4765,N_4685);
or U5935 (N_5935,N_4571,N_4412);
xor U5936 (N_5936,N_4606,N_4540);
xnor U5937 (N_5937,N_4479,N_4990);
nand U5938 (N_5938,N_4444,N_4219);
and U5939 (N_5939,N_4718,N_4167);
or U5940 (N_5940,N_4894,N_4274);
nand U5941 (N_5941,N_4738,N_4933);
xor U5942 (N_5942,N_4516,N_4215);
xor U5943 (N_5943,N_4296,N_4456);
nand U5944 (N_5944,N_4453,N_4956);
and U5945 (N_5945,N_4055,N_4457);
nand U5946 (N_5946,N_4212,N_4376);
and U5947 (N_5947,N_4254,N_4846);
nand U5948 (N_5948,N_4338,N_4641);
or U5949 (N_5949,N_4905,N_4303);
or U5950 (N_5950,N_4794,N_4720);
xor U5951 (N_5951,N_4383,N_4456);
or U5952 (N_5952,N_4408,N_4745);
and U5953 (N_5953,N_4441,N_4081);
or U5954 (N_5954,N_4848,N_4663);
nand U5955 (N_5955,N_4748,N_4816);
nor U5956 (N_5956,N_4396,N_4787);
or U5957 (N_5957,N_4243,N_4175);
or U5958 (N_5958,N_4079,N_4584);
nor U5959 (N_5959,N_4701,N_4738);
nor U5960 (N_5960,N_4176,N_4066);
nand U5961 (N_5961,N_4375,N_4944);
or U5962 (N_5962,N_4958,N_4675);
xor U5963 (N_5963,N_4614,N_4121);
nand U5964 (N_5964,N_4778,N_4540);
nand U5965 (N_5965,N_4377,N_4849);
nor U5966 (N_5966,N_4442,N_4420);
and U5967 (N_5967,N_4521,N_4137);
nor U5968 (N_5968,N_4653,N_4357);
or U5969 (N_5969,N_4727,N_4813);
nor U5970 (N_5970,N_4857,N_4337);
nand U5971 (N_5971,N_4896,N_4153);
nor U5972 (N_5972,N_4409,N_4662);
and U5973 (N_5973,N_4021,N_4551);
nand U5974 (N_5974,N_4801,N_4997);
and U5975 (N_5975,N_4667,N_4238);
nor U5976 (N_5976,N_4566,N_4132);
nor U5977 (N_5977,N_4112,N_4855);
and U5978 (N_5978,N_4201,N_4134);
or U5979 (N_5979,N_4169,N_4867);
or U5980 (N_5980,N_4376,N_4819);
nand U5981 (N_5981,N_4704,N_4303);
nor U5982 (N_5982,N_4428,N_4303);
nor U5983 (N_5983,N_4464,N_4160);
xnor U5984 (N_5984,N_4954,N_4492);
xor U5985 (N_5985,N_4110,N_4842);
or U5986 (N_5986,N_4380,N_4677);
and U5987 (N_5987,N_4686,N_4017);
nor U5988 (N_5988,N_4504,N_4292);
nor U5989 (N_5989,N_4516,N_4374);
and U5990 (N_5990,N_4193,N_4804);
or U5991 (N_5991,N_4531,N_4712);
nand U5992 (N_5992,N_4492,N_4761);
nor U5993 (N_5993,N_4128,N_4132);
or U5994 (N_5994,N_4541,N_4164);
and U5995 (N_5995,N_4373,N_4053);
nand U5996 (N_5996,N_4105,N_4577);
or U5997 (N_5997,N_4759,N_4726);
or U5998 (N_5998,N_4738,N_4521);
or U5999 (N_5999,N_4454,N_4615);
nand U6000 (N_6000,N_5856,N_5294);
xnor U6001 (N_6001,N_5829,N_5167);
nor U6002 (N_6002,N_5684,N_5103);
nor U6003 (N_6003,N_5094,N_5474);
nor U6004 (N_6004,N_5287,N_5008);
xnor U6005 (N_6005,N_5646,N_5476);
and U6006 (N_6006,N_5814,N_5597);
or U6007 (N_6007,N_5491,N_5468);
nand U6008 (N_6008,N_5300,N_5451);
nand U6009 (N_6009,N_5001,N_5582);
xor U6010 (N_6010,N_5198,N_5897);
xor U6011 (N_6011,N_5199,N_5720);
nor U6012 (N_6012,N_5450,N_5087);
xnor U6013 (N_6013,N_5818,N_5481);
or U6014 (N_6014,N_5953,N_5866);
and U6015 (N_6015,N_5955,N_5323);
xnor U6016 (N_6016,N_5742,N_5060);
xnor U6017 (N_6017,N_5432,N_5498);
xor U6018 (N_6018,N_5079,N_5281);
nor U6019 (N_6019,N_5427,N_5229);
nand U6020 (N_6020,N_5393,N_5091);
nor U6021 (N_6021,N_5022,N_5164);
and U6022 (N_6022,N_5739,N_5545);
nor U6023 (N_6023,N_5303,N_5993);
nand U6024 (N_6024,N_5553,N_5847);
nand U6025 (N_6025,N_5273,N_5762);
nand U6026 (N_6026,N_5188,N_5675);
or U6027 (N_6027,N_5196,N_5601);
nor U6028 (N_6028,N_5832,N_5958);
nand U6029 (N_6029,N_5013,N_5335);
nand U6030 (N_6030,N_5119,N_5066);
or U6031 (N_6031,N_5805,N_5666);
nand U6032 (N_6032,N_5678,N_5146);
xnor U6033 (N_6033,N_5193,N_5713);
nor U6034 (N_6034,N_5377,N_5584);
nor U6035 (N_6035,N_5685,N_5656);
and U6036 (N_6036,N_5072,N_5967);
xnor U6037 (N_6037,N_5279,N_5641);
or U6038 (N_6038,N_5497,N_5751);
or U6039 (N_6039,N_5041,N_5629);
and U6040 (N_6040,N_5373,N_5580);
and U6041 (N_6041,N_5268,N_5172);
and U6042 (N_6042,N_5746,N_5547);
nor U6043 (N_6043,N_5797,N_5860);
or U6044 (N_6044,N_5617,N_5435);
or U6045 (N_6045,N_5836,N_5098);
nor U6046 (N_6046,N_5006,N_5862);
and U6047 (N_6047,N_5980,N_5838);
and U6048 (N_6048,N_5423,N_5750);
xnor U6049 (N_6049,N_5525,N_5934);
xor U6050 (N_6050,N_5855,N_5467);
xnor U6051 (N_6051,N_5789,N_5674);
nor U6052 (N_6052,N_5744,N_5126);
nor U6053 (N_6053,N_5444,N_5181);
and U6054 (N_6054,N_5065,N_5891);
or U6055 (N_6055,N_5407,N_5833);
xnor U6056 (N_6056,N_5668,N_5526);
and U6057 (N_6057,N_5219,N_5489);
and U6058 (N_6058,N_5942,N_5364);
and U6059 (N_6059,N_5111,N_5705);
nor U6060 (N_6060,N_5828,N_5664);
or U6061 (N_6061,N_5345,N_5918);
and U6062 (N_6062,N_5056,N_5686);
nand U6063 (N_6063,N_5977,N_5113);
nor U6064 (N_6064,N_5716,N_5209);
nand U6065 (N_6065,N_5943,N_5027);
or U6066 (N_6066,N_5764,N_5213);
or U6067 (N_6067,N_5844,N_5286);
xor U6068 (N_6068,N_5023,N_5966);
nand U6069 (N_6069,N_5506,N_5654);
xnor U6070 (N_6070,N_5592,N_5975);
xor U6071 (N_6071,N_5090,N_5140);
nand U6072 (N_6072,N_5698,N_5817);
nor U6073 (N_6073,N_5941,N_5226);
and U6074 (N_6074,N_5773,N_5124);
nand U6075 (N_6075,N_5327,N_5661);
nand U6076 (N_6076,N_5125,N_5517);
nand U6077 (N_6077,N_5488,N_5996);
nand U6078 (N_6078,N_5558,N_5288);
xnor U6079 (N_6079,N_5243,N_5298);
nor U6080 (N_6080,N_5798,N_5130);
and U6081 (N_6081,N_5121,N_5433);
nand U6082 (N_6082,N_5142,N_5129);
xor U6083 (N_6083,N_5136,N_5080);
nor U6084 (N_6084,N_5640,N_5493);
nor U6085 (N_6085,N_5986,N_5988);
xnor U6086 (N_6086,N_5050,N_5346);
and U6087 (N_6087,N_5790,N_5403);
xor U6088 (N_6088,N_5203,N_5912);
and U6089 (N_6089,N_5340,N_5064);
or U6090 (N_6090,N_5551,N_5053);
or U6091 (N_6091,N_5852,N_5822);
or U6092 (N_6092,N_5054,N_5873);
or U6093 (N_6093,N_5510,N_5619);
xor U6094 (N_6094,N_5483,N_5304);
nor U6095 (N_6095,N_5183,N_5894);
or U6096 (N_6096,N_5033,N_5263);
nor U6097 (N_6097,N_5507,N_5767);
or U6098 (N_6098,N_5568,N_5003);
and U6099 (N_6099,N_5421,N_5449);
nand U6100 (N_6100,N_5613,N_5005);
and U6101 (N_6101,N_5715,N_5061);
or U6102 (N_6102,N_5906,N_5276);
xor U6103 (N_6103,N_5149,N_5959);
and U6104 (N_6104,N_5267,N_5907);
xnor U6105 (N_6105,N_5979,N_5439);
and U6106 (N_6106,N_5606,N_5448);
nand U6107 (N_6107,N_5443,N_5913);
nand U6108 (N_6108,N_5047,N_5143);
and U6109 (N_6109,N_5043,N_5075);
or U6110 (N_6110,N_5630,N_5480);
nor U6111 (N_6111,N_5555,N_5846);
and U6112 (N_6112,N_5028,N_5719);
and U6113 (N_6113,N_5952,N_5610);
nand U6114 (N_6114,N_5157,N_5595);
and U6115 (N_6115,N_5578,N_5824);
or U6116 (N_6116,N_5233,N_5440);
or U6117 (N_6117,N_5815,N_5154);
and U6118 (N_6118,N_5254,N_5224);
and U6119 (N_6119,N_5241,N_5880);
or U6120 (N_6120,N_5379,N_5903);
or U6121 (N_6121,N_5573,N_5712);
xor U6122 (N_6122,N_5886,N_5730);
xnor U6123 (N_6123,N_5973,N_5417);
nor U6124 (N_6124,N_5776,N_5777);
nor U6125 (N_6125,N_5337,N_5394);
and U6126 (N_6126,N_5778,N_5469);
nand U6127 (N_6127,N_5518,N_5357);
nand U6128 (N_6128,N_5564,N_5455);
nand U6129 (N_6129,N_5385,N_5946);
nand U6130 (N_6130,N_5914,N_5117);
or U6131 (N_6131,N_5348,N_5579);
nor U6132 (N_6132,N_5724,N_5634);
or U6133 (N_6133,N_5658,N_5332);
nand U6134 (N_6134,N_5519,N_5073);
xor U6135 (N_6135,N_5660,N_5312);
nand U6136 (N_6136,N_5296,N_5131);
or U6137 (N_6137,N_5158,N_5145);
xor U6138 (N_6138,N_5097,N_5275);
nand U6139 (N_6139,N_5479,N_5082);
and U6140 (N_6140,N_5883,N_5272);
nor U6141 (N_6141,N_5549,N_5347);
nor U6142 (N_6142,N_5736,N_5222);
or U6143 (N_6143,N_5513,N_5699);
nand U6144 (N_6144,N_5992,N_5755);
xnor U6145 (N_6145,N_5989,N_5301);
and U6146 (N_6146,N_5366,N_5763);
or U6147 (N_6147,N_5189,N_5232);
or U6148 (N_6148,N_5851,N_5714);
or U6149 (N_6149,N_5741,N_5826);
nand U6150 (N_6150,N_5620,N_5882);
nand U6151 (N_6151,N_5544,N_5342);
or U6152 (N_6152,N_5827,N_5037);
and U6153 (N_6153,N_5922,N_5933);
xnor U6154 (N_6154,N_5850,N_5672);
and U6155 (N_6155,N_5501,N_5425);
xnor U6156 (N_6156,N_5841,N_5169);
xor U6157 (N_6157,N_5960,N_5305);
nor U6158 (N_6158,N_5839,N_5138);
xor U6159 (N_6159,N_5995,N_5253);
nor U6160 (N_6160,N_5651,N_5593);
nand U6161 (N_6161,N_5105,N_5796);
nand U6162 (N_6162,N_5810,N_5076);
nand U6163 (N_6163,N_5255,N_5944);
nand U6164 (N_6164,N_5024,N_5919);
nand U6165 (N_6165,N_5878,N_5539);
nand U6166 (N_6166,N_5307,N_5358);
nor U6167 (N_6167,N_5529,N_5245);
xnor U6168 (N_6168,N_5144,N_5123);
or U6169 (N_6169,N_5530,N_5420);
and U6170 (N_6170,N_5494,N_5293);
nand U6171 (N_6171,N_5331,N_5864);
or U6172 (N_6172,N_5554,N_5905);
xor U6173 (N_6173,N_5228,N_5051);
or U6174 (N_6174,N_5831,N_5152);
nand U6175 (N_6175,N_5436,N_5676);
nand U6176 (N_6176,N_5095,N_5132);
nand U6177 (N_6177,N_5793,N_5689);
nor U6178 (N_6178,N_5260,N_5957);
xnor U6179 (N_6179,N_5632,N_5088);
or U6180 (N_6180,N_5608,N_5376);
nor U6181 (N_6181,N_5575,N_5457);
or U6182 (N_6182,N_5928,N_5819);
nand U6183 (N_6183,N_5354,N_5984);
xnor U6184 (N_6184,N_5461,N_5585);
or U6185 (N_6185,N_5801,N_5070);
xnor U6186 (N_6186,N_5035,N_5251);
and U6187 (N_6187,N_5004,N_5557);
and U6188 (N_6188,N_5156,N_5207);
or U6189 (N_6189,N_5625,N_5182);
and U6190 (N_6190,N_5478,N_5802);
and U6191 (N_6191,N_5422,N_5258);
xor U6192 (N_6192,N_5590,N_5548);
nand U6193 (N_6193,N_5236,N_5931);
nand U6194 (N_6194,N_5963,N_5502);
xnor U6195 (N_6195,N_5223,N_5218);
and U6196 (N_6196,N_5969,N_5133);
nand U6197 (N_6197,N_5534,N_5069);
and U6198 (N_6198,N_5752,N_5671);
and U6199 (N_6199,N_5285,N_5567);
nor U6200 (N_6200,N_5338,N_5127);
nand U6201 (N_6201,N_5441,N_5911);
nor U6202 (N_6202,N_5291,N_5092);
or U6203 (N_6203,N_5308,N_5187);
and U6204 (N_6204,N_5099,N_5700);
and U6205 (N_6205,N_5679,N_5411);
nor U6206 (N_6206,N_5353,N_5782);
nor U6207 (N_6207,N_5639,N_5418);
xnor U6208 (N_6208,N_5879,N_5367);
nor U6209 (N_6209,N_5197,N_5761);
xor U6210 (N_6210,N_5078,N_5760);
nand U6211 (N_6211,N_5779,N_5221);
nand U6212 (N_6212,N_5180,N_5375);
nand U6213 (N_6213,N_5701,N_5981);
nand U6214 (N_6214,N_5825,N_5572);
xnor U6215 (N_6215,N_5522,N_5540);
xor U6216 (N_6216,N_5310,N_5631);
and U6217 (N_6217,N_5192,N_5333);
or U6218 (N_6218,N_5800,N_5515);
xor U6219 (N_6219,N_5612,N_5032);
and U6220 (N_6220,N_5516,N_5437);
nor U6221 (N_6221,N_5854,N_5747);
nor U6222 (N_6222,N_5390,N_5754);
nand U6223 (N_6223,N_5871,N_5329);
nor U6224 (N_6224,N_5402,N_5570);
or U6225 (N_6225,N_5150,N_5527);
or U6226 (N_6226,N_5533,N_5278);
nor U6227 (N_6227,N_5615,N_5324);
or U6228 (N_6228,N_5175,N_5428);
xnor U6229 (N_6229,N_5721,N_5837);
nand U6230 (N_6230,N_5100,N_5677);
or U6231 (N_6231,N_5343,N_5128);
nand U6232 (N_6232,N_5514,N_5409);
xor U6233 (N_6233,N_5475,N_5165);
xor U6234 (N_6234,N_5982,N_5561);
nand U6235 (N_6235,N_5319,N_5234);
and U6236 (N_6236,N_5937,N_5148);
nor U6237 (N_6237,N_5994,N_5014);
xor U6238 (N_6238,N_5574,N_5045);
nor U6239 (N_6239,N_5673,N_5295);
nor U6240 (N_6240,N_5214,N_5642);
nand U6241 (N_6241,N_5991,N_5936);
and U6242 (N_6242,N_5650,N_5336);
nand U6243 (N_6243,N_5875,N_5780);
or U6244 (N_6244,N_5067,N_5737);
nor U6245 (N_6245,N_5453,N_5274);
nand U6246 (N_6246,N_5495,N_5857);
nor U6247 (N_6247,N_5247,N_5604);
nor U6248 (N_6248,N_5786,N_5265);
nand U6249 (N_6249,N_5044,N_5869);
nor U6250 (N_6250,N_5690,N_5283);
xnor U6251 (N_6251,N_5369,N_5821);
or U6252 (N_6252,N_5011,N_5589);
nand U6253 (N_6253,N_5624,N_5729);
and U6254 (N_6254,N_5473,N_5783);
xor U6255 (N_6255,N_5010,N_5999);
nor U6256 (N_6256,N_5904,N_5885);
xnor U6257 (N_6257,N_5531,N_5374);
xnor U6258 (N_6258,N_5397,N_5884);
or U6259 (N_6259,N_5868,N_5063);
nor U6260 (N_6260,N_5909,N_5983);
or U6261 (N_6261,N_5408,N_5297);
xnor U6262 (N_6262,N_5771,N_5965);
nand U6263 (N_6263,N_5788,N_5681);
or U6264 (N_6264,N_5770,N_5888);
xor U6265 (N_6265,N_5848,N_5636);
and U6266 (N_6266,N_5511,N_5723);
xor U6267 (N_6267,N_5381,N_5876);
and U6268 (N_6268,N_5361,N_5034);
nand U6269 (N_6269,N_5401,N_5482);
nand U6270 (N_6270,N_5052,N_5081);
or U6271 (N_6271,N_5466,N_5987);
and U6272 (N_6272,N_5018,N_5261);
nor U6273 (N_6273,N_5571,N_5220);
or U6274 (N_6274,N_5454,N_5021);
and U6275 (N_6275,N_5895,N_5104);
nor U6276 (N_6276,N_5732,N_5244);
or U6277 (N_6277,N_5176,N_5009);
xnor U6278 (N_6278,N_5315,N_5706);
or U6279 (N_6279,N_5692,N_5405);
xnor U6280 (N_6280,N_5485,N_5110);
or U6281 (N_6281,N_5161,N_5842);
xor U6282 (N_6282,N_5910,N_5598);
nor U6283 (N_6283,N_5849,N_5908);
nor U6284 (N_6284,N_5388,N_5787);
or U6285 (N_6285,N_5458,N_5599);
xnor U6286 (N_6286,N_5669,N_5252);
or U6287 (N_6287,N_5536,N_5865);
and U6288 (N_6288,N_5968,N_5626);
nand U6289 (N_6289,N_5362,N_5118);
and U6290 (N_6290,N_5093,N_5270);
and U6291 (N_6291,N_5687,N_5616);
and U6292 (N_6292,N_5622,N_5940);
xnor U6293 (N_6293,N_5368,N_5935);
and U6294 (N_6294,N_5807,N_5320);
nor U6295 (N_6295,N_5030,N_5330);
nor U6296 (N_6296,N_5947,N_5985);
xnor U6297 (N_6297,N_5670,N_5535);
or U6298 (N_6298,N_5945,N_5046);
or U6299 (N_6299,N_5108,N_5249);
nand U6300 (N_6300,N_5496,N_5434);
nand U6301 (N_6301,N_5726,N_5920);
nor U6302 (N_6302,N_5964,N_5059);
nand U6303 (N_6303,N_5753,N_5112);
nor U6304 (N_6304,N_5738,N_5899);
nor U6305 (N_6305,N_5107,N_5231);
xnor U6306 (N_6306,N_5185,N_5867);
or U6307 (N_6307,N_5404,N_5049);
nand U6308 (N_6308,N_5413,N_5872);
or U6309 (N_6309,N_5178,N_5976);
or U6310 (N_6310,N_5840,N_5282);
and U6311 (N_6311,N_5134,N_5521);
and U6312 (N_6312,N_5137,N_5808);
nand U6313 (N_6313,N_5302,N_5280);
nand U6314 (N_6314,N_5603,N_5204);
and U6315 (N_6315,N_5735,N_5902);
or U6316 (N_6316,N_5745,N_5649);
nand U6317 (N_6317,N_5722,N_5834);
nand U6318 (N_6318,N_5352,N_5812);
and U6319 (N_6319,N_5240,N_5292);
nand U6320 (N_6320,N_5384,N_5349);
and U6321 (N_6321,N_5925,N_5635);
or U6322 (N_6322,N_5765,N_5811);
or U6323 (N_6323,N_5299,N_5339);
nand U6324 (N_6324,N_5758,N_5471);
and U6325 (N_6325,N_5503,N_5365);
xnor U6326 (N_6326,N_5250,N_5256);
nor U6327 (N_6327,N_5160,N_5313);
or U6328 (N_6328,N_5392,N_5523);
nor U6329 (N_6329,N_5015,N_5877);
nand U6330 (N_6330,N_5962,N_5470);
nor U6331 (N_6331,N_5621,N_5637);
nand U6332 (N_6332,N_5900,N_5490);
xnor U6333 (N_6333,N_5628,N_5749);
nand U6334 (N_6334,N_5896,N_5201);
and U6335 (N_6335,N_5114,N_5707);
or U6336 (N_6336,N_5007,N_5215);
nand U6337 (N_6337,N_5101,N_5546);
nor U6338 (N_6338,N_5600,N_5926);
and U6339 (N_6339,N_5655,N_5016);
xnor U6340 (N_6340,N_5733,N_5644);
and U6341 (N_6341,N_5794,N_5520);
or U6342 (N_6342,N_5566,N_5356);
xor U6343 (N_6343,N_5084,N_5410);
nor U6344 (N_6344,N_5116,N_5717);
and U6345 (N_6345,N_5212,N_5326);
nand U6346 (N_6346,N_5089,N_5389);
or U6347 (N_6347,N_5806,N_5704);
xnor U6348 (N_6348,N_5487,N_5170);
xnor U6349 (N_6349,N_5923,N_5731);
or U6350 (N_6350,N_5057,N_5887);
or U6351 (N_6351,N_5970,N_5859);
or U6352 (N_6352,N_5031,N_5486);
xnor U6353 (N_6353,N_5665,N_5217);
nor U6354 (N_6354,N_5257,N_5835);
nor U6355 (N_6355,N_5205,N_5039);
nor U6356 (N_6356,N_5785,N_5077);
or U6357 (N_6357,N_5321,N_5951);
or U6358 (N_6358,N_5186,N_5820);
nand U6359 (N_6359,N_5162,N_5972);
nor U6360 (N_6360,N_5643,N_5442);
nand U6361 (N_6361,N_5492,N_5757);
nand U6362 (N_6362,N_5956,N_5916);
nor U6363 (N_6363,N_5317,N_5929);
nor U6364 (N_6364,N_5431,N_5718);
or U6365 (N_6365,N_5378,N_5759);
or U6366 (N_6366,N_5652,N_5858);
nand U6367 (N_6367,N_5823,N_5627);
or U6368 (N_6368,N_5932,N_5804);
nor U6369 (N_6369,N_5085,N_5845);
nand U6370 (N_6370,N_5924,N_5769);
and U6371 (N_6371,N_5216,N_5948);
or U6372 (N_6372,N_5269,N_5447);
nor U6373 (N_6373,N_5768,N_5153);
xor U6374 (N_6374,N_5618,N_5227);
and U6375 (N_6375,N_5784,N_5532);
or U6376 (N_6376,N_5195,N_5238);
or U6377 (N_6377,N_5371,N_5290);
nand U6378 (N_6378,N_5938,N_5708);
nand U6379 (N_6379,N_5355,N_5792);
or U6380 (N_6380,N_5576,N_5040);
nand U6381 (N_6381,N_5106,N_5974);
nand U6382 (N_6382,N_5562,N_5688);
or U6383 (N_6383,N_5556,N_5372);
or U6384 (N_6384,N_5237,N_5206);
or U6385 (N_6385,N_5863,N_5309);
and U6386 (N_6386,N_5605,N_5177);
nand U6387 (N_6387,N_5452,N_5505);
or U6388 (N_6388,N_5645,N_5775);
nor U6389 (N_6389,N_5843,N_5277);
nand U6390 (N_6390,N_5068,N_5772);
nor U6391 (N_6391,N_5416,N_5359);
nor U6392 (N_6392,N_5159,N_5591);
or U6393 (N_6393,N_5262,N_5200);
nand U6394 (N_6394,N_5102,N_5978);
nor U6395 (N_6395,N_5155,N_5194);
nor U6396 (N_6396,N_5813,N_5596);
xnor U6397 (N_6397,N_5399,N_5017);
and U6398 (N_6398,N_5950,N_5083);
or U6399 (N_6399,N_5509,N_5949);
xor U6400 (N_6400,N_5477,N_5874);
xnor U6401 (N_6401,N_5259,N_5391);
or U6402 (N_6402,N_5500,N_5246);
xnor U6403 (N_6403,N_5702,N_5048);
xor U6404 (N_6404,N_5171,N_5743);
or U6405 (N_6405,N_5693,N_5609);
and U6406 (N_6406,N_5774,N_5289);
and U6407 (N_6407,N_5998,N_5151);
and U6408 (N_6408,N_5799,N_5683);
or U6409 (N_6409,N_5710,N_5235);
and U6410 (N_6410,N_5042,N_5122);
or U6411 (N_6411,N_5202,N_5086);
nand U6412 (N_6412,N_5602,N_5893);
or U6413 (N_6413,N_5853,N_5424);
or U6414 (N_6414,N_5395,N_5036);
and U6415 (N_6415,N_5695,N_5537);
or U6416 (N_6416,N_5648,N_5429);
or U6417 (N_6417,N_5426,N_5248);
xor U6418 (N_6418,N_5406,N_5727);
or U6419 (N_6419,N_5344,N_5930);
nor U6420 (N_6420,N_5472,N_5415);
nor U6421 (N_6421,N_5583,N_5271);
nor U6422 (N_6422,N_5647,N_5055);
nor U6423 (N_6423,N_5939,N_5456);
xor U6424 (N_6424,N_5350,N_5543);
nand U6425 (N_6425,N_5328,N_5552);
nor U6426 (N_6426,N_5264,N_5954);
or U6427 (N_6427,N_5325,N_5139);
or U6428 (N_6428,N_5889,N_5166);
or U6429 (N_6429,N_5830,N_5311);
nand U6430 (N_6430,N_5019,N_5135);
nor U6431 (N_6431,N_5682,N_5581);
or U6432 (N_6432,N_5725,N_5460);
nor U6433 (N_6433,N_5242,N_5809);
nand U6434 (N_6434,N_5230,N_5306);
nand U6435 (N_6435,N_5538,N_5638);
nor U6436 (N_6436,N_5921,N_5816);
nor U6437 (N_6437,N_5382,N_5588);
xnor U6438 (N_6438,N_5318,N_5781);
and U6439 (N_6439,N_5446,N_5915);
xnor U6440 (N_6440,N_5898,N_5795);
nand U6441 (N_6441,N_5740,N_5109);
nor U6442 (N_6442,N_5711,N_5550);
xnor U6443 (N_6443,N_5890,N_5614);
nand U6444 (N_6444,N_5691,N_5587);
nor U6445 (N_6445,N_5012,N_5314);
and U6446 (N_6446,N_5062,N_5284);
and U6447 (N_6447,N_5071,N_5594);
xnor U6448 (N_6448,N_5901,N_5662);
nand U6449 (N_6449,N_5191,N_5029);
nand U6450 (N_6450,N_5748,N_5168);
xnor U6451 (N_6451,N_5559,N_5484);
and U6452 (N_6452,N_5210,N_5504);
nor U6453 (N_6453,N_5803,N_5380);
and U6454 (N_6454,N_5508,N_5586);
nor U6455 (N_6455,N_5208,N_5419);
nor U6456 (N_6456,N_5462,N_5115);
xor U6457 (N_6457,N_5623,N_5351);
nand U6458 (N_6458,N_5892,N_5512);
nor U6459 (N_6459,N_5560,N_5025);
nand U6460 (N_6460,N_5756,N_5000);
or U6461 (N_6461,N_5412,N_5541);
nor U6462 (N_6462,N_5163,N_5653);
nor U6463 (N_6463,N_5499,N_5569);
xnor U6464 (N_6464,N_5147,N_5542);
xnor U6465 (N_6465,N_5728,N_5611);
and U6466 (N_6466,N_5387,N_5663);
xnor U6467 (N_6467,N_5002,N_5703);
or U6468 (N_6468,N_5341,N_5791);
nor U6469 (N_6469,N_5463,N_5020);
nand U6470 (N_6470,N_5096,N_5563);
xor U6471 (N_6471,N_5459,N_5383);
nor U6472 (N_6472,N_5363,N_5577);
nor U6473 (N_6473,N_5386,N_5211);
nor U6474 (N_6474,N_5398,N_5607);
and U6475 (N_6475,N_5697,N_5633);
or U6476 (N_6476,N_5657,N_5414);
nor U6477 (N_6477,N_5173,N_5659);
or U6478 (N_6478,N_5360,N_5528);
or U6479 (N_6479,N_5709,N_5438);
nor U6480 (N_6480,N_5026,N_5174);
nor U6481 (N_6481,N_5734,N_5927);
or U6482 (N_6482,N_5990,N_5120);
and U6483 (N_6483,N_5179,N_5445);
nand U6484 (N_6484,N_5430,N_5766);
and U6485 (N_6485,N_5184,N_5881);
nand U6486 (N_6486,N_5370,N_5524);
nor U6487 (N_6487,N_5058,N_5961);
xnor U6488 (N_6488,N_5917,N_5971);
nand U6489 (N_6489,N_5997,N_5465);
nor U6490 (N_6490,N_5141,N_5694);
or U6491 (N_6491,N_5316,N_5074);
nor U6492 (N_6492,N_5861,N_5565);
or U6493 (N_6493,N_5396,N_5266);
or U6494 (N_6494,N_5239,N_5225);
nor U6495 (N_6495,N_5680,N_5400);
and U6496 (N_6496,N_5038,N_5870);
and U6497 (N_6497,N_5667,N_5190);
xnor U6498 (N_6498,N_5696,N_5464);
nand U6499 (N_6499,N_5334,N_5322);
xor U6500 (N_6500,N_5756,N_5207);
nand U6501 (N_6501,N_5056,N_5080);
xor U6502 (N_6502,N_5736,N_5075);
xor U6503 (N_6503,N_5315,N_5952);
nand U6504 (N_6504,N_5268,N_5650);
and U6505 (N_6505,N_5270,N_5097);
xnor U6506 (N_6506,N_5928,N_5749);
or U6507 (N_6507,N_5090,N_5369);
and U6508 (N_6508,N_5364,N_5538);
xnor U6509 (N_6509,N_5554,N_5557);
and U6510 (N_6510,N_5563,N_5377);
nand U6511 (N_6511,N_5492,N_5369);
nand U6512 (N_6512,N_5484,N_5952);
and U6513 (N_6513,N_5467,N_5716);
nand U6514 (N_6514,N_5480,N_5209);
xnor U6515 (N_6515,N_5963,N_5382);
nor U6516 (N_6516,N_5265,N_5257);
xnor U6517 (N_6517,N_5728,N_5792);
nand U6518 (N_6518,N_5304,N_5316);
or U6519 (N_6519,N_5876,N_5471);
xnor U6520 (N_6520,N_5632,N_5823);
nand U6521 (N_6521,N_5159,N_5442);
or U6522 (N_6522,N_5600,N_5301);
or U6523 (N_6523,N_5155,N_5703);
nor U6524 (N_6524,N_5709,N_5137);
or U6525 (N_6525,N_5517,N_5854);
xor U6526 (N_6526,N_5512,N_5737);
nand U6527 (N_6527,N_5075,N_5255);
and U6528 (N_6528,N_5005,N_5177);
and U6529 (N_6529,N_5902,N_5093);
nor U6530 (N_6530,N_5510,N_5332);
and U6531 (N_6531,N_5637,N_5022);
nor U6532 (N_6532,N_5835,N_5183);
nand U6533 (N_6533,N_5466,N_5938);
nand U6534 (N_6534,N_5257,N_5521);
nor U6535 (N_6535,N_5786,N_5921);
nand U6536 (N_6536,N_5286,N_5074);
nor U6537 (N_6537,N_5879,N_5985);
or U6538 (N_6538,N_5973,N_5486);
and U6539 (N_6539,N_5111,N_5528);
and U6540 (N_6540,N_5041,N_5509);
xnor U6541 (N_6541,N_5988,N_5164);
or U6542 (N_6542,N_5559,N_5325);
or U6543 (N_6543,N_5192,N_5851);
and U6544 (N_6544,N_5291,N_5855);
nand U6545 (N_6545,N_5065,N_5806);
xor U6546 (N_6546,N_5524,N_5193);
nand U6547 (N_6547,N_5773,N_5114);
and U6548 (N_6548,N_5774,N_5447);
nor U6549 (N_6549,N_5251,N_5028);
xor U6550 (N_6550,N_5345,N_5667);
or U6551 (N_6551,N_5201,N_5284);
xnor U6552 (N_6552,N_5431,N_5711);
xnor U6553 (N_6553,N_5180,N_5760);
nand U6554 (N_6554,N_5729,N_5351);
or U6555 (N_6555,N_5985,N_5122);
and U6556 (N_6556,N_5723,N_5853);
nand U6557 (N_6557,N_5797,N_5145);
nand U6558 (N_6558,N_5230,N_5485);
xnor U6559 (N_6559,N_5358,N_5377);
nand U6560 (N_6560,N_5290,N_5307);
and U6561 (N_6561,N_5355,N_5696);
nor U6562 (N_6562,N_5744,N_5178);
and U6563 (N_6563,N_5697,N_5799);
and U6564 (N_6564,N_5402,N_5079);
or U6565 (N_6565,N_5683,N_5648);
nor U6566 (N_6566,N_5228,N_5531);
nand U6567 (N_6567,N_5855,N_5069);
or U6568 (N_6568,N_5484,N_5596);
nand U6569 (N_6569,N_5514,N_5363);
nand U6570 (N_6570,N_5668,N_5356);
xor U6571 (N_6571,N_5958,N_5698);
xnor U6572 (N_6572,N_5356,N_5626);
nor U6573 (N_6573,N_5253,N_5163);
xor U6574 (N_6574,N_5678,N_5754);
and U6575 (N_6575,N_5363,N_5051);
or U6576 (N_6576,N_5611,N_5324);
nand U6577 (N_6577,N_5905,N_5565);
nand U6578 (N_6578,N_5482,N_5810);
nand U6579 (N_6579,N_5570,N_5056);
or U6580 (N_6580,N_5044,N_5918);
nor U6581 (N_6581,N_5633,N_5569);
nand U6582 (N_6582,N_5726,N_5747);
nand U6583 (N_6583,N_5456,N_5376);
xor U6584 (N_6584,N_5013,N_5752);
nand U6585 (N_6585,N_5549,N_5875);
or U6586 (N_6586,N_5364,N_5656);
xor U6587 (N_6587,N_5864,N_5075);
nand U6588 (N_6588,N_5522,N_5444);
or U6589 (N_6589,N_5752,N_5718);
nand U6590 (N_6590,N_5256,N_5793);
and U6591 (N_6591,N_5844,N_5054);
xor U6592 (N_6592,N_5907,N_5143);
or U6593 (N_6593,N_5935,N_5808);
xnor U6594 (N_6594,N_5814,N_5704);
xor U6595 (N_6595,N_5068,N_5670);
and U6596 (N_6596,N_5129,N_5508);
nand U6597 (N_6597,N_5172,N_5889);
or U6598 (N_6598,N_5764,N_5610);
xnor U6599 (N_6599,N_5019,N_5863);
nand U6600 (N_6600,N_5577,N_5188);
or U6601 (N_6601,N_5911,N_5531);
xor U6602 (N_6602,N_5976,N_5161);
and U6603 (N_6603,N_5222,N_5633);
nand U6604 (N_6604,N_5898,N_5143);
or U6605 (N_6605,N_5881,N_5358);
or U6606 (N_6606,N_5363,N_5718);
nand U6607 (N_6607,N_5893,N_5243);
or U6608 (N_6608,N_5115,N_5926);
xor U6609 (N_6609,N_5554,N_5083);
nand U6610 (N_6610,N_5981,N_5898);
nand U6611 (N_6611,N_5250,N_5503);
xnor U6612 (N_6612,N_5423,N_5206);
and U6613 (N_6613,N_5350,N_5604);
nor U6614 (N_6614,N_5357,N_5661);
nor U6615 (N_6615,N_5368,N_5988);
nand U6616 (N_6616,N_5698,N_5115);
xor U6617 (N_6617,N_5268,N_5167);
xnor U6618 (N_6618,N_5778,N_5905);
or U6619 (N_6619,N_5166,N_5070);
or U6620 (N_6620,N_5280,N_5927);
and U6621 (N_6621,N_5913,N_5105);
nor U6622 (N_6622,N_5296,N_5038);
nor U6623 (N_6623,N_5093,N_5432);
nor U6624 (N_6624,N_5359,N_5273);
nand U6625 (N_6625,N_5350,N_5454);
or U6626 (N_6626,N_5996,N_5187);
nand U6627 (N_6627,N_5117,N_5656);
nand U6628 (N_6628,N_5581,N_5769);
or U6629 (N_6629,N_5530,N_5037);
nand U6630 (N_6630,N_5777,N_5201);
xor U6631 (N_6631,N_5128,N_5724);
nor U6632 (N_6632,N_5753,N_5140);
nand U6633 (N_6633,N_5815,N_5387);
nand U6634 (N_6634,N_5580,N_5020);
nand U6635 (N_6635,N_5648,N_5891);
nand U6636 (N_6636,N_5627,N_5412);
and U6637 (N_6637,N_5592,N_5200);
nand U6638 (N_6638,N_5714,N_5718);
and U6639 (N_6639,N_5644,N_5994);
and U6640 (N_6640,N_5195,N_5851);
nand U6641 (N_6641,N_5614,N_5054);
and U6642 (N_6642,N_5591,N_5895);
xnor U6643 (N_6643,N_5537,N_5303);
nor U6644 (N_6644,N_5059,N_5595);
xnor U6645 (N_6645,N_5169,N_5382);
nor U6646 (N_6646,N_5875,N_5354);
and U6647 (N_6647,N_5036,N_5246);
nor U6648 (N_6648,N_5508,N_5463);
xnor U6649 (N_6649,N_5029,N_5553);
and U6650 (N_6650,N_5139,N_5388);
xnor U6651 (N_6651,N_5521,N_5659);
nand U6652 (N_6652,N_5077,N_5790);
and U6653 (N_6653,N_5490,N_5931);
or U6654 (N_6654,N_5162,N_5183);
xnor U6655 (N_6655,N_5944,N_5793);
nand U6656 (N_6656,N_5445,N_5008);
xor U6657 (N_6657,N_5894,N_5252);
or U6658 (N_6658,N_5558,N_5666);
and U6659 (N_6659,N_5437,N_5779);
nor U6660 (N_6660,N_5975,N_5816);
nor U6661 (N_6661,N_5738,N_5882);
and U6662 (N_6662,N_5011,N_5306);
or U6663 (N_6663,N_5909,N_5607);
xor U6664 (N_6664,N_5133,N_5441);
nor U6665 (N_6665,N_5629,N_5120);
xor U6666 (N_6666,N_5820,N_5444);
xor U6667 (N_6667,N_5308,N_5060);
xor U6668 (N_6668,N_5632,N_5188);
or U6669 (N_6669,N_5085,N_5150);
nand U6670 (N_6670,N_5014,N_5892);
nand U6671 (N_6671,N_5366,N_5034);
or U6672 (N_6672,N_5798,N_5153);
xor U6673 (N_6673,N_5468,N_5071);
nor U6674 (N_6674,N_5629,N_5285);
nand U6675 (N_6675,N_5450,N_5226);
and U6676 (N_6676,N_5969,N_5300);
xnor U6677 (N_6677,N_5264,N_5518);
nor U6678 (N_6678,N_5281,N_5600);
nor U6679 (N_6679,N_5410,N_5645);
nand U6680 (N_6680,N_5133,N_5229);
and U6681 (N_6681,N_5057,N_5856);
nor U6682 (N_6682,N_5619,N_5146);
or U6683 (N_6683,N_5394,N_5095);
xor U6684 (N_6684,N_5797,N_5296);
and U6685 (N_6685,N_5168,N_5217);
xnor U6686 (N_6686,N_5102,N_5900);
nor U6687 (N_6687,N_5497,N_5548);
nand U6688 (N_6688,N_5776,N_5381);
and U6689 (N_6689,N_5257,N_5313);
nor U6690 (N_6690,N_5425,N_5599);
nand U6691 (N_6691,N_5777,N_5176);
nor U6692 (N_6692,N_5706,N_5843);
nand U6693 (N_6693,N_5055,N_5702);
xnor U6694 (N_6694,N_5204,N_5398);
or U6695 (N_6695,N_5358,N_5933);
nor U6696 (N_6696,N_5026,N_5703);
and U6697 (N_6697,N_5308,N_5877);
or U6698 (N_6698,N_5012,N_5649);
or U6699 (N_6699,N_5884,N_5103);
and U6700 (N_6700,N_5777,N_5326);
nor U6701 (N_6701,N_5895,N_5858);
or U6702 (N_6702,N_5903,N_5582);
xor U6703 (N_6703,N_5514,N_5517);
and U6704 (N_6704,N_5578,N_5292);
nand U6705 (N_6705,N_5637,N_5609);
xor U6706 (N_6706,N_5303,N_5167);
or U6707 (N_6707,N_5535,N_5536);
nand U6708 (N_6708,N_5474,N_5435);
or U6709 (N_6709,N_5171,N_5228);
and U6710 (N_6710,N_5405,N_5785);
nor U6711 (N_6711,N_5157,N_5010);
nand U6712 (N_6712,N_5984,N_5097);
and U6713 (N_6713,N_5252,N_5317);
nor U6714 (N_6714,N_5955,N_5019);
nor U6715 (N_6715,N_5800,N_5143);
and U6716 (N_6716,N_5166,N_5262);
nand U6717 (N_6717,N_5128,N_5522);
or U6718 (N_6718,N_5498,N_5214);
nand U6719 (N_6719,N_5840,N_5368);
and U6720 (N_6720,N_5295,N_5404);
nand U6721 (N_6721,N_5902,N_5255);
or U6722 (N_6722,N_5307,N_5760);
xor U6723 (N_6723,N_5765,N_5706);
or U6724 (N_6724,N_5215,N_5035);
or U6725 (N_6725,N_5700,N_5293);
or U6726 (N_6726,N_5031,N_5388);
and U6727 (N_6727,N_5950,N_5720);
or U6728 (N_6728,N_5815,N_5017);
or U6729 (N_6729,N_5271,N_5820);
xnor U6730 (N_6730,N_5542,N_5151);
nor U6731 (N_6731,N_5002,N_5140);
nand U6732 (N_6732,N_5022,N_5439);
nor U6733 (N_6733,N_5994,N_5353);
nor U6734 (N_6734,N_5937,N_5582);
and U6735 (N_6735,N_5525,N_5043);
and U6736 (N_6736,N_5581,N_5121);
or U6737 (N_6737,N_5463,N_5184);
nor U6738 (N_6738,N_5812,N_5049);
and U6739 (N_6739,N_5663,N_5854);
and U6740 (N_6740,N_5697,N_5339);
xnor U6741 (N_6741,N_5728,N_5684);
and U6742 (N_6742,N_5600,N_5593);
nand U6743 (N_6743,N_5284,N_5878);
or U6744 (N_6744,N_5976,N_5096);
and U6745 (N_6745,N_5060,N_5393);
xor U6746 (N_6746,N_5515,N_5341);
nand U6747 (N_6747,N_5611,N_5687);
and U6748 (N_6748,N_5330,N_5293);
or U6749 (N_6749,N_5430,N_5931);
and U6750 (N_6750,N_5379,N_5842);
or U6751 (N_6751,N_5879,N_5709);
and U6752 (N_6752,N_5073,N_5621);
and U6753 (N_6753,N_5023,N_5738);
nor U6754 (N_6754,N_5706,N_5183);
and U6755 (N_6755,N_5392,N_5354);
and U6756 (N_6756,N_5787,N_5623);
and U6757 (N_6757,N_5189,N_5143);
or U6758 (N_6758,N_5585,N_5408);
xnor U6759 (N_6759,N_5499,N_5373);
nor U6760 (N_6760,N_5802,N_5096);
xnor U6761 (N_6761,N_5292,N_5938);
nor U6762 (N_6762,N_5120,N_5693);
xor U6763 (N_6763,N_5538,N_5602);
nor U6764 (N_6764,N_5820,N_5258);
or U6765 (N_6765,N_5590,N_5569);
nand U6766 (N_6766,N_5287,N_5589);
or U6767 (N_6767,N_5277,N_5983);
xnor U6768 (N_6768,N_5680,N_5549);
or U6769 (N_6769,N_5088,N_5813);
xor U6770 (N_6770,N_5873,N_5425);
and U6771 (N_6771,N_5194,N_5572);
xor U6772 (N_6772,N_5276,N_5468);
and U6773 (N_6773,N_5524,N_5412);
nand U6774 (N_6774,N_5928,N_5761);
nand U6775 (N_6775,N_5043,N_5787);
or U6776 (N_6776,N_5899,N_5782);
or U6777 (N_6777,N_5560,N_5318);
and U6778 (N_6778,N_5851,N_5026);
nand U6779 (N_6779,N_5396,N_5170);
and U6780 (N_6780,N_5141,N_5679);
xnor U6781 (N_6781,N_5099,N_5460);
or U6782 (N_6782,N_5377,N_5672);
and U6783 (N_6783,N_5956,N_5414);
nand U6784 (N_6784,N_5161,N_5511);
nor U6785 (N_6785,N_5377,N_5089);
nor U6786 (N_6786,N_5949,N_5588);
or U6787 (N_6787,N_5055,N_5245);
or U6788 (N_6788,N_5814,N_5910);
or U6789 (N_6789,N_5443,N_5631);
nor U6790 (N_6790,N_5849,N_5394);
nor U6791 (N_6791,N_5803,N_5444);
or U6792 (N_6792,N_5488,N_5853);
and U6793 (N_6793,N_5074,N_5157);
nand U6794 (N_6794,N_5088,N_5083);
or U6795 (N_6795,N_5073,N_5496);
nand U6796 (N_6796,N_5935,N_5408);
or U6797 (N_6797,N_5348,N_5004);
nand U6798 (N_6798,N_5185,N_5616);
nand U6799 (N_6799,N_5065,N_5316);
or U6800 (N_6800,N_5115,N_5914);
or U6801 (N_6801,N_5649,N_5751);
or U6802 (N_6802,N_5139,N_5091);
xor U6803 (N_6803,N_5320,N_5951);
nor U6804 (N_6804,N_5360,N_5390);
and U6805 (N_6805,N_5675,N_5517);
nor U6806 (N_6806,N_5379,N_5284);
nand U6807 (N_6807,N_5521,N_5608);
xor U6808 (N_6808,N_5524,N_5022);
xnor U6809 (N_6809,N_5222,N_5771);
nor U6810 (N_6810,N_5421,N_5368);
and U6811 (N_6811,N_5169,N_5190);
or U6812 (N_6812,N_5404,N_5885);
xor U6813 (N_6813,N_5258,N_5721);
nor U6814 (N_6814,N_5483,N_5586);
nand U6815 (N_6815,N_5727,N_5635);
and U6816 (N_6816,N_5129,N_5339);
or U6817 (N_6817,N_5207,N_5923);
nor U6818 (N_6818,N_5712,N_5451);
and U6819 (N_6819,N_5407,N_5408);
xnor U6820 (N_6820,N_5558,N_5385);
nor U6821 (N_6821,N_5408,N_5905);
or U6822 (N_6822,N_5518,N_5689);
and U6823 (N_6823,N_5265,N_5855);
nor U6824 (N_6824,N_5666,N_5975);
or U6825 (N_6825,N_5595,N_5574);
and U6826 (N_6826,N_5844,N_5181);
xnor U6827 (N_6827,N_5477,N_5005);
xnor U6828 (N_6828,N_5338,N_5243);
and U6829 (N_6829,N_5149,N_5595);
xor U6830 (N_6830,N_5292,N_5186);
or U6831 (N_6831,N_5785,N_5742);
nand U6832 (N_6832,N_5891,N_5137);
xor U6833 (N_6833,N_5026,N_5128);
nor U6834 (N_6834,N_5941,N_5553);
or U6835 (N_6835,N_5307,N_5161);
nor U6836 (N_6836,N_5168,N_5444);
nand U6837 (N_6837,N_5824,N_5503);
or U6838 (N_6838,N_5568,N_5229);
xnor U6839 (N_6839,N_5417,N_5264);
or U6840 (N_6840,N_5753,N_5764);
or U6841 (N_6841,N_5089,N_5942);
or U6842 (N_6842,N_5714,N_5711);
nor U6843 (N_6843,N_5146,N_5711);
and U6844 (N_6844,N_5573,N_5747);
nand U6845 (N_6845,N_5111,N_5717);
nor U6846 (N_6846,N_5118,N_5028);
nand U6847 (N_6847,N_5967,N_5627);
xor U6848 (N_6848,N_5157,N_5885);
and U6849 (N_6849,N_5501,N_5043);
and U6850 (N_6850,N_5260,N_5006);
and U6851 (N_6851,N_5355,N_5371);
or U6852 (N_6852,N_5172,N_5914);
xor U6853 (N_6853,N_5011,N_5360);
nand U6854 (N_6854,N_5711,N_5439);
nand U6855 (N_6855,N_5718,N_5151);
xor U6856 (N_6856,N_5912,N_5062);
xnor U6857 (N_6857,N_5253,N_5480);
or U6858 (N_6858,N_5303,N_5505);
nor U6859 (N_6859,N_5323,N_5314);
and U6860 (N_6860,N_5225,N_5192);
xnor U6861 (N_6861,N_5812,N_5577);
and U6862 (N_6862,N_5792,N_5687);
nor U6863 (N_6863,N_5077,N_5389);
nand U6864 (N_6864,N_5020,N_5320);
and U6865 (N_6865,N_5847,N_5194);
nand U6866 (N_6866,N_5688,N_5548);
and U6867 (N_6867,N_5748,N_5615);
or U6868 (N_6868,N_5589,N_5405);
and U6869 (N_6869,N_5038,N_5111);
xnor U6870 (N_6870,N_5240,N_5648);
or U6871 (N_6871,N_5778,N_5800);
xnor U6872 (N_6872,N_5556,N_5694);
xnor U6873 (N_6873,N_5556,N_5434);
xnor U6874 (N_6874,N_5088,N_5613);
xor U6875 (N_6875,N_5765,N_5655);
or U6876 (N_6876,N_5520,N_5934);
or U6877 (N_6877,N_5075,N_5435);
nand U6878 (N_6878,N_5389,N_5767);
and U6879 (N_6879,N_5399,N_5254);
and U6880 (N_6880,N_5526,N_5671);
xor U6881 (N_6881,N_5150,N_5115);
nor U6882 (N_6882,N_5452,N_5334);
and U6883 (N_6883,N_5639,N_5319);
nand U6884 (N_6884,N_5594,N_5527);
nand U6885 (N_6885,N_5568,N_5071);
nand U6886 (N_6886,N_5112,N_5937);
nor U6887 (N_6887,N_5284,N_5265);
nor U6888 (N_6888,N_5465,N_5211);
nand U6889 (N_6889,N_5058,N_5083);
nand U6890 (N_6890,N_5723,N_5359);
and U6891 (N_6891,N_5674,N_5635);
or U6892 (N_6892,N_5309,N_5115);
xor U6893 (N_6893,N_5834,N_5966);
or U6894 (N_6894,N_5743,N_5376);
xnor U6895 (N_6895,N_5397,N_5569);
nor U6896 (N_6896,N_5576,N_5991);
and U6897 (N_6897,N_5472,N_5231);
or U6898 (N_6898,N_5433,N_5514);
nand U6899 (N_6899,N_5556,N_5266);
and U6900 (N_6900,N_5494,N_5268);
nor U6901 (N_6901,N_5546,N_5580);
or U6902 (N_6902,N_5968,N_5873);
xnor U6903 (N_6903,N_5670,N_5869);
xnor U6904 (N_6904,N_5181,N_5652);
or U6905 (N_6905,N_5883,N_5181);
nand U6906 (N_6906,N_5144,N_5611);
and U6907 (N_6907,N_5385,N_5124);
nor U6908 (N_6908,N_5573,N_5429);
nor U6909 (N_6909,N_5482,N_5735);
and U6910 (N_6910,N_5868,N_5522);
and U6911 (N_6911,N_5810,N_5064);
xnor U6912 (N_6912,N_5148,N_5262);
and U6913 (N_6913,N_5572,N_5970);
and U6914 (N_6914,N_5176,N_5248);
xnor U6915 (N_6915,N_5552,N_5399);
and U6916 (N_6916,N_5030,N_5003);
xor U6917 (N_6917,N_5358,N_5638);
and U6918 (N_6918,N_5728,N_5947);
and U6919 (N_6919,N_5744,N_5601);
and U6920 (N_6920,N_5493,N_5937);
nor U6921 (N_6921,N_5689,N_5575);
nand U6922 (N_6922,N_5350,N_5825);
and U6923 (N_6923,N_5184,N_5680);
nand U6924 (N_6924,N_5941,N_5242);
and U6925 (N_6925,N_5630,N_5679);
or U6926 (N_6926,N_5226,N_5788);
nand U6927 (N_6927,N_5369,N_5904);
nor U6928 (N_6928,N_5979,N_5975);
nand U6929 (N_6929,N_5968,N_5475);
or U6930 (N_6930,N_5416,N_5853);
nor U6931 (N_6931,N_5902,N_5865);
or U6932 (N_6932,N_5994,N_5852);
and U6933 (N_6933,N_5948,N_5281);
or U6934 (N_6934,N_5591,N_5631);
xor U6935 (N_6935,N_5144,N_5127);
and U6936 (N_6936,N_5846,N_5585);
or U6937 (N_6937,N_5024,N_5460);
and U6938 (N_6938,N_5926,N_5802);
nor U6939 (N_6939,N_5034,N_5142);
nor U6940 (N_6940,N_5465,N_5651);
or U6941 (N_6941,N_5369,N_5579);
nor U6942 (N_6942,N_5148,N_5695);
xnor U6943 (N_6943,N_5379,N_5484);
nand U6944 (N_6944,N_5816,N_5644);
and U6945 (N_6945,N_5519,N_5239);
and U6946 (N_6946,N_5541,N_5257);
nand U6947 (N_6947,N_5941,N_5664);
or U6948 (N_6948,N_5354,N_5640);
and U6949 (N_6949,N_5628,N_5744);
and U6950 (N_6950,N_5589,N_5874);
nand U6951 (N_6951,N_5234,N_5471);
nor U6952 (N_6952,N_5774,N_5279);
xnor U6953 (N_6953,N_5801,N_5849);
nand U6954 (N_6954,N_5440,N_5569);
and U6955 (N_6955,N_5358,N_5701);
xor U6956 (N_6956,N_5342,N_5541);
xnor U6957 (N_6957,N_5047,N_5749);
nand U6958 (N_6958,N_5942,N_5190);
xor U6959 (N_6959,N_5461,N_5591);
nor U6960 (N_6960,N_5875,N_5467);
nor U6961 (N_6961,N_5050,N_5059);
nor U6962 (N_6962,N_5889,N_5263);
and U6963 (N_6963,N_5703,N_5859);
xnor U6964 (N_6964,N_5538,N_5927);
and U6965 (N_6965,N_5532,N_5646);
nand U6966 (N_6966,N_5514,N_5223);
nand U6967 (N_6967,N_5627,N_5974);
xnor U6968 (N_6968,N_5942,N_5772);
and U6969 (N_6969,N_5884,N_5583);
xor U6970 (N_6970,N_5536,N_5862);
xor U6971 (N_6971,N_5181,N_5691);
xnor U6972 (N_6972,N_5115,N_5916);
nand U6973 (N_6973,N_5211,N_5554);
nor U6974 (N_6974,N_5350,N_5411);
xnor U6975 (N_6975,N_5442,N_5115);
nor U6976 (N_6976,N_5196,N_5415);
nand U6977 (N_6977,N_5988,N_5048);
and U6978 (N_6978,N_5712,N_5277);
and U6979 (N_6979,N_5300,N_5914);
nor U6980 (N_6980,N_5379,N_5270);
nand U6981 (N_6981,N_5957,N_5408);
nor U6982 (N_6982,N_5212,N_5573);
and U6983 (N_6983,N_5161,N_5717);
nor U6984 (N_6984,N_5680,N_5331);
or U6985 (N_6985,N_5789,N_5330);
or U6986 (N_6986,N_5026,N_5481);
nor U6987 (N_6987,N_5064,N_5946);
xnor U6988 (N_6988,N_5321,N_5495);
nor U6989 (N_6989,N_5327,N_5503);
xnor U6990 (N_6990,N_5579,N_5238);
nor U6991 (N_6991,N_5087,N_5123);
nor U6992 (N_6992,N_5589,N_5233);
xor U6993 (N_6993,N_5154,N_5170);
nor U6994 (N_6994,N_5594,N_5243);
nor U6995 (N_6995,N_5928,N_5130);
nor U6996 (N_6996,N_5014,N_5267);
and U6997 (N_6997,N_5656,N_5525);
or U6998 (N_6998,N_5305,N_5125);
or U6999 (N_6999,N_5438,N_5866);
nor U7000 (N_7000,N_6918,N_6550);
nor U7001 (N_7001,N_6456,N_6050);
nand U7002 (N_7002,N_6540,N_6816);
or U7003 (N_7003,N_6254,N_6577);
xnor U7004 (N_7004,N_6804,N_6064);
xor U7005 (N_7005,N_6009,N_6093);
and U7006 (N_7006,N_6886,N_6291);
and U7007 (N_7007,N_6973,N_6857);
xnor U7008 (N_7008,N_6705,N_6891);
and U7009 (N_7009,N_6987,N_6028);
nor U7010 (N_7010,N_6189,N_6237);
nand U7011 (N_7011,N_6429,N_6232);
and U7012 (N_7012,N_6083,N_6689);
xor U7013 (N_7013,N_6764,N_6929);
or U7014 (N_7014,N_6304,N_6440);
nor U7015 (N_7015,N_6067,N_6605);
nor U7016 (N_7016,N_6353,N_6066);
nand U7017 (N_7017,N_6297,N_6059);
nor U7018 (N_7018,N_6972,N_6259);
nand U7019 (N_7019,N_6840,N_6514);
and U7020 (N_7020,N_6613,N_6938);
and U7021 (N_7021,N_6212,N_6681);
or U7022 (N_7022,N_6343,N_6846);
or U7023 (N_7023,N_6503,N_6906);
and U7024 (N_7024,N_6685,N_6608);
nor U7025 (N_7025,N_6321,N_6601);
xor U7026 (N_7026,N_6921,N_6867);
nor U7027 (N_7027,N_6197,N_6172);
or U7028 (N_7028,N_6024,N_6096);
or U7029 (N_7029,N_6777,N_6900);
and U7030 (N_7030,N_6757,N_6570);
or U7031 (N_7031,N_6080,N_6358);
or U7032 (N_7032,N_6731,N_6247);
and U7033 (N_7033,N_6650,N_6626);
nand U7034 (N_7034,N_6467,N_6325);
nor U7035 (N_7035,N_6296,N_6274);
nor U7036 (N_7036,N_6183,N_6854);
nor U7037 (N_7037,N_6193,N_6371);
xor U7038 (N_7038,N_6349,N_6547);
nor U7039 (N_7039,N_6801,N_6229);
nor U7040 (N_7040,N_6653,N_6436);
and U7041 (N_7041,N_6627,N_6907);
or U7042 (N_7042,N_6847,N_6497);
and U7043 (N_7043,N_6470,N_6735);
nor U7044 (N_7044,N_6622,N_6251);
xor U7045 (N_7045,N_6078,N_6772);
nand U7046 (N_7046,N_6831,N_6179);
nor U7047 (N_7047,N_6134,N_6961);
nor U7048 (N_7048,N_6173,N_6228);
xor U7049 (N_7049,N_6217,N_6563);
or U7050 (N_7050,N_6658,N_6700);
xor U7051 (N_7051,N_6925,N_6088);
nand U7052 (N_7052,N_6270,N_6382);
nand U7053 (N_7053,N_6344,N_6649);
and U7054 (N_7054,N_6401,N_6030);
nor U7055 (N_7055,N_6460,N_6094);
nand U7056 (N_7056,N_6486,N_6779);
and U7057 (N_7057,N_6124,N_6184);
and U7058 (N_7058,N_6359,N_6977);
nand U7059 (N_7059,N_6282,N_6071);
and U7060 (N_7060,N_6937,N_6081);
nand U7061 (N_7061,N_6654,N_6129);
and U7062 (N_7062,N_6722,N_6679);
or U7063 (N_7063,N_6375,N_6374);
nor U7064 (N_7064,N_6712,N_6288);
nand U7065 (N_7065,N_6231,N_6018);
and U7066 (N_7066,N_6742,N_6219);
xnor U7067 (N_7067,N_6781,N_6706);
or U7068 (N_7068,N_6607,N_6493);
and U7069 (N_7069,N_6561,N_6388);
nand U7070 (N_7070,N_6967,N_6277);
and U7071 (N_7071,N_6048,N_6453);
nor U7072 (N_7072,N_6373,N_6116);
nor U7073 (N_7073,N_6910,N_6533);
or U7074 (N_7074,N_6552,N_6487);
xor U7075 (N_7075,N_6743,N_6639);
and U7076 (N_7076,N_6203,N_6719);
nand U7077 (N_7077,N_6438,N_6598);
nor U7078 (N_7078,N_6174,N_6889);
and U7079 (N_7079,N_6959,N_6146);
nand U7080 (N_7080,N_6704,N_6955);
nand U7081 (N_7081,N_6152,N_6465);
xor U7082 (N_7082,N_6452,N_6348);
and U7083 (N_7083,N_6749,N_6796);
xnor U7084 (N_7084,N_6562,N_6167);
and U7085 (N_7085,N_6079,N_6095);
nor U7086 (N_7086,N_6943,N_6113);
and U7087 (N_7087,N_6769,N_6138);
xnor U7088 (N_7088,N_6107,N_6346);
xnor U7089 (N_7089,N_6481,N_6188);
nor U7090 (N_7090,N_6862,N_6790);
xor U7091 (N_7091,N_6177,N_6507);
xor U7092 (N_7092,N_6441,N_6058);
nor U7093 (N_7093,N_6306,N_6210);
xor U7094 (N_7094,N_6125,N_6870);
xnor U7095 (N_7095,N_6133,N_6301);
or U7096 (N_7096,N_6170,N_6276);
nor U7097 (N_7097,N_6407,N_6397);
xor U7098 (N_7098,N_6400,N_6157);
nor U7099 (N_7099,N_6462,N_6569);
and U7100 (N_7100,N_6839,N_6670);
and U7101 (N_7101,N_6333,N_6978);
nor U7102 (N_7102,N_6115,N_6912);
and U7103 (N_7103,N_6086,N_6084);
nand U7104 (N_7104,N_6750,N_6357);
nand U7105 (N_7105,N_6335,N_6305);
or U7106 (N_7106,N_6310,N_6381);
and U7107 (N_7107,N_6230,N_6338);
and U7108 (N_7108,N_6621,N_6027);
and U7109 (N_7109,N_6222,N_6711);
nand U7110 (N_7110,N_6329,N_6892);
and U7111 (N_7111,N_6826,N_6494);
or U7112 (N_7112,N_6145,N_6238);
or U7113 (N_7113,N_6383,N_6814);
xnor U7114 (N_7114,N_6198,N_6868);
xnor U7115 (N_7115,N_6039,N_6884);
or U7116 (N_7116,N_6015,N_6594);
xor U7117 (N_7117,N_6426,N_6005);
nand U7118 (N_7118,N_6127,N_6524);
xor U7119 (N_7119,N_6308,N_6240);
or U7120 (N_7120,N_6845,N_6806);
or U7121 (N_7121,N_6336,N_6614);
or U7122 (N_7122,N_6774,N_6794);
xnor U7123 (N_7123,N_6327,N_6528);
or U7124 (N_7124,N_6140,N_6418);
xor U7125 (N_7125,N_6758,N_6913);
or U7126 (N_7126,N_6454,N_6994);
and U7127 (N_7127,N_6459,N_6788);
nand U7128 (N_7128,N_6683,N_6474);
xor U7129 (N_7129,N_6733,N_6047);
xnor U7130 (N_7130,N_6098,N_6223);
nand U7131 (N_7131,N_6644,N_6315);
xnor U7132 (N_7132,N_6647,N_6444);
nor U7133 (N_7133,N_6478,N_6019);
or U7134 (N_7134,N_6110,N_6390);
nor U7135 (N_7135,N_6693,N_6392);
nand U7136 (N_7136,N_6143,N_6076);
nand U7137 (N_7137,N_6554,N_6490);
or U7138 (N_7138,N_6879,N_6933);
nand U7139 (N_7139,N_6661,N_6126);
and U7140 (N_7140,N_6620,N_6775);
xnor U7141 (N_7141,N_6021,N_6283);
nand U7142 (N_7142,N_6285,N_6334);
and U7143 (N_7143,N_6897,N_6419);
nand U7144 (N_7144,N_6461,N_6155);
or U7145 (N_7145,N_6160,N_6885);
nor U7146 (N_7146,N_6182,N_6952);
nor U7147 (N_7147,N_6549,N_6730);
or U7148 (N_7148,N_6209,N_6166);
and U7149 (N_7149,N_6196,N_6337);
nor U7150 (N_7150,N_6851,N_6416);
xor U7151 (N_7151,N_6709,N_6101);
nand U7152 (N_7152,N_6887,N_6350);
and U7153 (N_7153,N_6842,N_6384);
nor U7154 (N_7154,N_6111,N_6855);
or U7155 (N_7155,N_6164,N_6703);
nor U7156 (N_7156,N_6114,N_6150);
nor U7157 (N_7157,N_6515,N_6686);
or U7158 (N_7158,N_6206,N_6746);
or U7159 (N_7159,N_6587,N_6936);
xnor U7160 (N_7160,N_6828,N_6163);
nand U7161 (N_7161,N_6142,N_6483);
nand U7162 (N_7162,N_6819,N_6655);
or U7163 (N_7163,N_6762,N_6010);
nor U7164 (N_7164,N_6511,N_6850);
nand U7165 (N_7165,N_6396,N_6723);
nand U7166 (N_7166,N_6941,N_6108);
xnor U7167 (N_7167,N_6829,N_6032);
nand U7168 (N_7168,N_6034,N_6556);
nand U7169 (N_7169,N_6603,N_6187);
and U7170 (N_7170,N_6966,N_6249);
nand U7171 (N_7171,N_6747,N_6836);
nand U7172 (N_7172,N_6417,N_6871);
nor U7173 (N_7173,N_6070,N_6023);
xnor U7174 (N_7174,N_6506,N_6105);
nand U7175 (N_7175,N_6753,N_6378);
xnor U7176 (N_7176,N_6932,N_6861);
nor U7177 (N_7177,N_6199,N_6476);
xnor U7178 (N_7178,N_6568,N_6776);
or U7179 (N_7179,N_6011,N_6963);
nor U7180 (N_7180,N_6428,N_6602);
or U7181 (N_7181,N_6256,N_6266);
and U7182 (N_7182,N_6771,N_6741);
nand U7183 (N_7183,N_6944,N_6218);
nor U7184 (N_7184,N_6555,N_6402);
nor U7185 (N_7185,N_6089,N_6437);
nor U7186 (N_7186,N_6737,N_6983);
xor U7187 (N_7187,N_6948,N_6817);
and U7188 (N_7188,N_6877,N_6038);
nor U7189 (N_7189,N_6328,N_6962);
or U7190 (N_7190,N_6387,N_6702);
xor U7191 (N_7191,N_6643,N_6997);
nor U7192 (N_7192,N_6340,N_6158);
xor U7193 (N_7193,N_6097,N_6379);
xnor U7194 (N_7194,N_6539,N_6376);
and U7195 (N_7195,N_6976,N_6236);
nor U7196 (N_7196,N_6899,N_6316);
or U7197 (N_7197,N_6300,N_6457);
nor U7198 (N_7198,N_6181,N_6606);
nor U7199 (N_7199,N_6389,N_6707);
and U7200 (N_7200,N_6745,N_6638);
or U7201 (N_7201,N_6482,N_6235);
nand U7202 (N_7202,N_6245,N_6045);
nor U7203 (N_7203,N_6927,N_6754);
xor U7204 (N_7204,N_6420,N_6572);
or U7205 (N_7205,N_6560,N_6341);
or U7206 (N_7206,N_6536,N_6354);
and U7207 (N_7207,N_6433,N_6502);
nor U7208 (N_7208,N_6455,N_6844);
xnor U7209 (N_7209,N_6701,N_6551);
and U7210 (N_7210,N_6380,N_6789);
nand U7211 (N_7211,N_6248,N_6424);
xor U7212 (N_7212,N_6736,N_6399);
or U7213 (N_7213,N_6557,N_6633);
and U7214 (N_7214,N_6006,N_6975);
xor U7215 (N_7215,N_6782,N_6610);
xnor U7216 (N_7216,N_6153,N_6118);
xnor U7217 (N_7217,N_6532,N_6489);
nor U7218 (N_7218,N_6545,N_6136);
nor U7219 (N_7219,N_6284,N_6319);
nor U7220 (N_7220,N_6403,N_6544);
nand U7221 (N_7221,N_6599,N_6148);
nand U7222 (N_7222,N_6268,N_6641);
nand U7223 (N_7223,N_6596,N_6538);
nand U7224 (N_7224,N_6186,N_6950);
nor U7225 (N_7225,N_6054,N_6720);
and U7226 (N_7226,N_6660,N_6964);
xor U7227 (N_7227,N_6372,N_6109);
xor U7228 (N_7228,N_6629,N_6185);
xor U7229 (N_7229,N_6527,N_6667);
nor U7230 (N_7230,N_6953,N_6293);
and U7231 (N_7231,N_6911,N_6675);
xor U7232 (N_7232,N_6290,N_6810);
and U7233 (N_7233,N_6793,N_6471);
nand U7234 (N_7234,N_6016,N_6149);
nand U7235 (N_7235,N_6046,N_6202);
nand U7236 (N_7236,N_6980,N_6864);
and U7237 (N_7237,N_6904,N_6082);
xor U7238 (N_7238,N_6221,N_6242);
and U7239 (N_7239,N_6991,N_6044);
nor U7240 (N_7240,N_6154,N_6677);
nand U7241 (N_7241,N_6201,N_6585);
nor U7242 (N_7242,N_6224,N_6865);
nor U7243 (N_7243,N_6216,N_6664);
nand U7244 (N_7244,N_6367,N_6852);
xnor U7245 (N_7245,N_6824,N_6791);
or U7246 (N_7246,N_6571,N_6169);
or U7247 (N_7247,N_6207,N_6922);
xnor U7248 (N_7248,N_6908,N_6843);
nor U7249 (N_7249,N_6473,N_6993);
and U7250 (N_7250,N_6968,N_6979);
or U7251 (N_7251,N_6631,N_6519);
or U7252 (N_7252,N_6965,N_6175);
nor U7253 (N_7253,N_6355,N_6500);
xor U7254 (N_7254,N_6671,N_6513);
xnor U7255 (N_7255,N_6106,N_6688);
and U7256 (N_7256,N_6752,N_6618);
nor U7257 (N_7257,N_6074,N_6909);
nor U7258 (N_7258,N_6313,N_6530);
and U7259 (N_7259,N_6208,N_6104);
xnor U7260 (N_7260,N_6986,N_6567);
or U7261 (N_7261,N_6595,N_6008);
xnor U7262 (N_7262,N_6541,N_6930);
and U7263 (N_7263,N_6312,N_6065);
xor U7264 (N_7264,N_6682,N_6326);
and U7265 (N_7265,N_6529,N_6255);
and U7266 (N_7266,N_6499,N_6299);
or U7267 (N_7267,N_6468,N_6989);
and U7268 (N_7268,N_6784,N_6858);
xor U7269 (N_7269,N_6404,N_6369);
nor U7270 (N_7270,N_6652,N_6510);
or U7271 (N_7271,N_6269,N_6820);
and U7272 (N_7272,N_6443,N_6729);
nor U7273 (N_7273,N_6063,N_6368);
nand U7274 (N_7274,N_6496,N_6171);
or U7275 (N_7275,N_6841,N_6564);
and U7276 (N_7276,N_6365,N_6194);
nor U7277 (N_7277,N_6739,N_6036);
or U7278 (N_7278,N_6676,N_6425);
nand U7279 (N_7279,N_6002,N_6838);
nand U7280 (N_7280,N_6559,N_6225);
or U7281 (N_7281,N_6518,N_6120);
xor U7282 (N_7282,N_6874,N_6756);
or U7283 (N_7283,N_6581,N_6331);
nor U7284 (N_7284,N_6025,N_6665);
and U7285 (N_7285,N_6984,N_6226);
nand U7286 (N_7286,N_6694,N_6122);
and U7287 (N_7287,N_6439,N_6708);
nor U7288 (N_7288,N_6220,N_6013);
nand U7289 (N_7289,N_6695,N_6684);
nand U7290 (N_7290,N_6588,N_6717);
xor U7291 (N_7291,N_6636,N_6940);
nand U7292 (N_7292,N_6697,N_6692);
nor U7293 (N_7293,N_6345,N_6673);
or U7294 (N_7294,N_6783,N_6928);
nor U7295 (N_7295,N_6060,N_6413);
xor U7296 (N_7296,N_6446,N_6713);
or U7297 (N_7297,N_6632,N_6258);
and U7298 (N_7298,N_6159,N_6130);
and U7299 (N_7299,N_6935,N_6651);
xor U7300 (N_7300,N_6330,N_6077);
xor U7301 (N_7301,N_6469,N_6286);
nand U7302 (N_7302,N_6022,N_6916);
and U7303 (N_7303,N_6017,N_6934);
xor U7304 (N_7304,N_6195,N_6488);
and U7305 (N_7305,N_6766,N_6591);
or U7306 (N_7306,N_6798,N_6100);
or U7307 (N_7307,N_6263,N_6875);
nand U7308 (N_7308,N_6464,N_6640);
and U7309 (N_7309,N_6778,N_6718);
xnor U7310 (N_7310,N_6165,N_6479);
nor U7311 (N_7311,N_6053,N_6893);
and U7312 (N_7312,N_6725,N_6099);
nor U7313 (N_7313,N_6135,N_6289);
or U7314 (N_7314,N_6119,N_6128);
or U7315 (N_7315,N_6951,N_6947);
xnor U7316 (N_7316,N_6033,N_6190);
nor U7317 (N_7317,N_6307,N_6813);
xnor U7318 (N_7318,N_6537,N_6690);
xnor U7319 (N_7319,N_6821,N_6516);
nand U7320 (N_7320,N_6770,N_6003);
or U7321 (N_7321,N_6012,N_6575);
xor U7322 (N_7322,N_6168,N_6734);
xnor U7323 (N_7323,N_6767,N_6721);
nand U7324 (N_7324,N_6659,N_6205);
xor U7325 (N_7325,N_6147,N_6833);
nand U7326 (N_7326,N_6565,N_6410);
and U7327 (N_7327,N_6257,N_6409);
xnor U7328 (N_7328,N_6139,N_6710);
nor U7329 (N_7329,N_6141,N_6797);
or U7330 (N_7330,N_6637,N_6615);
and U7331 (N_7331,N_6026,N_6648);
nand U7332 (N_7332,N_6415,N_6020);
and U7333 (N_7333,N_6303,N_6377);
and U7334 (N_7334,N_6763,N_6969);
nand U7335 (N_7335,N_6272,N_6795);
and U7336 (N_7336,N_6787,N_6834);
xor U7337 (N_7337,N_6458,N_6475);
nor U7338 (N_7338,N_6958,N_6069);
xnor U7339 (N_7339,N_6342,N_6748);
xor U7340 (N_7340,N_6818,N_6724);
and U7341 (N_7341,N_6498,N_6432);
nand U7342 (N_7342,N_6830,N_6589);
nor U7343 (N_7343,N_6522,N_6508);
nand U7344 (N_7344,N_6759,N_6981);
or U7345 (N_7345,N_6954,N_6619);
nand U7346 (N_7346,N_6740,N_6996);
and U7347 (N_7347,N_6714,N_6234);
nor U7348 (N_7348,N_6394,N_6414);
xor U7349 (N_7349,N_6663,N_6121);
nand U7350 (N_7350,N_6674,N_6395);
nor U7351 (N_7351,N_6662,N_6043);
or U7352 (N_7352,N_6896,N_6520);
nor U7353 (N_7353,N_6447,N_6227);
nor U7354 (N_7354,N_6592,N_6573);
xor U7355 (N_7355,N_6137,N_6617);
nand U7356 (N_7356,N_6815,N_6999);
xor U7357 (N_7357,N_6347,N_6728);
nand U7358 (N_7358,N_6322,N_6785);
or U7359 (N_7359,N_6241,N_6584);
or U7360 (N_7360,N_6878,N_6988);
nor U7361 (N_7361,N_6485,N_6422);
or U7362 (N_7362,N_6691,N_6273);
and U7363 (N_7363,N_6985,N_6837);
xor U7364 (N_7364,N_6768,N_6042);
xor U7365 (N_7365,N_6324,N_6656);
xor U7366 (N_7366,N_6931,N_6657);
xnor U7367 (N_7367,N_6761,N_6872);
xnor U7368 (N_7368,N_6760,N_6809);
nor U7369 (N_7369,N_6668,N_6052);
or U7370 (N_7370,N_6463,N_6523);
xnor U7371 (N_7371,N_6477,N_6176);
or U7372 (N_7372,N_6856,N_6903);
nor U7373 (N_7373,N_6244,N_6509);
nand U7374 (N_7374,N_6253,N_6939);
and U7375 (N_7375,N_6616,N_6412);
and U7376 (N_7376,N_6888,N_6822);
and U7377 (N_7377,N_6215,N_6370);
nor U7378 (N_7378,N_6505,N_6957);
xor U7379 (N_7379,N_6430,N_6037);
nand U7380 (N_7380,N_6192,N_6534);
and U7381 (N_7381,N_6901,N_6531);
nand U7382 (N_7382,N_6512,N_6895);
nor U7383 (N_7383,N_6243,N_6558);
xnor U7384 (N_7384,N_6480,N_6068);
and U7385 (N_7385,N_6881,N_6261);
xor U7386 (N_7386,N_6687,N_6214);
and U7387 (N_7387,N_6323,N_6678);
or U7388 (N_7388,N_6859,N_6612);
and U7389 (N_7389,N_6727,N_6501);
or U7390 (N_7390,N_6451,N_6029);
nor U7391 (N_7391,N_6309,N_6213);
nor U7392 (N_7392,N_6366,N_6521);
or U7393 (N_7393,N_6073,N_6211);
nand U7394 (N_7394,N_6200,N_6869);
nand U7395 (N_7395,N_6574,N_6860);
or U7396 (N_7396,N_6298,N_6204);
xnor U7397 (N_7397,N_6880,N_6974);
or U7398 (N_7398,N_6287,N_6435);
and U7399 (N_7399,N_6112,N_6628);
nor U7400 (N_7400,N_6352,N_6669);
and U7401 (N_7401,N_6882,N_6905);
or U7402 (N_7402,N_6442,N_6807);
nor U7403 (N_7403,N_6385,N_6604);
or U7404 (N_7404,N_6946,N_6252);
or U7405 (N_7405,N_6295,N_6582);
nand U7406 (N_7406,N_6041,N_6262);
xor U7407 (N_7407,N_6630,N_6902);
nor U7408 (N_7408,N_6960,N_6265);
nor U7409 (N_7409,N_6040,N_6281);
nand U7410 (N_7410,N_6000,N_6472);
nand U7411 (N_7411,N_6786,N_6623);
nand U7412 (N_7412,N_6386,N_6625);
xor U7413 (N_7413,N_6853,N_6876);
xnor U7414 (N_7414,N_6866,N_6680);
nand U7415 (N_7415,N_6449,N_6131);
xor U7416 (N_7416,N_6696,N_6360);
nor U7417 (N_7417,N_6586,N_6590);
or U7418 (N_7418,N_6998,N_6491);
nand U7419 (N_7419,N_6624,N_6666);
nand U7420 (N_7420,N_6593,N_6191);
nand U7421 (N_7421,N_6546,N_6780);
nand U7422 (N_7422,N_6362,N_6970);
xor U7423 (N_7423,N_6332,N_6848);
nand U7424 (N_7424,N_6279,N_6364);
and U7425 (N_7425,N_6583,N_6090);
nand U7426 (N_7426,N_6091,N_6863);
or U7427 (N_7427,N_6835,N_6317);
and U7428 (N_7428,N_6894,N_6945);
xnor U7429 (N_7429,N_6151,N_6103);
xnor U7430 (N_7430,N_6949,N_6393);
and U7431 (N_7431,N_6832,N_6635);
and U7432 (N_7432,N_6014,N_6314);
nor U7433 (N_7433,N_6525,N_6578);
xnor U7434 (N_7434,N_6492,N_6576);
nor U7435 (N_7435,N_6007,N_6812);
nor U7436 (N_7436,N_6102,N_6356);
and U7437 (N_7437,N_6264,N_6406);
xor U7438 (N_7438,N_6411,N_6873);
nand U7439 (N_7439,N_6363,N_6239);
nand U7440 (N_7440,N_6178,N_6072);
or U7441 (N_7441,N_6942,N_6318);
or U7442 (N_7442,N_6914,N_6956);
nor U7443 (N_7443,N_6805,N_6075);
xor U7444 (N_7444,N_6004,N_6092);
nor U7445 (N_7445,N_6808,N_6995);
or U7446 (N_7446,N_6926,N_6611);
nor U7447 (N_7447,N_6275,N_6517);
and U7448 (N_7448,N_6755,N_6971);
nand U7449 (N_7449,N_6280,N_6504);
or U7450 (N_7450,N_6543,N_6448);
nor U7451 (N_7451,N_6117,N_6799);
or U7452 (N_7452,N_6278,N_6823);
and U7453 (N_7453,N_6919,N_6699);
and U7454 (N_7454,N_6716,N_6542);
nor U7455 (N_7455,N_6405,N_6920);
nand U7456 (N_7456,N_6566,N_6246);
or U7457 (N_7457,N_6849,N_6982);
nor U7458 (N_7458,N_6634,N_6398);
nor U7459 (N_7459,N_6535,N_6579);
nor U7460 (N_7460,N_6051,N_6738);
and U7461 (N_7461,N_6898,N_6434);
xor U7462 (N_7462,N_6597,N_6267);
and U7463 (N_7463,N_6990,N_6883);
or U7464 (N_7464,N_6645,N_6495);
xor U7465 (N_7465,N_6423,N_6055);
nand U7466 (N_7466,N_6726,N_6803);
xor U7467 (N_7467,N_6445,N_6123);
and U7468 (N_7468,N_6890,N_6087);
or U7469 (N_7469,N_6271,N_6061);
nand U7470 (N_7470,N_6292,N_6132);
nand U7471 (N_7471,N_6001,N_6031);
and U7472 (N_7472,N_6320,N_6351);
or U7473 (N_7473,N_6162,N_6361);
or U7474 (N_7474,N_6732,N_6915);
or U7475 (N_7475,N_6156,N_6773);
or U7476 (N_7476,N_6744,N_6311);
nor U7477 (N_7477,N_6765,N_6825);
or U7478 (N_7478,N_6580,N_6827);
nor U7479 (N_7479,N_6923,N_6924);
or U7480 (N_7480,N_6466,N_6035);
nor U7481 (N_7481,N_6715,N_6917);
and U7482 (N_7482,N_6600,N_6339);
or U7483 (N_7483,N_6294,N_6260);
xor U7484 (N_7484,N_6427,N_6144);
xnor U7485 (N_7485,N_6161,N_6800);
xnor U7486 (N_7486,N_6698,N_6751);
nor U7487 (N_7487,N_6421,N_6062);
and U7488 (N_7488,N_6672,N_6085);
or U7489 (N_7489,N_6548,N_6408);
or U7490 (N_7490,N_6233,N_6302);
nor U7491 (N_7491,N_6646,N_6484);
or U7492 (N_7492,N_6250,N_6391);
and U7493 (N_7493,N_6049,N_6057);
and U7494 (N_7494,N_6180,N_6642);
nand U7495 (N_7495,N_6450,N_6609);
nor U7496 (N_7496,N_6553,N_6811);
nor U7497 (N_7497,N_6802,N_6431);
nor U7498 (N_7498,N_6526,N_6792);
nor U7499 (N_7499,N_6056,N_6992);
nor U7500 (N_7500,N_6960,N_6617);
nand U7501 (N_7501,N_6443,N_6897);
or U7502 (N_7502,N_6573,N_6001);
nand U7503 (N_7503,N_6739,N_6851);
nor U7504 (N_7504,N_6627,N_6776);
xor U7505 (N_7505,N_6676,N_6801);
and U7506 (N_7506,N_6989,N_6097);
xnor U7507 (N_7507,N_6898,N_6063);
nand U7508 (N_7508,N_6955,N_6081);
xor U7509 (N_7509,N_6949,N_6137);
and U7510 (N_7510,N_6318,N_6745);
and U7511 (N_7511,N_6953,N_6490);
nor U7512 (N_7512,N_6849,N_6622);
nand U7513 (N_7513,N_6712,N_6035);
or U7514 (N_7514,N_6536,N_6391);
nand U7515 (N_7515,N_6046,N_6438);
xnor U7516 (N_7516,N_6274,N_6481);
xor U7517 (N_7517,N_6301,N_6880);
nor U7518 (N_7518,N_6503,N_6276);
or U7519 (N_7519,N_6715,N_6005);
and U7520 (N_7520,N_6867,N_6334);
or U7521 (N_7521,N_6001,N_6729);
nand U7522 (N_7522,N_6164,N_6707);
and U7523 (N_7523,N_6028,N_6312);
nor U7524 (N_7524,N_6553,N_6450);
and U7525 (N_7525,N_6286,N_6792);
and U7526 (N_7526,N_6202,N_6282);
or U7527 (N_7527,N_6466,N_6584);
nand U7528 (N_7528,N_6836,N_6703);
nand U7529 (N_7529,N_6873,N_6017);
xnor U7530 (N_7530,N_6499,N_6114);
and U7531 (N_7531,N_6058,N_6075);
nor U7532 (N_7532,N_6566,N_6360);
or U7533 (N_7533,N_6938,N_6707);
or U7534 (N_7534,N_6935,N_6918);
nand U7535 (N_7535,N_6773,N_6857);
or U7536 (N_7536,N_6686,N_6450);
and U7537 (N_7537,N_6381,N_6425);
or U7538 (N_7538,N_6683,N_6581);
or U7539 (N_7539,N_6667,N_6447);
or U7540 (N_7540,N_6761,N_6255);
xnor U7541 (N_7541,N_6603,N_6370);
xor U7542 (N_7542,N_6681,N_6277);
xnor U7543 (N_7543,N_6307,N_6150);
and U7544 (N_7544,N_6566,N_6839);
and U7545 (N_7545,N_6331,N_6683);
nand U7546 (N_7546,N_6502,N_6890);
nor U7547 (N_7547,N_6685,N_6978);
nand U7548 (N_7548,N_6671,N_6227);
and U7549 (N_7549,N_6350,N_6827);
and U7550 (N_7550,N_6692,N_6810);
or U7551 (N_7551,N_6720,N_6347);
or U7552 (N_7552,N_6775,N_6481);
or U7553 (N_7553,N_6054,N_6048);
nand U7554 (N_7554,N_6078,N_6172);
nand U7555 (N_7555,N_6809,N_6026);
xor U7556 (N_7556,N_6744,N_6997);
or U7557 (N_7557,N_6679,N_6058);
or U7558 (N_7558,N_6681,N_6367);
xnor U7559 (N_7559,N_6563,N_6983);
and U7560 (N_7560,N_6597,N_6246);
and U7561 (N_7561,N_6970,N_6693);
nand U7562 (N_7562,N_6493,N_6275);
and U7563 (N_7563,N_6592,N_6758);
or U7564 (N_7564,N_6610,N_6822);
nand U7565 (N_7565,N_6276,N_6090);
or U7566 (N_7566,N_6932,N_6789);
nor U7567 (N_7567,N_6137,N_6052);
nor U7568 (N_7568,N_6648,N_6907);
or U7569 (N_7569,N_6292,N_6623);
and U7570 (N_7570,N_6032,N_6052);
xnor U7571 (N_7571,N_6472,N_6621);
xor U7572 (N_7572,N_6233,N_6670);
nor U7573 (N_7573,N_6595,N_6618);
xor U7574 (N_7574,N_6813,N_6157);
nand U7575 (N_7575,N_6489,N_6315);
nor U7576 (N_7576,N_6199,N_6263);
and U7577 (N_7577,N_6086,N_6671);
or U7578 (N_7578,N_6967,N_6951);
or U7579 (N_7579,N_6407,N_6239);
nor U7580 (N_7580,N_6234,N_6822);
nor U7581 (N_7581,N_6206,N_6597);
and U7582 (N_7582,N_6107,N_6088);
or U7583 (N_7583,N_6148,N_6927);
nor U7584 (N_7584,N_6845,N_6149);
xor U7585 (N_7585,N_6968,N_6425);
nand U7586 (N_7586,N_6448,N_6628);
nand U7587 (N_7587,N_6659,N_6106);
nand U7588 (N_7588,N_6782,N_6066);
nand U7589 (N_7589,N_6523,N_6512);
nor U7590 (N_7590,N_6858,N_6844);
nor U7591 (N_7591,N_6831,N_6057);
or U7592 (N_7592,N_6301,N_6644);
or U7593 (N_7593,N_6714,N_6711);
nor U7594 (N_7594,N_6404,N_6383);
nor U7595 (N_7595,N_6637,N_6685);
nor U7596 (N_7596,N_6811,N_6286);
xor U7597 (N_7597,N_6457,N_6199);
and U7598 (N_7598,N_6928,N_6412);
nand U7599 (N_7599,N_6879,N_6289);
nand U7600 (N_7600,N_6593,N_6086);
and U7601 (N_7601,N_6667,N_6432);
and U7602 (N_7602,N_6765,N_6995);
or U7603 (N_7603,N_6567,N_6605);
nand U7604 (N_7604,N_6743,N_6769);
nand U7605 (N_7605,N_6920,N_6192);
nor U7606 (N_7606,N_6113,N_6518);
and U7607 (N_7607,N_6516,N_6524);
nor U7608 (N_7608,N_6524,N_6343);
or U7609 (N_7609,N_6269,N_6649);
and U7610 (N_7610,N_6896,N_6641);
and U7611 (N_7611,N_6659,N_6604);
nand U7612 (N_7612,N_6050,N_6382);
nor U7613 (N_7613,N_6653,N_6505);
and U7614 (N_7614,N_6455,N_6261);
xnor U7615 (N_7615,N_6502,N_6541);
nand U7616 (N_7616,N_6102,N_6831);
xnor U7617 (N_7617,N_6528,N_6568);
nand U7618 (N_7618,N_6089,N_6002);
xor U7619 (N_7619,N_6662,N_6272);
nor U7620 (N_7620,N_6509,N_6665);
nand U7621 (N_7621,N_6314,N_6004);
and U7622 (N_7622,N_6611,N_6367);
nand U7623 (N_7623,N_6236,N_6787);
or U7624 (N_7624,N_6450,N_6273);
nor U7625 (N_7625,N_6374,N_6126);
nand U7626 (N_7626,N_6514,N_6561);
nand U7627 (N_7627,N_6502,N_6107);
xor U7628 (N_7628,N_6125,N_6454);
nand U7629 (N_7629,N_6362,N_6539);
or U7630 (N_7630,N_6302,N_6397);
nand U7631 (N_7631,N_6669,N_6822);
xor U7632 (N_7632,N_6372,N_6470);
nor U7633 (N_7633,N_6375,N_6709);
or U7634 (N_7634,N_6948,N_6682);
xnor U7635 (N_7635,N_6931,N_6027);
and U7636 (N_7636,N_6937,N_6943);
and U7637 (N_7637,N_6810,N_6892);
and U7638 (N_7638,N_6806,N_6662);
or U7639 (N_7639,N_6151,N_6777);
or U7640 (N_7640,N_6036,N_6009);
nor U7641 (N_7641,N_6062,N_6717);
and U7642 (N_7642,N_6424,N_6498);
xor U7643 (N_7643,N_6068,N_6813);
nand U7644 (N_7644,N_6369,N_6434);
nand U7645 (N_7645,N_6975,N_6118);
or U7646 (N_7646,N_6187,N_6999);
nor U7647 (N_7647,N_6645,N_6456);
nand U7648 (N_7648,N_6613,N_6870);
nor U7649 (N_7649,N_6572,N_6767);
and U7650 (N_7650,N_6871,N_6708);
xor U7651 (N_7651,N_6188,N_6060);
and U7652 (N_7652,N_6777,N_6358);
nor U7653 (N_7653,N_6780,N_6895);
nor U7654 (N_7654,N_6504,N_6932);
and U7655 (N_7655,N_6045,N_6384);
or U7656 (N_7656,N_6140,N_6405);
and U7657 (N_7657,N_6160,N_6265);
nor U7658 (N_7658,N_6892,N_6439);
and U7659 (N_7659,N_6228,N_6896);
and U7660 (N_7660,N_6640,N_6917);
xor U7661 (N_7661,N_6497,N_6567);
nor U7662 (N_7662,N_6929,N_6321);
or U7663 (N_7663,N_6610,N_6525);
xor U7664 (N_7664,N_6300,N_6842);
or U7665 (N_7665,N_6437,N_6070);
xor U7666 (N_7666,N_6132,N_6778);
or U7667 (N_7667,N_6060,N_6178);
nand U7668 (N_7668,N_6849,N_6470);
or U7669 (N_7669,N_6257,N_6227);
xnor U7670 (N_7670,N_6201,N_6106);
xnor U7671 (N_7671,N_6849,N_6170);
and U7672 (N_7672,N_6843,N_6669);
xor U7673 (N_7673,N_6908,N_6747);
nor U7674 (N_7674,N_6196,N_6709);
or U7675 (N_7675,N_6370,N_6548);
nor U7676 (N_7676,N_6129,N_6160);
nor U7677 (N_7677,N_6439,N_6584);
xnor U7678 (N_7678,N_6648,N_6514);
xnor U7679 (N_7679,N_6359,N_6371);
nor U7680 (N_7680,N_6003,N_6949);
xnor U7681 (N_7681,N_6872,N_6392);
nand U7682 (N_7682,N_6152,N_6560);
nor U7683 (N_7683,N_6263,N_6578);
and U7684 (N_7684,N_6602,N_6983);
nor U7685 (N_7685,N_6259,N_6902);
nand U7686 (N_7686,N_6837,N_6708);
nor U7687 (N_7687,N_6174,N_6508);
and U7688 (N_7688,N_6469,N_6672);
nor U7689 (N_7689,N_6788,N_6895);
or U7690 (N_7690,N_6507,N_6455);
xor U7691 (N_7691,N_6362,N_6356);
xnor U7692 (N_7692,N_6151,N_6033);
or U7693 (N_7693,N_6553,N_6416);
and U7694 (N_7694,N_6250,N_6647);
or U7695 (N_7695,N_6243,N_6699);
nor U7696 (N_7696,N_6561,N_6501);
nand U7697 (N_7697,N_6463,N_6386);
nor U7698 (N_7698,N_6120,N_6378);
nor U7699 (N_7699,N_6796,N_6958);
nor U7700 (N_7700,N_6369,N_6335);
and U7701 (N_7701,N_6309,N_6960);
or U7702 (N_7702,N_6722,N_6210);
and U7703 (N_7703,N_6918,N_6891);
or U7704 (N_7704,N_6826,N_6954);
and U7705 (N_7705,N_6563,N_6821);
nor U7706 (N_7706,N_6515,N_6610);
nor U7707 (N_7707,N_6974,N_6544);
and U7708 (N_7708,N_6363,N_6079);
and U7709 (N_7709,N_6504,N_6299);
xor U7710 (N_7710,N_6598,N_6482);
and U7711 (N_7711,N_6077,N_6432);
or U7712 (N_7712,N_6683,N_6604);
or U7713 (N_7713,N_6604,N_6927);
and U7714 (N_7714,N_6919,N_6632);
or U7715 (N_7715,N_6098,N_6131);
and U7716 (N_7716,N_6587,N_6557);
xor U7717 (N_7717,N_6038,N_6615);
nand U7718 (N_7718,N_6867,N_6261);
nand U7719 (N_7719,N_6216,N_6267);
nand U7720 (N_7720,N_6858,N_6690);
nor U7721 (N_7721,N_6175,N_6785);
and U7722 (N_7722,N_6070,N_6036);
nor U7723 (N_7723,N_6036,N_6948);
xnor U7724 (N_7724,N_6903,N_6245);
or U7725 (N_7725,N_6695,N_6150);
nand U7726 (N_7726,N_6426,N_6130);
nand U7727 (N_7727,N_6084,N_6452);
and U7728 (N_7728,N_6979,N_6012);
or U7729 (N_7729,N_6951,N_6647);
or U7730 (N_7730,N_6238,N_6428);
nand U7731 (N_7731,N_6719,N_6471);
nor U7732 (N_7732,N_6289,N_6012);
nor U7733 (N_7733,N_6174,N_6726);
nor U7734 (N_7734,N_6172,N_6081);
nor U7735 (N_7735,N_6872,N_6602);
and U7736 (N_7736,N_6324,N_6181);
and U7737 (N_7737,N_6340,N_6191);
nor U7738 (N_7738,N_6163,N_6695);
and U7739 (N_7739,N_6319,N_6914);
nor U7740 (N_7740,N_6634,N_6955);
nand U7741 (N_7741,N_6261,N_6107);
xor U7742 (N_7742,N_6339,N_6251);
or U7743 (N_7743,N_6229,N_6671);
nor U7744 (N_7744,N_6624,N_6405);
xor U7745 (N_7745,N_6269,N_6425);
nor U7746 (N_7746,N_6900,N_6981);
nand U7747 (N_7747,N_6558,N_6351);
or U7748 (N_7748,N_6040,N_6947);
nor U7749 (N_7749,N_6602,N_6165);
nand U7750 (N_7750,N_6373,N_6608);
or U7751 (N_7751,N_6588,N_6731);
nand U7752 (N_7752,N_6347,N_6955);
and U7753 (N_7753,N_6244,N_6678);
nand U7754 (N_7754,N_6301,N_6805);
or U7755 (N_7755,N_6450,N_6867);
and U7756 (N_7756,N_6659,N_6771);
and U7757 (N_7757,N_6447,N_6778);
or U7758 (N_7758,N_6166,N_6921);
and U7759 (N_7759,N_6962,N_6321);
nor U7760 (N_7760,N_6849,N_6290);
and U7761 (N_7761,N_6781,N_6452);
xnor U7762 (N_7762,N_6135,N_6899);
or U7763 (N_7763,N_6157,N_6748);
and U7764 (N_7764,N_6366,N_6171);
and U7765 (N_7765,N_6588,N_6150);
or U7766 (N_7766,N_6409,N_6447);
xnor U7767 (N_7767,N_6725,N_6137);
nand U7768 (N_7768,N_6132,N_6829);
or U7769 (N_7769,N_6105,N_6642);
xnor U7770 (N_7770,N_6520,N_6933);
or U7771 (N_7771,N_6476,N_6483);
nand U7772 (N_7772,N_6808,N_6809);
nand U7773 (N_7773,N_6773,N_6531);
nand U7774 (N_7774,N_6715,N_6248);
xor U7775 (N_7775,N_6525,N_6770);
nor U7776 (N_7776,N_6559,N_6600);
or U7777 (N_7777,N_6504,N_6500);
or U7778 (N_7778,N_6812,N_6401);
or U7779 (N_7779,N_6736,N_6642);
nor U7780 (N_7780,N_6260,N_6369);
xor U7781 (N_7781,N_6125,N_6659);
xor U7782 (N_7782,N_6939,N_6062);
nor U7783 (N_7783,N_6320,N_6465);
and U7784 (N_7784,N_6709,N_6110);
and U7785 (N_7785,N_6541,N_6703);
xnor U7786 (N_7786,N_6139,N_6112);
or U7787 (N_7787,N_6382,N_6790);
xnor U7788 (N_7788,N_6371,N_6367);
nor U7789 (N_7789,N_6783,N_6104);
nor U7790 (N_7790,N_6554,N_6853);
nand U7791 (N_7791,N_6209,N_6081);
and U7792 (N_7792,N_6519,N_6750);
nor U7793 (N_7793,N_6336,N_6821);
nand U7794 (N_7794,N_6676,N_6949);
xor U7795 (N_7795,N_6087,N_6648);
nand U7796 (N_7796,N_6330,N_6388);
xnor U7797 (N_7797,N_6673,N_6172);
nand U7798 (N_7798,N_6459,N_6598);
nand U7799 (N_7799,N_6010,N_6497);
nor U7800 (N_7800,N_6930,N_6153);
and U7801 (N_7801,N_6755,N_6025);
xor U7802 (N_7802,N_6419,N_6876);
xor U7803 (N_7803,N_6400,N_6593);
nor U7804 (N_7804,N_6732,N_6193);
and U7805 (N_7805,N_6575,N_6445);
and U7806 (N_7806,N_6383,N_6232);
and U7807 (N_7807,N_6001,N_6422);
and U7808 (N_7808,N_6794,N_6273);
xor U7809 (N_7809,N_6906,N_6917);
and U7810 (N_7810,N_6771,N_6238);
nand U7811 (N_7811,N_6304,N_6347);
or U7812 (N_7812,N_6172,N_6287);
nand U7813 (N_7813,N_6754,N_6539);
and U7814 (N_7814,N_6679,N_6116);
nand U7815 (N_7815,N_6588,N_6925);
xor U7816 (N_7816,N_6707,N_6144);
or U7817 (N_7817,N_6746,N_6877);
and U7818 (N_7818,N_6426,N_6910);
nor U7819 (N_7819,N_6998,N_6952);
or U7820 (N_7820,N_6372,N_6833);
nand U7821 (N_7821,N_6279,N_6204);
nor U7822 (N_7822,N_6994,N_6746);
nor U7823 (N_7823,N_6980,N_6539);
or U7824 (N_7824,N_6919,N_6718);
nand U7825 (N_7825,N_6619,N_6328);
or U7826 (N_7826,N_6453,N_6634);
xnor U7827 (N_7827,N_6136,N_6471);
nor U7828 (N_7828,N_6236,N_6412);
nor U7829 (N_7829,N_6506,N_6966);
nand U7830 (N_7830,N_6066,N_6846);
and U7831 (N_7831,N_6314,N_6301);
nand U7832 (N_7832,N_6041,N_6412);
xnor U7833 (N_7833,N_6760,N_6987);
and U7834 (N_7834,N_6534,N_6323);
nor U7835 (N_7835,N_6080,N_6506);
xnor U7836 (N_7836,N_6001,N_6986);
and U7837 (N_7837,N_6144,N_6186);
and U7838 (N_7838,N_6225,N_6812);
nor U7839 (N_7839,N_6358,N_6926);
nand U7840 (N_7840,N_6058,N_6703);
and U7841 (N_7841,N_6793,N_6107);
and U7842 (N_7842,N_6676,N_6339);
xnor U7843 (N_7843,N_6480,N_6189);
and U7844 (N_7844,N_6605,N_6162);
nand U7845 (N_7845,N_6332,N_6520);
xnor U7846 (N_7846,N_6436,N_6541);
nand U7847 (N_7847,N_6914,N_6175);
xor U7848 (N_7848,N_6378,N_6019);
and U7849 (N_7849,N_6550,N_6853);
and U7850 (N_7850,N_6061,N_6430);
or U7851 (N_7851,N_6184,N_6552);
xnor U7852 (N_7852,N_6228,N_6346);
or U7853 (N_7853,N_6210,N_6228);
xnor U7854 (N_7854,N_6417,N_6540);
or U7855 (N_7855,N_6383,N_6560);
nor U7856 (N_7856,N_6346,N_6977);
nand U7857 (N_7857,N_6751,N_6947);
or U7858 (N_7858,N_6225,N_6933);
and U7859 (N_7859,N_6022,N_6143);
nor U7860 (N_7860,N_6037,N_6788);
and U7861 (N_7861,N_6600,N_6459);
or U7862 (N_7862,N_6276,N_6434);
xor U7863 (N_7863,N_6601,N_6322);
nand U7864 (N_7864,N_6896,N_6929);
xnor U7865 (N_7865,N_6570,N_6775);
nand U7866 (N_7866,N_6177,N_6867);
xor U7867 (N_7867,N_6444,N_6147);
nor U7868 (N_7868,N_6097,N_6201);
or U7869 (N_7869,N_6347,N_6128);
nand U7870 (N_7870,N_6128,N_6719);
nand U7871 (N_7871,N_6434,N_6122);
and U7872 (N_7872,N_6779,N_6393);
or U7873 (N_7873,N_6895,N_6476);
nor U7874 (N_7874,N_6506,N_6925);
nand U7875 (N_7875,N_6916,N_6089);
and U7876 (N_7876,N_6670,N_6323);
and U7877 (N_7877,N_6526,N_6768);
and U7878 (N_7878,N_6090,N_6715);
or U7879 (N_7879,N_6194,N_6228);
or U7880 (N_7880,N_6961,N_6519);
xor U7881 (N_7881,N_6666,N_6157);
xnor U7882 (N_7882,N_6694,N_6270);
and U7883 (N_7883,N_6293,N_6621);
nand U7884 (N_7884,N_6148,N_6249);
or U7885 (N_7885,N_6715,N_6992);
or U7886 (N_7886,N_6296,N_6380);
nand U7887 (N_7887,N_6202,N_6030);
xnor U7888 (N_7888,N_6163,N_6751);
nor U7889 (N_7889,N_6287,N_6788);
and U7890 (N_7890,N_6168,N_6609);
or U7891 (N_7891,N_6311,N_6889);
or U7892 (N_7892,N_6240,N_6820);
nor U7893 (N_7893,N_6777,N_6769);
xnor U7894 (N_7894,N_6340,N_6841);
nand U7895 (N_7895,N_6916,N_6717);
nand U7896 (N_7896,N_6186,N_6784);
and U7897 (N_7897,N_6685,N_6744);
nor U7898 (N_7898,N_6396,N_6188);
xnor U7899 (N_7899,N_6811,N_6177);
nand U7900 (N_7900,N_6437,N_6604);
nand U7901 (N_7901,N_6868,N_6675);
nor U7902 (N_7902,N_6436,N_6343);
and U7903 (N_7903,N_6572,N_6916);
nor U7904 (N_7904,N_6084,N_6573);
nand U7905 (N_7905,N_6786,N_6628);
and U7906 (N_7906,N_6341,N_6630);
xnor U7907 (N_7907,N_6600,N_6553);
nand U7908 (N_7908,N_6106,N_6323);
xor U7909 (N_7909,N_6251,N_6661);
xnor U7910 (N_7910,N_6400,N_6781);
nor U7911 (N_7911,N_6092,N_6941);
nor U7912 (N_7912,N_6609,N_6494);
nand U7913 (N_7913,N_6654,N_6253);
or U7914 (N_7914,N_6786,N_6486);
and U7915 (N_7915,N_6815,N_6273);
and U7916 (N_7916,N_6225,N_6451);
nor U7917 (N_7917,N_6168,N_6542);
or U7918 (N_7918,N_6053,N_6084);
and U7919 (N_7919,N_6300,N_6461);
xor U7920 (N_7920,N_6587,N_6464);
nor U7921 (N_7921,N_6614,N_6143);
and U7922 (N_7922,N_6734,N_6343);
or U7923 (N_7923,N_6382,N_6015);
xor U7924 (N_7924,N_6529,N_6940);
nor U7925 (N_7925,N_6964,N_6324);
xor U7926 (N_7926,N_6876,N_6453);
xor U7927 (N_7927,N_6582,N_6883);
or U7928 (N_7928,N_6637,N_6964);
and U7929 (N_7929,N_6468,N_6887);
nor U7930 (N_7930,N_6394,N_6786);
xor U7931 (N_7931,N_6019,N_6479);
nor U7932 (N_7932,N_6641,N_6288);
nand U7933 (N_7933,N_6880,N_6576);
nor U7934 (N_7934,N_6428,N_6310);
and U7935 (N_7935,N_6323,N_6205);
nor U7936 (N_7936,N_6378,N_6490);
and U7937 (N_7937,N_6066,N_6916);
xor U7938 (N_7938,N_6698,N_6382);
nand U7939 (N_7939,N_6289,N_6467);
nand U7940 (N_7940,N_6200,N_6005);
or U7941 (N_7941,N_6644,N_6380);
or U7942 (N_7942,N_6068,N_6486);
nand U7943 (N_7943,N_6998,N_6861);
or U7944 (N_7944,N_6418,N_6142);
nor U7945 (N_7945,N_6707,N_6657);
or U7946 (N_7946,N_6718,N_6736);
xnor U7947 (N_7947,N_6151,N_6042);
and U7948 (N_7948,N_6195,N_6305);
xor U7949 (N_7949,N_6980,N_6881);
or U7950 (N_7950,N_6498,N_6205);
xnor U7951 (N_7951,N_6422,N_6427);
nor U7952 (N_7952,N_6105,N_6949);
nand U7953 (N_7953,N_6419,N_6781);
or U7954 (N_7954,N_6597,N_6914);
or U7955 (N_7955,N_6785,N_6223);
or U7956 (N_7956,N_6431,N_6153);
or U7957 (N_7957,N_6431,N_6267);
or U7958 (N_7958,N_6628,N_6568);
or U7959 (N_7959,N_6904,N_6357);
and U7960 (N_7960,N_6124,N_6074);
or U7961 (N_7961,N_6130,N_6647);
or U7962 (N_7962,N_6952,N_6724);
nand U7963 (N_7963,N_6941,N_6841);
nand U7964 (N_7964,N_6318,N_6608);
xnor U7965 (N_7965,N_6399,N_6377);
xor U7966 (N_7966,N_6114,N_6928);
or U7967 (N_7967,N_6708,N_6544);
nor U7968 (N_7968,N_6076,N_6911);
and U7969 (N_7969,N_6025,N_6501);
nand U7970 (N_7970,N_6497,N_6593);
or U7971 (N_7971,N_6442,N_6619);
xor U7972 (N_7972,N_6049,N_6289);
xor U7973 (N_7973,N_6160,N_6493);
nand U7974 (N_7974,N_6220,N_6968);
and U7975 (N_7975,N_6874,N_6153);
nand U7976 (N_7976,N_6838,N_6892);
xnor U7977 (N_7977,N_6052,N_6476);
or U7978 (N_7978,N_6523,N_6688);
and U7979 (N_7979,N_6465,N_6199);
or U7980 (N_7980,N_6933,N_6493);
nand U7981 (N_7981,N_6184,N_6269);
and U7982 (N_7982,N_6038,N_6178);
nand U7983 (N_7983,N_6620,N_6310);
and U7984 (N_7984,N_6925,N_6240);
or U7985 (N_7985,N_6186,N_6229);
and U7986 (N_7986,N_6026,N_6134);
or U7987 (N_7987,N_6104,N_6860);
and U7988 (N_7988,N_6508,N_6293);
and U7989 (N_7989,N_6399,N_6194);
nor U7990 (N_7990,N_6096,N_6032);
nand U7991 (N_7991,N_6354,N_6797);
or U7992 (N_7992,N_6455,N_6067);
and U7993 (N_7993,N_6688,N_6159);
nand U7994 (N_7994,N_6110,N_6114);
nor U7995 (N_7995,N_6186,N_6121);
and U7996 (N_7996,N_6684,N_6079);
nand U7997 (N_7997,N_6643,N_6621);
and U7998 (N_7998,N_6341,N_6698);
and U7999 (N_7999,N_6982,N_6674);
nand U8000 (N_8000,N_7178,N_7074);
nor U8001 (N_8001,N_7329,N_7986);
nor U8002 (N_8002,N_7768,N_7731);
and U8003 (N_8003,N_7000,N_7494);
nand U8004 (N_8004,N_7645,N_7489);
or U8005 (N_8005,N_7369,N_7851);
nand U8006 (N_8006,N_7051,N_7314);
or U8007 (N_8007,N_7692,N_7355);
or U8008 (N_8008,N_7901,N_7853);
and U8009 (N_8009,N_7292,N_7516);
and U8010 (N_8010,N_7120,N_7041);
nand U8011 (N_8011,N_7023,N_7611);
nor U8012 (N_8012,N_7955,N_7211);
or U8013 (N_8013,N_7983,N_7043);
or U8014 (N_8014,N_7716,N_7264);
xnor U8015 (N_8015,N_7950,N_7831);
or U8016 (N_8016,N_7787,N_7810);
and U8017 (N_8017,N_7534,N_7490);
and U8018 (N_8018,N_7213,N_7911);
nand U8019 (N_8019,N_7166,N_7561);
nand U8020 (N_8020,N_7421,N_7048);
nand U8021 (N_8021,N_7339,N_7402);
xor U8022 (N_8022,N_7256,N_7274);
and U8023 (N_8023,N_7224,N_7958);
nand U8024 (N_8024,N_7728,N_7126);
or U8025 (N_8025,N_7954,N_7942);
and U8026 (N_8026,N_7107,N_7061);
xor U8027 (N_8027,N_7594,N_7883);
nand U8028 (N_8028,N_7872,N_7575);
nor U8029 (N_8029,N_7981,N_7888);
nand U8030 (N_8030,N_7485,N_7088);
nor U8031 (N_8031,N_7742,N_7801);
nor U8032 (N_8032,N_7448,N_7539);
xnor U8033 (N_8033,N_7610,N_7674);
xor U8034 (N_8034,N_7308,N_7142);
or U8035 (N_8035,N_7371,N_7102);
or U8036 (N_8036,N_7811,N_7838);
and U8037 (N_8037,N_7229,N_7583);
nor U8038 (N_8038,N_7342,N_7745);
xor U8039 (N_8039,N_7476,N_7457);
and U8040 (N_8040,N_7676,N_7190);
and U8041 (N_8041,N_7533,N_7303);
or U8042 (N_8042,N_7999,N_7245);
nor U8043 (N_8043,N_7825,N_7668);
or U8044 (N_8044,N_7125,N_7070);
nand U8045 (N_8045,N_7030,N_7722);
nor U8046 (N_8046,N_7311,N_7289);
nor U8047 (N_8047,N_7186,N_7093);
xnor U8048 (N_8048,N_7739,N_7297);
nand U8049 (N_8049,N_7702,N_7206);
nor U8050 (N_8050,N_7449,N_7138);
nand U8051 (N_8051,N_7390,N_7580);
or U8052 (N_8052,N_7977,N_7744);
and U8053 (N_8053,N_7760,N_7481);
or U8054 (N_8054,N_7252,N_7881);
nor U8055 (N_8055,N_7595,N_7972);
nor U8056 (N_8056,N_7115,N_7053);
and U8057 (N_8057,N_7149,N_7623);
nor U8058 (N_8058,N_7727,N_7600);
xnor U8059 (N_8059,N_7841,N_7748);
nand U8060 (N_8060,N_7531,N_7444);
nor U8061 (N_8061,N_7208,N_7873);
or U8062 (N_8062,N_7033,N_7124);
and U8063 (N_8063,N_7541,N_7191);
and U8064 (N_8064,N_7935,N_7067);
nand U8065 (N_8065,N_7202,N_7649);
or U8066 (N_8066,N_7767,N_7546);
nor U8067 (N_8067,N_7587,N_7525);
nand U8068 (N_8068,N_7424,N_7164);
and U8069 (N_8069,N_7968,N_7522);
or U8070 (N_8070,N_7473,N_7464);
xnor U8071 (N_8071,N_7903,N_7562);
and U8072 (N_8072,N_7528,N_7771);
nor U8073 (N_8073,N_7431,N_7076);
nor U8074 (N_8074,N_7374,N_7151);
xor U8075 (N_8075,N_7397,N_7871);
nor U8076 (N_8076,N_7082,N_7622);
nor U8077 (N_8077,N_7073,N_7215);
nor U8078 (N_8078,N_7543,N_7705);
nor U8079 (N_8079,N_7936,N_7244);
nand U8080 (N_8080,N_7313,N_7391);
or U8081 (N_8081,N_7930,N_7203);
xnor U8082 (N_8082,N_7373,N_7785);
nor U8083 (N_8083,N_7350,N_7666);
nor U8084 (N_8084,N_7634,N_7775);
or U8085 (N_8085,N_7773,N_7929);
nor U8086 (N_8086,N_7772,N_7301);
and U8087 (N_8087,N_7175,N_7226);
nand U8088 (N_8088,N_7018,N_7985);
or U8089 (N_8089,N_7196,N_7386);
and U8090 (N_8090,N_7209,N_7241);
nand U8091 (N_8091,N_7432,N_7309);
xor U8092 (N_8092,N_7167,N_7640);
nand U8093 (N_8093,N_7323,N_7334);
and U8094 (N_8094,N_7145,N_7212);
or U8095 (N_8095,N_7087,N_7777);
or U8096 (N_8096,N_7536,N_7804);
and U8097 (N_8097,N_7332,N_7358);
nand U8098 (N_8098,N_7139,N_7479);
xor U8099 (N_8099,N_7290,N_7752);
nand U8100 (N_8100,N_7195,N_7007);
nor U8101 (N_8101,N_7800,N_7267);
nand U8102 (N_8102,N_7571,N_7606);
nor U8103 (N_8103,N_7116,N_7460);
nand U8104 (N_8104,N_7419,N_7450);
or U8105 (N_8105,N_7480,N_7909);
nand U8106 (N_8106,N_7112,N_7598);
nor U8107 (N_8107,N_7524,N_7343);
or U8108 (N_8108,N_7009,N_7060);
or U8109 (N_8109,N_7592,N_7319);
nor U8110 (N_8110,N_7564,N_7637);
xnor U8111 (N_8111,N_7596,N_7751);
nand U8112 (N_8112,N_7140,N_7057);
nand U8113 (N_8113,N_7459,N_7130);
and U8114 (N_8114,N_7483,N_7345);
or U8115 (N_8115,N_7667,N_7101);
xor U8116 (N_8116,N_7133,N_7550);
and U8117 (N_8117,N_7786,N_7656);
nor U8118 (N_8118,N_7755,N_7947);
nand U8119 (N_8119,N_7188,N_7867);
nor U8120 (N_8120,N_7761,N_7613);
nor U8121 (N_8121,N_7884,N_7484);
nor U8122 (N_8122,N_7635,N_7478);
nand U8123 (N_8123,N_7512,N_7337);
nand U8124 (N_8124,N_7989,N_7643);
or U8125 (N_8125,N_7998,N_7732);
nor U8126 (N_8126,N_7495,N_7090);
xor U8127 (N_8127,N_7907,N_7700);
and U8128 (N_8128,N_7671,N_7978);
nand U8129 (N_8129,N_7890,N_7078);
xnor U8130 (N_8130,N_7180,N_7508);
nor U8131 (N_8131,N_7365,N_7664);
nand U8132 (N_8132,N_7326,N_7172);
nand U8133 (N_8133,N_7197,N_7919);
and U8134 (N_8134,N_7975,N_7399);
or U8135 (N_8135,N_7537,N_7520);
xnor U8136 (N_8136,N_7044,N_7654);
and U8137 (N_8137,N_7617,N_7582);
or U8138 (N_8138,N_7778,N_7880);
nor U8139 (N_8139,N_7819,N_7554);
xnor U8140 (N_8140,N_7136,N_7375);
nand U8141 (N_8141,N_7517,N_7360);
nand U8142 (N_8142,N_7774,N_7835);
nand U8143 (N_8143,N_7258,N_7718);
xor U8144 (N_8144,N_7361,N_7653);
xor U8145 (N_8145,N_7518,N_7660);
xor U8146 (N_8146,N_7430,N_7899);
or U8147 (N_8147,N_7754,N_7706);
nor U8148 (N_8148,N_7307,N_7222);
xor U8149 (N_8149,N_7847,N_7812);
nor U8150 (N_8150,N_7410,N_7865);
xor U8151 (N_8151,N_7458,N_7693);
and U8152 (N_8152,N_7927,N_7184);
xnor U8153 (N_8153,N_7058,N_7822);
nor U8154 (N_8154,N_7185,N_7472);
and U8155 (N_8155,N_7004,N_7788);
or U8156 (N_8156,N_7856,N_7670);
and U8157 (N_8157,N_7746,N_7165);
nor U8158 (N_8158,N_7372,N_7217);
or U8159 (N_8159,N_7945,N_7680);
or U8160 (N_8160,N_7148,N_7387);
nand U8161 (N_8161,N_7277,N_7367);
and U8162 (N_8162,N_7182,N_7262);
nor U8163 (N_8163,N_7796,N_7699);
and U8164 (N_8164,N_7563,N_7802);
and U8165 (N_8165,N_7734,N_7569);
or U8166 (N_8166,N_7228,N_7287);
or U8167 (N_8167,N_7500,N_7503);
or U8168 (N_8168,N_7254,N_7153);
nor U8169 (N_8169,N_7455,N_7552);
nand U8170 (N_8170,N_7515,N_7420);
nor U8171 (N_8171,N_7704,N_7336);
or U8172 (N_8172,N_7002,N_7905);
or U8173 (N_8173,N_7962,N_7615);
and U8174 (N_8174,N_7233,N_7527);
nor U8175 (N_8175,N_7282,N_7170);
xor U8176 (N_8176,N_7389,N_7694);
nor U8177 (N_8177,N_7408,N_7789);
and U8178 (N_8178,N_7817,N_7576);
nand U8179 (N_8179,N_7828,N_7176);
nand U8180 (N_8180,N_7870,N_7904);
nor U8181 (N_8181,N_7276,N_7965);
or U8182 (N_8182,N_7852,N_7377);
or U8183 (N_8183,N_7894,N_7510);
and U8184 (N_8184,N_7114,N_7366);
or U8185 (N_8185,N_7357,N_7032);
xnor U8186 (N_8186,N_7862,N_7349);
nor U8187 (N_8187,N_7467,N_7542);
nand U8188 (N_8188,N_7021,N_7493);
nand U8189 (N_8189,N_7348,N_7766);
or U8190 (N_8190,N_7123,N_7246);
nand U8191 (N_8191,N_7638,N_7984);
nand U8192 (N_8192,N_7902,N_7129);
or U8193 (N_8193,N_7687,N_7696);
nand U8194 (N_8194,N_7681,N_7996);
nand U8195 (N_8195,N_7616,N_7095);
xor U8196 (N_8196,N_7679,N_7255);
nor U8197 (N_8197,N_7299,N_7982);
or U8198 (N_8198,N_7143,N_7462);
or U8199 (N_8199,N_7220,N_7069);
nor U8200 (N_8200,N_7589,N_7625);
nand U8201 (N_8201,N_7415,N_7715);
xor U8202 (N_8202,N_7678,N_7118);
and U8203 (N_8203,N_7417,N_7280);
nand U8204 (N_8204,N_7216,N_7869);
nand U8205 (N_8205,N_7944,N_7733);
or U8206 (N_8206,N_7131,N_7497);
xnor U8207 (N_8207,N_7354,N_7317);
or U8208 (N_8208,N_7655,N_7709);
and U8209 (N_8209,N_7232,N_7097);
and U8210 (N_8210,N_7566,N_7347);
and U8211 (N_8211,N_7341,N_7187);
or U8212 (N_8212,N_7845,N_7557);
xnor U8213 (N_8213,N_7868,N_7505);
or U8214 (N_8214,N_7492,N_7221);
xnor U8215 (N_8215,N_7662,N_7293);
and U8216 (N_8216,N_7612,N_7991);
nor U8217 (N_8217,N_7895,N_7141);
nand U8218 (N_8218,N_7193,N_7511);
xnor U8219 (N_8219,N_7315,N_7647);
or U8220 (N_8220,N_7798,N_7234);
or U8221 (N_8221,N_7908,N_7194);
or U8222 (N_8222,N_7814,N_7128);
nand U8223 (N_8223,N_7414,N_7995);
nand U8224 (N_8224,N_7382,N_7750);
nand U8225 (N_8225,N_7049,N_7268);
xor U8226 (N_8226,N_7427,N_7703);
nor U8227 (N_8227,N_7532,N_7443);
and U8228 (N_8228,N_7012,N_7330);
xnor U8229 (N_8229,N_7891,N_7946);
nand U8230 (N_8230,N_7920,N_7017);
xnor U8231 (N_8231,N_7103,N_7558);
and U8232 (N_8232,N_7376,N_7629);
nor U8233 (N_8233,N_7691,N_7335);
nand U8234 (N_8234,N_7820,N_7031);
and U8235 (N_8235,N_7724,N_7833);
or U8236 (N_8236,N_7100,N_7501);
nor U8237 (N_8237,N_7207,N_7957);
nor U8238 (N_8238,N_7034,N_7108);
xnor U8239 (N_8239,N_7482,N_7475);
or U8240 (N_8240,N_7383,N_7723);
nand U8241 (N_8241,N_7837,N_7689);
xor U8242 (N_8242,N_7456,N_7370);
nor U8243 (N_8243,N_7089,N_7604);
nand U8244 (N_8244,N_7295,N_7028);
nand U8245 (N_8245,N_7111,N_7168);
or U8246 (N_8246,N_7618,N_7230);
nor U8247 (N_8247,N_7385,N_7834);
nand U8248 (N_8248,N_7675,N_7849);
or U8249 (N_8249,N_7970,N_7368);
or U8250 (N_8250,N_7897,N_7568);
xnor U8251 (N_8251,N_7974,N_7588);
and U8252 (N_8252,N_7488,N_7266);
or U8253 (N_8253,N_7914,N_7659);
xnor U8254 (N_8254,N_7949,N_7016);
or U8255 (N_8255,N_7218,N_7677);
nor U8256 (N_8256,N_7154,N_7923);
or U8257 (N_8257,N_7439,N_7401);
nand U8258 (N_8258,N_7306,N_7504);
or U8259 (N_8259,N_7393,N_7388);
or U8260 (N_8260,N_7614,N_7793);
and U8261 (N_8261,N_7782,N_7591);
xor U8262 (N_8262,N_7713,N_7286);
nand U8263 (N_8263,N_7379,N_7925);
or U8264 (N_8264,N_7827,N_7001);
xor U8265 (N_8265,N_7105,N_7840);
or U8266 (N_8266,N_7988,N_7338);
xnor U8267 (N_8267,N_7300,N_7658);
xnor U8268 (N_8268,N_7400,N_7413);
or U8269 (N_8269,N_7015,N_7565);
nand U8270 (N_8270,N_7036,N_7815);
or U8271 (N_8271,N_7199,N_7547);
nand U8272 (N_8272,N_7273,N_7506);
and U8273 (N_8273,N_7839,N_7863);
or U8274 (N_8274,N_7725,N_7816);
or U8275 (N_8275,N_7113,N_7310);
and U8276 (N_8276,N_7214,N_7045);
and U8277 (N_8277,N_7405,N_7607);
or U8278 (N_8278,N_7780,N_7875);
nand U8279 (N_8279,N_7066,N_7454);
or U8280 (N_8280,N_7447,N_7913);
or U8281 (N_8281,N_7010,N_7316);
nand U8282 (N_8282,N_7451,N_7227);
xor U8283 (N_8283,N_7509,N_7257);
or U8284 (N_8284,N_7271,N_7650);
xnor U8285 (N_8285,N_7085,N_7398);
nand U8286 (N_8286,N_7758,N_7673);
nor U8287 (N_8287,N_7624,N_7210);
and U8288 (N_8288,N_7896,N_7885);
or U8289 (N_8289,N_7738,N_7412);
nand U8290 (N_8290,N_7824,N_7491);
or U8291 (N_8291,N_7701,N_7325);
nand U8292 (N_8292,N_7452,N_7160);
and U8293 (N_8293,N_7247,N_7351);
nand U8294 (N_8294,N_7513,N_7364);
xor U8295 (N_8295,N_7380,N_7630);
nor U8296 (N_8296,N_7684,N_7079);
nand U8297 (N_8297,N_7205,N_7094);
nand U8298 (N_8298,N_7265,N_7423);
nand U8299 (N_8299,N_7327,N_7008);
and U8300 (N_8300,N_7850,N_7104);
or U8301 (N_8301,N_7577,N_7081);
or U8302 (N_8302,N_7642,N_7665);
xor U8303 (N_8303,N_7147,N_7469);
or U8304 (N_8304,N_7855,N_7470);
or U8305 (N_8305,N_7446,N_7039);
and U8306 (N_8306,N_7466,N_7052);
nor U8307 (N_8307,N_7019,N_7243);
nor U8308 (N_8308,N_7900,N_7599);
nor U8309 (N_8309,N_7685,N_7519);
nand U8310 (N_8310,N_7741,N_7163);
xor U8311 (N_8311,N_7238,N_7602);
or U8312 (N_8312,N_7915,N_7333);
nand U8313 (N_8313,N_7712,N_7340);
nand U8314 (N_8314,N_7931,N_7381);
and U8315 (N_8315,N_7156,N_7940);
xor U8316 (N_8316,N_7359,N_7169);
xor U8317 (N_8317,N_7086,N_7056);
nor U8318 (N_8318,N_7059,N_7632);
or U8319 (N_8319,N_7248,N_7378);
and U8320 (N_8320,N_7729,N_7445);
nor U8321 (N_8321,N_7441,N_7997);
and U8322 (N_8322,N_7652,N_7106);
xnor U8323 (N_8323,N_7235,N_7499);
or U8324 (N_8324,N_7545,N_7320);
nor U8325 (N_8325,N_7912,N_7553);
nor U8326 (N_8326,N_7826,N_7803);
and U8327 (N_8327,N_7468,N_7434);
and U8328 (N_8328,N_7943,N_7084);
xor U8329 (N_8329,N_7979,N_7759);
and U8330 (N_8330,N_7514,N_7821);
nand U8331 (N_8331,N_7783,N_7259);
nor U8332 (N_8332,N_7404,N_7861);
nand U8333 (N_8333,N_7726,N_7055);
nor U8334 (N_8334,N_7324,N_7077);
nor U8335 (N_8335,N_7302,N_7223);
or U8336 (N_8336,N_7174,N_7127);
and U8337 (N_8337,N_7876,N_7487);
nand U8338 (N_8338,N_7137,N_7710);
or U8339 (N_8339,N_7765,N_7934);
or U8340 (N_8340,N_7620,N_7179);
and U8341 (N_8341,N_7029,N_7590);
and U8342 (N_8342,N_7157,N_7964);
nor U8343 (N_8343,N_7062,N_7425);
and U8344 (N_8344,N_7922,N_7621);
nor U8345 (N_8345,N_7859,N_7858);
xor U8346 (N_8346,N_7406,N_7690);
and U8347 (N_8347,N_7047,N_7240);
and U8348 (N_8348,N_7608,N_7321);
xor U8349 (N_8349,N_7830,N_7892);
xor U8350 (N_8350,N_7776,N_7038);
xnor U8351 (N_8351,N_7416,N_7893);
or U8352 (N_8352,N_7721,N_7886);
nor U8353 (N_8353,N_7159,N_7743);
and U8354 (N_8354,N_7697,N_7763);
or U8355 (N_8355,N_7250,N_7969);
or U8356 (N_8356,N_7628,N_7540);
nor U8357 (N_8357,N_7961,N_7392);
or U8358 (N_8358,N_7987,N_7075);
and U8359 (N_8359,N_7025,N_7874);
or U8360 (N_8360,N_7132,N_7809);
and U8361 (N_8361,N_7993,N_7795);
nand U8362 (N_8362,N_7328,N_7204);
nand U8363 (N_8363,N_7570,N_7918);
nand U8364 (N_8364,N_7020,N_7657);
nand U8365 (N_8365,N_7296,N_7707);
and U8366 (N_8366,N_7578,N_7249);
and U8367 (N_8367,N_7072,N_7435);
nor U8368 (N_8368,N_7411,N_7219);
or U8369 (N_8369,N_7779,N_7555);
and U8370 (N_8370,N_7011,N_7263);
and U8371 (N_8371,N_7854,N_7152);
and U8372 (N_8372,N_7150,N_7080);
nor U8373 (N_8373,N_7573,N_7770);
nand U8374 (N_8374,N_7939,N_7792);
and U8375 (N_8375,N_7040,N_7322);
nand U8376 (N_8376,N_7474,N_7967);
xnor U8377 (N_8377,N_7737,N_7158);
nand U8378 (N_8378,N_7627,N_7708);
nand U8379 (N_8379,N_7046,N_7198);
nor U8380 (N_8380,N_7926,N_7281);
or U8381 (N_8381,N_7714,N_7272);
xnor U8382 (N_8382,N_7717,N_7122);
or U8383 (N_8383,N_7395,N_7110);
or U8384 (N_8384,N_7906,N_7636);
and U8385 (N_8385,N_7619,N_7994);
or U8386 (N_8386,N_7609,N_7284);
nor U8387 (N_8387,N_7866,N_7951);
nand U8388 (N_8388,N_7719,N_7022);
nand U8389 (N_8389,N_7161,N_7574);
nand U8390 (N_8390,N_7192,N_7442);
xor U8391 (N_8391,N_7720,N_7740);
nor U8392 (N_8392,N_7686,N_7261);
and U8393 (N_8393,N_7882,N_7980);
nor U8394 (N_8394,N_7769,N_7237);
or U8395 (N_8395,N_7529,N_7544);
or U8396 (N_8396,N_7035,N_7065);
nor U8397 (N_8397,N_7924,N_7878);
xnor U8398 (N_8398,N_7278,N_7312);
xnor U8399 (N_8399,N_7683,N_7933);
xor U8400 (N_8400,N_7027,N_7848);
or U8401 (N_8401,N_7806,N_7523);
xnor U8402 (N_8402,N_7502,N_7409);
and U8403 (N_8403,N_7037,N_7937);
xor U8404 (N_8404,N_7631,N_7530);
nor U8405 (N_8405,N_7135,N_7231);
xnor U8406 (N_8406,N_7889,N_7932);
xor U8407 (N_8407,N_7966,N_7938);
nand U8408 (N_8408,N_7356,N_7403);
nand U8409 (N_8409,N_7433,N_7794);
nor U8410 (N_8410,N_7661,N_7155);
nor U8411 (N_8411,N_7736,N_7548);
xor U8412 (N_8412,N_7465,N_7601);
or U8413 (N_8413,N_7836,N_7764);
or U8414 (N_8414,N_7916,N_7050);
and U8415 (N_8415,N_7024,N_7960);
nand U8416 (N_8416,N_7730,N_7711);
xor U8417 (N_8417,N_7560,N_7298);
nand U8418 (N_8418,N_7496,N_7183);
or U8419 (N_8419,N_7857,N_7797);
nor U8420 (N_8420,N_7887,N_7807);
xnor U8421 (N_8421,N_7042,N_7663);
xor U8422 (N_8422,N_7879,N_7526);
xor U8423 (N_8423,N_7846,N_7626);
xor U8424 (N_8424,N_7071,N_7651);
or U8425 (N_8425,N_7288,N_7790);
xor U8426 (N_8426,N_7362,N_7842);
or U8427 (N_8427,N_7091,N_7832);
and U8428 (N_8428,N_7805,N_7099);
nor U8429 (N_8429,N_7672,N_7275);
or U8430 (N_8430,N_7921,N_7682);
and U8431 (N_8431,N_7898,N_7603);
and U8432 (N_8432,N_7521,N_7236);
or U8433 (N_8433,N_7173,N_7633);
and U8434 (N_8434,N_7593,N_7781);
and U8435 (N_8435,N_7538,N_7860);
nor U8436 (N_8436,N_7762,N_7584);
and U8437 (N_8437,N_7461,N_7644);
nor U8438 (N_8438,N_7285,N_7953);
nand U8439 (N_8439,N_7352,N_7799);
xor U8440 (N_8440,N_7270,N_7003);
xor U8441 (N_8441,N_7877,N_7990);
nor U8442 (N_8442,N_7429,N_7064);
or U8443 (N_8443,N_7251,N_7477);
nand U8444 (N_8444,N_7586,N_7585);
xor U8445 (N_8445,N_7756,N_7269);
or U8446 (N_8446,N_7083,N_7201);
or U8447 (N_8447,N_7426,N_7639);
nand U8448 (N_8448,N_7535,N_7109);
nand U8449 (N_8449,N_7121,N_7641);
nand U8450 (N_8450,N_7418,N_7407);
xor U8451 (N_8451,N_7428,N_7463);
nor U8452 (N_8452,N_7959,N_7928);
xnor U8453 (N_8453,N_7422,N_7784);
xnor U8454 (N_8454,N_7551,N_7013);
or U8455 (N_8455,N_7146,N_7648);
xor U8456 (N_8456,N_7735,N_7749);
nand U8457 (N_8457,N_7498,N_7976);
and U8458 (N_8458,N_7177,N_7941);
xnor U8459 (N_8459,N_7823,N_7963);
nand U8460 (N_8460,N_7579,N_7006);
nand U8461 (N_8461,N_7572,N_7363);
nand U8462 (N_8462,N_7068,N_7092);
nor U8463 (N_8463,N_7956,N_7384);
and U8464 (N_8464,N_7556,N_7242);
nor U8465 (N_8465,N_7688,N_7394);
nand U8466 (N_8466,N_7181,N_7063);
nor U8467 (N_8467,N_7549,N_7597);
nand U8468 (N_8468,N_7864,N_7098);
nand U8469 (N_8469,N_7014,N_7605);
and U8470 (N_8470,N_7119,N_7283);
or U8471 (N_8471,N_7992,N_7471);
xnor U8472 (N_8472,N_7486,N_7507);
nand U8473 (N_8473,N_7695,N_7973);
nor U8474 (N_8474,N_7189,N_7026);
or U8475 (N_8475,N_7757,N_7747);
nand U8476 (N_8476,N_7829,N_7917);
or U8477 (N_8477,N_7910,N_7344);
xor U8478 (N_8478,N_7952,N_7440);
nand U8479 (N_8479,N_7559,N_7753);
and U8480 (N_8480,N_7005,N_7117);
nand U8481 (N_8481,N_7200,N_7162);
xor U8482 (N_8482,N_7436,N_7813);
nor U8483 (N_8483,N_7669,N_7396);
and U8484 (N_8484,N_7144,N_7134);
and U8485 (N_8485,N_7305,N_7225);
and U8486 (N_8486,N_7291,N_7437);
xnor U8487 (N_8487,N_7331,N_7279);
xnor U8488 (N_8488,N_7567,N_7294);
xor U8489 (N_8489,N_7438,N_7453);
xnor U8490 (N_8490,N_7239,N_7346);
nand U8491 (N_8491,N_7171,N_7096);
xnor U8492 (N_8492,N_7581,N_7791);
and U8493 (N_8493,N_7948,N_7260);
xor U8494 (N_8494,N_7304,N_7318);
xnor U8495 (N_8495,N_7818,N_7054);
nor U8496 (N_8496,N_7353,N_7698);
xor U8497 (N_8497,N_7844,N_7843);
nor U8498 (N_8498,N_7971,N_7808);
nor U8499 (N_8499,N_7253,N_7646);
xor U8500 (N_8500,N_7161,N_7610);
nand U8501 (N_8501,N_7871,N_7760);
and U8502 (N_8502,N_7937,N_7781);
and U8503 (N_8503,N_7098,N_7559);
nand U8504 (N_8504,N_7326,N_7256);
nand U8505 (N_8505,N_7012,N_7331);
and U8506 (N_8506,N_7909,N_7036);
nand U8507 (N_8507,N_7326,N_7484);
or U8508 (N_8508,N_7746,N_7682);
and U8509 (N_8509,N_7893,N_7088);
and U8510 (N_8510,N_7369,N_7937);
or U8511 (N_8511,N_7638,N_7983);
and U8512 (N_8512,N_7332,N_7526);
and U8513 (N_8513,N_7640,N_7791);
nor U8514 (N_8514,N_7249,N_7136);
xnor U8515 (N_8515,N_7964,N_7698);
nor U8516 (N_8516,N_7441,N_7857);
nor U8517 (N_8517,N_7121,N_7498);
nor U8518 (N_8518,N_7013,N_7240);
nand U8519 (N_8519,N_7304,N_7908);
nand U8520 (N_8520,N_7682,N_7911);
xor U8521 (N_8521,N_7486,N_7234);
or U8522 (N_8522,N_7652,N_7339);
or U8523 (N_8523,N_7234,N_7386);
or U8524 (N_8524,N_7441,N_7980);
xor U8525 (N_8525,N_7038,N_7782);
and U8526 (N_8526,N_7280,N_7657);
nor U8527 (N_8527,N_7290,N_7179);
xor U8528 (N_8528,N_7146,N_7060);
or U8529 (N_8529,N_7600,N_7968);
or U8530 (N_8530,N_7098,N_7566);
and U8531 (N_8531,N_7685,N_7171);
nor U8532 (N_8532,N_7949,N_7039);
or U8533 (N_8533,N_7937,N_7147);
xor U8534 (N_8534,N_7176,N_7219);
and U8535 (N_8535,N_7873,N_7460);
nand U8536 (N_8536,N_7520,N_7629);
and U8537 (N_8537,N_7460,N_7249);
xor U8538 (N_8538,N_7170,N_7145);
nand U8539 (N_8539,N_7640,N_7535);
and U8540 (N_8540,N_7231,N_7759);
nand U8541 (N_8541,N_7079,N_7679);
or U8542 (N_8542,N_7248,N_7770);
or U8543 (N_8543,N_7666,N_7937);
nor U8544 (N_8544,N_7583,N_7856);
and U8545 (N_8545,N_7572,N_7553);
or U8546 (N_8546,N_7381,N_7421);
xnor U8547 (N_8547,N_7392,N_7475);
nor U8548 (N_8548,N_7120,N_7409);
and U8549 (N_8549,N_7388,N_7837);
and U8550 (N_8550,N_7191,N_7674);
xor U8551 (N_8551,N_7321,N_7616);
or U8552 (N_8552,N_7079,N_7540);
nor U8553 (N_8553,N_7854,N_7962);
and U8554 (N_8554,N_7560,N_7001);
xor U8555 (N_8555,N_7316,N_7231);
xnor U8556 (N_8556,N_7908,N_7089);
or U8557 (N_8557,N_7716,N_7288);
xor U8558 (N_8558,N_7210,N_7995);
or U8559 (N_8559,N_7712,N_7096);
or U8560 (N_8560,N_7458,N_7083);
and U8561 (N_8561,N_7264,N_7695);
nor U8562 (N_8562,N_7704,N_7879);
and U8563 (N_8563,N_7728,N_7766);
xor U8564 (N_8564,N_7921,N_7555);
and U8565 (N_8565,N_7036,N_7411);
nor U8566 (N_8566,N_7058,N_7903);
or U8567 (N_8567,N_7070,N_7356);
and U8568 (N_8568,N_7060,N_7736);
or U8569 (N_8569,N_7822,N_7254);
xnor U8570 (N_8570,N_7248,N_7606);
and U8571 (N_8571,N_7786,N_7370);
and U8572 (N_8572,N_7734,N_7345);
nand U8573 (N_8573,N_7146,N_7551);
xnor U8574 (N_8574,N_7795,N_7969);
and U8575 (N_8575,N_7986,N_7782);
xnor U8576 (N_8576,N_7881,N_7292);
or U8577 (N_8577,N_7532,N_7004);
and U8578 (N_8578,N_7203,N_7071);
xnor U8579 (N_8579,N_7593,N_7775);
or U8580 (N_8580,N_7431,N_7990);
nor U8581 (N_8581,N_7013,N_7581);
xor U8582 (N_8582,N_7294,N_7352);
nor U8583 (N_8583,N_7828,N_7564);
nor U8584 (N_8584,N_7414,N_7697);
or U8585 (N_8585,N_7498,N_7029);
xnor U8586 (N_8586,N_7259,N_7073);
nor U8587 (N_8587,N_7649,N_7328);
or U8588 (N_8588,N_7723,N_7832);
and U8589 (N_8589,N_7814,N_7975);
or U8590 (N_8590,N_7189,N_7735);
nand U8591 (N_8591,N_7865,N_7178);
or U8592 (N_8592,N_7951,N_7438);
nand U8593 (N_8593,N_7392,N_7789);
nand U8594 (N_8594,N_7804,N_7063);
and U8595 (N_8595,N_7516,N_7801);
and U8596 (N_8596,N_7391,N_7592);
and U8597 (N_8597,N_7577,N_7405);
xor U8598 (N_8598,N_7488,N_7832);
or U8599 (N_8599,N_7705,N_7118);
nor U8600 (N_8600,N_7010,N_7394);
or U8601 (N_8601,N_7991,N_7422);
and U8602 (N_8602,N_7486,N_7694);
xor U8603 (N_8603,N_7349,N_7627);
xnor U8604 (N_8604,N_7650,N_7860);
nor U8605 (N_8605,N_7034,N_7800);
xor U8606 (N_8606,N_7161,N_7056);
nand U8607 (N_8607,N_7060,N_7684);
nor U8608 (N_8608,N_7392,N_7037);
xor U8609 (N_8609,N_7248,N_7290);
xnor U8610 (N_8610,N_7776,N_7880);
nand U8611 (N_8611,N_7432,N_7261);
xor U8612 (N_8612,N_7140,N_7028);
nor U8613 (N_8613,N_7293,N_7965);
xnor U8614 (N_8614,N_7015,N_7175);
or U8615 (N_8615,N_7622,N_7347);
xnor U8616 (N_8616,N_7656,N_7512);
nand U8617 (N_8617,N_7394,N_7864);
xor U8618 (N_8618,N_7806,N_7610);
and U8619 (N_8619,N_7809,N_7915);
and U8620 (N_8620,N_7846,N_7739);
nor U8621 (N_8621,N_7454,N_7384);
xor U8622 (N_8622,N_7224,N_7890);
or U8623 (N_8623,N_7668,N_7131);
and U8624 (N_8624,N_7180,N_7471);
and U8625 (N_8625,N_7373,N_7071);
or U8626 (N_8626,N_7751,N_7680);
nand U8627 (N_8627,N_7714,N_7694);
nor U8628 (N_8628,N_7720,N_7414);
and U8629 (N_8629,N_7382,N_7788);
and U8630 (N_8630,N_7175,N_7324);
or U8631 (N_8631,N_7846,N_7867);
and U8632 (N_8632,N_7789,N_7713);
nand U8633 (N_8633,N_7606,N_7992);
nand U8634 (N_8634,N_7937,N_7702);
xnor U8635 (N_8635,N_7162,N_7398);
xor U8636 (N_8636,N_7045,N_7425);
nor U8637 (N_8637,N_7402,N_7310);
xor U8638 (N_8638,N_7425,N_7964);
nand U8639 (N_8639,N_7561,N_7201);
nor U8640 (N_8640,N_7916,N_7862);
nor U8641 (N_8641,N_7666,N_7971);
and U8642 (N_8642,N_7325,N_7326);
nand U8643 (N_8643,N_7557,N_7855);
xor U8644 (N_8644,N_7276,N_7358);
nand U8645 (N_8645,N_7923,N_7366);
nand U8646 (N_8646,N_7469,N_7517);
or U8647 (N_8647,N_7794,N_7391);
and U8648 (N_8648,N_7062,N_7144);
and U8649 (N_8649,N_7253,N_7478);
nand U8650 (N_8650,N_7044,N_7474);
or U8651 (N_8651,N_7794,N_7642);
or U8652 (N_8652,N_7204,N_7181);
or U8653 (N_8653,N_7016,N_7058);
xor U8654 (N_8654,N_7502,N_7925);
xnor U8655 (N_8655,N_7276,N_7647);
and U8656 (N_8656,N_7206,N_7139);
xor U8657 (N_8657,N_7270,N_7368);
nor U8658 (N_8658,N_7020,N_7480);
nor U8659 (N_8659,N_7690,N_7270);
or U8660 (N_8660,N_7850,N_7737);
nor U8661 (N_8661,N_7506,N_7643);
or U8662 (N_8662,N_7272,N_7205);
xor U8663 (N_8663,N_7016,N_7365);
or U8664 (N_8664,N_7361,N_7127);
nand U8665 (N_8665,N_7742,N_7797);
nand U8666 (N_8666,N_7896,N_7431);
or U8667 (N_8667,N_7001,N_7466);
nor U8668 (N_8668,N_7634,N_7236);
nor U8669 (N_8669,N_7534,N_7980);
or U8670 (N_8670,N_7661,N_7947);
nor U8671 (N_8671,N_7066,N_7858);
nand U8672 (N_8672,N_7303,N_7963);
nand U8673 (N_8673,N_7687,N_7747);
nor U8674 (N_8674,N_7560,N_7393);
or U8675 (N_8675,N_7919,N_7370);
nand U8676 (N_8676,N_7793,N_7936);
nand U8677 (N_8677,N_7845,N_7644);
xor U8678 (N_8678,N_7992,N_7541);
nor U8679 (N_8679,N_7785,N_7588);
nor U8680 (N_8680,N_7340,N_7382);
xor U8681 (N_8681,N_7346,N_7278);
or U8682 (N_8682,N_7864,N_7159);
or U8683 (N_8683,N_7344,N_7278);
nor U8684 (N_8684,N_7396,N_7263);
and U8685 (N_8685,N_7994,N_7564);
or U8686 (N_8686,N_7610,N_7882);
and U8687 (N_8687,N_7716,N_7764);
or U8688 (N_8688,N_7561,N_7495);
xnor U8689 (N_8689,N_7771,N_7914);
nand U8690 (N_8690,N_7672,N_7428);
nand U8691 (N_8691,N_7710,N_7629);
nor U8692 (N_8692,N_7183,N_7191);
nand U8693 (N_8693,N_7063,N_7850);
or U8694 (N_8694,N_7698,N_7175);
nor U8695 (N_8695,N_7325,N_7750);
nor U8696 (N_8696,N_7936,N_7273);
or U8697 (N_8697,N_7871,N_7609);
nand U8698 (N_8698,N_7039,N_7844);
xor U8699 (N_8699,N_7824,N_7643);
and U8700 (N_8700,N_7497,N_7969);
nand U8701 (N_8701,N_7747,N_7471);
nand U8702 (N_8702,N_7896,N_7744);
and U8703 (N_8703,N_7544,N_7346);
xnor U8704 (N_8704,N_7632,N_7180);
or U8705 (N_8705,N_7793,N_7324);
nor U8706 (N_8706,N_7584,N_7390);
nor U8707 (N_8707,N_7255,N_7790);
nand U8708 (N_8708,N_7962,N_7814);
nand U8709 (N_8709,N_7167,N_7599);
nor U8710 (N_8710,N_7059,N_7845);
xnor U8711 (N_8711,N_7964,N_7973);
and U8712 (N_8712,N_7010,N_7180);
xnor U8713 (N_8713,N_7760,N_7286);
nand U8714 (N_8714,N_7505,N_7018);
xor U8715 (N_8715,N_7292,N_7309);
nor U8716 (N_8716,N_7054,N_7223);
or U8717 (N_8717,N_7001,N_7844);
xnor U8718 (N_8718,N_7252,N_7404);
or U8719 (N_8719,N_7728,N_7067);
and U8720 (N_8720,N_7086,N_7083);
or U8721 (N_8721,N_7801,N_7530);
nand U8722 (N_8722,N_7759,N_7016);
and U8723 (N_8723,N_7732,N_7653);
nand U8724 (N_8724,N_7101,N_7062);
and U8725 (N_8725,N_7385,N_7510);
xor U8726 (N_8726,N_7030,N_7865);
and U8727 (N_8727,N_7242,N_7017);
nand U8728 (N_8728,N_7860,N_7165);
xnor U8729 (N_8729,N_7110,N_7580);
nand U8730 (N_8730,N_7825,N_7236);
nand U8731 (N_8731,N_7677,N_7848);
and U8732 (N_8732,N_7242,N_7110);
and U8733 (N_8733,N_7893,N_7617);
and U8734 (N_8734,N_7394,N_7881);
nand U8735 (N_8735,N_7273,N_7904);
xnor U8736 (N_8736,N_7536,N_7601);
or U8737 (N_8737,N_7136,N_7830);
and U8738 (N_8738,N_7388,N_7135);
or U8739 (N_8739,N_7936,N_7738);
and U8740 (N_8740,N_7076,N_7655);
xnor U8741 (N_8741,N_7586,N_7848);
nand U8742 (N_8742,N_7435,N_7145);
xor U8743 (N_8743,N_7712,N_7607);
nor U8744 (N_8744,N_7622,N_7792);
or U8745 (N_8745,N_7232,N_7064);
nor U8746 (N_8746,N_7137,N_7417);
nor U8747 (N_8747,N_7128,N_7474);
xor U8748 (N_8748,N_7886,N_7496);
xor U8749 (N_8749,N_7374,N_7617);
or U8750 (N_8750,N_7708,N_7947);
and U8751 (N_8751,N_7207,N_7639);
or U8752 (N_8752,N_7258,N_7361);
xor U8753 (N_8753,N_7284,N_7016);
and U8754 (N_8754,N_7921,N_7345);
or U8755 (N_8755,N_7075,N_7461);
nand U8756 (N_8756,N_7114,N_7950);
nand U8757 (N_8757,N_7607,N_7891);
xor U8758 (N_8758,N_7621,N_7786);
xor U8759 (N_8759,N_7364,N_7616);
xnor U8760 (N_8760,N_7518,N_7255);
nand U8761 (N_8761,N_7070,N_7676);
and U8762 (N_8762,N_7255,N_7239);
nand U8763 (N_8763,N_7092,N_7399);
and U8764 (N_8764,N_7209,N_7212);
and U8765 (N_8765,N_7407,N_7579);
nand U8766 (N_8766,N_7201,N_7260);
and U8767 (N_8767,N_7383,N_7738);
or U8768 (N_8768,N_7555,N_7653);
nor U8769 (N_8769,N_7643,N_7287);
and U8770 (N_8770,N_7373,N_7923);
and U8771 (N_8771,N_7789,N_7787);
nand U8772 (N_8772,N_7445,N_7697);
nor U8773 (N_8773,N_7675,N_7842);
and U8774 (N_8774,N_7839,N_7083);
and U8775 (N_8775,N_7090,N_7857);
nor U8776 (N_8776,N_7501,N_7361);
nor U8777 (N_8777,N_7104,N_7666);
xnor U8778 (N_8778,N_7441,N_7344);
nand U8779 (N_8779,N_7839,N_7638);
xnor U8780 (N_8780,N_7635,N_7538);
nor U8781 (N_8781,N_7682,N_7498);
or U8782 (N_8782,N_7561,N_7884);
and U8783 (N_8783,N_7470,N_7841);
or U8784 (N_8784,N_7766,N_7921);
nor U8785 (N_8785,N_7051,N_7669);
nand U8786 (N_8786,N_7422,N_7797);
or U8787 (N_8787,N_7349,N_7354);
nor U8788 (N_8788,N_7884,N_7302);
or U8789 (N_8789,N_7444,N_7184);
xnor U8790 (N_8790,N_7892,N_7038);
xnor U8791 (N_8791,N_7520,N_7397);
or U8792 (N_8792,N_7547,N_7211);
and U8793 (N_8793,N_7948,N_7853);
nor U8794 (N_8794,N_7928,N_7503);
nor U8795 (N_8795,N_7631,N_7053);
or U8796 (N_8796,N_7460,N_7975);
and U8797 (N_8797,N_7948,N_7547);
nor U8798 (N_8798,N_7117,N_7213);
nand U8799 (N_8799,N_7850,N_7179);
and U8800 (N_8800,N_7580,N_7047);
nor U8801 (N_8801,N_7685,N_7308);
nor U8802 (N_8802,N_7947,N_7879);
nand U8803 (N_8803,N_7090,N_7601);
or U8804 (N_8804,N_7093,N_7891);
nand U8805 (N_8805,N_7888,N_7802);
nand U8806 (N_8806,N_7013,N_7452);
xnor U8807 (N_8807,N_7294,N_7948);
xor U8808 (N_8808,N_7020,N_7772);
nand U8809 (N_8809,N_7323,N_7277);
nand U8810 (N_8810,N_7666,N_7906);
and U8811 (N_8811,N_7544,N_7040);
nor U8812 (N_8812,N_7852,N_7960);
nand U8813 (N_8813,N_7657,N_7756);
xnor U8814 (N_8814,N_7188,N_7712);
and U8815 (N_8815,N_7743,N_7343);
or U8816 (N_8816,N_7399,N_7262);
and U8817 (N_8817,N_7343,N_7622);
xor U8818 (N_8818,N_7531,N_7432);
nand U8819 (N_8819,N_7521,N_7746);
or U8820 (N_8820,N_7819,N_7877);
nor U8821 (N_8821,N_7079,N_7111);
or U8822 (N_8822,N_7178,N_7821);
nand U8823 (N_8823,N_7471,N_7390);
nor U8824 (N_8824,N_7958,N_7768);
xor U8825 (N_8825,N_7865,N_7778);
nand U8826 (N_8826,N_7678,N_7136);
xnor U8827 (N_8827,N_7853,N_7941);
nor U8828 (N_8828,N_7785,N_7223);
and U8829 (N_8829,N_7313,N_7879);
or U8830 (N_8830,N_7512,N_7699);
xnor U8831 (N_8831,N_7135,N_7138);
nor U8832 (N_8832,N_7706,N_7275);
and U8833 (N_8833,N_7128,N_7598);
xnor U8834 (N_8834,N_7756,N_7301);
or U8835 (N_8835,N_7743,N_7546);
xor U8836 (N_8836,N_7159,N_7101);
xor U8837 (N_8837,N_7252,N_7049);
and U8838 (N_8838,N_7331,N_7417);
and U8839 (N_8839,N_7570,N_7727);
xor U8840 (N_8840,N_7596,N_7809);
xor U8841 (N_8841,N_7759,N_7269);
xnor U8842 (N_8842,N_7933,N_7911);
or U8843 (N_8843,N_7630,N_7990);
nand U8844 (N_8844,N_7264,N_7409);
nor U8845 (N_8845,N_7270,N_7987);
nor U8846 (N_8846,N_7992,N_7084);
nand U8847 (N_8847,N_7909,N_7269);
and U8848 (N_8848,N_7278,N_7256);
nor U8849 (N_8849,N_7547,N_7617);
or U8850 (N_8850,N_7477,N_7091);
or U8851 (N_8851,N_7531,N_7414);
xnor U8852 (N_8852,N_7587,N_7195);
and U8853 (N_8853,N_7943,N_7531);
or U8854 (N_8854,N_7771,N_7880);
nor U8855 (N_8855,N_7628,N_7685);
and U8856 (N_8856,N_7866,N_7132);
xnor U8857 (N_8857,N_7763,N_7729);
and U8858 (N_8858,N_7425,N_7316);
nand U8859 (N_8859,N_7656,N_7818);
nand U8860 (N_8860,N_7136,N_7398);
xnor U8861 (N_8861,N_7079,N_7708);
xor U8862 (N_8862,N_7356,N_7388);
xor U8863 (N_8863,N_7389,N_7870);
or U8864 (N_8864,N_7165,N_7850);
xnor U8865 (N_8865,N_7544,N_7156);
nand U8866 (N_8866,N_7002,N_7680);
nor U8867 (N_8867,N_7811,N_7173);
nor U8868 (N_8868,N_7065,N_7599);
or U8869 (N_8869,N_7495,N_7385);
and U8870 (N_8870,N_7064,N_7478);
nand U8871 (N_8871,N_7603,N_7992);
nand U8872 (N_8872,N_7755,N_7936);
xor U8873 (N_8873,N_7233,N_7515);
xor U8874 (N_8874,N_7488,N_7208);
or U8875 (N_8875,N_7646,N_7034);
xor U8876 (N_8876,N_7901,N_7408);
or U8877 (N_8877,N_7325,N_7053);
or U8878 (N_8878,N_7570,N_7711);
nor U8879 (N_8879,N_7592,N_7125);
and U8880 (N_8880,N_7690,N_7192);
and U8881 (N_8881,N_7486,N_7515);
xor U8882 (N_8882,N_7109,N_7849);
or U8883 (N_8883,N_7434,N_7579);
nor U8884 (N_8884,N_7309,N_7150);
and U8885 (N_8885,N_7017,N_7666);
or U8886 (N_8886,N_7235,N_7427);
and U8887 (N_8887,N_7385,N_7529);
or U8888 (N_8888,N_7207,N_7491);
xor U8889 (N_8889,N_7582,N_7799);
nand U8890 (N_8890,N_7511,N_7556);
nor U8891 (N_8891,N_7884,N_7183);
or U8892 (N_8892,N_7618,N_7398);
xor U8893 (N_8893,N_7119,N_7922);
nand U8894 (N_8894,N_7746,N_7102);
and U8895 (N_8895,N_7919,N_7995);
xnor U8896 (N_8896,N_7289,N_7497);
xnor U8897 (N_8897,N_7365,N_7348);
xnor U8898 (N_8898,N_7617,N_7424);
nand U8899 (N_8899,N_7561,N_7923);
nand U8900 (N_8900,N_7603,N_7735);
or U8901 (N_8901,N_7005,N_7502);
nand U8902 (N_8902,N_7748,N_7185);
nand U8903 (N_8903,N_7921,N_7847);
or U8904 (N_8904,N_7707,N_7644);
nand U8905 (N_8905,N_7212,N_7697);
xor U8906 (N_8906,N_7255,N_7602);
or U8907 (N_8907,N_7867,N_7216);
and U8908 (N_8908,N_7577,N_7548);
nor U8909 (N_8909,N_7106,N_7157);
nor U8910 (N_8910,N_7830,N_7845);
nor U8911 (N_8911,N_7012,N_7727);
or U8912 (N_8912,N_7047,N_7766);
and U8913 (N_8913,N_7751,N_7224);
nand U8914 (N_8914,N_7021,N_7788);
or U8915 (N_8915,N_7807,N_7639);
or U8916 (N_8916,N_7194,N_7864);
and U8917 (N_8917,N_7683,N_7428);
nand U8918 (N_8918,N_7183,N_7016);
xor U8919 (N_8919,N_7275,N_7524);
or U8920 (N_8920,N_7483,N_7528);
nor U8921 (N_8921,N_7172,N_7221);
and U8922 (N_8922,N_7016,N_7042);
and U8923 (N_8923,N_7915,N_7122);
xnor U8924 (N_8924,N_7958,N_7308);
xor U8925 (N_8925,N_7541,N_7570);
or U8926 (N_8926,N_7073,N_7866);
or U8927 (N_8927,N_7390,N_7101);
nor U8928 (N_8928,N_7745,N_7715);
xnor U8929 (N_8929,N_7821,N_7912);
nor U8930 (N_8930,N_7551,N_7156);
nand U8931 (N_8931,N_7546,N_7003);
xor U8932 (N_8932,N_7954,N_7842);
nand U8933 (N_8933,N_7824,N_7128);
and U8934 (N_8934,N_7004,N_7872);
or U8935 (N_8935,N_7582,N_7243);
nor U8936 (N_8936,N_7661,N_7541);
or U8937 (N_8937,N_7537,N_7797);
or U8938 (N_8938,N_7276,N_7139);
xnor U8939 (N_8939,N_7410,N_7032);
xnor U8940 (N_8940,N_7891,N_7835);
nor U8941 (N_8941,N_7820,N_7423);
or U8942 (N_8942,N_7470,N_7387);
xnor U8943 (N_8943,N_7818,N_7356);
and U8944 (N_8944,N_7789,N_7464);
or U8945 (N_8945,N_7721,N_7211);
or U8946 (N_8946,N_7981,N_7112);
or U8947 (N_8947,N_7600,N_7917);
nand U8948 (N_8948,N_7299,N_7673);
and U8949 (N_8949,N_7548,N_7933);
and U8950 (N_8950,N_7117,N_7024);
nand U8951 (N_8951,N_7313,N_7591);
nor U8952 (N_8952,N_7206,N_7768);
or U8953 (N_8953,N_7521,N_7630);
nand U8954 (N_8954,N_7974,N_7704);
nand U8955 (N_8955,N_7655,N_7950);
or U8956 (N_8956,N_7011,N_7716);
or U8957 (N_8957,N_7858,N_7831);
xnor U8958 (N_8958,N_7072,N_7769);
or U8959 (N_8959,N_7611,N_7386);
nand U8960 (N_8960,N_7518,N_7078);
and U8961 (N_8961,N_7446,N_7436);
or U8962 (N_8962,N_7192,N_7724);
nand U8963 (N_8963,N_7632,N_7077);
or U8964 (N_8964,N_7917,N_7200);
nor U8965 (N_8965,N_7756,N_7556);
nand U8966 (N_8966,N_7623,N_7651);
xnor U8967 (N_8967,N_7077,N_7483);
nand U8968 (N_8968,N_7393,N_7283);
or U8969 (N_8969,N_7107,N_7728);
or U8970 (N_8970,N_7730,N_7547);
or U8971 (N_8971,N_7769,N_7722);
and U8972 (N_8972,N_7307,N_7423);
xor U8973 (N_8973,N_7119,N_7484);
xnor U8974 (N_8974,N_7879,N_7646);
nor U8975 (N_8975,N_7408,N_7518);
and U8976 (N_8976,N_7751,N_7774);
nor U8977 (N_8977,N_7730,N_7173);
nor U8978 (N_8978,N_7804,N_7360);
or U8979 (N_8979,N_7091,N_7341);
xnor U8980 (N_8980,N_7971,N_7909);
xnor U8981 (N_8981,N_7450,N_7894);
nor U8982 (N_8982,N_7509,N_7009);
xor U8983 (N_8983,N_7732,N_7872);
xnor U8984 (N_8984,N_7062,N_7543);
xnor U8985 (N_8985,N_7731,N_7903);
xnor U8986 (N_8986,N_7428,N_7775);
or U8987 (N_8987,N_7927,N_7479);
nand U8988 (N_8988,N_7303,N_7039);
xnor U8989 (N_8989,N_7958,N_7343);
nor U8990 (N_8990,N_7208,N_7262);
xor U8991 (N_8991,N_7017,N_7157);
or U8992 (N_8992,N_7759,N_7055);
or U8993 (N_8993,N_7566,N_7475);
nand U8994 (N_8994,N_7520,N_7577);
xor U8995 (N_8995,N_7753,N_7606);
xor U8996 (N_8996,N_7865,N_7851);
nor U8997 (N_8997,N_7568,N_7920);
and U8998 (N_8998,N_7543,N_7028);
and U8999 (N_8999,N_7134,N_7719);
xor U9000 (N_9000,N_8980,N_8153);
nand U9001 (N_9001,N_8826,N_8578);
and U9002 (N_9002,N_8257,N_8147);
xnor U9003 (N_9003,N_8871,N_8188);
nor U9004 (N_9004,N_8545,N_8311);
or U9005 (N_9005,N_8315,N_8873);
nand U9006 (N_9006,N_8269,N_8998);
nand U9007 (N_9007,N_8466,N_8833);
and U9008 (N_9008,N_8403,N_8189);
or U9009 (N_9009,N_8222,N_8652);
and U9010 (N_9010,N_8192,N_8672);
and U9011 (N_9011,N_8174,N_8406);
nor U9012 (N_9012,N_8393,N_8777);
xor U9013 (N_9013,N_8896,N_8863);
or U9014 (N_9014,N_8358,N_8342);
nand U9015 (N_9015,N_8436,N_8558);
xor U9016 (N_9016,N_8015,N_8927);
nor U9017 (N_9017,N_8041,N_8682);
nor U9018 (N_9018,N_8533,N_8537);
nor U9019 (N_9019,N_8446,N_8650);
or U9020 (N_9020,N_8207,N_8888);
nor U9021 (N_9021,N_8542,N_8094);
or U9022 (N_9022,N_8331,N_8078);
nand U9023 (N_9023,N_8335,N_8547);
or U9024 (N_9024,N_8685,N_8474);
nor U9025 (N_9025,N_8934,N_8375);
or U9026 (N_9026,N_8908,N_8928);
and U9027 (N_9027,N_8017,N_8462);
nand U9028 (N_9028,N_8390,N_8302);
and U9029 (N_9029,N_8384,N_8572);
or U9030 (N_9030,N_8352,N_8385);
nand U9031 (N_9031,N_8540,N_8037);
nor U9032 (N_9032,N_8840,N_8471);
nor U9033 (N_9033,N_8936,N_8396);
or U9034 (N_9034,N_8503,N_8012);
or U9035 (N_9035,N_8283,N_8185);
nor U9036 (N_9036,N_8623,N_8963);
or U9037 (N_9037,N_8589,N_8664);
nand U9038 (N_9038,N_8325,N_8307);
nand U9039 (N_9039,N_8870,N_8782);
nor U9040 (N_9040,N_8836,N_8258);
or U9041 (N_9041,N_8292,N_8439);
and U9042 (N_9042,N_8831,N_8573);
or U9043 (N_9043,N_8250,N_8555);
or U9044 (N_9044,N_8932,N_8444);
nor U9045 (N_9045,N_8556,N_8778);
and U9046 (N_9046,N_8918,N_8214);
and U9047 (N_9047,N_8955,N_8075);
and U9048 (N_9048,N_8841,N_8148);
and U9049 (N_9049,N_8818,N_8554);
or U9050 (N_9050,N_8334,N_8628);
nand U9051 (N_9051,N_8365,N_8452);
nand U9052 (N_9052,N_8267,N_8971);
nand U9053 (N_9053,N_8590,N_8976);
nand U9054 (N_9054,N_8284,N_8518);
and U9055 (N_9055,N_8925,N_8990);
nor U9056 (N_9056,N_8392,N_8044);
or U9057 (N_9057,N_8100,N_8662);
and U9058 (N_9058,N_8988,N_8780);
nand U9059 (N_9059,N_8241,N_8160);
nand U9060 (N_9060,N_8536,N_8033);
nand U9061 (N_9061,N_8023,N_8411);
nor U9062 (N_9062,N_8900,N_8089);
nand U9063 (N_9063,N_8171,N_8243);
nor U9064 (N_9064,N_8730,N_8473);
or U9065 (N_9065,N_8637,N_8561);
xnor U9066 (N_9066,N_8395,N_8585);
xor U9067 (N_9067,N_8799,N_8217);
nor U9068 (N_9068,N_8176,N_8433);
xor U9069 (N_9069,N_8356,N_8271);
nand U9070 (N_9070,N_8613,N_8586);
or U9071 (N_9071,N_8909,N_8186);
xnor U9072 (N_9072,N_8801,N_8642);
xnor U9073 (N_9073,N_8931,N_8611);
nand U9074 (N_9074,N_8666,N_8180);
xor U9075 (N_9075,N_8118,N_8000);
nor U9076 (N_9076,N_8197,N_8600);
nor U9077 (N_9077,N_8061,N_8647);
nand U9078 (N_9078,N_8467,N_8839);
xor U9079 (N_9079,N_8592,N_8952);
xnor U9080 (N_9080,N_8701,N_8134);
and U9081 (N_9081,N_8301,N_8596);
or U9082 (N_9082,N_8785,N_8773);
or U9083 (N_9083,N_8454,N_8242);
nand U9084 (N_9084,N_8417,N_8743);
xor U9085 (N_9085,N_8654,N_8512);
and U9086 (N_9086,N_8245,N_8796);
xnor U9087 (N_9087,N_8762,N_8771);
and U9088 (N_9088,N_8622,N_8786);
or U9089 (N_9089,N_8373,N_8739);
or U9090 (N_9090,N_8420,N_8904);
nand U9091 (N_9091,N_8804,N_8032);
and U9092 (N_9092,N_8853,N_8725);
nor U9093 (N_9093,N_8665,N_8506);
xor U9094 (N_9094,N_8312,N_8294);
xnor U9095 (N_9095,N_8318,N_8101);
nor U9096 (N_9096,N_8351,N_8478);
and U9097 (N_9097,N_8337,N_8793);
nor U9098 (N_9098,N_8322,N_8570);
xor U9099 (N_9099,N_8391,N_8571);
nand U9100 (N_9100,N_8003,N_8475);
nand U9101 (N_9101,N_8263,N_8830);
and U9102 (N_9102,N_8499,N_8865);
nor U9103 (N_9103,N_8477,N_8768);
nor U9104 (N_9104,N_8869,N_8995);
xnor U9105 (N_9105,N_8155,N_8259);
or U9106 (N_9106,N_8149,N_8133);
or U9107 (N_9107,N_8750,N_8880);
xnor U9108 (N_9108,N_8047,N_8710);
nor U9109 (N_9109,N_8899,N_8834);
xnor U9110 (N_9110,N_8016,N_8889);
or U9111 (N_9111,N_8878,N_8563);
nand U9112 (N_9112,N_8868,N_8159);
or U9113 (N_9113,N_8681,N_8519);
and U9114 (N_9114,N_8922,N_8484);
xor U9115 (N_9115,N_8445,N_8265);
and U9116 (N_9116,N_8707,N_8313);
or U9117 (N_9117,N_8663,N_8615);
and U9118 (N_9118,N_8107,N_8150);
or U9119 (N_9119,N_8758,N_8703);
nand U9120 (N_9120,N_8848,N_8734);
nand U9121 (N_9121,N_8635,N_8143);
xor U9122 (N_9122,N_8125,N_8847);
nand U9123 (N_9123,N_8735,N_8168);
and U9124 (N_9124,N_8225,N_8116);
nand U9125 (N_9125,N_8923,N_8906);
and U9126 (N_9126,N_8961,N_8670);
xnor U9127 (N_9127,N_8949,N_8805);
and U9128 (N_9128,N_8985,N_8668);
or U9129 (N_9129,N_8208,N_8580);
and U9130 (N_9130,N_8689,N_8649);
xnor U9131 (N_9131,N_8993,N_8601);
nor U9132 (N_9132,N_8309,N_8915);
nor U9133 (N_9133,N_8086,N_8367);
nand U9134 (N_9134,N_8169,N_8942);
or U9135 (N_9135,N_8526,N_8718);
and U9136 (N_9136,N_8253,N_8146);
and U9137 (N_9137,N_8497,N_8212);
and U9138 (N_9138,N_8066,N_8442);
nor U9139 (N_9139,N_8014,N_8659);
xor U9140 (N_9140,N_8109,N_8708);
or U9141 (N_9141,N_8178,N_8379);
nand U9142 (N_9142,N_8717,N_8233);
and U9143 (N_9143,N_8280,N_8678);
nand U9144 (N_9144,N_8595,N_8428);
or U9145 (N_9145,N_8820,N_8553);
and U9146 (N_9146,N_8761,N_8053);
nand U9147 (N_9147,N_8892,N_8291);
xnor U9148 (N_9148,N_8073,N_8684);
xor U9149 (N_9149,N_8864,N_8527);
or U9150 (N_9150,N_8644,N_8330);
and U9151 (N_9151,N_8485,N_8509);
nor U9152 (N_9152,N_8803,N_8326);
nor U9153 (N_9153,N_8097,N_8005);
nand U9154 (N_9154,N_8562,N_8256);
nand U9155 (N_9155,N_8247,N_8369);
and U9156 (N_9156,N_8057,N_8631);
or U9157 (N_9157,N_8354,N_8093);
nor U9158 (N_9158,N_8103,N_8851);
nor U9159 (N_9159,N_8724,N_8597);
nor U9160 (N_9160,N_8599,N_8425);
nor U9161 (N_9161,N_8039,N_8106);
and U9162 (N_9162,N_8400,N_8190);
xor U9163 (N_9163,N_8310,N_8363);
and U9164 (N_9164,N_8860,N_8657);
xor U9165 (N_9165,N_8151,N_8494);
or U9166 (N_9166,N_8898,N_8164);
xor U9167 (N_9167,N_8856,N_8745);
nor U9168 (N_9168,N_8639,N_8544);
xnor U9169 (N_9169,N_8418,N_8779);
and U9170 (N_9170,N_8885,N_8756);
nand U9171 (N_9171,N_8386,N_8849);
and U9172 (N_9172,N_8062,N_8360);
nand U9173 (N_9173,N_8970,N_8121);
or U9174 (N_9174,N_8842,N_8213);
nor U9175 (N_9175,N_8574,N_8427);
xnor U9176 (N_9176,N_8809,N_8721);
xnor U9177 (N_9177,N_8587,N_8531);
nand U9178 (N_9178,N_8045,N_8127);
xor U9179 (N_9179,N_8646,N_8007);
xor U9180 (N_9180,N_8946,N_8626);
and U9181 (N_9181,N_8308,N_8316);
and U9182 (N_9182,N_8594,N_8472);
xnor U9183 (N_9183,N_8449,N_8429);
xnor U9184 (N_9184,N_8319,N_8832);
nand U9185 (N_9185,N_8481,N_8591);
xnor U9186 (N_9186,N_8953,N_8223);
nor U9187 (N_9187,N_8722,N_8054);
nor U9188 (N_9188,N_8002,N_8557);
nand U9189 (N_9189,N_8343,N_8237);
and U9190 (N_9190,N_8096,N_8763);
or U9191 (N_9191,N_8479,N_8432);
nor U9192 (N_9192,N_8890,N_8539);
and U9193 (N_9193,N_8364,N_8857);
nand U9194 (N_9194,N_8490,N_8397);
xor U9195 (N_9195,N_8877,N_8424);
and U9196 (N_9196,N_8059,N_8251);
nor U9197 (N_9197,N_8776,N_8177);
nor U9198 (N_9198,N_8610,N_8167);
or U9199 (N_9199,N_8549,N_8141);
nand U9200 (N_9200,N_8859,N_8683);
or U9201 (N_9201,N_8850,N_8104);
nand U9202 (N_9202,N_8112,N_8769);
or U9203 (N_9203,N_8951,N_8671);
nor U9204 (N_9204,N_8320,N_8691);
and U9205 (N_9205,N_8907,N_8117);
xor U9206 (N_9206,N_8370,N_8027);
or U9207 (N_9207,N_8731,N_8784);
and U9208 (N_9208,N_8248,N_8766);
and U9209 (N_9209,N_8366,N_8043);
and U9210 (N_9210,N_8607,N_8740);
xor U9211 (N_9211,N_8377,N_8145);
and U9212 (N_9212,N_8690,N_8273);
xor U9213 (N_9213,N_8938,N_8279);
xor U9214 (N_9214,N_8161,N_8108);
xnor U9215 (N_9215,N_8855,N_8119);
xor U9216 (N_9216,N_8618,N_8866);
xor U9217 (N_9217,N_8434,N_8088);
xnor U9218 (N_9218,N_8969,N_8426);
nand U9219 (N_9219,N_8603,N_8696);
nand U9220 (N_9220,N_8341,N_8838);
nor U9221 (N_9221,N_8193,N_8220);
nor U9222 (N_9222,N_8872,N_8825);
or U9223 (N_9223,N_8443,N_8297);
nand U9224 (N_9224,N_8797,N_8300);
nand U9225 (N_9225,N_8501,N_8902);
nand U9226 (N_9226,N_8021,N_8548);
or U9227 (N_9227,N_8939,N_8378);
and U9228 (N_9228,N_8276,N_8828);
nand U9229 (N_9229,N_8653,N_8688);
nand U9230 (N_9230,N_8274,N_8152);
and U9231 (N_9231,N_8465,N_8974);
nand U9232 (N_9232,N_8287,N_8566);
nand U9233 (N_9233,N_8964,N_8800);
nand U9234 (N_9234,N_8226,N_8254);
and U9235 (N_9235,N_8272,N_8440);
or U9236 (N_9236,N_8231,N_8099);
xnor U9237 (N_9237,N_8450,N_8098);
and U9238 (N_9238,N_8072,N_8741);
nor U9239 (N_9239,N_8948,N_8565);
xnor U9240 (N_9240,N_8867,N_8227);
or U9241 (N_9241,N_8068,N_8144);
xor U9242 (N_9242,N_8285,N_8264);
nor U9243 (N_9243,N_8410,N_8959);
nand U9244 (N_9244,N_8744,N_8447);
xnor U9245 (N_9245,N_8698,N_8030);
and U9246 (N_9246,N_8203,N_8543);
or U9247 (N_9247,N_8846,N_8401);
and U9248 (N_9248,N_8092,N_8598);
nand U9249 (N_9249,N_8994,N_8609);
or U9250 (N_9250,N_8667,N_8764);
nand U9251 (N_9251,N_8042,N_8581);
nand U9252 (N_9252,N_8306,N_8323);
xor U9253 (N_9253,N_8704,N_8064);
nor U9254 (N_9254,N_8338,N_8070);
or U9255 (N_9255,N_8055,N_8438);
nor U9256 (N_9256,N_8700,N_8984);
xor U9257 (N_9257,N_8945,N_8036);
or U9258 (N_9258,N_8051,N_8230);
nand U9259 (N_9259,N_8702,N_8920);
xnor U9260 (N_9260,N_8025,N_8448);
xnor U9261 (N_9261,N_8232,N_8669);
and U9262 (N_9262,N_8944,N_8034);
nor U9263 (N_9263,N_8175,N_8605);
or U9264 (N_9264,N_8077,N_8380);
or U9265 (N_9265,N_8080,N_8504);
nor U9266 (N_9266,N_8202,N_8720);
or U9267 (N_9267,N_8388,N_8480);
xnor U9268 (N_9268,N_8627,N_8024);
or U9269 (N_9269,N_8924,N_8625);
nand U9270 (N_9270,N_8071,N_8911);
xnor U9271 (N_9271,N_8339,N_8505);
nand U9272 (N_9272,N_8290,N_8960);
xor U9273 (N_9273,N_8975,N_8751);
nor U9274 (N_9274,N_8583,N_8421);
or U9275 (N_9275,N_8348,N_8435);
nand U9276 (N_9276,N_8852,N_8895);
nor U9277 (N_9277,N_8978,N_8018);
or U9278 (N_9278,N_8694,N_8082);
or U9279 (N_9279,N_8201,N_8063);
nor U9280 (N_9280,N_8381,N_8268);
nor U9281 (N_9281,N_8409,N_8602);
or U9282 (N_9282,N_8110,N_8011);
or U9283 (N_9283,N_8737,N_8333);
nand U9284 (N_9284,N_8496,N_8551);
xor U9285 (N_9285,N_8541,N_8755);
xor U9286 (N_9286,N_8712,N_8713);
and U9287 (N_9287,N_8382,N_8514);
and U9288 (N_9288,N_8136,N_8131);
nand U9289 (N_9289,N_8843,N_8781);
nand U9290 (N_9290,N_8619,N_8115);
nor U9291 (N_9291,N_8636,N_8977);
xnor U9292 (N_9292,N_8461,N_8759);
xnor U9293 (N_9293,N_8729,N_8965);
or U9294 (N_9294,N_8732,N_8726);
and U9295 (N_9295,N_8791,N_8753);
xnor U9296 (N_9296,N_8194,N_8087);
xnor U9297 (N_9297,N_8983,N_8022);
and U9298 (N_9298,N_8184,N_8124);
nor U9299 (N_9299,N_8216,N_8031);
nand U9300 (N_9300,N_8181,N_8821);
nor U9301 (N_9301,N_8522,N_8081);
nand U9302 (N_9302,N_8827,N_8048);
or U9303 (N_9303,N_8204,N_8822);
and U9304 (N_9304,N_8361,N_8026);
xor U9305 (N_9305,N_8001,N_8278);
and U9306 (N_9306,N_8930,N_8612);
nand U9307 (N_9307,N_8957,N_8742);
and U9308 (N_9308,N_8244,N_8028);
or U9309 (N_9309,N_8328,N_8530);
or U9310 (N_9310,N_8559,N_8486);
or U9311 (N_9311,N_8588,N_8065);
nor U9312 (N_9312,N_8170,N_8238);
nand U9313 (N_9313,N_8528,N_8714);
xnor U9314 (N_9314,N_8837,N_8643);
nand U9315 (N_9315,N_8538,N_8535);
xor U9316 (N_9316,N_8747,N_8288);
and U9317 (N_9317,N_8495,N_8673);
nor U9318 (N_9318,N_8933,N_8645);
and U9319 (N_9319,N_8638,N_8179);
nand U9320 (N_9320,N_8534,N_8329);
nor U9321 (N_9321,N_8355,N_8459);
and U9322 (N_9322,N_8376,N_8680);
nand U9323 (N_9323,N_8321,N_8138);
nor U9324 (N_9324,N_8058,N_8183);
and U9325 (N_9325,N_8723,N_8719);
nand U9326 (N_9326,N_8372,N_8236);
and U9327 (N_9327,N_8491,N_8399);
and U9328 (N_9328,N_8415,N_8277);
or U9329 (N_9329,N_8488,N_8286);
and U9330 (N_9330,N_8982,N_8861);
nor U9331 (N_9331,N_8903,N_8817);
and U9332 (N_9332,N_8529,N_8293);
or U9333 (N_9333,N_8234,N_8987);
nor U9334 (N_9334,N_8137,N_8757);
or U9335 (N_9335,N_8422,N_8575);
xnor U9336 (N_9336,N_8845,N_8387);
nand U9337 (N_9337,N_8733,N_8617);
xor U9338 (N_9338,N_8783,N_8517);
nand U9339 (N_9339,N_8897,N_8229);
and U9340 (N_9340,N_8416,N_8616);
xnor U9341 (N_9341,N_8568,N_8651);
xnor U9342 (N_9342,N_8324,N_8076);
and U9343 (N_9343,N_8632,N_8844);
nor U9344 (N_9344,N_8402,N_8235);
nand U9345 (N_9345,N_8196,N_8629);
and U9346 (N_9346,N_8887,N_8476);
or U9347 (N_9347,N_8489,N_8879);
nand U9348 (N_9348,N_8921,N_8579);
nand U9349 (N_9349,N_8430,N_8973);
and U9350 (N_9350,N_8981,N_8997);
xnor U9351 (N_9351,N_8139,N_8788);
nor U9352 (N_9352,N_8947,N_8345);
nor U9353 (N_9353,N_8128,N_8606);
nor U9354 (N_9354,N_8362,N_8413);
or U9355 (N_9355,N_8305,N_8508);
nor U9356 (N_9356,N_8327,N_8239);
and U9357 (N_9357,N_8687,N_8142);
and U9358 (N_9358,N_8130,N_8577);
or U9359 (N_9359,N_8035,N_8470);
nand U9360 (N_9360,N_8414,N_8648);
or U9361 (N_9361,N_8532,N_8266);
nor U9362 (N_9362,N_8102,N_8423);
nand U9363 (N_9363,N_8905,N_8198);
xor U9364 (N_9364,N_8736,N_8261);
xor U9365 (N_9365,N_8498,N_8738);
xnor U9366 (N_9366,N_8621,N_8754);
nor U9367 (N_9367,N_8219,N_8111);
nor U9368 (N_9368,N_8281,N_8770);
or U9369 (N_9369,N_8056,N_8716);
nor U9370 (N_9370,N_8968,N_8916);
nand U9371 (N_9371,N_8463,N_8711);
xor U9372 (N_9372,N_8950,N_8811);
or U9373 (N_9373,N_8966,N_8389);
nand U9374 (N_9374,N_8299,N_8040);
xnor U9375 (N_9375,N_8893,N_8344);
xnor U9376 (N_9376,N_8775,N_8810);
xnor U9377 (N_9377,N_8523,N_8749);
nand U9378 (N_9378,N_8912,N_8368);
nand U9379 (N_9379,N_8967,N_8069);
or U9380 (N_9380,N_8835,N_8765);
nand U9381 (N_9381,N_8210,N_8884);
nand U9382 (N_9382,N_8774,N_8608);
nand U9383 (N_9383,N_8914,N_8584);
nor U9384 (N_9384,N_8524,N_8067);
or U9385 (N_9385,N_8317,N_8383);
xor U9386 (N_9386,N_8469,N_8006);
or U9387 (N_9387,N_8090,N_8437);
and U9388 (N_9388,N_8582,N_8913);
nand U9389 (N_9389,N_8794,N_8252);
or U9390 (N_9390,N_8752,N_8640);
and U9391 (N_9391,N_8172,N_8812);
or U9392 (N_9392,N_8795,N_8894);
nor U9393 (N_9393,N_8419,N_8049);
and U9394 (N_9394,N_8956,N_8748);
xor U9395 (N_9395,N_8798,N_8824);
xor U9396 (N_9396,N_8019,N_8249);
xor U9397 (N_9397,N_8162,N_8569);
nor U9398 (N_9398,N_8862,N_8695);
or U9399 (N_9399,N_8295,N_8692);
and U9400 (N_9400,N_8520,N_8246);
nor U9401 (N_9401,N_8052,N_8705);
nand U9402 (N_9402,N_8709,N_8593);
or U9403 (N_9403,N_8340,N_8954);
and U9404 (N_9404,N_8886,N_8972);
and U9405 (N_9405,N_8516,N_8289);
xnor U9406 (N_9406,N_8802,N_8464);
xor U9407 (N_9407,N_8314,N_8521);
nor U9408 (N_9408,N_8876,N_8262);
and U9409 (N_9409,N_8020,N_8038);
xor U9410 (N_9410,N_8813,N_8374);
xnor U9411 (N_9411,N_8187,N_8943);
and U9412 (N_9412,N_8674,N_8050);
xor U9413 (N_9413,N_8398,N_8441);
nor U9414 (N_9414,N_8992,N_8567);
nand U9415 (N_9415,N_8206,N_8123);
or U9416 (N_9416,N_8760,N_8482);
xor U9417 (N_9417,N_8937,N_8166);
xnor U9418 (N_9418,N_8767,N_8046);
xnor U9419 (N_9419,N_8510,N_8173);
or U9420 (N_9420,N_8156,N_8641);
xnor U9421 (N_9421,N_8359,N_8468);
nand U9422 (N_9422,N_8336,N_8282);
xor U9423 (N_9423,N_8560,N_8221);
nor U9424 (N_9424,N_8431,N_8686);
and U9425 (N_9425,N_8679,N_8224);
xnor U9426 (N_9426,N_8456,N_8010);
nand U9427 (N_9427,N_8298,N_8693);
nand U9428 (N_9428,N_8550,N_8715);
nor U9429 (N_9429,N_8624,N_8515);
nor U9430 (N_9430,N_8660,N_8728);
nor U9431 (N_9431,N_8303,N_8408);
and U9432 (N_9432,N_8881,N_8091);
nand U9433 (N_9433,N_8999,N_8296);
and U9434 (N_9434,N_8120,N_8013);
nor U9435 (N_9435,N_8350,N_8487);
nor U9436 (N_9436,N_8129,N_8552);
and U9437 (N_9437,N_8346,N_8165);
or U9438 (N_9438,N_8407,N_8676);
and U9439 (N_9439,N_8304,N_8371);
or U9440 (N_9440,N_8191,N_8604);
nand U9441 (N_9441,N_8979,N_8576);
xnor U9442 (N_9442,N_8790,N_8655);
nand U9443 (N_9443,N_8260,N_8095);
nor U9444 (N_9444,N_8060,N_8215);
and U9445 (N_9445,N_8500,N_8772);
nor U9446 (N_9446,N_8935,N_8858);
nor U9447 (N_9447,N_8483,N_8140);
nor U9448 (N_9448,N_8829,N_8209);
nand U9449 (N_9449,N_8332,N_8564);
or U9450 (N_9450,N_8405,N_8929);
xor U9451 (N_9451,N_8882,N_8199);
nor U9452 (N_9452,N_8502,N_8814);
nor U9453 (N_9453,N_8460,N_8154);
and U9454 (N_9454,N_8727,N_8926);
and U9455 (N_9455,N_8789,N_8240);
nor U9456 (N_9456,N_8200,N_8218);
or U9457 (N_9457,N_8182,N_8492);
nand U9458 (N_9458,N_8630,N_8157);
or U9459 (N_9459,N_8275,N_8163);
xnor U9460 (N_9460,N_8453,N_8633);
or U9461 (N_9461,N_8658,N_8661);
or U9462 (N_9462,N_8806,N_8699);
nor U9463 (N_9463,N_8009,N_8807);
or U9464 (N_9464,N_8675,N_8819);
nand U9465 (N_9465,N_8792,N_8941);
and U9466 (N_9466,N_8228,N_8270);
xor U9467 (N_9467,N_8132,N_8958);
and U9468 (N_9468,N_8901,N_8083);
xor U9469 (N_9469,N_8823,N_8677);
nand U9470 (N_9470,N_8874,N_8507);
nand U9471 (N_9471,N_8883,N_8634);
nand U9472 (N_9472,N_8349,N_8074);
and U9473 (N_9473,N_8620,N_8989);
and U9474 (N_9474,N_8513,N_8004);
nand U9475 (N_9475,N_8126,N_8158);
or U9476 (N_9476,N_8891,N_8451);
xor U9477 (N_9477,N_8205,N_8546);
nor U9478 (N_9478,N_8084,N_8135);
and U9479 (N_9479,N_8008,N_8195);
nor U9480 (N_9480,N_8455,N_8347);
or U9481 (N_9481,N_8255,N_8412);
nor U9482 (N_9482,N_8211,N_8986);
nand U9483 (N_9483,N_8787,N_8815);
xor U9484 (N_9484,N_8962,N_8910);
or U9485 (N_9485,N_8394,N_8404);
and U9486 (N_9486,N_8940,N_8808);
or U9487 (N_9487,N_8706,N_8079);
nand U9488 (N_9488,N_8357,N_8353);
and U9489 (N_9489,N_8525,N_8114);
xnor U9490 (N_9490,N_8511,N_8875);
xor U9491 (N_9491,N_8917,N_8656);
xor U9492 (N_9492,N_8105,N_8697);
or U9493 (N_9493,N_8746,N_8458);
or U9494 (N_9494,N_8614,N_8029);
xnor U9495 (N_9495,N_8493,N_8113);
xor U9496 (N_9496,N_8122,N_8991);
nand U9497 (N_9497,N_8854,N_8085);
and U9498 (N_9498,N_8919,N_8816);
and U9499 (N_9499,N_8996,N_8457);
or U9500 (N_9500,N_8730,N_8776);
nor U9501 (N_9501,N_8131,N_8587);
or U9502 (N_9502,N_8175,N_8547);
or U9503 (N_9503,N_8866,N_8839);
nand U9504 (N_9504,N_8874,N_8457);
nor U9505 (N_9505,N_8509,N_8790);
xor U9506 (N_9506,N_8912,N_8875);
xor U9507 (N_9507,N_8316,N_8445);
or U9508 (N_9508,N_8380,N_8989);
and U9509 (N_9509,N_8256,N_8772);
nor U9510 (N_9510,N_8466,N_8277);
nand U9511 (N_9511,N_8529,N_8780);
xnor U9512 (N_9512,N_8475,N_8491);
xnor U9513 (N_9513,N_8354,N_8450);
and U9514 (N_9514,N_8116,N_8942);
and U9515 (N_9515,N_8428,N_8477);
nor U9516 (N_9516,N_8004,N_8005);
and U9517 (N_9517,N_8768,N_8574);
and U9518 (N_9518,N_8914,N_8444);
xor U9519 (N_9519,N_8955,N_8701);
xor U9520 (N_9520,N_8635,N_8115);
and U9521 (N_9521,N_8293,N_8566);
nor U9522 (N_9522,N_8781,N_8332);
xor U9523 (N_9523,N_8155,N_8399);
and U9524 (N_9524,N_8335,N_8341);
or U9525 (N_9525,N_8063,N_8839);
xnor U9526 (N_9526,N_8783,N_8224);
nor U9527 (N_9527,N_8115,N_8624);
nand U9528 (N_9528,N_8529,N_8591);
xor U9529 (N_9529,N_8700,N_8823);
nor U9530 (N_9530,N_8261,N_8748);
xnor U9531 (N_9531,N_8340,N_8125);
xnor U9532 (N_9532,N_8088,N_8850);
nand U9533 (N_9533,N_8214,N_8396);
and U9534 (N_9534,N_8633,N_8767);
or U9535 (N_9535,N_8828,N_8204);
xnor U9536 (N_9536,N_8225,N_8138);
nor U9537 (N_9537,N_8380,N_8621);
nor U9538 (N_9538,N_8042,N_8769);
nor U9539 (N_9539,N_8954,N_8009);
nor U9540 (N_9540,N_8629,N_8642);
nand U9541 (N_9541,N_8825,N_8578);
or U9542 (N_9542,N_8978,N_8521);
and U9543 (N_9543,N_8767,N_8788);
and U9544 (N_9544,N_8636,N_8385);
and U9545 (N_9545,N_8675,N_8312);
xor U9546 (N_9546,N_8326,N_8746);
and U9547 (N_9547,N_8954,N_8310);
and U9548 (N_9548,N_8272,N_8246);
xnor U9549 (N_9549,N_8319,N_8631);
or U9550 (N_9550,N_8610,N_8787);
nand U9551 (N_9551,N_8356,N_8328);
or U9552 (N_9552,N_8947,N_8354);
or U9553 (N_9553,N_8905,N_8350);
and U9554 (N_9554,N_8040,N_8130);
nand U9555 (N_9555,N_8617,N_8941);
or U9556 (N_9556,N_8789,N_8885);
xor U9557 (N_9557,N_8301,N_8461);
xnor U9558 (N_9558,N_8329,N_8684);
nand U9559 (N_9559,N_8077,N_8149);
xor U9560 (N_9560,N_8904,N_8958);
and U9561 (N_9561,N_8184,N_8156);
xor U9562 (N_9562,N_8720,N_8895);
nor U9563 (N_9563,N_8689,N_8839);
or U9564 (N_9564,N_8830,N_8137);
xnor U9565 (N_9565,N_8040,N_8906);
or U9566 (N_9566,N_8265,N_8522);
nand U9567 (N_9567,N_8789,N_8591);
or U9568 (N_9568,N_8511,N_8636);
and U9569 (N_9569,N_8862,N_8768);
xor U9570 (N_9570,N_8703,N_8011);
and U9571 (N_9571,N_8225,N_8038);
or U9572 (N_9572,N_8670,N_8238);
xor U9573 (N_9573,N_8032,N_8047);
nor U9574 (N_9574,N_8241,N_8504);
nor U9575 (N_9575,N_8950,N_8327);
and U9576 (N_9576,N_8693,N_8415);
nand U9577 (N_9577,N_8728,N_8258);
nor U9578 (N_9578,N_8380,N_8865);
and U9579 (N_9579,N_8870,N_8474);
nand U9580 (N_9580,N_8328,N_8355);
xnor U9581 (N_9581,N_8958,N_8807);
xor U9582 (N_9582,N_8729,N_8970);
and U9583 (N_9583,N_8094,N_8586);
or U9584 (N_9584,N_8032,N_8584);
nor U9585 (N_9585,N_8134,N_8099);
or U9586 (N_9586,N_8760,N_8006);
nand U9587 (N_9587,N_8265,N_8978);
nor U9588 (N_9588,N_8314,N_8828);
nand U9589 (N_9589,N_8281,N_8429);
xor U9590 (N_9590,N_8431,N_8690);
nor U9591 (N_9591,N_8200,N_8792);
and U9592 (N_9592,N_8139,N_8562);
nor U9593 (N_9593,N_8121,N_8211);
xnor U9594 (N_9594,N_8031,N_8987);
or U9595 (N_9595,N_8177,N_8638);
nand U9596 (N_9596,N_8467,N_8945);
and U9597 (N_9597,N_8080,N_8483);
nand U9598 (N_9598,N_8796,N_8121);
or U9599 (N_9599,N_8891,N_8188);
xnor U9600 (N_9600,N_8080,N_8519);
or U9601 (N_9601,N_8105,N_8836);
nor U9602 (N_9602,N_8449,N_8603);
and U9603 (N_9603,N_8086,N_8227);
xor U9604 (N_9604,N_8642,N_8344);
or U9605 (N_9605,N_8870,N_8494);
nand U9606 (N_9606,N_8504,N_8020);
and U9607 (N_9607,N_8472,N_8727);
nor U9608 (N_9608,N_8477,N_8026);
and U9609 (N_9609,N_8806,N_8346);
nand U9610 (N_9610,N_8054,N_8010);
nor U9611 (N_9611,N_8688,N_8983);
nor U9612 (N_9612,N_8498,N_8462);
xor U9613 (N_9613,N_8218,N_8881);
or U9614 (N_9614,N_8942,N_8472);
xor U9615 (N_9615,N_8334,N_8209);
nand U9616 (N_9616,N_8772,N_8348);
xnor U9617 (N_9617,N_8361,N_8876);
nand U9618 (N_9618,N_8685,N_8676);
and U9619 (N_9619,N_8474,N_8735);
and U9620 (N_9620,N_8708,N_8882);
or U9621 (N_9621,N_8839,N_8582);
and U9622 (N_9622,N_8095,N_8979);
or U9623 (N_9623,N_8627,N_8316);
xnor U9624 (N_9624,N_8200,N_8467);
and U9625 (N_9625,N_8411,N_8519);
nor U9626 (N_9626,N_8608,N_8266);
nand U9627 (N_9627,N_8846,N_8332);
nand U9628 (N_9628,N_8240,N_8916);
and U9629 (N_9629,N_8275,N_8806);
xor U9630 (N_9630,N_8737,N_8544);
nor U9631 (N_9631,N_8584,N_8907);
or U9632 (N_9632,N_8314,N_8871);
nor U9633 (N_9633,N_8425,N_8579);
xnor U9634 (N_9634,N_8042,N_8104);
nor U9635 (N_9635,N_8188,N_8260);
nand U9636 (N_9636,N_8920,N_8903);
xor U9637 (N_9637,N_8229,N_8192);
and U9638 (N_9638,N_8038,N_8715);
nand U9639 (N_9639,N_8987,N_8237);
and U9640 (N_9640,N_8795,N_8857);
or U9641 (N_9641,N_8793,N_8650);
or U9642 (N_9642,N_8643,N_8664);
xnor U9643 (N_9643,N_8847,N_8597);
or U9644 (N_9644,N_8626,N_8996);
nand U9645 (N_9645,N_8235,N_8744);
nand U9646 (N_9646,N_8027,N_8285);
and U9647 (N_9647,N_8163,N_8917);
or U9648 (N_9648,N_8476,N_8794);
xnor U9649 (N_9649,N_8614,N_8542);
or U9650 (N_9650,N_8652,N_8081);
nand U9651 (N_9651,N_8268,N_8640);
and U9652 (N_9652,N_8671,N_8975);
xor U9653 (N_9653,N_8488,N_8536);
and U9654 (N_9654,N_8485,N_8354);
or U9655 (N_9655,N_8620,N_8808);
or U9656 (N_9656,N_8676,N_8049);
nor U9657 (N_9657,N_8988,N_8863);
or U9658 (N_9658,N_8135,N_8654);
or U9659 (N_9659,N_8309,N_8315);
nor U9660 (N_9660,N_8111,N_8749);
nand U9661 (N_9661,N_8559,N_8461);
and U9662 (N_9662,N_8790,N_8505);
or U9663 (N_9663,N_8906,N_8914);
xor U9664 (N_9664,N_8526,N_8433);
xor U9665 (N_9665,N_8965,N_8903);
or U9666 (N_9666,N_8683,N_8625);
nor U9667 (N_9667,N_8372,N_8198);
and U9668 (N_9668,N_8982,N_8878);
nor U9669 (N_9669,N_8644,N_8935);
nand U9670 (N_9670,N_8094,N_8795);
and U9671 (N_9671,N_8628,N_8207);
and U9672 (N_9672,N_8142,N_8805);
xnor U9673 (N_9673,N_8935,N_8992);
xnor U9674 (N_9674,N_8776,N_8520);
nand U9675 (N_9675,N_8104,N_8843);
nand U9676 (N_9676,N_8005,N_8755);
xnor U9677 (N_9677,N_8456,N_8105);
and U9678 (N_9678,N_8514,N_8295);
xor U9679 (N_9679,N_8407,N_8691);
nor U9680 (N_9680,N_8416,N_8603);
xor U9681 (N_9681,N_8458,N_8644);
nor U9682 (N_9682,N_8652,N_8433);
and U9683 (N_9683,N_8550,N_8102);
or U9684 (N_9684,N_8596,N_8247);
nand U9685 (N_9685,N_8736,N_8262);
nand U9686 (N_9686,N_8729,N_8163);
and U9687 (N_9687,N_8016,N_8895);
xor U9688 (N_9688,N_8220,N_8924);
nor U9689 (N_9689,N_8124,N_8149);
xor U9690 (N_9690,N_8262,N_8360);
nor U9691 (N_9691,N_8781,N_8420);
and U9692 (N_9692,N_8781,N_8061);
and U9693 (N_9693,N_8990,N_8057);
xor U9694 (N_9694,N_8400,N_8938);
nand U9695 (N_9695,N_8338,N_8856);
nand U9696 (N_9696,N_8751,N_8951);
and U9697 (N_9697,N_8100,N_8476);
nand U9698 (N_9698,N_8648,N_8977);
xor U9699 (N_9699,N_8378,N_8786);
xnor U9700 (N_9700,N_8450,N_8930);
nor U9701 (N_9701,N_8295,N_8536);
xnor U9702 (N_9702,N_8788,N_8425);
xor U9703 (N_9703,N_8492,N_8241);
or U9704 (N_9704,N_8325,N_8424);
xnor U9705 (N_9705,N_8517,N_8652);
or U9706 (N_9706,N_8433,N_8715);
or U9707 (N_9707,N_8297,N_8392);
nor U9708 (N_9708,N_8780,N_8960);
nor U9709 (N_9709,N_8594,N_8443);
or U9710 (N_9710,N_8892,N_8315);
xor U9711 (N_9711,N_8960,N_8143);
nand U9712 (N_9712,N_8600,N_8792);
and U9713 (N_9713,N_8797,N_8375);
nand U9714 (N_9714,N_8806,N_8573);
or U9715 (N_9715,N_8203,N_8314);
xnor U9716 (N_9716,N_8717,N_8053);
nor U9717 (N_9717,N_8541,N_8174);
and U9718 (N_9718,N_8932,N_8686);
xnor U9719 (N_9719,N_8690,N_8348);
nor U9720 (N_9720,N_8332,N_8760);
and U9721 (N_9721,N_8609,N_8720);
nor U9722 (N_9722,N_8450,N_8796);
or U9723 (N_9723,N_8838,N_8580);
and U9724 (N_9724,N_8143,N_8090);
nand U9725 (N_9725,N_8807,N_8641);
xor U9726 (N_9726,N_8062,N_8717);
and U9727 (N_9727,N_8224,N_8995);
nand U9728 (N_9728,N_8873,N_8565);
nand U9729 (N_9729,N_8737,N_8188);
or U9730 (N_9730,N_8404,N_8539);
nand U9731 (N_9731,N_8207,N_8502);
nor U9732 (N_9732,N_8477,N_8659);
or U9733 (N_9733,N_8167,N_8871);
or U9734 (N_9734,N_8406,N_8373);
nor U9735 (N_9735,N_8832,N_8106);
or U9736 (N_9736,N_8287,N_8257);
xor U9737 (N_9737,N_8407,N_8842);
nor U9738 (N_9738,N_8575,N_8219);
nor U9739 (N_9739,N_8465,N_8261);
or U9740 (N_9740,N_8179,N_8323);
nor U9741 (N_9741,N_8104,N_8037);
and U9742 (N_9742,N_8517,N_8996);
or U9743 (N_9743,N_8662,N_8325);
nand U9744 (N_9744,N_8544,N_8201);
xnor U9745 (N_9745,N_8838,N_8853);
or U9746 (N_9746,N_8462,N_8014);
and U9747 (N_9747,N_8754,N_8162);
xnor U9748 (N_9748,N_8155,N_8099);
or U9749 (N_9749,N_8681,N_8809);
xor U9750 (N_9750,N_8252,N_8448);
or U9751 (N_9751,N_8539,N_8345);
nand U9752 (N_9752,N_8982,N_8767);
nand U9753 (N_9753,N_8457,N_8144);
or U9754 (N_9754,N_8931,N_8920);
or U9755 (N_9755,N_8683,N_8996);
or U9756 (N_9756,N_8822,N_8149);
nor U9757 (N_9757,N_8938,N_8412);
nor U9758 (N_9758,N_8189,N_8313);
and U9759 (N_9759,N_8484,N_8909);
xnor U9760 (N_9760,N_8060,N_8811);
and U9761 (N_9761,N_8482,N_8566);
xor U9762 (N_9762,N_8418,N_8299);
nand U9763 (N_9763,N_8030,N_8539);
nor U9764 (N_9764,N_8676,N_8141);
xor U9765 (N_9765,N_8463,N_8200);
or U9766 (N_9766,N_8048,N_8463);
or U9767 (N_9767,N_8552,N_8562);
or U9768 (N_9768,N_8533,N_8882);
xor U9769 (N_9769,N_8619,N_8112);
nor U9770 (N_9770,N_8513,N_8955);
and U9771 (N_9771,N_8068,N_8342);
and U9772 (N_9772,N_8794,N_8341);
nand U9773 (N_9773,N_8180,N_8756);
nor U9774 (N_9774,N_8802,N_8623);
and U9775 (N_9775,N_8464,N_8969);
xor U9776 (N_9776,N_8647,N_8217);
xnor U9777 (N_9777,N_8503,N_8137);
or U9778 (N_9778,N_8247,N_8896);
xnor U9779 (N_9779,N_8257,N_8096);
nand U9780 (N_9780,N_8637,N_8228);
xnor U9781 (N_9781,N_8242,N_8598);
nand U9782 (N_9782,N_8949,N_8797);
nand U9783 (N_9783,N_8342,N_8799);
or U9784 (N_9784,N_8501,N_8204);
nand U9785 (N_9785,N_8064,N_8256);
or U9786 (N_9786,N_8249,N_8796);
or U9787 (N_9787,N_8349,N_8672);
xor U9788 (N_9788,N_8539,N_8360);
or U9789 (N_9789,N_8746,N_8138);
xnor U9790 (N_9790,N_8556,N_8366);
xor U9791 (N_9791,N_8737,N_8444);
and U9792 (N_9792,N_8152,N_8547);
or U9793 (N_9793,N_8666,N_8226);
or U9794 (N_9794,N_8825,N_8259);
and U9795 (N_9795,N_8539,N_8990);
or U9796 (N_9796,N_8300,N_8335);
xnor U9797 (N_9797,N_8180,N_8126);
nand U9798 (N_9798,N_8268,N_8846);
nor U9799 (N_9799,N_8963,N_8613);
nand U9800 (N_9800,N_8845,N_8688);
or U9801 (N_9801,N_8022,N_8141);
nand U9802 (N_9802,N_8046,N_8173);
or U9803 (N_9803,N_8875,N_8046);
and U9804 (N_9804,N_8393,N_8631);
xor U9805 (N_9805,N_8518,N_8327);
and U9806 (N_9806,N_8470,N_8736);
and U9807 (N_9807,N_8127,N_8521);
and U9808 (N_9808,N_8386,N_8707);
or U9809 (N_9809,N_8599,N_8544);
xor U9810 (N_9810,N_8973,N_8671);
xor U9811 (N_9811,N_8107,N_8817);
or U9812 (N_9812,N_8782,N_8660);
nand U9813 (N_9813,N_8182,N_8615);
nand U9814 (N_9814,N_8868,N_8684);
and U9815 (N_9815,N_8418,N_8625);
and U9816 (N_9816,N_8553,N_8601);
xor U9817 (N_9817,N_8409,N_8912);
or U9818 (N_9818,N_8829,N_8226);
xor U9819 (N_9819,N_8864,N_8453);
nor U9820 (N_9820,N_8162,N_8035);
xor U9821 (N_9821,N_8314,N_8393);
or U9822 (N_9822,N_8487,N_8327);
xor U9823 (N_9823,N_8113,N_8409);
and U9824 (N_9824,N_8143,N_8464);
nand U9825 (N_9825,N_8358,N_8478);
nor U9826 (N_9826,N_8818,N_8849);
and U9827 (N_9827,N_8902,N_8334);
or U9828 (N_9828,N_8024,N_8666);
and U9829 (N_9829,N_8299,N_8330);
xnor U9830 (N_9830,N_8889,N_8368);
and U9831 (N_9831,N_8423,N_8879);
xor U9832 (N_9832,N_8183,N_8272);
and U9833 (N_9833,N_8953,N_8053);
and U9834 (N_9834,N_8912,N_8622);
xnor U9835 (N_9835,N_8205,N_8914);
nand U9836 (N_9836,N_8260,N_8110);
or U9837 (N_9837,N_8413,N_8784);
or U9838 (N_9838,N_8415,N_8815);
or U9839 (N_9839,N_8205,N_8600);
nand U9840 (N_9840,N_8096,N_8031);
nand U9841 (N_9841,N_8071,N_8456);
nor U9842 (N_9842,N_8435,N_8397);
or U9843 (N_9843,N_8245,N_8486);
and U9844 (N_9844,N_8108,N_8910);
xnor U9845 (N_9845,N_8846,N_8748);
and U9846 (N_9846,N_8296,N_8246);
nand U9847 (N_9847,N_8173,N_8770);
nor U9848 (N_9848,N_8522,N_8220);
nand U9849 (N_9849,N_8324,N_8299);
xor U9850 (N_9850,N_8423,N_8577);
or U9851 (N_9851,N_8829,N_8688);
or U9852 (N_9852,N_8628,N_8534);
and U9853 (N_9853,N_8918,N_8830);
nand U9854 (N_9854,N_8101,N_8446);
xor U9855 (N_9855,N_8912,N_8389);
xor U9856 (N_9856,N_8274,N_8477);
or U9857 (N_9857,N_8360,N_8920);
nor U9858 (N_9858,N_8828,N_8370);
or U9859 (N_9859,N_8637,N_8188);
nor U9860 (N_9860,N_8599,N_8369);
or U9861 (N_9861,N_8259,N_8958);
xnor U9862 (N_9862,N_8260,N_8755);
nor U9863 (N_9863,N_8553,N_8339);
nand U9864 (N_9864,N_8498,N_8550);
nand U9865 (N_9865,N_8253,N_8563);
nor U9866 (N_9866,N_8113,N_8689);
or U9867 (N_9867,N_8233,N_8845);
or U9868 (N_9868,N_8515,N_8834);
or U9869 (N_9869,N_8830,N_8193);
and U9870 (N_9870,N_8227,N_8237);
and U9871 (N_9871,N_8805,N_8597);
nor U9872 (N_9872,N_8053,N_8710);
or U9873 (N_9873,N_8976,N_8309);
and U9874 (N_9874,N_8567,N_8755);
nand U9875 (N_9875,N_8329,N_8384);
nand U9876 (N_9876,N_8176,N_8642);
and U9877 (N_9877,N_8780,N_8212);
or U9878 (N_9878,N_8001,N_8093);
nand U9879 (N_9879,N_8300,N_8378);
nor U9880 (N_9880,N_8181,N_8387);
xor U9881 (N_9881,N_8950,N_8965);
xor U9882 (N_9882,N_8730,N_8941);
and U9883 (N_9883,N_8303,N_8372);
nor U9884 (N_9884,N_8751,N_8527);
or U9885 (N_9885,N_8145,N_8660);
and U9886 (N_9886,N_8231,N_8846);
nor U9887 (N_9887,N_8925,N_8455);
and U9888 (N_9888,N_8940,N_8225);
nor U9889 (N_9889,N_8345,N_8743);
nand U9890 (N_9890,N_8971,N_8201);
or U9891 (N_9891,N_8357,N_8010);
xor U9892 (N_9892,N_8324,N_8651);
nand U9893 (N_9893,N_8576,N_8889);
and U9894 (N_9894,N_8748,N_8943);
or U9895 (N_9895,N_8024,N_8671);
or U9896 (N_9896,N_8529,N_8199);
nand U9897 (N_9897,N_8124,N_8947);
xor U9898 (N_9898,N_8721,N_8206);
or U9899 (N_9899,N_8697,N_8001);
nand U9900 (N_9900,N_8563,N_8933);
and U9901 (N_9901,N_8902,N_8964);
xor U9902 (N_9902,N_8822,N_8510);
xor U9903 (N_9903,N_8135,N_8288);
and U9904 (N_9904,N_8210,N_8865);
xor U9905 (N_9905,N_8522,N_8332);
and U9906 (N_9906,N_8210,N_8499);
or U9907 (N_9907,N_8423,N_8538);
nor U9908 (N_9908,N_8477,N_8444);
nor U9909 (N_9909,N_8257,N_8233);
nand U9910 (N_9910,N_8985,N_8224);
or U9911 (N_9911,N_8446,N_8788);
nand U9912 (N_9912,N_8856,N_8381);
nand U9913 (N_9913,N_8577,N_8535);
xnor U9914 (N_9914,N_8354,N_8949);
nor U9915 (N_9915,N_8005,N_8821);
or U9916 (N_9916,N_8593,N_8325);
nor U9917 (N_9917,N_8006,N_8671);
and U9918 (N_9918,N_8332,N_8227);
xnor U9919 (N_9919,N_8260,N_8359);
nor U9920 (N_9920,N_8751,N_8183);
or U9921 (N_9921,N_8777,N_8348);
or U9922 (N_9922,N_8786,N_8405);
nor U9923 (N_9923,N_8605,N_8125);
xnor U9924 (N_9924,N_8926,N_8849);
nor U9925 (N_9925,N_8624,N_8066);
xor U9926 (N_9926,N_8201,N_8922);
nand U9927 (N_9927,N_8533,N_8568);
or U9928 (N_9928,N_8746,N_8401);
or U9929 (N_9929,N_8463,N_8353);
or U9930 (N_9930,N_8405,N_8915);
xor U9931 (N_9931,N_8459,N_8241);
and U9932 (N_9932,N_8022,N_8090);
nor U9933 (N_9933,N_8965,N_8658);
xnor U9934 (N_9934,N_8705,N_8079);
xor U9935 (N_9935,N_8166,N_8085);
nand U9936 (N_9936,N_8084,N_8813);
xnor U9937 (N_9937,N_8176,N_8685);
and U9938 (N_9938,N_8975,N_8530);
xnor U9939 (N_9939,N_8297,N_8407);
or U9940 (N_9940,N_8671,N_8791);
nand U9941 (N_9941,N_8726,N_8852);
xnor U9942 (N_9942,N_8119,N_8677);
nand U9943 (N_9943,N_8284,N_8977);
and U9944 (N_9944,N_8283,N_8489);
nor U9945 (N_9945,N_8763,N_8746);
and U9946 (N_9946,N_8616,N_8726);
nor U9947 (N_9947,N_8782,N_8767);
nand U9948 (N_9948,N_8002,N_8259);
nand U9949 (N_9949,N_8167,N_8744);
and U9950 (N_9950,N_8012,N_8967);
and U9951 (N_9951,N_8599,N_8183);
xnor U9952 (N_9952,N_8911,N_8963);
or U9953 (N_9953,N_8373,N_8357);
and U9954 (N_9954,N_8212,N_8681);
nor U9955 (N_9955,N_8824,N_8953);
or U9956 (N_9956,N_8172,N_8589);
xnor U9957 (N_9957,N_8301,N_8133);
nor U9958 (N_9958,N_8595,N_8102);
nand U9959 (N_9959,N_8486,N_8231);
or U9960 (N_9960,N_8841,N_8621);
xor U9961 (N_9961,N_8321,N_8193);
xnor U9962 (N_9962,N_8486,N_8652);
nor U9963 (N_9963,N_8180,N_8773);
nor U9964 (N_9964,N_8808,N_8003);
xor U9965 (N_9965,N_8522,N_8667);
nor U9966 (N_9966,N_8590,N_8717);
nor U9967 (N_9967,N_8448,N_8161);
and U9968 (N_9968,N_8677,N_8645);
nor U9969 (N_9969,N_8083,N_8210);
nand U9970 (N_9970,N_8177,N_8794);
and U9971 (N_9971,N_8749,N_8341);
and U9972 (N_9972,N_8945,N_8854);
nor U9973 (N_9973,N_8410,N_8074);
nand U9974 (N_9974,N_8795,N_8374);
or U9975 (N_9975,N_8972,N_8237);
or U9976 (N_9976,N_8722,N_8433);
and U9977 (N_9977,N_8191,N_8803);
or U9978 (N_9978,N_8102,N_8402);
nand U9979 (N_9979,N_8008,N_8039);
nor U9980 (N_9980,N_8382,N_8437);
nor U9981 (N_9981,N_8568,N_8933);
xnor U9982 (N_9982,N_8197,N_8261);
nor U9983 (N_9983,N_8233,N_8301);
or U9984 (N_9984,N_8100,N_8391);
xnor U9985 (N_9985,N_8626,N_8248);
or U9986 (N_9986,N_8173,N_8817);
or U9987 (N_9987,N_8153,N_8041);
and U9988 (N_9988,N_8399,N_8732);
and U9989 (N_9989,N_8283,N_8713);
or U9990 (N_9990,N_8647,N_8335);
or U9991 (N_9991,N_8658,N_8899);
or U9992 (N_9992,N_8033,N_8602);
and U9993 (N_9993,N_8646,N_8176);
nor U9994 (N_9994,N_8378,N_8194);
or U9995 (N_9995,N_8770,N_8032);
or U9996 (N_9996,N_8289,N_8707);
or U9997 (N_9997,N_8621,N_8468);
nor U9998 (N_9998,N_8866,N_8576);
and U9999 (N_9999,N_8321,N_8580);
or UO_0 (O_0,N_9401,N_9449);
and UO_1 (O_1,N_9759,N_9425);
nor UO_2 (O_2,N_9155,N_9341);
nor UO_3 (O_3,N_9793,N_9665);
or UO_4 (O_4,N_9188,N_9097);
nand UO_5 (O_5,N_9932,N_9220);
xor UO_6 (O_6,N_9357,N_9326);
or UO_7 (O_7,N_9257,N_9271);
or UO_8 (O_8,N_9890,N_9804);
nor UO_9 (O_9,N_9572,N_9854);
and UO_10 (O_10,N_9429,N_9468);
nand UO_11 (O_11,N_9568,N_9356);
nor UO_12 (O_12,N_9632,N_9438);
or UO_13 (O_13,N_9725,N_9048);
or UO_14 (O_14,N_9721,N_9762);
xor UO_15 (O_15,N_9749,N_9594);
nand UO_16 (O_16,N_9872,N_9910);
and UO_17 (O_17,N_9314,N_9413);
xor UO_18 (O_18,N_9473,N_9720);
nor UO_19 (O_19,N_9618,N_9622);
xnor UO_20 (O_20,N_9095,N_9247);
xnor UO_21 (O_21,N_9833,N_9072);
xor UO_22 (O_22,N_9293,N_9988);
xnor UO_23 (O_23,N_9683,N_9682);
or UO_24 (O_24,N_9953,N_9621);
nand UO_25 (O_25,N_9135,N_9713);
nand UO_26 (O_26,N_9645,N_9339);
and UO_27 (O_27,N_9096,N_9007);
and UO_28 (O_28,N_9639,N_9724);
or UO_29 (O_29,N_9963,N_9969);
xnor UO_30 (O_30,N_9190,N_9411);
nor UO_31 (O_31,N_9422,N_9646);
nand UO_32 (O_32,N_9965,N_9525);
and UO_33 (O_33,N_9466,N_9433);
nor UO_34 (O_34,N_9921,N_9849);
nor UO_35 (O_35,N_9183,N_9671);
nor UO_36 (O_36,N_9458,N_9926);
or UO_37 (O_37,N_9016,N_9276);
or UO_38 (O_38,N_9968,N_9924);
nor UO_39 (O_39,N_9566,N_9669);
nand UO_40 (O_40,N_9308,N_9384);
xnor UO_41 (O_41,N_9363,N_9132);
xnor UO_42 (O_42,N_9636,N_9415);
and UO_43 (O_43,N_9011,N_9049);
and UO_44 (O_44,N_9191,N_9288);
nor UO_45 (O_45,N_9003,N_9487);
and UO_46 (O_46,N_9248,N_9131);
xnor UO_47 (O_47,N_9533,N_9589);
nand UO_48 (O_48,N_9094,N_9941);
and UO_49 (O_49,N_9014,N_9792);
and UO_50 (O_50,N_9586,N_9147);
and UO_51 (O_51,N_9838,N_9530);
or UO_52 (O_52,N_9554,N_9754);
and UO_53 (O_53,N_9571,N_9588);
xnor UO_54 (O_54,N_9635,N_9855);
nand UO_55 (O_55,N_9696,N_9630);
xnor UO_56 (O_56,N_9477,N_9939);
nand UO_57 (O_57,N_9858,N_9633);
or UO_58 (O_58,N_9758,N_9611);
xnor UO_59 (O_59,N_9087,N_9715);
xor UO_60 (O_60,N_9351,N_9602);
nand UO_61 (O_61,N_9175,N_9518);
nor UO_62 (O_62,N_9802,N_9840);
or UO_63 (O_63,N_9627,N_9428);
xor UO_64 (O_64,N_9142,N_9712);
nand UO_65 (O_65,N_9548,N_9836);
and UO_66 (O_66,N_9167,N_9181);
and UO_67 (O_67,N_9071,N_9416);
nand UO_68 (O_68,N_9763,N_9666);
or UO_69 (O_69,N_9361,N_9327);
or UO_70 (O_70,N_9911,N_9483);
or UO_71 (O_71,N_9563,N_9672);
or UO_72 (O_72,N_9524,N_9818);
or UO_73 (O_73,N_9610,N_9080);
and UO_74 (O_74,N_9005,N_9516);
nor UO_75 (O_75,N_9212,N_9006);
xnor UO_76 (O_76,N_9798,N_9209);
and UO_77 (O_77,N_9536,N_9151);
nand UO_78 (O_78,N_9812,N_9866);
and UO_79 (O_79,N_9277,N_9170);
and UO_80 (O_80,N_9026,N_9734);
nand UO_81 (O_81,N_9919,N_9527);
or UO_82 (O_82,N_9105,N_9883);
and UO_83 (O_83,N_9791,N_9644);
or UO_84 (O_84,N_9453,N_9219);
and UO_85 (O_85,N_9115,N_9534);
nor UO_86 (O_86,N_9591,N_9947);
nor UO_87 (O_87,N_9670,N_9502);
and UO_88 (O_88,N_9821,N_9021);
nor UO_89 (O_89,N_9598,N_9979);
or UO_90 (O_90,N_9182,N_9073);
xnor UO_91 (O_91,N_9814,N_9200);
nand UO_92 (O_92,N_9218,N_9723);
nor UO_93 (O_93,N_9169,N_9984);
xnor UO_94 (O_94,N_9454,N_9730);
xnor UO_95 (O_95,N_9058,N_9000);
and UO_96 (O_96,N_9399,N_9322);
and UO_97 (O_97,N_9587,N_9558);
nand UO_98 (O_98,N_9999,N_9279);
or UO_99 (O_99,N_9832,N_9189);
nor UO_100 (O_100,N_9726,N_9788);
nor UO_101 (O_101,N_9410,N_9579);
xnor UO_102 (O_102,N_9470,N_9262);
nand UO_103 (O_103,N_9737,N_9590);
or UO_104 (O_104,N_9060,N_9992);
nand UO_105 (O_105,N_9380,N_9834);
or UO_106 (O_106,N_9464,N_9997);
nor UO_107 (O_107,N_9280,N_9857);
nor UO_108 (O_108,N_9925,N_9124);
and UO_109 (O_109,N_9418,N_9180);
and UO_110 (O_110,N_9728,N_9013);
and UO_111 (O_111,N_9831,N_9837);
xnor UO_112 (O_112,N_9333,N_9229);
nand UO_113 (O_113,N_9227,N_9478);
and UO_114 (O_114,N_9557,N_9576);
or UO_115 (O_115,N_9597,N_9330);
nand UO_116 (O_116,N_9122,N_9120);
nor UO_117 (O_117,N_9196,N_9620);
or UO_118 (O_118,N_9030,N_9523);
xor UO_119 (O_119,N_9117,N_9868);
xor UO_120 (O_120,N_9938,N_9686);
and UO_121 (O_121,N_9017,N_9743);
or UO_122 (O_122,N_9661,N_9052);
nand UO_123 (O_123,N_9448,N_9900);
xor UO_124 (O_124,N_9972,N_9643);
and UO_125 (O_125,N_9908,N_9998);
or UO_126 (O_126,N_9395,N_9313);
xor UO_127 (O_127,N_9540,N_9581);
nor UO_128 (O_128,N_9511,N_9535);
xor UO_129 (O_129,N_9373,N_9368);
nand UO_130 (O_130,N_9830,N_9547);
or UO_131 (O_131,N_9442,N_9358);
nor UO_132 (O_132,N_9034,N_9657);
nor UO_133 (O_133,N_9647,N_9677);
nand UO_134 (O_134,N_9332,N_9844);
xnor UO_135 (O_135,N_9929,N_9741);
nand UO_136 (O_136,N_9393,N_9652);
or UO_137 (O_137,N_9264,N_9346);
nand UO_138 (O_138,N_9894,N_9617);
and UO_139 (O_139,N_9898,N_9430);
nor UO_140 (O_140,N_9867,N_9778);
xor UO_141 (O_141,N_9978,N_9889);
nor UO_142 (O_142,N_9084,N_9306);
or UO_143 (O_143,N_9660,N_9305);
or UO_144 (O_144,N_9826,N_9482);
nand UO_145 (O_145,N_9119,N_9417);
nand UO_146 (O_146,N_9396,N_9400);
xor UO_147 (O_147,N_9185,N_9782);
xnor UO_148 (O_148,N_9786,N_9769);
nand UO_149 (O_149,N_9971,N_9138);
nand UO_150 (O_150,N_9957,N_9905);
or UO_151 (O_151,N_9261,N_9027);
nor UO_152 (O_152,N_9824,N_9718);
and UO_153 (O_153,N_9962,N_9936);
and UO_154 (O_154,N_9675,N_9233);
nand UO_155 (O_155,N_9150,N_9378);
and UO_156 (O_156,N_9970,N_9560);
and UO_157 (O_157,N_9076,N_9452);
xor UO_158 (O_158,N_9771,N_9184);
nand UO_159 (O_159,N_9714,N_9435);
nand UO_160 (O_160,N_9192,N_9773);
xnor UO_161 (O_161,N_9809,N_9934);
and UO_162 (O_162,N_9063,N_9269);
and UO_163 (O_163,N_9053,N_9045);
nand UO_164 (O_164,N_9893,N_9110);
nand UO_165 (O_165,N_9044,N_9484);
xor UO_166 (O_166,N_9275,N_9684);
nor UO_167 (O_167,N_9056,N_9302);
nand UO_168 (O_168,N_9623,N_9210);
or UO_169 (O_169,N_9583,N_9592);
nor UO_170 (O_170,N_9995,N_9656);
xnor UO_171 (O_171,N_9197,N_9937);
nor UO_172 (O_172,N_9091,N_9785);
nand UO_173 (O_173,N_9272,N_9658);
nand UO_174 (O_174,N_9318,N_9492);
and UO_175 (O_175,N_9436,N_9852);
nor UO_176 (O_176,N_9223,N_9009);
or UO_177 (O_177,N_9245,N_9377);
and UO_178 (O_178,N_9334,N_9845);
nand UO_179 (O_179,N_9099,N_9555);
nor UO_180 (O_180,N_9043,N_9456);
nor UO_181 (O_181,N_9967,N_9575);
xnor UO_182 (O_182,N_9510,N_9878);
and UO_183 (O_183,N_9781,N_9237);
nand UO_184 (O_184,N_9580,N_9806);
xnor UO_185 (O_185,N_9899,N_9813);
xor UO_186 (O_186,N_9311,N_9895);
and UO_187 (O_187,N_9986,N_9480);
nor UO_188 (O_188,N_9427,N_9901);
xnor UO_189 (O_189,N_9663,N_9881);
and UO_190 (O_190,N_9001,N_9486);
xnor UO_191 (O_191,N_9465,N_9613);
or UO_192 (O_192,N_9940,N_9446);
and UO_193 (O_193,N_9153,N_9605);
nor UO_194 (O_194,N_9641,N_9154);
xnor UO_195 (O_195,N_9991,N_9186);
xnor UO_196 (O_196,N_9217,N_9710);
xnor UO_197 (O_197,N_9455,N_9985);
and UO_198 (O_198,N_9260,N_9816);
or UO_199 (O_199,N_9002,N_9199);
and UO_200 (O_200,N_9420,N_9692);
nand UO_201 (O_201,N_9942,N_9137);
or UO_202 (O_202,N_9093,N_9234);
and UO_203 (O_203,N_9437,N_9927);
and UO_204 (O_204,N_9216,N_9390);
xnor UO_205 (O_205,N_9061,N_9081);
or UO_206 (O_206,N_9325,N_9631);
nand UO_207 (O_207,N_9178,N_9561);
xor UO_208 (O_208,N_9461,N_9297);
and UO_209 (O_209,N_9931,N_9202);
and UO_210 (O_210,N_9161,N_9336);
or UO_211 (O_211,N_9177,N_9596);
or UO_212 (O_212,N_9372,N_9582);
nand UO_213 (O_213,N_9604,N_9015);
and UO_214 (O_214,N_9228,N_9441);
or UO_215 (O_215,N_9564,N_9873);
nand UO_216 (O_216,N_9168,N_9366);
or UO_217 (O_217,N_9176,N_9955);
and UO_218 (O_218,N_9208,N_9528);
or UO_219 (O_219,N_9655,N_9689);
xor UO_220 (O_220,N_9966,N_9603);
nor UO_221 (O_221,N_9023,N_9263);
or UO_222 (O_222,N_9127,N_9499);
or UO_223 (O_223,N_9139,N_9585);
and UO_224 (O_224,N_9827,N_9092);
or UO_225 (O_225,N_9029,N_9829);
and UO_226 (O_226,N_9164,N_9650);
and UO_227 (O_227,N_9757,N_9082);
and UO_228 (O_228,N_9907,N_9012);
xor UO_229 (O_229,N_9795,N_9805);
nor UO_230 (O_230,N_9847,N_9904);
nor UO_231 (O_231,N_9943,N_9038);
nor UO_232 (O_232,N_9545,N_9451);
xnor UO_233 (O_233,N_9123,N_9876);
nand UO_234 (O_234,N_9772,N_9206);
or UO_235 (O_235,N_9230,N_9386);
and UO_236 (O_236,N_9915,N_9162);
nor UO_237 (O_237,N_9800,N_9315);
xor UO_238 (O_238,N_9700,N_9078);
or UO_239 (O_239,N_9811,N_9748);
nor UO_240 (O_240,N_9698,N_9628);
nor UO_241 (O_241,N_9532,N_9619);
or UO_242 (O_242,N_9046,N_9116);
and UO_243 (O_243,N_9496,N_9387);
nand UO_244 (O_244,N_9779,N_9600);
nand UO_245 (O_245,N_9118,N_9498);
xnor UO_246 (O_246,N_9973,N_9982);
and UO_247 (O_247,N_9374,N_9459);
or UO_248 (O_248,N_9914,N_9961);
or UO_249 (O_249,N_9173,N_9066);
nor UO_250 (O_250,N_9808,N_9993);
xnor UO_251 (O_251,N_9828,N_9862);
nor UO_252 (O_252,N_9491,N_9529);
xor UO_253 (O_253,N_9193,N_9136);
or UO_254 (O_254,N_9152,N_9159);
xnor UO_255 (O_255,N_9794,N_9951);
xnor UO_256 (O_256,N_9394,N_9935);
or UO_257 (O_257,N_9426,N_9310);
xor UO_258 (O_258,N_9790,N_9243);
nand UO_259 (O_259,N_9148,N_9768);
and UO_260 (O_260,N_9909,N_9244);
nor UO_261 (O_261,N_9213,N_9214);
nor UO_262 (O_262,N_9507,N_9860);
or UO_263 (O_263,N_9556,N_9490);
nor UO_264 (O_264,N_9606,N_9803);
and UO_265 (O_265,N_9651,N_9974);
nand UO_266 (O_266,N_9392,N_9008);
xnor UO_267 (O_267,N_9166,N_9379);
and UO_268 (O_268,N_9050,N_9239);
nand UO_269 (O_269,N_9916,N_9106);
nand UO_270 (O_270,N_9917,N_9863);
and UO_271 (O_271,N_9694,N_9472);
or UO_272 (O_272,N_9928,N_9888);
xnor UO_273 (O_273,N_9292,N_9316);
xnor UO_274 (O_274,N_9140,N_9224);
or UO_275 (O_275,N_9842,N_9057);
and UO_276 (O_276,N_9887,N_9156);
and UO_277 (O_277,N_9874,N_9573);
xor UO_278 (O_278,N_9526,N_9740);
nand UO_279 (O_279,N_9807,N_9345);
xnor UO_280 (O_280,N_9296,N_9515);
xnor UO_281 (O_281,N_9419,N_9172);
nand UO_282 (O_282,N_9541,N_9514);
or UO_283 (O_283,N_9321,N_9559);
nor UO_284 (O_284,N_9764,N_9340);
xor UO_285 (O_285,N_9344,N_9077);
nor UO_286 (O_286,N_9031,N_9205);
nand UO_287 (O_287,N_9289,N_9668);
nand UO_288 (O_288,N_9171,N_9403);
nor UO_289 (O_289,N_9088,N_9975);
nand UO_290 (O_290,N_9949,N_9020);
nor UO_291 (O_291,N_9497,N_9839);
nor UO_292 (O_292,N_9735,N_9994);
nand UO_293 (O_293,N_9897,N_9817);
or UO_294 (O_294,N_9369,N_9756);
or UO_295 (O_295,N_9820,N_9447);
or UO_296 (O_296,N_9335,N_9989);
and UO_297 (O_297,N_9467,N_9320);
or UO_298 (O_298,N_9952,N_9780);
xor UO_299 (O_299,N_9918,N_9284);
xnor UO_300 (O_300,N_9215,N_9599);
or UO_301 (O_301,N_9637,N_9695);
or UO_302 (O_302,N_9294,N_9505);
and UO_303 (O_303,N_9408,N_9250);
xor UO_304 (O_304,N_9703,N_9291);
xnor UO_305 (O_305,N_9865,N_9103);
and UO_306 (O_306,N_9799,N_9381);
and UO_307 (O_307,N_9539,N_9475);
nand UO_308 (O_308,N_9355,N_9434);
xnor UO_309 (O_309,N_9542,N_9033);
nor UO_310 (O_310,N_9160,N_9246);
nor UO_311 (O_311,N_9954,N_9765);
xnor UO_312 (O_312,N_9144,N_9513);
nor UO_313 (O_313,N_9309,N_9520);
nand UO_314 (O_314,N_9688,N_9815);
or UO_315 (O_315,N_9933,N_9268);
nand UO_316 (O_316,N_9286,N_9512);
and UO_317 (O_317,N_9398,N_9457);
and UO_318 (O_318,N_9649,N_9543);
or UO_319 (O_319,N_9667,N_9450);
or UO_320 (O_320,N_9609,N_9242);
and UO_321 (O_321,N_9278,N_9179);
nor UO_322 (O_322,N_9365,N_9614);
nor UO_323 (O_323,N_9693,N_9307);
nor UO_324 (O_324,N_9328,N_9342);
xor UO_325 (O_325,N_9750,N_9653);
nand UO_326 (O_326,N_9086,N_9776);
and UO_327 (O_327,N_9755,N_9784);
and UO_328 (O_328,N_9295,N_9055);
and UO_329 (O_329,N_9360,N_9956);
or UO_330 (O_330,N_9040,N_9736);
or UO_331 (O_331,N_9508,N_9469);
nor UO_332 (O_332,N_9882,N_9550);
nand UO_333 (O_333,N_9789,N_9902);
nor UO_334 (O_334,N_9069,N_9626);
nor UO_335 (O_335,N_9143,N_9869);
or UO_336 (O_336,N_9987,N_9090);
nand UO_337 (O_337,N_9690,N_9553);
nand UO_338 (O_338,N_9019,N_9194);
nand UO_339 (O_339,N_9642,N_9367);
and UO_340 (O_340,N_9059,N_9648);
nor UO_341 (O_341,N_9343,N_9950);
nand UO_342 (O_342,N_9990,N_9825);
nand UO_343 (O_343,N_9462,N_9025);
nor UO_344 (O_344,N_9685,N_9959);
or UO_345 (O_345,N_9338,N_9746);
and UO_346 (O_346,N_9719,N_9409);
and UO_347 (O_347,N_9567,N_9896);
or UO_348 (O_348,N_9676,N_9522);
or UO_349 (O_349,N_9254,N_9036);
nand UO_350 (O_350,N_9766,N_9444);
and UO_351 (O_351,N_9370,N_9236);
nor UO_352 (O_352,N_9068,N_9221);
or UO_353 (O_353,N_9126,N_9265);
or UO_354 (O_354,N_9783,N_9673);
xor UO_355 (O_355,N_9112,N_9283);
or UO_356 (O_356,N_9382,N_9996);
xnor UO_357 (O_357,N_9312,N_9349);
nor UO_358 (O_358,N_9705,N_9493);
nand UO_359 (O_359,N_9070,N_9687);
nand UO_360 (O_360,N_9796,N_9331);
xnor UO_361 (O_361,N_9375,N_9850);
or UO_362 (O_362,N_9267,N_9412);
and UO_363 (O_363,N_9385,N_9738);
nor UO_364 (O_364,N_9035,N_9107);
or UO_365 (O_365,N_9531,N_9402);
and UO_366 (O_366,N_9324,N_9678);
xor UO_367 (O_367,N_9041,N_9266);
xor UO_368 (O_368,N_9299,N_9601);
and UO_369 (O_369,N_9912,N_9232);
and UO_370 (O_370,N_9891,N_9980);
and UO_371 (O_371,N_9722,N_9407);
and UO_372 (O_372,N_9285,N_9028);
nand UO_373 (O_373,N_9983,N_9981);
nor UO_374 (O_374,N_9108,N_9691);
nand UO_375 (O_375,N_9699,N_9752);
or UO_376 (O_376,N_9004,N_9240);
nand UO_377 (O_377,N_9463,N_9879);
nand UO_378 (O_378,N_9085,N_9707);
nor UO_379 (O_379,N_9679,N_9674);
xor UO_380 (O_380,N_9500,N_9625);
nand UO_381 (O_381,N_9075,N_9231);
xnor UO_382 (O_382,N_9846,N_9810);
and UO_383 (O_383,N_9774,N_9760);
nor UO_384 (O_384,N_9697,N_9823);
nand UO_385 (O_385,N_9253,N_9323);
xnor UO_386 (O_386,N_9282,N_9414);
and UO_387 (O_387,N_9241,N_9495);
nand UO_388 (O_388,N_9822,N_9195);
xnor UO_389 (O_389,N_9481,N_9853);
xor UO_390 (O_390,N_9024,N_9439);
nand UO_391 (O_391,N_9504,N_9359);
xnor UO_392 (O_392,N_9054,N_9880);
or UO_393 (O_393,N_9440,N_9303);
or UO_394 (O_394,N_9364,N_9258);
xnor UO_395 (O_395,N_9022,N_9501);
xnor UO_396 (O_396,N_9546,N_9371);
and UO_397 (O_397,N_9654,N_9074);
xnor UO_398 (O_398,N_9201,N_9141);
nor UO_399 (O_399,N_9775,N_9744);
nand UO_400 (O_400,N_9203,N_9083);
xor UO_401 (O_401,N_9624,N_9290);
xor UO_402 (O_402,N_9225,N_9851);
nor UO_403 (O_403,N_9319,N_9884);
nand UO_404 (O_404,N_9018,N_9109);
and UO_405 (O_405,N_9638,N_9709);
nand UO_406 (O_406,N_9859,N_9551);
nand UO_407 (O_407,N_9101,N_9383);
or UO_408 (O_408,N_9634,N_9389);
and UO_409 (O_409,N_9037,N_9047);
nand UO_410 (O_410,N_9406,N_9770);
nand UO_411 (O_411,N_9787,N_9569);
nand UO_412 (O_412,N_9424,N_9923);
and UO_413 (O_413,N_9204,N_9841);
nor UO_414 (O_414,N_9165,N_9128);
nor UO_415 (O_415,N_9945,N_9920);
nor UO_416 (O_416,N_9797,N_9347);
nor UO_417 (O_417,N_9042,N_9163);
nor UO_418 (O_418,N_9104,N_9064);
nor UO_419 (O_419,N_9348,N_9612);
xor UO_420 (O_420,N_9252,N_9570);
xnor UO_421 (O_421,N_9801,N_9509);
nor UO_422 (O_422,N_9174,N_9287);
nor UO_423 (O_423,N_9701,N_9871);
or UO_424 (O_424,N_9976,N_9747);
or UO_425 (O_425,N_9835,N_9886);
nand UO_426 (O_426,N_9727,N_9960);
nor UO_427 (O_427,N_9249,N_9664);
nand UO_428 (O_428,N_9304,N_9301);
and UO_429 (O_429,N_9708,N_9593);
and UO_430 (O_430,N_9479,N_9145);
or UO_431 (O_431,N_9877,N_9376);
xor UO_432 (O_432,N_9549,N_9111);
nor UO_433 (O_433,N_9616,N_9051);
and UO_434 (O_434,N_9716,N_9913);
xnor UO_435 (O_435,N_9100,N_9089);
nand UO_436 (O_436,N_9742,N_9629);
and UO_437 (O_437,N_9211,N_9751);
xnor UO_438 (O_438,N_9134,N_9711);
and UO_439 (O_439,N_9704,N_9039);
xnor UO_440 (O_440,N_9102,N_9875);
and UO_441 (O_441,N_9732,N_9198);
xor UO_442 (O_442,N_9944,N_9300);
nor UO_443 (O_443,N_9391,N_9114);
and UO_444 (O_444,N_9906,N_9607);
and UO_445 (O_445,N_9521,N_9517);
xnor UO_446 (O_446,N_9405,N_9471);
nor UO_447 (O_447,N_9354,N_9843);
nor UO_448 (O_448,N_9574,N_9930);
nand UO_449 (O_449,N_9270,N_9255);
xnor UO_450 (O_450,N_9552,N_9445);
xnor UO_451 (O_451,N_9133,N_9819);
xor UO_452 (O_452,N_9506,N_9544);
xnor UO_453 (O_453,N_9259,N_9238);
nor UO_454 (O_454,N_9731,N_9680);
nor UO_455 (O_455,N_9146,N_9353);
nand UO_456 (O_456,N_9432,N_9706);
nor UO_457 (O_457,N_9659,N_9753);
nor UO_458 (O_458,N_9130,N_9157);
and UO_459 (O_459,N_9098,N_9777);
xor UO_460 (O_460,N_9207,N_9538);
and UO_461 (O_461,N_9864,N_9729);
nand UO_462 (O_462,N_9958,N_9565);
and UO_463 (O_463,N_9494,N_9861);
nor UO_464 (O_464,N_9739,N_9519);
nor UO_465 (O_465,N_9274,N_9222);
and UO_466 (O_466,N_9251,N_9032);
or UO_467 (O_467,N_9273,N_9079);
or UO_468 (O_468,N_9578,N_9362);
or UO_469 (O_469,N_9149,N_9298);
or UO_470 (O_470,N_9562,N_9010);
xnor UO_471 (O_471,N_9640,N_9903);
xor UO_472 (O_472,N_9595,N_9702);
nor UO_473 (O_473,N_9584,N_9129);
and UO_474 (O_474,N_9489,N_9848);
nor UO_475 (O_475,N_9388,N_9187);
or UO_476 (O_476,N_9317,N_9226);
nor UO_477 (O_477,N_9948,N_9337);
nand UO_478 (O_478,N_9922,N_9281);
nor UO_479 (O_479,N_9503,N_9329);
nor UO_480 (O_480,N_9870,N_9885);
and UO_481 (O_481,N_9745,N_9977);
xnor UO_482 (O_482,N_9476,N_9460);
or UO_483 (O_483,N_9431,N_9577);
and UO_484 (O_484,N_9404,N_9397);
nor UO_485 (O_485,N_9946,N_9443);
and UO_486 (O_486,N_9062,N_9423);
xor UO_487 (O_487,N_9158,N_9485);
or UO_488 (O_488,N_9235,N_9352);
xnor UO_489 (O_489,N_9733,N_9892);
nand UO_490 (O_490,N_9662,N_9488);
or UO_491 (O_491,N_9256,N_9350);
nand UO_492 (O_492,N_9767,N_9421);
and UO_493 (O_493,N_9113,N_9067);
nor UO_494 (O_494,N_9761,N_9615);
or UO_495 (O_495,N_9537,N_9474);
xnor UO_496 (O_496,N_9608,N_9856);
nor UO_497 (O_497,N_9717,N_9065);
nand UO_498 (O_498,N_9681,N_9121);
xnor UO_499 (O_499,N_9964,N_9125);
nand UO_500 (O_500,N_9549,N_9025);
and UO_501 (O_501,N_9032,N_9774);
or UO_502 (O_502,N_9260,N_9237);
and UO_503 (O_503,N_9651,N_9858);
and UO_504 (O_504,N_9189,N_9510);
xor UO_505 (O_505,N_9113,N_9758);
and UO_506 (O_506,N_9106,N_9268);
or UO_507 (O_507,N_9845,N_9685);
nand UO_508 (O_508,N_9518,N_9569);
xor UO_509 (O_509,N_9360,N_9768);
or UO_510 (O_510,N_9229,N_9570);
xnor UO_511 (O_511,N_9390,N_9943);
xnor UO_512 (O_512,N_9981,N_9422);
xnor UO_513 (O_513,N_9044,N_9641);
and UO_514 (O_514,N_9376,N_9125);
nor UO_515 (O_515,N_9937,N_9906);
nand UO_516 (O_516,N_9047,N_9140);
nor UO_517 (O_517,N_9622,N_9531);
or UO_518 (O_518,N_9784,N_9628);
and UO_519 (O_519,N_9925,N_9090);
nand UO_520 (O_520,N_9481,N_9892);
nor UO_521 (O_521,N_9437,N_9136);
and UO_522 (O_522,N_9636,N_9119);
nand UO_523 (O_523,N_9876,N_9619);
or UO_524 (O_524,N_9725,N_9089);
nand UO_525 (O_525,N_9657,N_9494);
and UO_526 (O_526,N_9082,N_9504);
and UO_527 (O_527,N_9041,N_9141);
or UO_528 (O_528,N_9338,N_9741);
and UO_529 (O_529,N_9515,N_9370);
nand UO_530 (O_530,N_9100,N_9926);
nor UO_531 (O_531,N_9530,N_9921);
nand UO_532 (O_532,N_9179,N_9858);
nor UO_533 (O_533,N_9050,N_9531);
xnor UO_534 (O_534,N_9836,N_9198);
or UO_535 (O_535,N_9189,N_9325);
nand UO_536 (O_536,N_9078,N_9714);
nor UO_537 (O_537,N_9678,N_9413);
or UO_538 (O_538,N_9131,N_9080);
nand UO_539 (O_539,N_9727,N_9289);
xor UO_540 (O_540,N_9471,N_9731);
or UO_541 (O_541,N_9072,N_9884);
and UO_542 (O_542,N_9061,N_9247);
xor UO_543 (O_543,N_9740,N_9972);
xnor UO_544 (O_544,N_9770,N_9422);
or UO_545 (O_545,N_9498,N_9176);
and UO_546 (O_546,N_9455,N_9628);
nor UO_547 (O_547,N_9210,N_9334);
xnor UO_548 (O_548,N_9971,N_9687);
or UO_549 (O_549,N_9924,N_9437);
or UO_550 (O_550,N_9380,N_9528);
xnor UO_551 (O_551,N_9316,N_9853);
nor UO_552 (O_552,N_9799,N_9454);
and UO_553 (O_553,N_9799,N_9428);
and UO_554 (O_554,N_9034,N_9108);
xnor UO_555 (O_555,N_9631,N_9480);
xnor UO_556 (O_556,N_9093,N_9250);
xor UO_557 (O_557,N_9054,N_9412);
and UO_558 (O_558,N_9505,N_9224);
xor UO_559 (O_559,N_9121,N_9747);
nand UO_560 (O_560,N_9456,N_9498);
nor UO_561 (O_561,N_9032,N_9233);
xnor UO_562 (O_562,N_9376,N_9787);
xor UO_563 (O_563,N_9894,N_9767);
and UO_564 (O_564,N_9444,N_9818);
nor UO_565 (O_565,N_9267,N_9530);
xor UO_566 (O_566,N_9921,N_9739);
nor UO_567 (O_567,N_9923,N_9462);
nand UO_568 (O_568,N_9463,N_9160);
xor UO_569 (O_569,N_9978,N_9950);
xnor UO_570 (O_570,N_9568,N_9239);
or UO_571 (O_571,N_9345,N_9019);
nor UO_572 (O_572,N_9165,N_9879);
or UO_573 (O_573,N_9360,N_9212);
nor UO_574 (O_574,N_9234,N_9306);
xnor UO_575 (O_575,N_9546,N_9988);
nor UO_576 (O_576,N_9749,N_9784);
or UO_577 (O_577,N_9044,N_9065);
nand UO_578 (O_578,N_9250,N_9083);
or UO_579 (O_579,N_9593,N_9438);
or UO_580 (O_580,N_9538,N_9383);
xnor UO_581 (O_581,N_9287,N_9172);
nand UO_582 (O_582,N_9668,N_9039);
nand UO_583 (O_583,N_9400,N_9260);
xor UO_584 (O_584,N_9426,N_9448);
nand UO_585 (O_585,N_9930,N_9832);
and UO_586 (O_586,N_9865,N_9459);
and UO_587 (O_587,N_9950,N_9948);
xnor UO_588 (O_588,N_9881,N_9673);
or UO_589 (O_589,N_9656,N_9578);
nand UO_590 (O_590,N_9178,N_9804);
xor UO_591 (O_591,N_9084,N_9412);
nand UO_592 (O_592,N_9790,N_9463);
and UO_593 (O_593,N_9936,N_9895);
and UO_594 (O_594,N_9572,N_9218);
nand UO_595 (O_595,N_9099,N_9804);
and UO_596 (O_596,N_9775,N_9101);
nor UO_597 (O_597,N_9689,N_9862);
and UO_598 (O_598,N_9978,N_9070);
and UO_599 (O_599,N_9749,N_9610);
nor UO_600 (O_600,N_9349,N_9389);
or UO_601 (O_601,N_9928,N_9296);
nor UO_602 (O_602,N_9684,N_9322);
nor UO_603 (O_603,N_9959,N_9139);
and UO_604 (O_604,N_9708,N_9223);
and UO_605 (O_605,N_9082,N_9645);
nor UO_606 (O_606,N_9213,N_9480);
or UO_607 (O_607,N_9417,N_9464);
nand UO_608 (O_608,N_9888,N_9435);
xor UO_609 (O_609,N_9232,N_9972);
nand UO_610 (O_610,N_9766,N_9418);
xor UO_611 (O_611,N_9266,N_9014);
and UO_612 (O_612,N_9622,N_9297);
or UO_613 (O_613,N_9962,N_9780);
nor UO_614 (O_614,N_9288,N_9864);
xor UO_615 (O_615,N_9458,N_9689);
nand UO_616 (O_616,N_9414,N_9661);
nand UO_617 (O_617,N_9673,N_9938);
and UO_618 (O_618,N_9840,N_9951);
and UO_619 (O_619,N_9512,N_9214);
nor UO_620 (O_620,N_9287,N_9450);
nand UO_621 (O_621,N_9502,N_9229);
or UO_622 (O_622,N_9627,N_9006);
or UO_623 (O_623,N_9150,N_9903);
xnor UO_624 (O_624,N_9999,N_9952);
nand UO_625 (O_625,N_9698,N_9160);
nand UO_626 (O_626,N_9838,N_9916);
xor UO_627 (O_627,N_9763,N_9767);
and UO_628 (O_628,N_9485,N_9976);
nor UO_629 (O_629,N_9903,N_9165);
nor UO_630 (O_630,N_9886,N_9059);
or UO_631 (O_631,N_9508,N_9053);
xnor UO_632 (O_632,N_9883,N_9421);
and UO_633 (O_633,N_9313,N_9571);
nor UO_634 (O_634,N_9128,N_9004);
nand UO_635 (O_635,N_9406,N_9109);
nand UO_636 (O_636,N_9208,N_9455);
and UO_637 (O_637,N_9351,N_9300);
and UO_638 (O_638,N_9900,N_9301);
or UO_639 (O_639,N_9517,N_9262);
xor UO_640 (O_640,N_9886,N_9233);
or UO_641 (O_641,N_9211,N_9047);
xnor UO_642 (O_642,N_9545,N_9946);
or UO_643 (O_643,N_9885,N_9332);
xnor UO_644 (O_644,N_9485,N_9739);
nand UO_645 (O_645,N_9896,N_9278);
xnor UO_646 (O_646,N_9350,N_9170);
or UO_647 (O_647,N_9485,N_9489);
nand UO_648 (O_648,N_9132,N_9673);
xor UO_649 (O_649,N_9724,N_9121);
nor UO_650 (O_650,N_9180,N_9465);
nor UO_651 (O_651,N_9797,N_9607);
nor UO_652 (O_652,N_9321,N_9282);
and UO_653 (O_653,N_9031,N_9324);
and UO_654 (O_654,N_9590,N_9905);
nand UO_655 (O_655,N_9456,N_9720);
and UO_656 (O_656,N_9620,N_9116);
or UO_657 (O_657,N_9032,N_9886);
xor UO_658 (O_658,N_9455,N_9996);
or UO_659 (O_659,N_9320,N_9840);
xnor UO_660 (O_660,N_9655,N_9517);
nor UO_661 (O_661,N_9498,N_9984);
or UO_662 (O_662,N_9619,N_9558);
nand UO_663 (O_663,N_9202,N_9352);
xor UO_664 (O_664,N_9529,N_9473);
nand UO_665 (O_665,N_9408,N_9908);
xnor UO_666 (O_666,N_9728,N_9027);
or UO_667 (O_667,N_9266,N_9028);
xnor UO_668 (O_668,N_9414,N_9922);
nor UO_669 (O_669,N_9165,N_9275);
and UO_670 (O_670,N_9374,N_9664);
xor UO_671 (O_671,N_9921,N_9723);
nor UO_672 (O_672,N_9941,N_9466);
or UO_673 (O_673,N_9749,N_9210);
nor UO_674 (O_674,N_9899,N_9081);
or UO_675 (O_675,N_9218,N_9222);
or UO_676 (O_676,N_9001,N_9261);
nor UO_677 (O_677,N_9908,N_9700);
nand UO_678 (O_678,N_9889,N_9583);
nand UO_679 (O_679,N_9879,N_9984);
nor UO_680 (O_680,N_9865,N_9033);
or UO_681 (O_681,N_9227,N_9901);
nand UO_682 (O_682,N_9444,N_9675);
nor UO_683 (O_683,N_9122,N_9011);
nor UO_684 (O_684,N_9172,N_9595);
and UO_685 (O_685,N_9091,N_9691);
nand UO_686 (O_686,N_9570,N_9921);
nand UO_687 (O_687,N_9029,N_9220);
nand UO_688 (O_688,N_9774,N_9288);
nand UO_689 (O_689,N_9595,N_9755);
xnor UO_690 (O_690,N_9265,N_9536);
and UO_691 (O_691,N_9242,N_9728);
nor UO_692 (O_692,N_9328,N_9804);
and UO_693 (O_693,N_9713,N_9830);
nor UO_694 (O_694,N_9201,N_9282);
nor UO_695 (O_695,N_9433,N_9410);
or UO_696 (O_696,N_9467,N_9776);
xor UO_697 (O_697,N_9967,N_9881);
or UO_698 (O_698,N_9271,N_9312);
and UO_699 (O_699,N_9593,N_9373);
nand UO_700 (O_700,N_9307,N_9343);
nor UO_701 (O_701,N_9441,N_9037);
nor UO_702 (O_702,N_9356,N_9622);
xnor UO_703 (O_703,N_9910,N_9835);
xnor UO_704 (O_704,N_9594,N_9973);
or UO_705 (O_705,N_9341,N_9880);
and UO_706 (O_706,N_9069,N_9002);
nor UO_707 (O_707,N_9248,N_9657);
nor UO_708 (O_708,N_9810,N_9301);
nor UO_709 (O_709,N_9126,N_9792);
xor UO_710 (O_710,N_9234,N_9681);
or UO_711 (O_711,N_9597,N_9651);
nor UO_712 (O_712,N_9384,N_9919);
or UO_713 (O_713,N_9700,N_9940);
nand UO_714 (O_714,N_9497,N_9268);
or UO_715 (O_715,N_9075,N_9794);
or UO_716 (O_716,N_9665,N_9186);
and UO_717 (O_717,N_9382,N_9789);
nand UO_718 (O_718,N_9153,N_9119);
nor UO_719 (O_719,N_9625,N_9690);
xor UO_720 (O_720,N_9259,N_9998);
and UO_721 (O_721,N_9738,N_9485);
xnor UO_722 (O_722,N_9071,N_9323);
or UO_723 (O_723,N_9693,N_9242);
nor UO_724 (O_724,N_9901,N_9061);
and UO_725 (O_725,N_9803,N_9873);
or UO_726 (O_726,N_9296,N_9010);
nor UO_727 (O_727,N_9154,N_9059);
nor UO_728 (O_728,N_9212,N_9774);
or UO_729 (O_729,N_9860,N_9206);
nor UO_730 (O_730,N_9836,N_9546);
nand UO_731 (O_731,N_9861,N_9408);
nand UO_732 (O_732,N_9307,N_9177);
nor UO_733 (O_733,N_9378,N_9508);
nand UO_734 (O_734,N_9942,N_9685);
or UO_735 (O_735,N_9374,N_9651);
or UO_736 (O_736,N_9237,N_9486);
nand UO_737 (O_737,N_9708,N_9421);
nand UO_738 (O_738,N_9821,N_9202);
xnor UO_739 (O_739,N_9340,N_9538);
nand UO_740 (O_740,N_9506,N_9535);
nor UO_741 (O_741,N_9034,N_9945);
nand UO_742 (O_742,N_9102,N_9171);
xor UO_743 (O_743,N_9213,N_9323);
and UO_744 (O_744,N_9080,N_9400);
and UO_745 (O_745,N_9295,N_9022);
xor UO_746 (O_746,N_9733,N_9748);
nor UO_747 (O_747,N_9131,N_9382);
or UO_748 (O_748,N_9419,N_9131);
and UO_749 (O_749,N_9541,N_9638);
or UO_750 (O_750,N_9553,N_9030);
nand UO_751 (O_751,N_9261,N_9926);
or UO_752 (O_752,N_9815,N_9450);
xnor UO_753 (O_753,N_9067,N_9369);
nor UO_754 (O_754,N_9734,N_9759);
and UO_755 (O_755,N_9666,N_9219);
and UO_756 (O_756,N_9399,N_9461);
nand UO_757 (O_757,N_9829,N_9102);
xnor UO_758 (O_758,N_9833,N_9037);
xnor UO_759 (O_759,N_9020,N_9639);
and UO_760 (O_760,N_9074,N_9778);
nand UO_761 (O_761,N_9162,N_9728);
nor UO_762 (O_762,N_9836,N_9986);
and UO_763 (O_763,N_9801,N_9374);
or UO_764 (O_764,N_9229,N_9899);
nor UO_765 (O_765,N_9923,N_9170);
or UO_766 (O_766,N_9627,N_9337);
and UO_767 (O_767,N_9499,N_9153);
xnor UO_768 (O_768,N_9580,N_9565);
or UO_769 (O_769,N_9981,N_9444);
and UO_770 (O_770,N_9445,N_9821);
xor UO_771 (O_771,N_9608,N_9631);
xnor UO_772 (O_772,N_9226,N_9935);
xor UO_773 (O_773,N_9144,N_9910);
nand UO_774 (O_774,N_9753,N_9557);
nor UO_775 (O_775,N_9185,N_9917);
nor UO_776 (O_776,N_9978,N_9940);
and UO_777 (O_777,N_9350,N_9000);
xor UO_778 (O_778,N_9766,N_9831);
nand UO_779 (O_779,N_9221,N_9468);
xnor UO_780 (O_780,N_9027,N_9687);
or UO_781 (O_781,N_9959,N_9476);
xnor UO_782 (O_782,N_9221,N_9295);
xnor UO_783 (O_783,N_9420,N_9022);
nor UO_784 (O_784,N_9016,N_9951);
and UO_785 (O_785,N_9593,N_9627);
or UO_786 (O_786,N_9622,N_9689);
xnor UO_787 (O_787,N_9428,N_9796);
xnor UO_788 (O_788,N_9887,N_9858);
xnor UO_789 (O_789,N_9239,N_9681);
or UO_790 (O_790,N_9010,N_9294);
nor UO_791 (O_791,N_9640,N_9570);
nand UO_792 (O_792,N_9352,N_9795);
or UO_793 (O_793,N_9434,N_9909);
or UO_794 (O_794,N_9471,N_9377);
and UO_795 (O_795,N_9095,N_9848);
or UO_796 (O_796,N_9056,N_9761);
nand UO_797 (O_797,N_9899,N_9672);
nand UO_798 (O_798,N_9576,N_9392);
and UO_799 (O_799,N_9012,N_9752);
or UO_800 (O_800,N_9162,N_9274);
xnor UO_801 (O_801,N_9840,N_9400);
nor UO_802 (O_802,N_9093,N_9529);
xnor UO_803 (O_803,N_9522,N_9168);
and UO_804 (O_804,N_9420,N_9469);
nand UO_805 (O_805,N_9682,N_9283);
xnor UO_806 (O_806,N_9464,N_9965);
nand UO_807 (O_807,N_9873,N_9540);
or UO_808 (O_808,N_9726,N_9812);
nand UO_809 (O_809,N_9326,N_9184);
nor UO_810 (O_810,N_9658,N_9354);
nand UO_811 (O_811,N_9845,N_9533);
and UO_812 (O_812,N_9909,N_9710);
or UO_813 (O_813,N_9906,N_9301);
nand UO_814 (O_814,N_9964,N_9431);
xor UO_815 (O_815,N_9410,N_9955);
and UO_816 (O_816,N_9151,N_9014);
nor UO_817 (O_817,N_9844,N_9621);
nor UO_818 (O_818,N_9752,N_9404);
or UO_819 (O_819,N_9644,N_9105);
and UO_820 (O_820,N_9811,N_9226);
xor UO_821 (O_821,N_9990,N_9350);
nor UO_822 (O_822,N_9554,N_9201);
and UO_823 (O_823,N_9954,N_9565);
and UO_824 (O_824,N_9247,N_9008);
xor UO_825 (O_825,N_9303,N_9116);
nand UO_826 (O_826,N_9806,N_9102);
and UO_827 (O_827,N_9349,N_9642);
xor UO_828 (O_828,N_9466,N_9115);
or UO_829 (O_829,N_9321,N_9211);
nor UO_830 (O_830,N_9669,N_9562);
xor UO_831 (O_831,N_9303,N_9115);
or UO_832 (O_832,N_9807,N_9253);
nand UO_833 (O_833,N_9222,N_9912);
and UO_834 (O_834,N_9581,N_9943);
or UO_835 (O_835,N_9633,N_9432);
nand UO_836 (O_836,N_9754,N_9842);
nor UO_837 (O_837,N_9342,N_9524);
xor UO_838 (O_838,N_9309,N_9787);
nor UO_839 (O_839,N_9839,N_9011);
or UO_840 (O_840,N_9262,N_9469);
xor UO_841 (O_841,N_9321,N_9007);
or UO_842 (O_842,N_9354,N_9167);
and UO_843 (O_843,N_9226,N_9401);
xor UO_844 (O_844,N_9012,N_9543);
and UO_845 (O_845,N_9101,N_9312);
xor UO_846 (O_846,N_9804,N_9808);
nand UO_847 (O_847,N_9355,N_9693);
nand UO_848 (O_848,N_9701,N_9467);
or UO_849 (O_849,N_9000,N_9076);
nor UO_850 (O_850,N_9799,N_9159);
nor UO_851 (O_851,N_9124,N_9959);
nand UO_852 (O_852,N_9408,N_9254);
or UO_853 (O_853,N_9352,N_9673);
xor UO_854 (O_854,N_9928,N_9190);
nand UO_855 (O_855,N_9118,N_9342);
or UO_856 (O_856,N_9339,N_9486);
nor UO_857 (O_857,N_9682,N_9876);
and UO_858 (O_858,N_9463,N_9065);
nor UO_859 (O_859,N_9943,N_9987);
and UO_860 (O_860,N_9040,N_9740);
or UO_861 (O_861,N_9161,N_9767);
and UO_862 (O_862,N_9240,N_9012);
xnor UO_863 (O_863,N_9250,N_9008);
or UO_864 (O_864,N_9100,N_9902);
nor UO_865 (O_865,N_9364,N_9197);
or UO_866 (O_866,N_9444,N_9116);
nand UO_867 (O_867,N_9751,N_9791);
xor UO_868 (O_868,N_9448,N_9702);
xor UO_869 (O_869,N_9276,N_9639);
and UO_870 (O_870,N_9506,N_9015);
xnor UO_871 (O_871,N_9582,N_9556);
xnor UO_872 (O_872,N_9616,N_9795);
nand UO_873 (O_873,N_9442,N_9865);
xor UO_874 (O_874,N_9107,N_9566);
xor UO_875 (O_875,N_9084,N_9858);
and UO_876 (O_876,N_9973,N_9635);
or UO_877 (O_877,N_9143,N_9972);
and UO_878 (O_878,N_9940,N_9315);
xor UO_879 (O_879,N_9148,N_9281);
nor UO_880 (O_880,N_9114,N_9040);
or UO_881 (O_881,N_9356,N_9915);
xnor UO_882 (O_882,N_9314,N_9830);
and UO_883 (O_883,N_9302,N_9143);
and UO_884 (O_884,N_9494,N_9661);
nor UO_885 (O_885,N_9373,N_9989);
xnor UO_886 (O_886,N_9393,N_9465);
nor UO_887 (O_887,N_9045,N_9713);
and UO_888 (O_888,N_9287,N_9008);
or UO_889 (O_889,N_9057,N_9680);
or UO_890 (O_890,N_9821,N_9099);
xnor UO_891 (O_891,N_9178,N_9246);
and UO_892 (O_892,N_9074,N_9846);
nand UO_893 (O_893,N_9417,N_9471);
nand UO_894 (O_894,N_9382,N_9892);
xnor UO_895 (O_895,N_9043,N_9811);
or UO_896 (O_896,N_9549,N_9789);
nor UO_897 (O_897,N_9227,N_9378);
nand UO_898 (O_898,N_9400,N_9185);
nor UO_899 (O_899,N_9139,N_9374);
and UO_900 (O_900,N_9144,N_9625);
nand UO_901 (O_901,N_9832,N_9634);
nand UO_902 (O_902,N_9362,N_9615);
or UO_903 (O_903,N_9990,N_9213);
and UO_904 (O_904,N_9475,N_9003);
or UO_905 (O_905,N_9214,N_9992);
xnor UO_906 (O_906,N_9013,N_9688);
xor UO_907 (O_907,N_9330,N_9728);
and UO_908 (O_908,N_9033,N_9606);
nor UO_909 (O_909,N_9172,N_9586);
or UO_910 (O_910,N_9900,N_9869);
and UO_911 (O_911,N_9251,N_9055);
xor UO_912 (O_912,N_9921,N_9422);
or UO_913 (O_913,N_9459,N_9506);
and UO_914 (O_914,N_9793,N_9554);
xnor UO_915 (O_915,N_9407,N_9680);
and UO_916 (O_916,N_9174,N_9541);
or UO_917 (O_917,N_9109,N_9798);
nand UO_918 (O_918,N_9968,N_9305);
xor UO_919 (O_919,N_9639,N_9424);
and UO_920 (O_920,N_9609,N_9708);
or UO_921 (O_921,N_9155,N_9548);
or UO_922 (O_922,N_9680,N_9115);
xor UO_923 (O_923,N_9522,N_9701);
and UO_924 (O_924,N_9955,N_9124);
nand UO_925 (O_925,N_9092,N_9542);
or UO_926 (O_926,N_9803,N_9231);
or UO_927 (O_927,N_9086,N_9514);
or UO_928 (O_928,N_9089,N_9146);
nand UO_929 (O_929,N_9397,N_9611);
and UO_930 (O_930,N_9034,N_9263);
and UO_931 (O_931,N_9171,N_9745);
nor UO_932 (O_932,N_9065,N_9113);
xnor UO_933 (O_933,N_9649,N_9839);
nor UO_934 (O_934,N_9039,N_9846);
xor UO_935 (O_935,N_9582,N_9279);
xnor UO_936 (O_936,N_9386,N_9528);
nor UO_937 (O_937,N_9613,N_9207);
nor UO_938 (O_938,N_9048,N_9278);
xor UO_939 (O_939,N_9837,N_9729);
nor UO_940 (O_940,N_9359,N_9516);
xor UO_941 (O_941,N_9438,N_9356);
or UO_942 (O_942,N_9694,N_9997);
nand UO_943 (O_943,N_9666,N_9089);
and UO_944 (O_944,N_9332,N_9840);
or UO_945 (O_945,N_9747,N_9359);
or UO_946 (O_946,N_9795,N_9772);
xor UO_947 (O_947,N_9087,N_9792);
or UO_948 (O_948,N_9801,N_9187);
nand UO_949 (O_949,N_9107,N_9816);
or UO_950 (O_950,N_9010,N_9979);
or UO_951 (O_951,N_9531,N_9808);
and UO_952 (O_952,N_9299,N_9054);
nor UO_953 (O_953,N_9796,N_9548);
nor UO_954 (O_954,N_9642,N_9113);
and UO_955 (O_955,N_9818,N_9750);
nand UO_956 (O_956,N_9951,N_9789);
xnor UO_957 (O_957,N_9632,N_9327);
or UO_958 (O_958,N_9249,N_9359);
or UO_959 (O_959,N_9126,N_9924);
or UO_960 (O_960,N_9750,N_9351);
nor UO_961 (O_961,N_9473,N_9135);
or UO_962 (O_962,N_9087,N_9421);
nor UO_963 (O_963,N_9009,N_9274);
or UO_964 (O_964,N_9654,N_9710);
nand UO_965 (O_965,N_9574,N_9133);
nor UO_966 (O_966,N_9529,N_9031);
xor UO_967 (O_967,N_9187,N_9908);
nand UO_968 (O_968,N_9053,N_9267);
nand UO_969 (O_969,N_9327,N_9841);
nor UO_970 (O_970,N_9981,N_9056);
nor UO_971 (O_971,N_9329,N_9074);
nor UO_972 (O_972,N_9598,N_9941);
and UO_973 (O_973,N_9774,N_9833);
and UO_974 (O_974,N_9375,N_9909);
nor UO_975 (O_975,N_9856,N_9846);
nand UO_976 (O_976,N_9779,N_9041);
nor UO_977 (O_977,N_9265,N_9479);
nor UO_978 (O_978,N_9162,N_9187);
xor UO_979 (O_979,N_9843,N_9566);
nor UO_980 (O_980,N_9408,N_9622);
and UO_981 (O_981,N_9631,N_9069);
and UO_982 (O_982,N_9632,N_9030);
nand UO_983 (O_983,N_9062,N_9468);
nand UO_984 (O_984,N_9921,N_9358);
and UO_985 (O_985,N_9470,N_9209);
and UO_986 (O_986,N_9439,N_9498);
and UO_987 (O_987,N_9241,N_9513);
nand UO_988 (O_988,N_9036,N_9079);
and UO_989 (O_989,N_9693,N_9338);
and UO_990 (O_990,N_9430,N_9128);
nor UO_991 (O_991,N_9645,N_9399);
or UO_992 (O_992,N_9687,N_9751);
nand UO_993 (O_993,N_9809,N_9073);
nand UO_994 (O_994,N_9376,N_9722);
and UO_995 (O_995,N_9982,N_9719);
nor UO_996 (O_996,N_9575,N_9812);
and UO_997 (O_997,N_9896,N_9604);
nand UO_998 (O_998,N_9259,N_9847);
xnor UO_999 (O_999,N_9493,N_9842);
or UO_1000 (O_1000,N_9668,N_9061);
xor UO_1001 (O_1001,N_9953,N_9166);
and UO_1002 (O_1002,N_9301,N_9205);
and UO_1003 (O_1003,N_9002,N_9869);
xnor UO_1004 (O_1004,N_9653,N_9229);
xnor UO_1005 (O_1005,N_9599,N_9166);
and UO_1006 (O_1006,N_9582,N_9136);
and UO_1007 (O_1007,N_9850,N_9848);
and UO_1008 (O_1008,N_9081,N_9848);
and UO_1009 (O_1009,N_9546,N_9751);
and UO_1010 (O_1010,N_9153,N_9556);
and UO_1011 (O_1011,N_9672,N_9622);
xnor UO_1012 (O_1012,N_9615,N_9735);
nand UO_1013 (O_1013,N_9747,N_9572);
xnor UO_1014 (O_1014,N_9952,N_9400);
xnor UO_1015 (O_1015,N_9168,N_9921);
or UO_1016 (O_1016,N_9710,N_9884);
xor UO_1017 (O_1017,N_9158,N_9629);
xnor UO_1018 (O_1018,N_9343,N_9829);
xnor UO_1019 (O_1019,N_9537,N_9001);
or UO_1020 (O_1020,N_9047,N_9727);
nand UO_1021 (O_1021,N_9884,N_9719);
and UO_1022 (O_1022,N_9591,N_9890);
or UO_1023 (O_1023,N_9389,N_9437);
nand UO_1024 (O_1024,N_9528,N_9107);
or UO_1025 (O_1025,N_9004,N_9008);
or UO_1026 (O_1026,N_9459,N_9089);
nand UO_1027 (O_1027,N_9102,N_9604);
nor UO_1028 (O_1028,N_9953,N_9304);
or UO_1029 (O_1029,N_9397,N_9174);
nand UO_1030 (O_1030,N_9718,N_9535);
and UO_1031 (O_1031,N_9667,N_9303);
and UO_1032 (O_1032,N_9490,N_9518);
or UO_1033 (O_1033,N_9150,N_9253);
nor UO_1034 (O_1034,N_9750,N_9148);
and UO_1035 (O_1035,N_9538,N_9577);
nand UO_1036 (O_1036,N_9170,N_9352);
or UO_1037 (O_1037,N_9958,N_9249);
nor UO_1038 (O_1038,N_9629,N_9198);
or UO_1039 (O_1039,N_9077,N_9382);
or UO_1040 (O_1040,N_9352,N_9680);
and UO_1041 (O_1041,N_9289,N_9505);
xnor UO_1042 (O_1042,N_9599,N_9816);
xor UO_1043 (O_1043,N_9972,N_9692);
and UO_1044 (O_1044,N_9576,N_9258);
nor UO_1045 (O_1045,N_9038,N_9306);
and UO_1046 (O_1046,N_9468,N_9510);
xnor UO_1047 (O_1047,N_9629,N_9133);
xor UO_1048 (O_1048,N_9232,N_9003);
nand UO_1049 (O_1049,N_9568,N_9434);
xor UO_1050 (O_1050,N_9755,N_9986);
or UO_1051 (O_1051,N_9964,N_9692);
or UO_1052 (O_1052,N_9888,N_9714);
nand UO_1053 (O_1053,N_9537,N_9276);
or UO_1054 (O_1054,N_9079,N_9708);
nand UO_1055 (O_1055,N_9576,N_9811);
and UO_1056 (O_1056,N_9550,N_9881);
nor UO_1057 (O_1057,N_9146,N_9014);
nor UO_1058 (O_1058,N_9376,N_9495);
xnor UO_1059 (O_1059,N_9336,N_9368);
or UO_1060 (O_1060,N_9939,N_9259);
xnor UO_1061 (O_1061,N_9084,N_9939);
nor UO_1062 (O_1062,N_9734,N_9970);
or UO_1063 (O_1063,N_9223,N_9811);
and UO_1064 (O_1064,N_9475,N_9133);
nand UO_1065 (O_1065,N_9839,N_9875);
or UO_1066 (O_1066,N_9025,N_9505);
xnor UO_1067 (O_1067,N_9327,N_9505);
or UO_1068 (O_1068,N_9977,N_9535);
and UO_1069 (O_1069,N_9199,N_9637);
or UO_1070 (O_1070,N_9842,N_9405);
or UO_1071 (O_1071,N_9762,N_9794);
and UO_1072 (O_1072,N_9526,N_9542);
nand UO_1073 (O_1073,N_9971,N_9004);
nand UO_1074 (O_1074,N_9271,N_9432);
and UO_1075 (O_1075,N_9057,N_9416);
nor UO_1076 (O_1076,N_9042,N_9569);
nand UO_1077 (O_1077,N_9438,N_9512);
xor UO_1078 (O_1078,N_9270,N_9427);
and UO_1079 (O_1079,N_9522,N_9100);
nand UO_1080 (O_1080,N_9332,N_9771);
and UO_1081 (O_1081,N_9885,N_9044);
nand UO_1082 (O_1082,N_9572,N_9528);
nor UO_1083 (O_1083,N_9590,N_9588);
or UO_1084 (O_1084,N_9878,N_9615);
and UO_1085 (O_1085,N_9560,N_9318);
xnor UO_1086 (O_1086,N_9624,N_9031);
or UO_1087 (O_1087,N_9213,N_9719);
xor UO_1088 (O_1088,N_9263,N_9823);
xor UO_1089 (O_1089,N_9625,N_9919);
xnor UO_1090 (O_1090,N_9391,N_9412);
and UO_1091 (O_1091,N_9644,N_9834);
and UO_1092 (O_1092,N_9886,N_9013);
and UO_1093 (O_1093,N_9922,N_9326);
xnor UO_1094 (O_1094,N_9590,N_9429);
or UO_1095 (O_1095,N_9533,N_9804);
xnor UO_1096 (O_1096,N_9311,N_9655);
nor UO_1097 (O_1097,N_9671,N_9442);
nand UO_1098 (O_1098,N_9782,N_9023);
and UO_1099 (O_1099,N_9121,N_9982);
and UO_1100 (O_1100,N_9224,N_9920);
nor UO_1101 (O_1101,N_9231,N_9755);
or UO_1102 (O_1102,N_9211,N_9457);
and UO_1103 (O_1103,N_9214,N_9726);
and UO_1104 (O_1104,N_9512,N_9911);
nand UO_1105 (O_1105,N_9815,N_9430);
and UO_1106 (O_1106,N_9431,N_9377);
or UO_1107 (O_1107,N_9248,N_9630);
and UO_1108 (O_1108,N_9708,N_9006);
or UO_1109 (O_1109,N_9663,N_9625);
or UO_1110 (O_1110,N_9191,N_9713);
or UO_1111 (O_1111,N_9772,N_9655);
nor UO_1112 (O_1112,N_9484,N_9826);
or UO_1113 (O_1113,N_9342,N_9990);
and UO_1114 (O_1114,N_9303,N_9408);
and UO_1115 (O_1115,N_9236,N_9994);
nand UO_1116 (O_1116,N_9016,N_9057);
nand UO_1117 (O_1117,N_9380,N_9119);
nor UO_1118 (O_1118,N_9470,N_9731);
xnor UO_1119 (O_1119,N_9962,N_9394);
nor UO_1120 (O_1120,N_9434,N_9051);
nand UO_1121 (O_1121,N_9808,N_9052);
nor UO_1122 (O_1122,N_9655,N_9579);
or UO_1123 (O_1123,N_9855,N_9995);
xnor UO_1124 (O_1124,N_9913,N_9926);
nor UO_1125 (O_1125,N_9344,N_9852);
xor UO_1126 (O_1126,N_9752,N_9010);
or UO_1127 (O_1127,N_9580,N_9750);
nor UO_1128 (O_1128,N_9914,N_9745);
or UO_1129 (O_1129,N_9765,N_9704);
or UO_1130 (O_1130,N_9875,N_9484);
and UO_1131 (O_1131,N_9864,N_9363);
and UO_1132 (O_1132,N_9679,N_9722);
and UO_1133 (O_1133,N_9438,N_9704);
xnor UO_1134 (O_1134,N_9863,N_9152);
and UO_1135 (O_1135,N_9044,N_9361);
nand UO_1136 (O_1136,N_9882,N_9535);
or UO_1137 (O_1137,N_9772,N_9543);
or UO_1138 (O_1138,N_9625,N_9423);
and UO_1139 (O_1139,N_9318,N_9543);
nand UO_1140 (O_1140,N_9943,N_9320);
xor UO_1141 (O_1141,N_9858,N_9868);
nor UO_1142 (O_1142,N_9376,N_9724);
nor UO_1143 (O_1143,N_9816,N_9980);
or UO_1144 (O_1144,N_9453,N_9673);
xnor UO_1145 (O_1145,N_9221,N_9204);
xnor UO_1146 (O_1146,N_9082,N_9436);
or UO_1147 (O_1147,N_9074,N_9864);
or UO_1148 (O_1148,N_9351,N_9431);
nor UO_1149 (O_1149,N_9713,N_9224);
and UO_1150 (O_1150,N_9049,N_9346);
nor UO_1151 (O_1151,N_9149,N_9981);
xnor UO_1152 (O_1152,N_9693,N_9584);
or UO_1153 (O_1153,N_9188,N_9802);
xnor UO_1154 (O_1154,N_9772,N_9815);
and UO_1155 (O_1155,N_9451,N_9141);
xor UO_1156 (O_1156,N_9158,N_9337);
and UO_1157 (O_1157,N_9060,N_9921);
nor UO_1158 (O_1158,N_9403,N_9040);
xnor UO_1159 (O_1159,N_9218,N_9106);
xnor UO_1160 (O_1160,N_9004,N_9970);
nand UO_1161 (O_1161,N_9450,N_9474);
xor UO_1162 (O_1162,N_9226,N_9093);
and UO_1163 (O_1163,N_9982,N_9596);
nand UO_1164 (O_1164,N_9646,N_9260);
and UO_1165 (O_1165,N_9227,N_9847);
nand UO_1166 (O_1166,N_9837,N_9881);
nor UO_1167 (O_1167,N_9561,N_9384);
nor UO_1168 (O_1168,N_9664,N_9232);
xor UO_1169 (O_1169,N_9886,N_9458);
nand UO_1170 (O_1170,N_9567,N_9601);
or UO_1171 (O_1171,N_9287,N_9760);
nor UO_1172 (O_1172,N_9492,N_9886);
nand UO_1173 (O_1173,N_9572,N_9193);
xor UO_1174 (O_1174,N_9497,N_9558);
nand UO_1175 (O_1175,N_9272,N_9471);
nand UO_1176 (O_1176,N_9151,N_9517);
xnor UO_1177 (O_1177,N_9274,N_9760);
or UO_1178 (O_1178,N_9647,N_9485);
and UO_1179 (O_1179,N_9727,N_9097);
and UO_1180 (O_1180,N_9143,N_9467);
nand UO_1181 (O_1181,N_9502,N_9703);
or UO_1182 (O_1182,N_9840,N_9333);
xor UO_1183 (O_1183,N_9229,N_9210);
or UO_1184 (O_1184,N_9533,N_9424);
nor UO_1185 (O_1185,N_9202,N_9362);
xor UO_1186 (O_1186,N_9709,N_9983);
or UO_1187 (O_1187,N_9585,N_9851);
xnor UO_1188 (O_1188,N_9390,N_9286);
and UO_1189 (O_1189,N_9096,N_9282);
nand UO_1190 (O_1190,N_9904,N_9380);
and UO_1191 (O_1191,N_9975,N_9058);
nand UO_1192 (O_1192,N_9942,N_9447);
nor UO_1193 (O_1193,N_9279,N_9125);
and UO_1194 (O_1194,N_9641,N_9881);
and UO_1195 (O_1195,N_9177,N_9630);
and UO_1196 (O_1196,N_9794,N_9432);
xnor UO_1197 (O_1197,N_9438,N_9831);
nor UO_1198 (O_1198,N_9847,N_9676);
nor UO_1199 (O_1199,N_9632,N_9072);
and UO_1200 (O_1200,N_9192,N_9842);
and UO_1201 (O_1201,N_9585,N_9576);
nor UO_1202 (O_1202,N_9647,N_9994);
or UO_1203 (O_1203,N_9389,N_9878);
or UO_1204 (O_1204,N_9223,N_9952);
xnor UO_1205 (O_1205,N_9801,N_9012);
or UO_1206 (O_1206,N_9894,N_9546);
xnor UO_1207 (O_1207,N_9916,N_9463);
nand UO_1208 (O_1208,N_9507,N_9009);
or UO_1209 (O_1209,N_9037,N_9524);
xnor UO_1210 (O_1210,N_9366,N_9775);
nor UO_1211 (O_1211,N_9263,N_9540);
xor UO_1212 (O_1212,N_9261,N_9229);
and UO_1213 (O_1213,N_9467,N_9730);
xnor UO_1214 (O_1214,N_9880,N_9521);
nor UO_1215 (O_1215,N_9225,N_9099);
nor UO_1216 (O_1216,N_9498,N_9680);
xnor UO_1217 (O_1217,N_9805,N_9646);
nor UO_1218 (O_1218,N_9571,N_9221);
and UO_1219 (O_1219,N_9081,N_9196);
nand UO_1220 (O_1220,N_9303,N_9945);
xor UO_1221 (O_1221,N_9403,N_9644);
nand UO_1222 (O_1222,N_9009,N_9973);
and UO_1223 (O_1223,N_9749,N_9137);
nand UO_1224 (O_1224,N_9708,N_9640);
xnor UO_1225 (O_1225,N_9113,N_9098);
and UO_1226 (O_1226,N_9399,N_9046);
and UO_1227 (O_1227,N_9200,N_9563);
nand UO_1228 (O_1228,N_9187,N_9562);
xor UO_1229 (O_1229,N_9540,N_9103);
or UO_1230 (O_1230,N_9846,N_9525);
and UO_1231 (O_1231,N_9704,N_9600);
xor UO_1232 (O_1232,N_9829,N_9301);
nor UO_1233 (O_1233,N_9436,N_9287);
xor UO_1234 (O_1234,N_9071,N_9180);
nor UO_1235 (O_1235,N_9585,N_9734);
xnor UO_1236 (O_1236,N_9688,N_9108);
nor UO_1237 (O_1237,N_9789,N_9848);
and UO_1238 (O_1238,N_9497,N_9108);
nor UO_1239 (O_1239,N_9195,N_9337);
or UO_1240 (O_1240,N_9888,N_9261);
nand UO_1241 (O_1241,N_9619,N_9970);
nor UO_1242 (O_1242,N_9376,N_9535);
nor UO_1243 (O_1243,N_9911,N_9122);
or UO_1244 (O_1244,N_9799,N_9814);
xnor UO_1245 (O_1245,N_9596,N_9220);
and UO_1246 (O_1246,N_9045,N_9786);
or UO_1247 (O_1247,N_9836,N_9672);
xor UO_1248 (O_1248,N_9449,N_9152);
xor UO_1249 (O_1249,N_9153,N_9567);
xnor UO_1250 (O_1250,N_9795,N_9755);
nor UO_1251 (O_1251,N_9989,N_9498);
nand UO_1252 (O_1252,N_9675,N_9964);
and UO_1253 (O_1253,N_9746,N_9571);
nor UO_1254 (O_1254,N_9494,N_9655);
nor UO_1255 (O_1255,N_9154,N_9960);
nand UO_1256 (O_1256,N_9357,N_9419);
or UO_1257 (O_1257,N_9144,N_9991);
nand UO_1258 (O_1258,N_9119,N_9866);
or UO_1259 (O_1259,N_9154,N_9009);
or UO_1260 (O_1260,N_9868,N_9741);
nor UO_1261 (O_1261,N_9245,N_9700);
and UO_1262 (O_1262,N_9893,N_9833);
xor UO_1263 (O_1263,N_9925,N_9323);
and UO_1264 (O_1264,N_9854,N_9588);
nand UO_1265 (O_1265,N_9615,N_9886);
or UO_1266 (O_1266,N_9657,N_9539);
xnor UO_1267 (O_1267,N_9327,N_9336);
nand UO_1268 (O_1268,N_9255,N_9049);
nand UO_1269 (O_1269,N_9223,N_9108);
and UO_1270 (O_1270,N_9463,N_9585);
nand UO_1271 (O_1271,N_9258,N_9723);
or UO_1272 (O_1272,N_9484,N_9623);
or UO_1273 (O_1273,N_9788,N_9215);
xor UO_1274 (O_1274,N_9724,N_9005);
xnor UO_1275 (O_1275,N_9639,N_9697);
and UO_1276 (O_1276,N_9085,N_9438);
and UO_1277 (O_1277,N_9184,N_9600);
and UO_1278 (O_1278,N_9526,N_9815);
xnor UO_1279 (O_1279,N_9072,N_9364);
and UO_1280 (O_1280,N_9981,N_9989);
nor UO_1281 (O_1281,N_9414,N_9883);
nor UO_1282 (O_1282,N_9144,N_9444);
or UO_1283 (O_1283,N_9965,N_9119);
and UO_1284 (O_1284,N_9933,N_9013);
and UO_1285 (O_1285,N_9588,N_9713);
nor UO_1286 (O_1286,N_9304,N_9474);
nor UO_1287 (O_1287,N_9834,N_9299);
nand UO_1288 (O_1288,N_9478,N_9779);
nand UO_1289 (O_1289,N_9487,N_9133);
nand UO_1290 (O_1290,N_9835,N_9751);
and UO_1291 (O_1291,N_9670,N_9782);
or UO_1292 (O_1292,N_9229,N_9848);
and UO_1293 (O_1293,N_9536,N_9951);
xor UO_1294 (O_1294,N_9248,N_9449);
xor UO_1295 (O_1295,N_9183,N_9749);
and UO_1296 (O_1296,N_9456,N_9728);
nor UO_1297 (O_1297,N_9993,N_9026);
nor UO_1298 (O_1298,N_9632,N_9227);
nor UO_1299 (O_1299,N_9666,N_9316);
or UO_1300 (O_1300,N_9164,N_9268);
or UO_1301 (O_1301,N_9727,N_9954);
or UO_1302 (O_1302,N_9005,N_9907);
nand UO_1303 (O_1303,N_9242,N_9514);
xnor UO_1304 (O_1304,N_9632,N_9552);
or UO_1305 (O_1305,N_9113,N_9837);
nand UO_1306 (O_1306,N_9613,N_9112);
or UO_1307 (O_1307,N_9607,N_9065);
nand UO_1308 (O_1308,N_9825,N_9565);
or UO_1309 (O_1309,N_9342,N_9672);
or UO_1310 (O_1310,N_9899,N_9996);
nor UO_1311 (O_1311,N_9805,N_9191);
nor UO_1312 (O_1312,N_9713,N_9075);
or UO_1313 (O_1313,N_9643,N_9411);
or UO_1314 (O_1314,N_9164,N_9686);
nand UO_1315 (O_1315,N_9964,N_9302);
and UO_1316 (O_1316,N_9814,N_9584);
nor UO_1317 (O_1317,N_9492,N_9276);
nor UO_1318 (O_1318,N_9922,N_9255);
nor UO_1319 (O_1319,N_9034,N_9412);
or UO_1320 (O_1320,N_9651,N_9406);
nand UO_1321 (O_1321,N_9966,N_9333);
nand UO_1322 (O_1322,N_9293,N_9719);
and UO_1323 (O_1323,N_9519,N_9319);
nor UO_1324 (O_1324,N_9586,N_9435);
xnor UO_1325 (O_1325,N_9652,N_9361);
xnor UO_1326 (O_1326,N_9892,N_9020);
nand UO_1327 (O_1327,N_9522,N_9693);
or UO_1328 (O_1328,N_9457,N_9685);
nor UO_1329 (O_1329,N_9003,N_9652);
or UO_1330 (O_1330,N_9180,N_9388);
xor UO_1331 (O_1331,N_9007,N_9690);
and UO_1332 (O_1332,N_9204,N_9785);
nand UO_1333 (O_1333,N_9830,N_9852);
xnor UO_1334 (O_1334,N_9238,N_9245);
and UO_1335 (O_1335,N_9718,N_9908);
or UO_1336 (O_1336,N_9330,N_9775);
or UO_1337 (O_1337,N_9459,N_9773);
and UO_1338 (O_1338,N_9426,N_9695);
xor UO_1339 (O_1339,N_9312,N_9915);
nand UO_1340 (O_1340,N_9776,N_9093);
or UO_1341 (O_1341,N_9841,N_9690);
or UO_1342 (O_1342,N_9296,N_9834);
and UO_1343 (O_1343,N_9437,N_9903);
or UO_1344 (O_1344,N_9101,N_9853);
or UO_1345 (O_1345,N_9478,N_9188);
nor UO_1346 (O_1346,N_9881,N_9640);
xnor UO_1347 (O_1347,N_9659,N_9850);
or UO_1348 (O_1348,N_9238,N_9189);
nor UO_1349 (O_1349,N_9358,N_9773);
nand UO_1350 (O_1350,N_9356,N_9483);
xor UO_1351 (O_1351,N_9022,N_9804);
and UO_1352 (O_1352,N_9226,N_9544);
nor UO_1353 (O_1353,N_9863,N_9962);
xnor UO_1354 (O_1354,N_9558,N_9930);
xnor UO_1355 (O_1355,N_9509,N_9666);
xnor UO_1356 (O_1356,N_9435,N_9755);
or UO_1357 (O_1357,N_9809,N_9924);
nand UO_1358 (O_1358,N_9247,N_9647);
nor UO_1359 (O_1359,N_9164,N_9644);
or UO_1360 (O_1360,N_9117,N_9206);
or UO_1361 (O_1361,N_9188,N_9955);
nor UO_1362 (O_1362,N_9675,N_9536);
nand UO_1363 (O_1363,N_9243,N_9803);
xor UO_1364 (O_1364,N_9803,N_9508);
xnor UO_1365 (O_1365,N_9482,N_9538);
nor UO_1366 (O_1366,N_9645,N_9104);
nor UO_1367 (O_1367,N_9596,N_9371);
nor UO_1368 (O_1368,N_9479,N_9976);
nor UO_1369 (O_1369,N_9880,N_9969);
nand UO_1370 (O_1370,N_9338,N_9253);
xor UO_1371 (O_1371,N_9816,N_9183);
or UO_1372 (O_1372,N_9125,N_9229);
nor UO_1373 (O_1373,N_9599,N_9235);
nor UO_1374 (O_1374,N_9094,N_9480);
nand UO_1375 (O_1375,N_9784,N_9260);
xor UO_1376 (O_1376,N_9074,N_9360);
xor UO_1377 (O_1377,N_9774,N_9217);
xnor UO_1378 (O_1378,N_9981,N_9898);
nand UO_1379 (O_1379,N_9861,N_9803);
nand UO_1380 (O_1380,N_9267,N_9645);
xnor UO_1381 (O_1381,N_9198,N_9960);
xnor UO_1382 (O_1382,N_9394,N_9135);
and UO_1383 (O_1383,N_9184,N_9221);
nor UO_1384 (O_1384,N_9996,N_9122);
and UO_1385 (O_1385,N_9204,N_9186);
and UO_1386 (O_1386,N_9531,N_9195);
or UO_1387 (O_1387,N_9408,N_9113);
nor UO_1388 (O_1388,N_9406,N_9778);
and UO_1389 (O_1389,N_9433,N_9578);
or UO_1390 (O_1390,N_9702,N_9300);
nor UO_1391 (O_1391,N_9740,N_9033);
nor UO_1392 (O_1392,N_9953,N_9183);
and UO_1393 (O_1393,N_9838,N_9030);
nor UO_1394 (O_1394,N_9909,N_9241);
nand UO_1395 (O_1395,N_9167,N_9968);
nor UO_1396 (O_1396,N_9217,N_9612);
nand UO_1397 (O_1397,N_9461,N_9859);
nor UO_1398 (O_1398,N_9395,N_9622);
xnor UO_1399 (O_1399,N_9768,N_9760);
and UO_1400 (O_1400,N_9157,N_9973);
nor UO_1401 (O_1401,N_9477,N_9054);
nand UO_1402 (O_1402,N_9228,N_9189);
nand UO_1403 (O_1403,N_9144,N_9413);
nand UO_1404 (O_1404,N_9018,N_9677);
or UO_1405 (O_1405,N_9191,N_9827);
and UO_1406 (O_1406,N_9764,N_9369);
nand UO_1407 (O_1407,N_9460,N_9243);
and UO_1408 (O_1408,N_9118,N_9070);
and UO_1409 (O_1409,N_9816,N_9338);
xor UO_1410 (O_1410,N_9428,N_9360);
xnor UO_1411 (O_1411,N_9758,N_9891);
xnor UO_1412 (O_1412,N_9145,N_9021);
nor UO_1413 (O_1413,N_9481,N_9194);
nor UO_1414 (O_1414,N_9424,N_9845);
and UO_1415 (O_1415,N_9558,N_9946);
nand UO_1416 (O_1416,N_9758,N_9216);
or UO_1417 (O_1417,N_9914,N_9899);
and UO_1418 (O_1418,N_9343,N_9954);
xor UO_1419 (O_1419,N_9388,N_9020);
nor UO_1420 (O_1420,N_9471,N_9741);
nor UO_1421 (O_1421,N_9686,N_9940);
or UO_1422 (O_1422,N_9341,N_9242);
and UO_1423 (O_1423,N_9917,N_9206);
or UO_1424 (O_1424,N_9249,N_9760);
nor UO_1425 (O_1425,N_9540,N_9233);
xnor UO_1426 (O_1426,N_9975,N_9415);
nand UO_1427 (O_1427,N_9115,N_9530);
nor UO_1428 (O_1428,N_9046,N_9010);
nor UO_1429 (O_1429,N_9054,N_9208);
nor UO_1430 (O_1430,N_9286,N_9133);
nor UO_1431 (O_1431,N_9594,N_9159);
nand UO_1432 (O_1432,N_9700,N_9653);
xnor UO_1433 (O_1433,N_9407,N_9609);
nor UO_1434 (O_1434,N_9871,N_9105);
or UO_1435 (O_1435,N_9655,N_9460);
nand UO_1436 (O_1436,N_9060,N_9503);
or UO_1437 (O_1437,N_9944,N_9234);
nor UO_1438 (O_1438,N_9126,N_9659);
nor UO_1439 (O_1439,N_9871,N_9860);
nor UO_1440 (O_1440,N_9402,N_9081);
nor UO_1441 (O_1441,N_9979,N_9645);
nand UO_1442 (O_1442,N_9414,N_9647);
nand UO_1443 (O_1443,N_9472,N_9266);
or UO_1444 (O_1444,N_9331,N_9990);
xnor UO_1445 (O_1445,N_9373,N_9096);
nor UO_1446 (O_1446,N_9276,N_9407);
and UO_1447 (O_1447,N_9282,N_9246);
xnor UO_1448 (O_1448,N_9386,N_9028);
or UO_1449 (O_1449,N_9682,N_9084);
nand UO_1450 (O_1450,N_9810,N_9559);
and UO_1451 (O_1451,N_9347,N_9664);
nor UO_1452 (O_1452,N_9321,N_9809);
and UO_1453 (O_1453,N_9352,N_9492);
nand UO_1454 (O_1454,N_9141,N_9094);
and UO_1455 (O_1455,N_9771,N_9197);
nand UO_1456 (O_1456,N_9793,N_9847);
and UO_1457 (O_1457,N_9666,N_9608);
and UO_1458 (O_1458,N_9382,N_9802);
nand UO_1459 (O_1459,N_9335,N_9402);
xnor UO_1460 (O_1460,N_9696,N_9098);
nand UO_1461 (O_1461,N_9045,N_9759);
or UO_1462 (O_1462,N_9281,N_9035);
or UO_1463 (O_1463,N_9029,N_9295);
or UO_1464 (O_1464,N_9711,N_9720);
and UO_1465 (O_1465,N_9285,N_9503);
xnor UO_1466 (O_1466,N_9274,N_9742);
nor UO_1467 (O_1467,N_9591,N_9372);
xor UO_1468 (O_1468,N_9363,N_9034);
xor UO_1469 (O_1469,N_9025,N_9253);
and UO_1470 (O_1470,N_9155,N_9831);
nand UO_1471 (O_1471,N_9406,N_9184);
nand UO_1472 (O_1472,N_9602,N_9743);
or UO_1473 (O_1473,N_9800,N_9596);
nand UO_1474 (O_1474,N_9797,N_9937);
xor UO_1475 (O_1475,N_9039,N_9621);
xnor UO_1476 (O_1476,N_9797,N_9136);
or UO_1477 (O_1477,N_9246,N_9242);
and UO_1478 (O_1478,N_9590,N_9356);
or UO_1479 (O_1479,N_9140,N_9328);
xor UO_1480 (O_1480,N_9760,N_9957);
or UO_1481 (O_1481,N_9673,N_9799);
xnor UO_1482 (O_1482,N_9026,N_9095);
or UO_1483 (O_1483,N_9815,N_9886);
nand UO_1484 (O_1484,N_9427,N_9144);
xnor UO_1485 (O_1485,N_9830,N_9793);
xnor UO_1486 (O_1486,N_9173,N_9386);
nor UO_1487 (O_1487,N_9074,N_9458);
nand UO_1488 (O_1488,N_9849,N_9099);
nor UO_1489 (O_1489,N_9334,N_9399);
xnor UO_1490 (O_1490,N_9802,N_9463);
nor UO_1491 (O_1491,N_9660,N_9859);
nand UO_1492 (O_1492,N_9677,N_9523);
nand UO_1493 (O_1493,N_9351,N_9114);
nor UO_1494 (O_1494,N_9373,N_9569);
nor UO_1495 (O_1495,N_9668,N_9754);
nor UO_1496 (O_1496,N_9322,N_9493);
and UO_1497 (O_1497,N_9176,N_9715);
xor UO_1498 (O_1498,N_9092,N_9347);
or UO_1499 (O_1499,N_9895,N_9943);
endmodule